magic
tech sky130B
magscale 1 2
timestamp 1696637874
<< error_p >>
rect -29 1058 29 1064
rect -29 1024 -17 1058
rect -29 1018 29 1024
rect -29 693 29 699
rect -29 659 -17 693
rect -29 653 29 659
rect -29 70 29 76
rect -29 36 -17 70
rect -29 30 29 36
rect -33 20 33 21
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -402 29 -396
rect -29 -436 -17 -402
rect -29 -442 29 -436
rect -29 -767 29 -761
rect -29 -801 -17 -767
rect -29 -807 29 -801
<< nwell >>
rect -226 -1196 226 1196
<< pmos >>
rect -30 777 30 977
rect -30 412 30 612
rect -30 117 30 317
rect -30 -318 30 -118
rect -30 -683 30 -483
rect -30 -1048 30 -848
<< pdiff >>
rect -88 947 -30 977
rect -88 807 -76 947
rect -42 807 -30 947
rect -88 777 -30 807
rect 30 947 88 977
rect 30 807 42 947
rect 76 807 88 947
rect 30 777 88 807
rect -88 582 -30 612
rect -88 442 -76 582
rect -42 442 -30 582
rect -88 412 -30 442
rect 30 582 88 612
rect 30 442 42 582
rect 76 442 88 582
rect 30 412 88 442
rect -88 287 -30 317
rect -88 147 -76 287
rect -42 147 -30 287
rect -88 117 -30 147
rect 30 287 88 317
rect 30 147 42 287
rect 76 147 88 287
rect 30 117 88 147
rect -88 -148 -30 -118
rect -88 -288 -76 -148
rect -42 -288 -30 -148
rect -88 -318 -30 -288
rect 30 -148 88 -118
rect 30 -288 42 -148
rect 76 -288 88 -148
rect 30 -318 88 -288
rect -88 -513 -30 -483
rect -88 -653 -76 -513
rect -42 -653 -30 -513
rect -88 -683 -30 -653
rect 30 -513 88 -483
rect 30 -653 42 -513
rect 76 -653 88 -513
rect 30 -683 88 -653
rect -88 -878 -30 -848
rect -88 -1018 -76 -878
rect -42 -1018 -30 -878
rect -88 -1048 -30 -1018
rect 30 -878 88 -848
rect 30 -1018 42 -878
rect 76 -1018 88 -878
rect 30 -1048 88 -1018
<< pdiffc >>
rect -76 807 -42 947
rect 42 807 76 947
rect -76 442 -42 582
rect 42 442 76 582
rect -76 147 -42 287
rect 42 147 76 287
rect -76 -288 -42 -148
rect 42 -288 76 -148
rect -76 -653 -42 -513
rect 42 -653 76 -513
rect -76 -1018 -42 -878
rect 42 -1018 76 -878
<< nsubdiff >>
rect -190 1126 -75 1160
rect 75 1126 190 1160
rect -190 -1126 -156 1126
rect 156 -1126 190 1126
rect -190 -1160 -75 -1126
rect 75 -1160 190 -1126
<< nsubdiffcont >>
rect -75 1126 75 1160
rect -75 -1160 75 -1126
<< poly >>
rect -33 1058 33 1074
rect -33 1024 -17 1058
rect 17 1024 33 1058
rect -33 1008 33 1024
rect -30 977 30 1008
rect -30 751 30 777
rect -33 693 33 709
rect -33 659 -17 693
rect 17 659 33 693
rect -33 643 33 659
rect -30 612 30 643
rect -30 386 30 412
rect -30 317 30 343
rect -30 86 30 117
rect -33 70 33 86
rect -33 36 -17 70
rect 17 36 33 70
rect -33 20 33 36
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -30 -118 30 -87
rect -30 -344 30 -318
rect -33 -402 33 -386
rect -33 -436 -17 -402
rect 17 -436 33 -402
rect -33 -452 33 -436
rect -30 -483 30 -452
rect -30 -709 30 -683
rect -33 -767 33 -751
rect -33 -801 -17 -767
rect 17 -801 33 -767
rect -33 -817 33 -801
rect -30 -848 30 -817
rect -30 -1074 30 -1048
<< polycont >>
rect -17 1024 17 1058
rect -17 659 17 693
rect -17 36 17 70
rect -17 -71 17 -37
rect -17 -436 17 -402
rect -17 -801 17 -767
<< locali >>
rect -91 1126 -75 1160
rect 75 1126 91 1160
rect -33 1024 -17 1058
rect 17 1024 33 1058
rect -76 947 -42 963
rect -76 791 -42 807
rect 42 947 76 963
rect 42 791 76 807
rect -33 659 -17 693
rect 17 659 33 693
rect -76 582 -42 598
rect -76 426 -42 442
rect 42 582 76 598
rect 42 426 76 442
rect -76 287 -42 303
rect -76 131 -42 147
rect 42 287 76 303
rect 42 131 76 147
rect -33 36 -17 70
rect 17 36 33 70
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -76 -148 -42 -132
rect -76 -304 -42 -288
rect 42 -148 76 -132
rect 42 -304 76 -288
rect -33 -436 -17 -402
rect 17 -436 33 -402
rect -76 -513 -42 -497
rect -76 -669 -42 -653
rect 42 -513 76 -497
rect 42 -669 76 -653
rect -33 -801 -17 -767
rect 17 -801 33 -767
rect -76 -878 -42 -862
rect -76 -1034 -42 -1018
rect 42 -878 76 -862
rect 42 -1034 76 -1018
rect -91 -1160 -75 -1126
rect 75 -1160 91 -1126
<< viali >>
rect -17 1024 17 1058
rect -76 807 -42 947
rect 42 824 76 930
rect -17 659 17 693
rect -76 442 -42 582
rect 42 459 76 565
rect -76 147 -42 287
rect 42 164 76 270
rect -17 36 17 70
rect -17 -71 17 -37
rect -76 -288 -42 -148
rect 42 -271 76 -165
rect -17 -436 17 -402
rect -76 -653 -42 -513
rect 42 -636 76 -530
rect -17 -801 17 -767
rect -76 -1018 -42 -878
rect 42 -1001 76 -895
<< metal1 >>
rect -29 1058 29 1064
rect -29 1024 -17 1058
rect 17 1024 29 1058
rect -29 1018 29 1024
rect -82 947 -36 959
rect -82 807 -76 947
rect -42 807 -36 947
rect 36 930 82 942
rect 36 824 42 930
rect 76 824 82 930
rect 36 812 82 824
rect -82 795 -36 807
rect -29 693 29 699
rect -29 659 -17 693
rect 17 659 29 693
rect -29 653 29 659
rect -82 582 -36 594
rect -82 442 -76 582
rect -42 442 -36 582
rect 36 565 82 577
rect 36 459 42 565
rect 76 459 82 565
rect 36 447 82 459
rect -82 430 -36 442
rect -82 287 -36 299
rect -82 147 -76 287
rect -42 147 -36 287
rect 36 270 82 282
rect 36 164 42 270
rect 76 164 82 270
rect 36 152 82 164
rect -82 135 -36 147
rect -29 70 29 76
rect -29 36 -17 70
rect 17 36 29 70
rect -29 30 29 36
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -82 -148 -36 -136
rect -82 -288 -76 -148
rect -42 -288 -36 -148
rect 36 -165 82 -153
rect 36 -271 42 -165
rect 76 -271 82 -165
rect 36 -283 82 -271
rect -82 -300 -36 -288
rect -29 -402 29 -396
rect -29 -436 -17 -402
rect 17 -436 29 -402
rect -29 -442 29 -436
rect -82 -513 -36 -501
rect -82 -653 -76 -513
rect -42 -653 -36 -513
rect 36 -530 82 -518
rect 36 -636 42 -530
rect 76 -636 82 -530
rect 36 -648 82 -636
rect -82 -665 -36 -653
rect -29 -767 29 -761
rect -29 -801 -17 -767
rect 17 -801 29 -767
rect -29 -807 29 -801
rect -82 -878 -36 -866
rect -82 -1018 -76 -878
rect -42 -1018 -36 -878
rect 36 -895 82 -883
rect 36 -1001 42 -895
rect 76 -1001 82 -895
rect 36 -1013 82 -1001
rect -82 -1030 -36 -1018
<< properties >>
string FIXED_BBOX -173 -1143 173 1143
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.3 m 6 nf 1 diffcov 80 polycov 80 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 80 rlcov 80 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 60 viadrn 80 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
