* NGSPICE file created from dac.ext - technology: sky130B

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_FJK8MD m3_n386_n240# c1_n346_n200#
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt unitcap cp cn
Xsky130_fd_pr__cap_mim_m3_1_FJK8MD_0 cn cp sky130_fd_pr__cap_mim_m3_1_FJK8MD
.ends

.subckt carray n7 n6 n5 ndum n4 n3 n1 n0 unitcap_9/cp n2
Xunitcap_190 unitcap_9/cp n5 unitcap
Xunitcap_191 unitcap_9/cp unitcap_191/cn unitcap
Xunitcap_180 unitcap_9/cp n6 unitcap
Xunitcap_181 unitcap_9/cp n6 unitcap
Xunitcap_170 unitcap_9/cp n6 unitcap
Xunitcap_192 unitcap_9/cp unitcap_192/cn unitcap
Xunitcap_330 unitcap_9/cp unitcap_330/cn unitcap
Xunitcap_182 unitcap_9/cp n6 unitcap
Xunitcap_171 unitcap_9/cp n6 unitcap
Xunitcap_160 unitcap_9/cp unitcap_160/cn unitcap
Xunitcap_193 unitcap_9/cp n6 unitcap
Xunitcap_183 unitcap_9/cp unitcap_183/cn unitcap
Xunitcap_150 unitcap_9/cp n6 unitcap
Xunitcap_331 unitcap_9/cp unitcap_331/cn unitcap
Xunitcap_172 unitcap_9/cp n6 unitcap
Xunitcap_194 unitcap_9/cp n6 unitcap
Xunitcap_161 unitcap_9/cp n6 unitcap
Xunitcap_320 unitcap_9/cp unitcap_320/cn unitcap
Xunitcap_332 unitcap_9/cp n2 unitcap
Xunitcap_310 unitcap_9/cp n6 unitcap
Xunitcap_321 unitcap_9/cp unitcap_321/cn unitcap
Xunitcap_151 unitcap_9/cp unitcap_151/cn unitcap
Xunitcap_173 unitcap_9/cp n6 unitcap
Xunitcap_140 unitcap_9/cp n7 unitcap
Xunitcap_195 unitcap_9/cp n6 unitcap
Xunitcap_162 unitcap_9/cp n6 unitcap
Xunitcap_184 unitcap_9/cp unitcap_184/cn unitcap
Xunitcap_174 unitcap_9/cp n6 unitcap
Xunitcap_141 unitcap_9/cp n7 unitcap
Xunitcap_333 unitcap_9/cp n2 unitcap
Xunitcap_196 unitcap_9/cp n6 unitcap
Xunitcap_163 unitcap_9/cp n6 unitcap
Xunitcap_130 unitcap_9/cp n6 unitcap
Xunitcap_311 unitcap_9/cp n6 unitcap
Xunitcap_300 unitcap_9/cp n7 unitcap
Xunitcap_322 unitcap_9/cp unitcap_322/cn unitcap
Xunitcap_152 unitcap_9/cp unitcap_152/cn unitcap
Xunitcap_185 unitcap_9/cp n5 unitcap
Xunitcap_334 unitcap_9/cp unitcap_334/cn unitcap
Xunitcap_312 unitcap_9/cp n5 unitcap
Xunitcap_301 unitcap_9/cp n7 unitcap
Xunitcap_323 unitcap_9/cp n0 unitcap
Xunitcap_175 unitcap_9/cp unitcap_175/cn unitcap
Xunitcap_142 unitcap_9/cp n7 unitcap
Xunitcap_197 unitcap_9/cp n6 unitcap
Xunitcap_164 unitcap_9/cp n6 unitcap
Xunitcap_131 unitcap_9/cp n6 unitcap
Xunitcap_186 unitcap_9/cp n5 unitcap
Xunitcap_120 unitcap_9/cp unitcap_120/cn unitcap
Xunitcap_153 unitcap_9/cp n6 unitcap
Xunitcap_90 unitcap_9/cp n7 unitcap
Xunitcap_198 unitcap_9/cp n6 unitcap
Xunitcap_143 unitcap_9/cp unitcap_143/cn unitcap
Xunitcap_110 unitcap_9/cp n7 unitcap
Xunitcap_165 unitcap_9/cp n6 unitcap
Xunitcap_132 unitcap_9/cp n6 unitcap
Xunitcap_335 unitcap_9/cp n2 unitcap
Xunitcap_187 unitcap_9/cp n5 unitcap
Xunitcap_154 unitcap_9/cp n6 unitcap
Xunitcap_313 unitcap_9/cp n6 unitcap
Xunitcap_302 unitcap_9/cp n7 unitcap
Xunitcap_121 unitcap_9/cp n7 unitcap
Xunitcap_176 unitcap_9/cp unitcap_176/cn unitcap
Xunitcap_324 unitcap_9/cp unitcap_324/cn unitcap
Xunitcap_336 unitcap_9/cp unitcap_336/cn unitcap
Xunitcap_91 unitcap_9/cp n7 unitcap
Xunitcap_314 unitcap_9/cp n5 unitcap
Xunitcap_303 unitcap_9/cp n7 unitcap
Xunitcap_80 unitcap_9/cp unitcap_80/cn unitcap
Xunitcap_325 unitcap_9/cp ndum unitcap
Xunitcap_199 unitcap_9/cp unitcap_199/cn unitcap
Xunitcap_166 unitcap_9/cp n6 unitcap
Xunitcap_111 unitcap_9/cp unitcap_111/cn unitcap
Xunitcap_133 unitcap_9/cp n6 unitcap
Xunitcap_188 unitcap_9/cp n5 unitcap
Xunitcap_100 unitcap_9/cp n7 unitcap
Xunitcap_155 unitcap_9/cp n6 unitcap
Xunitcap_122 unitcap_9/cp n7 unitcap
Xunitcap_144 unitcap_9/cp unitcap_144/cn unitcap
Xunitcap_177 unitcap_9/cp n6 unitcap
Xunitcap_70 unitcap_9/cp n7 unitcap
Xunitcap_337 unitcap_9/cp unitcap_337/cn unitcap
Xunitcap_101 unitcap_9/cp n7 unitcap
Xunitcap_92 unitcap_9/cp n7 unitcap
Xunitcap_326 unitcap_9/cp unitcap_326/cn unitcap
Xunitcap_315 unitcap_9/cp n5 unitcap
Xunitcap_304 unitcap_9/cp n7 unitcap
Xunitcap_81 unitcap_9/cp n7 unitcap
Xunitcap_112 unitcap_9/cp unitcap_112/cn unitcap
Xunitcap_167 unitcap_9/cp unitcap_167/cn unitcap
Xunitcap_134 unitcap_9/cp n6 unitcap
Xunitcap_189 unitcap_9/cp n5 unitcap
Xunitcap_156 unitcap_9/cp n6 unitcap
Xunitcap_123 unitcap_9/cp n7 unitcap
Xunitcap_178 unitcap_9/cp n6 unitcap
Xunitcap_145 unitcap_9/cp n6 unitcap
Xunitcap_338 unitcap_9/cp unitcap_338/cn unitcap
Xunitcap_71 unitcap_9/cp unitcap_71/cn unitcap
Xunitcap_93 unitcap_9/cp n7 unitcap
Xunitcap_60 unitcap_9/cp n7 unitcap
Xunitcap_327 unitcap_9/cp n1 unitcap
Xunitcap_82 unitcap_9/cp n7 unitcap
Xunitcap_316 unitcap_9/cp n5 unitcap
Xunitcap_305 unitcap_9/cp n6 unitcap
Xunitcap_135 unitcap_9/cp unitcap_135/cn unitcap
Xunitcap_102 unitcap_9/cp n7 unitcap
Xunitcap_157 unitcap_9/cp n6 unitcap
Xunitcap_124 unitcap_9/cp n7 unitcap
Xunitcap_179 unitcap_9/cp n6 unitcap
Xunitcap_146 unitcap_9/cp n6 unitcap
Xunitcap_113 unitcap_9/cp n7 unitcap
Xunitcap_168 unitcap_9/cp unitcap_168/cn unitcap
Xunitcap_339 unitcap_9/cp n2 unitcap
Xunitcap_94 unitcap_9/cp n7 unitcap
Xunitcap_61 unitcap_9/cp n7 unitcap
Xunitcap_83 unitcap_9/cp n7 unitcap
Xunitcap_50 unitcap_9/cp n7 unitcap
Xunitcap_328 unitcap_9/cp unitcap_328/cn unitcap
Xunitcap_317 unitcap_9/cp n4 unitcap
Xunitcap_306 unitcap_9/cp n6 unitcap
Xunitcap_72 unitcap_9/cp unitcap_72/cn unitcap
Xunitcap_158 unitcap_9/cp n6 unitcap
Xunitcap_103 unitcap_9/cp unitcap_103/cn unitcap
Xunitcap_125 unitcap_9/cp n7 unitcap
Xunitcap_147 unitcap_9/cp n6 unitcap
Xunitcap_114 unitcap_9/cp n7 unitcap
Xunitcap_136 unitcap_9/cp unitcap_136/cn unitcap
Xunitcap_169 unitcap_9/cp n6 unitcap
Xunitcap_95 unitcap_9/cp unitcap_95/cn unitcap
Xunitcap_62 unitcap_9/cp n7 unitcap
Xunitcap_84 unitcap_9/cp n7 unitcap
Xunitcap_51 unitcap_9/cp n7 unitcap
Xunitcap_329 unitcap_9/cp n1 unitcap
Xunitcap_318 unitcap_9/cp n4 unitcap
Xunitcap_307 unitcap_9/cp n6 unitcap
Xunitcap_40 unitcap_9/cp unitcap_40/cn unitcap
Xunitcap_73 unitcap_9/cp n7 unitcap
Xunitcap_159 unitcap_9/cp unitcap_159/cn unitcap
Xunitcap_126 unitcap_9/cp n7 unitcap
Xunitcap_148 unitcap_9/cp n6 unitcap
Xunitcap_115 unitcap_9/cp n7 unitcap
Xunitcap_104 unitcap_9/cp unitcap_104/cn unitcap
Xunitcap_137 unitcap_9/cp n7 unitcap
Xunitcap_63 unitcap_9/cp unitcap_63/cn unitcap
Xunitcap_30 unitcap_9/cp n7 unitcap
Xunitcap_85 unitcap_9/cp n7 unitcap
Xunitcap_52 unitcap_9/cp n7 unitcap
Xunitcap_74 unitcap_9/cp n7 unitcap
Xunitcap_319 unitcap_9/cp n3 unitcap
Xunitcap_308 unitcap_9/cp n6 unitcap
Xunitcap_41 unitcap_9/cp n7 unitcap
Xunitcap_96 unitcap_9/cp unitcap_96/cn unitcap
Xunitcap_127 unitcap_9/cp unitcap_127/cn unitcap
Xunitcap_149 unitcap_9/cp n6 unitcap
Xunitcap_116 unitcap_9/cp n7 unitcap
Xunitcap_138 unitcap_9/cp n7 unitcap
Xunitcap_105 unitcap_9/cp n7 unitcap
Xunitcap_86 unitcap_9/cp n7 unitcap
Xunitcap_31 unitcap_9/cp unitcap_31/cn unitcap
Xunitcap_53 unitcap_9/cp n7 unitcap
Xunitcap_20 unitcap_9/cp n7 unitcap
Xunitcap_75 unitcap_9/cp n7 unitcap
Xunitcap_42 unitcap_9/cp n7 unitcap
Xunitcap_64 unitcap_9/cp unitcap_64/cn unitcap
Xunitcap_97 unitcap_9/cp n7 unitcap
Xunitcap_117 unitcap_9/cp n7 unitcap
Xunitcap_139 unitcap_9/cp n7 unitcap
Xunitcap_106 unitcap_9/cp n7 unitcap
Xunitcap_309 unitcap_9/cp n6 unitcap
Xunitcap_128 unitcap_9/cp unitcap_128/cn unitcap
Xunitcap_87 unitcap_9/cp unitcap_87/cn unitcap
Xunitcap_54 unitcap_9/cp n7 unitcap
Xunitcap_21 unitcap_9/cp n7 unitcap
Xunitcap_76 unitcap_9/cp n7 unitcap
Xunitcap_43 unitcap_9/cp n7 unitcap
Xunitcap_98 unitcap_9/cp n7 unitcap
Xunitcap_10 unitcap_9/cp unitcap_10/cn unitcap
Xunitcap_32 unitcap_9/cp unitcap_32/cn unitcap
Xunitcap_65 unitcap_9/cp n7 unitcap
Xunitcap_118 unitcap_9/cp n7 unitcap
Xunitcap_107 unitcap_9/cp n7 unitcap
Xunitcap_129 unitcap_9/cp n6 unitcap
Xunitcap_290 unitcap_9/cp n7 unitcap
Xunitcap_55 unitcap_9/cp unitcap_55/cn unitcap
Xunitcap_22 unitcap_9/cp n7 unitcap
Xunitcap_77 unitcap_9/cp n7 unitcap
Xunitcap_44 unitcap_9/cp n7 unitcap
Xunitcap_99 unitcap_9/cp n7 unitcap
Xunitcap_11 unitcap_9/cp unitcap_11/cn unitcap
Xunitcap_66 unitcap_9/cp n7 unitcap
Xunitcap_0 unitcap_9/cp unitcap_0/cn unitcap
Xunitcap_33 unitcap_9/cp n7 unitcap
Xunitcap_88 unitcap_9/cp unitcap_88/cn unitcap
Xunitcap_119 unitcap_9/cp unitcap_119/cn unitcap
Xunitcap_108 unitcap_9/cp n7 unitcap
Xunitcap_291 unitcap_9/cp n7 unitcap
Xunitcap_1 unitcap_9/cp n7 unitcap
Xunitcap_280 unitcap_9/cp n5 unitcap
Xunitcap_78 unitcap_9/cp n7 unitcap
Xunitcap_23 unitcap_9/cp unitcap_23/cn unitcap
Xunitcap_45 unitcap_9/cp n7 unitcap
Xunitcap_12 unitcap_9/cp unitcap_12/cn unitcap
Xunitcap_67 unitcap_9/cp n7 unitcap
Xunitcap_34 unitcap_9/cp n7 unitcap
Xunitcap_56 unitcap_9/cp unitcap_56/cn unitcap
Xunitcap_89 unitcap_9/cp n7 unitcap
Xunitcap_109 unitcap_9/cp n7 unitcap
Xunitcap_292 unitcap_9/cp n7 unitcap
Xunitcap_270 unitcap_9/cp n7 unitcap
Xunitcap_281 unitcap_9/cp n6 unitcap
Xunitcap_79 unitcap_9/cp unitcap_79/cn unitcap
Xunitcap_46 unitcap_9/cp n7 unitcap
Xunitcap_68 unitcap_9/cp n7 unitcap
Xunitcap_13 unitcap_9/cp unitcap_13/cn unitcap
Xunitcap_35 unitcap_9/cp n7 unitcap
Xunitcap_2 unitcap_9/cp n7 unitcap
Xunitcap_24 unitcap_9/cp unitcap_24/cn unitcap
Xunitcap_57 unitcap_9/cp n7 unitcap
Xunitcap_3 unitcap_9/cp n7 unitcap
Xunitcap_293 unitcap_9/cp n7 unitcap
Xunitcap_260 unitcap_9/cp n7 unitcap
Xunitcap_271 unitcap_9/cp n7 unitcap
Xunitcap_282 unitcap_9/cp n5 unitcap
Xunitcap_47 unitcap_9/cp unitcap_47/cn unitcap
Xunitcap_14 unitcap_9/cp unitcap_14/cn unitcap
Xunitcap_69 unitcap_9/cp n7 unitcap
Xunitcap_36 unitcap_9/cp n7 unitcap
Xunitcap_58 unitcap_9/cp n7 unitcap
Xunitcap_25 unitcap_9/cp n7 unitcap
Xunitcap_4 unitcap_9/cp n7 unitcap
Xunitcap_250 unitcap_9/cp n3 unitcap
Xunitcap_294 unitcap_9/cp n7 unitcap
Xunitcap_283 unitcap_9/cp n5 unitcap
Xunitcap_261 unitcap_9/cp n7 unitcap
Xunitcap_272 unitcap_9/cp n7 unitcap
Xunitcap_15 unitcap_9/cp unitcap_15/cn unitcap
Xunitcap_37 unitcap_9/cp n7 unitcap
Xunitcap_59 unitcap_9/cp n7 unitcap
Xunitcap_26 unitcap_9/cp n7 unitcap
Xunitcap_48 unitcap_9/cp unitcap_48/cn unitcap
Xunitcap_5 unitcap_9/cp n7 unitcap
Xunitcap_251 unitcap_9/cp n3 unitcap
Xunitcap_295 unitcap_9/cp n7 unitcap
Xunitcap_240 unitcap_9/cp unitcap_240/cn unitcap
Xunitcap_262 unitcap_9/cp n7 unitcap
Xunitcap_273 unitcap_9/cp n6 unitcap
Xunitcap_284 unitcap_9/cp n5 unitcap
Xunitcap_38 unitcap_9/cp n7 unitcap
Xunitcap_27 unitcap_9/cp n7 unitcap
Xunitcap_16 unitcap_9/cp unitcap_16/cn unitcap
Xunitcap_49 unitcap_9/cp n7 unitcap
Xunitcap_230 unitcap_9/cp n5 unitcap
Xunitcap_6 unitcap_9/cp n7 unitcap
Xunitcap_252 unitcap_9/cp n3 unitcap
Xunitcap_296 unitcap_9/cp n7 unitcap
Xunitcap_285 unitcap_9/cp n4 unitcap
Xunitcap_241 unitcap_9/cp n4 unitcap
Xunitcap_263 unitcap_9/cp n7 unitcap
Xunitcap_274 unitcap_9/cp n6 unitcap
Xunitcap_39 unitcap_9/cp unitcap_39/cn unitcap
Xunitcap_28 unitcap_9/cp n7 unitcap
Xunitcap_17 unitcap_9/cp n7 unitcap
Xunitcap_231 unitcap_9/cp unitcap_231/cn unitcap
Xunitcap_7 unitcap_9/cp unitcap_7/cn unitcap
Xunitcap_253 unitcap_9/cp n3 unitcap
Xunitcap_220 unitcap_9/cp n5 unitcap
Xunitcap_242 unitcap_9/cp n4 unitcap
Xunitcap_297 unitcap_9/cp n7 unitcap
Xunitcap_286 unitcap_9/cp n4 unitcap
Xunitcap_264 unitcap_9/cp n7 unitcap
Xunitcap_275 unitcap_9/cp n6 unitcap
Xunitcap_29 unitcap_9/cp n7 unitcap
Xunitcap_18 unitcap_9/cp n7 unitcap
Xunitcap_254 unitcap_9/cp n3 unitcap
Xunitcap_221 unitcap_9/cp n5 unitcap
Xunitcap_243 unitcap_9/cp n4 unitcap
Xunitcap_210 unitcap_9/cp n5 unitcap
Xunitcap_298 unitcap_9/cp n7 unitcap
Xunitcap_287 unitcap_9/cp n3 unitcap
Xunitcap_8 unitcap_9/cp unitcap_8/cn unitcap
Xunitcap_232 unitcap_9/cp unitcap_232/cn unitcap
Xunitcap_265 unitcap_9/cp n7 unitcap
Xunitcap_276 unitcap_9/cp n6 unitcap
Xunitcap_19 unitcap_9/cp n7 unitcap
Xunitcap_255 unitcap_9/cp unitcap_255/cn unitcap
Xunitcap_222 unitcap_9/cp n5 unitcap
Xunitcap_244 unitcap_9/cp n4 unitcap
Xunitcap_211 unitcap_9/cp n5 unitcap
Xunitcap_299 unitcap_9/cp n7 unitcap
Xunitcap_288 unitcap_9/cp unitcap_288/cn unitcap
Xunitcap_9 unitcap_9/cp unitcap_9/cn unitcap
Xunitcap_200 unitcap_9/cp unitcap_200/cn unitcap
Xunitcap_233 unitcap_9/cp n4 unitcap
Xunitcap_266 unitcap_9/cp n7 unitcap
Xunitcap_277 unitcap_9/cp n6 unitcap
Xunitcap_223 unitcap_9/cp unitcap_223/cn unitcap
Xunitcap_245 unitcap_9/cp n4 unitcap
Xunitcap_212 unitcap_9/cp n5 unitcap
Xunitcap_234 unitcap_9/cp n4 unitcap
Xunitcap_289 unitcap_9/cp n7 unitcap
Xunitcap_201 unitcap_9/cp n6 unitcap
Xunitcap_256 unitcap_9/cp unitcap_256/cn unitcap
Xunitcap_267 unitcap_9/cp n7 unitcap
Xunitcap_278 unitcap_9/cp n6 unitcap
Xunitcap_246 unitcap_9/cp n4 unitcap
Xunitcap_213 unitcap_9/cp n5 unitcap
Xunitcap_235 unitcap_9/cp n4 unitcap
Xunitcap_202 unitcap_9/cp n6 unitcap
Xunitcap_224 unitcap_9/cp unitcap_224/cn unitcap
Xunitcap_257 unitcap_9/cp n7 unitcap
Xunitcap_268 unitcap_9/cp n7 unitcap
Xunitcap_279 unitcap_9/cp n6 unitcap
Xunitcap_247 unitcap_9/cp unitcap_247/cn unitcap
Xunitcap_214 unitcap_9/cp n5 unitcap
Xunitcap_236 unitcap_9/cp n4 unitcap
Xunitcap_203 unitcap_9/cp n6 unitcap
Xunitcap_225 unitcap_9/cp n5 unitcap
Xunitcap_258 unitcap_9/cp n7 unitcap
Xunitcap_269 unitcap_9/cp n7 unitcap
Xunitcap_215 unitcap_9/cp unitcap_215/cn unitcap
Xunitcap_237 unitcap_9/cp n4 unitcap
Xunitcap_204 unitcap_9/cp n6 unitcap
Xunitcap_226 unitcap_9/cp n5 unitcap
Xunitcap_248 unitcap_9/cp unitcap_248/cn unitcap
Xunitcap_259 unitcap_9/cp n7 unitcap
Xunitcap_238 unitcap_9/cp n4 unitcap
Xunitcap_205 unitcap_9/cp n6 unitcap
Xunitcap_227 unitcap_9/cp n5 unitcap
Xunitcap_216 unitcap_9/cp unitcap_216/cn unitcap
Xunitcap_249 unitcap_9/cp n3 unitcap
Xunitcap_239 unitcap_9/cp unitcap_239/cn unitcap
Xunitcap_206 unitcap_9/cp n6 unitcap
Xunitcap_228 unitcap_9/cp n5 unitcap
Xunitcap_217 unitcap_9/cp n5 unitcap
Xunitcap_207 unitcap_9/cp unitcap_207/cn unitcap
Xunitcap_229 unitcap_9/cp n5 unitcap
Xunitcap_218 unitcap_9/cp n5 unitcap
Xunitcap_219 unitcap_9/cp n5 unitcap
Xunitcap_208 unitcap_9/cp unitcap_208/cn unitcap
Xunitcap_209 unitcap_9/cp n5 unitcap
.ends

.subckt sky130_fd_pr__pfet_01v8_VVAZD4 a_89_n136# a_n501_n136# a_26_95# a_561_n136#
+ a_n383_n136# a_n328_95# a_n446_95# w_n757_n284# a_443_n136# a_n265_n136# a_n210_95#
+ a_n619_n136# G0 a_325_n136# a_n147_n136# a_498_95# a_144_95# a_207_n136# a_262_95#
+ a_n29_n136# a_380_95# a_n92_95#
X0 a_443_n136# a_380_95# a_325_n136# w_n757_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 a_n383_n136# a_n446_95# a_n501_n136# w_n757_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 a_n29_n136# a_n92_95# a_n147_n136# w_n757_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 a_325_n136# a_262_95# a_207_n136# w_n757_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X4 a_561_n136# a_498_95# a_443_n136# w_n757_n284# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X5 a_n265_n136# a_n328_95# a_n383_n136# w_n757_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 a_89_n136# a_26_95# a_n29_n136# w_n757_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_207_n136# a_144_95# a_89_n136# w_n757_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X8 a_n501_n136# G0 a_n619_n136# w_n757_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X9 a_n147_n136# a_n210_95# a_n265_n136# w_n757_n284# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_pr__nfet_01v8_JJRV6Y a_n501_n131# a_561_n131# a_26_91# a_n383_n131#
+ a_n328_91# a_n446_91# a_n564_91# a_443_n131# a_n265_n131# a_n619_n131# a_n210_91#
+ a_n721_n243# a_325_n131# a_n147_n131# a_498_91# a_207_n131# a_144_91# a_262_91#
+ a_n29_n131# a_380_91# a_n92_91# a_89_n131#
X0 a_561_n131# a_498_91# a_443_n131# a_n721_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X1 a_n265_n131# a_n328_91# a_n383_n131# a_n721_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 a_89_n131# a_26_91# a_n29_n131# a_n721_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 a_207_n131# a_144_91# a_89_n131# a_n721_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X4 a_n501_n131# a_n564_91# a_n619_n131# a_n721_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X5 a_n147_n131# a_n210_91# a_n265_n131# a_n721_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 a_443_n131# a_380_91# a_325_n131# a_n721_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_n383_n131# a_n446_91# a_n501_n131# a_n721_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X8 a_n29_n131# a_n92_91# a_n147_n131# a_n721_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X9 a_325_n131# a_262_91# a_207_n131# a_n721_n243# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt sw_top out en in vdd vss
Xsky130_fd_pr__pfet_01v8_VVAZD4_0 in out en_buf in in en_buf en_buf vdd out out en_buf
+ in en_buf in in en_buf en_buf out en_buf out en_buf en_buf sky130_fd_pr__pfet_01v8_VVAZD4
Xsky130_fd_sc_hd__decap_3_0 vss vss vdd vdd sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__inv_4_0 en_buf vss vss vdd vdd net1 sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__inv_4_1 en vss vss vdd vdd en_buf sky130_fd_sc_hd__inv_4
Xsky130_fd_sc_hd__decap_8_0 vss vss vdd vdd sky130_fd_sc_hd__decap_8
Xsky130_fd_pr__nfet_01v8_JJRV6Y_0 out in net1 in net1 net1 net1 out out in net1 vss
+ in in net1 out net1 net1 out net1 net1 in sky130_fd_pr__nfet_01v8_JJRV6Y
.ends

.subckt dac ctl0 ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 dum vin vdd sample out vss
Xsky130_fd_sc_hd__inv_2_0 ctl5 vss vss sky130_fd_sc_hd__tap_2_1/VPB vdd carray_0/n5
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_1 ctl6 vss vss sky130_fd_sc_hd__tap_2_1/VPB vdd carray_0/n6
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_2 ctl7 vss vss sky130_fd_sc_hd__tap_2_1/VPB vdd carray_0/n7
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_3 ctl3 vss vss sky130_fd_sc_hd__tap_2_1/VPB vdd carray_0/n3
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_4 ctl1 vss vss sky130_fd_sc_hd__tap_2_1/VPB vdd carray_0/n1
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_6 ctl0 vss vss sky130_fd_sc_hd__tap_2_1/VPB vdd carray_0/n0
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_5 ctl2 vss vss sky130_fd_sc_hd__tap_2_1/VPB vdd carray_0/n2
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_7 dum vss vss sky130_fd_sc_hd__tap_2_1/VPB vdd carray_0/ndum
+ sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_8 ctl4 vss vss sky130_fd_sc_hd__tap_2_1/VPB vdd carray_0/n4
+ sky130_fd_sc_hd__inv_2
Xcarray_0 carray_0/n7 carray_0/n6 carray_0/n5 carray_0/ndum carray_0/n4 carray_0/n3
+ carray_0/n1 carray_0/n0 out carray_0/n2 carray
Xsw_top_0 out sample vin vdd vss sw_top
Xsw_top_1 out sample vin vdd vss sw_top
Xsw_top_2 out sample vin vdd vss sw_top
Xsw_top_3 out sample vin vdd vss sw_top
.ends

