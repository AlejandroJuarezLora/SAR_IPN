magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 406 542
<< pwell >>
rect 1 -19 367 163
rect 30 -57 64 -19
<< scnmos >>
rect 79 7 109 137
rect 175 7 205 137
rect 259 7 289 137
<< scpmoshvt >>
rect 79 257 109 457
rect 151 257 181 457
rect 259 317 289 457
<< ndiff >>
rect 27 63 79 137
rect 27 29 35 63
rect 69 29 79 63
rect 27 7 79 29
rect 109 49 175 137
rect 109 15 131 49
rect 165 15 175 49
rect 109 7 175 15
rect 205 72 259 137
rect 205 38 215 72
rect 249 38 259 72
rect 205 7 259 38
rect 289 88 341 137
rect 289 54 299 88
rect 333 54 341 88
rect 289 7 341 54
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 377 79 411
rect 27 343 35 377
rect 69 343 79 377
rect 27 309 79 343
rect 27 275 35 309
rect 69 275 79 309
rect 27 257 79 275
rect 109 257 151 457
rect 181 445 259 457
rect 181 411 209 445
rect 243 411 259 445
rect 181 377 259 411
rect 181 343 209 377
rect 243 343 259 377
rect 181 317 259 343
rect 289 445 341 457
rect 289 411 299 445
rect 333 411 341 445
rect 289 377 341 411
rect 289 343 299 377
rect 333 343 341 377
rect 289 317 341 343
rect 181 257 231 317
<< ndiffc >>
rect 35 29 69 63
rect 131 15 165 49
rect 215 38 249 72
rect 299 54 333 88
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 35 275 69 309
rect 209 411 243 445
rect 209 343 243 377
rect 299 411 333 445
rect 299 343 333 377
<< poly >>
rect 79 457 109 483
rect 151 457 181 483
rect 259 457 289 483
rect 259 285 289 317
rect 259 269 347 285
rect 79 225 109 257
rect 38 209 109 225
rect 38 175 48 209
rect 82 175 109 209
rect 38 159 109 175
rect 151 225 181 257
rect 259 235 303 269
rect 337 235 347 269
rect 151 209 207 225
rect 151 175 161 209
rect 195 175 207 209
rect 151 159 207 175
rect 259 219 347 235
rect 79 137 109 159
rect 175 137 205 159
rect 259 137 289 219
rect 79 -19 109 7
rect 175 -19 205 7
rect 259 -19 289 7
<< polycont >>
rect 48 175 82 209
rect 303 235 337 269
rect 161 175 195 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 368 521
rect 18 445 82 487
rect 18 411 35 445
rect 69 411 82 445
rect 193 445 259 453
rect 18 377 82 411
rect 18 343 35 377
rect 69 343 82 377
rect 18 309 82 343
rect 18 275 35 309
rect 69 275 82 309
rect 18 259 82 275
rect 118 225 157 435
rect 193 411 209 445
rect 243 411 259 445
rect 193 377 259 411
rect 193 343 209 377
rect 243 343 259 377
rect 193 317 259 343
rect 299 445 350 487
rect 333 411 350 445
rect 299 377 350 411
rect 333 343 350 377
rect 299 327 350 343
rect 193 261 263 317
rect 30 209 82 225
rect 30 175 48 209
rect 30 159 82 175
rect 118 209 195 225
rect 118 175 161 209
rect 118 159 195 175
rect 229 185 263 261
rect 301 269 350 291
rect 301 235 303 269
rect 337 235 350 269
rect 301 219 350 235
rect 229 151 333 185
rect 18 83 261 117
rect 18 63 76 83
rect 18 29 35 63
rect 69 29 76 63
rect 215 72 261 83
rect 18 13 76 29
rect 115 15 131 49
rect 165 15 181 49
rect 249 38 261 72
rect 299 88 333 151
rect 299 38 333 54
rect 215 22 261 38
rect 115 -23 181 15
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 368 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
<< metal1 >>
rect 0 521 368 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 368 521
rect 0 456 368 487
rect 0 -23 368 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 368 -23
rect 0 -88 368 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 o21ai_1
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 122 385 156 419 0 FreeSans 400 0 0 0 A2
port 7 nsew
flabel locali s 122 317 156 351 0 FreeSans 400 0 0 0 A2
port 7 nsew
flabel locali s 122 249 156 283 0 FreeSans 400 0 0 0 A2
port 7 nsew
flabel locali s 30 181 64 215 0 FreeSans 400 0 0 0 A1
port 10 nsew
flabel locali s 122 181 156 215 0 FreeSans 400 0 0 0 A2
port 7 nsew
flabel locali s 305 249 339 283 0 FreeSans 400 0 0 0 B1
port 8 nsew
flabel locali s 214 385 248 419 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel locali s 214 317 248 351 0 FreeSans 400 0 0 0 Y
port 9 nsew
<< properties >>
string FIXED_BBOX 0 -40 368 504
string path 0.000 12.600 9.200 12.600 
<< end >>
