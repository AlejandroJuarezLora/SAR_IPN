* NGSPICE file created from comparator.ext - technology: sky130B

.subckt sky130_fd_pr__pfet_01v8_QE5SNW a_n78_n136# a_n78_n437# a_n23_95# w_n226_n649#
+ a_n23_n534# a_40_n136# a_n23_460# a_40_n437# a_40_229# a_n78_229#
X0 a_40_n136# a_n23_95# a_n78_n136# w_n226_n649# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X1 a_40_n437# a_n23_n534# a_n78_n437# w_n226_n649# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X2 a_40_229# a_n23_460# a_n78_229# w_n226_n649# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_763N5J D S G B
X0 S G D B sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_FJK8MD m3_n386_n240# c1_n346_n200#
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt trimcap m1_179_405# m1_176_1185#
Xsky130_fd_pr__cap_mim_m3_1_FJK8MD_0 m1_179_405# m1_176_1185# sky130_fd_pr__cap_mim_m3_1_FJK8MD
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_3SNHZA a_n501_n131# a_26_91# a_n383_n131# a_n328_91#
+ a_n446_91# a_443_n131# a_n265_n131# a_n210_91# a_325_n131# a_n147_n131# a_n603_n243#
+ a_207_n131# a_144_91# a_262_91# a_n29_n131# a_380_91# a_n92_91# a_89_n131#
X0 a_n265_n131# a_n328_91# a_n383_n131# a_n603_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 a_89_n131# a_26_91# a_n29_n131# a_n603_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 a_207_n131# a_144_91# a_89_n131# a_n603_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 a_n147_n131# a_n210_91# a_n265_n131# a_n603_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X4 a_443_n131# a_380_91# a_325_n131# a_n603_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X5 a_n383_n131# a_n446_91# a_n501_n131# a_n603_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X6 a_n29_n131# a_n92_91# a_n147_n131# a_n603_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_325_n131# a_262_91# a_207_n131# a_n603_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_FS2HZA a_n367_n243# a_26_91# a_n265_n131# a_n210_91#
+ a_n147_n131# a_207_n131# a_144_91# a_n29_n131# a_n92_91# a_89_n131#
X0 a_89_n131# a_26_91# a_n29_n131# a_n367_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 a_207_n131# a_144_91# a_89_n131# a_n367_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X2 a_n147_n131# a_n210_91# a_n265_n131# a_n367_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X3 a_n29_n131# a_n92_91# a_n147_n131# a_n367_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_THUHZA a_n249_n243# a_26_91# a_n147_n131# a_n29_n131#
+ a_n92_91# a_89_n131#
X0 a_89_n131# a_26_91# a_n29_n131# a_n249_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X1 a_n29_n131# a_n92_91# a_n147_n131# a_n249_n243# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt trim drain d_4_ d_3_ d_2_ d_1_ d_0_ vss
Xsky130_fd_pr__nfet_01v8_lvt_763N5J_0 n1 vss d_1_ vss sky130_fd_pr__nfet_01v8_lvt_763N5J
Xtrimcap_12 n4 drain trimcap
Xtrimcap_11 n4 drain trimcap
Xsky130_fd_pr__nfet_01v8_lvt_763N5J_1 n0 vss d_0_ vss sky130_fd_pr__nfet_01v8_lvt_763N5J
Xtrimcap_13 n4 drain trimcap
Xtrimcap_14 n4 drain trimcap
Xtrimcap_15 n4 drain trimcap
Xsky130_fd_pr__nfet_01v8_lvt_3SNHZA_0 n4 d_4_ vss d_4_ d_4_ n4 n4 d_4_ vss vss vss
+ n4 d_4_ d_4_ n4 d_4_ d_4_ vss sky130_fd_pr__nfet_01v8_lvt_3SNHZA
Xsky130_fd_pr__nfet_01v8_lvt_FS2HZA_0 vss d_3_ n3 d_3_ vss n3 d_3_ n3 d_3_ vss sky130_fd_pr__nfet_01v8_lvt_FS2HZA
Xsky130_fd_pr__nfet_01v8_lvt_THUHZA_0 vss d_2_ n2 vss d_2_ n2 sky130_fd_pr__nfet_01v8_lvt_THUHZA
Xtrimcap_0 n3 drain trimcap
Xtrimcap_2 n3 drain trimcap
Xtrimcap_1 n3 drain trimcap
Xtrimcap_3 n3 drain trimcap
Xtrimcap_4 n2 drain trimcap
Xtrimcap_5 n2 drain trimcap
Xtrimcap_6 n1 drain trimcap
Xtrimcap_7 n0 drain trimcap
Xtrimcap_8 n4 drain trimcap
Xtrimcap_9 n4 drain trimcap
Xtrimcap_10 n4 drain trimcap
.ends

.subckt sky130_fd_pr__nfet_01v8_7UX3DE a_n33_n87# a_30_117# a_30_n309# a_n88_n309#
+ a_n88_117# a_n33_29# a_n190_n421#
X0 a_30_n309# a_n33_n87# a_n88_n309# a_n190_n421# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X1 a_30_117# a_n33_29# a_n88_117# a_n190_n421# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt comparator clk vdd vss outp outn trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ trimb_4_
+ trimb_3_ trimb_2_ trimb_1_ trimb_0_
Xsky130_fd_pr__pfet_01v8_QE5SNW_0 outp outp clk vdd outn vdd clk vdd vdd ip sky130_fd_pr__pfet_01v8_QE5SNW
Xsky130_fd_pr__pfet_01v8_QE5SNW_1 outn outn clk vdd outp vdd clk vdd vdd in sky130_fd_pr__pfet_01v8_QE5SNW
Xtrim_0 in trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ vss trim
Xtrim_1 ip trimb_4_ trimb_3_ trimb_2_ trimb_1_ trimb_0_ vss trim
Xsky130_fd_pr__nfet_01v8_7UX3DE_0 clk vss vss diff diff clk vss sky130_fd_pr__nfet_01v8_7UX3DE
Xsky130_fd_pr__nfet_01v8_7UX3DE_1 outp ip in outn outp outn vss sky130_fd_pr__nfet_01v8_7UX3DE
Xsky130_fd_pr__nfet_01v8_7UX3DE_2 sky130_fd_pr__nfet_01v8_7UX3DE_2/a_n33_n87# diff
+ diff in ip sky130_fd_pr__nfet_01v8_7UX3DE_2/a_n33_29# vss sky130_fd_pr__nfet_01v8_7UX3DE
.ends

