magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 774 542
<< pwell >>
rect 1 -19 735 143
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 657 117
<< scpmoshvt >>
rect 79 283 657 457
<< ndiff >>
rect 27 72 79 117
rect 27 38 35 72
rect 69 38 79 72
rect 27 7 79 38
rect 657 72 709 117
rect 657 38 667 72
rect 701 38 709 72
rect 657 7 709 38
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 343 79 411
rect 27 309 35 343
rect 69 309 79 343
rect 27 283 79 309
rect 657 445 709 457
rect 657 411 667 445
rect 701 411 709 445
rect 657 343 709 411
rect 657 309 667 343
rect 701 309 709 343
rect 657 283 709 309
<< ndiffc >>
rect 35 38 69 72
rect 667 38 701 72
<< pdiffc >>
rect 35 411 69 445
rect 35 309 69 343
rect 667 411 701 445
rect 667 309 701 343
<< poly >>
rect 79 457 657 483
rect 79 257 657 283
rect 79 235 343 257
rect 79 201 95 235
rect 129 201 194 235
rect 228 201 293 235
rect 327 201 343 235
rect 79 185 343 201
rect 385 199 657 215
rect 385 165 401 199
rect 435 165 504 199
rect 538 165 607 199
rect 641 165 657 199
rect 385 143 657 165
rect 79 117 657 143
rect 79 -19 657 7
<< polycont >>
rect 95 201 129 235
rect 194 201 228 235
rect 293 201 327 235
rect 401 165 435 199
rect 504 165 538 199
rect 607 165 641 199
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 17 445 719 487
rect 17 411 35 445
rect 69 411 667 445
rect 701 411 719 445
rect 17 343 719 411
rect 17 309 35 343
rect 69 309 667 343
rect 701 309 719 343
rect 17 269 719 309
rect 17 201 95 235
rect 129 201 194 235
rect 228 201 293 235
rect 327 201 347 235
rect 17 131 347 201
rect 381 199 719 269
rect 381 165 401 199
rect 435 165 504 199
rect 538 165 607 199
rect 641 165 719 199
rect 17 72 719 131
rect 17 38 35 72
rect 69 38 667 72
rect 701 38 719 72
rect 17 -23 719 38
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
<< metal1 >>
rect 0 521 736 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 0 456 736 487
rect 0 -23 736 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
rect 0 -88 736 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 decap_8
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
<< properties >>
string FIXED_BBOX 0 -40 736 504
string path 0.000 -1.000 18.400 -1.000 
<< end >>
