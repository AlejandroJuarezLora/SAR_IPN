magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 406 542
<< pwell >>
rect 4 -19 367 163
rect 29 -57 63 -19
<< scnmos >>
rect 83 7 113 137
rect 169 7 199 137
rect 258 7 288 137
<< scpmoshvt >>
rect 83 257 113 457
rect 169 257 199 457
rect 258 257 288 457
<< ndiff >>
rect 30 53 83 137
rect 30 19 38 53
rect 72 19 83 53
rect 30 7 83 19
rect 113 87 169 137
rect 113 53 124 87
rect 158 53 169 87
rect 113 7 169 53
rect 199 7 258 137
rect 288 83 341 137
rect 288 49 299 83
rect 333 49 341 83
rect 288 7 341 49
<< pdiff >>
rect 30 413 83 457
rect 30 379 38 413
rect 72 379 83 413
rect 30 339 83 379
rect 30 305 38 339
rect 72 305 83 339
rect 30 257 83 305
rect 113 435 169 457
rect 113 401 124 435
rect 158 401 169 435
rect 113 367 169 401
rect 113 333 124 367
rect 158 333 169 367
rect 113 257 169 333
rect 199 449 258 457
rect 199 415 210 449
rect 244 415 258 449
rect 199 257 258 415
rect 288 443 341 457
rect 288 409 299 443
rect 333 409 341 443
rect 288 375 341 409
rect 288 341 299 375
rect 333 341 341 375
rect 288 307 341 341
rect 288 273 299 307
rect 333 273 341 307
rect 288 257 341 273
<< ndiffc >>
rect 38 19 72 53
rect 124 53 158 87
rect 299 49 333 83
<< pdiffc >>
rect 38 379 72 413
rect 38 305 72 339
rect 124 401 158 435
rect 124 333 158 367
rect 210 415 244 449
rect 299 409 333 443
rect 299 341 333 375
rect 299 273 333 307
<< poly >>
rect 83 457 113 483
rect 169 457 199 483
rect 258 457 288 483
rect 83 225 113 257
rect 169 225 199 257
rect 258 225 288 257
rect 21 209 113 225
rect 21 175 31 209
rect 65 175 113 209
rect 21 159 113 175
rect 162 209 216 225
rect 162 175 172 209
rect 206 175 216 209
rect 162 159 216 175
rect 258 209 342 225
rect 258 175 298 209
rect 332 175 342 209
rect 258 159 342 175
rect 83 137 113 159
rect 169 137 199 159
rect 258 137 288 159
rect 83 -19 113 7
rect 169 -19 199 7
rect 258 -19 288 7
<< polycont >>
rect 31 175 65 209
rect 172 175 206 209
rect 298 175 332 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 368 521
rect 19 413 74 451
rect 19 379 38 413
rect 72 379 74 413
rect 19 339 74 379
rect 19 305 38 339
rect 72 305 74 339
rect 108 435 174 451
rect 108 401 124 435
rect 158 401 174 435
rect 108 367 174 401
rect 208 449 247 487
rect 208 415 210 449
rect 244 415 247 449
rect 208 399 247 415
rect 283 443 349 451
rect 283 409 299 443
rect 333 409 349 443
rect 108 333 124 367
rect 158 365 174 367
rect 283 375 349 409
rect 283 365 299 375
rect 158 341 299 365
rect 333 341 349 375
rect 158 333 349 341
rect 108 331 349 333
rect 19 297 74 305
rect 170 307 349 331
rect 19 259 136 297
rect 170 273 299 307
rect 333 273 349 307
rect 170 265 349 273
rect 19 209 67 225
rect 19 175 31 209
rect 65 175 67 209
rect 19 95 67 175
rect 101 125 136 259
rect 170 209 253 225
rect 170 175 172 209
rect 206 175 253 209
rect 170 159 253 175
rect 289 209 348 225
rect 289 175 298 209
rect 332 175 348 209
rect 289 159 348 175
rect 101 89 167 125
rect 122 87 167 89
rect 22 53 88 55
rect 22 19 38 53
rect 72 19 88 53
rect 22 -23 88 19
rect 122 53 124 87
rect 158 53 167 87
rect 122 13 167 53
rect 207 35 253 159
rect 289 83 349 123
rect 289 49 299 83
rect 333 49 349 83
rect 289 -23 349 49
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 368 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
<< metal1 >>
rect 0 521 368 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 368 521
rect 0 456 368 487
rect 0 -23 368 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 368 -23
rect 0 -88 368 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 a21oi_1
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 213 181 247 215 0 FreeSans 200 0 0 0 A1
port 8 nsew
flabel locali s 29 113 63 147 0 FreeSans 200 0 0 0 B1
port 9 nsew
flabel locali s 213 113 247 147 0 FreeSans 200 0 0 0 A1
port 8 nsew
flabel locali s 213 45 247 79 0 FreeSans 200 0 0 0 A1
port 8 nsew
flabel locali s 29 385 63 419 0 FreeSans 200 0 0 0 Y
port 10 nsew
flabel locali s 29 181 63 215 0 FreeSans 200 0 0 0 B1
port 9 nsew
flabel locali s 29 317 63 351 0 FreeSans 200 0 0 0 Y
port 10 nsew
flabel locali s 305 181 339 215 0 FreeSans 200 0 0 0 A2
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 368 504
string path 0.000 12.600 9.200 12.600 
<< end >>
