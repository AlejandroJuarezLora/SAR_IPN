** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/dac/dac.sch
.subckt dac vin sample out ctl_7_,ctl_6_,ctl_5_,ctl_4_,ctl_3_,ctl_2_,ctl_1_,ctl_0_ dum vdd vss
*.ipin vin
*.ipin sample
*.opin out
*.ipin ctl_7_,ctl_6_,ctl_5_,ctl_4_,ctl_3_,ctl_2_,ctl_1_,ctl_0_
*.ipin dum
*.iopin vdd
*.iopin vss
xca out n6 n0 n5 n4 n2 ndum n3 n1 n7 carray
xi6 ctl_6_ vss vss vdd vdd n6 sky130_fd_sc_hd__inv_2
xi5 ctl_5_ vss vss vdd vdd n5 sky130_fd_sc_hd__inv_2
xi4 ctl_4_ vss vss vdd vdd n4 sky130_fd_sc_hd__inv_2
xi3 ctl_3_ vss vss vdd vdd n3 sky130_fd_sc_hd__inv_2
xi2 ctl_2_ vss vss vdd vdd n2 sky130_fd_sc_hd__inv_2
xi1 ctl_1_ vss vss vdd vdd n1 sky130_fd_sc_hd__inv_2
xi0 ctl_0_ vss vss vdd vdd n0 sky130_fd_sc_hd__inv_2
xidum dum vss vss vdd vdd ndum sky130_fd_sc_hd__inv_2
xi7 ctl_7_ vss vss vdd vdd n7 sky130_fd_sc_hd__inv_2
xswt out sample vdd vin vss sw_top
.ends

* expanding   symbol:  sar/dac/carray.sym # of pins=10
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/dac/carray.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/dac/carray.sch
.subckt carray top n6 n0 n5 n4 n2 ndum n3 n1 n7
*.iopin top
*.iopin n7
*.iopin n6
*.iopin n5
*.iopin n4
*.iopin n2
*.iopin n0
*.iopin ndum
*.iopin n3
*.iopin n1
xcdum top ndum unitcap
xc0 top n0 unitcap
xc1_1_ top n1 unitcap
xc1_0_ top n1 unitcap
xc2_3_ top n2 unitcap
xc2_2_ top n2 unitcap
xc2_1_ top n2 unitcap
xc2_0_ top n2 unitcap
xc3_7_ top n3 unitcap
xc3_6_ top n3 unitcap
xc3_5_ top n3 unitcap
xc3_4_ top n3 unitcap
xc3_3_ top n3 unitcap
xc3_2_ top n3 unitcap
xc3_1_ top n3 unitcap
xc3_0_ top n3 unitcap
xc4_15_ top n4 unitcap
xc4_14_ top n4 unitcap
xc4_13_ top n4 unitcap
xc4_12_ top n4 unitcap
xc4_11_ top n4 unitcap
xc4_10_ top n4 unitcap
xc4_9_ top n4 unitcap
xc4_8_ top n4 unitcap
xc4_7_ top n4 unitcap
xc4_6_ top n4 unitcap
xc4_5_ top n4 unitcap
xc4_4_ top n4 unitcap
xc4_3_ top n4 unitcap
xc4_2_ top n4 unitcap
xc4_1_ top n4 unitcap
xc4_0_ top n4 unitcap
xc5_31_ top n5 unitcap
xc5_30_ top n5 unitcap
xc5_29_ top n5 unitcap
xc5_28_ top n5 unitcap
xc5_27_ top n5 unitcap
xc5_26_ top n5 unitcap
xc5_25_ top n5 unitcap
xc5_24_ top n5 unitcap
xc5_23_ top n5 unitcap
xc5_22_ top n5 unitcap
xc5_21_ top n5 unitcap
xc5_20_ top n5 unitcap
xc5_19_ top n5 unitcap
xc5_18_ top n5 unitcap
xc5_17_ top n5 unitcap
xc5_16_ top n5 unitcap
xc5_15_ top n5 unitcap
xc5_14_ top n5 unitcap
xc5_13_ top n5 unitcap
xc5_12_ top n5 unitcap
xc5_11_ top n5 unitcap
xc5_10_ top n5 unitcap
xc5_9_ top n5 unitcap
xc5_8_ top n5 unitcap
xc5_7_ top n5 unitcap
xc5_6_ top n5 unitcap
xc5_5_ top n5 unitcap
xc5_4_ top n5 unitcap
xc5_3_ top n5 unitcap
xc5_2_ top n5 unitcap
xc5_1_ top n5 unitcap
xc5_0_ top n5 unitcap
xc6_63_ top n6 unitcap
xc6_62_ top n6 unitcap
xc6_61_ top n6 unitcap
xc6_60_ top n6 unitcap
xc6_59_ top n6 unitcap
xc6_58_ top n6 unitcap
xc6_57_ top n6 unitcap
xc6_56_ top n6 unitcap
xc6_55_ top n6 unitcap
xc6_54_ top n6 unitcap
xc6_53_ top n6 unitcap
xc6_52_ top n6 unitcap
xc6_51_ top n6 unitcap
xc6_50_ top n6 unitcap
xc6_49_ top n6 unitcap
xc6_48_ top n6 unitcap
xc6_47_ top n6 unitcap
xc6_46_ top n6 unitcap
xc6_45_ top n6 unitcap
xc6_44_ top n6 unitcap
xc6_43_ top n6 unitcap
xc6_42_ top n6 unitcap
xc6_41_ top n6 unitcap
xc6_40_ top n6 unitcap
xc6_39_ top n6 unitcap
xc6_38_ top n6 unitcap
xc6_37_ top n6 unitcap
xc6_36_ top n6 unitcap
xc6_35_ top n6 unitcap
xc6_34_ top n6 unitcap
xc6_33_ top n6 unitcap
xc6_32_ top n6 unitcap
xc6_31_ top n6 unitcap
xc6_30_ top n6 unitcap
xc6_29_ top n6 unitcap
xc6_28_ top n6 unitcap
xc6_27_ top n6 unitcap
xc6_26_ top n6 unitcap
xc6_25_ top n6 unitcap
xc6_24_ top n6 unitcap
xc6_23_ top n6 unitcap
xc6_22_ top n6 unitcap
xc6_21_ top n6 unitcap
xc6_20_ top n6 unitcap
xc6_19_ top n6 unitcap
xc6_18_ top n6 unitcap
xc6_17_ top n6 unitcap
xc6_16_ top n6 unitcap
xc6_15_ top n6 unitcap
xc6_14_ top n6 unitcap
xc6_13_ top n6 unitcap
xc6_12_ top n6 unitcap
xc6_11_ top n6 unitcap
xc6_10_ top n6 unitcap
xc6_9_ top n6 unitcap
xc6_8_ top n6 unitcap
xc6_7_ top n6 unitcap
xc6_6_ top n6 unitcap
xc6_5_ top n6 unitcap
xc6_4_ top n6 unitcap
xc6_3_ top n6 unitcap
xc6_2_ top n6 unitcap
xc6_1_ top n6 unitcap
xc6_0_ top n6 unitcap
xc7_127_ top n7 unitcap
xc7_126_ top n7 unitcap
xc7_125_ top n7 unitcap
xc7_124_ top n7 unitcap
xc7_123_ top n7 unitcap
xc7_122_ top n7 unitcap
xc7_121_ top n7 unitcap
xc7_120_ top n7 unitcap
xc7_119_ top n7 unitcap
xc7_118_ top n7 unitcap
xc7_117_ top n7 unitcap
xc7_116_ top n7 unitcap
xc7_115_ top n7 unitcap
xc7_114_ top n7 unitcap
xc7_113_ top n7 unitcap
xc7_112_ top n7 unitcap
xc7_111_ top n7 unitcap
xc7_110_ top n7 unitcap
xc7_109_ top n7 unitcap
xc7_108_ top n7 unitcap
xc7_107_ top n7 unitcap
xc7_106_ top n7 unitcap
xc7_105_ top n7 unitcap
xc7_104_ top n7 unitcap
xc7_103_ top n7 unitcap
xc7_102_ top n7 unitcap
xc7_101_ top n7 unitcap
xc7_100_ top n7 unitcap
xc7_99_ top n7 unitcap
xc7_98_ top n7 unitcap
xc7_97_ top n7 unitcap
xc7_96_ top n7 unitcap
xc7_95_ top n7 unitcap
xc7_94_ top n7 unitcap
xc7_93_ top n7 unitcap
xc7_92_ top n7 unitcap
xc7_91_ top n7 unitcap
xc7_90_ top n7 unitcap
xc7_89_ top n7 unitcap
xc7_88_ top n7 unitcap
xc7_87_ top n7 unitcap
xc7_86_ top n7 unitcap
xc7_85_ top n7 unitcap
xc7_84_ top n7 unitcap
xc7_83_ top n7 unitcap
xc7_82_ top n7 unitcap
xc7_81_ top n7 unitcap
xc7_80_ top n7 unitcap
xc7_79_ top n7 unitcap
xc7_78_ top n7 unitcap
xc7_77_ top n7 unitcap
xc7_76_ top n7 unitcap
xc7_75_ top n7 unitcap
xc7_74_ top n7 unitcap
xc7_73_ top n7 unitcap
xc7_72_ top n7 unitcap
xc7_71_ top n7 unitcap
xc7_70_ top n7 unitcap
xc7_69_ top n7 unitcap
xc7_68_ top n7 unitcap
xc7_67_ top n7 unitcap
xc7_66_ top n7 unitcap
xc7_65_ top n7 unitcap
xc7_64_ top n7 unitcap
xc7_63_ top n7 unitcap
xc7_62_ top n7 unitcap
xc7_61_ top n7 unitcap
xc7_60_ top n7 unitcap
xc7_59_ top n7 unitcap
xc7_58_ top n7 unitcap
xc7_57_ top n7 unitcap
xc7_56_ top n7 unitcap
xc7_55_ top n7 unitcap
xc7_54_ top n7 unitcap
xc7_53_ top n7 unitcap
xc7_52_ top n7 unitcap
xc7_51_ top n7 unitcap
xc7_50_ top n7 unitcap
xc7_49_ top n7 unitcap
xc7_48_ top n7 unitcap
xc7_47_ top n7 unitcap
xc7_46_ top n7 unitcap
xc7_45_ top n7 unitcap
xc7_44_ top n7 unitcap
xc7_43_ top n7 unitcap
xc7_42_ top n7 unitcap
xc7_41_ top n7 unitcap
xc7_40_ top n7 unitcap
xc7_39_ top n7 unitcap
xc7_38_ top n7 unitcap
xc7_37_ top n7 unitcap
xc7_36_ top n7 unitcap
xc7_35_ top n7 unitcap
xc7_34_ top n7 unitcap
xc7_33_ top n7 unitcap
xc7_32_ top n7 unitcap
xc7_31_ top n7 unitcap
xc7_30_ top n7 unitcap
xc7_29_ top n7 unitcap
xc7_28_ top n7 unitcap
xc7_27_ top n7 unitcap
xc7_26_ top n7 unitcap
xc7_25_ top n7 unitcap
xc7_24_ top n7 unitcap
xc7_23_ top n7 unitcap
xc7_22_ top n7 unitcap
xc7_21_ top n7 unitcap
xc7_20_ top n7 unitcap
xc7_19_ top n7 unitcap
xc7_18_ top n7 unitcap
xc7_17_ top n7 unitcap
xc7_16_ top n7 unitcap
xc7_15_ top n7 unitcap
xc7_14_ top n7 unitcap
xc7_13_ top n7 unitcap
xc7_12_ top n7 unitcap
xc7_11_ top n7 unitcap
xc7_10_ top n7 unitcap
xc7_9_ top n7 unitcap
xc7_8_ top n7 unitcap
xc7_7_ top n7 unitcap
xc7_6_ top n7 unitcap
xc7_5_ top n7 unitcap
xc7_4_ top n7 unitcap
xc7_3_ top n7 unitcap
xc7_2_ top n7 unitcap
xc7_1_ top n7 unitcap
xc7_0_ top n7 unitcap
xdummy_83_ top dum_bot_83_ unitcap
xdummy_82_ top dum_bot_82_ unitcap
xdummy_81_ top dum_bot_81_ unitcap
xdummy_80_ top dum_bot_80_ unitcap
xdummy_79_ top dum_bot_79_ unitcap
xdummy_78_ top dum_bot_78_ unitcap
xdummy_77_ top dum_bot_77_ unitcap
xdummy_76_ top dum_bot_76_ unitcap
xdummy_75_ top dum_bot_75_ unitcap
xdummy_74_ top dum_bot_74_ unitcap
xdummy_73_ top dum_bot_73_ unitcap
xdummy_72_ top dum_bot_72_ unitcap
xdummy_71_ top dum_bot_71_ unitcap
xdummy_70_ top dum_bot_70_ unitcap
xdummy_69_ top dum_bot_69_ unitcap
xdummy_68_ top dum_bot_68_ unitcap
xdummy_67_ top dum_bot_67_ unitcap
xdummy_66_ top dum_bot_66_ unitcap
xdummy_65_ top dum_bot_65_ unitcap
xdummy_64_ top dum_bot_64_ unitcap
xdummy_63_ top dum_bot_63_ unitcap
xdummy_62_ top dum_bot_62_ unitcap
xdummy_61_ top dum_bot_61_ unitcap
xdummy_60_ top dum_bot_60_ unitcap
xdummy_59_ top dum_bot_59_ unitcap
xdummy_58_ top dum_bot_58_ unitcap
xdummy_57_ top dum_bot_57_ unitcap
xdummy_56_ top dum_bot_56_ unitcap
xdummy_55_ top dum_bot_55_ unitcap
xdummy_54_ top dum_bot_54_ unitcap
xdummy_53_ top dum_bot_53_ unitcap
xdummy_52_ top dum_bot_52_ unitcap
xdummy_51_ top dum_bot_51_ unitcap
xdummy_50_ top dum_bot_50_ unitcap
xdummy_49_ top dum_bot_49_ unitcap
xdummy_48_ top dum_bot_48_ unitcap
xdummy_47_ top dum_bot_47_ unitcap
xdummy_46_ top dum_bot_46_ unitcap
xdummy_45_ top dum_bot_45_ unitcap
xdummy_44_ top dum_bot_44_ unitcap
xdummy_43_ top dum_bot_43_ unitcap
xdummy_42_ top dum_bot_42_ unitcap
xdummy_41_ top dum_bot_41_ unitcap
xdummy_40_ top dum_bot_40_ unitcap
xdummy_39_ top dum_bot_39_ unitcap
xdummy_38_ top dum_bot_38_ unitcap
xdummy_37_ top dum_bot_37_ unitcap
xdummy_36_ top dum_bot_36_ unitcap
xdummy_35_ top dum_bot_35_ unitcap
xdummy_34_ top dum_bot_34_ unitcap
xdummy_33_ top dum_bot_33_ unitcap
xdummy_32_ top dum_bot_32_ unitcap
xdummy_31_ top dum_bot_31_ unitcap
xdummy_30_ top dum_bot_30_ unitcap
xdummy_29_ top dum_bot_29_ unitcap
xdummy_28_ top dum_bot_28_ unitcap
xdummy_27_ top dum_bot_27_ unitcap
xdummy_26_ top dum_bot_26_ unitcap
xdummy_25_ top dum_bot_25_ unitcap
xdummy_24_ top dum_bot_24_ unitcap
xdummy_23_ top dum_bot_23_ unitcap
xdummy_22_ top dum_bot_22_ unitcap
xdummy_21_ top dum_bot_21_ unitcap
xdummy_20_ top dum_bot_20_ unitcap
xdummy_19_ top dum_bot_19_ unitcap
xdummy_18_ top dum_bot_18_ unitcap
xdummy_17_ top dum_bot_17_ unitcap
xdummy_16_ top dum_bot_16_ unitcap
xdummy_15_ top dum_bot_15_ unitcap
xdummy_14_ top dum_bot_14_ unitcap
xdummy_13_ top dum_bot_13_ unitcap
xdummy_12_ top dum_bot_12_ unitcap
xdummy_11_ top dum_bot_11_ unitcap
xdummy_10_ top dum_bot_10_ unitcap
xdummy_9_ top dum_bot_9_ unitcap
xdummy_8_ top dum_bot_8_ unitcap
xdummy_7_ top dum_bot_7_ unitcap
xdummy_6_ top dum_bot_6_ unitcap
xdummy_5_ top dum_bot_5_ unitcap
xdummy_4_ top dum_bot_4_ unitcap
xdummy_3_ top dum_bot_3_ unitcap
xdummy_2_ top dum_bot_2_ unitcap
xdummy_1_ top dum_bot_1_ unitcap
xdummy_0_ top dum_bot_0_ unitcap
.ends


* expanding   symbol:  sar/sw/sw_top.sym # of pins=5
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/sw/sw_top.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/sw/sw_top.sch
.subckt sw_top out en vdd in vss
*.iopin out
*.ipin en
*.iopin vss
*.iopin vdd
*.iopin in
x2 vss vss vdd vdd sky130_fd_sc_hd__decap_8
x4 en vss vss vdd vdd en_buf sky130_fd_sc_hd__inv_4
x1 VGND VNB VPB VPWR sky130_fd_sc_hd__decap_3
XM1 in en out vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM2 in en_buf out vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
.ends


* expanding   symbol:  sar/unitcap/unitcap.sym # of pins=2
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/unitcap/unitcap.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/unitcap/unitcap.sch
.subckt unitcap cp cn
*.iopin cp
*.iopin cn
XC2 cp cn sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=1 m=1
.ends

.end
