magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 682 542
<< pwell >>
rect 1 -19 585 163
rect 30 -57 64 -19
<< scnmos >>
rect 80 7 110 137
rect 179 7 209 137
rect 273 7 303 137
rect 369 7 399 137
rect 465 7 495 137
<< scpmoshvt >>
rect 80 257 110 457
rect 179 257 209 457
rect 273 257 303 457
rect 369 257 399 457
rect 465 257 495 457
<< ndiff >>
rect 27 122 80 137
rect 27 88 35 122
rect 69 88 80 122
rect 27 54 80 88
rect 27 20 35 54
rect 69 20 80 54
rect 27 7 80 20
rect 110 57 179 137
rect 110 23 135 57
rect 169 23 179 57
rect 110 7 179 23
rect 209 7 273 137
rect 303 7 369 137
rect 399 125 465 137
rect 399 91 411 125
rect 445 91 465 125
rect 399 57 465 91
rect 399 23 411 57
rect 445 23 465 57
rect 399 7 465 23
rect 495 57 559 137
rect 495 23 511 57
rect 545 23 559 57
rect 495 7 559 23
<< pdiff >>
rect 27 445 80 457
rect 27 411 35 445
rect 69 411 80 445
rect 27 377 80 411
rect 27 343 35 377
rect 69 343 80 377
rect 27 309 80 343
rect 27 275 35 309
rect 69 275 80 309
rect 27 257 80 275
rect 110 445 179 457
rect 110 411 127 445
rect 161 411 179 445
rect 110 377 179 411
rect 110 343 127 377
rect 161 343 179 377
rect 110 309 179 343
rect 110 275 127 309
rect 161 275 179 309
rect 110 257 179 275
rect 209 427 273 457
rect 209 393 223 427
rect 257 393 273 427
rect 209 359 273 393
rect 209 325 223 359
rect 257 325 273 359
rect 209 257 273 325
rect 303 427 369 457
rect 303 393 319 427
rect 353 393 369 427
rect 303 257 369 393
rect 399 427 465 457
rect 399 393 415 427
rect 449 393 465 427
rect 399 359 465 393
rect 399 325 415 359
rect 449 325 465 359
rect 399 257 465 325
rect 495 445 559 457
rect 495 411 517 445
rect 551 411 559 445
rect 495 359 559 411
rect 495 325 517 359
rect 551 325 559 359
rect 495 257 559 325
<< ndiffc >>
rect 35 88 69 122
rect 35 20 69 54
rect 135 23 169 57
rect 411 91 445 125
rect 411 23 445 57
rect 511 23 545 57
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 35 275 69 309
rect 127 411 161 445
rect 127 343 161 377
rect 127 275 161 309
rect 223 393 257 427
rect 223 325 257 359
rect 319 393 353 427
rect 415 393 449 427
rect 415 325 449 359
rect 517 411 551 445
rect 517 325 551 359
<< poly >>
rect 80 457 110 483
rect 179 457 209 483
rect 273 457 303 483
rect 369 457 399 483
rect 465 457 495 483
rect 80 225 110 257
rect 179 225 209 257
rect 273 225 303 257
rect 369 225 399 257
rect 465 225 495 257
rect 80 209 135 225
rect 80 175 91 209
rect 125 175 135 209
rect 80 159 135 175
rect 177 209 231 225
rect 177 175 187 209
rect 221 175 231 209
rect 177 159 231 175
rect 273 209 327 225
rect 273 175 283 209
rect 317 175 327 209
rect 273 159 327 175
rect 369 209 423 225
rect 369 175 379 209
rect 413 175 423 209
rect 369 159 423 175
rect 465 209 519 225
rect 465 175 475 209
rect 509 175 519 209
rect 465 159 519 175
rect 80 137 110 159
rect 179 137 209 159
rect 273 137 303 159
rect 369 137 399 159
rect 465 137 495 159
rect 80 -19 110 7
rect 179 -19 209 7
rect 273 -19 303 7
rect 369 -19 399 7
rect 465 -19 495 7
<< polycont >>
rect 91 175 125 209
rect 187 175 221 209
rect 283 175 317 209
rect 379 175 413 209
rect 475 175 509 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 644 521
rect 119 445 169 487
rect 19 411 35 445
rect 69 411 85 445
rect 19 377 85 411
rect 19 343 35 377
rect 69 343 85 377
rect 19 309 85 343
rect 19 275 35 309
rect 69 275 85 309
rect 119 411 127 445
rect 161 411 169 445
rect 119 377 169 411
rect 119 343 127 377
rect 161 343 169 377
rect 119 309 169 343
rect 207 427 257 443
rect 207 393 223 427
rect 303 427 369 487
rect 303 393 319 427
rect 353 393 369 427
rect 415 427 465 443
rect 449 393 465 427
rect 207 359 257 393
rect 415 359 465 393
rect 207 325 223 359
rect 257 325 415 359
rect 449 325 465 359
rect 501 411 517 445
rect 551 411 567 445
rect 501 359 567 411
rect 501 325 517 359
rect 551 325 592 359
rect 119 275 127 309
rect 161 275 169 309
rect 19 122 57 275
rect 119 259 169 275
rect 205 225 248 291
rect 91 209 153 225
rect 125 175 153 209
rect 91 159 153 175
rect 187 209 248 225
rect 221 175 248 209
rect 187 159 248 175
rect 283 209 340 291
rect 317 175 340 209
rect 283 159 340 175
rect 379 209 432 291
rect 413 175 432 209
rect 379 159 432 175
rect 475 209 524 291
rect 509 175 524 209
rect 475 159 524 175
rect 119 125 153 159
rect 558 125 592 325
rect 19 88 35 122
rect 69 88 85 122
rect 119 91 411 125
rect 445 91 592 125
rect 19 54 85 88
rect 395 57 461 91
rect 19 20 35 54
rect 69 20 85 54
rect 119 23 135 57
rect 169 23 185 57
rect 395 23 411 57
rect 445 23 461 57
rect 495 23 511 57
rect 545 23 561 57
rect 119 -23 185 23
rect 495 -23 561 23
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 644 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
<< metal1 >>
rect 0 521 644 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 644 521
rect 0 456 644 487
rect 0 -23 644 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 644 -23
rect 0 -88 644 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 a31o_1
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 306 249 340 283 0 FreeSans 200 0 0 0 A2
port 9 nsew
flabel locali s 490 249 524 283 0 FreeSans 200 0 0 0 B1
port 11 nsew
flabel locali s 398 181 432 215 0 FreeSans 200 0 0 0 A1
port 10 nsew
flabel locali s 214 249 248 283 0 FreeSans 200 0 0 0 A3
port 8 nsew
flabel locali s 306 181 340 215 0 FreeSans 200 0 0 0 A2
port 9 nsew
flabel locali s 214 181 248 215 0 FreeSans 200 0 0 0 A3
port 8 nsew
flabel locali s 30 385 64 419 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 398 249 432 283 0 FreeSans 200 0 0 0 A1
port 10 nsew
flabel locali s 30 317 64 351 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 30 45 64 79 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 490 181 524 215 0 FreeSans 200 0 0 0 B1
port 11 nsew
<< properties >>
string FIXED_BBOX 0 -40 644 504
string path 0.000 -1.000 16.100 -1.000 
<< end >>
