* SPICE3 file created from SAR.ext - technology: sky130B

.subckt SAR comp ctln1 ctln0 ctlp1 ctlp0 ctln7 ctln6 ctln5 ctln4 ctln3 ctln2 trim4
+ trim1 trim0 trim2 trim3 trimb3 trimb2 trimb0 trimb1 trimb4 ctlp2 ctlp3 ctlp4 ctlp5
+ ctlp6 ctlp7 clkc result7 result6 result5 result4 rstn result3 result2 result1 result0
+ valid cal en clk dvdd avdd avss vinp vinn
X0 avss avdd avss avss sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=260 ps=2.74k w=0.55 l=0.59
X1 avdd avss avdd avdd sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=31.7 ps=307 w=0.87 l=0.59
C0 DAC_1/out DAC_1/carray_0/n4 12.2f
C1 DAC_0/carray_0/m3_26900_1156# DAC_0/carray_0/m3_27100_1156# 3.35f
C2 sarlogic_0/_341_/Q dvdd 2.26f
C3 DAC_1/carray_0/m3_34700_1156# DAC_1/carray_0/n7 4.08f
C4 DAC_0/carray_0/m2_16400_1156# DAC_0/carray_0/n5 2.39f
C5 sarlogic_0/_297_/Y dvdd 2.88f
C6 DAC_1/carray_0/m2_29800_1156# DAC_1/carray_0/n7 3.52f
C7 DAC_0/carray_0/m3_8700_1156# DAC_0/carray_0/n7 2.16f
C8 vinn avdd 3.42f
C9 DAC_0/carray_0/m3_16500_1156# DAC_0/carray_0/m3_16700_1156# 3.35f
C10 sarlogic_0/_188_/S dvdd 2.15f
C11 comparator_0/trim_1/drain comparator_0/trim_1/n3 3.41f
C12 DAC_0/carray_0/m3_7400_1156# DAC_0/carray_0/m3_7600_1156# 3.35f
C13 DAC_0/carray_0/m3_18000_1156# DAC_0/carray_0/n7 3.1f
C14 sarlogic_0/_263_/B dvdd 2.11f
C15 DAC_0/carray_0/m2_13800_1156# DAC_0/carray_0/n7 3.52f
C16 DAC_1/carray_0/m3_37300_1156# DAC_1/carray_0/n6 4.09f
C17 sarlogic_0/_298_/C dvdd 2.1f
C18 DAC_1/carray_0/m3_39900_1156# DAC_1/carray_0/m3_40100_1156# 3.35f
C19 DAC_1/carray_0/m2_37600_1156# DAC_1/carray_0/m3_37500_1156# 2.11f
C20 DAC_0/carray_0/m3_29500_1156# DAC_0/carray_0/n7 3.1f
C21 DAC_1/carray_0/m3_36000_1156# DAC_1/carray_0/n7 4.08f
C22 DAC_1/carray_0/m3_30800_1156# DAC_1/carray_0/m3_31000_1156# 3.35f
C23 DAC_0/carray_0/m2_24600_1156# DAC_0/carray_0/m3_24500_1156# 2.11f
C24 DAC_0/out DAC_0/carray_0/n7 97.2f
C25 DAC_1/carray_0/m2_28500_1156# DAC_1/carray_0/m3_28400_1156# 2.11f
C26 DAC_1/carray_0/m3_10200_1156# DAC_1/carray_0/n5 4.08f
C27 DAC_1/out DAC_1/carray_0/n5 24.3f
C28 sample DAC_1/carray_0/n7 4.96f
C29 DAC_0/carray_0/m2_15100_1156# DAC_0/carray_0/m3_15200_1156# 2.11f
C30 sample DAC_1/carray_0/ndum 11.1f
C31 DAC_0/carray_0/m3_38800_1156# DAC_0/carray_0/n7 2.16f
C32 sarlogic_0/_286_/B sarlogic_0/_306_/S 3.15f
C33 DAC_0/carray_0/m3_33400_1156# DAC_0/carray_0/n5 4.08f
C34 DAC_0/carray_0/m3_2400_1156# DAC_0/carray_0/n6 4.08f
C35 avdd DAC_1/sw_top_3/m2_1158_361# 2.15f
C36 DAC_1/carray_0/m3_11300_1156# DAC_1/carray_0/m3_11500_1156# 3.35f
C37 DAC_0/carray_0/n5 DAC_0/carray_0/n6 17.4f
C38 DAC_0/carray_0/n3 DAC_0/carray_0/n1 3.36f
C39 DAC_1/carray_0/m2_2100_1156# DAC_1/carray_0/m3_2200_1156# 2.11f
C40 DAC_0/carray_0/m3_32100_1156# DAC_0/carray_0/n6 4.08f
C41 DAC_0/carray_0/m2_15100_1156# DAC_0/carray_0/n7 2.39f
C42 DAC_0/carray_0/m2_20300_1156# DAC_0/carray_0/m3_20400_1156# 2.11f
C43 ctlp6 ctlp5 2.33f
C44 DAC_0/carray_0/m3_37300_1156# DAC_0/carray_0/m3_37500_1156# 3.35f
C45 DAC_1/carray_0/m3_2200_1156# DAC_1/carray_0/m3_2400_1156# 3.35f
C46 DAC_0/carray_0/m3_1100_1156# DAC_0/carray_0/n7 4.08f
C47 DAC_0/carray_0/m2_35000_1156# DAC_0/carray_0/m3_34900_1156# 2.11f
C48 avdd DAC_1/sw_top_0/m2_1158_361# 2.15f
C49 DAC_1/carray_0/m3_7600_1156# DAC_1/carray_0/n7 4.08f
C50 DAC_1/carray_0/n7 DAC_1/carray_0/n1 11.4f
C51 DAC_1/carray_0/ndum DAC_1/carray_0/n1 3.54f
C52 DAC_0/carray_0/m2_7300_1156# DAC_0/carray_0/m3_7400_1156# 2.11f
C53 DAC_0/carray_0/m3_30800_1156# DAC_0/carray_0/n7 3.14f
C54 vinp avdd 3.42f
C55 DAC_0/carray_0/m3_28200_1156# DAC_0/carray_0/m3_28400_1156# 3.35f
C56 DAC_0/carray_0/m2_24600_1156# DAC_0/carray_0/n7 2.39f
C57 sarlogic_0/_216_/A sarlogic_0/_215_/A 2.43f
C58 DAC_1/carray_0/m2_7300_1156# DAC_1/carray_0/n6 2.39f
C59 DAC_0/carray_0/m3_17800_1156# DAC_0/carray_0/m3_18000_1156# 3.35f
C60 DAC_1/carray_0/m3_24300_1156# DAC_1/carray_0/n4 4.08f
C61 DAC_1/carray_0/m2_6000_1156# DAC_1/carray_0/n7 2.39f
C62 DAC_0/carray_0/m2_3400_1156# DAC_0/carray_0/n6 2.39f
C63 DAC_0/carray_0/m3_8700_1156# DAC_0/carray_0/m3_8900_1156# 3.35f
C64 DAC_1/carray_0/n2 DAC_1/carray_0/n1 2.02f
C65 DAC_1/out DAC_1/carray_0/n6 48.6f
C66 DAC_1/carray_0/m2_9900_1156# DAC_1/carray_0/m3_10000_1156# 2.11f
C67 DAC_0/carray_0/m2_2100_1156# DAC_0/carray_0/n7 2.39f
C68 sarlogic_0/_160_/X dvdd 3.77f
C69 DAC_1/carray_0/m3_41200_1156# DAC_1/carray_0/m3_41400_1156# 3.35f
C70 comparator_0/trim_1/drain comparator_0/trim_1/n4 6.89f
C71 DAC_1/carray_0/m3_8900_1156# DAC_1/carray_0/n7 4.08f
C72 sarlogic_0/_172_/A dvdd 6.02f
C73 DAC_1/carray_0/m2_38900_1156# DAC_1/carray_0/m3_38800_1156# 2.11f
C74 sarlogic_0/_246_/B dvdd 2.08f
C75 DAC_0/carray_0/m2_8600_1156# DAC_0/carray_0/n7 3.52f
C76 DAC_0/carray_0/n2 DAC_0/carray_0/n3 20.7f
C77 DAC_1/carray_0/m3_38600_1156# DAC_1/carray_0/n7 4.08f
C78 clk rstn 3.17f
C79 DAC_1/carray_0/m3_32100_1156# DAC_1/carray_0/m3_32300_1156# 3.35f
C80 DAC_1/carray_0/m2_33700_1156# DAC_1/carray_0/n7 2.39f
C81 DAC_1/carray_0/m2_27200_1156# DAC_1/carray_0/n5 2.39f
C82 DAC_1/carray_0/m2_29800_1156# DAC_1/carray_0/m3_29700_1156# 2.11f
C83 DAC_0/carray_0/m2_16400_1156# DAC_0/carray_0/m3_16500_1156# 2.11f
C84 avdd DAC_1/enb 4.27f
C85 result5 result6 2.6f
C86 DAC_1/carray_0/m2_25900_1156# DAC_1/carray_0/n6 2.39f
C87 DAC_1/carray_0/m2_20300_1156# DAC_1/carray_0/n4 2.39f
C88 result4 result5 2.32f
C89 DAC_0/sw_top_0/m2_1158_361# avdd 2.15f
C90 DAC_1/carray_0/m3_12600_1156# DAC_1/carray_0/m3_12800_1156# 3.35f
C91 DAC_1/carray_0/m3_11500_1156# DAC_1/carray_0/n6 4.08f
C92 DAC_1/carray_0/m3_29700_1156# DAC_1/carray_0/n7 2.16f
C93 sarlogic_0/_191_/B dvdd 2.19f
C94 DAC_1/carray_0/m2_3400_1156# DAC_1/carray_0/m3_3500_1156# 2.11f
C95 ctlp0 ctlp1 3.52f
C96 DAC_1/carray_0/m3_41200_1156# DAC_1/carray_0/n6 4.08f
C97 DAC_0/carray_0/m3_38600_1156# DAC_0/carray_0/m3_38800_1156# 3.35f
C98 sarlogic_0/_306_/S dvdd 3.44f
C99 DAC_1/carray_0/m3_3500_1156# DAC_1/carray_0/m3_3700_1156# 3.35f
C100 DAC_0/out DAC_0/carray_0/n2 3.35f
C101 DAC_0/carray_0/m3_3700_1156# DAC_0/carray_0/n7 4.08f
C102 DAC_0/carray_0/m2_36300_1156# DAC_0/carray_0/m3_36200_1156# 2.11f
C103 sarlogic_0/_248_/B dvdd 3.2f
C104 DAC_1/out DAC_1/carray_0/n7 97.2f
C105 sarlogic_0/_215_/A dvdd 4.19f
C106 DAC_0/carray_0/m3_29500_1156# DAC_0/carray_0/m3_29700_1156# 3.35f
C107 DAC_1/carray_0/m3_39900_1156# DAC_1/carray_0/n7 4.08f
C108 DAC_1/carray_0/m2_17700_1156# DAC_1/carray_0/n6 2.39f
C109 DAC_0/carray_0/m2_28500_1156# DAC_0/carray_0/n7 2.42f
C110 DAC_1/carray_0/m2_35000_1156# DAC_1/carray_0/n7 3.52f
C111 DAC_0/carray_0/m3_13900_1156# DAC_0/carray_0/n7 2.16f
C112 DAC_0/carray_0/n6 DAC_0/carray_0/n7 22.1f
C113 DAC_0/carray_0/m3_19100_1156# DAC_0/carray_0/m3_19300_1156# 3.35f
C114 sarlogic_0/_297_/B dvdd 5.86f
C115 DAC_0/carray_0/m2_4700_1156# DAC_0/carray_0/m3_4800_1156# 2.11f
C116 sarlogic_0/_318_/Q dvdd 2.49f
C117 sarlogic_0/_286_/B dvdd 3.19f
C118 DAC_0/carray_0/m2_32400_1156# DAC_0/carray_0/n5 2.39f
C119 DAC_0/carray_0/m3_10000_1156# DAC_0/carray_0/m3_10200_1156# 3.35f
C120 sarlogic_0/repeater43/X dvdd 6.68f
C121 DAC_1/out DAC_1/carray_0/n2 3.35f
C122 DAC_0/carray_0/m3_6300_1156# DAC_0/carray_0/n6 4.08f
C123 DAC_1/carray_0/m2_11200_1156# DAC_1/carray_0/m3_11300_1156# 2.11f
C124 sarlogic_0/_194_/A dvdd 2.15f
C125 sarlogic_0/_331_/CLK dvdd 8.04f
C126 DAC_0/carray_0/m3_900_1156# DAC_0/carray_0/m3_1100_1156# 3.35f
C127 DAC_0/carray_0/m2_31100_1156# DAC_0/carray_0/n6 2.39f
C128 DAC_1/carray_0/m2_25900_1156# DAC_1/carray_0/m3_25800_1156# 2.11f
C129 DAC_0/carray_0/m3_5000_1156# DAC_0/carray_0/n7 4.08f
C130 DAC_1/carray_0/m3_42500_1156# DAC_1/carray_0/m3_42700_1156# 3.35f
C131 sarlogic_0/_324_/Q dvdd 2.94f
C132 DAC_1/carray_0/n2 DAC_1/carray_0/m3_20400_1156# 3.43f
C133 DAC_1/carray_0/m2_40200_1156# DAC_1/carray_0/m3_40100_1156# 2.11f
C134 DAC_0/carray_0/m3_34700_1156# DAC_0/carray_0/n7 4.08f
C135 DAC_0/carray_0/m2_29800_1156# DAC_0/carray_0/n7 3.52f
C136 DAC_1/carray_0/m3_33400_1156# DAC_1/carray_0/m3_33600_1156# 3.35f
C137 sarlogic_0/_267_/A dvdd 2.48f
C138 DAC_1/carray_0/m2_31100_1156# DAC_1/carray_0/m3_31000_1156# 2.11f
C139 DAC_1/carray_0/m3_15400_1156# DAC_1/carray_0/n5 4.08f
C140 DAC_1/carray_0/m3_24300_1156# DAC_1/carray_0/m3_24500_1156# 3.35f
C141 result6 result7 3.09f
C142 sarlogic_0/_255_/B dvdd 2.22f
C143 DAC_1/carray_0/m3_13900_1156# DAC_1/carray_0/m3_14100_1156# 3.35f
C144 DAC_0/carray_0/m3_37300_1156# DAC_0/carray_0/n6 4.09f
C145 DAC_1/carray_0/n3 DAC_1/carray_0/n4 12.1f
C146 sarlogic_0/_196_/A dvdd 3.27f
C147 DAC_0/carray_0/m3_39900_1156# DAC_0/carray_0/m3_40100_1156# 3.35f
C148 DAC_1/carray_0/m3_4800_1156# DAC_1/carray_0/m3_5000_1156# 3.35f
C149 DAC_0/carray_0/m2_37600_1156# DAC_0/carray_0/m3_37500_1156# 2.11f
C150 DAC_1/carray_0/m3_12800_1156# DAC_1/carray_0/n7 4.08f
C151 DAC_0/carray_0/m3_36000_1156# DAC_0/carray_0/n7 4.08f
C152 DAC_1/carray_0/m2_800_1156# DAC_1/carray_0/m3_900_1156# 2.11f
C153 DAC_0/carray_0/m3_30800_1156# DAC_0/carray_0/m3_31000_1156# 3.35f
C154 DAC_1/carray_0/m3_42500_1156# DAC_1/carray_0/n7 4.08f
C155 DAC_0/carray_0/m2_28500_1156# DAC_0/carray_0/m3_28400_1156# 2.11f
C156 sarlogic_0/_332_/Q dvdd 2.8f
C157 DAC_1/carray_0/m2_37600_1156# DAC_1/carray_0/n7 2.39f
C158 DAC_0/carray_0/m3_10200_1156# DAC_0/carray_0/n5 4.08f
C159 sarlogic_0/_327_/Q dvdd 2.22f
C160 sarlogic_0/_192_/B dvdd 2.35f
C161 DAC_0/carray_0/n2 DAC_0/carray_0/m3_23200_1156# 3.4f
C162 DAC_1/carray_0/m2_19000_1156# DAC_1/carray_0/n7 2.42f
C163 avdd DAC_0/enb 4.27f
C164 DAC_1/carray_0/m2_23300_1156# DAC_1/carray_0/n4 2.39f
C165 DAC_0/carray_0/m3_11300_1156# DAC_0/carray_0/m3_11500_1156# 3.35f
C166 DAC_1/carray_0/m3_4800_1156# DAC_1/carray_0/n7 2.16f
C167 sarlogic_0/clkbuf_2_1_0_clk/A dvdd 4.64f
C168 DAC_0/carray_0/m2_2100_1156# DAC_0/carray_0/m3_2200_1156# 2.11f
C169 DAC_1/carray_0/m2_12500_1156# DAC_1/carray_0/m3_12600_1156# 2.11f
C170 DAC_1/carray_0/m3_28200_1156# DAC_1/carray_0/n5 4.09f
C171 DAC_0/carray_0/m3_2200_1156# DAC_0/carray_0/m3_2400_1156# 3.35f
C172 sarlogic_0/_319_/Q dvdd 4.95f
C173 DAC_1/carray_0/m2_27200_1156# DAC_1/carray_0/m3_27100_1156# 2.11f
C174 DAC_1/carray_0/m2_40200_1156# DAC_1/carray_0/n6 2.39f
C175 DAC_0/carray_0/m3_7600_1156# DAC_0/carray_0/n7 4.08f
C176 DAC_0/carray_0/n7 DAC_0/carray_0/n1 11.4f
C177 DAC_1/carray_0/m3_14100_1156# DAC_1/carray_0/n7 4.08f
C178 DAC_1/carray_0/m2_41500_1156# DAC_1/carray_0/m3_41400_1156# 2.11f
C179 DAC_1/carray_0/m2_8600_1156# DAC_1/carray_0/m3_8700_1156# 2.11f
C180 DAC_1/carray_0/m3_26900_1156# DAC_1/carray_0/n6 4.08f
C181 DAC_0/carray_0/n0 DAC_0/carray_0/n1 14.5f
C182 DAC_1/carray_0/m2_9900_1156# DAC_1/carray_0/n7 2.39f
C183 DAC_1/carray_0/m3_19300_1156# DAC_1/carray_0/n4 4.08f
C184 DAC_0/carray_0/m2_7300_1156# DAC_0/carray_0/n6 2.39f
C185 DAC_1/carray_0/m2_17700_1156# DAC_1/carray_0/m3_17800_1156# 2.11f
C186 DAC_1/carray_0/m3_34700_1156# DAC_1/carray_0/m3_34900_1156# 3.35f
C187 DAC_1/carray_0/m2_38900_1156# DAC_1/carray_0/n7 3.52f
C188 DAC_1/carray_0/m2_32400_1156# DAC_1/carray_0/m3_32300_1156# 2.11f
C189 sarlogic_0/_346_/SET_B dvdd 7.91f
C190 DAC_1/carray_0/m3_25600_1156# DAC_1/carray_0/n7 4.08f
C191 DAC_0/carray_0/m3_24300_1156# DAC_0/carray_0/n4 4.08f
C192 DAC_0/carray_0/m2_6000_1156# DAC_0/carray_0/n7 2.39f
C193 DAC_1/carray_0/m3_25600_1156# DAC_1/carray_0/m3_25800_1156# 3.35f
C194 DAC_1/carray_0/ndum DAC_1/carray_0/n0 14.5f
C195 sarlogic_0/_343_/CLK dvdd 4.6f
C196 sarlogic_0/_279_/Y dvdd 2.16f
C197 DAC_1/carray_0/m3_15200_1156# DAC_1/carray_0/m3_15400_1156# 3.35f
C198 DAC_0/carray_0/m2_9900_1156# DAC_0/carray_0/m3_10000_1156# 2.11f
C199 DAC_1/carray_0/m3_16700_1156# DAC_1/carray_0/n6 3.14f
C200 DAC_1/carray_0/m2_12500_1156# DAC_1/carray_0/n6 2.39f
C201 DAC_1/carray_0/m2_4700_1156# DAC_1/carray_0/n7 3.52f
C202 DAC_0/carray_0/m3_41200_1156# DAC_0/carray_0/m3_41400_1156# 3.35f
C203 DAC_1/carray_0/m3_6100_1156# DAC_1/carray_0/m3_6300_1156# 3.35f
C204 DAC_0/carray_0/ndum DAC_0/carray_0/n0 14.5f
C205 DAC_0/carray_0/m3_8900_1156# DAC_0/carray_0/n7 4.08f
C206 DAC_0/carray_0/m2_38900_1156# DAC_0/carray_0/m3_38800_1156# 2.11f
C207 ctln1 ctln0 3.52f
C208 DAC_0/carray_0/m3_38600_1156# DAC_0/carray_0/n7 4.08f
C209 DAC_0/carray_0/m3_32100_1156# DAC_0/carray_0/m3_32300_1156# 3.35f
C210 DAC_0/carray_0/m2_33700_1156# DAC_0/carray_0/n7 2.39f
C211 sarlogic_0/_342_/Q dvdd 3.01f
C212 DAC_0/carray_0/m2_27200_1156# DAC_0/carray_0/n5 2.39f
C213 DAC_0/carray_0/m2_29800_1156# DAC_0/carray_0/m3_29700_1156# 2.11f
C214 ctlp6 ctlp7 2.73f
C215 sarlogic_0/_258_/S dvdd 3.42f
C216 vinn DAC_1/out 21.5f
C217 DAC_1/carray_0/n4 DAC_1/carray_0/n5 12.7f
C218 DAC_0/carray_0/m2_25900_1156# DAC_0/carray_0/n6 2.39f
C219 DAC_0/carray_0/m2_20300_1156# DAC_0/carray_0/n4 2.39f
C220 DAC_1/carray_0/m2_23300_1156# DAC_1/carray_0/m3_23200_1156# 2.11f
C221 DAC_0/carray_0/m3_12600_1156# DAC_0/carray_0/m3_12800_1156# 3.35f
C222 DAC_0/carray_0/m3_11500_1156# DAC_0/carray_0/n6 4.08f
C223 DAC_1/carray_0/n0 DAC_1/carray_0/n1 14.5f
C224 DAC_0/carray_0/m3_29700_1156# DAC_0/carray_0/n7 2.16f
C225 sarlogic_0/_304_/S dvdd 2.79f
C226 DAC_0/carray_0/m2_3400_1156# DAC_0/carray_0/m3_3500_1156# 2.11f
C227 sarlogic_0/input4/X dvdd 4.66f
C228 DAC_1/carray_0/m2_13800_1156# DAC_1/carray_0/m3_13900_1156# 2.11f
C229 DAC_0/carray_0/m3_41200_1156# DAC_0/carray_0/n6 4.08f
C230 clk dvdd 3.2f
C231 DAC_0/carray_0/m3_3500_1156# DAC_0/carray_0/m3_3700_1156# 3.35f
C232 sarlogic_0/_217_/X dvdd 3.5f
C233 DAC_1/carray_0/m2_42800_1156# DAC_1/carray_0/m3_42700_1156# 2.11f
C234 DAC_0/carray_0/m3_39900_1156# DAC_0/carray_0/n7 4.08f
C235 DAC_0/carray_0/ndum DAC_0/carray_0/n1 3.54f
C236 DAC_0/carray_0/m2_17700_1156# DAC_0/carray_0/n6 2.39f
C237 sarlogic_0/_242_/A dvdd 3.85f
C238 DAC_1/carray_0/m2_19000_1156# DAC_1/carray_0/m3_19100_1156# 2.11f
C239 ctln5 ctln6 2.34f
C240 DAC_0/out DAC_1/out 10.2f
C241 DAC_0/carray_0/m2_35000_1156# DAC_0/carray_0/n7 3.52f
C242 DAC_1/carray_0/m3_36000_1156# DAC_1/carray_0/m3_36200_1156# 3.35f
C243 DAC_1/carray_0/m2_41500_1156# DAC_1/carray_0/n7 2.39f
C244 sarlogic_0/input4/X sarlogic_0/_343_/CLK 3.47f
C245 DAC_1/carray_0/m2_33700_1156# DAC_1/carray_0/m3_33600_1156# 2.11f
C246 sarlogic_0/_271_/A dvdd 2.81f
C247 DAC_1/carray_0/m2_6000_1156# DAC_1/carray_0/m3_6100_1156# 2.11f
C248 sarlogic_0/_298_/A dvdd 3.4f
C249 DAC_1/carray_0/m3_26900_1156# DAC_1/carray_0/m3_27100_1156# 3.35f
C250 DAC_1/carray_0/m2_16400_1156# DAC_1/carray_0/n5 2.39f
C251 DAC_1/carray_0/m3_8700_1156# DAC_1/carray_0/n7 2.16f
C252 DAC_0/carray_0/n2 DAC_0/carray_0/n1 2.02f
C253 DAC_1/carray_0/m3_16500_1156# DAC_1/carray_0/m3_16700_1156# 3.35f
C254 sarlogic_0/_162_/X dvdd 6.56f
C255 DAC_0/carray_0/m2_11200_1156# DAC_0/carray_0/m3_11300_1156# 2.11f
C256 DAC_0/carray_0/m2_25900_1156# DAC_0/carray_0/m3_25800_1156# 2.11f
C257 DAC_0/carray_0/m3_42500_1156# DAC_0/carray_0/m3_42700_1156# 3.35f
C258 DAC_1/carray_0/m3_7400_1156# DAC_1/carray_0/m3_7600_1156# 3.35f
C259 sarlogic_0/_340_/CLK dvdd 5.49f
C260 DAC_0/carray_0/m2_40200_1156# DAC_0/carray_0/m3_40100_1156# 2.11f
C261 DAC_1/carray_0/m3_18000_1156# DAC_1/carray_0/n7 3.1f
C262 DAC_1/carray_0/m2_13800_1156# DAC_1/carray_0/n7 3.52f
C263 DAC_0/carray_0/m3_33400_1156# DAC_0/carray_0/m3_33600_1156# 3.35f
C264 cal dvdd 5.37f
C265 DAC_0/carray_0/m2_31100_1156# DAC_0/carray_0/m3_31000_1156# 2.11f
C266 DAC_0/out DAC_0/carray_0/n3 6.38f
C267 DAC_0/carray_0/m3_15400_1156# DAC_0/carray_0/n5 4.08f
C268 DAC_1/carray_0/n2 DAC_1/carray_0/n3 20.7f
C269 DAC_0/carray_0/m3_24300_1156# DAC_0/carray_0/m3_24500_1156# 3.35f
C270 DAC_1/carray_0/m3_29500_1156# DAC_1/carray_0/n7 3.1f
C271 comparator_0/trim_0/n3 comparator_0/trim_0/drain 3.41f
C272 DAC_1/carray_0/m2_24600_1156# DAC_1/carray_0/m3_24500_1156# 2.11f
C273 DAC_0/carray_0/m3_13900_1156# DAC_0/carray_0/m3_14100_1156# 3.35f
C274 DAC_1/carray_0/m2_15100_1156# DAC_1/carray_0/m3_15200_1156# 2.11f
C275 DAC_1/carray_0/m3_38800_1156# DAC_1/carray_0/n7 2.16f
C276 DAC_1/carray_0/m3_33400_1156# DAC_1/carray_0/n5 4.08f
C277 DAC_0/carray_0/n3 DAC_0/carray_0/n4 12.1f
C278 sarlogic_0/_217_/A dvdd 2.36f
C279 DAC_0/carray_0/m3_4800_1156# DAC_0/carray_0/m3_5000_1156# 3.35f
C280 sample avdd 13.4f
C281 DAC_1/carray_0/m3_2400_1156# DAC_1/carray_0/n6 4.08f
C282 DAC_0/carray_0/m3_12800_1156# DAC_0/carray_0/n7 4.08f
C283 sample DAC_0/carray_0/n7 4.96f
C284 DAC_0/carray_0/m2_800_1156# DAC_0/carray_0/m3_900_1156# 2.11f
C285 DAC_1/carray_0/n5 DAC_1/carray_0/n6 17.4f
C286 DAC_1/carray_0/n3 DAC_1/carray_0/n1 3.36f
C287 DAC_1/carray_0/m3_32100_1156# DAC_1/carray_0/n6 4.08f
C288 DAC_0/carray_0/m3_42500_1156# DAC_0/carray_0/n7 4.08f
C289 DAC_1/carray_0/m2_15100_1156# DAC_1/carray_0/n7 2.39f
C290 DAC_1/carray_0/m2_20300_1156# DAC_1/carray_0/m3_20400_1156# 2.11f
C291 DAC_0/carray_0/m2_37600_1156# DAC_0/carray_0/n7 2.39f
C292 DAC_1/carray_0/m3_37300_1156# DAC_1/carray_0/m3_37500_1156# 3.35f
C293 avdd DAC_0/sw_top_3/m2_1158_361# 2.15f
C294 DAC_1/carray_0/m3_1100_1156# DAC_1/carray_0/n7 4.08f
C295 ctlp1 ctlp7 3.12f
C296 DAC_1/carray_0/m2_35000_1156# DAC_1/carray_0/m3_34900_1156# 2.11f
C297 DAC_1/carray_0/m2_7300_1156# DAC_1/carray_0/m3_7400_1156# 2.11f
C298 DAC_1/carray_0/m3_30800_1156# DAC_1/carray_0/n7 3.14f
C299 DAC_0/carray_0/m2_19000_1156# DAC_0/carray_0/n7 2.42f
C300 sarlogic_0/clkbuf_0_clk/X dvdd 3.63f
C301 DAC_1/carray_0/m3_28200_1156# DAC_1/carray_0/m3_28400_1156# 3.35f
C302 comparator_0/trim_0/drain comparator_0/trim_0/n4 6.89f
C303 sarlogic_0/input1/X dvdd 3.35f
C304 DAC_1/carray_0/m2_24600_1156# DAC_1/carray_0/n7 2.39f
C305 DAC_0/carray_0/m2_23300_1156# DAC_0/carray_0/n4 2.39f
C306 sarlogic_0/_275_/A dvdd 2.97f
C307 DAC_0/out DAC_0/carray_0/n4 12.2f
C308 DAC_0/carray_0/m3_4800_1156# DAC_0/carray_0/n7 2.16f
C309 DAC_1/carray_0/m3_17800_1156# DAC_1/carray_0/m3_18000_1156# 3.35f
C310 DAC_0/carray_0/m2_12500_1156# DAC_0/carray_0/m3_12600_1156# 2.11f
C311 DAC_0/carray_0/m3_28200_1156# DAC_0/carray_0/n5 4.09f
C312 DAC_1/carray_0/m2_3400_1156# DAC_1/carray_0/n6 2.39f
C313 DAC_0/carray_0/m2_27200_1156# DAC_0/carray_0/m3_27100_1156# 2.11f
C314 DAC_0/carray_0/m2_40200_1156# DAC_0/carray_0/n6 2.39f
C315 DAC_1/carray_0/m3_8700_1156# DAC_1/carray_0/m3_8900_1156# 3.35f
C316 DAC_0/carray_0/m3_14100_1156# DAC_0/carray_0/n7 4.08f
C317 DAC_0/carray_0/m2_41500_1156# DAC_0/carray_0/m3_41400_1156# 2.11f
C318 DAC_0/carray_0/n2 DAC_0/carray_0/m3_20400_1156# 3.43f
C319 DAC_0/carray_0/m2_8600_1156# DAC_0/carray_0/m3_8700_1156# 2.11f
C320 DAC_0/carray_0/m3_26900_1156# DAC_0/carray_0/n6 4.08f
C321 DAC_0/carray_0/m2_9900_1156# DAC_0/carray_0/n7 2.39f
C322 DAC_0/carray_0/m3_19300_1156# DAC_0/carray_0/n4 4.08f
C323 vinp DAC_0/out 21.5f
C324 DAC_0/carray_0/m2_17700_1156# DAC_0/carray_0/m3_17800_1156# 2.11f
C325 DAC_1/carray_0/m2_2100_1156# DAC_1/carray_0/n7 2.39f
C326 DAC_0/carray_0/m3_34700_1156# DAC_0/carray_0/m3_34900_1156# 3.35f
C327 DAC_0/carray_0/m2_38900_1156# DAC_0/carray_0/n7 3.52f
C328 DAC_0/carray_0/m2_32400_1156# DAC_0/carray_0/m3_32300_1156# 2.11f
C329 DAC_0/carray_0/m3_25600_1156# DAC_0/carray_0/n7 4.08f
C330 clk en 2.63f
C331 DAC_0/carray_0/m3_25600_1156# DAC_0/carray_0/m3_25800_1156# 3.35f
C332 DAC_1/carray_0/m2_8600_1156# DAC_1/carray_0/n7 3.52f
C333 sarlogic_0/_248_/A dvdd 4.56f
C334 DAC_0/carray_0/m3_15200_1156# DAC_0/carray_0/m3_15400_1156# 3.35f
C335 DAC_0/carray_0/m3_16700_1156# DAC_0/carray_0/n6 3.14f
C336 sarlogic_0/_339_/Q dvdd 3.02f
C337 DAC_0/carray_0/m2_12500_1156# DAC_0/carray_0/n6 2.39f
C338 DAC_0/carray_0/m2_4700_1156# DAC_0/carray_0/n7 3.52f
C339 DAC_1/carray_0/m2_16400_1156# DAC_1/carray_0/m3_16500_1156# 2.11f
C340 DAC_0/carray_0/m3_6100_1156# DAC_0/carray_0/m3_6300_1156# 3.35f
C341 DAC_0/out DAC_0/carray_0/n5 24.3f
C342 DAC_1/out DAC_1/carray_0/n3 6.38f
C343 DAC_0/carray_0/ndum sample 11.1f
C344 DAC_1/carray_0/m3_38600_1156# DAC_1/carray_0/m3_38800_1156# 3.35f
C345 ctln7 ctln1 3.13f
C346 DAC_1/carray_0/m3_3700_1156# DAC_1/carray_0/n7 4.08f
C347 DAC_1/carray_0/m2_36300_1156# DAC_1/carray_0/m3_36200_1156# 2.11f
C348 DAC_0/carray_0/n4 DAC_0/carray_0/n5 12.7f
C349 DAC_1/carray_0/m3_29500_1156# DAC_1/carray_0/m3_29700_1156# 3.35f
C350 DAC_0/carray_0/m2_23300_1156# DAC_0/carray_0/m3_23200_1156# 2.11f
C351 DAC_1/carray_0/m2_28500_1156# DAC_1/carray_0/n7 2.42f
C352 DAC_1/carray_0/n2 DAC_1/carray_0/m3_23200_1156# 3.4f
C353 DAC_1/carray_0/m3_13900_1156# DAC_1/carray_0/n7 2.16f
C354 DAC_1/carray_0/n6 DAC_1/carray_0/n7 22.1f
C355 DAC_1/carray_0/m3_19100_1156# DAC_1/carray_0/m3_19300_1156# 3.35f
C356 sarlogic_0/_320_/Q dvdd 6.63f
C357 DAC_0/carray_0/m2_13800_1156# DAC_0/carray_0/m3_13900_1156# 2.11f
C358 cal en 2.22f
C359 DAC_1/carray_0/m2_4700_1156# DAC_1/carray_0/m3_4800_1156# 2.11f
C360 sarlogic_0/_273_/A dvdd 5.67f
C361 ctln7 ctln6 2.73f
C362 DAC_1/carray_0/m2_32400_1156# DAC_1/carray_0/n5 2.39f
C363 DAC_1/carray_0/m3_10000_1156# DAC_1/carray_0/m3_10200_1156# 3.35f
C364 DAC_1/carray_0/m3_6300_1156# DAC_1/carray_0/n6 4.08f
C365 DAC_0/carray_0/m2_42800_1156# DAC_0/carray_0/m3_42700_1156# 2.11f
C366 ctln7 dvdd 2.13f
C367 DAC_0/carray_0/m2_19000_1156# DAC_0/carray_0/m3_19100_1156# 2.11f
C368 sarlogic_0/_225_/X dvdd 2.8f
C369 DAC_0/carray_0/m3_36000_1156# DAC_0/carray_0/m3_36200_1156# 3.35f
C370 DAC_1/carray_0/m3_900_1156# DAC_1/carray_0/m3_1100_1156# 3.35f
C371 DAC_0/out DAC_0/carray_0/n6 48.6f
C372 DAC_1/carray_0/m2_31100_1156# DAC_1/carray_0/n6 2.39f
C373 DAC_0/carray_0/m2_41500_1156# DAC_0/carray_0/n7 2.39f
C374 DAC_0/carray_0/m2_33700_1156# DAC_0/carray_0/m3_33600_1156# 2.11f
C375 DAC_1/carray_0/m3_5000_1156# DAC_1/carray_0/n7 4.08f
C376 sarlogic_0/_283_/Y sarlogic_0/_343_/CLK 4.37f
C377 DAC_0/carray_0/m2_6000_1156# DAC_0/carray_0/m3_6100_1156# 2.11f
Xlatch_0 avdd avss latch_0/Qn latch_0/S latch_0/R comp latch
XDAC_0 DAC_0/enb DAC_0/en_buf ctlp1 ctlp0 avdd ctlp3 ctlp4 ctlp5 ctlp6 ctlp7 ctlp2
+ avdd avss sample DAC_0/out vinp DAC
XDAC_1 DAC_1/enb DAC_1/en_buf ctln1 ctln0 avss ctln3 ctln4 ctln5 ctln6 ctln7 ctln2
+ avdd avss sample DAC_1/out vinn DAC
Xcomparator_0 trim3 trim2 trim0 trim1 trim4 trimb4 trimb1 trimb0 trimb2 trimb3 latch_0/R
+ latch_0/S clkc avdd avss DAC_1/out DAC_0/out comparator
Xsarlogic_0 ctln0 ctln1 ctln2 ctln3 ctln4 ctln5 ctln6 ctln7 ctlp0 ctlp1 ctlp2 ctlp3
+ ctlp4 ctlp5 ctlp6 ctlp7 cal clk clkc comp en result0 result1 result2 result3 result4
+ result5 result6 result7 rstn sample trim0 trim1 trim2 trim3 trim4 trimb0 trimb1
+ trimb2 trimb3 trimb4 valid dvdd avss sarlogic
C378 sarlogic_0/_286_/Y avss 4.3f
C379 dvdd avss 5.48p
C380 sarlogic_0/_284_/A avss 2.54f
C381 sarlogic_0/_147_/Y avss 3.97f
C382 sarlogic_0/_190_/A avss 2.2f
C383 sarlogic_0/_333_/Q avss 2.02f
C384 sarlogic_0/_328_/Q avss 3.67f
C385 sarlogic_0/_212_/X avss 3.15f
C386 sarlogic_0/_327_/Q avss 2.34f
C387 sarlogic_0/_207_/C avss 3.47f
C388 sarlogic_0/_254_/B avss 5.11f
C389 sarlogic_0/_304_/X avss 2.93f
C390 sarlogic_0/_147_/A avss 6.15f
C391 sarlogic_0/_192_/B avss 3.21f
C392 sarlogic_0/_267_/A avss 3.45f
C393 sarlogic_0/_228_/A avss 3.19f
C394 sarlogic_0/_297_/B avss 3.05f
C395 sarlogic_0/_248_/A avss 2.92f
C396 sarlogic_0/_315_/D avss 3.89f
C397 sarlogic_0/_340_/CLK avss 4.88f
C398 sarlogic_0/_281_/A avss 2.48f
C399 sarlogic_0/_331_/CLK avss 4.41f
C400 sarlogic_0/_306_/S avss 4.04f
C401 sarlogic_0/_340_/Q avss 2.1f
C402 sarlogic_0/_343_/CLK avss 3.82f
C403 sarlogic_0/_283_/A avss 5.42f
C404 sarlogic_0/_346_/SET_B avss 13.8f
C405 sarlogic_0/_197_/X avss 2.47f
C406 rstn avss 4.06f
C407 sarlogic_0/_227_/A avss 5.07f
C408 sarlogic_0/_161_/Y avss 2.08f
C409 sarlogic_0/_242_/A avss 3f
C410 sarlogic_0/_304_/S avss 2.49f
C411 sarlogic_0/_215_/A avss 2.2f
C412 sarlogic_0/_232_/X avss 2.7f
C413 sarlogic_0/_216_/A avss 2.36f
C414 result7 avss 3.01f
C415 sarlogic_0/_181_/X avss 2.07f
C416 sarlogic_0/_196_/A avss 4.84f
C417 sarlogic_0/_286_/B avss 3.17f
C418 sarlogic_0/_330_/Q avss 2.6f
C419 sarlogic_0/_321_/Q avss 2.62f
C420 sarlogic_0/_324_/Q avss 2.79f
C421 sarlogic_0/_157_/A avss 2.21f
C422 sarlogic_0/clkbuf_0_clk/X avss 2.8f
C423 clk avss 2.71f
C424 sarlogic_0/clkbuf_0_clk/a_110_7# avss 2.34f **FLOATING
C425 sarlogic_0/_325_/Q avss 3.5f
C426 sarlogic_0/_329_/Q avss 2.08f
C427 sarlogic_0/_254_/A avss 2.28f
C428 sarlogic_0/_172_/A avss 3.15f
C429 sarlogic_0/repeater43/X avss 15.7f
C430 sarlogic_0/_273_/A avss 2.25f
C431 sarlogic_0/_316_/Q avss 2.05f
C432 sarlogic_0/_258_/S avss 3.05f
C433 sarlogic_0/_285_/A avss 2.14f
C434 sarlogic_0/_294_/A avss 3.28f
C435 clkc avss 5.93f
C436 latch_0/R avss 3.17f
C437 comparator_0/comparator_core_0/w_302_2337# avss 4.58f **FLOATING
C438 latch_0/S avss 3.34f
C439 comparator_0/trim_1/drain avss 4.12f
C440 comparator_0/trim_1/n3 avss 2.65f
C441 trimb3 avss 3.92f
C442 comparator_0/trim_1/n4 avss 4.07f
C443 trimb4 avss 4f
C444 comparator_0/trim_0/drain avss 4.09f
C445 comparator_0/trim_0/n3 avss 2.65f
C446 trim3 avss 3.65f
C447 comparator_0/trim_0/n4 avss 4.07f
C448 trim4 avss 4.06f
C449 ctln7 avss 2.07f
C450 ctln2 avss 2.07f
C451 DAC_1/sw_top_3/m2_990_200# avss 2.32f **FLOATING
C452 DAC_1/sw_top_3/m2_1158_361# avss 2.14f
C453 DAC_1/en_buf avss 4.5f
C454 DAC_1/enb avss 4.07f
C455 DAC_1/carray_0/n1 avss 4.16f
C456 DAC_1/carray_0/n7 avss 65.7f
C457 DAC_1/carray_0/n6 avss 32.3f
C458 DAC_1/carray_0/n5 avss 17.4f
C459 DAC_1/carray_0/n4 avss 8.63f
C460 DAC_1/carray_0/n3 avss 6.31f
C461 DAC_1/carray_0/m2_42800_1156# avss 2.03f
C462 DAC_1/carray_0/m2_800_1156# avss 2.03f
C463 DAC_1/carray_0/n0 avss 3.21f
C464 DAC_1/carray_0/n2 avss 8.22f
C465 DAC_1/out avss 35.8f
C466 DAC_1/carray_0/ndum avss 6.89f
C467 sample avss 64.6f
C468 DAC_1/sw_top_0/m2_990_200# avss 2.32f **FLOATING
C469 vinn avss 7.69f
C470 DAC_1/sw_top_0/m2_1158_361# avss 2.14f
C471 avdd avss 12.3p
C472 ctln0 avss 2.58f
C473 ctln6 avss 2.33f
C474 ctlp7 avss 2.49f
C475 ctlp2 avss 2.28f
C476 DAC_0/sw_top_3/m2_990_200# avss 2.32f **FLOATING
C477 DAC_0/sw_top_3/m2_1158_361# avss 2.14f
C478 DAC_0/en_buf avss 4.5f
C479 DAC_0/enb avss 4.07f
C480 DAC_0/carray_0/n1 avss 4.16f
C481 DAC_0/carray_0/n7 avss 65.7f
C482 DAC_0/carray_0/n6 avss 32.3f
C483 DAC_0/carray_0/n5 avss 17.4f
C484 DAC_0/carray_0/n4 avss 8.63f
C485 DAC_0/carray_0/n3 avss 6.31f
C486 DAC_0/carray_0/m2_42800_1156# avss 2.03f
C487 DAC_0/carray_0/m2_800_1156# avss 2.03f
C488 DAC_0/carray_0/n0 avss 3.19f
C489 DAC_0/carray_0/n2 avss 8.22f
C490 DAC_0/out avss 35.8f
C491 DAC_0/carray_0/ndum avss 6.77f
C492 ctlp4 avss 2.34f
C493 DAC_0/sw_top_0/m2_990_200# avss 2.32f **FLOATING
C494 vinp avss 7.69f
C495 DAC_0/sw_top_0/m2_1158_361# avss 2.14f
C496 ctlp5 avss 2.55f
C497 ctlp1 avss 2.75f
C498 ctlp0 avss 3.52f
C499 ctlp6 avss 2.28f
C500 comp avss 3.03f
.ends
