** sch_path: /home/alex/Desktop/SAR_IPN/xschem/tb/sar/tr_sar.sch

.include /home/alex/pdk/sky130B/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
*.include /home/alex/pdk/sky130B/libs.ref/sky130_fd_sc_hd/spice/cells/inv/sky130_fd_sc_hd__inv_4.spice
*.include /home/alex/pdk/sky130B/libs.ref/sky130_fd_sc_hd/spice/cells/decap/sky130_fd_sc_hd__decap_8.spice
*.include /home/alex/pdk/sky130B/libs.ref/sky130_fd_sc_hd/spice/cells/decap/sky130_fd_sc_hd__decap_3.spice
*.include /home/alex/pdk/sky130B/libs.ref/sky130_fd_sc_hd/spice/cells/buf/sky130_fd_sc_hd__buf_1.spice
*.include /home/alex/pdk/sky130B/libs.ref/sky130_fd_sc_hd/spice/cells/inv/sky130_fd_sc_hd__inv_1.spice
*.include /home/alex/pdk/sky130B/libs.ref/sky130_fd_sc_hd/spice/cells/inv/sky130_fd_sc_hd__inv_2.spice
*.include /home/alex/pdk/sky130B/libs.ref/sky130_fd_sc_hd/spice/cells/tap/sky130_fd_sc_hd__tap_2.spice


.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/alex/pdk/sky130B/libs.tech/ngspice/corners/tt.spice
.include /home/alex/pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/alex/pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/alex/pdk/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice

**.subckt tr_sar
V1 vss GND 0
.save i(v1)
V2 vdd GND 1.4
.save i(v2)
V4 vinn GND vsign
.save i(v4)
V5 vinp GND vsigp
.save i(v5)
Vclk clk GND PULSE(0 1 1e-9 1e-9 1e-9 2e-6 4e-6)
.save i(vclk)
Ven en GND 1.4
.save i(ven)
V3 cal GND 0
.save i(v3)
xsar vdd vdd vss result_7_ result_6_ result_5_ result_4_ result_3_ result_2_ result_1_ result_0_
+ vinn vss clk vinp en valid cal rstn sar
V7 rstn GND PWL(0 0 4e-6 0 4.001e-6 1.4)
.save i(v7)
**.ends

* expanding   symbol:  sar/sar/sar.sym # of pins=12
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/sar/sar.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/sar/sar.sch
.subckt sar avdd dvdd dvss result_7_ result_6_ result_5_ result_4_ result_3_ result_2_ result_1_
+ result_0_ vinn avss clk vinp en valid cal rstn
*.iopin avss
*.iopin avdd
*.iopin dvss
*.iopin dvdd
*.ipin vinp
*.ipin vinn
*.opin result_7_,result_6_,result_5_,result_4_,result_3_,result_2_,result_1_,result_0_
*.ipin clk
*.ipin en
*.opin valid
*.ipin cal
*.ipin rstn
xlat avdd comp net1 avss outn outp latch
**** begin user architecture code

.include /home/alex/Desktop/SAR_IPN/xschem/sar/control/cmos_cells_digital.sp
.include /home/alex/Desktop/SAR_IPN/xschem/sar/control/sar_logic.sp

**** end user architecture code
xdn vn sample avdd avss vinn ctln_7_ ctln_6_ ctln_5_ ctln_4_ ctln_3_ ctln_2_ ctln_1_ ctln_0_ avss
+ dac
xdp vp sample avdd avss vinp ctlp_7_ ctlp_6_ ctlp_5_ ctlp_4_ ctlp_3_ ctlp_2_ ctlp_1_ ctlp_0_ avdd
+ dac
xcom avss avdd clkc outp vp outn vn trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ trimb_4_ trimb_3_
+ trimb_2_ trimb_1_ trimb_0_ comparator
**** begin user architecture code


Xuut dclk drstn den dcomp dcal dvalid dres0 dres1 dres2 dres3 dres4 dres5 dres6 dres7 dsamp dctlp0
+ dctlp1 dctlp2 dctlp3 dctlp4 dctlp5 dctlp6 dctlp7 dctln0 dctln1 dctln2 dctln3 dctln4 dctln5 dctln6 dctln7
+ dtrim0 dtrim1 dtrim2 dtrim3 dtrim4 dtrimb0 dtrimb1 dtrimb2 dtrimb3 dtrimb4 dclkc sar_logic

.model adc_buff adc_bridge(in_low = 0.2 in_high=0.8)
.model dac_buff dac_bridge(out_high = 1.2)

Aad [clk rstn en comp cal] [dclk drstn den dcomp dcal] adc_buff
Ada [dctlp0 dctlp1 dctlp2 dctlp3 dctlp4 dctlp5 dctlp6 dctlp7 dctln0 dctln1 dctln2 dctln3 dctln4
+ dctln5 dctln6 dctln7 dres0 dres1 dres2 dres3 dres4 dres5 dres6 dres7 dsamp dclkc] [ctlp_0_ ctlp_1_ ctlp_2_
+ ctlp_3_ ctlp_4_ ctlp_5_ ctlp_6_ ctlp_7_ ctln_0_ ctln_1_ ctln_2_ ctln_3_ ctln_4_ ctln_5_ ctln_6_ ctln_7_
+ res0 res1 res2 res3 res4 res5 res6 res7 sample clkc] dac_buff
Ada2 [dtrim4 dtrim3 dtrim2 dtrim1 dtrim0 dtrimb4 dtrimb3 dtrimb2 dtrimb1 dtrimb0] [trim_4_ trim_3_
+ trim_2_ trim_1_ trim_0_ trimb_4_ trimb_3_ trimb_2_ trimb_1_ trimb_0_ ] dac_buff



**** end user architecture code
.ends


* expanding   symbol:  sar/latch/latch.sym # of pins=6
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/latch/latch.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/latch/latch.sch
.subckt latch vdd Q Qn vss R S
*.ipin S
*.ipin R
*.iopin vss
*.iopin vdd
*.opin Q
*.opin Qn
x1 vdd Qn Q vss inv_lvt
x2 vdd Q Qn vss inv_lvt
x3 vdd R net2 vss inv_lvt
x4 vdd S net1 vss inv_lvt
XM4 Q net2 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 Qn net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sar/dac/dac.sym # of pins=7
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/dac/dac.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/dac/dac.sch
.subckt dac out sample vdd vss vin ctl_7_ ctl_6_ ctl_5_ ctl_4_ ctl_3_ ctl_2_ ctl_1_ ctl_0_ dum
*.ipin vin
*.ipin sample
*.opin out
*.ipin ctl_7_,ctl_6_,ctl_5_,ctl_4_,ctl_3_,ctl_2_,ctl_1_,ctl_0_
*.ipin dum
*.iopin vdd
*.iopin vss
xca out n6 n0 n5 n4 n2 ndum n3 n1 n7 carray
xi6 ctl_6_ vss vss vdd vdd n6 sky130_fd_sc_hd__inv_2
xi5 ctl_5_ vss vss vdd vdd n5 sky130_fd_sc_hd__inv_2
xi4 ctl_4_ vss vss vdd vdd n4 sky130_fd_sc_hd__inv_2
xi3 ctl_3_ vss vss vdd vdd n3 sky130_fd_sc_hd__inv_2
xi2 ctl_2_ vss vss vdd vdd n2 sky130_fd_sc_hd__inv_2
xi1 ctl_1_ vss vss vdd vdd n1 sky130_fd_sc_hd__inv_2
xi0 ctl_0_ vss vss vdd vdd n0 sky130_fd_sc_hd__inv_2
xidum dum vss vss vdd vdd ndum sky130_fd_sc_hd__inv_2
xi7 ctl_7_ vss vss vdd vdd n7 sky130_fd_sc_hd__inv_2
xswt out sample vdd vin vss sw_top
.ends


* expanding   symbol:  sar/comparator/comparator.sym # of pins=9
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/comparator.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/comparator.sch
.subckt comparator vss vdd clk outp vp outn vn trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ trimb_4_
+ trimb_3_ trimb_2_ trimb_1_ trimb_0_
*.ipin vn
*.ipin vp
*.ipin clk
*.iopin vdd
*.iopin vss
*.opin outp
*.opin outn
*.ipin trim_4_,trim_3_,trim_2_,trim_1_,trim_0_
*.ipin trimb_4_,trimb_3_,trimb_2_,trimb_1_,trimb_0_
x2 in trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ vss trim
x3 ip trimb_4_ trimb_3_ trimb_2_ trimb_1_ trimb_0_ vss trim
XM1 in clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 outn clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 outn outp vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMl4 outp outn vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 outp clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 ip clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMl2 outp outn ip vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMl1 outn outp in vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMinn in vn diff vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMinp ip vp diff vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMdiff diff clk vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  logic/inv_lvt.sym # of pins=4
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/logic/inv_lvt.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/logic/inv_lvt.sch
.subckt inv_lvt vdd in out vss
*.iopin vdd
*.iopin vss
*.ipin in
*.opin out
XM3 out in vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 out in vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sar/dac/carray.sym # of pins=10
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/dac/carray.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/dac/carray.sch
.subckt carray top n6 n0 n5 n4 n2 ndum n3 n1 n7
*.iopin top
*.iopin n7
*.iopin n6
*.iopin n5
*.iopin n4
*.iopin n2
*.iopin n0
*.iopin ndum
*.iopin n3
*.iopin n1
xcdum top ndum unitcap
xc0 top n0 unitcap
xc1_1_ top n1 unitcap
xc1_0_ top n1 unitcap
xc2_3_ top n2 unitcap
xc2_2_ top n2 unitcap
xc2_1_ top n2 unitcap
xc2_0_ top n2 unitcap
xc3_7_ top n3 unitcap
xc3_6_ top n3 unitcap
xc3_5_ top n3 unitcap
xc3_4_ top n3 unitcap
xc3_3_ top n3 unitcap
xc3_2_ top n3 unitcap
xc3_1_ top n3 unitcap
xc3_0_ top n3 unitcap
xc4_15_ top n4 unitcap
xc4_14_ top n4 unitcap
xc4_13_ top n4 unitcap
xc4_12_ top n4 unitcap
xc4_11_ top n4 unitcap
xc4_10_ top n4 unitcap
xc4_9_ top n4 unitcap
xc4_8_ top n4 unitcap
xc4_7_ top n4 unitcap
xc4_6_ top n4 unitcap
xc4_5_ top n4 unitcap
xc4_4_ top n4 unitcap
xc4_3_ top n4 unitcap
xc4_2_ top n4 unitcap
xc4_1_ top n4 unitcap
xc4_0_ top n4 unitcap
xc5_31_ top n5 unitcap
xc5_30_ top n5 unitcap
xc5_29_ top n5 unitcap
xc5_28_ top n5 unitcap
xc5_27_ top n5 unitcap
xc5_26_ top n5 unitcap
xc5_25_ top n5 unitcap
xc5_24_ top n5 unitcap
xc5_23_ top n5 unitcap
xc5_22_ top n5 unitcap
xc5_21_ top n5 unitcap
xc5_20_ top n5 unitcap
xc5_19_ top n5 unitcap
xc5_18_ top n5 unitcap
xc5_17_ top n5 unitcap
xc5_16_ top n5 unitcap
xc5_15_ top n5 unitcap
xc5_14_ top n5 unitcap
xc5_13_ top n5 unitcap
xc5_12_ top n5 unitcap
xc5_11_ top n5 unitcap
xc5_10_ top n5 unitcap
xc5_9_ top n5 unitcap
xc5_8_ top n5 unitcap
xc5_7_ top n5 unitcap
xc5_6_ top n5 unitcap
xc5_5_ top n5 unitcap
xc5_4_ top n5 unitcap
xc5_3_ top n5 unitcap
xc5_2_ top n5 unitcap
xc5_1_ top n5 unitcap
xc5_0_ top n5 unitcap
xc6_63_ top n6 unitcap
xc6_62_ top n6 unitcap
xc6_61_ top n6 unitcap
xc6_60_ top n6 unitcap
xc6_59_ top n6 unitcap
xc6_58_ top n6 unitcap
xc6_57_ top n6 unitcap
xc6_56_ top n6 unitcap
xc6_55_ top n6 unitcap
xc6_54_ top n6 unitcap
xc6_53_ top n6 unitcap
xc6_52_ top n6 unitcap
xc6_51_ top n6 unitcap
xc6_50_ top n6 unitcap
xc6_49_ top n6 unitcap
xc6_48_ top n6 unitcap
xc6_47_ top n6 unitcap
xc6_46_ top n6 unitcap
xc6_45_ top n6 unitcap
xc6_44_ top n6 unitcap
xc6_43_ top n6 unitcap
xc6_42_ top n6 unitcap
xc6_41_ top n6 unitcap
xc6_40_ top n6 unitcap
xc6_39_ top n6 unitcap
xc6_38_ top n6 unitcap
xc6_37_ top n6 unitcap
xc6_36_ top n6 unitcap
xc6_35_ top n6 unitcap
xc6_34_ top n6 unitcap
xc6_33_ top n6 unitcap
xc6_32_ top n6 unitcap
xc6_31_ top n6 unitcap
xc6_30_ top n6 unitcap
xc6_29_ top n6 unitcap
xc6_28_ top n6 unitcap
xc6_27_ top n6 unitcap
xc6_26_ top n6 unitcap
xc6_25_ top n6 unitcap
xc6_24_ top n6 unitcap
xc6_23_ top n6 unitcap
xc6_22_ top n6 unitcap
xc6_21_ top n6 unitcap
xc6_20_ top n6 unitcap
xc6_19_ top n6 unitcap
xc6_18_ top n6 unitcap
xc6_17_ top n6 unitcap
xc6_16_ top n6 unitcap
xc6_15_ top n6 unitcap
xc6_14_ top n6 unitcap
xc6_13_ top n6 unitcap
xc6_12_ top n6 unitcap
xc6_11_ top n6 unitcap
xc6_10_ top n6 unitcap
xc6_9_ top n6 unitcap
xc6_8_ top n6 unitcap
xc6_7_ top n6 unitcap
xc6_6_ top n6 unitcap
xc6_5_ top n6 unitcap
xc6_4_ top n6 unitcap
xc6_3_ top n6 unitcap
xc6_2_ top n6 unitcap
xc6_1_ top n6 unitcap
xc6_0_ top n6 unitcap
xc7_127_ top n7 unitcap
xc7_126_ top n7 unitcap
xc7_125_ top n7 unitcap
xc7_124_ top n7 unitcap
xc7_123_ top n7 unitcap
xc7_122_ top n7 unitcap
xc7_121_ top n7 unitcap
xc7_120_ top n7 unitcap
xc7_119_ top n7 unitcap
xc7_118_ top n7 unitcap
xc7_117_ top n7 unitcap
xc7_116_ top n7 unitcap
xc7_115_ top n7 unitcap
xc7_114_ top n7 unitcap
xc7_113_ top n7 unitcap
xc7_112_ top n7 unitcap
xc7_111_ top n7 unitcap
xc7_110_ top n7 unitcap
xc7_109_ top n7 unitcap
xc7_108_ top n7 unitcap
xc7_107_ top n7 unitcap
xc7_106_ top n7 unitcap
xc7_105_ top n7 unitcap
xc7_104_ top n7 unitcap
xc7_103_ top n7 unitcap
xc7_102_ top n7 unitcap
xc7_101_ top n7 unitcap
xc7_100_ top n7 unitcap
xc7_99_ top n7 unitcap
xc7_98_ top n7 unitcap
xc7_97_ top n7 unitcap
xc7_96_ top n7 unitcap
xc7_95_ top n7 unitcap
xc7_94_ top n7 unitcap
xc7_93_ top n7 unitcap
xc7_92_ top n7 unitcap
xc7_91_ top n7 unitcap
xc7_90_ top n7 unitcap
xc7_89_ top n7 unitcap
xc7_88_ top n7 unitcap
xc7_87_ top n7 unitcap
xc7_86_ top n7 unitcap
xc7_85_ top n7 unitcap
xc7_84_ top n7 unitcap
xc7_83_ top n7 unitcap
xc7_82_ top n7 unitcap
xc7_81_ top n7 unitcap
xc7_80_ top n7 unitcap
xc7_79_ top n7 unitcap
xc7_78_ top n7 unitcap
xc7_77_ top n7 unitcap
xc7_76_ top n7 unitcap
xc7_75_ top n7 unitcap
xc7_74_ top n7 unitcap
xc7_73_ top n7 unitcap
xc7_72_ top n7 unitcap
xc7_71_ top n7 unitcap
xc7_70_ top n7 unitcap
xc7_69_ top n7 unitcap
xc7_68_ top n7 unitcap
xc7_67_ top n7 unitcap
xc7_66_ top n7 unitcap
xc7_65_ top n7 unitcap
xc7_64_ top n7 unitcap
xc7_63_ top n7 unitcap
xc7_62_ top n7 unitcap
xc7_61_ top n7 unitcap
xc7_60_ top n7 unitcap
xc7_59_ top n7 unitcap
xc7_58_ top n7 unitcap
xc7_57_ top n7 unitcap
xc7_56_ top n7 unitcap
xc7_55_ top n7 unitcap
xc7_54_ top n7 unitcap
xc7_53_ top n7 unitcap
xc7_52_ top n7 unitcap
xc7_51_ top n7 unitcap
xc7_50_ top n7 unitcap
xc7_49_ top n7 unitcap
xc7_48_ top n7 unitcap
xc7_47_ top n7 unitcap
xc7_46_ top n7 unitcap
xc7_45_ top n7 unitcap
xc7_44_ top n7 unitcap
xc7_43_ top n7 unitcap
xc7_42_ top n7 unitcap
xc7_41_ top n7 unitcap
xc7_40_ top n7 unitcap
xc7_39_ top n7 unitcap
xc7_38_ top n7 unitcap
xc7_37_ top n7 unitcap
xc7_36_ top n7 unitcap
xc7_35_ top n7 unitcap
xc7_34_ top n7 unitcap
xc7_33_ top n7 unitcap
xc7_32_ top n7 unitcap
xc7_31_ top n7 unitcap
xc7_30_ top n7 unitcap
xc7_29_ top n7 unitcap
xc7_28_ top n7 unitcap
xc7_27_ top n7 unitcap
xc7_26_ top n7 unitcap
xc7_25_ top n7 unitcap
xc7_24_ top n7 unitcap
xc7_23_ top n7 unitcap
xc7_22_ top n7 unitcap
xc7_21_ top n7 unitcap
xc7_20_ top n7 unitcap
xc7_19_ top n7 unitcap
xc7_18_ top n7 unitcap
xc7_17_ top n7 unitcap
xc7_16_ top n7 unitcap
xc7_15_ top n7 unitcap
xc7_14_ top n7 unitcap
xc7_13_ top n7 unitcap
xc7_12_ top n7 unitcap
xc7_11_ top n7 unitcap
xc7_10_ top n7 unitcap
xc7_9_ top n7 unitcap
xc7_8_ top n7 unitcap
xc7_7_ top n7 unitcap
xc7_6_ top n7 unitcap
xc7_5_ top n7 unitcap
xc7_4_ top n7 unitcap
xc7_3_ top n7 unitcap
xc7_2_ top n7 unitcap
xc7_1_ top n7 unitcap
xc7_0_ top n7 unitcap
.ends


* expanding   symbol:  sar/sw/sw_top.sym # of pins=5
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/sw/sw_top.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/sw/sw_top.sch
.subckt sw_top out en vdd in vss
*.iopin out
*.ipin en
*.iopin vss
*.iopin vdd
*.iopin in
x2 vss vss vdd vdd sky130_fd_sc_hd__decap_8
x4 en vss vss vdd vdd en_buf sky130_fd_sc_hd__inv_4
x1 VGND VNB VPB VPWR sky130_fd_sc_hd__decap_3
XM1 in en out vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM2 in en_buf out vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
.ends


* expanding   symbol:  sar/comparator/trim.sym # of pins=3
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/trim.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/trim.sch
.subckt trim drain d_4_ d_3_ d_2_ d_1_ d_0_ vss
*.iopin vss
*.ipin d_4_,d_3_,d_2_,d_1_,d_0_
*.opin drain
x4_7_ drain n4 trimcap
x4_6_ drain n4 trimcap
x4_5_ drain n4 trimcap
x4_4_ drain n4 trimcap
x4_3_ drain n4 trimcap
x4_2_ drain n4 trimcap
x4_1_ drain n4 trimcap
x4_0_ drain n4 trimcap
x3_3_ drain n3 trimcap
x3_2_ drain n3 trimcap
x3_1_ drain n3 trimcap
x3_0_ drain n3 trimcap
x2_1_ drain n2 trimcap
x2_0_ drain n2 trimcap
x1 drain n1 trimcap
x0 drain n0 trimcap
XM4_7_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_6_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_5_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_4_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_3_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_2_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_1_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_0_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3_3_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3_2_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3_1_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3_0_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2_1_ n2 d_2_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2_0_ n2 d_2_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 n1 d_1_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 n0 d_0_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sar/unitcap/unitcap.sym # of pins=2
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/unitcap/unitcap.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/unitcap/unitcap.sch
.subckt unitcap cp cn
*.iopin cp
*.iopin cn
XC2 cp cn sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=1 m=1
.ends


* expanding   symbol:  sar/comparator/trimcap.sym # of pins=2
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/trimcap.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/trimcap.sch
.subckt trimcap cp cn
*.iopin cp
*.iopin cn
C1 cp cn 2f m=1
.ends

.GLOBAL GND
**** begin user architecture code

.options method trap
*.options method gear
.options gmin 1e-15
.options abstol 1e-15
.options reltol 0.0001
.options vntol 0.1e-6
.options warn 1

.param MC_SWITCH=0
.param vin=0.1
.param vcm=0.7
.param vsigp={vcm + vin/2}
.param vsign={vcm - vin/2}

.tran 100e-9 48e-6
.save all
.control

run
write tr_sar.raw
meas tran d0 find v(xsar.res0) at=47e-6
meas tran d1 find v(xsar.res1) at=47e-6
meas tran d2 find v(xsar.res2) at=47e-6
meas tran d3 find v(xsar.res3) at=47e-6
meas tran d4 find v(xsar.res4) at=47e-6
meas tran d5 find v(xsar.res5) at=47e-6
meas tran d6 find v(xsar.res6) at=47e-6
meas tran d7 find v(xsar.res7) at=47e-6

* meas tran d0 find v(xsar.result0) at=47e-6
* meas tran d1 find v(xsar.result1) at=47e-6
* meas tran d2 find v(xsar.result2) at=47e-6
* meas tran d3 find v(xsar.result3) at=47e-6
* meas tran d4 find v(xsar.result4) at=47e-6
* meas tran d5 find v(xsar.result5) at=47e-6
* meas tran d6 find v(xsar.result6) at=47e-6
* meas tran d7 find v(xsar.result7) at=47e-6

meas tran vpmax max xsar.vp
meas tran vpmin min xsar.vp
meas tran vpend find v(xsar.vp) at=39e-6

meas tran vnmax max xsar.vn
meas tran vnmin min xsar.vn
meas tran vnend find v(xsar.vn) at=39e-6

print d0
print d1
print d2
print d3
print d4
print d5
print d6
print d7

print vpmax
print vpmin

print vnmax
print vnmin

print vpend
print vnend

.endc


**** end user architecture code
.end
