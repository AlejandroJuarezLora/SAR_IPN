magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_p >>
rect 6 214 40 248
rect 6 142 40 176
rect 6 70 40 104
rect 6 -2 40 32
<< viali >>
rect 6 214 40 248
rect 6 142 40 176
rect 6 70 40 104
rect 6 -2 40 32
<< metal1 >>
rect 0 248 46 295
rect 0 214 6 248
rect 40 214 46 248
rect 0 176 46 214
rect 0 142 6 176
rect 40 142 46 176
rect 0 104 46 142
rect 0 70 6 104
rect 40 70 46 104
rect 0 32 46 70
rect 0 -2 6 32
rect 40 -2 46 32
rect 0 -40 46 -2
<< properties >>
string path 0.575 6.800 0.575 -0.425 
<< end >>
