magic
tech sky130B
magscale 1 2
timestamp 1696623031
<< pwell >>
rect -285 -279 285 279
<< nmoslvt >>
rect -89 -131 -29 69
rect 29 -131 89 69
<< ndiff >>
rect -147 39 -89 69
rect -147 -101 -135 39
rect -101 -101 -89 39
rect -147 -131 -89 -101
rect -29 39 29 69
rect -29 -101 -17 39
rect 17 -101 29 39
rect -29 -131 29 -101
rect 89 39 147 69
rect 89 -101 101 39
rect 135 -101 147 39
rect 89 -131 147 -101
<< ndiffc >>
rect -135 -101 -101 39
rect -17 -101 17 39
rect 101 -101 135 39
<< psubdiff >>
rect -249 209 249 243
rect -249 -209 -215 209
rect 215 -209 249 209
rect -249 -243 -122 -209
rect 122 -243 249 -209
<< psubdiffcont >>
rect -122 -243 122 -209
<< poly >>
rect -92 141 -26 157
rect -92 107 -76 141
rect -42 107 -26 141
rect -92 91 -26 107
rect 26 141 92 157
rect 26 107 42 141
rect 76 107 92 141
rect 26 91 92 107
rect -89 69 -29 91
rect 29 69 89 91
rect -89 -157 -29 -131
rect 29 -157 89 -131
<< polycont >>
rect -76 107 -42 141
rect 42 107 76 141
<< locali >>
rect -92 107 -76 141
rect -42 107 -26 141
rect 26 107 42 141
rect 76 107 92 141
rect -135 39 -101 55
rect -135 -117 -101 -101
rect -17 39 17 55
rect -17 -117 17 -101
rect 101 39 135 55
rect 101 -117 135 -101
rect -138 -243 -122 -209
rect 122 -243 138 -209
<< viali >>
rect -76 107 -42 141
rect 42 107 76 141
rect -135 -101 -101 39
rect -17 -84 17 22
rect 101 -101 135 39
<< metal1 >>
rect -90 141 -29 154
rect -90 107 -76 141
rect -42 107 -29 141
rect -90 94 -29 107
rect 28 141 89 155
rect 28 107 42 141
rect 76 107 89 141
rect 28 95 89 107
rect -141 39 -95 51
rect -141 -101 -135 39
rect -101 -101 -95 39
rect 95 39 141 51
rect -23 22 23 34
rect -23 -84 -17 22
rect 17 -84 23 22
rect -23 -96 23 -84
rect -141 -113 -95 -101
rect 95 -101 101 39
rect 135 -101 141 39
rect 95 -113 141 -101
<< properties >>
string FIXED_BBOX -232 -226 232 226
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1 l 0.3 m 1 nf 2 diffcov 80 polycov 80 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 80 rlcov 80 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 60 viadrn 80 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
