magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_p >>
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect -29 -187 29 -181
<< pwell >>
rect -114 -135 114 117
<< nmoslvt >>
rect -30 -109 30 91
<< ndiff >>
rect -88 76 -30 91
rect -88 42 -76 76
rect -42 42 -30 76
rect -88 8 -30 42
rect -88 -26 -76 8
rect -42 -26 -30 8
rect -88 -60 -30 -26
rect -88 -94 -76 -60
rect -42 -94 -30 -60
rect -88 -109 -30 -94
rect 30 76 88 91
rect 30 42 42 76
rect 76 42 88 76
rect 30 8 88 42
rect 30 -26 42 8
rect 76 -26 88 8
rect 30 -60 88 -26
rect 30 -94 42 -60
rect 76 -94 88 -60
rect 30 -109 88 -94
<< ndiffc >>
rect -76 42 -42 76
rect -76 -26 -42 8
rect -76 -94 -42 -60
rect 42 42 76 76
rect 42 -26 76 8
rect 42 -94 76 -60
<< poly >>
rect -30 91 30 117
rect -30 -131 30 -109
rect -33 -147 33 -131
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -197 33 -181
<< polycont >>
rect -17 -181 17 -147
<< locali >>
rect -76 76 -42 95
rect -76 8 -42 10
rect -76 -28 -42 -26
rect -76 -113 -42 -94
rect 42 76 76 95
rect 42 8 76 10
rect 42 -28 76 -26
rect 42 -113 76 -94
rect -33 -181 -17 -147
rect 17 -181 33 -147
<< viali >>
rect -76 42 -42 44
rect -76 10 -42 42
rect -76 -60 -42 -28
rect -76 -62 -42 -60
rect 42 42 76 44
rect 42 10 76 42
rect 42 -60 76 -28
rect 42 -62 76 -60
rect -17 -181 17 -147
<< metal1 >>
rect -82 44 -36 91
rect -82 10 -76 44
rect -42 10 -36 44
rect -82 -28 -36 10
rect -82 -62 -76 -28
rect -42 -62 -36 -28
rect -82 -109 -36 -62
rect 36 44 82 91
rect 36 10 42 44
rect 76 10 82 44
rect 36 -28 82 10
rect 36 -62 42 -28
rect 76 -62 82 -28
rect 36 -109 82 -62
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect 17 -181 29 -147
rect -29 -187 29 -181
<< end >>
