magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_s >>
rect 3962 3476 6134 3562
rect 3962 2972 4048 3476
rect 6048 2972 6134 3476
rect 3962 2886 6134 2972
<< metal1 >>
rect 3350 1365 3909 1411
rect 6195 1365 6754 1411
rect 5022 448 5082 559
rect 3512 388 5082 448
rect 3512 -40 3572 388
<< metal2 >>
rect 140 2907 690 2967
rect 9414 2907 9964 2967
rect 140 -40 200 2907
rect 260 2362 690 2422
rect 9414 2362 9844 2422
rect 260 -40 320 2362
rect 380 2086 690 2146
rect 9414 2086 9724 2146
rect 380 -40 440 2086
rect 500 1784 690 1844
rect 9414 1784 9604 1844
rect 500 -40 560 1784
rect 620 1154 768 1214
rect 9336 1154 9484 1214
rect 620 -40 680 1154
rect 1249 34 1309 624
rect 4555 -40 4635 579
rect 5012 34 5092 579
rect 5469 -40 5549 579
rect 8795 34 8855 624
rect 9424 -40 9484 1154
rect 9544 -40 9604 1784
rect 9664 -40 9724 2086
rect 9784 -40 9844 2362
rect 9904 -40 9964 2907
<< metal3 >>
rect 0 3690 10104 3770
rect 0 274 80 3690
rect 10024 274 10104 3690
rect 0 194 10104 274
rect 0 34 10104 114
<< metal4 >>
rect 4802 3970 4902 4020
rect 5202 3970 5302 4020
use comparator_core  comparator_core_0
timestamp 1696364841
transform 1 0 3650 0 1 539
box 0 -40 2804 3481
use trim  trim_0
timestamp 1696364841
transform 0 1 730 -1 0 3332
box -1 -83 2781 2620
use trim  trim_1
timestamp 1696364841
transform 0 -1 9374 -1 0 3332
box -1 -83 2781 2620
use via2_1  via2_1_0
timestamp 1696364841
transform 0 1 3380 -1 0 1458
box 0 -40 140 40
use via2_1  via2_1_1
timestamp 1696364841
transform 0 1 6724 1 0 1318
box 0 -40 140 40
use via23  via23_0
timestamp 1696364841
transform 1 0 1198 0 1 -6
box 1 40 161 120
use via23  via23_1
timestamp 1696364841
transform 1 0 4971 0 1 -6
box 1 40 161 120
use via23  via23_2
timestamp 1696364841
transform 1 0 8744 0 1 -6
box 1 40 161 120
use via23  via23_3
timestamp 1696364841
transform 1 0 4972 0 1 3650
box 1 40 161 120
<< labels >>
flabel metal2 s 140 -40 200 -10 1 FreeSans 44 0 0 0 trim_3
port 2 nsew
flabel metal2 s 260 -40 320 -10 1 FreeSans 44 0 0 0 trim_2
port 3 nsew
flabel metal2 s 380 -40 440 -10 1 FreeSans 44 0 0 0 trim_0
port 4 nsew
flabel metal2 s 500 -40 560 -10 1 FreeSans 44 0 0 0 trim_1
port 5 nsew
flabel metal2 s 620 -40 680 -10 1 FreeSans 44 0 0 0 trim_4
port 6 nsew
flabel metal2 s 9424 -40 9484 -10 1 FreeSans 44 0 0 0 trimb_4
port 7 nsew
flabel metal2 s 9544 -40 9604 -10 1 FreeSans 44 0 0 0 trimb_1
port 8 nsew
flabel metal2 s 9664 -40 9724 -10 1 FreeSans 44 0 0 0 trimb_0
port 9 nsew
flabel metal2 s 9784 -40 9844 -10 1 FreeSans 44 0 0 0 trimb_2
port 10 nsew
flabel metal2 s 9904 -40 9964 -10 1 FreeSans 44 0 0 0 trimb_3
port 11 nsew
flabel metal2 s 4555 -40 4635 0 1 FreeSans 44 0 0 0 outn
port 12 nsew
flabel metal2 s 5469 -40 5549 0 1 FreeSans 44 0 0 0 outp
port 13 nsew
flabel metal1 s 3512 -40 3572 -10 1 FreeSans 44 0 0 0 clk
port 14 nsew
flabel metal3 s 0 194 80 274 1 FreeSans 96 0 0 0 vdd
port 16 nsew
flabel metal3 s 0 34 80 114 1 FreeSans 96 0 0 0 vss
port 17 nsew
flabel metal4 s 4802 3970 4902 4020 1 FreeSans 96 0 0 0 vn
port 19 nsew
flabel metal4 s 5202 3970 5302 4020 1 FreeSans 96 0 0 0 vp
port 20 nsew
<< properties >>
string FIXED_BBOX 0 -40 10104 4020
string path 248.100 5.850 4.500 5.850 
<< end >>
