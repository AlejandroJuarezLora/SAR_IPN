* SPICE3 file created from comparator_flat.ext - technology: sky130B

.subckt comparator_flat trim_4 trim_3 trim_2 trim_1 vp vn outp outn clk vdd trimb_1
+ trimb_2 trimb_3 trimb_4 trimb_0 trim_0 vss
X0 trim_1.n4.t11 trimb_4.t0 vss.t46 vss.t45 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 ip.t3 trim_1.n4.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 vss.t7 trim_3.t0 trim_0.n3.t5 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X3 vss.t44 trimb_4.t1 trim_1.n4.t10 vss.t43 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X4 vdd.t6 clk.t0 in.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X5 vss.t9 trim_4.t0 trim_0.n4.t15 vss.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 in.t3 trim_0.n1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 diff clk.t1 vss.t64 vss.t63 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X8 vdd.t5 clk.t2 outn.t2 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X9 vss.t50 trim_4.t1 trim_0.n4.t14 vss.t49 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X10 trim_1.n4.t9 trimb_4.t2 vss.t42 vss.t41 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X11 vss.t58 trim_2.t0 trim_0.n2 vss.t57 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X12 ip.t4 trim_1.n4.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 trim_0.n4.t13 trim_4.t2 vss.t54 vss.t53 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X14 ip.t5 trim_1.n4.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 ip.t6 trim_1.n4.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 in.t4 trim_0.n3.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 diff clk.t3 vss.t62 vss.t61 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X18 ip.t7 trim_1.n1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 ip.t8 trim_1.n3.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 ip.t9 trim_1.n3.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 trim_1.n3.t6 trimb_3.t0 vss.t52 vss.t51 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X22 vss.t40 trimb_4.t3 trim_1.n4.t8 vss.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X23 in.t5 trim_0.n4.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 trim_1.n1 trimb_1.t0 vss.t68 vss.t67 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X25 trim_0.n3.t4 trim_3.t1 vss.t3 vss.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X26 outn.t0 outp.t3 in.t0 vss.t19 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X27 trim_1.n4.t7 trimb_4.t4 vss.t38 vss.t37 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X28 vss.t13 trimb_3.t1 trim_1.n3.t1 vss.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X29 trim_0.n4.t12 trim_4.t3 vss.t48 vss.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X30 in.t6 trim_0.n3.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 ip.t10 trim_1.n4.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 vss.t36 trimb_4.t5 trim_1.n4.t6 vss.t35 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X33 in.t7 trim_0.n0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 in.t8 trim_0.n4.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 in.t9 trim_0.n4.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 ip.t11 trim_1.n3.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 ip.t2 clk.t4 vdd.t4 vdd.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X38 outp.t1 outn.t3 vdd.t7 vdd.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X39 ip.t12 trim_1.n4.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 ip.t13 trim_1.n3.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 in.t10 trim_0.n3.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 trim_0.n2 trim_2.t1 vss.t28 vss.t27 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X43 vss.t56 trimb_2.t0 trim_1.n2 vss.t55 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X44 trim_1.n3.t7 trimb_3.t2 vss.t66 vss.t65 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X45 in.t2 vn.t0 diff vss.t69 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X46 vss.t71 trim_4.t4 trim_0.n4.t11 vss.t70 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X47 in.t11 trim_0.n4.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 ip.t14 trim_1.n4.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 outp.t2 clk.t5 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X50 vss.t34 trimb_4.t6 trim_1.n4.t5 vss.t33 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X51 in.t12 trim_0.n2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 in.t13 trim_0.n4.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 trim_0.n4.t10 trim_4.t5 vss.t18 vss.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X54 in.t14 trim_0.n4.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 vss.t23 trim_0.t0 trim_0.n0 vss.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X56 vss.t16 trim_1.t0 trim_0.n1 vss.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X57 trim_1.n0 trimb_0.t0 vss.t30 vss.t29 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X58 trim_1.n2 trimb_2.t1 vss.t60 vss.t59 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X59 ip.t1 vp.t0 diff vss.t24 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X60 trim_0.n4.t9 trim_4.t6 vss.t1 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X61 ip.t15 trim_1.n2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 ip.t16 trim_1.n2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 in.t15 trim_0.n3.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 outp.t0 outn.t4 ip.t0 vss.t14 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X65 in.t16 trim_0.n4.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 vss.t26 trim_3.t2 trim_0.n3.t3 vss.t25 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X67 in.t17 trim_0.n2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 vdd.t1 outp.t4 outn.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X69 vss.t21 trim_4.t7 trim_0.n4.t8 vss.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X70 ip.t17 trim_1.n0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 in.t18 trim_0.n4.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 ip.t18 trim_1.n4.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 trim_0.n3.t2 trim_3.t3 vss.t5 vss.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X74 trim_1.n4.t4 trimb_4.t7 vss.t32 vss.t31 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X75 vss.t11 trimb_3.t3 trim_1.n3.t0 vss.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
R0 trimb_4 trimb_4.n6 281.043
R1 trimb_4.n0 trimb_4.t7 135.841
R2 trimb_4.n2 trimb_4.t5 135.841
R3 trimb_4.n2 trimb_4.t2 135.52
R4 trimb_4.n3 trimb_4.t3 135.52
R5 trimb_4.n4 trimb_4.t0 135.52
R6 trimb_4.n5 trimb_4.t6 135.52
R7 trimb_4.n1 trimb_4.t4 135.52
R8 trimb_4.n0 trimb_4.t1 135.52
R9 trimb_4.n1 trimb_4.n0 0.321152
R10 trimb_4.n5 trimb_4.n4 0.321152
R11 trimb_4.n4 trimb_4.n3 0.321152
R12 trimb_4.n3 trimb_4.n2 0.321152
R13 trimb_4.n6 trimb_4.n1 0.101043
R14 trimb_4.n6 trimb_4.n5 0.0956087
R15 vss.t61 vss.t19 716.199
R16 vss.n13 vss.t67 594.287
R17 vss.t15 vss.n37 577.361
R18 vss.n26 vss.n0 567.549
R19 vss.n26 vss.n1 563.729
R20 vss vss.n60 553.972
R21 vss.n12 vss.t59 543.674
R22 vss.t27 vss.n40 528.191
R23 vss.n23 vss.t14 346.106
R24 vss.n60 vss.n28 332.8
R25 vss.n27 vss.n26 330.272
R26 vss.n21 vss.n20 325.935
R27 vss.n49 vss.n48 325.935
R28 vss.t67 vss.n12 318.368
R29 vss.n40 vss.t15 309.301
R30 vss.n53 vss.n28 302.625
R31 vss.n60 vss 300.057
R32 vss.n36 vss.n32 271.844
R33 vss.n15 vss.n14 271.844
R34 vss.n17 vss.n16 267.671
R35 vss.n44 vss.n42 267.671
R36 vss.n34 vss.t22 237.924
R37 vss.n11 vss.t29 207.347
R38 vss.t10 vss.t51 192.654
R39 vss.t65 vss.t12 192.654
R40 vss.t43 vss.t31 192.654
R41 vss.t37 vss.t43 192.654
R42 vss.t45 vss.t39 192.654
R43 vss.t39 vss.t41 192.654
R44 vss.t41 vss.t35 192.654
R45 vss.t25 vss.t4 187.167
R46 vss.t2 vss.t6 187.167
R47 vss.t8 vss.t17 187.167
R48 vss.t47 vss.t8 187.167
R49 vss.t20 vss.t47 187.167
R50 vss.t0 vss.t49 187.167
R51 vss.t49 vss.t53 187.167
R52 vss.t53 vss.t70 187.167
R53 vss.n29 vss.t62 184.464
R54 vss.n23 vss.t37 158.368
R55 vss.n42 vss.n32 134.4
R56 vss.n16 vss.n15 134.4
R57 vss.n13 vss.n11 111.02
R58 vss.t59 vss.n7 96.327
R59 vss.n7 vss.t55 96.327
R60 vss.n18 vss.t10 96.327
R61 vss.n18 vss.t65 96.327
R62 vss.n24 vss.t33 96.327
R63 vss.n24 vss.t45 96.327
R64 vss.n41 vss.t27 93.5838
R65 vss.n41 vss.t57 93.5838
R66 vss.n45 vss.t25 93.5838
R67 vss.n45 vss.t2 93.5838
R68 vss.n56 vss.t0 93.5838
R69 vss.n57 vss.n56 90.4115
R70 vss.n22 vss.n21 73.4481
R71 vss.n50 vss.n49 73.4481
R72 vss.n26 vss.n25 71.9243
R73 vss.n37 vss.n34 71.3776
R74 vss.n48 vss.n47 69.3723
R75 vss.n44 vss.n43 69.3467
R76 vss.n42 vss.n33 69.3126
R77 vss.n20 vss.n4 69.2957
R78 vss.n17 vss.n5 69.2702
R79 vss.n16 vss.n6 69.2363
R80 vss.n39 vss.n32 67.7652
R81 vss.n15 vss.n9 67.7652
R82 vss.n54 vss.n53 67.4138
R83 vss.n39 vss.n38 64.3972
R84 vss.n36 vss.n35 64.3972
R85 vss.n9 vss.n8 64.3972
R86 vss.n14 vss.n10 64.3972
R87 vss.n50 vss.n30 60.4824
R88 vss.n22 vss.n2 60.4093
R89 vss.n53 vss.n52 60.3406
R90 vss.n49 vss.n31 60.0765
R91 vss.n21 vss.n3 60.0059
R92 vss.n54 vss.n51 59.8927
R93 vss.n29 vss.t64 58.6822
R94 vss vss.n59 44.6517
R95 vss.n59 vss.n58 44.2758
R96 vss.n59 vss.n29 39.8889
R97 vss.n20 vss.n19 38.024
R98 vss.n48 vss.n46 38.024
R99 vss.n19 vss.n17 37.6476
R100 vss.n46 vss.n44 37.6476
R101 vss.n25 vss.n22 35.3529
R102 vss.n55 vss.n50 35.3529
R103 vss.n55 vss.n54 35.3122
R104 vss.t33 vss.n23 34.2862
R105 vss vss.n39 21.4593
R106 vss vss.n9 21.4593
R107 vss vss.n36 21.0506
R108 vss.n14 vss 21.0506
R109 vss.n38 vss.t16 17.4059
R110 vss.n35 vss.t23 17.4059
R111 vss.n8 vss.t68 17.4059
R112 vss.n10 vss.t30 17.4059
R113 vss.n52 vss.t54 17.4005
R114 vss.n52 vss.t71 17.4005
R115 vss.n51 vss.t1 17.4005
R116 vss.n51 vss.t50 17.4005
R117 vss.n30 vss.t48 17.4005
R118 vss.n30 vss.t21 17.4005
R119 vss.n31 vss.t18 17.4005
R120 vss.n31 vss.t9 17.4005
R121 vss.n3 vss.t32 17.4005
R122 vss.n3 vss.t44 17.4005
R123 vss.n2 vss.t38 17.4005
R124 vss.n2 vss.t34 17.4005
R125 vss.n0 vss.t46 17.4005
R126 vss.n0 vss.t40 17.4005
R127 vss.n1 vss.t42 17.4005
R128 vss.n1 vss.t36 17.4005
R129 vss.n4 vss.t66 17.4005
R130 vss.n4 vss.t13 17.4005
R131 vss.n5 vss.t52 17.4005
R132 vss.n5 vss.t11 17.4005
R133 vss.n6 vss.t60 17.4005
R134 vss.n6 vss.t56 17.4005
R135 vss.n33 vss.t28 17.4005
R136 vss.n33 vss.t58 17.4005
R137 vss.n43 vss.t5 17.4005
R138 vss.n43 vss.t26 17.4005
R139 vss.n47 vss.t3 17.4005
R140 vss.n47 vss.t7 17.4005
R141 vss.t24 vss.t61 8.56748
R142 vss.t69 vss.t63 8.56748
R143 vss.n27 vss 7.52991
R144 vss.t14 vss.t24 5.14069
R145 vss.t19 vss.t69 5.14069
R146 vss vss.n27 5.06097
R147 vss.n28 vss 5.06097
R148 vss.n57 vss.t20 3.17281
R149 vss.n40 vss 0.986602
R150 vss.n37 vss 0.986602
R151 vss vss.n13 0.986602
R152 vss.n12 vss 0.986602
R153 vss.n16 vss.n7 0.129298
R154 vss.n42 vss.n41 0.129298
R155 vss.n19 vss.n18 0.0681222
R156 vss.n46 vss.n45 0.0681222
R157 vss.n25 vss.n24 0.0352676
R158 vss.n56 vss.n55 0.0352676
R159 vss.n58 vss.n57 0.0147549
R160 vss.n38 vss 0.00766301
R161 vss.n35 vss 0.00766301
R162 vss.n8 vss 0.00766301
R163 vss.n10 vss 0.00766301
R164 trim_1.n4.n9 trim_1.n4.t4 18.7888
R165 trim_1.n4.n6 trim_1.n4.t6 17.6293
R166 trim_1.n4.n7 trim_1.n4.t8 17.4005
R167 trim_1.n4.n7 trim_1.n4.t9 17.4005
R168 trim_1.n4.n8 trim_1.n4.t10 17.4005
R169 trim_1.n4.n8 trim_1.n4.t7 17.4005
R170 trim_1.n4.n10 trim_1.n4.t5 17.4005
R171 trim_1.n4.n10 trim_1.n4.t11 17.4005
R172 trim_1.n4.n0 trim_1.n4.t12 2.32631
R173 trim_1.n4.n2 trim_1.n4.n1 2.23987
R174 trim_1.n4.n4 trim_1.n4.n3 2.23987
R175 trim_1.n4.n1 trim_1.n4.n0 2.22263
R176 trim_1.n4.n5 trim_1.n4.n4 2.22263
R177 trim_1.n4.n3 trim_1.n4.n2 2.18815
R178 trim_1.n4.n14 trim_1.n4.t1 1.31613
R179 trim_1.n4.n11 trim_1.n4.n9 0.909983
R180 trim_1.n4.n13 trim_1.n4.n12 0.888431
R181 trim_1.n4.n14 trim_1.n4.n5 0.884681
R182 trim_1.n4.n12 trim_1.n4.n11 0.884121
R183 trim_1.n4.n14 trim_1.n4.n13 0.828086
R184 trim_1.n4.n6 trim_1.n4 0.731478
R185 trim_1.n4.n11 trim_1.n4.n10 0.500883
R186 trim_1.n4.n12 trim_1.n4.n7 0.500883
R187 trim_1.n4.n9 trim_1.n4.n8 0.500883
R188 trim_1.n4.n13 trim_1.n4.n6 0.272052
R189 trim_1.n4.n5 trim_1.n4.t3 0.0869351
R190 trim_1.n4.n4 trim_1.n4.t0 0.0869351
R191 trim_1.n4.n3 trim_1.n4.t15 0.0869351
R192 trim_1.n4.n2 trim_1.n4.t13 0.0869351
R193 trim_1.n4.n1 trim_1.n4.t14 0.0869351
R194 trim_1.n4.n0 trim_1.n4.t2 0.0869351
R195 trim_1.n4 trim_1.n4.n14 0.0608448
R196 ip.n0 ip.t2 29.756
R197 ip.n2 ip.t0 17.4313
R198 ip ip.t1 17.4118
R199 ip.t7 ip 16.6643
R200 ip.t16 ip 14.0781
R201 ip.t15 ip 11.4574
R202 ip.t10 ip 10.4971
R203 ip.t13 ip 8.89705
R204 ip.t9 ip 6.28498
R205 ip.t17 ip 4.94368
R206 ip.t7 ip 4.25505
R207 ip.t11 ip 3.69016
R208 ip.t16 ip 3.57323
R209 ip.t15 ip 2.88232
R210 ip.t4 ip.t5 2.35391
R211 ip.t15 ip.t16 2.23518
R212 ip.t3 ip.t6 2.22656
R213 ip.t7 ip.t17 2.22656
R214 ip.t14 ip.t18 2.20931
R215 ip.t13 ip 2.20732
R216 ip.t16 ip.t7 2.20069
R217 ip.t12 ip.t3 2.17483
R218 ip.t13 ip.t15 2.17483
R219 ip.t9 ip.t13 2.08671
R220 ip.t8 ip.t11 2.08671
R221 ip.t11 ip.t9 2.06947
R222 ip.t18 ip.t10 2.06178
R223 ip.t12 ip.t14 1.83768
R224 ip.t9 ip 1.65853
R225 ip.n0 ip.t4 1.6092
R226 ip.n1 ip.t12 1.50144
R227 ip.t8 ip 1.07809
R228 ip.t11 ip 0.97444
R229 ip.n2 ip.n1 0.556421
R230 ip.t6 ip.n0 0.475611
R231 ip ip.t8 0.427224
R232 ip.n1 ip 0.418263
R233 ip ip.n2 0.3005
R234 ip.t8 ip 0.285803
R235 trim_3.n0 trim_3.t3 135.841
R236 trim_3.n1 trim_3.t0 135.841
R237 trim_3.n1 trim_3.t1 135.52
R238 trim_3.n0 trim_3.t2 135.52
R239 trim_3 trim_3.n2 69.1659
R240 trim_3.n2 trim_3.n0 0.106478
R241 trim_3.n2 trim_3.n1 0.0901739
R242 trim_0.n3.n3 trim_0.n3.t2 18.7775
R243 trim_0.n3.n4 trim_0.n3.t5 17.8604
R244 trim_0.n3.n2 trim_0.n3.t3 17.4005
R245 trim_0.n3.n2 trim_0.n3.t4 17.4005
R246 trim_0.n3 trim_0.n3.n4 3.34964
R247 trim_0.n3.n0 trim_0.n3.t7 2.32531
R248 trim_0.n3.n1 trim_0.n3.n0 2.22263
R249 trim_0.n3 trim_0.n3.n1 1.78672
R250 trim_0.n3.n4 trim_0.n3.n3 0.901362
R251 trim_0.n3.n3 trim_0.n3.n2 0.459422
R252 trim_0.n3 trim_0.n3.t0 0.415082
R253 trim_0.n3.n1 trim_0.n3.t1 0.0869351
R254 trim_0.n3.n0 trim_0.n3.t6 0.0869351
R255 clk.n3 clk.t4 144.121
R256 clk.n1 clk.t5 144.065
R257 clk.n3 clk.t0 142.686
R258 clk.n1 clk.t2 142.675
R259 clk.n0 clk.t3 135.874
R260 clk.n0 clk.t1 135.453
R261 clk.n2 clk.n0 10.8293
R262 clk.n4 clk.n3 2.42642
R263 clk.n2 clk.n1 2.42528
R264 clk clk.n4 1.50467
R265 clk.n4 clk.n2 1.38383
R266 in.n0 in.t1 30.0626
R267 in.n2 in.t0 17.4313
R268 in in.t2 17.431
R269 in.t3 in 16.6643
R270 in.t12 in 14.0781
R271 in.t17 in 11.4574
R272 in.t5 in 10.5575
R273 in.t15 in 8.89705
R274 in.t4 in 6.28498
R275 in.t7 in 4.94368
R276 in.t3 in 4.25505
R277 in.t6 in 3.69016
R278 in.t12 in 3.57323
R279 in.t17 in 2.88232
R280 in.t13 in.t11 2.35491
R281 in.t17 in.t12 2.23518
R282 in.t9 in.t8 2.22656
R283 in.t3 in.t7 2.22656
R284 in.t16 in.t14 2.20931
R285 in.t15 in 2.20732
R286 in.t12 in.t3 2.20069
R287 in.t18 in.t9 2.17483
R288 in.t15 in.t17 2.17483
R289 in.t4 in.t15 2.08671
R290 in.t10 in.t6 2.08671
R291 in.t6 in.t4 2.06947
R292 in.t14 in.t5 2.06178
R293 in.t18 in.t16 1.85061
R294 in.n1 in.t18 1.73851
R295 in.n0 in.t13 1.68679
R296 in.t4 in 1.65853
R297 in.t10 in 1.07809
R298 in.t6 in 0.97444
R299 in.n1 in 0.503789
R300 in.n2 in.n1 0.470895
R301 in in.t10 0.427224
R302 in.t8 in.n0 0.398025
R303 in in.n2 0.297615
R304 in.t10 in 0.285803
R305 vdd.n0 vdd.t2 134.669
R306 vdd.n0 vdd.t0 128.083
R307 vdd vdd.n4 79.3384
R308 vdd.n4 vdd.n3 69.9591
R309 vdd.n2 vdd.n1 68.0792
R310 vdd.n2 vdd.t3 51.9559
R311 vdd.n4 vdd.t4 51.9559
R312 vdd.n1 vdd.t7 51.9559
R313 vdd.n1 vdd.t1 51.2175
R314 vdd.n2 vdd.t5 50.2329
R315 vdd.n4 vdd.t6 50.2329
R316 vdd.n3 vdd.n2 11.2557
R317 vdd.n3 vdd.n0 0.000773431
R318 trim_4 trim_4.n6 281.05
R319 trim_4.n0 trim_4.t5 135.841
R320 trim_4.n2 trim_4.t4 135.841
R321 trim_4.n2 trim_4.t2 135.52
R322 trim_4.n3 trim_4.t1 135.52
R323 trim_4.n4 trim_4.t6 135.52
R324 trim_4.n5 trim_4.t7 135.52
R325 trim_4.n1 trim_4.t3 135.52
R326 trim_4.n0 trim_4.t0 135.52
R327 trim_4.n1 trim_4.n0 0.321152
R328 trim_4.n5 trim_4.n4 0.321152
R329 trim_4.n4 trim_4.n3 0.321152
R330 trim_4.n3 trim_4.n2 0.321152
R331 trim_4.n6 trim_4.n1 0.101043
R332 trim_4.n6 trim_4.n5 0.0956087
R333 trim_0.n4.n8 trim_0.n4.t10 18.7845
R334 trim_0.n4 trim_0.n4.t11 17.4527
R335 trim_0.n4.n7 trim_0.n4.t15 17.4005
R336 trim_0.n4.n7 trim_0.n4.t12 17.4005
R337 trim_0.n4.n9 trim_0.n4.t8 17.4005
R338 trim_0.n4.n9 trim_0.n4.t9 17.4005
R339 trim_0.n4.n11 trim_0.n4.t14 17.4005
R340 trim_0.n4.n11 trim_0.n4.t13 17.4005
R341 trim_0.n4.n0 trim_0.n4.t4 2.32675
R342 trim_0.n4.n2 trim_0.n4.n1 2.23987
R343 trim_0.n4.n4 trim_0.n4.n3 2.23987
R344 trim_0.n4.n1 trim_0.n4.n0 2.22263
R345 trim_0.n4.n5 trim_0.n4.n4 2.22263
R346 trim_0.n4.n3 trim_0.n4.n2 2.18815
R347 trim_0.n4.n6 trim_0.n4.t7 1.31656
R348 trim_0.n4.n10 trim_0.n4.n8 0.909983
R349 trim_0.n4.n13 trim_0.n4.n12 0.888431
R350 trim_0.n4.n6 trim_0.n4.n5 0.884681
R351 trim_0.n4.n12 trim_0.n4.n10 0.884121
R352 trim_0.n4.n13 trim_0.n4.n6 0.828086
R353 trim_0.n4.n12 trim_0.n4.n11 0.496573
R354 trim_0.n4.n8 trim_0.n4.n7 0.496573
R355 trim_0.n4.n10 trim_0.n4.n9 0.496573
R356 trim_0.n4 trim_0.n4.n14 0.280672
R357 trim_0.n4.n14 trim_0.n4.n13 0.267741
R358 trim_0.n4.n14 trim_0.n4 0.17713
R359 trim_0.n4.n5 trim_0.n4.t2 0.0873744
R360 trim_0.n4.n4 trim_0.n4.t1 0.0873744
R361 trim_0.n4.n3 trim_0.n4.t0 0.0873744
R362 trim_0.n4.n2 trim_0.n4.t5 0.0873744
R363 trim_0.n4.n1 trim_0.n4.t6 0.0873744
R364 trim_0.n4.n0 trim_0.n4.t3 0.0873744
R365 outn.n5 outn.t3 143.925
R366 outn.n5 outn.t4 136.066
R367 outn.n0 outn.t2 28.7495
R368 outn.n2 outn.t1 28.5716
R369 outn.n8 outn.t0 17.5641
R370 outn.n6 outn.n5 10.2168
R371 outn.n1 outn 2.2505
R372 outn.n0 outn 1.25578
R373 outn.n4 outn.n3 1.04738
R374 outn.n3 outn 0.725852
R375 outn.n4 outn 0.563
R376 outn.n1 outn.n0 0.535656
R377 outn.n8 outn.n7 0.203625
R378 outn.n7 outn 0.192808
R379 outn.n2 outn.n1 0.144866
R380 outn.n3 outn.n2 0.144866
R381 outn outn.n8 0.109875
R382 outn.n6 outn.n4 0.0774231
R383 outn.n7 outn.n6 0.0774231
R384 outn.n8 outn 0.0439783
R385 trim_2 trim_2.n0 146.404
R386 trim_2.n0 trim_2.t0 135.803
R387 trim_2.n0 trim_2.t1 135.52
R388 trim_1.n3.n2 trim_1.n3.t6 18.7818
R389 trim_1.n3.n1 trim_1.n3.t0 17.4005
R390 trim_1.n3.n1 trim_1.n3.t7 17.4005
R391 trim_1.n3 trim_1.n3.n0 2.3324
R392 trim_1.n3.t3 trim_1.n3.t5 2.32575
R393 trim_1.n3.t4 trim_1.n3.t3 2.22263
R394 trim_1.n3.n0 trim_1.n3.t4 1.78672
R395 trim_1.n3 trim_1.n3.t1 1.01774
R396 trim_1.n3.t1 trim_1.n3.n2 0.901362
R397 trim_1.n3.n2 trim_1.n3.n1 0.464714
R398 trim_1.n3.n0 trim_1.n3.t2 0.415521
R399 trimb_3.n0 trimb_3.t0 135.841
R400 trimb_3.n1 trimb_3.t1 135.841
R401 trimb_3.n1 trimb_3.t2 135.52
R402 trimb_3.n0 trimb_3.t3 135.52
R403 trimb_3 trimb_3.n2 69.1347
R404 trimb_3.n2 trimb_3.n0 0.106478
R405 trimb_3.n2 trimb_3.n1 0.0901739
R406 trimb_1 trimb_1.t0 135.52
R407 outp.n5 outp.t4 143.425
R408 outp.n5 outp.t3 136.528
R409 outp.n0 outp.t2 28.7517
R410 outp.n2 outp.t1 28.5716
R411 outp outp.t0 17.4935
R412 outp.n6 outp.n5 10.1595
R413 outp.n1 outp 2.21144
R414 outp.n0 outp 1.41784
R415 outp.n4 outp 0.961438
R416 outp.n3 outp 0.810984
R417 outp.n8 outp.n7 0.688
R418 outp.n4 outp.n3 0.609875
R419 outp.n1 outp.n0 0.535656
R420 outp.n7 outp 0.379406
R421 outp.n2 outp.n1 0.165823
R422 outp.n3 outp.n2 0.165823
R423 outp outp.n8 0.0708125
R424 outp.n6 outp.n4 0.0512812
R425 outp.n7 outp.n6 0.0512812
R426 outp.n8 outp 0.0439783
R427 trimb_2 trimb_2.n0 146.279
R428 trimb_2.n0 trimb_2.t0 135.803
R429 trimb_2.n0 trimb_2.t1 135.52
R430 vn vn.t0 132.754
R431 trim_0 trim_0.t0 135.525
R432 trim_1 trim_1.t0 135.52
R433 trimb_0 trimb_0.t0 135.525
R434 vp vp.t0 133.359
C0 trim_3 vdd 3.79e-19
C1 trim_2 trim_0 7.61e-19
C2 trim_2 in 0.0958f
C3 trim_0 trim_0.n4 0.0101f
C4 trim_3 trim_0.n3 0.231f
C5 vdd diff 0.00122f
C6 trim_0.n4 in 4.88f
C7 trim_1.n3 ip 2.47f
C8 trimb_2 clk 4.96e-19
C9 ip outp 0.266f
C10 trim_2 clk 6.22e-19
C11 trim_0.n0 trim_0.n2 1.16e-19
C12 ip vn 0.0069f
C13 vp in 2.54e-19
C14 trim_0.n4 clk 0.0697f
C15 ip outn 0.0303f
C16 trim_2 trim_0.n4 0.0234f
C17 vdd in 0.257f
C18 trim_1.n4 trim_1.n2 0.187f
C19 trim_3 outp 4.66e-19
C20 vp clk 0.01f
C21 trim_1.n2 trim_1.n1 0.217f
C22 in trim_0.n3 2.47f
C23 diff outp 0.00287f
C24 trim_0.n0 trim_1 0.0594f
C25 trim_0.n4 vp 0.00105f
C26 vdd trimb_2 4.99e-19
C27 diff vn 0.0177f
C28 trim_3 outn 9.68e-20
C29 vdd clk 0.896f
C30 diff outn 0.00328f
C31 trim_0.n3 clk 6.61e-19
C32 trim_2 vdd 4.71e-19
C33 trim_3 trim_0.n2 0.127f
C34 trim_2 trim_0.n3 0.00123f
C35 trimb_0 trim_1.n2 9.83e-19
C36 vdd trim_0.n4 0.0514f
C37 trim_0.n4 trim_0.n3 0.461f
C38 trim_1.n2 ip 1.18f
C39 trim_1.n4 trim_1.n1 0.0527f
C40 trim_0.n2 trim_0.n1 0.217f
C41 in outp 0.026f
C42 vdd vp 3.91e-19
C43 in vn 0.0349f
C44 trim_1.n3 trimb_2 0.00123f
C45 trim_3 trim_1 7.6e-20
C46 in outn 0.239f
C47 clk outp 0.0741f
C48 trimb_0 trim_1.n4 0.0101f
C49 trimb_0 trim_1.n1 0.00397f
C50 trim_1.n4 ip 4.88f
C51 trim_0 trim_0.n2 9.83e-19
C52 trim_1 trim_0.n1 0.183f
C53 vn clk 0.0119f
C54 ip trim_1.n1 0.578f
C55 in trim_0.n2 1.18f
C56 trim_1.n2 trim_1.n0 1.16e-19
C57 trim_0.n4 outp 0.0098f
C58 clk outn 0.122f
C59 trim_3 trim_4 0.016f
C60 diff trim_4 4.62e-20
C61 trim_0.n4 vn 0.00127f
C62 trim_0.n4 outn 0.00841f
C63 trim_0.n2 clk 5.42e-19
C64 vp outp 8.08e-19
C65 trim_1 trim_0 0.0416f
C66 trim_1 in 0.0877f
C67 trimb_0 ip 0.0297f
C68 trim_2 trim_0.n2 0.243f
C69 trim_1.n4 diff 0.00626f
C70 vp vn 0.0631f
C71 trim_0.n4 trim_0.n2 0.187f
C72 trim_1.n4 trim_1.n0 0.052f
C73 vdd outp 0.489f
C74 vp outn 0.0123f
C75 trim_1.n1 trim_1.n0 0.207f
C76 trim_0.n3 outp 5.99e-20
C77 vdd vn 3.39e-19
C78 trim_1 clk 1.34e-19
C79 trim_0.n0 trim_0.n1 0.207f
C80 in trim_4 0.104f
C81 trim_1.n2 trimb_2 0.243f
C82 vdd outn 0.469f
C83 trim_1.n2 clk 5.88e-20
C84 trim_2 trim_1 0.0693f
C85 trim_1 trim_0.n4 0.0154f
C86 diff ip 0.158f
C87 trim_1.n4 in 0.0156f
C88 trimb_0 trim_1.n0 0.117f
C89 trim_4 clk 0.00154f
C90 trim_0.n3 trim_0.n2 0.264f
C91 ip trim_1.n0 0.556f
C92 trim_1.n3 outp 1.93e-20
C93 trim_0.n0 trim_0 0.117f
C94 trim_0.n0 in 0.556f
C95 trim_1.n4 trimb_2 0.0234f
C96 trim_0.n4 trim_4 0.359f
C97 trim_1.n4 clk 0.0233f
C98 trim_1.n1 trimb_2 0.0715f
C99 trim_1.n3 outn 9.64e-20
C100 vn outp 0.013f
C101 outn outp 0.619f
C102 trim_1 trim_0.n3 4.9e-20
C103 trim_3 trim_0.n1 0.00122f
C104 trim_1.n4 trim_0.n4 0.12f
C105 ip in 0.295f
C106 vn outn 0.00126f
C107 trim_0.n0 trim_2 2.84e-19
C108 trim_0.n0 trim_0.n4 0.052f
C109 trimb_0 trimb_2 0.00129f
C110 trim_1.n4 vp 0.00193f
C111 trim_0.n3 trim_4 0.319f
C112 ip trimb_2 0.0958f
C113 ip clk 0.0863f
C114 vdd trim_1.n4 0.0573f
C115 trim_3 in 0.102f
C116 trim_1.n3 trim_1.n2 0.264f
C117 trim_0.n4 ip 0.0152f
C118 diff in 0.148f
C119 trim_0 trim_0.n1 0.00397f
C120 in trim_0.n1 0.578f
C121 trim_3 clk 0.00176f
C122 ip vp 0.0206f
C123 diff clk 0.104f
C124 trim_3 trim_2 0.0317f
C125 trim_0.n1 clk 5.25e-20
C126 trimb_2 trim_1.n0 2.84e-19
C127 trim_3 trim_0.n4 0.0166f
C128 trim_1.n4 trim_1.n3 0.461f
C129 vdd ip 0.289f
C130 diff trim_0.n4 0.00539f
C131 trim_1 trim_0.n2 0.0074f
C132 trim_2 trim_0.n1 0.0715f
C133 trim_0 in 0.0297f
C134 trim_0.n4 trim_0.n1 0.0527f
C135 trim_1.n4 outp 0.0114f
C136 diff vp 0.0486f
C137 trim_1.n4 vn 2.73e-20
C138 trim_4 trim_0.n2 0.00188f
C139 trim_1.n4 outn 0.011f
C140 in clk 0.326f
.ends

