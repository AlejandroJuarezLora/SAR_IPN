magic
tech sky130B
timestamp 1696364841
<< error_p >>
rect -548 136 548 154
rect -548 -176 -530 136
rect -513 101 513 119
rect -513 -141 -495 101
rect 495 -141 513 101
rect -513 -159 513 -141
rect 530 -176 548 136
rect -548 -194 548 -176
<< pwell >>
rect -543 106 543 149
rect -543 -146 -500 106
rect 500 -146 543 106
rect -543 -189 543 -146
<< nsubdiff >>
rect -530 119 530 136
rect -530 -159 -513 119
rect 513 -159 530 119
rect -530 -176 530 -159
<< locali >>
rect -530 119 530 136
rect -530 -159 -513 119
rect 513 -159 530 119
rect -530 -176 530 -159
<< properties >>
string FIXED_BBOX -521 -167 521 127
<< end >>
