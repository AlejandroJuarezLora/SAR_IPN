magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 774 542
<< pwell >>
rect 1 -19 696 163
rect 30 -57 64 -19
<< scnmos >>
rect 79 7 109 137
rect 267 7 297 137
rect 362 7 392 137
rect 480 7 510 137
rect 580 7 610 137
<< scpmoshvt >>
rect 79 257 109 457
rect 267 257 297 457
rect 362 257 392 457
rect 480 257 510 457
rect 580 257 610 457
<< ndiff >>
rect 27 121 79 137
rect 27 87 35 121
rect 69 87 79 121
rect 27 53 79 87
rect 27 19 35 53
rect 69 19 79 53
rect 27 7 79 19
rect 109 121 161 137
rect 109 87 119 121
rect 153 87 161 121
rect 109 53 161 87
rect 109 19 119 53
rect 153 19 161 53
rect 109 7 161 19
rect 215 121 267 137
rect 215 87 223 121
rect 257 87 267 121
rect 215 53 267 87
rect 215 19 223 53
rect 257 19 267 53
rect 215 7 267 19
rect 297 53 362 137
rect 297 19 313 53
rect 347 19 362 53
rect 297 7 362 19
rect 392 121 480 137
rect 392 87 402 121
rect 436 87 480 121
rect 392 53 480 87
rect 392 19 402 53
rect 436 19 480 53
rect 392 7 480 19
rect 510 7 580 137
rect 610 121 670 137
rect 610 87 628 121
rect 662 87 670 121
rect 610 53 670 87
rect 610 19 628 53
rect 662 19 670 53
rect 610 7 670 19
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 377 79 411
rect 27 343 35 377
rect 69 343 79 377
rect 27 309 79 343
rect 27 275 35 309
rect 69 275 79 309
rect 27 257 79 275
rect 109 445 161 457
rect 109 411 119 445
rect 153 411 161 445
rect 109 377 161 411
rect 109 343 119 377
rect 153 343 161 377
rect 109 309 161 343
rect 109 275 119 309
rect 153 275 161 309
rect 109 257 161 275
rect 215 445 267 457
rect 215 411 223 445
rect 257 411 267 445
rect 215 377 267 411
rect 215 343 223 377
rect 257 343 267 377
rect 215 257 267 343
rect 297 257 362 457
rect 392 445 480 457
rect 392 411 402 445
rect 436 411 480 445
rect 392 377 480 411
rect 392 343 402 377
rect 436 343 480 377
rect 392 309 480 343
rect 392 275 402 309
rect 436 275 480 309
rect 392 257 480 275
rect 510 445 580 457
rect 510 411 528 445
rect 562 411 580 445
rect 510 377 580 411
rect 510 343 528 377
rect 562 343 580 377
rect 510 257 580 343
rect 610 445 670 457
rect 610 411 628 445
rect 662 411 670 445
rect 610 377 670 411
rect 610 343 628 377
rect 662 343 670 377
rect 610 309 670 343
rect 610 275 628 309
rect 662 275 670 309
rect 610 257 670 275
<< ndiffc >>
rect 35 87 69 121
rect 35 19 69 53
rect 119 87 153 121
rect 119 19 153 53
rect 223 87 257 121
rect 223 19 257 53
rect 313 19 347 53
rect 402 87 436 121
rect 402 19 436 53
rect 628 87 662 121
rect 628 19 662 53
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 35 275 69 309
rect 119 411 153 445
rect 119 343 153 377
rect 119 275 153 309
rect 223 411 257 445
rect 223 343 257 377
rect 402 411 436 445
rect 402 343 436 377
rect 402 275 436 309
rect 528 411 562 445
rect 528 343 562 377
rect 628 411 662 445
rect 628 343 662 377
rect 628 275 662 309
<< poly >>
rect 79 457 109 483
rect 267 457 297 483
rect 362 457 392 483
rect 480 457 510 483
rect 580 457 610 483
rect 79 219 109 257
rect 267 225 297 257
rect 362 225 392 257
rect 480 225 510 257
rect 580 225 610 257
rect 79 209 152 219
rect 79 175 102 209
rect 136 175 152 209
rect 79 165 152 175
rect 266 209 320 225
rect 266 175 276 209
rect 310 175 320 209
rect 79 137 109 165
rect 266 159 320 175
rect 362 209 438 225
rect 362 175 394 209
rect 428 175 438 209
rect 362 159 438 175
rect 480 209 538 225
rect 480 175 494 209
rect 528 175 538 209
rect 480 159 538 175
rect 580 209 715 225
rect 580 175 665 209
rect 699 175 715 209
rect 580 159 715 175
rect 267 137 297 159
rect 362 137 392 159
rect 480 137 510 159
rect 580 137 610 159
rect 79 -19 109 7
rect 267 -19 297 7
rect 362 -19 392 7
rect 480 -19 510 7
rect 580 -19 610 7
<< polycont >>
rect 102 175 136 209
rect 276 175 310 209
rect 394 175 428 209
rect 494 175 528 209
rect 665 175 699 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 17 445 85 453
rect 17 411 35 445
rect 69 411 85 445
rect 17 377 85 411
rect 17 343 35 377
rect 69 343 85 377
rect 17 309 85 343
rect 17 275 35 309
rect 69 275 85 309
rect 17 259 85 275
rect 119 445 153 487
rect 119 377 153 411
rect 119 309 153 343
rect 207 445 257 487
rect 207 411 223 445
rect 207 377 257 411
rect 207 343 223 377
rect 207 327 257 343
rect 386 445 452 453
rect 386 411 402 445
rect 436 411 452 445
rect 386 377 452 411
rect 386 343 402 377
rect 436 343 452 377
rect 386 309 452 343
rect 512 445 578 487
rect 512 411 528 445
rect 562 411 578 445
rect 512 377 578 411
rect 512 343 528 377
rect 562 343 578 377
rect 512 327 578 343
rect 612 445 678 453
rect 612 411 628 445
rect 662 411 678 445
rect 612 377 678 411
rect 612 343 628 377
rect 662 343 678 377
rect 386 293 402 309
rect 119 259 153 275
rect 191 275 402 293
rect 436 293 452 309
rect 612 309 678 343
rect 612 293 628 309
rect 436 275 628 293
rect 662 275 678 309
rect 191 259 678 275
rect 17 137 52 259
rect 191 209 225 259
rect 86 175 102 209
rect 136 175 225 209
rect 260 209 344 215
rect 260 175 276 209
rect 310 175 344 209
rect 378 209 444 215
rect 378 175 394 209
rect 428 175 444 209
rect 478 209 544 215
rect 478 175 494 209
rect 528 175 544 209
rect 17 121 85 137
rect 17 87 35 121
rect 69 87 85 121
rect 17 53 85 87
rect 17 19 35 53
rect 69 19 85 53
rect 17 11 85 19
rect 119 121 169 137
rect 153 87 169 121
rect 119 53 169 87
rect 153 19 169 53
rect 119 -23 169 19
rect 207 121 452 141
rect 207 87 223 121
rect 257 107 402 121
rect 257 87 273 107
rect 207 53 273 87
rect 386 87 402 107
rect 436 87 452 121
rect 207 19 223 53
rect 257 19 273 53
rect 207 11 273 19
rect 307 53 352 69
rect 307 19 313 53
rect 347 19 352 53
rect 307 -23 352 19
rect 386 53 452 87
rect 386 19 402 53
rect 436 19 452 53
rect 386 11 452 19
rect 578 133 612 259
rect 649 209 719 225
rect 649 175 665 209
rect 699 175 719 209
rect 578 121 678 133
rect 578 87 628 121
rect 662 87 678 121
rect 578 53 678 87
rect 578 19 628 53
rect 662 19 678 53
rect 578 11 678 19
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
<< metal1 >>
rect 0 521 736 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 0 456 736 487
rect 0 -23 736 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
rect 0 -88 736 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 o211a_1
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 673 181 707 215 0 FreeSans 250 0 0 0 C1
port 11 nsew
flabel locali s 494 181 528 215 0 FreeSans 250 0 0 0 B1
port 10 nsew
flabel locali s 402 181 436 215 0 FreeSans 250 0 0 0 A2
port 9 nsew
flabel locali s 310 181 344 215 0 FreeSans 250 0 0 0 A1
port 8 nsew
flabel locali s 30 45 64 79 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 30 385 64 419 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 30 317 64 351 0 FreeSans 250 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 736 504
string path 0.000 -1.000 18.400 -1.000 
<< end >>
