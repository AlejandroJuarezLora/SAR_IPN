magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 2154 542
<< pwell >>
rect 903 117 1089 161
rect 1633 117 2075 163
rect 1 -19 2075 117
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 109 91
rect 163 7 193 91
rect 418 7 448 91
rect 513 7 543 79
rect 609 7 639 79
rect 775 7 805 91
rect 847 7 877 91
rect 979 7 1009 135
rect 1078 7 1108 79
rect 1187 7 1217 79
rect 1283 7 1313 91
rect 1432 7 1462 91
rect 1523 7 1553 91
rect 1711 7 1741 137
rect 1795 7 1825 137
rect 1879 7 1909 137
rect 1963 7 1993 137
<< scpmoshvt >>
rect 79 323 109 451
rect 163 323 193 451
rect 430 373 460 457
rect 522 373 552 457
rect 621 373 651 457
rect 761 373 791 457
rect 858 373 888 457
rect 1055 289 1085 457
rect 1154 373 1184 457
rect 1240 373 1270 457
rect 1324 373 1354 457
rect 1432 373 1462 457
rect 1516 373 1546 457
rect 1711 257 1741 457
rect 1795 257 1825 457
rect 1879 257 1909 457
rect 1963 257 1993 457
<< ndiff >>
rect 27 79 79 91
rect 27 45 35 79
rect 69 45 79 79
rect 27 7 79 45
rect 109 53 163 91
rect 109 19 119 53
rect 153 19 163 53
rect 109 7 163 19
rect 193 79 245 91
rect 193 45 203 79
rect 237 45 245 79
rect 193 7 245 45
rect 313 49 418 91
rect 313 15 325 49
rect 359 15 418 49
rect 313 7 418 15
rect 448 79 498 91
rect 929 91 979 135
rect 657 79 775 91
rect 448 55 513 79
rect 448 21 458 55
rect 492 21 513 55
rect 448 7 513 21
rect 543 55 609 79
rect 543 21 565 55
rect 599 21 609 55
rect 543 7 609 21
rect 639 7 775 79
rect 805 7 847 91
rect 877 53 979 91
rect 877 19 911 53
rect 945 19 979 53
rect 877 7 979 19
rect 1009 79 1063 135
rect 1659 123 1711 137
rect 1233 79 1283 91
rect 1009 49 1078 79
rect 1009 15 1023 49
rect 1057 15 1078 49
rect 1009 7 1078 15
rect 1108 53 1187 79
rect 1108 19 1133 53
rect 1167 19 1187 53
rect 1108 7 1187 19
rect 1217 7 1283 79
rect 1313 49 1432 91
rect 1313 15 1345 49
rect 1379 15 1432 49
rect 1313 7 1432 15
rect 1462 7 1523 91
rect 1553 69 1605 91
rect 1553 35 1563 69
rect 1597 35 1605 69
rect 1553 7 1605 35
rect 1659 89 1667 123
rect 1701 89 1711 123
rect 1659 55 1711 89
rect 1659 21 1667 55
rect 1701 21 1711 55
rect 1659 7 1711 21
rect 1741 123 1795 137
rect 1741 89 1751 123
rect 1785 89 1795 123
rect 1741 55 1795 89
rect 1741 21 1751 55
rect 1785 21 1795 55
rect 1741 7 1795 21
rect 1825 55 1879 137
rect 1825 21 1835 55
rect 1869 21 1879 55
rect 1825 7 1879 21
rect 1909 123 1963 137
rect 1909 89 1919 123
rect 1953 89 1963 123
rect 1909 55 1963 89
rect 1909 21 1919 55
rect 1953 21 1963 55
rect 1909 7 1963 21
rect 1993 55 2049 137
rect 1993 21 2003 55
rect 2037 21 2049 55
rect 1993 7 2049 21
<< pdiff >>
rect 27 437 79 451
rect 27 403 35 437
rect 69 403 79 437
rect 27 369 79 403
rect 27 335 35 369
rect 69 335 79 369
rect 27 323 79 335
rect 109 421 163 451
rect 109 387 119 421
rect 153 387 163 421
rect 109 323 163 387
rect 193 437 245 451
rect 193 403 203 437
rect 237 403 245 437
rect 193 369 245 403
rect 378 445 430 457
rect 378 411 386 445
rect 420 411 430 445
rect 378 373 430 411
rect 460 437 522 457
rect 460 403 470 437
rect 504 403 522 437
rect 460 373 522 403
rect 552 443 621 457
rect 552 409 563 443
rect 597 409 621 443
rect 552 373 621 409
rect 651 419 761 457
rect 651 385 717 419
rect 751 385 761 419
rect 651 373 761 385
rect 791 435 858 457
rect 791 401 814 435
rect 848 401 858 435
rect 791 373 858 401
rect 888 419 940 457
rect 888 385 898 419
rect 932 385 940 419
rect 888 373 940 385
rect 1003 445 1055 457
rect 1003 411 1011 445
rect 1045 411 1055 445
rect 193 335 203 369
rect 237 335 245 369
rect 193 323 245 335
rect 1003 289 1055 411
rect 1085 437 1154 457
rect 1085 403 1099 437
rect 1133 403 1154 437
rect 1085 373 1154 403
rect 1184 444 1240 457
rect 1184 410 1196 444
rect 1230 410 1240 444
rect 1184 373 1240 410
rect 1270 373 1324 457
rect 1354 445 1432 457
rect 1354 411 1388 445
rect 1422 411 1432 445
rect 1354 373 1432 411
rect 1462 419 1516 457
rect 1462 385 1472 419
rect 1506 385 1516 419
rect 1462 373 1516 385
rect 1546 445 1600 457
rect 1546 411 1558 445
rect 1592 411 1600 445
rect 1546 373 1600 411
rect 1659 445 1711 457
rect 1659 411 1667 445
rect 1701 411 1711 445
rect 1659 377 1711 411
rect 1085 289 1139 373
rect 1659 343 1667 377
rect 1701 343 1711 377
rect 1659 257 1711 343
rect 1741 437 1795 457
rect 1741 403 1751 437
rect 1785 403 1795 437
rect 1741 369 1795 403
rect 1741 335 1751 369
rect 1785 335 1795 369
rect 1741 301 1795 335
rect 1741 267 1751 301
rect 1785 267 1795 301
rect 1741 257 1795 267
rect 1825 437 1879 457
rect 1825 403 1835 437
rect 1869 403 1879 437
rect 1825 369 1879 403
rect 1825 335 1835 369
rect 1869 335 1879 369
rect 1825 257 1879 335
rect 1909 437 1963 457
rect 1909 403 1919 437
rect 1953 403 1963 437
rect 1909 369 1963 403
rect 1909 335 1919 369
rect 1953 335 1963 369
rect 1909 301 1963 335
rect 1909 267 1919 301
rect 1953 267 1963 301
rect 1909 257 1963 267
rect 1993 437 2054 457
rect 1993 403 2003 437
rect 2037 403 2054 437
rect 1993 369 2054 403
rect 1993 335 2003 369
rect 2037 335 2054 369
rect 1993 257 2054 335
<< ndiffc >>
rect 35 45 69 79
rect 119 19 153 53
rect 203 45 237 79
rect 325 15 359 49
rect 458 21 492 55
rect 565 21 599 55
rect 911 19 945 53
rect 1023 15 1057 49
rect 1133 19 1167 53
rect 1345 15 1379 49
rect 1563 35 1597 69
rect 1667 89 1701 123
rect 1667 21 1701 55
rect 1751 89 1785 123
rect 1751 21 1785 55
rect 1835 21 1869 55
rect 1919 89 1953 123
rect 1919 21 1953 55
rect 2003 21 2037 55
<< pdiffc >>
rect 35 403 69 437
rect 35 335 69 369
rect 119 387 153 421
rect 203 403 237 437
rect 386 411 420 445
rect 470 403 504 437
rect 563 409 597 443
rect 717 385 751 419
rect 814 401 848 435
rect 898 385 932 419
rect 1011 411 1045 445
rect 203 335 237 369
rect 1099 403 1133 437
rect 1196 410 1230 444
rect 1388 411 1422 445
rect 1472 385 1506 419
rect 1558 411 1592 445
rect 1667 411 1701 445
rect 1667 343 1701 377
rect 1751 403 1785 437
rect 1751 335 1785 369
rect 1751 267 1785 301
rect 1835 403 1869 437
rect 1835 335 1869 369
rect 1919 403 1953 437
rect 1919 335 1953 369
rect 1919 267 1953 301
rect 2003 403 2037 437
rect 2003 335 2037 369
<< poly >>
rect 79 451 109 477
rect 163 451 193 477
rect 430 457 460 483
rect 522 457 552 483
rect 621 457 651 483
rect 761 457 791 483
rect 858 457 888 483
rect 1055 457 1085 483
rect 1154 457 1184 483
rect 1240 457 1270 483
rect 1324 457 1354 483
rect 1432 457 1462 483
rect 1516 457 1546 483
rect 1711 457 1741 483
rect 1795 457 1825 483
rect 1879 457 1909 483
rect 1963 457 1993 483
rect 79 308 109 323
rect 46 278 109 308
rect 46 225 76 278
rect 163 234 193 323
rect 430 286 460 373
rect 522 335 552 373
rect 22 209 76 225
rect 22 175 32 209
rect 66 175 76 209
rect 118 224 193 234
rect 118 190 134 224
rect 168 190 193 224
rect 331 270 460 286
rect 506 325 572 335
rect 506 291 522 325
rect 556 291 572 325
rect 506 281 572 291
rect 331 236 341 270
rect 375 256 460 270
rect 375 236 448 256
rect 621 239 651 373
rect 761 315 791 373
rect 761 299 816 315
rect 761 265 771 299
rect 805 265 816 299
rect 761 249 816 265
rect 331 220 448 236
rect 118 180 193 190
rect 22 159 76 175
rect 46 136 76 159
rect 46 106 109 136
rect 79 91 109 106
rect 163 91 193 180
rect 418 91 448 220
rect 513 209 651 239
rect 513 179 544 209
rect 490 163 544 179
rect 490 129 500 163
rect 534 129 544 163
rect 490 113 544 129
rect 586 157 652 167
rect 586 123 602 157
rect 636 123 652 157
rect 586 113 652 123
rect 513 79 543 113
rect 609 79 639 113
rect 775 91 805 249
rect 858 179 888 373
rect 1055 274 1085 289
rect 979 244 1085 274
rect 979 227 1009 244
rect 943 211 1009 227
rect 847 163 901 179
rect 847 129 857 163
rect 891 129 901 163
rect 943 177 953 211
rect 987 177 1009 211
rect 1154 239 1184 373
rect 1240 341 1270 373
rect 1226 325 1280 341
rect 1226 291 1236 325
rect 1270 291 1280 325
rect 1226 275 1280 291
rect 1154 227 1204 239
rect 1154 215 1217 227
rect 1154 209 1241 215
rect 1175 199 1241 209
rect 1175 197 1197 199
rect 943 161 1009 177
rect 979 135 1009 161
rect 1078 151 1145 167
rect 847 113 901 129
rect 847 91 877 113
rect 1078 117 1101 151
rect 1135 117 1145 151
rect 1078 101 1145 117
rect 1187 165 1197 197
rect 1231 165 1241 199
rect 1187 149 1241 165
rect 1324 189 1354 373
rect 1432 217 1462 373
rect 1516 325 1546 373
rect 1504 309 1558 325
rect 1504 275 1514 309
rect 1548 275 1558 309
rect 1504 259 1558 275
rect 1427 201 1481 217
rect 1324 173 1385 189
rect 1324 153 1341 173
rect 1078 79 1108 101
rect 1187 79 1217 149
rect 1283 139 1341 153
rect 1375 139 1385 173
rect 1427 167 1437 201
rect 1471 167 1481 201
rect 1427 151 1481 167
rect 1283 123 1385 139
rect 1283 91 1313 123
rect 1432 91 1462 151
rect 1523 91 1553 259
rect 1711 225 1741 257
rect 1795 225 1825 257
rect 1879 225 1909 257
rect 1963 225 1993 257
rect 1699 209 1993 225
rect 1699 175 1715 209
rect 1749 175 1783 209
rect 1817 175 1851 209
rect 1885 175 1919 209
rect 1953 175 1993 209
rect 1699 159 1993 175
rect 1711 137 1741 159
rect 1795 137 1825 159
rect 1879 137 1909 159
rect 1963 137 1993 159
rect 79 -19 109 7
rect 163 -19 193 7
rect 418 -19 448 7
rect 513 -19 543 7
rect 609 -19 639 7
rect 775 -19 805 7
rect 847 -19 877 7
rect 979 -19 1009 7
rect 1078 -19 1108 7
rect 1187 -19 1217 7
rect 1283 -19 1313 7
rect 1432 -19 1462 7
rect 1523 -19 1553 7
rect 1711 -19 1741 7
rect 1795 -19 1825 7
rect 1879 -19 1909 7
rect 1963 -19 1993 7
<< polycont >>
rect 32 175 66 209
rect 134 190 168 224
rect 522 291 556 325
rect 341 236 375 270
rect 771 265 805 299
rect 500 129 534 163
rect 602 123 636 157
rect 857 129 891 163
rect 953 177 987 211
rect 1236 291 1270 325
rect 1101 117 1135 151
rect 1197 165 1231 199
rect 1514 275 1548 309
rect 1341 139 1375 173
rect 1437 167 1471 201
rect 1715 175 1749 209
rect 1783 175 1817 209
rect 1851 175 1885 209
rect 1919 175 1953 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1133 521
rect 1167 487 1225 521
rect 1259 487 1317 521
rect 1351 487 1409 521
rect 1443 487 1501 521
rect 1535 487 1593 521
rect 1627 487 1685 521
rect 1719 487 1777 521
rect 1811 487 1869 521
rect 1903 487 1961 521
rect 1995 487 2053 521
rect 2087 487 2116 521
rect 18 437 69 453
rect 18 403 35 437
rect 18 369 69 403
rect 103 421 169 487
rect 103 387 119 421
rect 153 387 169 421
rect 203 437 237 453
rect 18 335 35 369
rect 203 369 237 403
rect 69 335 168 353
rect 18 319 168 335
rect 18 209 88 285
rect 18 175 32 209
rect 66 175 88 209
rect 18 155 88 175
rect 122 224 168 319
rect 122 215 134 224
rect 156 181 168 190
rect 122 121 168 181
rect 18 87 168 121
rect 18 79 69 87
rect 18 45 35 79
rect 203 79 237 317
rect 271 293 336 450
rect 370 445 420 487
rect 370 411 386 445
rect 370 395 420 411
rect 454 437 504 453
rect 454 403 470 437
rect 454 387 504 403
rect 547 443 683 453
rect 547 409 563 443
rect 597 409 683 443
rect 798 435 864 487
rect 991 445 1065 487
rect 547 387 683 409
rect 454 361 488 387
rect 409 327 488 361
rect 522 351 615 353
rect 283 270 375 293
rect 283 236 341 270
rect 283 83 375 236
rect 18 29 69 45
rect 103 19 119 53
rect 153 19 169 53
rect 409 55 443 327
rect 522 325 581 351
rect 556 317 581 325
rect 556 291 615 317
rect 522 275 615 291
rect 477 215 547 237
rect 477 181 489 215
rect 523 181 547 215
rect 477 163 547 181
rect 477 129 500 163
rect 534 129 547 163
rect 477 113 547 129
rect 581 157 615 275
rect 649 231 683 387
rect 717 419 751 435
rect 798 401 814 435
rect 848 401 864 435
rect 898 419 932 435
rect 717 367 751 385
rect 991 411 1011 445
rect 1045 411 1065 445
rect 991 395 1065 411
rect 1099 437 1133 453
rect 898 367 932 385
rect 717 333 932 367
rect 1099 361 1133 403
rect 1180 444 1354 453
rect 1180 410 1196 444
rect 1230 410 1354 444
rect 1180 385 1354 410
rect 1388 445 1438 487
rect 1422 411 1438 445
rect 1542 445 1608 487
rect 1388 395 1438 411
rect 1472 419 1506 435
rect 1021 327 1133 361
rect 1021 299 1055 327
rect 755 265 771 299
rect 805 265 1055 299
rect 1194 317 1205 351
rect 1239 325 1286 351
rect 1194 293 1236 317
rect 649 211 987 231
rect 649 197 953 211
rect 581 123 602 157
rect 636 123 652 157
rect 581 113 652 123
rect 686 55 720 197
rect 761 147 857 163
rect 795 113 833 147
rect 891 129 919 163
rect 953 161 987 177
rect 867 113 919 129
rect 1021 127 1055 265
rect 203 29 237 45
rect 103 -23 169 19
rect 309 15 325 49
rect 359 15 375 49
rect 409 21 458 55
rect 492 21 508 55
rect 549 21 565 55
rect 599 21 720 55
rect 895 53 961 69
rect 309 -23 375 15
rect 895 19 911 53
rect 945 19 961 53
rect 895 -23 961 19
rect 1003 49 1055 127
rect 1093 291 1236 293
rect 1270 291 1286 325
rect 1320 309 1354 385
rect 1542 411 1558 445
rect 1592 411 1608 445
rect 1667 445 1701 487
rect 1472 377 1506 385
rect 1667 377 1701 411
rect 1472 343 1632 377
rect 1093 259 1228 291
rect 1320 275 1514 309
rect 1548 275 1564 309
rect 1093 151 1135 259
rect 1320 257 1354 275
rect 1093 117 1101 151
rect 1093 101 1135 117
rect 1169 215 1239 225
rect 1169 199 1205 215
rect 1169 165 1197 199
rect 1231 165 1239 181
rect 1169 101 1239 165
rect 1273 223 1354 257
rect 1273 67 1307 223
rect 1421 210 1529 241
rect 1598 219 1632 343
rect 1667 275 1701 343
rect 1743 437 1801 453
rect 1743 403 1751 437
rect 1785 403 1801 437
rect 1743 369 1801 403
rect 1743 335 1751 369
rect 1785 335 1801 369
rect 1743 301 1801 335
rect 1835 437 1869 487
rect 1835 369 1869 403
rect 1835 319 1869 335
rect 1911 437 1961 453
rect 1911 403 1919 437
rect 1953 403 1961 437
rect 1911 369 1961 403
rect 1911 335 1919 369
rect 1953 335 1961 369
rect 1743 267 1751 301
rect 1785 285 1801 301
rect 1911 301 1961 335
rect 2003 437 2037 487
rect 2003 369 2037 403
rect 2003 319 2037 335
rect 1911 285 1919 301
rect 1785 267 1919 285
rect 1953 285 1961 301
rect 1953 267 2088 285
rect 1743 251 2088 267
rect 1455 201 1529 210
rect 1341 173 1385 189
rect 1375 139 1385 173
rect 1421 167 1437 176
rect 1471 167 1529 201
rect 1341 133 1385 139
rect 1481 147 1529 167
rect 1341 99 1447 133
rect 1117 53 1307 67
rect 1003 15 1023 49
rect 1057 15 1073 49
rect 1117 19 1133 53
rect 1167 19 1307 53
rect 1117 11 1307 19
rect 1341 49 1379 65
rect 1341 15 1345 49
rect 1413 53 1447 99
rect 1515 113 1529 147
rect 1481 87 1529 113
rect 1563 217 1632 219
rect 1563 209 1969 217
rect 1563 175 1715 209
rect 1749 175 1783 209
rect 1817 175 1851 209
rect 1885 175 1919 209
rect 1953 175 1969 209
rect 1563 124 1628 175
rect 2006 141 2088 251
rect 1563 69 1627 124
rect 1413 35 1563 53
rect 1597 35 1627 69
rect 1413 19 1627 35
rect 1667 123 1701 139
rect 1667 55 1701 89
rect 1341 -23 1379 15
rect 1667 -23 1701 21
rect 1735 123 2088 141
rect 1735 89 1751 123
rect 1785 107 1919 123
rect 1785 89 1801 107
rect 1735 55 1801 89
rect 1903 89 1919 107
rect 1953 107 2088 123
rect 1953 89 1969 107
rect 1735 21 1751 55
rect 1785 21 1801 55
rect 1735 11 1801 21
rect 1835 55 1869 71
rect 1835 -23 1869 21
rect 1903 55 1969 89
rect 1903 21 1919 55
rect 1953 21 1969 55
rect 1903 11 1969 21
rect 2003 55 2037 71
rect 2003 -23 2037 21
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1133 -23
rect 1167 -57 1225 -23
rect 1259 -57 1317 -23
rect 1351 -57 1409 -23
rect 1443 -57 1501 -23
rect 1535 -57 1593 -23
rect 1627 -57 1685 -23
rect 1719 -57 1777 -23
rect 1811 -57 1869 -23
rect 1903 -57 1961 -23
rect 1995 -57 2053 -23
rect 2087 -57 2116 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 857 487 891 521
rect 949 487 983 521
rect 1041 487 1075 521
rect 1133 487 1167 521
rect 1225 487 1259 521
rect 1317 487 1351 521
rect 1409 487 1443 521
rect 1501 487 1535 521
rect 1593 487 1627 521
rect 1685 487 1719 521
rect 1777 487 1811 521
rect 1869 487 1903 521
rect 1961 487 1995 521
rect 2053 487 2087 521
rect 122 190 134 215
rect 134 190 156 215
rect 122 181 156 190
rect 203 335 237 351
rect 203 317 237 335
rect 581 317 615 351
rect 489 181 523 215
rect 1205 325 1239 351
rect 1205 317 1236 325
rect 1236 317 1239 325
rect 761 113 795 147
rect 833 129 857 147
rect 857 129 867 147
rect 833 113 867 129
rect 1205 199 1239 215
rect 1205 181 1231 199
rect 1231 181 1239 199
rect 1421 201 1455 210
rect 1421 176 1437 201
rect 1437 176 1455 201
rect 1481 113 1515 147
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
rect 857 -57 891 -23
rect 949 -57 983 -23
rect 1041 -57 1075 -23
rect 1133 -57 1167 -23
rect 1225 -57 1259 -23
rect 1317 -57 1351 -23
rect 1409 -57 1443 -23
rect 1501 -57 1535 -23
rect 1593 -57 1627 -23
rect 1685 -57 1719 -23
rect 1777 -57 1811 -23
rect 1869 -57 1903 -23
rect 1961 -57 1995 -23
rect 2053 -57 2087 -23
<< metal1 >>
rect 0 521 2116 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1133 521
rect 1167 487 1225 521
rect 1259 487 1317 521
rect 1351 487 1409 521
rect 1443 487 1501 521
rect 1535 487 1593 521
rect 1627 487 1685 521
rect 1719 487 1777 521
rect 1811 487 1869 521
rect 1903 487 1961 521
rect 1995 487 2053 521
rect 2087 487 2116 521
rect 0 456 2116 487
rect 191 351 249 357
rect 191 317 203 351
rect 237 348 249 351
rect 569 351 627 357
rect 569 348 581 351
rect 237 320 581 348
rect 237 317 249 320
rect 191 311 249 317
rect 569 317 581 320
rect 615 348 627 351
rect 1193 351 1251 357
rect 1193 348 1205 351
rect 615 320 1205 348
rect 615 317 627 320
rect 569 311 627 317
rect 1193 317 1205 320
rect 1239 317 1251 351
rect 1193 311 1251 317
rect 110 215 168 221
rect 110 181 122 215
rect 156 212 168 215
rect 477 215 535 221
rect 477 212 489 215
rect 156 184 489 212
rect 156 181 168 184
rect 110 175 168 181
rect 477 181 489 184
rect 523 212 535 215
rect 1193 215 1251 221
rect 1193 212 1205 215
rect 523 184 1205 212
rect 523 181 535 184
rect 477 175 535 181
rect 1193 181 1205 184
rect 1239 181 1251 215
rect 1193 175 1251 181
rect 1409 210 1467 216
rect 1409 176 1421 210
rect 1455 176 1467 210
rect 1409 153 1467 176
rect 749 147 879 153
rect 749 113 761 147
rect 795 113 833 147
rect 867 144 879 147
rect 1409 147 1527 153
rect 1409 144 1481 147
rect 867 116 1481 144
rect 867 113 879 116
rect 749 107 879 113
rect 1469 113 1481 116
rect 1515 113 1527 147
rect 1469 107 1527 113
rect 0 -23 2116 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1133 -23
rect 1167 -57 1225 -23
rect 1259 -57 1317 -23
rect 1351 -57 1409 -23
rect 1443 -57 1501 -23
rect 1535 -57 1593 -23
rect 1627 -57 1685 -23
rect 1719 -57 1777 -23
rect 1811 -57 1869 -23
rect 1903 -57 1961 -23
rect 1995 -57 2053 -23
rect 2087 -57 2116 -23
rect 0 -88 2116 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 dfrtp_4
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 2042 181 2076 215 0 FreeSans 400 0 0 0 Q
port 11 nsew
flabel locali s 2042 249 2076 283 0 FreeSans 400 0 0 0 Q
port 11 nsew
flabel locali s 1481 113 1515 147 0 FreeSans 400 0 0 0 RESET_B
port 9 nsew
flabel locali s 305 249 339 283 0 FreeSans 400 0 0 0 D
port 8 nsew
flabel locali s 30 249 64 283 0 FreeSans 400 0 0 0 CLK
port 7 nsew
flabel locali s 30 181 64 215 0 FreeSans 400 0 0 0 CLK
port 7 nsew
flabel locali s 1481 181 1515 215 0 FreeSans 400 0 0 0 RESET_B
port 9 nsew
<< properties >>
string FIXED_BBOX 0 -40 2116 504
string path 48.300 12.600 50.600 12.600 
<< end >>
