magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 774 542
<< pwell >>
rect 17 -19 707 163
rect 29 -57 63 -19
<< scnmos >>
rect 95 7 125 137
rect 192 53 222 137
rect 418 7 448 137
rect 514 7 544 137
rect 598 7 628 137
<< scpmoshvt >>
rect 79 257 109 457
rect 192 257 222 341
rect 418 257 448 457
rect 514 257 544 457
rect 586 257 616 457
<< ndiff >>
rect 43 109 95 137
rect 43 75 51 109
rect 85 75 95 109
rect 43 7 95 75
rect 125 109 192 137
rect 125 75 142 109
rect 176 75 192 109
rect 125 53 192 75
rect 222 109 274 137
rect 222 75 232 109
rect 266 75 274 109
rect 222 53 274 75
rect 366 91 418 137
rect 366 57 374 91
rect 408 57 418 91
rect 125 7 177 53
rect 366 7 418 57
rect 448 123 514 137
rect 448 89 470 123
rect 504 89 514 123
rect 448 55 514 89
rect 448 21 470 55
rect 504 21 514 55
rect 448 7 514 21
rect 544 55 598 137
rect 544 21 554 55
rect 588 21 598 55
rect 544 7 598 21
rect 628 123 681 137
rect 628 89 638 123
rect 672 89 681 123
rect 628 55 681 89
rect 628 21 638 55
rect 672 21 681 55
rect 628 7 681 21
<< pdiff >>
rect 27 442 79 457
rect 27 408 35 442
rect 69 408 79 442
rect 27 374 79 408
rect 27 340 35 374
rect 69 340 79 374
rect 27 306 79 340
rect 27 272 35 306
rect 69 272 79 306
rect 27 257 79 272
rect 109 435 177 457
rect 109 401 135 435
rect 169 401 177 435
rect 109 341 177 401
rect 358 437 418 457
rect 358 403 366 437
rect 400 403 418 437
rect 109 257 192 341
rect 222 299 278 341
rect 222 265 232 299
rect 266 265 278 299
rect 222 257 278 265
rect 358 257 418 403
rect 448 437 514 457
rect 448 403 470 437
rect 504 403 514 437
rect 448 369 514 403
rect 448 335 470 369
rect 504 335 514 369
rect 448 301 514 335
rect 448 267 470 301
rect 504 267 514 301
rect 448 257 514 267
rect 544 257 586 457
rect 616 437 672 457
rect 616 403 626 437
rect 660 403 672 437
rect 616 369 672 403
rect 616 335 626 369
rect 660 335 672 369
rect 616 301 672 335
rect 616 267 626 301
rect 660 267 672 301
rect 616 257 672 267
<< ndiffc >>
rect 51 75 85 109
rect 142 75 176 109
rect 232 75 266 109
rect 374 57 408 91
rect 470 89 504 123
rect 470 21 504 55
rect 554 21 588 55
rect 638 89 672 123
rect 638 21 672 55
<< pdiffc >>
rect 35 408 69 442
rect 35 340 69 374
rect 35 272 69 306
rect 135 401 169 435
rect 366 403 400 437
rect 232 265 266 299
rect 470 403 504 437
rect 470 335 504 369
rect 470 267 504 301
rect 626 403 660 437
rect 626 335 660 369
rect 626 267 660 301
<< poly >>
rect 79 457 109 483
rect 418 457 448 483
rect 514 457 544 483
rect 586 457 616 483
rect 192 341 222 367
rect 79 225 109 257
rect 192 225 222 257
rect 418 225 448 257
rect 514 225 544 257
rect 79 209 146 225
rect 79 175 102 209
rect 136 175 146 209
rect 79 159 146 175
rect 192 209 254 225
rect 192 175 210 209
rect 244 175 254 209
rect 192 159 254 175
rect 296 209 448 225
rect 296 175 306 209
rect 340 175 448 209
rect 296 159 448 175
rect 490 209 544 225
rect 490 175 500 209
rect 534 175 544 209
rect 490 159 544 175
rect 586 225 616 257
rect 586 209 656 225
rect 586 175 606 209
rect 640 175 656 209
rect 586 159 656 175
rect 95 137 125 159
rect 192 137 222 159
rect 418 137 448 159
rect 514 137 544 159
rect 598 137 628 159
rect 192 27 222 53
rect 95 -19 125 7
rect 418 -19 448 7
rect 514 -19 544 7
rect 598 -19 628 7
<< polycont >>
rect 102 175 136 209
rect 210 175 244 209
rect 306 175 340 209
rect 500 175 534 209
rect 606 175 640 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 17 442 85 453
rect 17 408 35 442
rect 69 408 85 442
rect 17 374 85 408
rect 119 435 201 487
rect 119 401 135 435
rect 169 401 201 435
rect 350 437 416 487
rect 350 403 366 437
rect 400 403 416 437
rect 450 437 515 453
rect 450 403 470 437
rect 504 403 515 437
rect 17 340 35 374
rect 69 340 85 374
rect 450 369 515 403
rect 450 367 470 369
rect 17 306 85 340
rect 17 272 35 306
rect 69 272 85 306
rect 17 256 85 272
rect 119 335 470 367
rect 504 335 515 369
rect 119 333 515 335
rect 17 125 68 256
rect 119 225 172 333
rect 374 301 515 333
rect 215 265 232 299
rect 266 265 340 299
rect 102 209 172 225
rect 136 175 172 209
rect 102 159 172 175
rect 206 209 272 225
rect 206 175 210 209
rect 244 175 272 209
rect 206 159 272 175
rect 306 209 340 265
rect 306 125 340 175
rect 17 109 89 125
rect 17 75 51 109
rect 85 75 89 109
rect 17 50 89 75
rect 142 109 176 125
rect 142 -23 176 75
rect 232 109 340 125
rect 266 91 340 109
rect 374 267 470 301
rect 504 267 515 301
rect 610 437 676 487
rect 610 403 626 437
rect 660 403 676 437
rect 610 369 676 403
rect 610 335 626 369
rect 660 335 676 369
rect 610 301 676 335
rect 610 267 626 301
rect 660 267 676 301
rect 374 251 515 267
rect 374 91 408 251
rect 442 209 556 217
rect 442 175 500 209
rect 534 175 556 209
rect 590 209 719 217
rect 590 175 606 209
rect 640 175 719 209
rect 232 50 266 75
rect 374 11 408 57
rect 454 123 688 141
rect 454 89 470 123
rect 504 107 638 123
rect 504 89 520 107
rect 454 55 520 89
rect 622 89 638 107
rect 672 89 688 123
rect 454 21 470 55
rect 504 21 520 55
rect 454 11 520 21
rect 554 55 588 71
rect 554 -23 588 21
rect 622 55 688 89
rect 622 21 638 55
rect 672 21 688 55
rect 622 14 688 21
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
<< metal1 >>
rect 0 521 736 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 0 456 736 487
rect 0 -23 736 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
rect 0 -88 736 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 o21ba_1
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 213 181 247 215 0 FreeSans 400 0 0 0 B1_N
port 7 nsew
flabel locali s 673 181 707 215 0 FreeSans 400 0 0 0 A1
port 8 nsew
flabel locali s 29 385 63 419 0 FreeSans 400 0 0 0 X
port 10 nsew
flabel locali s 489 181 523 215 0 FreeSans 400 0 0 0 A2
port 9 nsew
<< properties >>
string FIXED_BBOX 0 -40 736 504
string path 0.000 -1.000 18.400 -1.000 
<< end >>
