magic
tech sky130B
magscale 1 2
timestamp 1697659686
<< viali >>
rect 28179 2935 28219 2975
rect 28179 2836 28219 2876
rect 28181 2661 28221 2701
rect 28182 2562 28222 2602
rect 28185 2382 28225 2422
rect 28180 2287 28220 2327
rect 28185 2111 28225 2151
rect 28179 2011 28219 2051
rect 28180 1833 28220 1873
rect 28180 1736 28220 1776
rect 28179 1559 28219 1599
rect 28180 1462 28220 1502
rect 28186 1281 28226 1321
rect 28180 1185 28220 1225
rect 28183 1011 28223 1051
rect 28183 914 28223 954
rect 28185 734 28225 774
rect 28183 636 28223 676
<< metal1 >>
rect 27080 4112 27086 4175
rect 27149 4112 27155 4175
rect 27085 3511 27091 3595
rect 27175 3511 27181 3595
rect 636 3422 6538 3458
rect 636 2871 672 3422
rect -234 2835 769 2871
rect 2654 2836 2690 3422
rect 4578 2836 4614 3422
rect 6502 2836 6538 3422
rect 28173 2981 28225 2987
rect 27071 2892 27077 2976
rect 27161 2892 27167 2976
rect 28173 2923 28225 2929
rect 28173 2882 28225 2888
rect 28173 2824 28225 2830
rect 28175 2707 28227 2713
rect 28175 2649 28227 2655
rect 28176 2608 28228 2614
rect 28176 2550 28228 2556
rect 28179 2428 28231 2434
rect 28179 2370 28231 2376
rect 28174 2333 28226 2339
rect 28174 2275 28226 2281
rect -232 2110 626 2204
rect 8228 2112 8230 2200
rect 28179 2157 28231 2163
rect 28179 2099 28231 2105
rect 28173 2057 28225 2063
rect 28173 1999 28225 2005
rect 28174 1879 28226 1885
rect 28174 1821 28226 1827
rect 28174 1782 28226 1788
rect 28174 1724 28226 1730
rect -280 1572 578 1666
rect 28173 1605 28225 1611
rect 28173 1547 28225 1553
rect 28174 1508 28226 1514
rect 28174 1450 28226 1456
rect 28180 1327 28232 1333
rect 28180 1269 28232 1275
rect 28174 1231 28226 1237
rect 28174 1173 28226 1179
rect 28177 1057 28229 1063
rect 28177 999 28229 1005
rect 28177 960 28229 966
rect 28177 902 28229 908
rect 28179 780 28231 786
rect 28179 722 28231 728
rect 28177 682 28229 688
rect 28177 624 28229 630
rect 27913 342 28008 492
rect 28459 340 28554 490
<< via1 >>
rect 27086 4112 27149 4175
rect 27091 3511 27175 3595
rect 27077 2892 27161 2976
rect 28173 2975 28225 2981
rect 28173 2935 28179 2975
rect 28179 2935 28219 2975
rect 28219 2935 28225 2975
rect 28173 2929 28225 2935
rect 28173 2876 28225 2882
rect 28173 2836 28179 2876
rect 28179 2836 28219 2876
rect 28219 2836 28225 2876
rect 28173 2830 28225 2836
rect 28175 2701 28227 2707
rect 28175 2661 28181 2701
rect 28181 2661 28221 2701
rect 28221 2661 28227 2701
rect 28175 2655 28227 2661
rect 28176 2602 28228 2608
rect 28176 2562 28182 2602
rect 28182 2562 28222 2602
rect 28222 2562 28228 2602
rect 28176 2556 28228 2562
rect 28179 2422 28231 2428
rect 28179 2382 28185 2422
rect 28185 2382 28225 2422
rect 28225 2382 28231 2422
rect 28179 2376 28231 2382
rect 28174 2327 28226 2333
rect 28174 2287 28180 2327
rect 28180 2287 28220 2327
rect 28220 2287 28226 2327
rect 28174 2281 28226 2287
rect 28179 2151 28231 2157
rect 28179 2111 28185 2151
rect 28185 2111 28225 2151
rect 28225 2111 28231 2151
rect 28179 2105 28231 2111
rect 28173 2051 28225 2057
rect 28173 2011 28179 2051
rect 28179 2011 28219 2051
rect 28219 2011 28225 2051
rect 28173 2005 28225 2011
rect 28174 1873 28226 1879
rect 28174 1833 28180 1873
rect 28180 1833 28220 1873
rect 28220 1833 28226 1873
rect 28174 1827 28226 1833
rect 28174 1776 28226 1782
rect 28174 1736 28180 1776
rect 28180 1736 28220 1776
rect 28220 1736 28226 1776
rect 28174 1730 28226 1736
rect 28173 1599 28225 1605
rect 28173 1559 28179 1599
rect 28179 1559 28219 1599
rect 28219 1559 28225 1599
rect 28173 1553 28225 1559
rect 28174 1502 28226 1508
rect 28174 1462 28180 1502
rect 28180 1462 28220 1502
rect 28220 1462 28226 1502
rect 28174 1456 28226 1462
rect 28180 1321 28232 1327
rect 28180 1281 28186 1321
rect 28186 1281 28226 1321
rect 28226 1281 28232 1321
rect 28180 1275 28232 1281
rect 28174 1225 28226 1231
rect 28174 1185 28180 1225
rect 28180 1185 28220 1225
rect 28220 1185 28226 1225
rect 28174 1179 28226 1185
rect 28177 1051 28229 1057
rect 28177 1011 28183 1051
rect 28183 1011 28223 1051
rect 28223 1011 28229 1051
rect 28177 1005 28229 1011
rect 28177 954 28229 960
rect 28177 914 28183 954
rect 28183 914 28223 954
rect 28223 914 28229 954
rect 28177 908 28229 914
rect 28179 774 28231 780
rect 28179 734 28185 774
rect 28185 734 28225 774
rect 28225 734 28231 774
rect 28179 728 28231 734
rect 28177 676 28229 682
rect 28177 636 28183 676
rect 28183 636 28223 676
rect 28223 636 28229 676
rect 28177 630 28229 636
<< metal2 >>
rect 27071 5310 27875 5399
rect 27079 4696 27750 4772
rect 27086 4175 27149 4181
rect 27149 4112 27646 4175
rect 27086 4106 27149 4112
rect 3020 3666 3080 3675
rect 3020 3597 3080 3606
rect 3031 3515 3069 3597
rect 27091 3595 27175 3601
rect 2451 3477 8211 3515
rect 27175 3511 27550 3595
rect 27091 3505 27175 3511
rect 2451 2875 2489 3477
rect 2321 2837 2489 2875
rect 4361 2873 4399 3477
rect 6245 2875 6283 3477
rect 4243 2835 4399 2873
rect 6163 2837 6283 2875
rect 8173 2873 8211 3477
rect 27077 2976 27161 2982
rect 27161 2892 27438 2976
rect 27077 2886 27161 2892
rect 8095 2835 8211 2873
rect 27093 2313 27325 2395
rect -232 1504 7194 1545
rect 27095 1325 27176 1801
rect 27243 1603 27325 2313
rect 27354 1877 27438 2892
rect 27466 2156 27550 3511
rect 27583 2424 27646 4112
rect 27674 2704 27750 4696
rect 27786 2980 27875 5310
rect 28167 2980 28173 2981
rect 27786 2929 28173 2980
rect 28225 2929 28231 2981
rect 27786 2928 27875 2929
rect 28167 2830 28173 2882
rect 28225 2873 28231 2882
rect 28225 2839 28662 2873
rect 28225 2830 28231 2839
rect 28169 2704 28175 2707
rect 27674 2657 28175 2704
rect 27674 2656 27750 2657
rect 28169 2655 28175 2657
rect 28227 2655 28233 2707
rect 28170 2556 28176 2608
rect 28228 2599 28234 2608
rect 28228 2565 28659 2599
rect 28228 2556 28234 2565
rect 28173 2424 28179 2428
rect 27583 2381 28179 2424
rect 27675 2380 28179 2381
rect 28173 2376 28179 2380
rect 28231 2376 28237 2428
rect 28168 2281 28174 2333
rect 28226 2324 28232 2333
rect 28226 2290 28660 2324
rect 28226 2281 28232 2290
rect 28173 2156 28179 2157
rect 27466 2105 28179 2156
rect 28231 2105 28237 2157
rect 27466 2104 27550 2105
rect 28167 2005 28173 2057
rect 28225 2048 28231 2057
rect 28225 2014 28662 2048
rect 28225 2005 28231 2014
rect 28168 1877 28174 1879
rect 27354 1829 28174 1877
rect 28168 1827 28174 1829
rect 28226 1827 28232 1879
rect 28168 1730 28174 1782
rect 28226 1773 28232 1782
rect 28226 1739 28663 1773
rect 28226 1730 28232 1739
rect 28167 1603 28173 1605
rect 27243 1555 28173 1603
rect 27243 1552 27325 1555
rect 28167 1553 28173 1555
rect 28225 1553 28231 1605
rect 28168 1456 28174 1508
rect 28226 1499 28232 1508
rect 28226 1465 28660 1499
rect 28226 1456 28232 1465
rect 28174 1325 28180 1327
rect 27095 1277 28180 1325
rect 27095 1276 27176 1277
rect 28174 1275 28180 1277
rect 28232 1275 28238 1327
rect 28168 1179 28174 1231
rect 28226 1222 28232 1231
rect 28226 1188 28660 1222
rect 28226 1179 28232 1188
rect 27094 1052 27167 1167
rect 28171 1052 28177 1057
rect 27094 1009 28177 1052
rect 27094 994 27167 1009
rect 28171 1005 28177 1009
rect 28229 1005 28235 1057
rect 28171 908 28177 960
rect 28229 951 28235 960
rect 28229 917 28662 951
rect 28229 908 28235 917
rect 27087 775 27150 786
rect 28173 775 28179 780
rect 27087 733 28179 775
rect 27087 525 27150 733
rect 28173 728 28179 733
rect 28231 728 28237 780
rect 28171 630 28177 682
rect 28229 673 28235 682
rect 28229 639 28662 673
rect 28229 630 28235 639
<< via2 >>
rect 3020 3606 3080 3666
<< metal3 >>
rect 2998 3671 3098 3686
rect 2998 3601 3015 3671
rect 3085 3601 3098 3671
rect 2998 3582 3098 3601
<< via3 >>
rect 3015 3666 3085 3671
rect 3015 3606 3020 3666
rect 3020 3606 3080 3666
rect 3080 3606 3085 3666
rect 3015 3601 3085 3606
<< metal4 >>
rect 3020 3672 3080 3794
rect 3014 3671 3086 3672
rect 3014 3601 3015 3671
rect 3085 3601 3086 3671
rect 3014 3600 3086 3601
use carray  carray_0
timestamp 1697065033
transform 1 0 -62 0 1 5400
box 62 -5400 27238 480
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1693170804
transform 0 1 27963 1 0 2261
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1693170804
transform 0 1 27963 1 0 2535
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_2
timestamp 1693170804
transform 0 1 27963 1 0 2810
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_3
timestamp 1693170804
transform 0 1 27963 1 0 1711
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_4
timestamp 1693170804
transform 0 1 27963 1 0 1160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_5
timestamp 1693170804
transform 0 1 27963 1 0 1435
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_6
timestamp 1693170804
transform 0 1 27963 1 0 886
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_7
timestamp 1693170804
transform 0 1 27963 1 0 611
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_8
timestamp 1693170804
transform 0 1 27963 1 0 1986
box -38 -48 314 592
use sky130_fd_sc_hd__tap_2  sky130_fd_sc_hd__tap_2_0
timestamp 1693170804
transform 0 1 27963 -1 0 614
box -38 -48 222 592
use sky130_fd_sc_hd__tap_2  sky130_fd_sc_hd__tap_2_1
timestamp 1693170804
transform 0 1 27963 -1 0 3267
box -38 -48 222 592
use sky130_fd_sc_hd__tap_2  sky130_fd_sc_hd__tap_2_2
timestamp 1693170804
transform 1 0 428 0 1 1616
box -38 -48 222 592
use sky130_fd_sc_hd__tap_2  sky130_fd_sc_hd__tap_2_3
timestamp 1693170804
transform 1 0 8304 0 1 1616
box -38 -48 222 592
use sw_top  sw_top_0
timestamp 1697571680
transform 1 0 6753 0 1 2396
box -410 -892 1590 1027
use sw_top  sw_top_1
timestamp 1697571680
transform 1 0 4830 0 1 2396
box -410 -892 1590 1027
use sw_top  sw_top_2
timestamp 1697571680
transform 1 0 984 0 1 2396
box -410 -892 1590 1027
use sw_top  sw_top_3
timestamp 1697571680
transform 1 0 2907 0 1 2396
box -410 -892 1590 1027
<< labels >>
flabel metal2 -232 1504 -191 1545 0 FreeSans 800 0 0 0 sample
port 11 nsew
flabel metal1 -224 2835 -188 2871 0 FreeSans 800 0 0 0 vin
port 9 nsew
flabel metal2 2451 3477 8211 3515 0 FreeSans 1600 0 0 0 out
port 12 nsew
flabel metal1 s -232 2110 -138 2204 0 FreeSans 640 0 0 0 vdd
port 10 nsew
flabel metal1 28459 340 28554 490 0 FreeSans 800 0 0 0 vdd
port 10 nsew
flabel metal2 28229 639 28662 673 0 FreeSans 800 0 0 0 dum
port 8 nsew
flabel metal2 28229 917 28662 951 0 FreeSans 800 0 0 0 ctl0
port 0 nsew
flabel metal2 28226 1188 28660 1222 0 FreeSans 800 0 0 0 ctl1
port 1 nsew
flabel metal2 28226 1465 28660 1499 0 FreeSans 800 0 0 0 ctl2
port 2 nsew
flabel metal2 28226 1739 28663 1773 0 FreeSans 800 0 0 0 ctl3
port 3 nsew
flabel metal2 28225 2014 28662 2048 0 FreeSans 800 0 0 0 ctl4
port 4 nsew
flabel metal2 28226 2290 28660 2324 0 FreeSans 800 0 0 0 ctl5
port 5 nsew
flabel metal2 28228 2565 28659 2599 0 FreeSans 800 0 0 0 ctl6
port 6 nsew
flabel metal2 28225 2839 28662 2873 0 FreeSans 800 0 0 0 ctl7
port 7 nsew
flabel metal1 27913 342 28008 492 0 FreeSans 800 0 0 0 vss
port 13 nsew
flabel metal1 -280 1572 578 1666 0 FreeSans 800 0 0 0 vss
port 13 nsew
<< end >>
