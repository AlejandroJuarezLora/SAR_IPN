magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 498 542
<< pwell >>
rect 211 117 397 163
rect 30 -19 397 117
rect 30 -23 63 -19
rect 29 -57 63 -23
<< scnmos >>
rect 108 7 138 91
rect 192 7 222 91
rect 289 7 319 137
<< scpmoshvt >>
rect 120 257 150 341
rect 192 257 222 341
rect 289 257 319 457
<< ndiff >>
rect 237 91 289 137
rect 56 63 108 91
rect 56 29 64 63
rect 98 29 108 63
rect 56 7 108 29
rect 138 63 192 91
rect 138 29 148 63
rect 182 29 192 63
rect 138 7 192 29
rect 222 63 289 91
rect 222 29 244 63
rect 278 29 289 63
rect 222 7 289 29
rect 319 123 371 137
rect 319 89 329 123
rect 363 89 371 123
rect 319 55 371 89
rect 319 21 329 55
rect 363 21 371 55
rect 319 7 371 21
<< pdiff >>
rect 237 429 289 457
rect 237 395 245 429
rect 279 395 289 429
rect 237 361 289 395
rect 237 341 245 361
rect 68 309 120 341
rect 68 275 76 309
rect 110 275 120 309
rect 68 257 120 275
rect 150 257 192 341
rect 222 327 245 341
rect 279 327 289 361
rect 222 257 289 327
rect 319 445 387 457
rect 319 411 345 445
rect 379 411 387 445
rect 319 377 387 411
rect 319 343 345 377
rect 379 343 387 377
rect 319 257 387 343
<< ndiffc >>
rect 64 29 98 63
rect 148 29 182 63
rect 244 29 278 63
rect 329 89 363 123
rect 329 21 363 55
<< pdiffc >>
rect 245 395 279 429
rect 76 275 110 309
rect 245 327 279 361
rect 345 411 379 445
rect 345 343 379 377
<< poly >>
rect 289 457 319 483
rect 120 341 150 367
rect 192 341 222 367
rect 120 225 150 257
rect 50 209 150 225
rect 50 175 66 209
rect 100 175 150 209
rect 50 159 150 175
rect 192 225 222 257
rect 289 225 319 257
rect 192 209 246 225
rect 192 175 202 209
rect 236 175 246 209
rect 192 159 246 175
rect 289 209 355 225
rect 289 175 305 209
rect 339 175 355 209
rect 289 159 355 175
rect 108 91 138 159
rect 192 91 222 159
rect 289 137 319 159
rect 108 -19 138 7
rect 192 -19 222 7
rect 289 -19 319 7
<< polycont >>
rect 66 175 100 209
rect 202 175 236 209
rect 305 175 339 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 229 429 295 487
rect 229 395 245 429
rect 279 395 295 429
rect 229 361 295 395
rect 54 309 132 328
rect 229 327 245 361
rect 279 327 295 361
rect 329 445 436 453
rect 329 411 345 445
rect 379 411 436 445
rect 329 377 436 411
rect 329 343 345 377
rect 379 343 436 377
rect 329 329 436 343
rect 54 275 76 309
rect 110 293 132 309
rect 110 275 339 293
rect 54 259 339 275
rect 29 209 100 225
rect 29 175 66 209
rect 29 113 100 175
rect 134 79 168 259
rect 202 209 255 225
rect 236 175 255 209
rect 202 113 255 175
rect 305 209 339 259
rect 305 159 339 175
rect 373 125 436 329
rect 313 123 436 125
rect 313 89 329 123
rect 363 89 436 123
rect 50 63 98 79
rect 50 29 64 63
rect 50 -23 98 29
rect 134 63 190 79
rect 134 29 148 63
rect 182 29 190 63
rect 134 13 190 29
rect 236 63 279 79
rect 236 29 244 63
rect 278 29 279 63
rect 236 -23 279 29
rect 313 55 436 89
rect 313 21 329 55
rect 363 21 436 55
rect 313 11 436 21
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
<< metal1 >>
rect 0 521 460 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 0 456 460 487
rect 0 -23 460 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
rect 0 -88 460 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 or2_1
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 213 181 247 215 0 FreeSans 200 0 0 0 A
port 8 nsew
flabel locali s 397 317 431 351 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 29 181 63 215 0 FreeSans 200 0 0 0 B
port 9 nsew
<< properties >>
string FIXED_BBOX 0 -40 460 504
string path 0.000 -1.000 11.500 -1.000 
<< end >>
