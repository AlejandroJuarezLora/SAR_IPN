VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO comparator
  CLASS BLOCK ;
  FOREIGN comparator ;
  ORIGIN 0.000 0.200 ;
  SIZE 50.520 BY 20.300 ;
  PIN trim_3
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 4.335 15.405 4.505 15.735 ;
        RECT 4.335 14.815 4.505 15.145 ;
        RECT 4.335 14.225 4.505 14.555 ;
        RECT 4.335 13.635 4.505 13.965 ;
      LAYER mcon ;
        RECT 4.335 15.485 4.505 15.655 ;
        RECT 4.335 14.895 4.505 15.065 ;
        RECT 4.335 14.305 4.505 14.475 ;
        RECT 4.335 13.715 4.505 13.885 ;
      LAYER met1 ;
        RECT 4.305 14.835 4.535 15.715 ;
        RECT 3.605 14.535 4.535 14.835 ;
        RECT 4.305 13.655 4.535 14.535 ;
      LAYER via ;
        RECT 3.665 14.555 3.925 14.815 ;
        RECT 3.985 14.555 4.245 14.815 ;
      LAYER met2 ;
        RECT 3.655 14.835 4.255 14.885 ;
        RECT 0.700 14.535 4.255 14.835 ;
        RECT 0.700 -0.200 1.000 14.535 ;
        RECT 3.655 14.485 4.255 14.535 ;
    END
  END trim_3
  PIN trim_2
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 4.335 12.090 4.505 12.420 ;
        RECT 4.335 11.500 4.505 11.830 ;
      LAYER mcon ;
        RECT 4.335 12.170 4.505 12.340 ;
        RECT 4.335 11.580 4.505 11.750 ;
      LAYER met1 ;
        RECT 4.305 12.110 4.535 12.400 ;
        RECT 3.605 11.810 4.535 12.110 ;
        RECT 4.305 11.520 4.535 11.810 ;
      LAYER via ;
        RECT 3.665 11.830 3.925 12.090 ;
        RECT 3.985 11.830 4.245 12.090 ;
      LAYER met2 ;
        RECT 3.655 12.110 4.255 12.160 ;
        RECT 1.300 11.810 4.255 12.110 ;
        RECT 1.300 -0.200 1.600 11.810 ;
        RECT 3.655 11.760 4.255 11.810 ;
    END
  END trim_2
  PIN trim_0
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 4.335 9.955 4.505 10.285 ;
      LAYER mcon ;
        RECT 4.335 10.035 4.505 10.205 ;
      LAYER met1 ;
        RECT 3.605 10.430 4.535 10.730 ;
        RECT 4.305 9.975 4.535 10.430 ;
      LAYER via ;
        RECT 3.665 10.450 3.925 10.710 ;
        RECT 3.985 10.450 4.245 10.710 ;
      LAYER met2 ;
        RECT 3.655 10.730 4.255 10.780 ;
        RECT 1.900 10.430 4.255 10.730 ;
        RECT 1.900 -0.200 2.200 10.430 ;
        RECT 3.655 10.380 4.255 10.430 ;
    END
  END trim_0
  PIN trim_1
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 4.335 9.365 4.505 9.695 ;
      LAYER mcon ;
        RECT 4.335 9.445 4.505 9.615 ;
      LAYER met1 ;
        RECT 4.305 9.220 4.535 9.675 ;
        RECT 3.605 8.920 4.535 9.220 ;
      LAYER via ;
        RECT 3.665 8.940 3.925 9.200 ;
        RECT 3.985 8.940 4.245 9.200 ;
      LAYER met2 ;
        RECT 3.655 9.220 4.255 9.270 ;
        RECT 2.500 8.920 4.255 9.220 ;
        RECT 2.500 -0.200 2.800 8.920 ;
        RECT 3.655 8.870 4.255 8.920 ;
    END
  END trim_1
  PIN trim_4
    ANTENNAGATEAREA 2.400000 ;
    PORT
      LAYER li1 ;
        RECT 4.335 7.820 4.505 8.150 ;
        RECT 4.335 7.230 4.505 7.560 ;
        RECT 4.335 6.640 4.505 6.970 ;
        RECT 4.335 6.050 4.505 6.380 ;
        RECT 4.335 5.460 4.505 5.790 ;
        RECT 4.335 4.870 4.505 5.200 ;
        RECT 4.335 4.280 4.505 4.610 ;
        RECT 4.335 3.690 4.505 4.020 ;
      LAYER mcon ;
        RECT 4.335 7.900 4.505 8.070 ;
        RECT 4.335 7.310 4.505 7.480 ;
        RECT 4.335 6.720 4.505 6.890 ;
        RECT 4.335 6.130 4.505 6.300 ;
        RECT 4.335 5.540 4.505 5.710 ;
        RECT 4.335 4.950 4.505 5.120 ;
        RECT 4.335 4.360 4.505 4.530 ;
        RECT 4.335 3.770 4.505 3.940 ;
      LAYER met1 ;
        RECT 4.305 6.070 4.535 8.130 ;
        RECT 3.605 5.770 4.535 6.070 ;
        RECT 4.305 3.710 4.535 5.770 ;
      LAYER via ;
        RECT 3.665 5.790 3.925 6.050 ;
        RECT 3.985 5.790 4.245 6.050 ;
      LAYER met2 ;
        RECT 3.655 6.070 4.255 6.120 ;
        RECT 3.100 5.770 4.255 6.070 ;
        RECT 3.100 -0.200 3.400 5.770 ;
        RECT 3.655 5.720 4.255 5.770 ;
    END
  END trim_4
  PIN trimb_4
    ANTENNAGATEAREA 2.400000 ;
    PORT
      LAYER li1 ;
        RECT 46.015 7.820 46.185 8.150 ;
        RECT 46.015 7.230 46.185 7.560 ;
        RECT 46.015 6.640 46.185 6.970 ;
        RECT 46.015 6.050 46.185 6.380 ;
        RECT 46.015 5.460 46.185 5.790 ;
        RECT 46.015 4.870 46.185 5.200 ;
        RECT 46.015 4.280 46.185 4.610 ;
        RECT 46.015 3.690 46.185 4.020 ;
      LAYER mcon ;
        RECT 46.015 7.900 46.185 8.070 ;
        RECT 46.015 7.310 46.185 7.480 ;
        RECT 46.015 6.720 46.185 6.890 ;
        RECT 46.015 6.130 46.185 6.300 ;
        RECT 46.015 5.540 46.185 5.710 ;
        RECT 46.015 4.950 46.185 5.120 ;
        RECT 46.015 4.360 46.185 4.530 ;
        RECT 46.015 3.770 46.185 3.940 ;
      LAYER met1 ;
        RECT 45.985 6.070 46.215 8.130 ;
        RECT 45.985 5.770 46.915 6.070 ;
        RECT 45.985 3.710 46.215 5.770 ;
      LAYER via ;
        RECT 46.275 5.790 46.535 6.050 ;
        RECT 46.595 5.790 46.855 6.050 ;
      LAYER met2 ;
        RECT 46.265 6.070 46.865 6.120 ;
        RECT 46.265 5.770 47.420 6.070 ;
        RECT 46.265 5.720 46.865 5.770 ;
        RECT 47.120 -0.200 47.420 5.770 ;
    END
  END trimb_4
  PIN trimb_1
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 46.015 9.365 46.185 9.695 ;
      LAYER mcon ;
        RECT 46.015 9.445 46.185 9.615 ;
      LAYER met1 ;
        RECT 45.985 9.220 46.215 9.675 ;
        RECT 45.985 8.920 46.915 9.220 ;
      LAYER via ;
        RECT 46.275 8.940 46.535 9.200 ;
        RECT 46.595 8.940 46.855 9.200 ;
      LAYER met2 ;
        RECT 46.265 9.220 46.865 9.270 ;
        RECT 46.265 8.920 48.020 9.220 ;
        RECT 46.265 8.870 46.865 8.920 ;
        RECT 47.720 -0.200 48.020 8.920 ;
    END
  END trimb_1
  PIN trimb_0
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 46.015 9.955 46.185 10.285 ;
      LAYER mcon ;
        RECT 46.015 10.035 46.185 10.205 ;
      LAYER met1 ;
        RECT 45.985 10.430 46.915 10.730 ;
        RECT 45.985 9.975 46.215 10.430 ;
      LAYER via ;
        RECT 46.275 10.450 46.535 10.710 ;
        RECT 46.595 10.450 46.855 10.710 ;
      LAYER met2 ;
        RECT 46.265 10.730 46.865 10.780 ;
        RECT 46.265 10.430 48.620 10.730 ;
        RECT 46.265 10.380 46.865 10.430 ;
        RECT 48.320 -0.200 48.620 10.430 ;
    END
  END trimb_0
  PIN trimb_2
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER li1 ;
        RECT 46.015 12.090 46.185 12.420 ;
        RECT 46.015 11.500 46.185 11.830 ;
      LAYER mcon ;
        RECT 46.015 12.170 46.185 12.340 ;
        RECT 46.015 11.580 46.185 11.750 ;
      LAYER met1 ;
        RECT 45.985 12.110 46.215 12.400 ;
        RECT 45.985 11.810 46.915 12.110 ;
        RECT 45.985 11.520 46.215 11.810 ;
      LAYER via ;
        RECT 46.275 11.830 46.535 12.090 ;
        RECT 46.595 11.830 46.855 12.090 ;
      LAYER met2 ;
        RECT 46.265 12.110 46.865 12.160 ;
        RECT 46.265 11.810 49.220 12.110 ;
        RECT 46.265 11.760 46.865 11.810 ;
        RECT 48.920 -0.200 49.220 11.810 ;
    END
  END trimb_2
  PIN trimb_3
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER li1 ;
        RECT 46.015 15.405 46.185 15.735 ;
        RECT 46.015 14.815 46.185 15.145 ;
        RECT 46.015 14.225 46.185 14.555 ;
        RECT 46.015 13.635 46.185 13.965 ;
      LAYER mcon ;
        RECT 46.015 15.485 46.185 15.655 ;
        RECT 46.015 14.895 46.185 15.065 ;
        RECT 46.015 14.305 46.185 14.475 ;
        RECT 46.015 13.715 46.185 13.885 ;
      LAYER met1 ;
        RECT 45.985 14.835 46.215 15.715 ;
        RECT 45.985 14.535 46.915 14.835 ;
        RECT 45.985 13.655 46.215 14.535 ;
      LAYER via ;
        RECT 46.275 14.555 46.535 14.815 ;
        RECT 46.595 14.555 46.855 14.815 ;
      LAYER met2 ;
        RECT 46.265 14.835 46.865 14.885 ;
        RECT 46.265 14.535 49.820 14.835 ;
        RECT 46.265 14.485 46.865 14.535 ;
        RECT 49.520 -0.200 49.820 14.535 ;
    END
  END trimb_3
  PIN outn
    ANTENNAGATEAREA 0.600000 ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER li1 ;
        RECT 21.825 15.685 21.995 16.725 ;
        RECT 24.590 15.685 24.760 16.725 ;
        RECT 25.395 15.300 25.725 15.470 ;
        RECT 25.980 9.135 26.310 9.305 ;
        RECT 23.995 7.925 24.165 8.965 ;
      LAYER mcon ;
        RECT 21.825 16.300 21.995 16.470 ;
        RECT 21.825 15.940 21.995 16.110 ;
        RECT 24.590 16.300 24.760 16.470 ;
        RECT 24.590 15.940 24.760 16.110 ;
        RECT 25.475 15.300 25.645 15.470 ;
        RECT 26.060 9.135 26.230 9.305 ;
        RECT 23.995 8.540 24.165 8.710 ;
        RECT 23.995 8.180 24.165 8.350 ;
      LAYER met1 ;
        RECT 21.795 16.345 22.025 16.705 ;
        RECT 22.825 16.345 23.125 16.545 ;
        RECT 24.560 16.345 24.790 16.705 ;
        RECT 21.795 16.045 24.790 16.345 ;
        RECT 21.795 15.705 22.025 16.045 ;
        RECT 22.825 15.845 23.125 16.045 ;
        RECT 24.560 15.705 24.790 16.045 ;
        RECT 25.415 15.270 26.260 15.500 ;
        RECT 26.030 14.250 26.260 15.270 ;
        RECT 25.995 13.550 26.295 14.250 ;
        RECT 26.030 13.525 26.260 13.550 ;
        RECT 23.460 12.680 26.260 12.910 ;
        RECT 22.620 12.135 23.320 12.170 ;
        RECT 23.460 12.135 23.690 12.680 ;
        RECT 26.030 12.375 26.260 12.680 ;
        RECT 22.620 11.905 23.690 12.135 ;
        RECT 22.620 11.870 23.320 11.905 ;
        RECT 25.995 11.675 26.295 12.375 ;
        RECT 25.995 9.335 26.295 10.035 ;
        RECT 26.000 9.105 26.290 9.335 ;
        RECT 23.965 8.645 24.195 8.945 ;
        RECT 22.825 7.945 24.195 8.645 ;
      LAYER via ;
        RECT 22.845 16.225 23.105 16.485 ;
        RECT 22.845 15.905 23.105 16.165 ;
        RECT 26.015 13.930 26.275 14.190 ;
        RECT 26.015 13.610 26.275 13.870 ;
        RECT 22.680 11.890 22.940 12.150 ;
        RECT 23.000 11.890 23.260 12.150 ;
        RECT 26.015 12.055 26.275 12.315 ;
        RECT 26.015 11.735 26.275 11.995 ;
        RECT 26.015 9.715 26.275 9.975 ;
        RECT 26.015 9.395 26.275 9.655 ;
        RECT 22.845 8.325 23.105 8.585 ;
        RECT 22.845 8.005 23.105 8.265 ;
      LAYER met2 ;
        RECT 22.775 12.220 23.175 16.495 ;
        RECT 25.995 14.200 26.295 14.250 ;
        RECT 25.945 13.600 26.345 14.200 ;
        RECT 25.995 12.325 26.295 13.600 ;
        RECT 22.670 11.820 23.270 12.220 ;
        RECT 22.775 -0.200 23.175 11.820 ;
        RECT 25.945 11.725 26.345 12.325 ;
        RECT 25.995 9.985 26.295 11.725 ;
        RECT 25.945 9.385 26.345 9.985 ;
    END
  END outn
  PIN outp
    ANTENNAGATEAREA 0.600000 ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER li1 ;
        RECT 25.770 15.685 25.940 16.725 ;
        RECT 28.485 15.685 28.655 16.725 ;
        RECT 24.805 15.300 25.135 15.470 ;
        RECT 24.210 9.135 24.540 9.305 ;
        RECT 26.355 7.925 26.525 8.965 ;
      LAYER mcon ;
        RECT 25.770 16.300 25.940 16.470 ;
        RECT 25.770 15.940 25.940 16.110 ;
        RECT 28.485 16.300 28.655 16.470 ;
        RECT 28.485 15.940 28.655 16.110 ;
        RECT 24.885 15.300 25.055 15.470 ;
        RECT 24.290 9.135 24.460 9.305 ;
        RECT 26.355 8.540 26.525 8.710 ;
        RECT 26.355 8.180 26.525 8.350 ;
      LAYER met1 ;
        RECT 25.740 16.345 25.970 16.705 ;
        RECT 27.395 16.345 27.695 16.545 ;
        RECT 28.455 16.345 28.685 16.705 ;
        RECT 25.740 16.045 28.685 16.345 ;
        RECT 25.740 15.705 25.970 16.045 ;
        RECT 27.395 15.845 27.695 16.045 ;
        RECT 28.455 15.705 28.685 16.045 ;
        RECT 24.260 15.270 25.115 15.500 ;
        RECT 24.260 14.250 24.490 15.270 ;
        RECT 24.225 13.550 24.525 14.250 ;
        RECT 24.225 11.675 24.525 12.375 ;
        RECT 27.200 12.135 27.900 12.170 ;
        RECT 26.830 11.905 27.900 12.135 ;
        RECT 24.260 11.370 24.490 11.675 ;
        RECT 26.830 11.370 27.060 11.905 ;
        RECT 27.200 11.870 27.900 11.905 ;
        RECT 24.260 11.140 27.060 11.370 ;
        RECT 24.225 9.335 24.525 10.035 ;
        RECT 24.230 9.105 24.520 9.335 ;
        RECT 26.325 8.645 26.555 8.945 ;
        RECT 26.325 7.945 27.695 8.645 ;
      LAYER via ;
        RECT 27.415 16.225 27.675 16.485 ;
        RECT 27.415 15.905 27.675 16.165 ;
        RECT 24.245 13.930 24.505 14.190 ;
        RECT 24.245 13.610 24.505 13.870 ;
        RECT 24.245 12.055 24.505 12.315 ;
        RECT 24.245 11.735 24.505 11.995 ;
        RECT 27.260 11.890 27.520 12.150 ;
        RECT 27.580 11.890 27.840 12.150 ;
        RECT 24.245 9.715 24.505 9.975 ;
        RECT 24.245 9.395 24.505 9.655 ;
        RECT 27.415 8.325 27.675 8.585 ;
        RECT 27.415 8.005 27.675 8.265 ;
      LAYER met2 ;
        RECT 24.225 14.200 24.525 14.250 ;
        RECT 24.175 13.600 24.575 14.200 ;
        RECT 24.225 12.325 24.525 13.600 ;
        RECT 24.175 11.725 24.575 12.325 ;
        RECT 27.345 12.220 27.745 16.495 ;
        RECT 27.250 11.820 27.850 12.220 ;
        RECT 24.225 9.985 24.525 11.725 ;
        RECT 24.175 9.385 24.575 9.985 ;
        RECT 27.345 -0.200 27.745 11.820 ;
    END
  END outp
  PIN clk
    ANTENNAGATEAREA 1.800000 ;
    PORT
      LAYER li1 ;
        RECT 20.860 15.300 21.190 15.470 ;
        RECT 21.450 15.300 21.780 15.470 ;
        RECT 28.700 15.300 29.030 15.470 ;
        RECT 29.290 15.300 29.620 15.470 ;
        RECT 24.800 4.435 25.130 4.605 ;
        RECT 25.390 4.435 25.720 4.605 ;
      LAYER mcon ;
        RECT 20.940 15.300 21.110 15.470 ;
        RECT 21.530 15.300 21.700 15.470 ;
        RECT 28.780 15.300 28.950 15.470 ;
        RECT 29.370 15.300 29.540 15.470 ;
        RECT 24.880 4.435 25.050 4.605 ;
        RECT 25.470 4.435 25.640 4.605 ;
      LAYER met1 ;
        RECT 20.880 15.270 21.800 15.500 ;
        RECT 28.720 15.270 29.640 15.500 ;
        RECT 21.205 11.665 21.435 15.270 ;
        RECT 20.080 11.435 21.435 11.665 ;
        RECT 29.055 11.665 29.285 15.270 ;
        RECT 29.055 11.435 30.440 11.665 ;
        RECT 20.080 8.645 20.310 11.435 ;
        RECT 30.210 8.645 30.440 11.435 ;
        RECT 20.045 7.945 20.345 8.645 ;
        RECT 30.175 7.945 30.475 8.645 ;
        RECT 20.045 4.980 20.345 5.680 ;
        RECT 30.175 4.980 30.475 5.680 ;
        RECT 20.080 4.635 20.310 4.980 ;
        RECT 30.210 4.635 30.440 4.980 ;
        RECT 20.080 4.405 30.440 4.635 ;
        RECT 25.110 2.240 25.410 4.405 ;
        RECT 17.560 1.940 25.410 2.240 ;
        RECT 17.560 -0.200 17.860 1.940 ;
      LAYER via ;
        RECT 20.065 8.325 20.325 8.585 ;
        RECT 20.065 8.005 20.325 8.265 ;
        RECT 30.195 8.325 30.455 8.585 ;
        RECT 30.195 8.005 30.455 8.265 ;
        RECT 20.065 5.360 20.325 5.620 ;
        RECT 20.065 5.040 20.325 5.300 ;
        RECT 30.195 5.360 30.455 5.620 ;
        RECT 30.195 5.040 30.455 5.300 ;
      LAYER met2 ;
        RECT 19.995 5.030 20.395 8.595 ;
        RECT 30.125 5.030 30.525 8.595 ;
    END
  END clk
  PIN vdd
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER li1 ;
        RECT 19.940 17.510 30.540 17.680 ;
        RECT 19.940 14.730 20.110 17.510 ;
        RECT 21.235 15.685 21.405 16.725 ;
        RECT 25.180 15.685 25.350 16.725 ;
        RECT 29.075 15.685 29.245 16.725 ;
        RECT 30.370 14.730 30.540 17.510 ;
        RECT 19.940 14.560 30.540 14.730 ;
      LAYER mcon ;
        RECT 22.510 17.510 22.680 17.680 ;
        RECT 22.870 17.510 23.040 17.680 ;
        RECT 23.230 17.510 23.400 17.680 ;
        RECT 23.590 17.510 23.760 17.680 ;
        RECT 26.730 17.510 26.900 17.680 ;
        RECT 27.090 17.510 27.260 17.680 ;
        RECT 27.450 17.510 27.620 17.680 ;
        RECT 27.810 17.510 27.980 17.680 ;
        RECT 21.235 16.300 21.405 16.470 ;
        RECT 21.235 15.940 21.405 16.110 ;
        RECT 25.180 16.300 25.350 16.470 ;
        RECT 25.180 15.940 25.350 16.110 ;
        RECT 29.075 16.300 29.245 16.470 ;
        RECT 29.075 15.940 29.245 16.110 ;
      LAYER met1 ;
        RECT 20.970 18.500 21.670 18.800 ;
        RECT 22.825 18.500 23.525 18.800 ;
        RECT 24.915 18.500 25.615 18.800 ;
        RECT 27.045 18.500 27.745 18.800 ;
        RECT 28.810 18.500 29.510 18.800 ;
        RECT 21.205 15.705 21.435 18.500 ;
        RECT 23.060 17.710 23.290 18.500 ;
        RECT 22.320 17.480 23.995 17.710 ;
        RECT 25.150 15.705 25.380 18.500 ;
        RECT 27.280 17.710 27.510 18.500 ;
        RECT 26.540 17.480 28.215 17.710 ;
        RECT 29.045 15.705 29.275 18.500 ;
      LAYER via ;
        RECT 21.030 18.520 21.290 18.780 ;
        RECT 21.350 18.520 21.610 18.780 ;
        RECT 22.885 18.520 23.145 18.780 ;
        RECT 23.205 18.520 23.465 18.780 ;
        RECT 24.975 18.520 25.235 18.780 ;
        RECT 25.295 18.520 25.555 18.780 ;
        RECT 27.105 18.520 27.365 18.780 ;
        RECT 27.425 18.520 27.685 18.780 ;
        RECT 28.870 18.520 29.130 18.780 ;
        RECT 29.190 18.520 29.450 18.780 ;
      LAYER met2 ;
        RECT 21.020 18.450 29.460 18.850 ;
      LAYER via2 ;
        RECT 24.925 18.510 25.205 18.790 ;
        RECT 25.325 18.510 25.605 18.790 ;
      LAYER met3 ;
        RECT 0.000 18.450 50.520 18.850 ;
        RECT 0.000 1.370 0.400 18.450 ;
        RECT 50.120 1.370 50.520 18.450 ;
        RECT 0.000 0.970 50.520 1.370 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 20.448900 ;
    PORT
      LAYER pwell ;
        RECT 3.630 16.235 6.520 16.665 ;
        RECT 3.630 3.185 4.060 16.235 ;
        RECT 6.090 3.185 6.520 16.235 ;
        RECT 44.000 16.235 46.890 16.665 ;
        RECT 23.180 9.585 27.340 10.015 ;
        RECT 23.180 7.615 23.610 9.585 ;
        RECT 26.910 7.615 27.340 9.585 ;
        RECT 23.180 7.185 27.340 7.615 ;
        RECT 23.670 6.145 26.850 6.575 ;
        RECT 23.670 4.250 24.100 6.145 ;
        RECT 26.420 4.250 26.850 6.145 ;
        RECT 23.670 3.820 26.850 4.250 ;
        RECT 3.630 2.755 6.520 3.185 ;
        RECT 44.000 3.185 44.430 16.235 ;
        RECT 46.460 3.185 46.890 16.235 ;
        RECT 44.000 2.755 46.890 3.185 ;
      LAYER li1 ;
        RECT 3.760 16.365 6.390 16.535 ;
        RECT 3.760 3.055 3.930 16.365 ;
        RECT 4.675 15.190 5.715 15.360 ;
        RECT 4.675 14.010 5.715 14.180 ;
        RECT 4.675 11.875 5.715 12.045 ;
        RECT 4.675 9.740 5.715 9.910 ;
        RECT 4.675 8.195 5.715 8.365 ;
        RECT 4.675 7.015 5.715 7.185 ;
        RECT 4.675 5.835 5.715 6.005 ;
        RECT 4.675 4.655 5.715 4.825 ;
        RECT 4.675 3.475 5.715 3.645 ;
        RECT 6.220 3.055 6.390 16.365 ;
        RECT 44.130 16.365 46.760 16.535 ;
        RECT 23.310 9.715 27.210 9.885 ;
        RECT 23.310 7.485 23.480 9.715 ;
        RECT 27.040 7.485 27.210 9.715 ;
        RECT 23.310 7.315 27.210 7.485 ;
        RECT 23.800 6.275 26.720 6.445 ;
        RECT 23.800 4.120 23.970 6.275 ;
        RECT 24.585 4.775 24.755 5.815 ;
        RECT 25.765 4.775 25.935 5.815 ;
        RECT 26.550 4.120 26.720 6.275 ;
        RECT 23.800 3.950 26.720 4.120 ;
        RECT 3.760 2.885 6.390 3.055 ;
        RECT 44.130 3.055 44.300 16.365 ;
        RECT 44.805 15.190 45.845 15.360 ;
        RECT 44.805 14.010 45.845 14.180 ;
        RECT 44.805 11.875 45.845 12.045 ;
        RECT 44.805 9.740 45.845 9.910 ;
        RECT 44.805 8.195 45.845 8.365 ;
        RECT 44.805 7.015 45.845 7.185 ;
        RECT 44.805 5.835 45.845 6.005 ;
        RECT 44.805 4.655 45.845 4.825 ;
        RECT 44.805 3.475 45.845 3.645 ;
        RECT 46.590 3.055 46.760 16.365 ;
        RECT 44.130 2.885 46.760 3.055 ;
      LAYER mcon ;
        RECT 5.025 16.365 5.195 16.535 ;
        RECT 5.385 16.365 5.555 16.535 ;
        RECT 4.930 15.190 5.100 15.360 ;
        RECT 5.290 15.190 5.460 15.360 ;
        RECT 4.930 14.010 5.100 14.180 ;
        RECT 5.290 14.010 5.460 14.180 ;
        RECT 4.930 11.875 5.100 12.045 ;
        RECT 5.290 11.875 5.460 12.045 ;
        RECT 4.930 9.740 5.100 9.910 ;
        RECT 5.290 9.740 5.460 9.910 ;
        RECT 4.930 8.195 5.100 8.365 ;
        RECT 5.290 8.195 5.460 8.365 ;
        RECT 4.930 7.015 5.100 7.185 ;
        RECT 5.290 7.015 5.460 7.185 ;
        RECT 4.930 5.835 5.100 6.005 ;
        RECT 5.290 5.835 5.460 6.005 ;
        RECT 4.930 4.655 5.100 4.825 ;
        RECT 5.290 4.655 5.460 4.825 ;
        RECT 4.930 3.475 5.100 3.645 ;
        RECT 5.290 3.475 5.460 3.645 ;
        RECT 44.965 16.365 45.135 16.535 ;
        RECT 45.325 16.365 45.495 16.535 ;
        RECT 23.620 7.315 23.790 7.485 ;
        RECT 23.980 7.315 24.150 7.485 ;
        RECT 26.370 7.315 26.540 7.485 ;
        RECT 26.730 7.315 26.900 7.485 ;
        RECT 23.800 5.390 23.970 5.560 ;
        RECT 23.800 5.030 23.970 5.200 ;
        RECT 24.585 5.390 24.755 5.560 ;
        RECT 24.585 5.030 24.755 5.200 ;
        RECT 25.765 5.390 25.935 5.560 ;
        RECT 25.765 5.030 25.935 5.200 ;
        RECT 26.550 5.390 26.720 5.560 ;
        RECT 26.550 5.030 26.720 5.200 ;
        RECT 5.025 2.885 5.195 3.055 ;
        RECT 5.385 2.885 5.555 3.055 ;
        RECT 45.060 15.190 45.230 15.360 ;
        RECT 45.420 15.190 45.590 15.360 ;
        RECT 45.060 14.010 45.230 14.180 ;
        RECT 45.420 14.010 45.590 14.180 ;
        RECT 45.060 11.875 45.230 12.045 ;
        RECT 45.420 11.875 45.590 12.045 ;
        RECT 45.060 9.740 45.230 9.910 ;
        RECT 45.420 9.740 45.590 9.910 ;
        RECT 45.060 8.195 45.230 8.365 ;
        RECT 45.420 8.195 45.590 8.365 ;
        RECT 45.060 7.015 45.230 7.185 ;
        RECT 45.420 7.015 45.590 7.185 ;
        RECT 45.060 5.835 45.230 6.005 ;
        RECT 45.420 5.835 45.590 6.005 ;
        RECT 45.060 4.655 45.230 4.825 ;
        RECT 45.420 4.655 45.590 4.825 ;
        RECT 45.060 3.475 45.230 3.645 ;
        RECT 45.420 3.475 45.590 3.645 ;
        RECT 44.965 2.885 45.135 3.055 ;
        RECT 45.325 2.885 45.495 3.055 ;
      LAYER met1 ;
        RECT 4.940 16.300 5.640 16.600 ;
        RECT 44.880 16.300 45.580 16.600 ;
        RECT 6.045 15.390 6.745 15.425 ;
        RECT 4.695 15.160 6.745 15.390 ;
        RECT 6.045 15.125 6.745 15.160 ;
        RECT 43.775 15.390 44.475 15.425 ;
        RECT 43.775 15.160 45.825 15.390 ;
        RECT 43.775 15.125 44.475 15.160 ;
        RECT 6.045 14.210 6.745 14.245 ;
        RECT 4.695 13.980 6.745 14.210 ;
        RECT 6.045 13.945 6.745 13.980 ;
        RECT 43.775 14.210 44.475 14.245 ;
        RECT 43.775 13.980 45.825 14.210 ;
        RECT 43.775 13.945 44.475 13.980 ;
        RECT 6.045 12.075 6.745 12.110 ;
        RECT 4.695 11.845 6.745 12.075 ;
        RECT 6.045 11.810 6.745 11.845 ;
        RECT 43.775 12.075 44.475 12.110 ;
        RECT 43.775 11.845 45.825 12.075 ;
        RECT 43.775 11.810 44.475 11.845 ;
        RECT 6.045 9.940 6.745 9.975 ;
        RECT 4.695 9.710 6.745 9.940 ;
        RECT 6.045 9.675 6.745 9.710 ;
        RECT 43.775 9.940 44.475 9.975 ;
        RECT 43.775 9.710 45.825 9.940 ;
        RECT 43.775 9.675 44.475 9.710 ;
        RECT 6.045 8.395 6.745 8.430 ;
        RECT 4.695 8.165 6.745 8.395 ;
        RECT 6.045 8.130 6.745 8.165 ;
        RECT 43.775 8.395 44.475 8.430 ;
        RECT 43.775 8.165 45.825 8.395 ;
        RECT 43.775 8.130 44.475 8.165 ;
        RECT 23.535 7.250 24.235 7.550 ;
        RECT 26.285 7.250 26.985 7.550 ;
        RECT 6.045 7.215 6.745 7.250 ;
        RECT 4.695 6.985 6.745 7.215 ;
        RECT 6.045 6.950 6.745 6.985 ;
        RECT 43.775 7.215 44.475 7.250 ;
        RECT 43.775 6.985 45.825 7.215 ;
        RECT 43.775 6.950 44.475 6.985 ;
        RECT 6.045 6.035 6.745 6.070 ;
        RECT 4.695 5.805 6.745 6.035 ;
        RECT 6.045 5.770 6.745 5.805 ;
        RECT 43.775 6.035 44.475 6.070 ;
        RECT 43.775 5.805 45.825 6.035 ;
        RECT 24.555 5.645 24.785 5.795 ;
        RECT 23.735 4.945 24.785 5.645 ;
        RECT 6.045 4.855 6.745 4.890 ;
        RECT 4.695 4.625 6.745 4.855 ;
        RECT 24.555 4.795 24.785 4.945 ;
        RECT 25.735 5.645 25.965 5.795 ;
        RECT 43.775 5.770 44.475 5.805 ;
        RECT 25.735 4.945 26.785 5.645 ;
        RECT 25.735 4.795 25.965 4.945 ;
        RECT 43.775 4.855 44.475 4.890 ;
        RECT 6.045 4.590 6.745 4.625 ;
        RECT 43.775 4.625 45.825 4.855 ;
        RECT 43.775 4.590 44.475 4.625 ;
        RECT 6.045 3.675 6.745 3.710 ;
        RECT 4.695 3.445 6.745 3.675 ;
        RECT 6.045 3.410 6.745 3.445 ;
        RECT 43.775 3.675 44.475 3.710 ;
        RECT 43.775 3.445 45.825 3.675 ;
        RECT 43.775 3.410 44.475 3.445 ;
        RECT 4.940 2.820 5.640 3.120 ;
        RECT 44.880 2.820 45.580 3.120 ;
      LAYER via ;
        RECT 5.000 16.320 5.260 16.580 ;
        RECT 5.320 16.320 5.580 16.580 ;
        RECT 44.940 16.320 45.200 16.580 ;
        RECT 45.260 16.320 45.520 16.580 ;
        RECT 6.105 15.145 6.365 15.405 ;
        RECT 6.425 15.145 6.685 15.405 ;
        RECT 43.835 15.145 44.095 15.405 ;
        RECT 44.155 15.145 44.415 15.405 ;
        RECT 6.105 13.965 6.365 14.225 ;
        RECT 6.425 13.965 6.685 14.225 ;
        RECT 43.835 13.965 44.095 14.225 ;
        RECT 44.155 13.965 44.415 14.225 ;
        RECT 6.105 11.830 6.365 12.090 ;
        RECT 6.425 11.830 6.685 12.090 ;
        RECT 43.835 11.830 44.095 12.090 ;
        RECT 44.155 11.830 44.415 12.090 ;
        RECT 6.105 9.695 6.365 9.955 ;
        RECT 6.425 9.695 6.685 9.955 ;
        RECT 43.835 9.695 44.095 9.955 ;
        RECT 44.155 9.695 44.415 9.955 ;
        RECT 6.105 8.150 6.365 8.410 ;
        RECT 6.425 8.150 6.685 8.410 ;
        RECT 43.835 8.150 44.095 8.410 ;
        RECT 44.155 8.150 44.415 8.410 ;
        RECT 23.595 7.270 23.855 7.530 ;
        RECT 23.915 7.270 24.175 7.530 ;
        RECT 26.345 7.270 26.605 7.530 ;
        RECT 26.665 7.270 26.925 7.530 ;
        RECT 6.105 6.970 6.365 7.230 ;
        RECT 6.425 6.970 6.685 7.230 ;
        RECT 43.835 6.970 44.095 7.230 ;
        RECT 44.155 6.970 44.415 7.230 ;
        RECT 6.105 5.790 6.365 6.050 ;
        RECT 6.425 5.790 6.685 6.050 ;
        RECT 23.755 5.325 24.015 5.585 ;
        RECT 23.755 5.005 24.015 5.265 ;
        RECT 6.105 4.610 6.365 4.870 ;
        RECT 6.425 4.610 6.685 4.870 ;
        RECT 43.835 5.790 44.095 6.050 ;
        RECT 44.155 5.790 44.415 6.050 ;
        RECT 26.505 5.325 26.765 5.585 ;
        RECT 26.505 5.005 26.765 5.265 ;
        RECT 43.835 4.610 44.095 4.870 ;
        RECT 44.155 4.610 44.415 4.870 ;
        RECT 6.105 3.430 6.365 3.690 ;
        RECT 6.425 3.430 6.685 3.690 ;
        RECT 43.835 3.430 44.095 3.690 ;
        RECT 44.155 3.430 44.415 3.690 ;
        RECT 5.000 2.840 5.260 3.100 ;
        RECT 5.320 2.840 5.580 3.100 ;
        RECT 44.940 2.840 45.200 3.100 ;
        RECT 45.260 2.840 45.520 3.100 ;
      LAYER met2 ;
        RECT 4.990 16.600 5.590 16.650 ;
        RECT 44.930 16.600 45.530 16.650 ;
        RECT 4.990 16.565 6.545 16.600 ;
        RECT 43.975 16.565 45.530 16.600 ;
        RECT 4.990 16.335 12.275 16.565 ;
        RECT 4.990 16.300 6.545 16.335 ;
        RECT 4.990 16.250 5.590 16.300 ;
        RECT 6.245 15.475 6.545 16.300 ;
        RECT 6.095 15.075 6.695 15.475 ;
        RECT 6.245 14.295 6.545 15.075 ;
        RECT 12.045 14.700 12.275 16.335 ;
        RECT 38.245 16.335 45.530 16.565 ;
        RECT 38.245 14.700 38.475 16.335 ;
        RECT 43.975 16.300 45.530 16.335 ;
        RECT 43.975 15.475 44.275 16.300 ;
        RECT 44.930 16.250 45.530 16.300 ;
        RECT 43.825 15.075 44.425 15.475 ;
        RECT 12.045 14.655 12.480 14.700 ;
        RECT 38.040 14.655 38.475 14.700 ;
        RECT 12.045 14.515 16.290 14.655 ;
        RECT 34.230 14.515 38.475 14.655 ;
        RECT 12.045 14.470 12.480 14.515 ;
        RECT 38.040 14.470 38.475 14.515 ;
        RECT 43.975 14.295 44.275 15.075 ;
        RECT 6.095 13.895 6.695 14.295 ;
        RECT 43.825 13.895 44.425 14.295 ;
        RECT 6.245 12.160 6.545 13.895 ;
        RECT 43.975 12.160 44.275 13.895 ;
        RECT 6.095 11.760 6.695 12.160 ;
        RECT 43.825 11.760 44.425 12.160 ;
        RECT 6.245 10.025 6.545 11.760 ;
        RECT 43.975 10.025 44.275 11.760 ;
        RECT 6.095 9.625 6.695 10.025 ;
        RECT 43.825 9.625 44.425 10.025 ;
        RECT 6.245 8.480 6.545 9.625 ;
        RECT 43.975 8.480 44.275 9.625 ;
        RECT 6.095 8.080 6.695 8.480 ;
        RECT 43.825 8.080 44.425 8.480 ;
        RECT 6.245 7.300 6.545 8.080 ;
        RECT 6.095 6.900 6.695 7.300 ;
        RECT 23.585 7.200 24.185 7.600 ;
        RECT 26.335 7.200 26.935 7.600 ;
        RECT 43.975 7.300 44.275 8.080 ;
        RECT 6.245 6.120 6.545 6.900 ;
        RECT 6.095 5.720 6.695 6.120 ;
        RECT 6.245 4.940 6.545 5.720 ;
        RECT 12.045 5.135 12.480 5.180 ;
        RECT 12.045 4.995 16.290 5.135 ;
        RECT 12.045 4.950 12.480 4.995 ;
        RECT 6.095 4.540 6.695 4.940 ;
        RECT 6.245 3.760 6.545 4.540 ;
        RECT 6.095 3.360 6.695 3.760 ;
        RECT 4.990 3.120 5.590 3.170 ;
        RECT 6.245 3.120 6.545 3.360 ;
        RECT 4.990 3.085 6.545 3.120 ;
        RECT 12.045 3.085 12.275 4.950 ;
        RECT 23.685 4.235 24.085 7.200 ;
        RECT 26.435 4.235 26.835 7.200 ;
        RECT 43.825 6.900 44.425 7.300 ;
        RECT 43.975 6.120 44.275 6.900 ;
        RECT 43.825 5.720 44.425 6.120 ;
        RECT 38.040 5.135 38.475 5.180 ;
        RECT 34.230 4.995 38.475 5.135 ;
        RECT 38.040 4.950 38.475 4.995 ;
        RECT 23.685 3.835 26.835 4.235 ;
        RECT 4.990 2.855 12.275 3.085 ;
        RECT 4.990 2.820 6.545 2.855 ;
        RECT 4.990 2.770 5.590 2.820 ;
        RECT 6.245 0.570 6.545 2.820 ;
        RECT 25.060 0.570 25.460 3.835 ;
        RECT 38.245 3.085 38.475 4.950 ;
        RECT 43.975 4.940 44.275 5.720 ;
        RECT 43.825 4.540 44.425 4.940 ;
        RECT 43.975 3.760 44.275 4.540 ;
        RECT 43.825 3.360 44.425 3.760 ;
        RECT 43.975 3.120 44.275 3.360 ;
        RECT 44.930 3.120 45.530 3.170 ;
        RECT 43.975 3.085 45.530 3.120 ;
        RECT 38.245 2.855 45.530 3.085 ;
        RECT 43.975 2.820 45.530 2.855 ;
        RECT 43.975 0.570 44.275 2.820 ;
        RECT 44.930 2.770 45.530 2.820 ;
        RECT 5.995 0.170 6.795 0.570 ;
        RECT 24.860 0.170 25.660 0.570 ;
        RECT 43.725 0.170 44.525 0.570 ;
      LAYER via2 ;
        RECT 6.055 0.230 6.335 0.510 ;
        RECT 6.455 0.230 6.735 0.510 ;
        RECT 24.920 0.230 25.200 0.510 ;
        RECT 25.320 0.230 25.600 0.510 ;
        RECT 43.785 0.230 44.065 0.510 ;
        RECT 44.185 0.230 44.465 0.510 ;
      LAYER met3 ;
        RECT 0.000 0.170 50.520 0.570 ;
    END
  END vss
  PIN vn
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 24.800 9.135 25.130 9.305 ;
      LAYER mcon ;
        RECT 24.880 9.135 25.050 9.305 ;
      LAYER met1 ;
        RECT 21.125 10.555 21.825 10.590 ;
        RECT 21.125 10.325 25.080 10.555 ;
        RECT 21.125 10.290 21.825 10.325 ;
        RECT 24.850 9.335 25.080 10.325 ;
        RECT 24.820 9.105 25.110 9.335 ;
      LAYER via ;
        RECT 21.185 10.310 21.445 10.570 ;
        RECT 21.505 10.310 21.765 10.570 ;
      LAYER met2 ;
        RECT 21.075 10.240 21.875 10.640 ;
      LAYER via2 ;
        RECT 21.135 10.300 21.415 10.580 ;
        RECT 21.535 10.300 21.815 10.580 ;
      LAYER met3 ;
        RECT 20.970 10.240 21.980 10.640 ;
      LAYER via3 ;
        RECT 21.115 10.280 21.435 10.600 ;
        RECT 21.515 10.280 21.835 10.600 ;
      LAYER met4 ;
        RECT 24.010 19.850 24.510 20.100 ;
        RECT 18.250 19.350 24.510 19.850 ;
        RECT 18.250 10.690 18.750 19.350 ;
        RECT 18.250 10.190 21.990 10.690 ;
    END
  END vn
  PIN vp
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 25.390 9.135 25.720 9.305 ;
      LAYER mcon ;
        RECT 25.470 9.135 25.640 9.305 ;
      LAYER met1 ;
        RECT 28.695 10.555 29.395 10.590 ;
        RECT 25.440 10.325 29.395 10.555 ;
        RECT 25.440 9.335 25.670 10.325 ;
        RECT 28.695 10.290 29.395 10.325 ;
        RECT 25.410 9.105 25.700 9.335 ;
      LAYER via ;
        RECT 28.755 10.310 29.015 10.570 ;
        RECT 29.075 10.310 29.335 10.570 ;
      LAYER met2 ;
        RECT 28.645 10.240 29.445 10.640 ;
      LAYER via2 ;
        RECT 28.705 10.300 28.985 10.580 ;
        RECT 29.105 10.300 29.385 10.580 ;
      LAYER met3 ;
        RECT 28.540 10.240 29.550 10.640 ;
      LAYER via3 ;
        RECT 28.685 10.280 29.005 10.600 ;
        RECT 29.085 10.280 29.405 10.600 ;
      LAYER met4 ;
        RECT 26.010 19.850 26.510 20.100 ;
        RECT 26.010 19.350 32.270 19.850 ;
        RECT 31.770 10.690 32.270 19.350 ;
        RECT 28.530 10.190 32.270 10.690 ;
    END
  END vp
  OBS
      LAYER nwell ;
        RECT 19.760 17.810 30.720 17.860 ;
      LAYER pwell ;
        RECT 4.565 13.230 5.825 16.140 ;
      LAYER nwell ;
        RECT 19.760 14.430 19.810 17.810 ;
      LAYER pwell ;
        RECT 19.810 17.380 30.670 17.810 ;
        RECT 19.810 14.860 20.240 17.380 ;
      LAYER nwell ;
        RECT 20.240 14.860 30.240 17.380 ;
      LAYER pwell ;
        RECT 30.240 14.860 30.670 17.380 ;
        RECT 19.810 14.430 30.670 14.860 ;
      LAYER nwell ;
        RECT 30.670 14.430 30.720 17.810 ;
        RECT 19.760 14.380 30.720 14.430 ;
      LAYER pwell ;
        RECT 44.695 13.230 45.955 16.140 ;
        RECT 4.565 11.095 5.825 12.825 ;
        RECT 44.695 11.095 45.955 12.825 ;
        RECT 4.565 8.960 5.825 10.690 ;
        RECT 4.565 3.285 5.825 8.555 ;
        RECT 23.805 7.815 26.715 9.075 ;
        RECT 44.695 8.960 45.955 10.690 ;
        RECT 24.395 4.665 26.125 5.925 ;
        RECT 44.695 3.285 45.955 8.555 ;
      LAYER li1 ;
        RECT 4.675 15.780 5.715 15.950 ;
        RECT 20.645 15.685 20.815 16.725 ;
        RECT 29.665 15.685 29.835 16.725 ;
        RECT 44.805 15.780 45.845 15.950 ;
        RECT 4.675 14.600 5.715 14.770 ;
        RECT 44.805 14.600 45.845 14.770 ;
        RECT 4.675 13.420 5.715 13.590 ;
        RECT 44.805 13.420 45.845 13.590 ;
        RECT 4.675 12.465 5.715 12.635 ;
        RECT 44.805 12.465 45.845 12.635 ;
        RECT 4.675 11.285 5.715 11.455 ;
        RECT 44.805 11.285 45.845 11.455 ;
        RECT 4.675 10.330 5.715 10.500 ;
        RECT 44.805 10.330 45.845 10.500 ;
        RECT 4.675 9.150 5.715 9.320 ;
        RECT 44.805 9.150 45.845 9.320 ;
        RECT 24.585 7.925 24.755 8.965 ;
        RECT 25.175 7.925 25.345 8.965 ;
        RECT 25.765 7.925 25.935 8.965 ;
        RECT 4.675 7.605 5.715 7.775 ;
        RECT 44.805 7.605 45.845 7.775 ;
        RECT 4.675 6.425 5.715 6.595 ;
        RECT 44.805 6.425 45.845 6.595 ;
        RECT 4.675 5.245 5.715 5.415 ;
        RECT 25.175 4.775 25.345 5.815 ;
        RECT 44.805 5.245 45.845 5.415 ;
        RECT 4.675 4.065 5.715 4.235 ;
        RECT 44.805 4.065 45.845 4.235 ;
      LAYER mcon ;
        RECT 20.645 16.300 20.815 16.470 ;
        RECT 4.930 15.780 5.100 15.950 ;
        RECT 5.290 15.780 5.460 15.950 ;
        RECT 20.645 15.940 20.815 16.110 ;
        RECT 29.665 16.300 29.835 16.470 ;
        RECT 29.665 15.940 29.835 16.110 ;
        RECT 45.060 15.780 45.230 15.950 ;
        RECT 45.420 15.780 45.590 15.950 ;
        RECT 4.930 14.600 5.100 14.770 ;
        RECT 5.290 14.600 5.460 14.770 ;
        RECT 45.060 14.600 45.230 14.770 ;
        RECT 45.420 14.600 45.590 14.770 ;
        RECT 4.930 13.420 5.100 13.590 ;
        RECT 5.290 13.420 5.460 13.590 ;
        RECT 45.060 13.420 45.230 13.590 ;
        RECT 45.420 13.420 45.590 13.590 ;
        RECT 4.930 12.465 5.100 12.635 ;
        RECT 5.290 12.465 5.460 12.635 ;
        RECT 45.060 12.465 45.230 12.635 ;
        RECT 45.420 12.465 45.590 12.635 ;
        RECT 4.930 11.285 5.100 11.455 ;
        RECT 5.290 11.285 5.460 11.455 ;
        RECT 45.060 11.285 45.230 11.455 ;
        RECT 45.420 11.285 45.590 11.455 ;
        RECT 4.930 10.330 5.100 10.500 ;
        RECT 5.290 10.330 5.460 10.500 ;
        RECT 45.060 10.330 45.230 10.500 ;
        RECT 45.420 10.330 45.590 10.500 ;
        RECT 4.930 9.150 5.100 9.320 ;
        RECT 5.290 9.150 5.460 9.320 ;
        RECT 45.060 9.150 45.230 9.320 ;
        RECT 45.420 9.150 45.590 9.320 ;
        RECT 24.585 8.540 24.755 8.710 ;
        RECT 24.585 8.180 24.755 8.350 ;
        RECT 25.175 8.540 25.345 8.710 ;
        RECT 25.175 8.180 25.345 8.350 ;
        RECT 25.765 8.540 25.935 8.710 ;
        RECT 25.765 8.180 25.935 8.350 ;
        RECT 4.930 7.605 5.100 7.775 ;
        RECT 5.290 7.605 5.460 7.775 ;
        RECT 45.060 7.605 45.230 7.775 ;
        RECT 45.420 7.605 45.590 7.775 ;
        RECT 4.930 6.425 5.100 6.595 ;
        RECT 5.290 6.425 5.460 6.595 ;
        RECT 45.060 6.425 45.230 6.595 ;
        RECT 45.420 6.425 45.590 6.595 ;
        RECT 4.930 5.245 5.100 5.415 ;
        RECT 5.290 5.245 5.460 5.415 ;
        RECT 25.175 5.390 25.345 5.560 ;
        RECT 45.060 5.245 45.230 5.415 ;
        RECT 45.420 5.245 45.590 5.415 ;
        RECT 25.175 5.030 25.345 5.200 ;
        RECT 4.930 4.065 5.100 4.235 ;
        RECT 5.290 4.065 5.460 4.235 ;
        RECT 45.060 4.065 45.230 4.235 ;
        RECT 45.420 4.065 45.590 4.235 ;
      LAYER met1 ;
        RECT 20.615 16.320 20.845 16.705 ;
        RECT 19.315 16.090 20.845 16.320 ;
        RECT 4.695 15.750 9.985 15.980 ;
        RECT 7.195 14.800 7.425 15.750 ;
        RECT 4.695 14.570 7.425 14.800 ;
        RECT 7.195 13.620 7.425 14.570 ;
        RECT 4.695 13.390 7.425 13.620 ;
        RECT 9.755 13.615 9.985 15.750 ;
        RECT 11.130 13.875 11.830 14.175 ;
        RECT 9.755 13.315 10.455 13.615 ;
        RECT 4.695 12.495 8.790 12.665 ;
        RECT 4.695 12.435 9.260 12.495 ;
        RECT 7.195 11.485 7.425 12.435 ;
        RECT 4.695 11.255 7.425 11.485 ;
        RECT 8.560 12.195 9.260 12.435 ;
        RECT 4.695 10.300 7.755 10.530 ;
        RECT 7.525 10.255 7.755 10.300 ;
        RECT 7.525 9.955 8.225 10.255 ;
        RECT 7.525 9.395 8.225 9.695 ;
        RECT 7.525 9.350 7.755 9.395 ;
        RECT 4.695 9.120 7.755 9.350 ;
        RECT 4.695 7.575 7.425 7.805 ;
        RECT 7.195 6.625 7.425 7.575 ;
        RECT 8.560 7.455 8.790 12.195 ;
        RECT 9.755 11.375 9.985 13.315 ;
        RECT 11.130 13.055 11.360 13.875 ;
        RECT 11.130 12.755 11.830 13.055 ;
        RECT 11.130 11.935 11.360 12.755 ;
        RECT 11.130 11.635 11.830 11.935 ;
        RECT 9.755 11.075 10.455 11.375 ;
        RECT 9.755 8.575 9.985 11.075 ;
        RECT 11.130 10.815 11.360 11.635 ;
        RECT 11.130 10.515 11.830 10.815 ;
        RECT 11.130 9.135 11.360 10.515 ;
        RECT 11.130 8.835 11.830 9.135 ;
        RECT 9.755 8.275 10.455 8.575 ;
        RECT 8.560 7.155 9.260 7.455 ;
        RECT 4.695 6.395 7.425 6.625 ;
        RECT 7.195 5.445 7.425 6.395 ;
        RECT 9.755 6.335 9.985 8.275 ;
        RECT 11.130 8.015 11.360 8.835 ;
        RECT 11.130 7.715 11.830 8.015 ;
        RECT 11.130 6.895 11.360 7.715 ;
        RECT 16.750 7.055 17.050 7.290 ;
        RECT 19.315 7.055 19.545 16.090 ;
        RECT 20.615 15.705 20.845 16.090 ;
        RECT 29.635 16.320 29.865 16.705 ;
        RECT 29.635 16.090 31.205 16.320 ;
        RECT 29.635 15.705 29.865 16.090 ;
        RECT 24.555 7.055 24.785 8.945 ;
        RECT 11.130 6.595 11.830 6.895 ;
        RECT 16.750 6.825 24.785 7.055 ;
        RECT 9.755 6.035 10.455 6.335 ;
        RECT 4.695 5.215 7.425 5.445 ;
        RECT 7.195 4.265 7.425 5.215 ;
        RECT 11.130 5.775 11.360 6.595 ;
        RECT 16.750 6.590 17.050 6.825 ;
        RECT 11.130 5.475 11.830 5.775 ;
        RECT 11.130 4.265 11.360 5.475 ;
        RECT 25.145 4.795 25.375 8.945 ;
        RECT 25.735 7.055 25.965 8.945 ;
        RECT 30.975 7.055 31.205 16.090 ;
        RECT 40.535 15.750 45.825 15.980 ;
        RECT 38.690 13.875 39.390 14.175 ;
        RECT 39.160 13.055 39.390 13.875 ;
        RECT 40.535 13.615 40.765 15.750 ;
        RECT 40.065 13.315 40.765 13.615 ;
        RECT 43.095 14.800 43.325 15.750 ;
        RECT 43.095 14.570 45.825 14.800 ;
        RECT 43.095 13.620 43.325 14.570 ;
        RECT 43.095 13.390 45.825 13.620 ;
        RECT 38.690 12.755 39.390 13.055 ;
        RECT 39.160 11.935 39.390 12.755 ;
        RECT 38.690 11.635 39.390 11.935 ;
        RECT 39.160 10.815 39.390 11.635 ;
        RECT 40.535 11.375 40.765 13.315 ;
        RECT 41.730 12.495 45.825 12.665 ;
        RECT 41.260 12.435 45.825 12.495 ;
        RECT 41.260 12.195 41.960 12.435 ;
        RECT 40.065 11.075 40.765 11.375 ;
        RECT 38.690 10.515 39.390 10.815 ;
        RECT 39.160 9.135 39.390 10.515 ;
        RECT 38.690 8.835 39.390 9.135 ;
        RECT 39.160 8.015 39.390 8.835 ;
        RECT 40.535 8.575 40.765 11.075 ;
        RECT 40.065 8.275 40.765 8.575 ;
        RECT 38.690 7.715 39.390 8.015 ;
        RECT 33.470 7.055 33.770 7.290 ;
        RECT 25.735 6.825 33.770 7.055 ;
        RECT 39.160 6.895 39.390 7.715 ;
        RECT 33.470 6.590 33.770 6.825 ;
        RECT 38.690 6.595 39.390 6.895 ;
        RECT 39.160 5.775 39.390 6.595 ;
        RECT 40.535 6.335 40.765 8.275 ;
        RECT 41.730 7.455 41.960 12.195 ;
        RECT 43.095 11.485 43.325 12.435 ;
        RECT 43.095 11.255 45.825 11.485 ;
        RECT 42.765 10.300 45.825 10.530 ;
        RECT 42.765 10.255 42.995 10.300 ;
        RECT 42.295 9.955 42.995 10.255 ;
        RECT 42.295 9.395 42.995 9.695 ;
        RECT 42.765 9.350 42.995 9.395 ;
        RECT 42.765 9.120 45.825 9.350 ;
        RECT 41.260 7.155 41.960 7.455 ;
        RECT 43.095 7.575 45.825 7.805 ;
        RECT 40.065 6.035 40.765 6.335 ;
        RECT 43.095 6.625 43.325 7.575 ;
        RECT 43.095 6.395 45.825 6.625 ;
        RECT 38.690 5.475 39.390 5.775 ;
        RECT 4.695 4.035 11.360 4.265 ;
        RECT 39.160 4.265 39.390 5.475 ;
        RECT 43.095 5.445 43.325 6.395 ;
        RECT 43.095 5.215 45.825 5.445 ;
        RECT 43.095 4.265 43.325 5.215 ;
        RECT 39.160 4.035 45.825 4.265 ;
      LAYER via ;
        RECT 11.190 13.895 11.450 14.155 ;
        RECT 11.510 13.895 11.770 14.155 ;
        RECT 9.815 13.335 10.075 13.595 ;
        RECT 10.135 13.335 10.395 13.595 ;
        RECT 8.620 12.215 8.880 12.475 ;
        RECT 8.940 12.215 9.200 12.475 ;
        RECT 7.585 9.975 7.845 10.235 ;
        RECT 7.905 9.975 8.165 10.235 ;
        RECT 7.585 9.415 7.845 9.675 ;
        RECT 7.905 9.415 8.165 9.675 ;
        RECT 11.190 12.775 11.450 13.035 ;
        RECT 11.510 12.775 11.770 13.035 ;
        RECT 11.190 11.655 11.450 11.915 ;
        RECT 11.510 11.655 11.770 11.915 ;
        RECT 9.815 11.095 10.075 11.355 ;
        RECT 10.135 11.095 10.395 11.355 ;
        RECT 11.190 10.535 11.450 10.795 ;
        RECT 11.510 10.535 11.770 10.795 ;
        RECT 11.190 8.855 11.450 9.115 ;
        RECT 11.510 8.855 11.770 9.115 ;
        RECT 9.815 8.295 10.075 8.555 ;
        RECT 10.135 8.295 10.395 8.555 ;
        RECT 8.620 7.175 8.880 7.435 ;
        RECT 8.940 7.175 9.200 7.435 ;
        RECT 11.190 7.735 11.450 7.995 ;
        RECT 11.510 7.735 11.770 7.995 ;
        RECT 16.770 6.970 17.030 7.230 ;
        RECT 11.190 6.615 11.450 6.875 ;
        RECT 11.510 6.615 11.770 6.875 ;
        RECT 16.770 6.650 17.030 6.910 ;
        RECT 9.815 6.055 10.075 6.315 ;
        RECT 10.135 6.055 10.395 6.315 ;
        RECT 11.190 5.495 11.450 5.755 ;
        RECT 11.510 5.495 11.770 5.755 ;
        RECT 38.750 13.895 39.010 14.155 ;
        RECT 39.070 13.895 39.330 14.155 ;
        RECT 40.125 13.335 40.385 13.595 ;
        RECT 40.445 13.335 40.705 13.595 ;
        RECT 38.750 12.775 39.010 13.035 ;
        RECT 39.070 12.775 39.330 13.035 ;
        RECT 38.750 11.655 39.010 11.915 ;
        RECT 39.070 11.655 39.330 11.915 ;
        RECT 41.320 12.215 41.580 12.475 ;
        RECT 41.640 12.215 41.900 12.475 ;
        RECT 40.125 11.095 40.385 11.355 ;
        RECT 40.445 11.095 40.705 11.355 ;
        RECT 38.750 10.535 39.010 10.795 ;
        RECT 39.070 10.535 39.330 10.795 ;
        RECT 38.750 8.855 39.010 9.115 ;
        RECT 39.070 8.855 39.330 9.115 ;
        RECT 40.125 8.295 40.385 8.555 ;
        RECT 40.445 8.295 40.705 8.555 ;
        RECT 38.750 7.735 39.010 7.995 ;
        RECT 39.070 7.735 39.330 7.995 ;
        RECT 33.490 6.970 33.750 7.230 ;
        RECT 33.490 6.650 33.750 6.910 ;
        RECT 38.750 6.615 39.010 6.875 ;
        RECT 39.070 6.615 39.330 6.875 ;
        RECT 42.355 9.975 42.615 10.235 ;
        RECT 42.675 9.975 42.935 10.235 ;
        RECT 42.355 9.415 42.615 9.675 ;
        RECT 42.675 9.415 42.935 9.675 ;
        RECT 41.320 7.175 41.580 7.435 ;
        RECT 41.640 7.175 41.900 7.435 ;
        RECT 40.125 6.055 40.385 6.315 ;
        RECT 40.445 6.055 40.705 6.315 ;
        RECT 38.750 5.495 39.010 5.755 ;
        RECT 39.070 5.495 39.330 5.755 ;
      LAYER met2 ;
        RECT 16.430 14.935 16.750 15.375 ;
        RECT 12.620 14.795 16.750 14.935 ;
        RECT 16.430 14.375 16.750 14.795 ;
        RECT 12.620 14.235 16.750 14.375 ;
        RECT 11.180 14.140 11.780 14.225 ;
        RECT 11.180 14.095 12.480 14.140 ;
        RECT 11.180 13.955 16.290 14.095 ;
        RECT 11.180 13.910 12.480 13.955 ;
        RECT 11.180 13.825 11.780 13.910 ;
        RECT 16.430 13.815 16.750 14.235 ;
        RECT 12.620 13.675 16.750 13.815 ;
        RECT 9.805 13.580 10.405 13.665 ;
        RECT 9.805 13.535 12.480 13.580 ;
        RECT 9.805 13.395 16.290 13.535 ;
        RECT 9.805 13.350 12.480 13.395 ;
        RECT 9.805 13.265 10.405 13.350 ;
        RECT 16.430 13.255 16.750 13.675 ;
        RECT 12.620 13.115 16.750 13.255 ;
        RECT 11.180 13.020 11.780 13.105 ;
        RECT 11.180 12.975 12.480 13.020 ;
        RECT 11.180 12.835 16.290 12.975 ;
        RECT 11.180 12.790 12.480 12.835 ;
        RECT 11.180 12.705 11.780 12.790 ;
        RECT 16.430 12.695 16.750 13.115 ;
        RECT 12.620 12.555 16.750 12.695 ;
        RECT 8.610 12.460 9.210 12.545 ;
        RECT 8.610 12.415 12.480 12.460 ;
        RECT 8.610 12.275 16.290 12.415 ;
        RECT 8.610 12.230 12.480 12.275 ;
        RECT 8.610 12.145 9.210 12.230 ;
        RECT 16.430 12.135 16.750 12.555 ;
        RECT 12.620 11.995 16.750 12.135 ;
        RECT 11.180 11.900 11.780 11.985 ;
        RECT 11.180 11.855 12.480 11.900 ;
        RECT 11.180 11.715 16.290 11.855 ;
        RECT 11.180 11.670 12.480 11.715 ;
        RECT 11.180 11.585 11.780 11.670 ;
        RECT 16.430 11.575 16.750 11.995 ;
        RECT 12.620 11.435 16.750 11.575 ;
        RECT 9.805 11.340 10.405 11.425 ;
        RECT 9.805 11.295 12.480 11.340 ;
        RECT 9.805 11.155 16.290 11.295 ;
        RECT 9.805 11.110 12.480 11.155 ;
        RECT 9.805 11.025 10.405 11.110 ;
        RECT 16.430 11.015 16.750 11.435 ;
        RECT 12.620 10.875 16.750 11.015 ;
        RECT 11.180 10.780 11.780 10.865 ;
        RECT 11.180 10.735 12.480 10.780 ;
        RECT 11.180 10.595 16.290 10.735 ;
        RECT 11.180 10.550 12.480 10.595 ;
        RECT 11.180 10.465 11.780 10.550 ;
        RECT 16.430 10.455 16.750 10.875 ;
        RECT 12.620 10.315 16.750 10.455 ;
        RECT 7.575 10.220 8.175 10.305 ;
        RECT 7.575 10.175 12.480 10.220 ;
        RECT 7.575 10.035 16.290 10.175 ;
        RECT 7.575 9.990 12.480 10.035 ;
        RECT 7.575 9.905 8.175 9.990 ;
        RECT 16.430 9.895 16.750 10.315 ;
        RECT 12.620 9.755 16.750 9.895 ;
        RECT 7.575 9.660 8.175 9.745 ;
        RECT 7.575 9.615 12.480 9.660 ;
        RECT 7.575 9.475 16.290 9.615 ;
        RECT 7.575 9.430 12.480 9.475 ;
        RECT 7.575 9.345 8.175 9.430 ;
        RECT 16.430 9.335 16.750 9.755 ;
        RECT 12.620 9.195 16.750 9.335 ;
        RECT 11.180 9.100 11.780 9.185 ;
        RECT 11.180 9.055 12.480 9.100 ;
        RECT 11.180 8.915 16.290 9.055 ;
        RECT 11.180 8.870 12.480 8.915 ;
        RECT 11.180 8.785 11.780 8.870 ;
        RECT 16.430 8.775 16.750 9.195 ;
        RECT 12.620 8.635 16.750 8.775 ;
        RECT 9.805 8.540 10.405 8.625 ;
        RECT 9.805 8.495 12.480 8.540 ;
        RECT 9.805 8.355 16.290 8.495 ;
        RECT 9.805 8.310 12.480 8.355 ;
        RECT 9.805 8.225 10.405 8.310 ;
        RECT 16.430 8.215 16.750 8.635 ;
        RECT 12.620 8.075 16.750 8.215 ;
        RECT 11.180 7.980 11.780 8.065 ;
        RECT 11.180 7.935 12.480 7.980 ;
        RECT 11.180 7.795 16.290 7.935 ;
        RECT 11.180 7.750 12.480 7.795 ;
        RECT 11.180 7.665 11.780 7.750 ;
        RECT 16.430 7.655 16.750 8.075 ;
        RECT 12.620 7.515 16.750 7.655 ;
        RECT 8.610 7.420 9.210 7.505 ;
        RECT 8.610 7.375 12.480 7.420 ;
        RECT 8.610 7.235 16.290 7.375 ;
        RECT 16.430 7.240 16.750 7.515 ;
        RECT 33.770 14.935 34.090 15.375 ;
        RECT 33.770 14.795 37.900 14.935 ;
        RECT 33.770 14.375 34.090 14.795 ;
        RECT 33.770 14.235 37.900 14.375 ;
        RECT 33.770 13.815 34.090 14.235 ;
        RECT 38.740 14.140 39.340 14.225 ;
        RECT 38.040 14.095 39.340 14.140 ;
        RECT 34.230 13.955 39.340 14.095 ;
        RECT 38.040 13.910 39.340 13.955 ;
        RECT 38.740 13.825 39.340 13.910 ;
        RECT 33.770 13.675 37.900 13.815 ;
        RECT 33.770 13.255 34.090 13.675 ;
        RECT 40.115 13.580 40.715 13.665 ;
        RECT 38.040 13.535 40.715 13.580 ;
        RECT 34.230 13.395 40.715 13.535 ;
        RECT 38.040 13.350 40.715 13.395 ;
        RECT 40.115 13.265 40.715 13.350 ;
        RECT 33.770 13.115 37.900 13.255 ;
        RECT 33.770 12.695 34.090 13.115 ;
        RECT 38.740 13.020 39.340 13.105 ;
        RECT 38.040 12.975 39.340 13.020 ;
        RECT 34.230 12.835 39.340 12.975 ;
        RECT 38.040 12.790 39.340 12.835 ;
        RECT 38.740 12.705 39.340 12.790 ;
        RECT 33.770 12.555 37.900 12.695 ;
        RECT 33.770 12.135 34.090 12.555 ;
        RECT 41.310 12.460 41.910 12.545 ;
        RECT 38.040 12.415 41.910 12.460 ;
        RECT 34.230 12.275 41.910 12.415 ;
        RECT 38.040 12.230 41.910 12.275 ;
        RECT 41.310 12.145 41.910 12.230 ;
        RECT 33.770 11.995 37.900 12.135 ;
        RECT 33.770 11.575 34.090 11.995 ;
        RECT 38.740 11.900 39.340 11.985 ;
        RECT 38.040 11.855 39.340 11.900 ;
        RECT 34.230 11.715 39.340 11.855 ;
        RECT 38.040 11.670 39.340 11.715 ;
        RECT 38.740 11.585 39.340 11.670 ;
        RECT 33.770 11.435 37.900 11.575 ;
        RECT 33.770 11.015 34.090 11.435 ;
        RECT 40.115 11.340 40.715 11.425 ;
        RECT 38.040 11.295 40.715 11.340 ;
        RECT 34.230 11.155 40.715 11.295 ;
        RECT 38.040 11.110 40.715 11.155 ;
        RECT 40.115 11.025 40.715 11.110 ;
        RECT 33.770 10.875 37.900 11.015 ;
        RECT 33.770 10.455 34.090 10.875 ;
        RECT 38.740 10.780 39.340 10.865 ;
        RECT 38.040 10.735 39.340 10.780 ;
        RECT 34.230 10.595 39.340 10.735 ;
        RECT 38.040 10.550 39.340 10.595 ;
        RECT 38.740 10.465 39.340 10.550 ;
        RECT 33.770 10.315 37.900 10.455 ;
        RECT 33.770 9.895 34.090 10.315 ;
        RECT 42.345 10.220 42.945 10.305 ;
        RECT 38.040 10.175 42.945 10.220 ;
        RECT 34.230 10.035 42.945 10.175 ;
        RECT 38.040 9.990 42.945 10.035 ;
        RECT 42.345 9.905 42.945 9.990 ;
        RECT 33.770 9.755 37.900 9.895 ;
        RECT 33.770 9.335 34.090 9.755 ;
        RECT 42.345 9.660 42.945 9.745 ;
        RECT 38.040 9.615 42.945 9.660 ;
        RECT 34.230 9.475 42.945 9.615 ;
        RECT 38.040 9.430 42.945 9.475 ;
        RECT 42.345 9.345 42.945 9.430 ;
        RECT 33.770 9.195 37.900 9.335 ;
        RECT 33.770 8.775 34.090 9.195 ;
        RECT 38.740 9.100 39.340 9.185 ;
        RECT 38.040 9.055 39.340 9.100 ;
        RECT 34.230 8.915 39.340 9.055 ;
        RECT 38.040 8.870 39.340 8.915 ;
        RECT 38.740 8.785 39.340 8.870 ;
        RECT 33.770 8.635 37.900 8.775 ;
        RECT 33.770 8.215 34.090 8.635 ;
        RECT 40.115 8.540 40.715 8.625 ;
        RECT 38.040 8.495 40.715 8.540 ;
        RECT 34.230 8.355 40.715 8.495 ;
        RECT 38.040 8.310 40.715 8.355 ;
        RECT 40.115 8.225 40.715 8.310 ;
        RECT 33.770 8.075 37.900 8.215 ;
        RECT 33.770 7.655 34.090 8.075 ;
        RECT 38.740 7.980 39.340 8.065 ;
        RECT 38.040 7.935 39.340 7.980 ;
        RECT 34.230 7.795 39.340 7.935 ;
        RECT 38.040 7.750 39.340 7.795 ;
        RECT 38.740 7.665 39.340 7.750 ;
        RECT 33.770 7.515 37.900 7.655 ;
        RECT 33.770 7.240 34.090 7.515 ;
        RECT 41.310 7.420 41.910 7.505 ;
        RECT 38.040 7.375 41.910 7.420 ;
        RECT 8.610 7.190 12.480 7.235 ;
        RECT 8.610 7.105 9.210 7.190 ;
        RECT 16.430 7.095 17.100 7.240 ;
        RECT 12.620 6.955 17.100 7.095 ;
        RECT 11.180 6.860 11.780 6.945 ;
        RECT 11.180 6.815 12.480 6.860 ;
        RECT 11.180 6.675 16.290 6.815 ;
        RECT 11.180 6.630 12.480 6.675 ;
        RECT 16.430 6.640 17.100 6.955 ;
        RECT 33.420 7.095 34.090 7.240 ;
        RECT 34.230 7.235 41.910 7.375 ;
        RECT 38.040 7.190 41.910 7.235 ;
        RECT 41.310 7.105 41.910 7.190 ;
        RECT 33.420 6.955 37.900 7.095 ;
        RECT 33.420 6.640 34.090 6.955 ;
        RECT 38.740 6.860 39.340 6.945 ;
        RECT 38.040 6.815 39.340 6.860 ;
        RECT 34.230 6.675 39.340 6.815 ;
        RECT 11.180 6.545 11.780 6.630 ;
        RECT 16.430 6.535 16.750 6.640 ;
        RECT 12.620 6.395 16.750 6.535 ;
        RECT 9.805 6.300 10.405 6.385 ;
        RECT 9.805 6.255 12.480 6.300 ;
        RECT 9.805 6.115 16.290 6.255 ;
        RECT 9.805 6.070 12.480 6.115 ;
        RECT 9.805 5.985 10.405 6.070 ;
        RECT 16.430 5.975 16.750 6.395 ;
        RECT 12.620 5.835 16.750 5.975 ;
        RECT 11.180 5.740 11.780 5.825 ;
        RECT 11.180 5.695 12.480 5.740 ;
        RECT 11.180 5.555 16.290 5.695 ;
        RECT 11.180 5.510 12.480 5.555 ;
        RECT 11.180 5.425 11.780 5.510 ;
        RECT 16.430 5.415 16.750 5.835 ;
        RECT 12.620 5.275 16.750 5.415 ;
        RECT 16.430 4.855 16.750 5.275 ;
        RECT 12.620 4.715 16.750 4.855 ;
        RECT 16.430 4.275 16.750 4.715 ;
        RECT 33.770 6.535 34.090 6.640 ;
        RECT 38.040 6.630 39.340 6.675 ;
        RECT 38.740 6.545 39.340 6.630 ;
        RECT 33.770 6.395 37.900 6.535 ;
        RECT 33.770 5.975 34.090 6.395 ;
        RECT 40.115 6.300 40.715 6.385 ;
        RECT 38.040 6.255 40.715 6.300 ;
        RECT 34.230 6.115 40.715 6.255 ;
        RECT 38.040 6.070 40.715 6.115 ;
        RECT 40.115 5.985 40.715 6.070 ;
        RECT 33.770 5.835 37.900 5.975 ;
        RECT 33.770 5.415 34.090 5.835 ;
        RECT 38.740 5.740 39.340 5.825 ;
        RECT 38.040 5.695 39.340 5.740 ;
        RECT 34.230 5.555 39.340 5.695 ;
        RECT 38.040 5.510 39.340 5.555 ;
        RECT 38.740 5.425 39.340 5.510 ;
        RECT 33.770 5.275 37.900 5.415 ;
        RECT 33.770 4.855 34.090 5.275 ;
        RECT 33.770 4.715 37.900 4.855 ;
        RECT 33.770 4.275 34.090 4.715 ;
  END
END comparator
END LIBRARY

