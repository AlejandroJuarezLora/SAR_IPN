magic
tech sky130B
magscale 1 2
timestamp 1696285618
<< nwell >>
rect -226 -284 226 284
<< pmos >>
rect -30 -136 30 64
<< pdiff >>
rect -88 34 -30 64
rect -88 -106 -76 34
rect -42 -106 -30 34
rect -88 -136 -30 -106
rect 30 34 88 64
rect 30 -106 42 34
rect 76 -106 88 34
rect 30 -136 88 -106
<< pdiffc >>
rect -76 -106 -42 34
rect 42 -106 76 34
<< nsubdiff >>
rect -190 214 190 248
rect -190 -214 -156 214
rect 156 -214 190 214
rect -190 -248 -75 -214
rect 75 -248 190 -214
<< nsubdiffcont >>
rect -75 -248 75 -214
<< poly >>
rect -33 145 33 161
rect -33 111 -17 145
rect 17 111 33 145
rect -33 95 33 111
rect -30 64 30 95
rect -30 -162 30 -136
<< polycont >>
rect -17 111 17 145
<< locali >>
rect -33 111 -17 145
rect 17 111 33 145
rect -76 34 -42 50
rect -76 -122 -42 -106
rect 42 34 76 50
rect 42 -122 76 -106
rect -91 -248 -75 -214
rect 75 -248 91 -214
<< viali >>
rect -17 111 17 145
rect -76 -106 -42 34
rect 42 -89 76 17
<< metal1 >>
rect -30 145 30 156
rect -30 111 -17 145
rect 17 111 30 145
rect -30 100 30 111
rect -82 34 -36 46
rect -82 -106 -76 34
rect -42 -106 -36 34
rect 36 17 82 29
rect 36 -89 42 17
rect 76 -89 82 17
rect 36 -101 82 -89
rect -82 -118 -36 -106
<< labels >>
flabel viali -58 -34 -58 -34 0 FreeSans 480 0 0 0 D
port 0 nsew
flabel viali 60 -36 60 -36 0 FreeSans 480 0 0 0 S
port 1 nsew
flabel viali 0 128 0 128 0 FreeSans 480 0 0 0 G
port 2 nsew
flabel nwell -108 -262 114 -200 0 FreeSans 480 0 0 0 B
port 3 nsew
<< end >>
