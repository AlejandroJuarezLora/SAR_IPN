* NGSPICE file created from latch_temp.ext - technology: sky130B

.subckt latch vdd vss Qn S R Q
X0 Q.t0 Qn.t3 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X1 Qn.t2 a_329_215# vss.t9 vss.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X2 vss.t3 Q.t3 Qn.t0 vss.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X3 vss.t5 R.t0 a_1663_189# vss.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X4 a_329_215# S.t0 vss.t7 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X5 Q.t1 Qn.t4 vss.t1 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X6 vdd.t3 Q.t4 Qn.t1 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X7 vdd.t7 R.t1 a_1663_189# vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X8 vss.t11 a_1663_189# Q.t2 vss.t10 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
X9 a_329_215# S.t1 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
* R0 Qn.n49 Qn.t3 112.543
* R1 Qn.n50 Qn.t4 106.802
* R2 Qn.n15 Qn.t1 28.5655
* R3 Qn.n49 Qn.t2 24.7676
* R4 Qn.n39 Qn.t0 17.4005
* R5 Qn.n11 Qn.n10 13.177
* R6 Qn.n35 Qn.n34 13.177
* R7 Qn.n17 Qn.n16 9.32733
* R8 Qn.n41 Qn.n40 9.32596
* R9 Qn.n12 Qn.n11 9.3005
* R10 Qn.n5 Qn.n4 9.3005
* R11 Qn.n2 Qn.n1 9.3005
* R12 Qn.n25 Qn.n24 9.3005
* R13 Qn.n36 Qn.n35 9.3005
* R14 Qn.n29 Qn.n28 9.3005
* R15 Qn.n16 Qn.n15 9.02061
* R16 Qn.n3 Qn.n0 9.0005
* R17 Qn.n14 Qn.n13 9.0005
* R18 Qn.n38 Qn.n37 9.0005
* R19 Qn.n27 Qn.n26 9.0005
* R20 Qn.n40 Qn.n39 8.50001
* R21 Qn Qn.n48 2.98602
* R22 Qn.n42 Qn.n41 2.2535
* R23 Qn.n18 Qn.n17 2.25346
* R24 Qn.n48 Qn.n23 0.68449
* R25 Qn.n48 Qn.n47 0.660418
* R26 Qn Qn.n50 0.410826
* R27 Qn.n50 Qn.n49 0.318208
* R28 Qn.n8 Qn.n7 0.0525833
* R29 Qn.n32 Qn.n31 0.0525833
* R30 Qn.n9 Qn.n8 0.0421667
* R31 Qn.n31 Qn.n30 0.0421667
* R32 Qn.n7 Qn.n6 0.0400833
* R33 Qn.n33 Qn.n32 0.0400833
* R34 Qn.n20 Qn.n19 0.0395625
* R35 Qn.n44 Qn.n43 0.0395625
* R36 Qn.n3 Qn.n2 0.0338333
* R37 Qn.n27 Qn.n25 0.0338333
* R38 Qn.n19 Qn.n18 0.03175
* R39 Qn.n23 Qn.n22 0.03175
* R40 Qn.n45 Qn.n44 0.03175
* R41 Qn.n21 Qn.n20 0.0301875
* R42 Qn.n47 Qn.n46 0.0301875
* R43 Qn.n43 Qn.n42 0.0301875
* R44 Qn.n17 Qn.n14 0.00990809
* R45 Qn.n41 Qn.n38 0.009283
* R46 Qn.n12 Qn.n9 0.00675
* R47 Qn.n6 Qn.n5 0.00675
* R48 Qn.n22 Qn.n21 0.00675
* R49 Qn.n30 Qn.n29 0.00675
* R50 Qn.n36 Qn.n33 0.00675
* R51 Qn.n46 Qn.n45 0.00675
* R52 Qn.n14 Qn.n12 0.00258333
* R53 Qn.n5 Qn.n3 0.00258333
* R54 Qn.n29 Qn.n27 0.00258333
* R55 Qn.n38 Qn.n36 0.00258333
* R56 vdd.n125 vdd.n121 99.0123
* R57 vdd.n92 vdd.n90 95.8462
* R58 vdd.n37 vdd.n35 95.8462
* R59 vdd.n170 vdd.n168 95.8462
* R60 vdd.n171 vdd.n170 93.0272
* R61 vdd.n256 vdd.n246 92.5005
* R62 vdd.n246 vdd.n245 92.5005
* R63 vdd.n255 vdd.n254 92.5005
* R64 vdd.n252 vdd.n251 92.5005
* R65 vdd.n250 vdd.n249 92.5005
* R66 vdd.n248 vdd.n247 92.5005
* R67 vdd.n261 vdd.n260 92.5005
* R68 vdd.n235 vdd.n234 92.5005
* R69 vdd.n237 vdd.n236 92.5005
* R70 vdd.n232 vdd.n231 92.5005
* R71 vdd.n233 vdd.n232 92.5005
* R72 vdd.n213 vdd.n212 92.5005
* R73 vdd.n214 vdd.n213 92.5005
* R74 vdd.n195 vdd.n194 92.5005
* R75 vdd.n192 vdd.n191 92.5005
* R76 vdd.n193 vdd.n192 92.5005
* R77 vdd.n179 vdd.n178 92.5005
* R78 vdd.n180 vdd.n179 92.5005
* R79 vdd.n170 vdd.n169 92.5005
* R80 vdd.n168 vdd.n167 92.5005
* R81 vdd.n156 vdd.n155 92.5005
* R82 vdd.n152 vdd.n151 92.5005
* R83 vdd.n148 vdd.n147 92.5005
* R84 vdd.n144 vdd.n143 92.5005
* R85 vdd.n3 vdd.n2 92.5005
* R86 vdd.n7 vdd.n6 92.5005
* R87 vdd.n11 vdd.n10 92.5005
* R88 vdd.n15 vdd.n14 92.5005
* R89 vdd.n35 vdd.n34 92.5005
* R90 vdd.n37 vdd.n36 92.5005
* R91 vdd.n33 vdd.n32 92.5005
* R92 vdd.n39 vdd.n33 92.5005
* R93 vdd.n55 vdd.n54 92.5005
* R94 vdd.n57 vdd.n55 92.5005
* R95 vdd.n53 vdd.n52 92.5005
* R96 vdd.n74 vdd.n73 92.5005
* R97 vdd.n76 vdd.n74 92.5005
* R98 vdd.n98 vdd.n97 92.5005
* R99 vdd.n100 vdd.n98 92.5005
* R100 vdd.n92 vdd.n91 92.5005
* R101 vdd.n90 vdd.n89 92.5005
* R102 vdd.n127 vdd.n126 92.5005
* R103 vdd.n123 vdd.n122 92.5005
* R104 vdd.n108 vdd.n107 92.5005
* R105 vdd.n110 vdd.n109 92.5005
* R106 vdd.n113 vdd.n112 92.5005
* R107 vdd.n116 vdd.n115 92.5005
* R108 vdd.n121 vdd.n120 92.5005
* R109 vdd.n125 vdd.n124 92.5005
* R110 vdd.n124 vdd.n123 92.5005
* R111 vdd.n129 vdd.n128 92.5005
* R112 vdd.n128 vdd.n127 92.5005
* R113 vdd.n131 vdd.n130 92.5005
* R114 vdd.n133 vdd.n132 92.5005
* R115 vdd.n65 vdd.n64 92.5005
* R116 vdd.n21 vdd.n20 92.5005
* R117 vdd.n19 vdd.n18 92.5005
* R118 vdd.n17 vdd.n16 92.5005
* R119 vdd.n16 vdd.n15 92.5005
* R120 vdd.n13 vdd.n12 92.5005
* R121 vdd.n12 vdd.n11 92.5005
* R122 vdd.n9 vdd.n8 92.5005
* R123 vdd.n8 vdd.n7 92.5005
* R124 vdd.n5 vdd.n4 92.5005
* R125 vdd.n4 vdd.n3 92.5005
* R126 vdd.n146 vdd.n145 92.5005
* R127 vdd.n145 vdd.n144 92.5005
* R128 vdd.n150 vdd.n149 92.5005
* R129 vdd.n149 vdd.n148 92.5005
* R130 vdd.n154 vdd.n153 92.5005
* R131 vdd.n153 vdd.n152 92.5005
* R132 vdd.n158 vdd.n157 92.5005
* R133 vdd.n157 vdd.n156 92.5005
* R134 vdd.n160 vdd.n159 92.5005
* R135 vdd.n162 vdd.n161 92.5005
* R136 vdd.n203 vdd.n202 92.5005
* R137 vdd.n267 vdd.n266 92.5005
* R138 vdd.n265 vdd.n264 92.5005
* R139 vdd.n263 vdd.n262 92.5005
* R140 vdd.n262 vdd.n261 92.5005
* R141 vdd.n259 vdd.n258 92.5005
* R142 vdd.n258 vdd.n257 92.5005
* R143 vdd.n101 vdd.n92 85.9797
* R144 vdd.n58 vdd.n53 83.1607
* R145 vdd.n38 vdd.n37 81.7512
* R146 vdd.n259 vdd.n256 79.4358
* R147 vdd.n237 vdd.t4 78.9322
* R148 vdd.n238 vdd.n237 74.7038
* R149 vdd.n112 vdd.n111 72.7879
* R150 vdd.n115 vdd.n114 72.7879
* R151 vdd.n196 vdd.n195 71.8848
* R152 vdd.n35 vdd.t2 62.0183
* R153 vdd.n197 vdd.n190 60.0005
* R154 vdd.n90 vdd.t6 56.3803
* R155 vdd.n182 vdd.n166 52.9417
* R156 vdd.n239 vdd.n226 52.9417
* R157 vdd.n254 vdd.n253 52.2363
* R158 vdd.n216 vdd.n209 45.8829
* R159 vdd.n120 vdd.n119 42.8997
* R160 vdd.n71 vdd.n70 42.3534
* R161 vdd.n156 vdd.t0 39.4664
* R162 vdd.n136 vdd.t7 36.0998
* R163 vdd.n272 vdd.t5 36.065
* R164 vdd.n140 vdd.t1 36.065
* R165 vdd.n0 vdd.t3 36.065
* R166 vdd.n88 vdd.n87 35.2946
* R167 vdd.n25 vdd.n24 35.2946
* R168 vdd.n119 vdd.n118 33.0688
* R169 vdd.n118 vdd.n117 33.0686
* R170 vdd.n59 vdd.n51 31.7652
* R171 vdd.n51 vdd.n50 28.2358
* R172 vdd.n256 vdd.n255 25.6005
* R173 vdd.n255 vdd.n252 25.6005
* R174 vdd.n252 vdd.n250 25.6005
* R175 vdd.n250 vdd.n248 25.6005
* R176 vdd.n94 vdd.n93 25.6005
* R177 vdd.n95 vdd.n94 25.6005
* R178 vdd.n96 vdd.n95 25.6005
* R179 vdd.n97 vdd.n96 25.6005
* R180 vdd.n73 vdd.n72 25.6005
* R181 vdd.n32 vdd.n31 25.6005
* R182 vdd.n31 vdd.n30 25.6005
* R183 vdd.n30 vdd.n29 25.6005
* R184 vdd.n29 vdd.n28 25.6005
* R185 vdd.n28 vdd.n27 25.6005
* R186 vdd.n27 vdd.n26 25.6005
* R187 vdd.n173 vdd.n172 25.6005
* R188 vdd.n174 vdd.n173 25.6005
* R189 vdd.n175 vdd.n174 25.6005
* R190 vdd.n176 vdd.n175 25.6005
* R191 vdd.n177 vdd.n176 25.6005
* R192 vdd.n178 vdd.n177 25.6005
* R193 vdd.n212 vdd.n211 25.6005
* R194 vdd.n231 vdd.n230 25.6005
* R195 vdd.n230 vdd.n229 25.6005
* R196 vdd.n229 vdd.n228 25.6005
* R197 vdd.n121 vdd.n116 25.6005
* R198 vdd.n116 vdd.n113 25.6005
* R199 vdd.n113 vdd.n110 25.6005
* R200 vdd.n110 vdd.n108 25.6005
* R201 vdd.n129 vdd.n125 25.6005
* R202 vdd.n131 vdd.n129 25.6005
* R203 vdd.n133 vdd.n131 25.6005
* R204 vdd.n21 vdd.n19 25.6005
* R205 vdd.n19 vdd.n17 25.6005
* R206 vdd.n17 vdd.n13 25.6005
* R207 vdd.n13 vdd.n9 25.6005
* R208 vdd.n9 vdd.n5 25.6005
* R209 vdd.n150 vdd.n146 25.6005
* R210 vdd.n154 vdd.n150 25.6005
* R211 vdd.n158 vdd.n154 25.6005
* R212 vdd.n160 vdd.n158 25.6005
* R213 vdd.n162 vdd.n160 25.6005
* R214 vdd.n267 vdd.n265 25.6005
* R215 vdd.n265 vdd.n263 25.6005
* R216 vdd.n263 vdd.n259 25.6005
* R217 vdd.n163 vdd.n162 24.8476
* R218 vdd.n102 vdd.n88 24.7064
* R219 vdd.n41 vdd.n25 24.7064
* R220 vdd.n196 vdd.n193 23.9619
* R221 vdd.n22 vdd.n21 21.8358
* R222 vdd.n181 vdd.n180 21.1429
* R223 vdd.n238 vdd.n233 21.1429
* R224 vdd.n245 vdd.n244 20.1334
* R225 vdd.n215 vdd.n214 18.3239
* R226 vdd.n78 vdd.n71 17.6476
* R227 vdd.n76 vdd.n75 16.9144
* R228 vdd.t4 vdd.n235 16.9144
* R229 vdd.n134 vdd.n133 16.5652
* R230 vdd.n66 vdd.n65 15.8123
* R231 vdd.n209 vdd.n208 14.1181
* R232 vdd.n100 vdd.n99 14.0955
* R233 vdd.n39 vdd.n38 14.0955
* R234 vdd.n268 vdd.n267 13.5534
* R235 vdd.n204 vdd.n203 12.8005
* R236 vdd.n58 vdd.n57 12.686
* R237 vdd.n57 vdd.n56 11.2765
* R238 vdd.n101 vdd.n100 9.86697
* R239 vdd.n40 vdd.n39 9.86697
* R240 vdd.n269 vdd.n268 9.3005
* R241 vdd.n199 vdd.n198 9.3005
* R242 vdd.n198 vdd.n197 9.3005
* R243 vdd.n197 vdd.n196 9.3005
* R244 vdd.n184 vdd.n183 9.3005
* R245 vdd.n183 vdd.n182 9.3005
* R246 vdd.n182 vdd.n181 9.3005
* R247 vdd.n188 vdd.n187 9.3005
* R248 vdd.n186 vdd.n185 9.3005
* R249 vdd.n201 vdd.n200 9.3005
* R250 vdd.n205 vdd.n204 9.3005
* R251 vdd.n218 vdd.n217 9.3005
* R252 vdd.n217 vdd.n216 9.3005
* R253 vdd.n216 vdd.n215 9.3005
* R254 vdd.n222 vdd.n221 9.3005
* R255 vdd.n220 vdd.n219 9.3005
* R256 vdd.n243 vdd.n242 9.3005
* R257 vdd.n241 vdd.n240 9.3005
* R258 vdd.n240 vdd.n239 9.3005
* R259 vdd.n239 vdd.n238 9.3005
* R260 vdd.n47 vdd.n46 9.3005
* R261 vdd.n67 vdd.n66 9.3005
* R262 vdd.n80 vdd.n79 9.3005
* R263 vdd.n79 vdd.n78 9.3005
* R264 vdd.n78 vdd.n77 9.3005
* R265 vdd.n84 vdd.n83 9.3005
* R266 vdd.n135 vdd.n134 9.3005
* R267 vdd.n82 vdd.n81 9.3005
* R268 vdd.n106 vdd.n105 9.3005
* R269 vdd.n104 vdd.n103 9.3005
* R270 vdd.n103 vdd.n102 9.3005
* R271 vdd.n102 vdd.n101 9.3005
* R272 vdd.n61 vdd.n60 9.3005
* R273 vdd.n60 vdd.n59 9.3005
* R274 vdd.n59 vdd.n58 9.3005
* R275 vdd.n63 vdd.n62 9.3005
* R276 vdd.n45 vdd.n44 9.3005
* R277 vdd.n43 vdd.n42 9.3005
* R278 vdd.n42 vdd.n41 9.3005
* R279 vdd.n41 vdd.n40 9.3005
* R280 vdd.n166 vdd.n165 7.05932
* R281 vdd.n226 vdd.n225 7.05932
* R282 vdd.n77 vdd.n76 7.04798
* R283 vdd.n198 vdd.n189 6.4005
* R284 vdd.n183 vdd.n164 5.64756
* R285 vdd.n240 vdd.n224 5.64756
* R286 vdd.n214 vdd.n210 5.63848
* R287 vdd.n217 vdd.n207 4.89462
* R288 vdd.n273 vdd.n272 4.56717
* R289 vdd.n69 vdd.n68 4.51815
* R290 vdd.n142 vdd.n141 4.5005
* R291 vdd.n271 vdd.n270 4.5005
* R292 vdd.n86 vdd.n85 3.76521
* R293 vdd.n23 vdd.n22 3.76521
* R294 vdd.n60 vdd.n49 3.38874
* R295 vdd.n137 vdd.n136 3.1568
* R296 vdd.n49 vdd.n48 3.01226
* R297 vdd.n180 vdd.n171 2.81949
* R298 vdd.n233 vdd.n227 2.81949
* R299 vdd.n103 vdd.n86 2.63579
* R300 vdd.n42 vdd.n23 2.63579
* R301 vdd.n79 vdd.n69 1.88285
* R302 vdd.n207 vdd.n206 1.50638
* R303 vdd.n271 vdd.n142 0.88175
* R304 vdd.n139 vdd.n138 0.853625
* R305 vdd.n164 vdd.n163 0.753441
* R306 vdd.n224 vdd.n223 0.753441
* R307 vdd.n136 vdd.n135 0.42761
* R308 vdd.n270 vdd.n269 0.26925
* R309 vdd.n218 vdd.n205 0.240083
* R310 vdd.n80 vdd.n67 0.240083
* R311 vdd.n43 vdd.n1 0.179667
* R312 vdd.n199 vdd.n188 0.110917
* R313 vdd.n241 vdd.n222 0.110917
* R314 vdd.n104 vdd.n84 0.110917
* R315 vdd.n61 vdd.n47 0.110917
* R316 vdd.n138 vdd.n137 0.1005
* R317 vdd.n142 vdd.n139 0.1005
* R318 vdd.n273 vdd.n271 0.1005
* R319 vdd.n141 vdd.n140 0.0671667
* R320 vdd.n1 vdd.n0 0.0671667
* R321 vdd vdd.n273 0.04425
* R322 vdd.n201 vdd.n199 0.0338333
* R323 vdd.n186 vdd.n184 0.0296667
* R324 vdd.n243 vdd.n241 0.0296667
* R325 vdd.n220 vdd.n218 0.0255
* R326 vdd.n84 vdd.n82 0.0234167
* R327 vdd.n63 vdd.n61 0.0213333
* R328 vdd.n135 vdd.n106 0.01925
* R329 vdd.n47 vdd.n45 0.01925
* R330 vdd.n106 vdd.n104 0.0171667
* R331 vdd.n45 vdd.n43 0.0171667
* R332 vdd.n67 vdd.n63 0.0150833
* R333 vdd.n82 vdd.n80 0.013
* R334 vdd.n222 vdd.n220 0.0109167
* R335 vdd.n188 vdd.n186 0.00675
* R336 vdd.n269 vdd.n243 0.00675
* R337 vdd.n205 vdd.n201 0.00258333
* R338 Q.n50 Q.t4 112.225
* R339 Q.n49 Q.t3 107.12
* R340 Q.n15 Q.t0 28.5655
* R341 Q.n49 Q.t2 24.7676
* R342 Q.n39 Q.t1 17.4005
* R343 Q.n11 Q.n10 13.177
* R344 Q.n35 Q.n34 13.177
* R345 Q.n17 Q.n16 9.32733
* R346 Q.n41 Q.n40 9.32596
* R347 Q.n12 Q.n11 9.3005
* R348 Q.n5 Q.n4 9.3005
* R349 Q.n2 Q.n1 9.3005
* R350 Q.n25 Q.n24 9.3005
* R351 Q.n36 Q.n35 9.3005
* R352 Q.n29 Q.n28 9.3005
* R353 Q.n16 Q.n15 9.02061
* R354 Q.n3 Q.n0 9.0005
* R355 Q.n14 Q.n13 9.0005
* R356 Q.n38 Q.n37 9.0005
* R357 Q.n27 Q.n26 9.0005
* R358 Q.n40 Q.n39 8.50001
* R359 Q.n51 Q.n48 2.77388
* R360 Q.n42 Q.n41 2.2535
* R361 Q.n18 Q.n17 2.25346
* R362 Q Q.n51 1.00467
* R363 Q.n48 Q.n23 0.682942
* R364 Q.n48 Q.n47 0.660969
* R365 Q.n51 Q.n50 0.462457
* R366 Q.n50 Q.n49 0.318208
* R367 Q.n8 Q.n7 0.0525833
* R368 Q.n32 Q.n31 0.0525833
* R369 Q.n9 Q.n8 0.0421667
* R370 Q.n31 Q.n30 0.0421667
* R371 Q.n7 Q.n6 0.0400833
* R372 Q.n33 Q.n32 0.0400833
* R373 Q.n20 Q.n19 0.0395625
* R374 Q.n44 Q.n43 0.0395625
* R375 Q.n3 Q.n2 0.0338333
* R376 Q.n27 Q.n25 0.0338333
* R377 Q.n19 Q.n18 0.03175
* R378 Q.n23 Q.n22 0.03175
* R379 Q.n45 Q.n44 0.03175
* R380 Q.n21 Q.n20 0.0301875
* R381 Q.n47 Q.n46 0.0301875
* R382 Q.n43 Q.n42 0.0301875
* R383 Q.n17 Q.n14 0.00990809
* R384 Q.n41 Q.n38 0.009283
* R385 Q.n12 Q.n9 0.00675
* R386 Q.n6 Q.n5 0.00675
* R387 Q.n22 Q.n21 0.00675
* R388 Q.n30 Q.n29 0.00675
* R389 Q.n36 Q.n33 0.00675
* R390 Q.n46 Q.n45 0.00675
* R391 Q.n14 Q.n12 0.00258333
* R392 Q.n5 Q.n3 0.00258333
* R393 Q.n29 Q.n27 0.00258333
* R394 Q.n38 Q.n36 0.00258333
* R395 vss.n12 vss.n11 403.438
* R396 vss.n143 vss.n142 403.438
* R397 vss.n14 vss.n13 394
* R398 vss.n147 vss.n144 394
* R399 vss.n324 vss.n323 371.921
* R400 vss.n245 vss.n244 359.312
* R401 vss.n204 vss.n203 346.705
* R402 vss.n34 vss.n30 334.098
* R403 vss.n97 vss.n93 334.098
* R404 vss.n124 vss.n123 334.098
* R405 vss.n167 vss.n166 334.098
* R406 vss.n62 vss.n61 292.5
* R407 vss.n60 vss.n59 292.5
* R408 vss.n56 vss.n55 292.5
* R409 vss.n54 vss.n53 292.5
* R410 vss.n52 vss.n51 292.5
* R411 vss.n50 vss.n49 292.5
* R412 vss.n48 vss.n47 292.5
* R413 vss.n30 vss.n29 292.5
* R414 vss.n33 vss.n32 292.5
* R415 vss.n15 vss.n14 292.5
* R416 vss.n93 vss.n92 292.5
* R417 vss.n96 vss.n95 292.5
* R418 vss.n120 vss.n119 292.5
* R419 vss.n121 vss.n120 292.5
* R420 vss.n123 vss.n122 292.5
* R421 vss.n147 vss.n146 292.5
* R422 vss.n148 vss.n147 292.5
* R423 vss.n163 vss.n162 292.5
* R424 vss.n164 vss.n163 292.5
* R425 vss.n166 vss.n165 292.5
* R426 vss.n184 vss.n183 292.5
* R427 vss.n185 vss.n184 292.5
* R428 vss.n201 vss.n200 292.5
* R429 vss.n203 vss.n202 292.5
* R430 vss.n227 vss.n226 292.5
* R431 vss.n242 vss.n241 292.5
* R432 vss.n244 vss.n243 292.5
* R433 vss.n267 vss.n266 292.5
* R434 vss.n321 vss.n320 292.5
* R435 vss.n323 vss.n322 292.5
* R436 vss.n290 vss.n289 292.5
* R437 vss.n292 vss.n291 292.5
* R438 vss.n295 vss.n294 292.5
* R439 vss.n294 vss.n293 292.5
* R440 vss.n298 vss.n297 292.5
* R441 vss.n300 vss.n299 292.5
* R442 vss.n304 vss.n303 292.5
* R443 vss.n307 vss.n306 292.5
* R444 vss.n306 vss.n305 292.5
* R445 vss.n310 vss.n309 292.5
* R446 vss.n309 vss.n308 292.5
* R447 vss.n312 vss.n311 292.5
* R448 vss.n252 vss.n251 292.5
* R449 vss.n133 vss.n132 292.5
* R450 vss.n4 vss.n3 292.5
* R451 vss.n2 vss.n1 292.5
* R452 vss.n135 vss.n134 292.5
* R453 vss.n174 vss.n173 292.5
* R454 vss.n210 vss.n209 292.5
* R455 vss.n76 vss.n75 292.5
* R456 vss.n74 vss.n73 292.5
* R457 vss.n73 vss.n72 292.5
* R458 vss.n71 vss.n70 292.5
* R459 vss.n70 vss.n69 292.5
* R460 vss.n68 vss.n67 292.5
* R461 vss.n67 vss.n66 292.5
* R462 vss.n65 vss.n64 292.5
* R463 vss.n64 vss.n63 292.5
* R464 vss.n265 vss.t8 226.935
* R465 vss.n66 vss.t4 201.72
* R466 vss.n56 vss.n54 156.236
* R467 vss.n307 vss.n304 156.236
* R468 vss.n65 vss.n62 144.189
* R469 vss.n298 vss.n295 142.683
* R470 vss.n302 vss.n301 134.577
* R471 vss.n59 vss.n58 117.719
* R472 vss.n199 vss.t0 100.861
* R473 vss.n34 vss.n33 94.5564
* R474 vss.n97 vss.n96 94.5564
* R475 vss.n124 vss.n121 94.5564
* R476 vss.n167 vss.n164 94.5564
* R477 vss.n297 vss.n296 90.6381
* R478 vss.n303 vss.n302 90.6381
* R479 vss.n117 vss.t2 88.2527
* R480 vss.n58 vss.n57 87.3925
* R481 vss.n35 vss.n28 86.9123
* R482 vss.n98 vss.n91 86.9123
* R483 vss.n125 vss.n116 86.9123
* R484 vss.n168 vss.n160 86.9123
* R485 vss.n16 vss.n15 81.9489
* R486 vss.n149 vss.n148 81.9489
* R487 vss.n204 vss.n201 81.9489
* R488 vss.n17 vss.n10 75.324
* R489 vss.n150 vss.n141 75.324
* R490 vss.n205 vss.n198 75.324
* R491 vss.n186 vss.n185 69.3415
* R492 vss.n245 vss.n242 69.3415
* R493 vss.n187 vss.n180 63.7358
* R494 vss.n246 vss.n239 63.7358
* R495 vss.n267 vss.n265 63.0378
* R496 vss.n264 vss.n263 57.9417
* R497 vss.n228 vss.n227 56.734
* R498 vss.n324 vss.n321 56.734
* R499 vss.n229 vss.n224 52.1476
* R500 vss.n325 vss.n318 52.1476
* R501 vss.n31 vss.t10 50.4303
* R502 vss.n227 vss.n225 50.4303
* R503 vss.n321 vss.n319 50.4303
* R504 vss.n224 vss.n223 46.3534
* R505 vss.n318 vss.n317 46.3534
* R506 vss.n268 vss.n267 44.1266
* R507 vss.n269 vss.n264 40.5593
* R508 vss.n185 vss.n181 37.8228
* R509 vss.n242 vss.n240 37.8228
* R510 vss.n180 vss.n179 34.7652
* R511 vss.n239 vss.n238 34.7652
* R512 vss.n60 vss.n56 25.6005
* R513 vss.n62 vss.n60 25.6005
* R514 vss.n54 vss.n52 25.6005
* R515 vss.n52 vss.n50 25.6005
* R516 vss.n50 vss.n48 25.6005
* R517 vss.n48 vss.n46 25.6005
* R518 vss.n46 vss.n45 25.6005
* R519 vss.n45 vss.n44 25.6005
* R520 vss.n44 vss.n43 25.6005
* R521 vss.n43 vss.n42 25.6005
* R522 vss.n42 vss.n41 25.6005
* R523 vss.n119 vss.n118 25.6005
* R524 vss.n146 vss.n145 25.6005
* R525 vss.n183 vss.n182 25.6005
* R526 vss.n282 vss.n281 25.6005
* R527 vss.n283 vss.n282 25.6005
* R528 vss.n284 vss.n283 25.6005
* R529 vss.n285 vss.n284 25.6005
* R530 vss.n286 vss.n285 25.6005
* R531 vss.n287 vss.n286 25.6005
* R532 vss.n288 vss.n287 25.6005
* R533 vss.n290 vss.n288 25.6005
* R534 vss.n292 vss.n290 25.6005
* R535 vss.n295 vss.n292 25.6005
* R536 vss.n300 vss.n298 25.6005
* R537 vss.n304 vss.n300 25.6005
* R538 vss.n68 vss.n65 25.6005
* R539 vss.n71 vss.n68 25.6005
* R540 vss.n74 vss.n71 25.6005
* R541 vss.n76 vss.n74 25.6005
* R542 vss.n312 vss.n310 25.6005
* R543 vss.n310 vss.n307 25.6005
* R544 vss.n15 vss.n12 25.2154
* R545 vss.n148 vss.n143 25.2154
* R546 vss.n201 vss.n199 25.2154
* R547 vss.n305 vss.t6 25.2154
* R548 vss.n81 vss.t5 24.7712
* R549 vss.n273 vss.t9 24.5445
* R550 vss.n80 vss.t11 24.5445
* R551 vss.n101 vss.t3 24.5445
* R552 vss.n208 vss.t1 24.5445
* R553 vss.n279 vss.t7 24.5445
* R554 vss.n10 vss.n9 23.177
* R555 vss.n141 vss.n140 23.177
* R556 vss.n198 vss.n197 23.177
* R557 vss.n313 vss.n312 15.8123
* R558 vss.n253 vss.n252 15.0593
* R559 vss.n211 vss.n210 14.3064
* R560 vss.n77 vss.n76 13.5534
* R561 vss.n175 vss.n174 13.5534
* R562 vss.n5 vss.n2 12.8005
* R563 vss.n5 vss.n4 12.8005
* R564 vss.n136 vss.n133 12.8005
* R565 vss.n136 vss.n135 12.8005
* R566 vss.n33 vss.n31 12.608
* R567 vss.n96 vss.n94 12.608
* R568 vss.n121 vss.n117 12.608
* R569 vss.n164 vss.n161 12.608
* R570 vss.n28 vss.n27 11.5887
* R571 vss.n91 vss.n90 11.5887
* R572 vss.n116 vss.n115 11.5887
* R573 vss.n160 vss.n159 11.5887
* R574 vss.n78 vss.n77 9.3005
* R575 vss.n275 vss.n274 9.3005
* R576 vss.n273 vss.n272 9.3005
* R577 vss.n235 vss.n234 9.3005
* R578 vss.n212 vss.n211 9.3005
* R579 vss.n170 vss.n169 9.3005
* R580 vss.n169 vss.n168 9.3005
* R581 vss.n168 vss.n167 9.3005
* R582 vss.n105 vss.n104 9.3005
* R583 vss.n23 vss.n22 9.3005
* R584 vss.n21 vss.n20 9.3005
* R585 vss.n19 vss.n18 9.3005
* R586 vss.n18 vss.n17 9.3005
* R587 vss.n17 vss.n16 9.3005
* R588 vss.n103 vss.n102 9.3005
* R589 vss.n100 vss.n99 9.3005
* R590 vss.n99 vss.n98 9.3005
* R591 vss.n98 vss.n97 9.3005
* R592 vss.n127 vss.n126 9.3005
* R593 vss.n126 vss.n125 9.3005
* R594 vss.n125 vss.n124 9.3005
* R595 vss.n131 vss.n130 9.3005
* R596 vss.n129 vss.n128 9.3005
* R597 vss.n152 vss.n151 9.3005
* R598 vss.n151 vss.n150 9.3005
* R599 vss.n150 vss.n149 9.3005
* R600 vss.n156 vss.n155 9.3005
* R601 vss.n154 vss.n153 9.3005
* R602 vss.n172 vss.n171 9.3005
* R603 vss.n176 vss.n175 9.3005
* R604 vss.n189 vss.n188 9.3005
* R605 vss.n188 vss.n187 9.3005
* R606 vss.n187 vss.n186 9.3005
* R607 vss.n193 vss.n192 9.3005
* R608 vss.n191 vss.n190 9.3005
* R609 vss.n207 vss.n206 9.3005
* R610 vss.n206 vss.n205 9.3005
* R611 vss.n205 vss.n204 9.3005
* R612 vss.n233 vss.n232 9.3005
* R613 vss.n231 vss.n230 9.3005
* R614 vss.n230 vss.n229 9.3005
* R615 vss.n229 vss.n228 9.3005
* R616 vss.n248 vss.n247 9.3005
* R617 vss.n247 vss.n246 9.3005
* R618 vss.n246 vss.n245 9.3005
* R619 vss.n254 vss.n253 9.3005
* R620 vss.n250 vss.n249 9.3005
* R621 vss.n270 vss.n269 9.3005
* R622 vss.n269 vss.n268 9.3005
* R623 vss.n327 vss.n326 9.3005
* R624 vss.n326 vss.n325 9.3005
* R625 vss.n325 vss.n324 9.3005
* R626 vss.n314 vss.n313 9.3005
* R627 vss.n316 vss.n315 9.3005
* R628 vss.n37 vss.n36 9.3005
* R629 vss.n36 vss.n35 9.3005
* R630 vss.n35 vss.n34 9.3005
* R631 vss.n331 vss.n330 9.0005
* R632 vss.n277 vss.n276 9.0005
* R633 vss.n107 vss.n106 9.0005
* R634 vss.n214 vss.n213 9.0005
* R635 vss.n40 vss.n39 9.0005
* R636 vss.n36 vss.n26 5.64756
* R637 vss.n99 vss.n89 5.64756
* R638 vss.n126 vss.n114 5.64756
* R639 vss.n169 vss.n158 5.64756
* R640 vss.n18 vss.n8 4.89462
* R641 vss.n151 vss.n139 4.89462
* R642 vss.n206 vss.n196 4.89462
* R643 vss.n6 vss.n5 4.6505
* R644 vss.n137 vss.n136 4.6505
* R645 vss.n271 vss.n270 4.57427
* R646 vss.n188 vss.n178 4.14168
* R647 vss.n247 vss.n237 4.14168
* R648 vss.n262 vss.n261 3.76521
* R649 vss.n230 vss.n222 3.38874
* R650 vss.n222 vss.n221 3.01226
* R651 vss.n329 vss.n328 3.01226
* R652 vss.n109 vss.n108 3.0005
* R653 vss.n216 vss.n215 3.0005
* R654 vss.n257 vss.n256 3.0005
* R655 vss.n333 vss.n332 3.0005
* R656 vss.n270 vss.n262 2.63579
* R657 vss.n330 vss.n329 2.63579
* R658 vss.n178 vss.n177 2.25932
* R659 vss.n237 vss.n236 2.25932
* R660 vss.n82 vss.n81 1.61892
* R661 vss.n8 vss.n7 1.50638
* R662 vss.n139 vss.n138 1.50638
* R663 vss.n196 vss.n195 1.50638
* R664 vss.n112 vss.n111 0.827063
* R665 vss.n26 vss.n25 0.753441
* R666 vss.n89 vss.n88 0.753441
* R667 vss.n114 vss.n113 0.753441
* R668 vss.n158 vss.n157 0.753441
* R669 vss.n314 vss.n280 0.440083
* R670 vss.n81 vss.n80 0.390712
* R671 vss.n219 vss.n218 0.3755
* R672 vss.n335 vss.n334 0.359875
* R673 vss.n86 vss.n85 0.341125
* R674 vss.n19 vss.n6 0.240083
* R675 vss.n152 vss.n137 0.240083
* R676 vss.n189 vss.n176 0.240083
* R677 vss.n255 vss.n254 0.185917
* R678 vss.n137 vss.n131 0.146333
* R679 vss.n231 vss.n220 0.133833
* R680 vss.n170 vss.n156 0.110917
* R681 vss.n248 vss.n235 0.110917
* R682 vss.n336 vss.n335 0.1005
* R683 vss.n24 vss.n23 0.09425
* R684 vss.n218 vss.n217 0.0864375
* R685 vss.n6 vss.n0 0.0859167
* R686 vss.n194 vss.n193 0.0838333
* R687 vss.n111 vss.n110 0.078625
* R688 vss.n280 vss.n279 0.0671667
* R689 vss.n100 vss.n87 0.063
* R690 vss vss.n336 0.04425
* R691 vss.n278 vss.n277 0.0421667
* R692 vss.n332 vss.n331 0.0421667
* R693 vss.n212 vss.n208 0.0400833
* R694 vss.n79 vss.n78 0.038
* R695 vss.n259 vss.n258 0.0364375
* R696 vss.n273 vss.n271 0.0338333
* R697 vss.n129 vss.n127 0.03175
* R698 vss.n172 vss.n170 0.03175
* R699 vss.n327 vss.n316 0.03175
* R700 vss.n83 vss.n82 0.03175
* R701 vss.n85 vss.n84 0.03175
* R702 vss.n260 vss.n259 0.03175
* R703 vss.n334 vss.n333 0.03175
* R704 vss.n108 vss.n107 0.0296667
* R705 vss.n105 vss.n103 0.0296667
* R706 vss.n21 vss.n19 0.0275833
* R707 vss.n154 vss.n152 0.0275833
* R708 vss.n207 vss.n194 0.0275833
* R709 vss.n216 vss.n112 0.0270625
* R710 vss.n38 vss.n37 0.0255
* R711 vss.n258 vss.n257 0.0255
* R712 vss.n191 vss.n189 0.0234167
* R713 vss.n250 vss.n248 0.0234167
* R714 vss.n110 vss.n109 0.022375
* R715 vss.n256 vss.n255 0.0213333
* R716 vss.n80 vss.n79 0.01925
* R717 vss.n215 vss.n214 0.01925
* R718 vss.n233 vss.n231 0.01925
* R719 vss.n109 vss.n86 0.01925
* R720 vss.n37 vss.n24 0.0171667
* R721 vss.n235 vss.n233 0.0171667
* R722 vss.n257 vss.n219 0.016125
* R723 vss.n217 vss.n216 0.0145625
* R724 vss.n193 vss.n191 0.013
* R725 vss.n254 vss.n250 0.013
* R726 vss.n277 vss.n275 0.013
* R727 vss.n332 vss.n278 0.0109167
* R728 vss.n23 vss.n21 0.00883333
* R729 vss.n156 vss.n154 0.00883333
* R730 vss.n215 vss.n207 0.00883333
* R731 vss.n214 vss.n212 0.00883333
* R732 vss.n333 vss.n260 0.0083125
* R733 vss.n40 vss.n38 0.00675
* R734 vss.n107 vss.n105 0.00675
* R735 vss.n84 vss.n83 0.0051875
* R736 vss.n78 vss.n40 0.00466667
* R737 vss.n101 vss.n100 0.00466667
* R738 vss.n131 vss.n129 0.00466667
* R739 vss.n176 vss.n172 0.00466667
* R740 vss.n331 vss.n327 0.00466667
* R741 vss.n316 vss.n314 0.00466667
* R742 vss.n103 vss.n101 0.00258333
* R743 vss.n275 vss.n273 0.00258333
* R744 R.n0 R.t1 112.543
* R745 R.n0 R.t0 107.12
* R746 R R.n0 0.354667
* R747 S.n0 S.t1 112.543
* R748 S.n0 S.t0 107.12
* R749 S S.n0 0.417167
* C0 Q a_329_215# 0.0695f
* C1 Qn S 0.0154f
* C2 vdd a_1663_189# 0.382f
* C3 R vdd 0.319f
* C4 Qn vdd 0.55f
* C5 Qn a_329_215# 0.117f
* C6 vdd S 0.321f
* C7 Q a_1663_189# 0.117f
* C8 R Q 0.0155f
* C9 Qn Q 0.827f
* C10 S a_329_215# 0.149f
* C11 vdd a_329_215# 0.381f
* C12 R a_1663_189# 0.149f
* C13 Qn a_1663_189# 0.0695f
* C14 Q S 1.46e-19
* C15 Q vdd 0.815f
.ends

