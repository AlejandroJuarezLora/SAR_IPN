magic
tech sky130B
timestamp 1696364841
<< metal4 >>
rect -5 119 315 140
rect -5 1 16 119
rect 134 1 176 119
rect 294 1 315 119
rect -5 -20 315 1
<< via4 >>
rect 16 1 134 119
rect 176 1 294 119
<< metal5 >>
rect -5 119 315 140
rect -5 1 16 119
rect 134 1 176 119
rect 294 1 315 119
rect -5 -20 315 1
<< end >>
