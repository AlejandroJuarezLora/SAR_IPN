magic
tech sky130B
magscale 1 2
timestamp 1697741630
<< pwell >>
rect 1564 -377 1600 -133
rect 1144 -411 1602 -377
rect 1564 -468 1600 -411
<< nsubdiffcont >>
rect 1362 915 1398 1660
<< locali >>
rect 1358 1660 1410 2120
rect 1358 1630 1362 1660
rect 1252 1578 1362 1630
rect 1352 1262 1362 1578
rect 1252 1210 1362 1262
rect 1356 973 1362 1210
rect 1256 921 1362 973
rect 1358 915 1362 921
rect 1398 1630 1410 1660
rect 1398 1578 1520 1630
rect 1398 1262 1410 1578
rect 1398 1210 1516 1262
rect 1398 973 1410 1210
rect 1398 921 1512 973
rect 1398 915 1410 921
rect 1358 867 1410 915
rect 950 -682 993 353
rect 1307 -109 1341 -41
rect 1424 -111 1459 -43
rect 1084 -682 1127 -577
rect 1503 -682 1546 -582
rect 950 -725 1546 -682
rect 950 -1883 993 -725
rect -169 -1926 2869 -1883
<< metal1 >>
rect -1769 2956 -1677 3006
rect 4384 2933 4495 2983
rect -1776 2222 -1686 2266
rect 4392 2199 4474 2243
rect 1181 1784 1233 1790
rect -1805 1703 -1690 1749
rect 1233 1743 1594 1773
rect 1181 1726 1233 1732
rect 4392 1680 4489 1726
rect 782 1614 1159 1643
rect 1621 1609 1920 1638
rect 1178 1422 1230 1428
rect 1230 1381 1601 1411
rect 1178 1364 1230 1370
rect -1772 615 -1686 659
rect 1098 582 1130 1198
rect 1630 882 1662 1212
rect 1616 852 1662 882
rect 1620 850 1662 852
rect 1172 752 1340 786
rect 1430 784 1462 786
rect 1428 754 1582 784
rect 1308 700 1340 752
rect 1298 694 1350 700
rect 1298 636 1350 642
rect 1088 576 1140 582
rect 1088 518 1140 524
rect 1098 438 1130 518
rect 1308 374 1340 636
rect 1430 582 1462 754
rect 1630 694 1662 850
rect 1614 642 1620 694
rect 1672 642 1678 694
rect 1424 576 1476 582
rect 1424 518 1476 524
rect 1430 352 1462 518
rect 1630 448 1662 642
rect 4382 592 4466 636
rect 1141 174 1179 331
rect 782 145 1179 174
rect 1580 148 1618 328
rect 1141 -7 1179 145
rect 1566 119 1920 148
rect 1580 -10 1618 119
rect 1142 -377 1178 -130
rect 1564 -377 1600 -133
rect 1142 -411 1602 -377
rect 1142 -465 1178 -411
rect 1564 -468 1600 -411
rect 1293 -512 1345 -506
rect 1345 -553 1453 -523
rect 1293 -570 1345 -564
rect -1775 -627 -1690 -581
rect 4391 -650 4477 -604
<< via1 >>
rect 1181 1732 1233 1784
rect 1178 1370 1230 1422
rect 1298 642 1350 694
rect 1088 524 1140 576
rect 1620 642 1672 694
rect 1424 524 1476 576
rect 1293 -564 1345 -512
<< metal2 >>
rect 951 1773 981 2164
rect 1175 1773 1181 1784
rect 951 1743 1181 1773
rect 951 1411 981 1743
rect 1175 1732 1181 1743
rect 1233 1732 1239 1784
rect 1172 1411 1178 1422
rect 951 1381 1178 1411
rect 951 -523 981 1381
rect 1172 1370 1178 1381
rect 1230 1370 1236 1422
rect 1620 694 1672 700
rect 1292 642 1298 694
rect 1350 684 1356 694
rect 1350 652 1620 684
rect 1350 642 1356 652
rect 1620 636 1672 642
rect 1082 524 1088 576
rect 1140 566 1146 576
rect 1418 566 1424 576
rect 1140 534 1424 566
rect 1140 524 1146 534
rect 1418 524 1424 534
rect 1476 524 1482 576
rect 1287 -523 1293 -512
rect 951 -553 1293 -523
rect 1287 -564 1293 -553
rect 1345 -564 1351 -512
use sky130_fd_pr__nfet_01v8_7UX3DE  sky130_fd_pr__nfet_01v8_7UX3DE_0
timestamp 1696715056
transform 0 1 1373 -1 0 -534
box -226 -457 226 457
use sky130_fd_pr__nfet_01v8_7UX3DE  sky130_fd_pr__nfet_01v8_7UX3DE_1
timestamp 1696715056
transform 0 1 1381 -1 0 384
box -226 -457 226 457
use sky130_fd_pr__nfet_01v8_7UX3DE  sky130_fd_pr__nfet_01v8_7UX3DE_2
timestamp 1696715056
transform 0 1 1378 -1 0 -76
box -226 -457 226 457
use sky130_fd_pr__pfet_01v8_QE5SNW  sky130_fd_pr__pfet_01v8_QE5SNW_0
timestamp 1696717065
transform -1 0 1574 0 1 1269
box -226 -649 226 649
use sky130_fd_pr__pfet_01v8_QE5SNW  sky130_fd_pr__pfet_01v8_QE5SNW_1
timestamp 1696717065
transform 1 0 1195 0 1 1269
box -226 -649 226 649
use trim  trim_0
timestamp 1696628412
transform 0 -1 -677 1 0 2433
box -4358 -1541 573 1059
use trim  trim_1
timestamp 1696628412
transform 0 1 3379 1 0 2410
box -4358 -1541 573 1059
<< labels >>
flabel metal1 1098 438 1130 1198 0 FreeSans 640 0 0 0 outn
port 13 nsew
flabel metal1 1630 448 1662 1212 0 FreeSans 640 0 0 0 outp
port 12 nsew
flabel metal1 1580 -10 1618 328 0 FreeSans 640 0 0 0 ip
flabel metal1 1141 -7 1179 331 0 FreeSans 640 0 0 0 in
flabel metal1 1144 -411 1602 -377 0 FreeSans 640 0 0 0 diff
flabel locali 950 -875 993 -832 0 FreeSans 640 0 0 0 vss
port 16 nsew
flabel locali 1358 1929 1410 1981 0 FreeSans 640 0 0 0 vdd
port 15 nsew
flabel metal2 951 2134 981 2164 0 FreeSans 640 0 0 0 clk
port 14 nsew
flabel locali 1440 -83 1440 -83 0 FreeSans 640 0 0 0 vp
port 10 nsew
flabel locali 1322 -81 1322 -81 0 FreeSans 640 0 0 0 vn
port 11 nsew
flabel metal1 -1775 -627 -1690 -581 0 FreeSans 800 0 0 0 trim_4
port 0 nsew
flabel metal1 -1772 615 -1728 659 0 FreeSans 800 0 0 0 trim_3
port 1 nsew
flabel metal1 -1805 1703 -1759 1749 0 FreeSans 800 0 0 0 trim_2
port 2 nsew
flabel metal1 -1776 2222 -1732 2266 0 FreeSans 800 0 0 0 trim_1
port 3 nsew
flabel metal1 -1769 2956 -1719 3006 0 FreeSans 800 0 0 0 trim_0
port 4 nsew
flabel metal1 4431 -650 4477 -604 0 FreeSans 800 0 0 0 trimb_4
port 5 nsew
flabel metal1 4422 592 4466 636 0 FreeSans 800 0 0 0 trimb_3
port 6 nsew
flabel metal1 4443 1680 4489 1726 0 FreeSans 800 0 0 0 trimb_2
port 7 nsew
flabel metal1 4430 2199 4474 2243 0 FreeSans 800 0 0 0 trimb_1
port 8 nsew
flabel metal1 4445 2933 4495 2983 0 FreeSans 800 0 0 0 trimb_0
port 9 nsew
<< end >>
