* SPICE3 file created from comparator.ext - technology: sky130B

.subckt M1_1 a_30_n109# a_n88_n109# a_n33_n197# VSUBS
X0 a_30_n109# a_n33_n197# a_n88_n109# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n109# a_n88_n109# 0.121f
C1 a_30_n109# a_n33_n197# 0.0116f
C2 a_n88_n109# a_n33_n197# 0.0116f
C3 a_30_n109# VSUBS 0.121f
C4 a_n88_n109# VSUBS 0.121f
C5 a_n33_n197# VSUBS 0.227f
.ends

.subckt trim_sw d_0 d_1 d_2 d_3 d_4 m1_1462_409# m1_1771_409# m1_799_409# m1_1226_409#
+ m1_136_409# vss
XM1_1_14 vss m1_799_409# d_2 vss M1_1
XM1_1_15 m1_799_409# vss d_2 vss M1_1
XM1_1_0 vss m1_1226_409# d_0 vss M1_1
XM1_1_1 vss m1_1771_409# d_4 vss M1_1
XM1_1_2 m1_1771_409# vss d_4 vss M1_1
XM1_1_3 vss m1_1771_409# d_4 vss M1_1
XM1_1_4 m1_1771_409# vss d_4 vss M1_1
XM1_1_5 m1_1771_409# vss d_4 vss M1_1
XM1_1_6 vss m1_1771_409# d_4 vss M1_1
XM1_1_7 vss m1_1771_409# d_4 vss M1_1
XM1_1_8 m1_1771_409# vss d_4 vss M1_1
XM1_1_9 m1_1462_409# vss d_1 vss M1_1
XM1_1_10 m1_136_409# vss d_3 vss M1_1
XM1_1_11 vss m1_136_409# d_3 vss M1_1
XM1_1_12 m1_136_409# vss d_3 vss M1_1
XM1_1_13 vss m1_136_409# d_3 vss M1_1
C0 d_3 m1_799_409# 1.67e-19
C1 m1_1226_409# m1_1462_409# 0.0249f
C2 d_0 m1_799_409# 1.67e-19
C3 m1_1226_409# d_0 0.0315f
C4 vss m1_136_409# 0.662f
C5 m1_136_409# m1_799_409# 0.153f
C6 m1_136_409# d_3 0.067f
C7 d_4 m1_1771_409# 0.165f
C8 vss m1_1771_409# 0.926f
C9 vss d_2 0.146f
C10 m1_1462_409# m1_1771_409# 0.0191f
C11 d_2 m1_799_409# 0.0168f
C12 m1_1226_409# d_2 1.67e-19
C13 d_3 d_2 0.0446f
C14 d_4 d_1 0.0454f
C15 d_4 vss 0.446f
C16 vss d_1 0.0796f
C17 d_0 d_2 0.0764f
C18 vss m1_799_409# 0.297f
C19 m1_1226_409# vss 0.133f
C20 m1_136_409# d_2 1.67e-19
C21 d_4 m1_1462_409# 1.67e-19
C22 vss d_3 0.262f
C23 m1_1462_409# d_1 0.0315f
C24 vss m1_1462_409# 0.259f
C25 d_1 d_0 0.113f
C26 vss d_0 0.0759f
C27 m1_1226_409# m1_799_409# 0.153f
C28 d_2 0 0.362f
C29 m1_136_409# 0 0.38f
C30 vss 0 1f
C31 d_3 0 0.702f
C32 m1_1462_409# 0 0.0797f
C33 d_1 0 0.239f
C34 m1_1771_409# 0 0.401f
C35 d_4 0 1.29f
C36 m1_1226_409# 0 0.0757f
C37 d_0 0 0.227f
C38 m1_799_409# 0 0.219f
.ends

.subckt trim n1 n0 trim_sw_0/d_4 trim_sw_0/d_3 trim_sw_0/d_2 trim_sw_0/d_1 trim_sw_0/d_0
+ n2 n4 VSUBS drain n3
Xtrim_sw_0 trim_sw_0/d_0 trim_sw_0/d_1 trim_sw_0/d_2 trim_sw_0/d_3 trim_sw_0/d_4 n1
+ n4 n2 n0 n3 VSUBS trim_sw
C0 n3 trim_sw_0/d_2 9.86e-20
C1 n3 VSUBS 0.112f
C2 trim_sw_0/d_1 n2 0.00217f
C3 n4 drain 6.84f
C4 n1 drain 0.851f
C5 n3 drain 3.41f
C6 n2 n0 0.0935f
C7 trim_sw_0/d_0 n0 0.0074f
C8 n4 trim_sw_0/d_1 2.85e-20
C9 n1 trim_sw_0/d_1 0.0074f
C10 n4 trim_sw_0/d_3 6.08e-20
C11 n3 trim_sw_0/d_1 4.93e-20
C12 n4 n0 0.138f
C13 n1 n0 0.482f
C14 n3 trim_sw_0/d_3 2.03e-19
C15 drain trim_sw_0/d_2 2.61e-20
C16 n3 n0 0.077f
C17 drain VSUBS 1.76f
C18 n2 trim_sw_0/d_4 0.00497f
C19 n2 trim_sw_0/d_0 0.00217f
C20 trim_sw_0/d_3 VSUBS 6.59e-20
C21 n4 trim_sw_0/d_4 5.87e-19
C22 VSUBS n0 0.0281f
C23 trim_sw_0/d_3 drain 1.1e-19
C24 n3 trim_sw_0/d_4 4.9e-19
C25 n4 n2 0.551f
C26 n1 n2 0.0775f
C27 drain n0 0.851f
C28 n3 n2 0.517f
C29 n4 trim_sw_0/d_0 2.85e-20
C30 n3 trim_sw_0/d_0 4.93e-20
C31 n4 n1 0.145f
C32 n3 n4 1.35f
C33 n3 n1 0.0769f
C34 VSUBS trim_sw_0/d_4 1.43e-19
C35 n2 trim_sw_0/d_2 6e-19
C36 n2 VSUBS 0.0679f
C37 drain trim_sw_0/d_4 2.61e-20
C38 n2 drain 1.7f
C39 n4 trim_sw_0/d_2 1.61e-19
C40 n4 VSUBS 0.192f
C41 n1 VSUBS 0.0284f
C42 n1 0 0.237f
C43 n0 0 0.224f
C44 drain 0 -4.84f
C45 trim_sw_0/d_2 0 0.362f
C46 n3 0 1.39f
C47 VSUBS 0 1.65f
C48 trim_sw_0/d_3 0 0.702f
C49 trim_sw_0/d_1 0 0.239f
C50 n4 0 1.98f
C51 trim_sw_0/d_4 0 1.29f
C52 trim_sw_0/d_0 0 0.227f
C53 n2 0 0.746f
.ends

.subckt Mdiff a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n171# a_n33_51# 0.0116f
C1 a_30_n171# a_n88_n171# 0.121f
C2 a_n88_n171# a_n33_51# 0.0116f
C3 a_30_n171# VSUBS 0.121f
C4 a_n88_n171# VSUBS 0.121f
C5 a_n33_51# VSUBS 0.227f
.ends

.subckt M3 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n33_55# a_30_n176# 0.0116f
C1 a_n88_n176# w_n124_n238# 0.00827f
C2 a_n88_n176# a_n33_55# 0.0116f
C3 a_n33_55# w_n124_n238# 0.0663f
C4 a_n88_n176# a_30_n176# 0.121f
C5 a_30_n176# w_n124_n238# 0.00827f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt Ml1 a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n171# a_n33_51# 0.0116f
C1 a_30_n171# a_n88_n171# 0.121f
C2 a_n88_n171# a_n33_51# 0.0116f
C3 a_30_n171# VSUBS 0.121f
C4 a_n88_n171# VSUBS 0.121f
C5 a_n33_51# VSUBS 0.227f
.ends

.subckt Minp a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n171# a_n33_51# 0.0116f
C1 a_30_n171# a_n88_n171# 0.121f
C2 a_n88_n171# a_n33_51# 0.0116f
C3 a_30_n171# VSUBS 0.121f
C4 a_n88_n171# VSUBS 0.121f
C5 a_n33_51# VSUBS 0.227f
.ends

.subckt M1 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n33_55# a_30_n176# 0.0116f
C1 a_n88_n176# w_n124_n238# 0.00827f
C2 a_n88_n176# a_n33_55# 0.0116f
C3 a_n33_55# w_n124_n238# 0.0663f
C4 a_n88_n176# a_30_n176# 0.121f
C5 a_30_n176# w_n124_n238# 0.00827f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt Minn a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n171# a_n33_51# 0.0116f
C1 a_30_n171# a_n88_n171# 0.121f
C2 a_n88_n171# a_n33_51# 0.0116f
C3 a_30_n171# VSUBS 0.121f
C4 a_n88_n171# VSUBS 0.121f
C5 a_n33_51# VSUBS 0.227f
.ends

.subckt Ml4 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n33_55# a_30_n176# 0.0116f
C1 a_n88_n176# w_n124_n238# 0.00827f
C2 a_n88_n176# a_n33_55# 0.0116f
C3 a_n33_55# w_n124_n238# 0.0663f
C4 a_n88_n176# a_30_n176# 0.121f
C5 a_30_n176# w_n124_n238# 0.00827f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt M4 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n33_55# a_30_n176# 0.0116f
C1 a_n88_n176# w_n124_n238# 0.00827f
C2 a_n88_n176# a_n33_55# 0.0116f
C3 a_n33_55# w_n124_n238# 0.0663f
C4 a_n88_n176# a_30_n176# 0.121f
C5 a_30_n176# w_n124_n238# 0.00827f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt Ml2 a_n33_51# a_30_n171# a_n88_n171# VSUBS
X0 a_30_n171# a_n33_51# a_n88_n171# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_30_n171# a_n33_51# 0.0116f
C1 a_30_n171# a_n88_n171# 0.121f
C2 a_n88_n171# a_n33_51# 0.0116f
C3 a_30_n171# VSUBS 0.121f
C4 a_n88_n171# VSUBS 0.121f
C5 a_n33_51# VSUBS 0.227f
.ends

.subckt M2 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n33_55# a_30_n176# 0.0116f
C1 a_n88_n176# w_n124_n238# 0.00827f
C2 a_n88_n176# a_n33_55# 0.0116f
C3 a_n33_55# w_n124_n238# 0.0663f
C4 a_n88_n176# a_30_n176# 0.121f
C5 a_30_n176# w_n124_n238# 0.00827f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt Ml3 a_n88_n176# a_n33_55# w_n124_n238# a_30_n176# VSUBS
X0 a_30_n176# a_n33_55# a_n88_n176# w_n124_n238# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
C0 a_n33_55# a_30_n176# 0.0116f
C1 a_n88_n176# w_n124_n238# 0.00827f
C2 a_n88_n176# a_n33_55# 0.0116f
C3 a_n33_55# w_n124_n238# 0.0663f
C4 a_n88_n176# a_30_n176# 0.121f
C5 a_30_n176# w_n124_n238# 0.00827f
C6 a_30_n176# VSUBS 0.113f
C7 a_n88_n176# VSUBS 0.113f
C8 a_n33_55# VSUBS 0.167f
C9 w_n124_n238# VSUBS 0.269f
.ends

.subckt comparator_core outn clk ip in diff outp w_302_2337# vdd vn vp vss
XMdiff_0 clk vss diff vss Mdiff
XMdiff_1 clk diff vss vss Mdiff
XM3_0 outp clk w_302_2337# vdd vss M3
XMl1_0 outp outn in vss Ml1
XMinp_0 vp ip diff vss Minp
XM1_0 in clk w_302_2337# vdd vss M1
XMinn_0 vn diff in vss Minn
XMl4_0 vdd outn w_302_2337# outp vss Ml4
XM4_0 vdd clk w_302_2337# ip vss M4
XMl2_0 outn ip outp vss Ml2
XM2_0 vdd clk w_302_2337# outn vss M2
XMl3_0 outn outp w_302_2337# vdd vss Ml3
C0 vdd vn 0.0761f
C1 in vdd 0.111f
C2 vdd vp 0.0755f
C3 outp diff 0.00669f
C4 outp outn 1.02f
C5 ip diff 0.0808f
C6 outp vn 0.223f
C7 ip outn 0.0133f
C8 outp in 0.0133f
C9 outp vp 0.236f
C10 outn w_302_2337# 0.304f
C11 diff clk 0.0314f
C12 outn clk 0.215f
C13 w_302_2337# vn 0.0775f
C14 ip vp 0.0723f
C15 clk vn 0.0937f
C16 outp vdd 0.204f
C17 w_302_2337# in 0.0589f
C18 w_302_2337# vp 0.0765f
C19 ip vdd 0.11f
C20 in clk 0.436f
C21 clk vp 0.0951f
C22 w_302_2337# vdd 1.17f
C23 clk vdd 0.276f
C24 outn diff 0.00221f
C25 outp ip 0.0618f
C26 diff vn 0.00126f
C27 outn vn 0.167f
C28 outp w_302_2337# 0.291f
C29 outp clk 0.21f
C30 in diff 0.0808f
C31 diff vp 0.00126f
C32 outn in 0.0617f
C33 ip w_302_2337# 0.0584f
C34 outn vp 0.178f
C35 ip clk 0.436f
C36 in vn 0.0722f
C37 vp vn 0.202f
C38 outn vdd 0.211f
C39 w_302_2337# clk 0.222f
C40 clk vss 3.13f
C41 vdd vss 2.09f
C42 outn vss 1.77f
C43 w_302_2337# vss 4.58f
C44 vn vss 1.7f
C45 ip vss 1.16f
C46 vp vss 1.69f
C47 in vss 1.16f
C48 outp vss 1.76f
C49 diff vss 0.226f
.ends

.subckt comparator trim_3 trim_2 trim_0 trim_1 trim_4 trimb_4 trimb_1 trimb_0 trimb_2
+ trimb_3 outn outp clk vdd vss vn vp
Xtrim_0 trim_0/n1 trim_0/n0 trim_4 trim_3 trim_2 trim_1 trim_0 trim_0/n2 trim_0/n4
+ vss trim_0/drain trim_0/n3 trim
Xtrim_1 trim_1/n1 trim_1/n0 trimb_4 trimb_3 trimb_2 trimb_1 trimb_0 trim_1/n2 trim_1/n4
+ vss trim_1/drain trim_1/n3 trim
Xcomparator_core_0 outn clk trim_1/drain trim_0/drain comparator_core_0/diff outp
+ comparator_core_0/w_302_2337# vdd vn vp vss comparator_core
X0 trim_0/n4 trim_4.t7 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X1 trim_0/n3 trim_3.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X2 vss trimb_3.t3 trim_1/n3 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X3 trim_1/n3 trimb_3.t2 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X4 trim_0/n4 trim_4.t4 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X5 trim_1/n4 trimb_4.t4 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X6 trim_0/n4 trim_4.t1 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X7 vss trim_3.t1 trim_0/n3 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X8 trim_1/n4 trimb_4.t1 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X9 vss trimb_3.t1 trim_1/n3 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X10 trim_0/n2 trim_2.t1 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X11 trim_1/drain vp.t0 comparator_core_0/diff vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X12 comparator_core_0/diff vn.t0 trim_0/drain vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X13 vss trim_4.t6 trim_0/n4 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X14 trim_1/n2 trimb_2.t1 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X15 vss trimb_4.t6 trim_1/n4 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X16 vss trimb_4.t5 trim_1/n4 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X17 comparator_core_0/diff clk.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X18 trim_1/drain clk.t4 vdd comparator_core_0/w_302_2337# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X19 vss trim_4.t5 trim_0/n4 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X20 outp outn.t0 vdd comparator_core_0/w_302_2337# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X21 vdd outp.t1 outn comparator_core_0/w_302_2337# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X22 outn clk.t5 vdd comparator_core_0/w_302_2337# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X23 trim_0/n3 trim_3.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X24 outn outp.t0 trim_0/drain vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X25 trim_1/n3 trimb_3.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X26 trim_0/n1 trim_1.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X27 vss trim_2.t0 trim_0/n2 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X28 trim_1/n1 trimb_1.t0 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X29 trim_1/drain outn.t1 outp vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X30 trim_0/n4 trim_4.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X31 vss trimb_2.t0 trim_1/n2 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X32 trim_1/n4 trimb_4.t3 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X33 vdd clk.t2 outp comparator_core_0/w_302_2337# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X34 vss trim_4.t2 trim_0/n4 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X35 vss trimb_4.t2 trim_1/n4 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X36 vdd clk.t3 trim_0/drain comparator_core_0/w_302_2337# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X37 vss trimb_4.t0 trim_1/n4 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X38 vss clk.t0 comparator_core_0/diff vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X39 vss trim_4.t0 trim_0/n4 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X40 trim_1/n4 trimb_4.t7 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X41 vss trim_0.t0 trim_0/n0 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X42 vss trim_3.t3 trim_0/n3 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X43 vss trimb_0.t0 trim_1/n0 vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
R0 trim_2.n0 trim_2.t0 135.6
R1 trim_2.n0 trim_2.t1 135.6
R2 trim_2 trim_2 5.838
R3 trim_2 trim_2.n0 2.56687
R4 vss.n168 vss.n119 2916.35
R5 vss.n483 vss.n482 1084.91
R6 vss.n220 vss.n171 833.399
R7 vss.n109 vss.n108 292.5
R8 vss.n107 vss.n106 292.5
R9 vss.n105 vss.n104 292.5
R10 vss.n103 vss.n102 292.5
R11 vss.n101 vss.n100 292.5
R12 vss.n99 vss.n98 292.5
R13 vss.n97 vss.n96 292.5
R14 vss.n95 vss.n94 292.5
R15 vss.n93 vss.n92 292.5
R16 vss.n91 vss.n90 292.5
R17 vss.n89 vss.n88 292.5
R18 vss.n88 vss.n87 292.5
R19 vss.n86 vss.n85 292.5
R20 vss.n85 vss.n84 292.5
R21 vss.n83 vss.n82 292.5
R22 vss.n82 vss.n81 292.5
R23 vss.n80 vss.n79 292.5
R24 vss.n79 vss.n78 292.5
R25 vss.n77 vss.n76 292.5
R26 vss.n76 vss.n75 292.5
R27 vss.n74 vss.n73 292.5
R28 vss.n73 vss.n72 292.5
R29 vss.n71 vss.n70 292.5
R30 vss.n70 vss.n69 292.5
R31 vss.n68 vss.n67 292.5
R32 vss.n67 vss.n66 292.5
R33 vss.n511 vss.n510 292.5
R34 vss.n510 vss.n509 292.5
R35 vss.n514 vss.n513 292.5
R36 vss.n513 vss.n512 292.5
R37 vss.n517 vss.n516 292.5
R38 vss.n516 vss.n515 292.5
R39 vss.n520 vss.n519 292.5
R40 vss.n519 vss.n518 292.5
R41 vss.n523 vss.n522 292.5
R42 vss.n522 vss.n521 292.5
R43 vss.n526 vss.n525 292.5
R44 vss.n525 vss.n524 292.5
R45 vss.n529 vss.n528 292.5
R46 vss.n528 vss.n527 292.5
R47 vss.n531 vss.n530 292.5
R48 vss.n533 vss.n532 292.5
R49 vss.n535 vss.n534 292.5
R50 vss.n537 vss.n536 292.5
R51 vss.n539 vss.n538 292.5
R52 vss.n541 vss.n540 292.5
R53 vss.n543 vss.n542 292.5
R54 vss.n545 vss.n544 292.5
R55 vss.n547 vss.n546 292.5
R56 vss.n549 vss.n548 292.5
R57 vss.n379 vss.n378 292.5
R58 vss.n377 vss.n376 292.5
R59 vss.n375 vss.n374 292.5
R60 vss.n373 vss.n372 292.5
R61 vss.n371 vss.n370 292.5
R62 vss.n369 vss.n368 292.5
R63 vss.n367 vss.n366 292.5
R64 vss.n365 vss.n364 292.5
R65 vss.n363 vss.n362 292.5
R66 vss.n361 vss.n360 292.5
R67 vss.n359 vss.n358 292.5
R68 vss.n357 vss.n356 292.5
R69 vss.n355 vss.n354 292.5
R70 vss.n353 vss.n352 292.5
R71 vss.n351 vss.n350 292.5
R72 vss.n349 vss.n348 292.5
R73 vss.n347 vss.n346 292.5
R74 vss.n1 vss.n0 292.5
R75 vss.n3 vss.n2 292.5
R76 vss.n5 vss.n4 292.5
R77 vss.n7 vss.n6 292.5
R78 vss.n9 vss.n8 292.5
R79 vss.n11 vss.n10 292.5
R80 vss.n13 vss.n12 292.5
R81 vss.n15 vss.n14 292.5
R82 vss.n17 vss.n16 292.5
R83 vss.n19 vss.n18 292.5
R84 vss.n21 vss.n20 292.5
R85 vss.n23 vss.n22 292.5
R86 vss.n25 vss.n24 292.5
R87 vss.n27 vss.n26 292.5
R88 vss.n29 vss.n28 292.5
R89 vss.n31 vss.n30 292.5
R90 vss.n33 vss.n32 292.5
R91 vss.n472 vss.n471 292.5
R92 vss.n470 vss.n469 292.5
R93 vss.n428 vss.n427 292.5
R94 vss.n406 vss.n405 292.5
R95 vss.n399 vss.n398 292.5
R96 vss.n401 vss.n400 292.5
R97 vss.n419 vss.n418 292.5
R98 vss.n417 vss.n416 292.5
R99 vss.n438 vss.n437 292.5
R100 vss.n453 vss.n452 292.5
R101 vss.n391 vss.n390 292.5
R102 vss.n393 vss.n392 292.5
R103 vss.n463 vss.n462 292.5
R104 vss.n461 vss.n460 292.5
R105 vss.n459 vss.n458 292.5
R106 vss.n432 vss.n431 292.5
R107 vss.n434 vss.n433 292.5
R108 vss.n436 vss.n435 292.5
R109 vss.n335 vss.n334 292.5
R110 vss.n333 vss.n332 292.5
R111 vss.n331 vss.n330 292.5
R112 vss.n263 vss.n262 292.5
R113 vss.n243 vss.n242 292.5
R114 vss.n300 vss.n299 292.5
R115 vss.n302 vss.n301 292.5
R116 vss.n304 vss.n303 292.5
R117 vss.n306 vss.n305 292.5
R118 vss.n169 vss.n168 233.006
R119 vss.n494 vss.n493 222.222
R120 vss.n221 vss.n220 216.75
R121 vss.n54 vss.n53 204.445
R122 vss.n34 vss.n33 163.766
R123 vss.n243 vss.n241 163.766
R124 vss.n424 vss.n419 162.964
R125 vss.n496 vss.n495 157.778
R126 vss.n56 vss.n55 157.778
R127 vss.n407 vss.n406 155.482
R128 vss.n478 vss.n393 153.91
R129 vss.n402 vss.n401 150.213
R130 vss.n482 vss.n478 147.875
R131 vss.n424 vss.n423 147.875
R132 vss.n441 vss.n440 146.447
R133 vss.n456 vss.n455 144.189
R134 vss.n380 vss.n379 144.189
R135 vss.n306 vss.n304 144.189
R136 vss.n429 vss.n428 140.968
R137 vss.n473 vss.n472 135.697
R138 vss.n550 vss.n549 131.766
R139 vss.n336 vss.n335 131.766
R140 vss.n110 vss.n109 125.742
R141 vss.n264 vss.n263 125.742
R142 vss.n422 vss.n420 117.719
R143 vss.n481 vss.n479 117.719
R144 vss.n219 vss.n218 117.719
R145 vss.n219 vss.n217 117.719
R146 vss.n422 vss.n421 117.719
R147 vss.n481 vss.n480 117.719
R148 vss.n216 vss.n214 117.719
R149 vss.n213 vss.n211 117.719
R150 vss.n210 vss.n208 117.719
R151 vss.n207 vss.n205 117.719
R152 vss.n204 vss.n202 117.719
R153 vss.n201 vss.n199 117.719
R154 vss.n198 vss.n196 117.719
R155 vss.n195 vss.n193 117.719
R156 vss.n192 vss.n190 117.719
R157 vss.n189 vss.n187 117.719
R158 vss.n186 vss.n184 117.719
R159 vss.n183 vss.n181 117.719
R160 vss.n180 vss.n178 117.719
R161 vss.n177 vss.n175 117.719
R162 vss.n124 vss.n122 117.719
R163 vss.n127 vss.n125 117.719
R164 vss.n130 vss.n128 117.719
R165 vss.n133 vss.n131 117.719
R166 vss.n136 vss.n134 117.719
R167 vss.n139 vss.n137 117.719
R168 vss.n142 vss.n140 117.719
R169 vss.n145 vss.n143 117.719
R170 vss.n148 vss.n146 117.719
R171 vss.n151 vss.n149 117.719
R172 vss.n154 vss.n152 117.719
R173 vss.n157 vss.n155 117.719
R174 vss.n160 vss.n158 117.719
R175 vss.n163 vss.n161 117.719
R176 vss.n166 vss.n164 117.719
R177 vss.n166 vss.n165 117.719
R178 vss.n163 vss.n162 117.719
R179 vss.n160 vss.n159 117.719
R180 vss.n157 vss.n156 117.719
R181 vss.n154 vss.n153 117.719
R182 vss.n151 vss.n150 117.719
R183 vss.n148 vss.n147 117.719
R184 vss.n145 vss.n144 117.719
R185 vss.n142 vss.n141 117.719
R186 vss.n139 vss.n138 117.719
R187 vss.n136 vss.n135 117.719
R188 vss.n133 vss.n132 117.719
R189 vss.n130 vss.n129 117.719
R190 vss.n127 vss.n126 117.719
R191 vss.n124 vss.n123 117.719
R192 vss.n121 vss.n120 117.719
R193 vss.n216 vss.n215 117.719
R194 vss.n213 vss.n212 117.719
R195 vss.n210 vss.n209 117.719
R196 vss.n207 vss.n206 117.719
R197 vss.n204 vss.n203 117.719
R198 vss.n201 vss.n200 117.719
R199 vss.n198 vss.n197 117.719
R200 vss.n195 vss.n194 117.719
R201 vss.n192 vss.n191 117.719
R202 vss.n189 vss.n188 117.719
R203 vss.n186 vss.n185 117.719
R204 vss.n183 vss.n182 117.719
R205 vss.n180 vss.n179 117.719
R206 vss.n177 vss.n176 117.719
R207 vss.n174 vss.n173 117.719
R208 vss.n393 vss.n391 102.606
R209 vss.n419 vss.n417 102.606
R210 vss.n464 vss.n457 100.216
R211 vss.n443 vss.n442 100.216
R212 vss.n220 vss.n219 87.3927
R213 vss.n423 vss.n422 87.3927
R214 vss.n482 vss.n481 87.3927
R215 vss.n168 vss.n167 87.3925
R216 vss.n168 vss.n166 87.3925
R217 vss.n168 vss.n163 87.3925
R218 vss.n168 vss.n160 87.3925
R219 vss.n168 vss.n157 87.3925
R220 vss.n168 vss.n154 87.3925
R221 vss.n168 vss.n151 87.3925
R222 vss.n168 vss.n148 87.3925
R223 vss.n168 vss.n145 87.3925
R224 vss.n168 vss.n142 87.3925
R225 vss.n168 vss.n139 87.3925
R226 vss.n168 vss.n136 87.3925
R227 vss.n168 vss.n133 87.3925
R228 vss.n168 vss.n130 87.3925
R229 vss.n168 vss.n127 87.3925
R230 vss.n168 vss.n124 87.3925
R231 vss.n168 vss.n121 87.3925
R232 vss.n220 vss.n216 87.3925
R233 vss.n220 vss.n213 87.3925
R234 vss.n220 vss.n210 87.3925
R235 vss.n220 vss.n207 87.3925
R236 vss.n220 vss.n204 87.3925
R237 vss.n220 vss.n201 87.3925
R238 vss.n220 vss.n198 87.3925
R239 vss.n220 vss.n195 87.3925
R240 vss.n220 vss.n192 87.3925
R241 vss.n220 vss.n189 87.3925
R242 vss.n220 vss.n186 87.3925
R243 vss.n220 vss.n183 87.3925
R244 vss.n220 vss.n180 87.3925
R245 vss.n220 vss.n177 87.3925
R246 vss.n220 vss.n174 87.3925
R247 vss.n220 vss.n172 87.3925
R248 vss.n53 vss.n52 75.5561
R249 vss.n52 vss.n51 75.5561
R250 vss.n51 vss.n50 75.5561
R251 vss.n50 vss.n49 75.5561
R252 vss.n49 vss.n48 75.5561
R253 vss.n48 vss.n47 75.5561
R254 vss.n47 vss.n46 75.5561
R255 vss.n46 vss.n45 75.5561
R256 vss.n45 vss.n44 75.5561
R257 vss.n485 vss.n484 75.5561
R258 vss.n486 vss.n485 75.5561
R259 vss.n487 vss.n486 75.5561
R260 vss.n488 vss.n487 75.5561
R261 vss.n489 vss.n488 75.5561
R262 vss.n490 vss.n489 75.5561
R263 vss.n491 vss.n490 75.5561
R264 vss.n492 vss.n491 75.5561
R265 vss.n493 vss.n492 75.5561
R266 vss.n280 vss.n221 65.0251
R267 vss.n425 vss.n413 63.7358
R268 vss.n477 vss.n396 63.7358
R269 vss.n389 vss.n388 57.3393
R270 vss.n417 vss.n415 57.3393
R271 vss.n223 vss.n222 52.1476
R272 vss.n118 vss.n117 52.1476
R273 vss.n279 vss.n223 46.3534
R274 vss.n281 vss.n118 46.3534
R275 vss.n391 vss.n389 45.268
R276 vss.n388 vss.n387 45.268
R277 vss.n415 vss.n414 45.268
R278 vss.n500 vss.n499 40.5593
R279 vss.n57 vss.n43 40.5593
R280 vss.n443 vss.n436 30.5684
R281 vss.n464 vss.n463 28.3093
R282 vss.n498 vss.n497 27.6046
R283 vss.n42 vss.n41 27.6046
R284 vss.n499 vss.n498 27.6046
R285 vss.n43 vss.n42 27.6046
R286 vss.n457 vss.n456 25.6005
R287 vss.n455 vss.n454 25.6005
R288 vss.n454 vss.n453 25.6005
R289 vss.n439 vss.n438 25.6005
R290 vss.n440 vss.n439 25.6005
R291 vss.n442 vss.n441 25.6005
R292 vss.n463 vss.n461 25.6005
R293 vss.n461 vss.n459 25.6005
R294 vss.n434 vss.n432 25.6005
R295 vss.n436 vss.n434 25.6005
R296 vss.n472 vss.n470 25.6005
R297 vss.n401 vss.n399 25.6005
R298 vss.n109 vss.n107 25.6005
R299 vss.n107 vss.n105 25.6005
R300 vss.n105 vss.n103 25.6005
R301 vss.n103 vss.n101 25.6005
R302 vss.n101 vss.n99 25.6005
R303 vss.n99 vss.n97 25.6005
R304 vss.n97 vss.n95 25.6005
R305 vss.n95 vss.n93 25.6005
R306 vss.n93 vss.n91 25.6005
R307 vss.n91 vss.n89 25.6005
R308 vss.n89 vss.n86 25.6005
R309 vss.n86 vss.n83 25.6005
R310 vss.n83 vss.n80 25.6005
R311 vss.n80 vss.n77 25.6005
R312 vss.n77 vss.n74 25.6005
R313 vss.n74 vss.n71 25.6005
R314 vss.n71 vss.n68 25.6005
R315 vss.n514 vss.n511 25.6005
R316 vss.n517 vss.n514 25.6005
R317 vss.n520 vss.n517 25.6005
R318 vss.n523 vss.n520 25.6005
R319 vss.n526 vss.n523 25.6005
R320 vss.n529 vss.n526 25.6005
R321 vss.n531 vss.n529 25.6005
R322 vss.n533 vss.n531 25.6005
R323 vss.n535 vss.n533 25.6005
R324 vss.n537 vss.n535 25.6005
R325 vss.n539 vss.n537 25.6005
R326 vss.n541 vss.n539 25.6005
R327 vss.n543 vss.n541 25.6005
R328 vss.n545 vss.n543 25.6005
R329 vss.n547 vss.n545 25.6005
R330 vss.n549 vss.n547 25.6005
R331 vss.n33 vss.n31 25.6005
R332 vss.n31 vss.n29 25.6005
R333 vss.n29 vss.n27 25.6005
R334 vss.n27 vss.n25 25.6005
R335 vss.n25 vss.n23 25.6005
R336 vss.n23 vss.n21 25.6005
R337 vss.n21 vss.n19 25.6005
R338 vss.n19 vss.n17 25.6005
R339 vss.n17 vss.n15 25.6005
R340 vss.n15 vss.n13 25.6005
R341 vss.n13 vss.n11 25.6005
R342 vss.n11 vss.n9 25.6005
R343 vss.n9 vss.n7 25.6005
R344 vss.n7 vss.n5 25.6005
R345 vss.n5 vss.n3 25.6005
R346 vss.n3 vss.n1 25.6005
R347 vss.n349 vss.n347 25.6005
R348 vss.n351 vss.n349 25.6005
R349 vss.n353 vss.n351 25.6005
R350 vss.n355 vss.n353 25.6005
R351 vss.n357 vss.n355 25.6005
R352 vss.n359 vss.n357 25.6005
R353 vss.n361 vss.n359 25.6005
R354 vss.n363 vss.n361 25.6005
R355 vss.n365 vss.n363 25.6005
R356 vss.n367 vss.n365 25.6005
R357 vss.n369 vss.n367 25.6005
R358 vss.n371 vss.n369 25.6005
R359 vss.n373 vss.n371 25.6005
R360 vss.n375 vss.n373 25.6005
R361 vss.n377 vss.n375 25.6005
R362 vss.n379 vss.n377 25.6005
R363 vss.n263 vss.n261 25.6005
R364 vss.n261 vss.n260 25.6005
R365 vss.n260 vss.n259 25.6005
R366 vss.n259 vss.n258 25.6005
R367 vss.n258 vss.n257 25.6005
R368 vss.n257 vss.n256 25.6005
R369 vss.n256 vss.n255 25.6005
R370 vss.n255 vss.n254 25.6005
R371 vss.n254 vss.n253 25.6005
R372 vss.n253 vss.n252 25.6005
R373 vss.n252 vss.n251 25.6005
R374 vss.n251 vss.n250 25.6005
R375 vss.n250 vss.n249 25.6005
R376 vss.n249 vss.n248 25.6005
R377 vss.n248 vss.n247 25.6005
R378 vss.n247 vss.n246 25.6005
R379 vss.n316 vss.n315 25.6005
R380 vss.n317 vss.n316 25.6005
R381 vss.n318 vss.n317 25.6005
R382 vss.n319 vss.n318 25.6005
R383 vss.n320 vss.n319 25.6005
R384 vss.n321 vss.n320 25.6005
R385 vss.n322 vss.n321 25.6005
R386 vss.n323 vss.n322 25.6005
R387 vss.n324 vss.n323 25.6005
R388 vss.n325 vss.n324 25.6005
R389 vss.n326 vss.n325 25.6005
R390 vss.n327 vss.n326 25.6005
R391 vss.n328 vss.n327 25.6005
R392 vss.n329 vss.n328 25.6005
R393 vss.n331 vss.n329 25.6005
R394 vss.n333 vss.n331 25.6005
R395 vss.n335 vss.n333 25.6005
R396 vss.n241 vss.n240 25.6005
R397 vss.n240 vss.n239 25.6005
R398 vss.n239 vss.n238 25.6005
R399 vss.n238 vss.n237 25.6005
R400 vss.n237 vss.n236 25.6005
R401 vss.n236 vss.n235 25.6005
R402 vss.n235 vss.n234 25.6005
R403 vss.n234 vss.n233 25.6005
R404 vss.n233 vss.n232 25.6005
R405 vss.n232 vss.n231 25.6005
R406 vss.n231 vss.n230 25.6005
R407 vss.n230 vss.n229 25.6005
R408 vss.n229 vss.n228 25.6005
R409 vss.n228 vss.n227 25.6005
R410 vss.n227 vss.n226 25.6005
R411 vss.n285 vss.n284 25.6005
R412 vss.n286 vss.n285 25.6005
R413 vss.n287 vss.n286 25.6005
R414 vss.n288 vss.n287 25.6005
R415 vss.n289 vss.n288 25.6005
R416 vss.n290 vss.n289 25.6005
R417 vss.n291 vss.n290 25.6005
R418 vss.n292 vss.n291 25.6005
R419 vss.n293 vss.n292 25.6005
R420 vss.n294 vss.n293 25.6005
R421 vss.n295 vss.n294 25.6005
R422 vss.n296 vss.n295 25.6005
R423 vss.n297 vss.n296 25.6005
R424 vss.n298 vss.n297 25.6005
R425 vss.n300 vss.n298 25.6005
R426 vss.n302 vss.n300 25.6005
R427 vss.n304 vss.n302 25.6005
R428 vss.n412 vss.n411 16.8818
R429 vss.n395 vss.n394 16.8818
R430 vss.n413 vss.n412 16.8818
R431 vss.n396 vss.n395 16.8818
R432 vss.n381 vss.n380 16.5652
R433 vss.n35 vss.n34 16.5652
R434 vss.n244 vss.n243 16.1887
R435 vss.n307 vss.n306 16.1887
R436 vss.n484 vss.n483 13.3338
R437 vss.n170 vss.n169 9.75419
R438 vss.n308 vss.n307 9.31144
R439 vss.n36 vss.n35 9.31039
R440 vss.n382 vss.n381 9.31039
R441 vss.n502 vss.n501 9.3005
R442 vss.n501 vss.n500 9.3005
R443 vss.n59 vss.n58 9.3005
R444 vss.n58 vss.n57 9.3005
R445 vss.n426 vss.n425 9.3005
R446 vss.n425 vss.n424 9.3005
R447 vss.n477 vss.n476 9.3005
R448 vss.n478 vss.n477 9.3005
R449 vss.n278 vss.n277 9.3005
R450 vss.n279 vss.n278 9.3005
R451 vss.n280 vss.n279 9.3005
R452 vss.n283 vss.n282 9.3005
R453 vss.n282 vss.n281 9.3005
R454 vss.n281 vss.n280 9.3005
R455 vss.n384 vss.n383 9.0005
R456 vss.n38 vss.n37 9.0005
R457 vss.n310 vss.n309 9.0005
R458 vss.n280 vss.n170 8.67045
R459 vss.n500 vss.n496 5.01811
R460 vss.n57 vss.n56 5.01748
R461 vss.n343 vss 4.80467
R462 vss.n556 vss.n555 4.74217
R463 vss.n430 vss.n407 4.57427
R464 vss.n468 vss.n402 4.57427
R465 vss.n551 vss.n550 4.57427
R466 vss.n111 vss.n110 4.57427
R467 vss.n265 vss.n264 4.57427
R468 vss.n337 vss.n336 4.57427
R469 vss.n496 vss.n494 4.15288
R470 vss.n56 vss.n54 4.15252
R471 vss.n426 vss.n410 4.14168
R472 vss.n476 vss.n475 4.14168
R473 vss.n555 vss.n345 4.02849
R474 vss.n386 vss.n385 3.76521
R475 vss.n40 vss.n39 3.76521
R476 vss.n245 vss.n244 3.76521
R477 vss.n225 vss.n224 3.38874
R478 vss.n116 vss.n115 3.38874
R479 vss.n278 vss.n225 3.01226
R480 vss.n282 vss.n116 3.01226
R481 vss.n276 vss.n275 3.0005
R482 vss.n61 vss.n60 3.0005
R483 vss.n113 vss.n112 3.0005
R484 vss.n504 vss.n503 3.0005
R485 vss.n553 vss.n552 3.0005
R486 vss.n312 vss.n311 3.0005
R487 vss.n341 vss.n340 3.0005
R488 vss.n429 vss.n426 2.65111
R489 vss.n476 vss.n473 2.65111
R490 vss.n501 vss.n386 2.63579
R491 vss.n58 vss.n40 2.63579
R492 vss.n278 vss.n245 2.63579
R493 vss.n410 vss.n409 2.25932
R494 vss.n475 vss.n474 2.25932
R495 vss.n345 vss.n344 2.21752
R496 vss.n430 vss.n429 2.05223
R497 vss.n473 vss.n468 2.05223
R498 vss.n465 vss.n464 1.84239
R499 vss.n444 vss.n443 1.84237
R500 vss.n344 vss.n343 1.81065
R501 vss.n468 vss.n467 1.77862
R502 vss.n446 vss.n430 1.4761
R503 vss vss.n345 1.47472
R504 vss.n344 vss 0.752104
R505 vss.n450 vss.n449 0.673937
R506 vss.n449 vss.n448 0.673937
R507 vss.n449 vss 0.41925
R508 vss.n343 vss.n342 0.359081
R509 vss.n556 vss.n114 0.358301
R510 vss.n555 vss.n554 0.358301
R511 vss.n271 vss 0.296581
R512 vss.n467 vss.n466 0.0697748
R513 vss vss.n556 0.063
R514 vss.n446 vss.n445 0.0589808
R515 vss.n447 vss.n446 0.0581328
R516 vss.n268 vss.n267 0.0525833
R517 vss.n65 vss.n64 0.0525833
R518 vss.n508 vss.n507 0.0525833
R519 vss.n339 vss.n338 0.0525833
R520 vss.n467 vss.n451 0.0467812
R521 vss.n267 vss.n266 0.0421667
R522 vss.n340 vss.n339 0.0421667
R523 vss.n112 vss.n65 0.0400833
R524 vss.n552 vss.n508 0.0400833
R525 vss.n274 vss.n273 0.0395625
R526 vss.n63 vss.n62 0.0395625
R527 vss.n506 vss.n505 0.0395625
R528 vss.n314 vss.n313 0.0395625
R529 vss.n277 vss.n268 0.0338333
R530 vss.n273 vss.n272 0.03175
R531 vss.n451 vss.n450 0.03175
R532 vss.n448 vss.n447 0.03175
R533 vss.n62 vss.n61 0.03175
R534 vss.n505 vss.n504 0.03175
R535 vss.n341 vss.n314 0.03175
R536 vss.n275 vss.n274 0.0301875
R537 vss.n466 vss.n465 0.0301875
R538 vss.n445 vss.n444 0.0301875
R539 vss.n113 vss.n63 0.0301875
R540 vss.n553 vss.n506 0.0301875
R541 vss.n313 vss.n312 0.0301875
R542 vss.n114 vss.n113 0.022812
R543 vss.n554 vss.n553 0.022812
R544 vss.n272 vss.n271 0.0220368
R545 vss.n342 vss.n341 0.0220368
R546 vss.n468 vss.n403 0.0201429
R547 vss.n430 vss.n408 0.0201429
R548 vss.n430 vss.n404 0.01925
R549 vss.n270 vss.n269 0.0113746
R550 vss.n310 vss.n308 0.0113746
R551 vss.n468 vss.n397 0.0103652
R552 vss.n38 vss.n36 0.0103391
R553 vss.n384 vss.n382 0.0103391
R554 vss.n266 vss.n265 0.00883333
R555 vss.n276 vss.n270 0.00883333
R556 vss.n60 vss.n38 0.00883333
R557 vss.n60 vss.n59 0.00883333
R558 vss.n112 vss.n111 0.00883333
R559 vss.n503 vss.n384 0.00883333
R560 vss.n503 vss.n502 0.00883333
R561 vss.n552 vss.n551 0.00883333
R562 vss.n340 vss.n337 0.00883333
R563 vss.n311 vss.n310 0.00883333
R564 vss.n277 vss.n276 0.00675
R565 vss.n311 vss.n283 0.00675
R566 trim_0 trim_0.t0 138.256
R567 trim_0 trim_0 5.013
R568 trim_4.n0 trim_4.t1 135.841
R569 trim_4.n3 trim_4.t0 135.841
R570 trim_4.n3 trim_4.t7 135.52
R571 trim_4.n4 trim_4.t5 135.52
R572 trim_4.n5 trim_4.t4 135.52
R573 trim_4.n2 trim_4.t6 135.52
R574 trim_4.n1 trim_4.t3 135.52
R575 trim_4.n0 trim_4.t2 135.52
R576 trim_4 trim_4 2.57133
R577 trim_4 trim_4.n6 2.56687
R578 trim_4.n1 trim_4.n0 0.321152
R579 trim_4.n2 trim_4.n1 0.321152
R580 trim_4.n5 trim_4.n4 0.321152
R581 trim_4.n4 trim_4.n3 0.321152
R582 trim_4.n6 trim_4.n2 0.0793043
R583 trim_4.n6 trim_4.n5 0.0793043
R584 trim_1 trim_1.t0 138.256
R585 trim_1 trim_1 4.13383
R586 trim_3.n0 trim_3.t3 135.841
R587 trim_3.n1 trim_3.t2 135.841
R588 trim_3.n1 trim_3.t1 135.52
R589 trim_3.n0 trim_3.t0 135.52
R590 trim_3 trim_3 7.22342
R591 trim_3 trim_3.n2 2.56687
R592 trim_3.n2 trim_3.n0 0.0793043
R593 trim_3.n2 trim_3.n1 0.0793043
R594 trimb_2.n0 trimb_2.t0 135.6
R595 trimb_2.n0 trimb_2.t1 135.6
R596 trimb_2 trimb_2 5.92342
R597 trimb_2 trimb_2.n0 2.48064
R598 trimb_0 trimb_0.t0 138.169
R599 trimb_0 trimb_0 5.09842
R600 trimb_4.n0 trimb_4.t1 135.841
R601 trimb_4.n3 trimb_4.t0 135.841
R602 trimb_4.n3 trimb_4.t7 135.52
R603 trimb_4.n4 trimb_4.t5 135.52
R604 trimb_4.n5 trimb_4.t4 135.52
R605 trimb_4.n2 trimb_4.t6 135.52
R606 trimb_4.n1 trimb_4.t3 135.52
R607 trimb_4.n0 trimb_4.t2 135.52
R608 trimb_4 trimb_4 2.65675
R609 trimb_4 trimb_4.n6 2.48064
R610 trimb_4.n1 trimb_4.n0 0.321152
R611 trimb_4.n2 trimb_4.n1 0.321152
R612 trimb_4.n5 trimb_4.n4 0.321152
R613 trimb_4.n4 trimb_4.n3 0.321152
R614 trimb_4.n6 trimb_4.n2 0.0793043
R615 trimb_4.n6 trimb_4.n5 0.0793043
R616 trimb_1 trimb_1.t0 138.169
R617 trimb_1 trimb_1 4.21925
R618 trimb_3.n0 trimb_3.t3 135.841
R619 trimb_3.n1 trimb_3.t2 135.841
R620 trimb_3.n1 trimb_3.t1 135.52
R621 trimb_3.n0 trimb_3.t0 135.52
R622 trimb_3 trimb_3 7.30883
R623 trimb_3 trimb_3.n2 2.48064
R624 trimb_3.n2 trimb_3.n0 0.0793043
R625 trimb_3.n2 trimb_3.n1 0.0793043
R626 clk.n2 clk.t2 142.917
R627 clk.n0 clk.t5 142.911
R628 clk.n0 clk.t3 142.911
R629 clk.n2 clk.t4 142.905
R630 clk.n3 clk.t0 135.52
R631 clk.n1 clk.t1 135.52
R632 clk.n3 clk.n2 12.4888
R633 clk.n1 clk.n0 12.4715
R634 clk clk 4.14425
R635 clk clk.n4 0.84425
R636 clk.n4 clk.n1 0.0793043
R637 clk.n4 clk.n3 0.0793043
R638 outp.n0 outp.t1 146.688
R639 outp.n0 outp.t0 138.821
R640 outp outp.n0 9.64859
R641 outp outp 0.842688
R642 vdd.n9 vdd.n8 4.91552
R643 vdd.n11 vdd.n10 1.13717
R644 vdd vdd.n13 0.674808
R645 vdd.n13 vdd.n12 0.555146
R646 vdd.n3 vdd.n2 0.112557
R647 vdd.n7 vdd.n6 0.041625
R648 vdd.n1 vdd.n0 0.0364375
R649 vdd.n12 vdd.n11 0.0364375
R650 vdd.n8 vdd 0.024
R651 vdd.n5 vdd.n4 0.0140125
R652 vdd.n10 vdd.n9 0.0140125
R653 vdd.n2 vdd.n1 0.0083125
R654 vdd.n11 vdd.n3 0.0083125
R655 vdd.n6 vdd.n5 0.0034375
R656 vdd.n10 vdd.n7 0.0034375
R657 outn.n0 outn.t0 146.68
R658 outn.n0 outn.t1 138.822
R659 outn outn.n0 9.65222
R660 outn outn 0.842688
R661 vp.n1 vp.t0 138.87
R662 vp vp.n7 1.64973
R663 vp.n5 vp.n1 0.751481
R664 vp.n6 vp.n5 0.512485
R665 vp.n1 vp.n0 0.0589631
R666 vp.n5 vp.n4 0.0390429
R667 vp.n7 vp.n6 0.0146
R668 vp.n3 vp.n2 0.00458983
R669 vp.n4 vp.n3 0.0034375
R670 vn.n1 vn.t0 138.87
R671 vn vn.n7 1.64973
R672 vn.n5 vn.n1 0.750898
R673 vn.n6 vn.n5 0.513756
R674 vn.n1 vn.n0 0.0589632
R675 vn.n5 vn.n4 0.0392964
R676 vn.n7 vn.n6 0.0146
R677 vn.n3 vn.n2 0.00434178
R678 vn.n4 vn.n3 0.0034375
C0 vn trim_0/n0 9.27e-20
C1 trim_1/n1 vss 4.27e-20
C2 outn outp 0.00414f
C3 trim_2 trim_4 0.00265f
C4 vdd trim_0 0.0784f
C5 trim_1/n0 trim_1/n4 0.0442f
C6 trim_0/n2 trim_3 6.02e-19
C7 vdd trim_0/n3 0.0253f
C8 trim_1/drain outn 4.78e-20
C9 vdd trim_1 0.0649f
C10 trim_0/drain vn 0.0539f
C11 trim_0/n4 trim_0/n3 0.354f
C12 trim_0/n4 trim_1 0.00216f
C13 vdd trim_3 0.435f
C14 trimb_4 trimb_1 0.546f
C15 trim_0 vss 0.0573f
C16 vdd trimb_3 0.435f
C17 trim_0/n3 vss 2.61e-20
C18 trim_0/drain outp 4.78e-20
C19 vdd vp 0.221f
C20 vss trim_1 0.0863f
C21 trim_1/drain trim_1/n2 1.7f
C22 trim_3 vss 0.0691f
C23 trimb_3 vss 0.0691f
C24 trim_1/n1 trim_1/n4 0.0442f
C25 vp vss 0.00394f
C26 trim_0/n1 trim_0 2.97e-19
C27 trimb_3 trimb_2 1.07f
C28 trimb_0 trim_1/n2 3.92e-20
C29 comparator_core_0/w_302_2337# outp 5.68e-32
C30 trim_1/n3 trim_1/drain 3.41f
C31 trim_4 trim_0 0.0039f
C32 comparator_core_0/diff trim_1/drain -2.84e-32
C33 comparator_core_0/w_302_2337# trim_1/drain 0.00474f
C34 trimb_0 trimb_1 0.82f
C35 trim_4 trim_1 0.546f
C36 trim_4 trim_3 0.00191f
C37 trim_0 trim_0/n0 2.97e-19
C38 vdd clk 0.104f
C39 vp trim_1/n4 0.0126f
C40 vdd trim_0/n2 0.00772f
C41 trim_1/drain outp 0.0565f
C42 trim_0/n4 clk 2.01e-19
C43 trim_0/n4 trim_0/n2 0.177f
C44 trim_0/drain trim_0/n3 3.41f
C45 trim_1/n0 trim_1/drain 0.851f
C46 trimb_4 trimb_0 0.0039f
C47 vss clk 0.0684f
C48 trim_0/n2 vss 1.83e-20
C49 vdd trim_0/n4 0.0293f
C50 trimb_3 trim_1/n2 6.02e-19
C51 vp trim_1/n2 0.00276f
C52 vdd vss 5.14f
C53 trimb_0 trim_1/n0 2.97e-19
C54 trimb_3 trimb_1 3.33e-19
C55 trim_0/n4 vss 0.0914f
C56 vdd trimb_2 0.12f
C57 trim_1/n1 trim_1/drain 0.851f
C58 trimb_3 trim_1/n3 4.9e-19
C59 trim_1/n1 trim_1/n0 0.0442f
C60 vp trim_1/n3 0.00558f
C61 vn trim_0/n3 0.00558f
C62 trim_1/n4 clk 2.01e-19
C63 vdd trim_0/n1 0.00179f
C64 trimb_2 vss 0.0525f
C65 outn clk 0.0392f
C66 trim_0/n1 trim_0/n4 0.0442f
C67 vdd trim_4 0.103f
C68 trim_1/n1 trimb_0 2.97e-19
C69 trimb_4 trimb_3 0.00191f
C70 vdd trim_1/n4 0.0293f
C71 trim_0/n4 trim_4 0.00329f
C72 trim_2 trim_0 0.969f
C73 trim_0/n1 vss 4.27e-20
C74 vdd outn 0.102f
C75 trim_2 trim_1 4.8e-19
C76 vp outp 5.68e-32
C77 trim_4 vss 0.156f
C78 trim_0/drain clk 0.0801f
C79 trim_0/drain trim_0/n2 1.7f
C80 vdd trim_0/n0 0.00143f
C81 vp trim_1/drain 0.0539f
C82 trim_1/n4 vss 0.0914f
C83 trim_2 trim_3 1.07f
C84 vp trim_1/n0 9.27e-20
C85 trim_0/n4 trim_0/n0 0.0442f
C86 vss outn 0.12f
C87 trim_0/drain vdd 0.03f
C88 vdd trim_1/n2 0.00772f
C89 trimb_3 trimb_0 3.33e-19
C90 vdd trimb_1 0.0649f
C91 trim_0/drain trim_0/n4 6.86f
C92 trim_0/drain vss 1.71f
C93 vss trim_1/n2 1.83e-20
C94 vdd trim_1/n3 0.0253f
C95 vss trimb_1 0.0863f
C96 vdd comparator_core_0/diff 0.0019f
C97 vn clk 2.17e-19
C98 vdd comparator_core_0/w_302_2337# 0.346f
C99 trim_0/n2 vn 0.00276f
C100 trimb_2 trim_1/n2 7.08e-19
C101 trim_0/n1 trim_0/n0 0.0442f
C102 trim_0 trim_1 0.82f
C103 trim_1/n4 outn 3.12e-21
C104 trimb_2 trimb_1 4.8e-19
C105 outp clk 0.00182f
C106 trim_1/n3 vss 2.61e-20
C107 vdd trimb_4 0.103f
C108 trim_0 trim_3 3.33e-19
C109 vdd vn 0.221f
C110 trim_1/drain clk 0.0575f
C111 trim_0/drain trim_0/n1 0.851f
C112 trim_0/n3 trim_3 4.9e-19
C113 comparator_core_0/diff vss -5.68e-32
C114 comparator_core_0/w_302_2337# vss 6.22e-19
C115 trim_3 trim_1 3.33e-19
C116 trim_0/n4 vn 0.0126f
C117 trim_2 trim_0/n2 7.08e-19
C118 vdd outp 0.102f
C119 vdd trim_1/drain 0.0307f
C120 trim_1/n4 trim_1/n2 0.177f
C121 trimb_4 vss 0.156f
C122 vn vss 0.00394f
C123 trim_0/n4 outp 3.12e-21
C124 vdd trim_1/n0 0.00143f
C125 trim_1/n4 trimb_1 0.00216f
C126 trim_0/drain outn 0.0565f
C127 trim_2 vdd 0.12f
C128 trimb_4 trimb_2 0.00265f
C129 vss outp 0.12f
C130 trim_0/drain trim_0/n0 0.851f
C131 vss trim_1/drain 1.71f
C132 trim_1/n3 trim_1/n4 0.354f
C133 vdd trimb_0 0.0784f
C134 trim_2 vss 0.0525f
C135 comparator_core_0/w_302_2337# outn 5.68e-32
C136 trim_1/n2 trimb_1 4.74e-20
C137 trimb_0 vss 0.0573f
C138 vdd trim_1/n1 0.00179f
C139 trimb_4 trim_1/n4 0.00329f
C140 trim_0/n2 trim_0 3.92e-20
C141 vn outn 2.49e-32
C142 trimb_0 trimb_2 0.969f
C143 trim_0/n2 trim_1 4.74e-20
C144 trim_0/drain comparator_core_0/diff -2.84e-32
C145 trim_0/drain comparator_core_0/w_302_2337# 0.00484f
C146 trim_1/n4 trim_1/drain 6.86f
C147 vdd.n0 0 0.457f
C148 vdd.n1 0 0.00216f
C149 vdd.n2 0 0.0575f
C150 vdd.n3 0 0.0557f
C151 vdd.n4 0 1.43f
C152 vdd.n5 0 0.00216f
C153 vdd.n6 0 0.00578f
C154 vdd.n7 0 0.00578f
C155 vdd.n8 0 2.07f
C156 vdd.n9 0 0.649f
C157 vdd.n10 0 0.00216f
C158 vdd.n11 0 0.00216f
C159 vdd.n12 0 0.0293f
C160 vdd.n13 0 0.31f
C161 vss.n0 0 5.02e-19
C162 vss.n1 0 5.02e-19
C163 vss.n2 0 5.02e-19
C164 vss.n3 0 5.02e-19
C165 vss.n4 0 5.02e-19
C166 vss.n5 0 5.02e-19
C167 vss.n6 0 5.02e-19
C168 vss.n7 0 5.02e-19
C169 vss.n8 0 5.02e-19
C170 vss.n9 0 5.02e-19
C171 vss.n10 0 5.02e-19
C172 vss.n11 0 5.02e-19
C173 vss.n12 0 5.02e-19
C174 vss.n13 0 5.02e-19
C175 vss.n14 0 5.02e-19
C176 vss.n15 0 5.02e-19
C177 vss.n16 0 5.02e-19
C178 vss.n17 0 5.02e-19
C179 vss.n18 0 5.02e-19
C180 vss.n19 0 5.02e-19
C181 vss.n20 0 5.02e-19
C182 vss.n21 0 5.02e-19
C183 vss.n22 0 5.02e-19
C184 vss.n23 0 5.02e-19
C185 vss.n24 0 5.02e-19
C186 vss.n25 0 5.02e-19
C187 vss.n26 0 5.02e-19
C188 vss.n27 0 5.02e-19
C189 vss.n28 0 5.02e-19
C190 vss.n29 0 5.02e-19
C191 vss.n30 0 5.02e-19
C192 vss.n31 0 5.02e-19
C193 vss.n32 0 0.00191f
C194 vss.n33 0 0.00191f
C195 vss.n34 0 0.00183f
C196 vss.n35 0 1.96e-19
C197 vss.n36 0 3.84e-19
C198 vss.n37 0 6.27e-20
C199 vss.n38 0 8.46e-20
C200 vss.n39 0 2.1e-19
C201 vss.n40 0 6.27e-20
C202 vss.n41 0 0.0015f
C203 vss.n43 0 6.27e-20
C204 vss.n44 0 0.0584f
C205 vss.n45 0 0.0584f
C206 vss.n46 0 0.0584f
C207 vss.n47 0 0.0584f
C208 vss.n48 0 0.0584f
C209 vss.n49 0 0.0584f
C210 vss.n50 0 0.0584f
C211 vss.n51 0 0.0584f
C212 vss.n52 0 0.0584f
C213 vss.n53 0 0.108f
C214 vss.n54 0 0.8f
C215 vss.n55 0 0.0019f
C216 vss.n57 0 2.51e-19
C217 vss.n58 0 5.53e-20
C218 vss.n59 0 1.3e-19
C219 vss.n60 0 5.21e-20
C220 vss.n61 0 6.59e-19
C221 vss.n62 0 3.9e-19
C222 vss.n63 0 3.82e-19
C223 vss.n64 0 2.67e-19
C224 vss.n65 0 2.86e-19
C225 vss.n66 0 0.0584f
C226 vss.n67 0 5.02e-19
C227 vss.n68 0 5.02e-19
C228 vss.n69 0 0.0584f
C229 vss.n70 0 5.02e-19
C230 vss.n71 0 5.02e-19
C231 vss.n72 0 0.0584f
C232 vss.n73 0 5.02e-19
C233 vss.n74 0 5.02e-19
C234 vss.n75 0 0.0584f
C235 vss.n76 0 5.02e-19
C236 vss.n77 0 5.02e-19
C237 vss.n78 0 0.0584f
C238 vss.n79 0 5.02e-19
C239 vss.n80 0 5.02e-19
C240 vss.n81 0 0.0584f
C241 vss.n82 0 5.02e-19
C242 vss.n83 0 5.02e-19
C243 vss.n84 0 0.0584f
C244 vss.n85 0 5.02e-19
C245 vss.n86 0 5.02e-19
C246 vss.n87 0 0.0584f
C247 vss.n88 0 5.02e-19
C248 vss.n89 0 5.02e-19
C249 vss.n90 0 5.02e-19
C250 vss.n91 0 5.02e-19
C251 vss.n92 0 5.02e-19
C252 vss.n93 0 5.02e-19
C253 vss.n94 0 5.02e-19
C254 vss.n95 0 5.02e-19
C255 vss.n96 0 5.02e-19
C256 vss.n97 0 5.02e-19
C257 vss.n98 0 5.02e-19
C258 vss.n99 0 5.02e-19
C259 vss.n100 0 5.02e-19
C260 vss.n101 0 5.02e-19
C261 vss.n102 0 5.02e-19
C262 vss.n103 0 5.02e-19
C263 vss.n104 0 5.02e-19
C264 vss.n105 0 5.02e-19
C265 vss.n106 0 5.02e-19
C266 vss.n107 0 5.02e-19
C267 vss.n108 0 0.00173f
C268 vss.n109 0 0.00155f
C269 vss.n110 0 0.00147f
C270 vss.n111 0 4.67e-19
C271 vss.n112 0 1.5e-19
C272 vss.n113 0 3.5e-19
C273 vss.n114 0 0.00127f
C274 vss.n115 0 2.1e-19
C275 vss.n116 0 6.27e-20
C276 vss.n117 0 0.00156f
C277 vss.n118 0 6.27e-20
C278 vss.n119 0 1.53f
C279 vss.n120 0 5.02e-19
C280 vss.n122 0 5.02e-19
C281 vss.n123 0 5.02e-19
C282 vss.n125 0 5.02e-19
C283 vss.n126 0 5.02e-19
C284 vss.n128 0 5.02e-19
C285 vss.n129 0 5.02e-19
C286 vss.n131 0 5.02e-19
C287 vss.n132 0 5.02e-19
C288 vss.n134 0 5.02e-19
C289 vss.n135 0 5.02e-19
C290 vss.n137 0 5.02e-19
C291 vss.n138 0 5.02e-19
C292 vss.n140 0 5.02e-19
C293 vss.n141 0 5.02e-19
C294 vss.n143 0 5.02e-19
C295 vss.n144 0 5.02e-19
C296 vss.n146 0 5.02e-19
C297 vss.n147 0 5.02e-19
C298 vss.n149 0 5.02e-19
C299 vss.n150 0 5.02e-19
C300 vss.n152 0 5.02e-19
C301 vss.n153 0 5.02e-19
C302 vss.n155 0 5.02e-19
C303 vss.n156 0 5.02e-19
C304 vss.n158 0 5.02e-19
C305 vss.n159 0 5.02e-19
C306 vss.n161 0 5.02e-19
C307 vss.n162 0 5.02e-19
C308 vss.n164 0 5.02e-19
C309 vss.n165 0 5.02e-19
C310 vss.n168 0 1.28f
C311 vss.n169 0 0.0986f
C312 vss.n170 0 0.00749f
C313 vss.n171 0 0.339f
C314 vss.n173 0 5.02e-19
C315 vss.n175 0 5.02e-19
C316 vss.n176 0 5.02e-19
C317 vss.n178 0 5.02e-19
C318 vss.n179 0 5.02e-19
C319 vss.n181 0 5.02e-19
C320 vss.n182 0 5.02e-19
C321 vss.n184 0 5.02e-19
C322 vss.n185 0 5.02e-19
C323 vss.n187 0 5.02e-19
C324 vss.n188 0 5.02e-19
C325 vss.n190 0 5.02e-19
C326 vss.n191 0 5.02e-19
C327 vss.n193 0 5.02e-19
C328 vss.n194 0 5.02e-19
C329 vss.n196 0 5.02e-19
C330 vss.n197 0 5.02e-19
C331 vss.n199 0 5.02e-19
C332 vss.n200 0 5.02e-19
C333 vss.n202 0 5.02e-19
C334 vss.n203 0 5.02e-19
C335 vss.n205 0 5.02e-19
C336 vss.n206 0 5.02e-19
C337 vss.n208 0 5.02e-19
C338 vss.n209 0 5.02e-19
C339 vss.n211 0 5.02e-19
C340 vss.n212 0 5.02e-19
C341 vss.n214 0 5.02e-19
C342 vss.n215 0 5.02e-19
C343 vss.n217 0 5.02e-19
C344 vss.n218 0 0.00191f
C345 vss.n220 0 0.427f
C346 vss.n221 0 0.114f
C347 vss.n222 0 0.0015f
C348 vss.n223 0 6.27e-20
C349 vss.n224 0 2.1e-19
C350 vss.n225 0 6.27e-20
C351 vss.n226 0 5.02e-19
C352 vss.n227 0 5.02e-19
C353 vss.n228 0 5.02e-19
C354 vss.n229 0 5.02e-19
C355 vss.n230 0 5.02e-19
C356 vss.n231 0 5.02e-19
C357 vss.n232 0 5.02e-19
C358 vss.n233 0 5.02e-19
C359 vss.n234 0 5.02e-19
C360 vss.n235 0 5.02e-19
C361 vss.n236 0 5.02e-19
C362 vss.n237 0 5.02e-19
C363 vss.n238 0 5.02e-19
C364 vss.n239 0 5.02e-19
C365 vss.n240 0 5.02e-19
C366 vss.n241 0 0.00191f
C367 vss.n242 0 0.00189f
C368 vss.n243 0 0.00183f
C369 vss.n244 0 1.96e-19
C370 vss.n245 0 6.27e-20
C371 vss.n246 0 5.02e-19
C372 vss.n247 0 5.02e-19
C373 vss.n248 0 5.02e-19
C374 vss.n249 0 5.02e-19
C375 vss.n250 0 5.02e-19
C376 vss.n251 0 5.02e-19
C377 vss.n252 0 5.02e-19
C378 vss.n253 0 5.02e-19
C379 vss.n254 0 5.02e-19
C380 vss.n255 0 5.02e-19
C381 vss.n256 0 5.02e-19
C382 vss.n257 0 5.02e-19
C383 vss.n258 0 5.02e-19
C384 vss.n259 0 5.02e-19
C385 vss.n260 0 5.02e-19
C386 vss.n261 0 5.02e-19
C387 vss.n262 0 0.00173f
C388 vss.n263 0 0.00155f
C389 vss.n264 0 0.00147f
C390 vss.n265 0 4.67e-19
C391 vss.n266 0 1.56e-19
C392 vss.n267 0 2.93e-19
C393 vss.n268 0 2.67e-19
C394 vss.n269 0 3.78e-19
C395 vss.n270 0 9.11e-20
C396 vss.n271 0 0.00108f
C397 vss.n272 0 3.5e-19
C398 vss.n273 0 3.9e-19
C399 vss.n274 0 3.82e-19
C400 vss.n275 0 6.5e-19
C401 vss.n276 0 4.56e-20
C402 vss.n277 0 1.24e-19
C403 vss.n278 0 5.53e-20
C404 vss.n279 0 2.51e-19
C405 vss.n280 0 0.0299f
C406 vss.n281 0 2.51e-19
C407 vss.n282 0 5.53e-20
C408 vss.n283 0 1.24e-19
C409 vss.n284 0 5.02e-19
C410 vss.n285 0 5.02e-19
C411 vss.n286 0 5.02e-19
C412 vss.n287 0 5.02e-19
C413 vss.n288 0 5.02e-19
C414 vss.n289 0 5.02e-19
C415 vss.n290 0 5.02e-19
C416 vss.n291 0 5.02e-19
C417 vss.n292 0 5.02e-19
C418 vss.n293 0 5.02e-19
C419 vss.n294 0 5.02e-19
C420 vss.n295 0 5.02e-19
C421 vss.n296 0 5.02e-19
C422 vss.n297 0 5.02e-19
C423 vss.n298 0 5.02e-19
C424 vss.n299 0 5.02e-19
C425 vss.n300 0 5.02e-19
C426 vss.n301 0 5.02e-19
C427 vss.n302 0 5.02e-19
C428 vss.n303 0 0.00173f
C429 vss.n304 0 0.00173f
C430 vss.n305 0 0.00169f
C431 vss.n306 0 0.00163f
C432 vss.n307 0 1.96e-19
C433 vss.n308 0 3.78e-19
C434 vss.n309 0 6.27e-20
C435 vss.n310 0 9.11e-20
C436 vss.n311 0 4.56e-20
C437 vss.n312 0 6.5e-19
C438 vss.n313 0 3.82e-19
C439 vss.n314 0 3.9e-19
C440 vss.n315 0 5.02e-19
C441 vss.n316 0 5.02e-19
C442 vss.n317 0 5.02e-19
C443 vss.n318 0 5.02e-19
C444 vss.n319 0 5.02e-19
C445 vss.n320 0 5.02e-19
C446 vss.n321 0 5.02e-19
C447 vss.n322 0 5.02e-19
C448 vss.n323 0 5.02e-19
C449 vss.n324 0 5.02e-19
C450 vss.n325 0 5.02e-19
C451 vss.n326 0 5.02e-19
C452 vss.n327 0 5.02e-19
C453 vss.n328 0 5.02e-19
C454 vss.n329 0 5.02e-19
C455 vss.n330 0 5.02e-19
C456 vss.n331 0 5.02e-19
C457 vss.n332 0 5.02e-19
C458 vss.n333 0 5.02e-19
C459 vss.n334 0 0.00179f
C460 vss.n335 0 0.0016f
C461 vss.n336 0 0.00153f
C462 vss.n337 0 4.67e-19
C463 vss.n338 0 2.67e-19
C464 vss.n339 0 2.93e-19
C465 vss.n340 0 1.56e-19
C466 vss.n341 0 3.5e-19
C467 vss.n342 0 0.00128f
C468 vss.n343 0 0.0857f
C469 vss.n344 0 0.0468f
C470 vss.n345 0 0.0941f
C471 vss.n346 0 5.02e-19
C472 vss.n347 0 5.02e-19
C473 vss.n348 0 5.02e-19
C474 vss.n349 0 5.02e-19
C475 vss.n350 0 5.02e-19
C476 vss.n351 0 5.02e-19
C477 vss.n352 0 5.02e-19
C478 vss.n353 0 5.02e-19
C479 vss.n354 0 5.02e-19
C480 vss.n355 0 5.02e-19
C481 vss.n356 0 5.02e-19
C482 vss.n357 0 5.02e-19
C483 vss.n358 0 5.02e-19
C484 vss.n359 0 5.02e-19
C485 vss.n360 0 5.02e-19
C486 vss.n361 0 5.02e-19
C487 vss.n362 0 5.02e-19
C488 vss.n363 0 5.02e-19
C489 vss.n364 0 5.02e-19
C490 vss.n365 0 5.02e-19
C491 vss.n366 0 5.02e-19
C492 vss.n367 0 5.02e-19
C493 vss.n368 0 5.02e-19
C494 vss.n369 0 5.02e-19
C495 vss.n370 0 5.02e-19
C496 vss.n371 0 5.02e-19
C497 vss.n372 0 5.02e-19
C498 vss.n373 0 5.02e-19
C499 vss.n374 0 5.02e-19
C500 vss.n375 0 5.02e-19
C501 vss.n376 0 5.02e-19
C502 vss.n377 0 5.02e-19
C503 vss.n378 0 0.00173f
C504 vss.n379 0 0.00173f
C505 vss.n380 0 0.00163f
C506 vss.n381 0 1.96e-19
C507 vss.n382 0 3.84e-19
C508 vss.n383 0 6.27e-20
C509 vss.n384 0 8.46e-20
C510 vss.n385 0 2.1e-19
C511 vss.n386 0 6.27e-20
C512 vss.n387 0 0.0215f
C513 vss.n388 0 0.0215f
C514 vss.n389 0 0.0215f
C515 vss.n390 0 5.02e-19
C516 vss.n391 0 0.031f
C517 vss.n392 0 0.00172f
C518 vss.n393 0 0.0538f
C519 vss.n394 0 0.00171f
C520 vss.n396 0 6.27e-20
C521 vss.n397 0 5.92e-19
C522 vss.n398 0 5.02e-19
C523 vss.n399 0 5.02e-19
C524 vss.n400 0 0.00195f
C525 vss.n401 0 0.00178f
C526 vss.n402 0 0.00169f
C527 vss.n403 0 0.00858f
C528 vss.n404 0 0.0086f
C529 vss.n405 0 0.002f
C530 vss.n406 0 0.00183f
C531 vss.n407 0 0.00175f
C532 vss.n408 0 5.77e-19
C533 vss.n409 0 1.81e-19
C534 vss.n410 0 6.27e-20
C535 vss.n411 0 0.00176f
C536 vss.n413 0 6.27e-20
C537 vss.n414 0 0.0215f
C538 vss.n415 0 0.0215f
C539 vss.n416 0 5.02e-19
C540 vss.n417 0 0.0335f
C541 vss.n418 0 0.00174f
C542 vss.n419 0 0.0557f
C543 vss.n420 0 0.00179f
C544 vss.n421 0 0.00175f
C545 vss.n423 0 0.261f
C546 vss.n424 0 0.0652f
C547 vss.n425 0 0.00153f
C548 vss.n426 0 9.46e-20
C549 vss.n427 0 0.00173f
C550 vss.n428 0 0.00169f
C551 vss.n429 0 0.00148f
C552 vss.n430 0 6.53e-19
C553 vss.n431 0 5.02e-19
C554 vss.n432 0 5.02e-19
C555 vss.n433 0 5.02e-19
C556 vss.n434 0 5.02e-19
C557 vss.n435 0 0.00179f
C558 vss.n436 0 5.78e-19
C559 vss.n437 0 5.02e-19
C560 vss.n438 0 5.02e-19
C561 vss.n439 0 5.02e-19
C562 vss.n440 0 0.00174f
C563 vss.n441 0 0.00175f
C564 vss.n442 0 0.00127f
C565 vss.n443 0 0.00435f
C566 vss.n444 0 0.00711f
C567 vss.n445 0 6.71e-19
C568 vss.n446 0 2.36e-19
C569 vss.n447 0 6.81e-19
C570 vss.n448 0 0.00436f
C571 vss.n449 0 0.0103f
C572 vss.n450 0 0.00436f
C573 vss.n451 0 6.24e-19
C574 vss.n452 0 5.02e-19
C575 vss.n453 0 5.02e-19
C576 vss.n454 0 5.02e-19
C577 vss.n455 0 0.00172f
C578 vss.n456 0 0.00173f
C579 vss.n457 0 0.00127f
C580 vss.n458 0 5.02e-19
C581 vss.n459 0 5.02e-19
C582 vss.n460 0 5.02e-19
C583 vss.n461 0 5.02e-19
C584 vss.n462 0 0.00177f
C585 vss.n463 0 5.58e-19
C586 vss.n464 0 0.00433f
C587 vss.n465 0 0.00711f
C588 vss.n466 0 6.79e-19
C589 vss.n467 0 2.85e-19
C590 vss.n468 0 6.53e-19
C591 vss.n469 0 5.02e-19
C592 vss.n470 0 5.02e-19
C593 vss.n471 0 0.00168f
C594 vss.n472 0 0.00164f
C595 vss.n473 0 0.00143f
C596 vss.n474 0 1.81e-19
C597 vss.n475 0 6.27e-20
C598 vss.n476 0 9.46e-20
C599 vss.n477 0 0.00148f
C600 vss.n478 0 0.0633f
C601 vss.n479 0 0.00173f
C602 vss.n480 0 0.00177f
C603 vss.n482 0 0.258f
C604 vss.n483 0 0.257f
C605 vss.n484 0 0.0344f
C606 vss.n485 0 0.0584f
C607 vss.n486 0 0.0584f
C608 vss.n487 0 0.0584f
C609 vss.n488 0 0.0584f
C610 vss.n489 0 0.0584f
C611 vss.n490 0 0.0584f
C612 vss.n491 0 0.0584f
C613 vss.n492 0 0.0584f
C614 vss.n493 0 0.115f
C615 vss.n494 0 0.631f
C616 vss.n495 0 0.0017f
C617 vss.n497 0 0.00156f
C618 vss.n499 0 6.27e-20
C619 vss.n500 0 2.51e-19
C620 vss.n501 0 5.53e-20
C621 vss.n502 0 1.3e-19
C622 vss.n503 0 5.21e-20
C623 vss.n504 0 6.59e-19
C624 vss.n505 0 3.9e-19
C625 vss.n506 0 3.82e-19
C626 vss.n507 0 2.67e-19
C627 vss.n508 0 2.86e-19
C628 vss.n509 0 0.0584f
C629 vss.n510 0 5.02e-19
C630 vss.n511 0 5.02e-19
C631 vss.n512 0 0.0584f
C632 vss.n513 0 5.02e-19
C633 vss.n514 0 5.02e-19
C634 vss.n515 0 0.0584f
C635 vss.n516 0 5.02e-19
C636 vss.n517 0 5.02e-19
C637 vss.n518 0 0.0584f
C638 vss.n519 0 5.02e-19
C639 vss.n520 0 5.02e-19
C640 vss.n521 0 0.0584f
C641 vss.n522 0 5.02e-19
C642 vss.n523 0 5.02e-19
C643 vss.n524 0 0.0584f
C644 vss.n525 0 5.02e-19
C645 vss.n526 0 5.02e-19
C646 vss.n527 0 0.0533f
C647 vss.n528 0 5.02e-19
C648 vss.n529 0 5.02e-19
C649 vss.n530 0 5.02e-19
C650 vss.n531 0 5.02e-19
C651 vss.n532 0 5.02e-19
C652 vss.n533 0 5.02e-19
C653 vss.n534 0 5.02e-19
C654 vss.n535 0 5.02e-19
C655 vss.n536 0 5.02e-19
C656 vss.n537 0 5.02e-19
C657 vss.n538 0 5.02e-19
C658 vss.n539 0 5.02e-19
C659 vss.n540 0 5.02e-19
C660 vss.n541 0 5.02e-19
C661 vss.n542 0 5.02e-19
C662 vss.n543 0 5.02e-19
C663 vss.n544 0 5.02e-19
C664 vss.n545 0 5.02e-19
C665 vss.n546 0 5.02e-19
C666 vss.n547 0 5.02e-19
C667 vss.n548 0 0.00178f
C668 vss.n549 0 0.0016f
C669 vss.n550 0 0.00153f
C670 vss.n551 0 4.67e-19
C671 vss.n552 0 1.5e-19
C672 vss.n553 0 3.5e-19
C673 vss.n554 0 0.00127f
C674 vss.n555 0 0.117f
C675 vss.n556 0 0.0558f
C676 clk 0 3.16f
C677 vdd 0 6.93f
C678 outn 0 1.31f
C679 comparator_core_0/w_302_2337# 0 4.58f
C680 vn 0 1.56f
C681 vp 0 1.55f
C682 outp 0 1.31f
C683 comparator_core_0/diff 0 0.13f
C684 trim_1/n1 0 0.237f
C685 trim_1/n0 0 0.224f
C686 trim_1/drain 0 -3.83f
C687 trimb_2 0 0.531f
C688 trim_1/n3 0 1.39f
C689 trimb_3 0 1.47f
C690 trimb_1 0 0.359f
C691 trim_1/n4 0 1.98f
C692 trimb_4 0 1.4f
C693 trimb_0 0 0.357f
C694 trim_1/n2 0 0.746f
C695 trim_0/n1 0 0.237f
C696 trim_0/n0 0 0.224f
C697 trim_0/drain 0 -3.86f
C698 trim_2 0 0.531f
C699 trim_0/n3 0 1.39f
C700 vss 0 5.64f
C701 trim_3 0 1.47f
C702 trim_1 0 0.359f
C703 trim_0/n4 0 1.98f
C704 trim_4 0 1.4f
C705 trim_0 0 0.357f
C706 trim_0/n2 0 0.746f
.ends

