* SPICE3 file created from DAC.ext - technology: sky130B

.subckt inv2 w_0_269# a_67_305# a_59_207# a_149_55# a_67_55# VSUBS
X0 a_67_55# a_59_207# a_149_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_149_55# a_59_207# a_67_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_67_305# a_59_207# a_149_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_149_55# a_59_207# a_67_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
C0 w_0_269# a_67_305# 0.0521f
C1 w_0_269# a_149_55# 0.0061f
C2 a_59_207# a_67_55# 0.0638f
C3 a_59_207# a_67_305# 0.0631f
C4 a_59_207# a_149_55# 0.0894f
C5 a_59_207# w_0_269# 0.0742f
C6 a_67_55# a_67_305# 0.0423f
C7 a_67_55# a_149_55# 0.155f
C8 a_149_55# a_67_305# 0.209f
C9 a_67_55# w_0_269# 0.00649f
C10 a_67_55# VSUBS 0.266f
C11 a_149_55# VSUBS 0.0332f
C12 a_67_305# VSUBS 0.246f
C13 a_59_207# VSUBS 0.263f
C14 w_0_269# VSUBS 0.339f
.ends

.subckt decap_8 a_65_55# a_65_331# w_0_269# VSUBS
X0 a_65_55# a_65_331# a_65_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
X1 a_65_331# a_65_55# a_65_331# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=2.89
C0 a_65_55# a_65_331# 1.27f
C1 a_65_55# w_0_269# 0.22f
C2 a_65_331# w_0_269# 0.105f
C3 a_65_331# VSUBS 1.14f
C4 a_65_55# VSUBS 0.992f
C5 w_0_269# VSUBS 0.782f
.ends

.subckt M1_3 a_207_n176# a_n29_n176# a_26_55# a_n328_55# a_89_n176# a_n446_55# a_n564_55#
+ a_n210_55# a_n501_n176# a_561_n176# a_n383_n176# a_498_55# a_144_55# a_443_n176#
+ a_n265_n176# a_262_55# a_380_55# a_n619_n176# a_n92_55# w_n757_n324# a_325_n176#
+ a_n147_n176# VSUBS
X0 a_n383_n176# a_n446_55# a_n501_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 a_n29_n176# a_n92_55# a_n147_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 a_325_n176# a_262_55# a_207_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 a_561_n176# a_498_55# a_443_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X4 a_n265_n176# a_n328_55# a_n383_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X5 a_89_n176# a_26_55# a_n29_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 a_207_n176# a_144_55# a_89_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_n501_n176# a_n564_55# a_n619_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X8 a_n147_n176# a_n210_55# a_n265_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X9 a_443_n176# a_380_55# a_325_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
C0 a_n147_n176# a_n210_55# 0.0116f
C1 a_n564_55# a_n501_n176# 0.0116f
C2 w_n757_n324# a_207_n176# 0.0274f
C3 w_n757_n324# a_380_55# 0.105f
C4 a_325_n176# a_443_n176# 0.121f
C5 a_89_n176# a_207_n176# 0.121f
C6 w_n757_n324# a_26_55# 0.105f
C7 a_89_n176# a_26_55# 0.0116f
C8 a_n446_55# a_n383_n176# 0.0116f
C9 w_n757_n324# a_144_55# 0.104f
C10 w_n757_n324# a_325_n176# 0.0258f
C11 a_89_n176# a_144_55# 0.0116f
C12 a_262_55# a_207_n176# 0.0116f
C13 a_n92_55# a_n29_n176# 0.0116f
C14 a_262_55# a_380_55# 0.0657f
C15 a_n564_55# a_n446_55# 0.0657f
C16 a_n501_n176# a_n619_n176# 0.121f
C17 w_n757_n324# a_443_n176# 0.0247f
C18 w_n757_n324# a_n29_n176# 0.0238f
C19 w_n757_n324# a_n92_55# 0.105f
C20 a_n29_n176# a_89_n176# 0.121f
C21 a_262_55# a_144_55# 0.0657f
C22 a_262_55# a_325_n176# 0.0116f
C23 a_n265_n176# a_n328_55# 0.0116f
C24 a_n147_n176# a_n29_n176# 0.121f
C25 w_n757_n324# a_89_n176# 0.0258f
C26 a_n147_n176# a_n92_55# 0.0116f
C27 a_498_55# a_380_55# 0.0657f
C28 a_n265_n176# a_n210_55# 0.0116f
C29 a_n147_n176# w_n757_n324# 0.0258f
C30 w_n757_n324# a_262_55# 0.104f
C31 a_n383_n176# w_n757_n324# 0.0258f
C32 a_n446_55# a_n501_n176# 0.0116f
C33 a_n210_55# a_n328_55# 0.0657f
C34 a_n446_55# a_n328_55# 0.0657f
C35 a_n564_55# w_n757_n324# 0.13f
C36 a_498_55# a_443_n176# 0.0116f
C37 a_561_n176# a_443_n176# 0.121f
C38 w_n757_n324# a_498_55# 0.13f
C39 w_n757_n324# a_561_n176# 0.0913f
C40 w_n757_n324# a_n619_n176# 0.0913f
C41 a_n265_n176# w_n757_n324# 0.0274f
C42 a_n501_n176# w_n757_n324# 0.0247f
C43 a_n265_n176# a_n147_n176# 0.121f
C44 w_n757_n324# a_n328_55# 0.104f
C45 a_207_n176# a_144_55# 0.0116f
C46 a_207_n176# a_325_n176# 0.121f
C47 a_380_55# a_325_n176# 0.0116f
C48 a_n210_55# a_n92_55# 0.0657f
C49 a_n265_n176# a_n383_n176# 0.121f
C50 a_144_55# a_26_55# 0.0657f
C51 a_n564_55# a_n619_n176# 0.0116f
C52 w_n757_n324# a_n210_55# 0.104f
C53 a_n446_55# w_n757_n324# 0.105f
C54 a_n501_n176# a_n383_n176# 0.121f
C55 a_380_55# a_443_n176# 0.0116f
C56 a_498_55# a_561_n176# 0.0116f
C57 a_n29_n176# a_26_55# 0.0116f
C58 a_n383_n176# a_n328_55# 0.0116f
C59 a_n92_55# a_26_55# 0.0657f
C60 a_561_n176# VSUBS 0.056f
C61 a_443_n176# VSUBS 0.0249f
C62 a_325_n176# VSUBS 0.0249f
C63 a_207_n176# VSUBS 0.0249f
C64 a_89_n176# VSUBS 0.0249f
C65 a_n29_n176# VSUBS 0.0249f
C66 a_n147_n176# VSUBS 0.0249f
C67 a_n265_n176# VSUBS 0.0249f
C68 a_n383_n176# VSUBS 0.0249f
C69 a_n501_n176# VSUBS 0.0249f
C70 a_n619_n176# VSUBS 0.056f
C71 a_498_55# VSUBS 0.0832f
C72 a_380_55# VSUBS 0.0669f
C73 a_262_55# VSUBS 0.0669f
C74 a_144_55# VSUBS 0.0669f
C75 a_26_55# VSUBS 0.0669f
C76 a_n92_55# VSUBS 0.0669f
C77 a_n210_55# VSUBS 0.0669f
C78 a_n328_55# VSUBS 0.0669f
C79 a_n446_55# VSUBS 0.0669f
C80 a_n564_55# VSUBS 0.0832f
C81 w_n757_n324# VSUBS 3.39f
.ends

.subckt M2_2 a_26_51# a_89_n171# a_n328_51# a_n446_51# a_n564_51# a_n501_n171# a_n210_51#
+ a_561_n171# a_n383_n171# a_498_51# a_443_n171# a_144_51# a_n265_n171# a_262_51#
+ a_n619_n171# a_380_51# a_n92_51# a_n721_n283# a_325_n171# a_n147_n171# a_207_n171#
+ a_n29_n171#
X0 a_89_n171# a_26_51# a_n29_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 a_207_n171# a_144_51# a_89_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 a_n147_n171# a_n210_51# a_n265_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 a_n501_n171# a_n564_51# a_n619_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X4 a_443_n171# a_380_51# a_325_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X5 a_n383_n171# a_n446_51# a_n501_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 a_n29_n171# a_n92_51# a_n147_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_325_n171# a_262_51# a_207_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X8 a_561_n171# a_498_51# a_443_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X9 a_n265_n171# a_n328_51# a_n383_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
C0 a_26_51# a_n29_n171# 0.0116f
C1 a_n210_51# a_n92_51# 0.0633f
C2 a_n446_51# a_n328_51# 0.0633f
C3 a_207_n171# a_262_51# 0.0116f
C4 a_n501_n171# a_n446_51# 0.0116f
C5 a_n265_n171# a_n383_n171# 0.121f
C6 a_144_51# a_26_51# 0.0633f
C7 a_498_51# a_561_n171# 0.0116f
C8 a_n619_n171# a_n501_n171# 0.121f
C9 a_n564_51# a_n446_51# 0.0633f
C10 a_144_51# a_262_51# 0.0633f
C11 a_n147_n171# a_n29_n171# 0.121f
C12 a_n383_n171# a_n328_51# 0.0116f
C13 a_207_n171# a_325_n171# 0.121f
C14 a_n619_n171# a_n564_51# 0.0116f
C15 a_n383_n171# a_n501_n171# 0.121f
C16 a_n147_n171# a_n265_n171# 0.121f
C17 a_380_51# a_262_51# 0.0633f
C18 a_207_n171# a_89_n171# 0.121f
C19 a_n265_n171# a_n328_51# 0.0116f
C20 a_n92_51# a_n29_n171# 0.0116f
C21 a_26_51# a_n92_51# 0.0633f
C22 a_n383_n171# a_n446_51# 0.0116f
C23 a_n265_n171# a_n210_51# 0.0116f
C24 a_89_n171# a_n29_n171# 0.121f
C25 a_262_51# a_325_n171# 0.0116f
C26 a_89_n171# a_26_51# 0.0116f
C27 a_380_51# a_443_n171# 0.0116f
C28 a_144_51# a_89_n171# 0.0116f
C29 a_380_51# a_325_n171# 0.0116f
C30 a_n147_n171# a_n210_51# 0.0116f
C31 a_n328_51# a_n210_51# 0.0633f
C32 a_380_51# a_498_51# 0.0633f
C33 a_n147_n171# a_n92_51# 0.0116f
C34 a_325_n171# a_443_n171# 0.121f
C35 a_561_n171# a_443_n171# 0.121f
C36 a_207_n171# a_144_51# 0.0116f
C37 a_n501_n171# a_n564_51# 0.0116f
C38 a_498_51# a_443_n171# 0.0116f
C39 a_561_n171# a_n721_n283# 0.148f
C40 a_443_n171# a_n721_n283# 0.0499f
C41 a_325_n171# a_n721_n283# 0.051f
C42 a_207_n171# a_n721_n283# 0.0526f
C43 a_89_n171# a_n721_n283# 0.051f
C44 a_n29_n171# a_n721_n283# 0.0489f
C45 a_n147_n171# a_n721_n283# 0.051f
C46 a_n265_n171# a_n721_n283# 0.0526f
C47 a_n383_n171# a_n721_n283# 0.051f
C48 a_n501_n171# a_n721_n283# 0.0499f
C49 a_n619_n171# a_n721_n283# 0.148f
C50 a_498_51# a_n721_n283# 0.208f
C51 a_380_51# a_n721_n283# 0.169f
C52 a_262_51# a_n721_n283# 0.168f
C53 a_144_51# a_n721_n283# 0.168f
C54 a_26_51# a_n721_n283# 0.169f
C55 a_n92_51# a_n721_n283# 0.169f
C56 a_n210_51# a_n721_n283# 0.168f
C57 a_n328_51# a_n721_n283# 0.168f
C58 a_n446_51# a_n721_n283# 0.169f
C59 a_n564_51# a_n721_n283# 0.208f
.ends

.subckt inv_4 w_0_269# a_59_207# a_75_55# a_75_305# a_157_55# VSUBS
X0 a_75_55# a_59_207# a_157_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_75_305# a_59_207# a_157_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_157_55# a_59_207# a_75_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_157_55# a_59_207# a_75_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_157_55# a_59_207# a_75_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_75_305# a_59_207# a_157_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_75_55# a_59_207# a_157_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_157_55# a_59_207# a_75_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
C0 a_75_55# w_0_269# 0.00667f
C1 w_0_269# a_75_305# 0.0654f
C2 a_75_55# a_59_207# 0.0819f
C3 a_59_207# a_75_305# 0.0982f
C4 a_59_207# w_0_269# 0.142f
C5 a_75_55# a_157_55# 0.263f
C6 a_157_55# a_75_305# 0.362f
C7 w_0_269# a_157_55# 0.0159f
C8 a_75_55# a_75_305# 0.0501f
C9 a_59_207# a_157_55# 0.36f
C10 a_75_55# VSUBS 0.327f
C11 a_157_55# VSUBS 0.0849f
C12 a_75_305# VSUBS 0.296f
C13 a_59_207# VSUBS 0.452f
C14 w_0_269# VSUBS 0.516f
.ends

.subckt decap_3 a_65_55# a_65_331# w_0_269# VSUBS
X0 a_65_55# a_65_331# a_65_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
X1 a_65_331# a_65_55# a_65_331# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
C0 a_65_55# w_0_269# 0.0797f
C1 a_65_331# w_0_269# 0.0625f
C2 a_65_55# a_65_331# 0.353f
C3 a_65_331# VSUBS 0.47f
C4 a_65_55# VSUBS 0.427f
C5 w_0_269# VSUBS 0.339f
.ends

.subckt sw_top en m2_1158_361# inv_4_1/w_0_269# out vdd in m2_990_200# vss
Xdecap_8_0 vss vdd inv_4_1/w_0_269# vss decap_8
XM1_3_0 out out m2_1158_361# m2_1158_361# in m2_1158_361# m2_1158_361# m2_1158_361#
+ out in in m2_1158_361# m2_1158_361# out out m2_1158_361# m2_1158_361# in m2_1158_361#
+ vdd in in vss M1_3
XM2_2_0 m2_990_200# in m2_990_200# m2_990_200# m2_990_200# out m2_990_200# in in m2_990_200#
+ out m2_990_200# out m2_990_200# in m2_990_200# m2_990_200# vss in in out out M2_2
Xinv_4_0 inv_4_1/w_0_269# m2_1158_361# vss vdd m2_990_200# vss inv_4
Xinv_4_1 inv_4_1/w_0_269# en vss vdd m2_1158_361# vss inv_4
Xdecap_3_0 vss vdd inv_4_1/w_0_269# vss decap_3
C0 inv_4_1/w_0_269# in 0.00429f
C1 en out 0.00102f
C2 en m2_1158_361# 0.0462f
C3 m2_990_200# inv_4_1/w_0_269# 0.0334f
C4 en vdd 0.0728f
C5 in out 2.9f
C6 in m2_1158_361# 0.348f
C7 m2_990_200# out 0.165f
C8 m2_990_200# m2_1158_361# 0.421f
C9 vdd in 0.42f
C10 inv_4_1/w_0_269# m2_1158_361# 0.0248f
C11 vdd m2_990_200# 0.35f
C12 vdd inv_4_1/w_0_269# -0.0142f
C13 en in 0.0109f
C14 out m2_1158_361# 0.307f
C15 en m2_990_200# 0.0721f
C16 vdd out 0.218f
C17 en inv_4_1/w_0_269# 0.00729f
C18 vdd m2_1158_361# 0.374f
C19 m2_990_200# in 0.249f
C20 en vss 0.581f
C21 vdd vss 5.69f
C22 m2_990_200# vss 2.04f
C23 out vss 0.723f
C24 in vss 1.55f
C25 m2_1158_361# vss 1.76f
C26 inv_4_1/w_0_269# vss 1.95f
.ends

.subckt C7 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 m3_n450_n340# c1_n250_n240# 0.503f
C1 c1_n250_n240# VSUBS 0.199f
C2 m3_n450_n340# VSUBS 0.653f
.ends

.subckt DUMMY m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 m3_n450_n340# c1_n250_n240# 0.503f
C1 c1_n250_n240# VSUBS 0.199f
C2 m3_n450_n340# VSUBS 0.653f
.ends

.subckt C6 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 m3_n450_n340# c1_n250_n240# 0.503f
C1 c1_n250_n240# VSUBS 0.199f
C2 m3_n450_n340# VSUBS 0.653f
.ends

.subckt CDUM m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 m3_n450_n340# c1_n250_n240# 0.503f
C1 c1_n250_n240# VSUBS 0.199f
C2 m3_n450_n340# VSUBS 0.653f
.ends

.subckt C4 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 m3_n450_n340# c1_n250_n240# 0.503f
C1 c1_n250_n240# VSUBS 0.199f
C2 m3_n450_n340# VSUBS 0.653f
.ends

.subckt C2 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 m3_n450_n340# c1_n250_n240# 0.503f
C1 c1_n250_n240# VSUBS 0.199f
C2 m3_n450_n340# VSUBS 0.653f
.ends

.subckt C5 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 m3_n450_n340# c1_n250_n240# 0.503f
C1 c1_n250_n240# VSUBS 0.199f
C2 m3_n450_n340# VSUBS 0.653f
.ends

.subckt C3 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 m3_n450_n340# c1_n250_n240# 0.503f
C1 c1_n250_n240# VSUBS 0.199f
C2 m3_n450_n340# VSUBS 0.653f
.ends

.subckt C1 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 m3_n450_n340# c1_n250_n240# 0.503f
C1 c1_n250_n240# VSUBS 0.199f
C2 m3_n450_n340# VSUBS 0.653f
.ends

.subckt C0_1 m3_n450_n340# c1_n250_n240# VSUBS
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
C0 m3_n450_n340# c1_n250_n240# 0.503f
C1 c1_n250_n240# VSUBS 0.199f
C2 m3_n450_n340# VSUBS 0.653f
.ends

.subckt carray n2 n3 n0 via23_4_702/m2_1_40# m2_800_1156# via23_4_459/m2_1_40# m2_27200_1156#
+ m2_23300_1156# m2_28500_1156# via23_4_447/m2_1_40# m2_24600_1156# m2_29800_1156#
+ m2_35000_1156# m2_31100_1156# m2_25900_1156# via23_4_369/m2_1_40# m2_36300_1156#
+ via23_4_379/m2_1_40# m2_32400_1156# m2_37600_1156# m3_42700_1156# m2_33700_1156#
+ m2_38900_1156# m3_900_1156# via23_4_635/m2_1_40# via23_4_455/m2_1_40# via23_4_414/m2_1_40#
+ via23_4_439/m2_1_40# m2_40200_1156# via23_4_460/m2_1_40# via23_4_704/m2_1_40# m2_41500_1156#
+ via23_4_366/m2_1_40# via23_4_429/m2_1_40# m2_42800_1156# n4 via23_4_128/m2_1_40#
+ via23_4_458/m2_1_40# ndum via23_4_381/m2_1_40# via23_4_419/m2_1_40# via23_4_449/m2_1_40#
+ via23_4_641/m2_1_40# via23_4_378/m2_1_40# n1 n6 via23_4_642/m2_1_40# via23_4_368/m2_1_40#
+ via23_4_705/m2_1_40# via23_4_446/m2_1_40# via23_4_96/m2_1_40# top n5 via23_4_448/m2_1_40#
+ m3_42500_1156# VSUBS via23_4_380/m2_1_40# n7 via23_4_367/m2_1_40#
XC7_121 n7 top VSUBS C7
XC7_110 n7 top VSUBS C7
XDUMMY_80 via23_4_712/m2_1_40# top VSUBS DUMMY
XC6_20 n6 top VSUBS C6
XC6_53 n6 top VSUBS C6
XC6_31 n6 top VSUBS C6
XC6_42 n6 top VSUBS C6
XC7_122 n7 top VSUBS C7
XC7_100 n7 top VSUBS C7
XC7_111 n7 top VSUBS C7
XDUMMY_81 via23_4_709/m2_1_40# top VSUBS DUMMY
XDUMMY_70 via23_4_642/m2_1_40# top VSUBS DUMMY
XC6_21 n6 top VSUBS C6
XC6_10 n6 top VSUBS C6
XC6_54 n6 top VSUBS C6
XC6_32 n6 top VSUBS C6
XC6_43 n6 top VSUBS C6
XC6_0 n6 top VSUBS C6
XC7_123 n7 top VSUBS C7
XC7_101 n7 top VSUBS C7
XC7_112 n7 top VSUBS C7
XDUMMY_71 via23_4_641/m2_1_40# top VSUBS DUMMY
XDUMMY_82 via23_4_439/m2_1_40# top VSUBS DUMMY
XDUMMY_60 via23_4_448/m2_1_40# top VSUBS DUMMY
XC6_44 n6 top VSUBS C6
XC6_22 n6 top VSUBS C6
XC6_55 n6 top VSUBS C6
XC6_11 n6 top VSUBS C6
XC6_33 n6 top VSUBS C6
XC6_1 n6 top VSUBS C6
XC7_124 n7 top VSUBS C7
XC7_102 n7 top VSUBS C7
XC7_113 n7 top VSUBS C7
XDUMMY_72 via23_4_676/m2_1_40# top VSUBS DUMMY
XDUMMY_83 via23_4_675/m2_1_40# top VSUBS DUMMY
XDUMMY_61 via23_4_588/m2_1_40# top VSUBS DUMMY
XDUMMY_50 via23_4_429/m2_1_40# top VSUBS DUMMY
XC6_56 n6 top VSUBS C6
XC6_12 n6 top VSUBS C6
XC6_45 n6 top VSUBS C6
XC6_23 n6 top VSUBS C6
XC6_34 n6 top VSUBS C6
XC6_2 n6 top VSUBS C6
XCDUM_0 ndum top VSUBS CDUM
XC7_103 n7 top VSUBS C7
XC7_125 n7 top VSUBS C7
XC7_114 n7 top VSUBS C7
XDUMMY_73 via23_4_677/m2_1_40# top VSUBS DUMMY
XDUMMY_62 via23_4_589/m2_1_40# top VSUBS DUMMY
XDUMMY_40 via23_4_326/m2_1_40# top VSUBS DUMMY
XDUMMY_51 via23_4_414/m2_1_40# top VSUBS DUMMY
XC6_57 n6 top VSUBS C6
XC6_24 n6 top VSUBS C6
XC6_46 n6 top VSUBS C6
XC6_13 n6 top VSUBS C6
XC6_35 n6 top VSUBS C6
XDUMMY_0 via23_4_3/m2_1_40# top VSUBS DUMMY
XC6_3 n6 top VSUBS C6
XC4_0 n4 top VSUBS C4
XC7_104 n7 top VSUBS C7
XC7_115 n7 top VSUBS C7
XC7_126 n7 top VSUBS C7
XDUMMY_74 via23_4_678/m2_1_40# top VSUBS DUMMY
XDUMMY_63 via23_4_590/m2_1_40# top VSUBS DUMMY
XDUMMY_30 via23_4_251/m2_1_40# top VSUBS DUMMY
XDUMMY_52 via23_4_381/m2_1_40# top VSUBS DUMMY
XDUMMY_41 via23_4_89/m2_1_40# top VSUBS DUMMY
XC6_47 n6 top VSUBS C6
XC6_14 n6 top VSUBS C6
XC6_58 n6 top VSUBS C6
XC6_25 n6 top VSUBS C6
XC6_36 n6 top VSUBS C6
XDUMMY_1 via23_4_9/m2_1_40# top VSUBS DUMMY
XC7_90 n7 top VSUBS C7
XC6_4 n6 top VSUBS C6
XC4_1 n4 top VSUBS C4
XC7_116 n7 top VSUBS C7
XC7_105 n7 top VSUBS C7
XC7_127 n7 top VSUBS C7
XDUMMY_20 via23_4_199/m2_1_40# top VSUBS DUMMY
XDUMMY_64 via23_4_584/m2_1_40# top VSUBS DUMMY
XDUMMY_31 via23_4_245/m2_1_40# top VSUBS DUMMY
XDUMMY_75 via23_4_704/m2_1_40# top VSUBS DUMMY
XDUMMY_42 via23_4_366/m2_1_40# top VSUBS DUMMY
XDUMMY_53 via23_4_449/m2_1_40# top VSUBS DUMMY
XC6_26 n6 top VSUBS C6
XC6_15 n6 top VSUBS C6
XC6_59 n6 top VSUBS C6
XC6_48 n6 top VSUBS C6
XDUMMY_2 via23_4_1/m2_1_40# top VSUBS DUMMY
XC6_37 n6 top VSUBS C6
XC7_91 n7 top VSUBS C7
XC7_80 n7 top VSUBS C7
XC6_5 n6 top VSUBS C6
XC4_2 n4 top VSUBS C4
XC7_117 n7 top VSUBS C7
XC7_106 n7 top VSUBS C7
XDUMMY_76 via23_4_702/m2_1_40# top VSUBS DUMMY
XDUMMY_65 via23_4_600/m2_1_40# top VSUBS DUMMY
XDUMMY_32 via23_4_331/m2_1_40# top VSUBS DUMMY
XDUMMY_21 via23_4_198/m2_1_40# top VSUBS DUMMY
XDUMMY_43 via23_4_367/m2_1_40# top VSUBS DUMMY
XDUMMY_54 via23_4_446/m2_1_40# top VSUBS DUMMY
XDUMMY_10 via23_4_90/m2_1_40# top VSUBS DUMMY
XC6_27 n6 top VSUBS C6
XC6_16 n6 top VSUBS C6
XC6_49 n6 top VSUBS C6
XC6_38 n6 top VSUBS C6
XDUMMY_3 via23_4_2/m2_1_40# top VSUBS DUMMY
XC7_92 n7 top VSUBS C7
XC7_81 n7 top VSUBS C7
XC7_70 n7 top VSUBS C7
XC6_6 n6 top VSUBS C6
XC4_3 n4 top VSUBS C4
XC7_118 n7 top VSUBS C7
XC7_107 n7 top VSUBS C7
XC2_0 n2 top VSUBS C2
XDUMMY_66 via23_4_601/m2_1_40# top VSUBS DUMMY
XDUMMY_33 via23_4_332/m2_1_40# top VSUBS DUMMY
XDUMMY_22 via23_4_220/m2_1_40# top VSUBS DUMMY
XDUMMY_77 via23_4_705/m2_1_40# top VSUBS DUMMY
XDUMMY_44 via23_4_368/m2_1_40# top VSUBS DUMMY
XDUMMY_55 via23_4_447/m2_1_40# top VSUBS DUMMY
XDUMMY_11 via23_4_96/m2_1_40# top VSUBS DUMMY
XC6_28 n6 top VSUBS C6
XC6_17 n6 top VSUBS C6
XC6_39 n6 top VSUBS C6
XDUMMY_4 via23_4_20/m2_1_40# top VSUBS DUMMY
XC7_60 n7 top VSUBS C7
XC7_93 n7 top VSUBS C7
XC7_82 n7 top VSUBS C7
XC7_71 n7 top VSUBS C7
XC6_7 n6 top VSUBS C6
XC4_4 n4 top VSUBS C4
XC7_119 n7 top VSUBS C7
XC7_108 n7 top VSUBS C7
XC2_1 n2 top VSUBS C2
XDUMMY_78 via23_4_710/m2_1_40# top VSUBS DUMMY
XDUMMY_67 via23_4_599/m2_1_40# top VSUBS DUMMY
XDUMMY_34 via23_4_333/m2_1_40# top VSUBS DUMMY
XDUMMY_23 via23_4_213/m2_1_40# top VSUBS DUMMY
XDUMMY_45 via23_4_369/m2_1_40# top VSUBS DUMMY
XDUMMY_56 via23_4_458/m2_1_40# top VSUBS DUMMY
XDUMMY_12 via23_4_103/m2_1_40# top VSUBS DUMMY
XC6_18 n6 top VSUBS C6
XC6_29 n6 top VSUBS C6
XDUMMY_5 via23_4_21/m2_1_40# top VSUBS DUMMY
XC7_61 n7 top VSUBS C7
XC7_94 n7 top VSUBS C7
XC7_50 n7 top VSUBS C7
XC7_72 n7 top VSUBS C7
XC7_83 n7 top VSUBS C7
XC6_8 n6 top VSUBS C6
XC4_5 n4 top VSUBS C4
XC7_109 n7 top VSUBS C7
XC2_2 n2 top VSUBS C2
XDUMMY_79 via23_4_711/m2_1_40# top VSUBS DUMMY
XDUMMY_68 via23_4_598/m2_1_40# top VSUBS DUMMY
XDUMMY_35 via23_4_347/m2_1_40# top VSUBS DUMMY
XDUMMY_24 via23_4_229/m2_1_40# top VSUBS DUMMY
XDUMMY_46 via23_4_378/m2_1_40# top VSUBS DUMMY
XDUMMY_57 via23_4_455/m2_1_40# top VSUBS DUMMY
XDUMMY_13 via23_4_91/m2_1_40# top VSUBS DUMMY
XC6_19 n6 top VSUBS C6
XDUMMY_6 via23_4_22/m2_1_40# top VSUBS DUMMY
XC7_62 n7 top VSUBS C7
XC7_40 n7 top VSUBS C7
XC7_95 n7 top VSUBS C7
XC7_51 n7 top VSUBS C7
XC7_73 n7 top VSUBS C7
XC7_84 n7 top VSUBS C7
XC6_9 n6 top VSUBS C6
XC4_6 n4 top VSUBS C4
XC2_3 n2 top VSUBS C2
XDUMMY_36 via23_4_354/m2_1_40# top VSUBS DUMMY
XDUMMY_25 via23_4_228/m2_1_40# top VSUBS DUMMY
XDUMMY_14 via23_4_94/m2_1_40# top VSUBS DUMMY
XDUMMY_69 via23_4_635/m2_1_40# top VSUBS DUMMY
XDUMMY_47 via23_4_379/m2_1_40# top VSUBS DUMMY
XDUMMY_58 via23_4_459/m2_1_40# top VSUBS DUMMY
XDUMMY_7 via23_4_23/m2_1_40# top VSUBS DUMMY
XC7_41 n7 top VSUBS C7
XC7_63 n7 top VSUBS C7
XC7_96 n7 top VSUBS C7
XC7_52 n7 top VSUBS C7
XC7_30 n7 top VSUBS C7
XC7_74 n7 top VSUBS C7
XC7_85 n7 top VSUBS C7
XC4_7 n4 top VSUBS C4
XDUMMY_37 via23_4_345/m2_1_40# top VSUBS DUMMY
XDUMMY_26 via23_4_230/m2_1_40# top VSUBS DUMMY
XDUMMY_48 via23_4_380/m2_1_40# top VSUBS DUMMY
XDUMMY_59 via23_4_460/m2_1_40# top VSUBS DUMMY
XDUMMY_15 via23_4_117/m2_1_40# top VSUBS DUMMY
XDUMMY_8 via23_4_87/m2_1_40# top VSUBS DUMMY
XC7_97 n7 top VSUBS C7
XC7_42 n7 top VSUBS C7
XC7_53 n7 top VSUBS C7
XC7_31 n7 top VSUBS C7
XC7_86 n7 top VSUBS C7
XC7_20 n7 top VSUBS C7
XC7_64 n7 top VSUBS C7
XC7_75 n7 top VSUBS C7
XC4_10 n4 top VSUBS C4
XC4_8 n4 top VSUBS C4
XDUMMY_38 via23_4_346/m2_1_40# top VSUBS DUMMY
XDUMMY_27 via23_4_218/m2_1_40# top VSUBS DUMMY
XDUMMY_16 via23_4_111/m2_1_40# top VSUBS DUMMY
XDUMMY_49 via23_4_419/m2_1_40# top VSUBS DUMMY
XDUMMY_9 via23_4_88/m2_1_40# top VSUBS DUMMY
XC7_98 n7 top VSUBS C7
XC7_43 n7 top VSUBS C7
XC7_54 n7 top VSUBS C7
XC7_32 n7 top VSUBS C7
XC7_87 n7 top VSUBS C7
XC7_65 n7 top VSUBS C7
XC7_10 n7 top VSUBS C7
XC7_21 n7 top VSUBS C7
XC7_76 n7 top VSUBS C7
XC4_11 n4 top VSUBS C4
XC4_9 n4 top VSUBS C4
XDUMMY_39 via23_4_334/m2_1_40# top VSUBS DUMMY
XDUMMY_28 via23_4_249/m2_1_40# top VSUBS DUMMY
XDUMMY_17 via23_4_128/m2_1_40# top VSUBS DUMMY
XC7_99 n7 top VSUBS C7
XC7_33 n7 top VSUBS C7
XC7_88 n7 top VSUBS C7
XC7_55 n7 top VSUBS C7
XC7_44 n7 top VSUBS C7
XC7_66 n7 top VSUBS C7
XC7_11 n7 top VSUBS C7
XC7_77 n7 top VSUBS C7
XC7_22 n7 top VSUBS C7
XC4_12 n4 top VSUBS C4
XDUMMY_29 via23_4_250/m2_1_40# top VSUBS DUMMY
XDUMMY_18 via23_4_95/m2_1_40# top VSUBS DUMMY
XC7_45 n7 top VSUBS C7
XC7_56 n7 top VSUBS C7
XC7_34 n7 top VSUBS C7
XC7_89 n7 top VSUBS C7
XC7_12 n7 top VSUBS C7
XC7_23 n7 top VSUBS C7
XC7_78 n7 top VSUBS C7
XC7_67 n7 top VSUBS C7
XC4_13 n4 top VSUBS C4
XDUMMY_19 via23_4_200/m2_1_40# top VSUBS DUMMY
XC7_46 n7 top VSUBS C7
XC7_57 n7 top VSUBS C7
XC7_24 n7 top VSUBS C7
XC7_35 n7 top VSUBS C7
XC7_13 n7 top VSUBS C7
XC7_79 n7 top VSUBS C7
XC7_68 n7 top VSUBS C7
XC4_14 n4 top VSUBS C4
XC7_36 n7 top VSUBS C7
XC7_58 n7 top VSUBS C7
XC7_47 n7 top VSUBS C7
XC7_25 n7 top VSUBS C7
XC7_14 n7 top VSUBS C7
XC7_69 n7 top VSUBS C7
XC4_15 n4 top VSUBS C4
XC7_0 n7 top VSUBS C7
XC7_37 n7 top VSUBS C7
XC7_59 n7 top VSUBS C7
XC7_26 n7 top VSUBS C7
XC7_48 n7 top VSUBS C7
XC7_15 n7 top VSUBS C7
XC7_1 n7 top VSUBS C7
XC7_38 n7 top VSUBS C7
XC7_27 n7 top VSUBS C7
XC7_49 n7 top VSUBS C7
XC7_16 n7 top VSUBS C7
XC7_2 n7 top VSUBS C7
XC7_39 n7 top VSUBS C7
XC7_28 n7 top VSUBS C7
XC7_17 n7 top VSUBS C7
XC7_3 n7 top VSUBS C7
XC5_0 n5 top VSUBS C5
XC7_29 n7 top VSUBS C7
XC7_18 n7 top VSUBS C7
XC7_4 n7 top VSUBS C7
XC5_1 n5 top VSUBS C5
XC7_19 n7 top VSUBS C7
XC5_30 n5 top VSUBS C5
XC7_5 n7 top VSUBS C7
XC5_2 n5 top VSUBS C5
XC5_31 n5 top VSUBS C5
XC5_20 n5 top VSUBS C5
XC7_6 n7 top VSUBS C7
XC5_3 n5 top VSUBS C5
XC3_0 n3 top VSUBS C3
XC5_10 n5 top VSUBS C5
XC5_21 n5 top VSUBS C5
XC7_7 n7 top VSUBS C7
XC5_4 n5 top VSUBS C5
XC3_1 n3 top VSUBS C3
XC5_22 n5 top VSUBS C5
XC5_11 n5 top VSUBS C5
XC7_8 n7 top VSUBS C7
XC5_5 n5 top VSUBS C5
XC3_2 n3 top VSUBS C3
XC5_23 n5 top VSUBS C5
XC7_9 n7 top VSUBS C7
XC5_12 n5 top VSUBS C5
XC5_6 n5 top VSUBS C5
XC3_3 n3 top VSUBS C3
XC1_0 n1 top VSUBS C1
XC5_24 n5 top VSUBS C5
XC5_13 n5 top VSUBS C5
XC5_7 n5 top VSUBS C5
XC3_4 n3 top VSUBS C3
XC1_1 n1 top VSUBS C1
XC5_25 n5 top VSUBS C5
XC5_14 n5 top VSUBS C5
XC5_8 n5 top VSUBS C5
XC3_5 n3 top VSUBS C3
XC5_15 n5 top VSUBS C5
XC5_26 n5 top VSUBS C5
XC5_9 n5 top VSUBS C5
XC3_6 n3 top VSUBS C3
XC5_16 n5 top VSUBS C5
XC5_27 n5 top VSUBS C5
XC3_7 n3 top VSUBS C3
XC0_1_0 n0 top VSUBS C0_1
XC5_28 n5 top VSUBS C5
XC5_17 n5 top VSUBS C5
XC6_60 n6 top VSUBS C6
XC5_29 n5 top VSUBS C5
XC5_18 n5 top VSUBS C5
XC6_61 n6 top VSUBS C6
XC6_50 n6 top VSUBS C6
XC5_19 n5 top VSUBS C5
XC6_51 n6 top VSUBS C6
XC6_62 n6 top VSUBS C6
XC6_40 n6 top VSUBS C6
XC7_120 n7 top VSUBS C7
XC6_63 n6 top VSUBS C6
XC6_52 n6 top VSUBS C6
XC6_30 n6 top VSUBS C6
XC6_41 n6 top VSUBS C6
C0 ndum via23_4_584/m2_1_40# 0.247f
C1 via23_4_589/m2_1_40# n7 0.452f
C2 n6 m2_31100_1156# 2.39f
C3 top m2_15100_1156# 0.267f
C4 m3_16500_1156# m3_16700_1156# 3.35f
C5 via23_4_449/m2_1_40# n5 0.0714f
C6 top m3_34900_1156# 0.221f
C7 m3_32100_1156# via23_4_446/m2_1_40# 0.247f
C8 m2_16400_1156# m3_16500_1156# 2.11f
C9 m3_24500_1156# m3_25600_1156# 0.148f
C10 n2 m3_20400_1156# 3.43f
C11 m3_900_1156# via23_4_213/m2_1_40# 0.247f
C12 m2_25900_1156# m3_25800_1156# 2.11f
C13 m3_900_1156# via23_4_200/m2_1_40# 0.247f
C14 ndum m2_15100_1156# 3.15e-20
C15 m3_5000_1156# m3_4800_1156# 3.35f
C16 via23_4_368/m2_1_40# n7 0.452f
C17 m3_900_1156# via23_4_220/m2_1_40# 0.247f
C18 m3_7600_1156# n2 0.021f
C19 m2_23300_1156# m3_23200_1156# 2.11f
C20 top via23_4_331/m2_1_40# 0.347f
C21 top via23_4_334/m2_1_40# 0.347f
C22 m2_15100_1156# m3_15200_1156# 2.11f
C23 via23_4_91/m2_1_40# n5 2.03e-19
C24 top via23_4_705/m2_1_40# 0.216f
C25 top via23_4_230/m2_1_40# 0.347f
C26 m3_39900_1156# n6 0.00746f
C27 n7 n1 10.3f
C28 m2_42800_1156# via23_4_641/m2_1_40# 0.251f
C29 via23_4_378/m2_1_40# m2_33700_1156# 0.251f
C30 n4 n1 0.0766f
C31 n2 via23_4_2/m2_1_40# 0.352f
C32 via23_4_448/m2_1_40# m3_27100_1156# 0.247f
C33 via23_4_229/m2_1_40# m3_1100_1156# 0.247f
C34 top m2_29800_1156# 0.267f
C35 m3_10000_1156# n5 0.181f
C36 via23_4_128/m2_1_40# via23_4_117/m2_1_40# 0.199f
C37 m3_41200_1156# m2_41500_1156# 0.181f
C38 m2_12500_1156# n7 1.13f
C39 m3_32100_1156# n6 4.08f
C40 via23_4_460/m2_1_40# n7 0.452f
C41 top via23_4_346/m2_1_40# 0.347f
C42 via23_4_117/m2_1_40# via23_4_111/m2_1_40# 0.199f
C43 m3_4800_1156# n7 2.16f
C44 m2_12500_1156# n4 3.19e-19
C45 m3_29500_1156# n5 0.00889f
C46 via23_4_455/m2_1_40# n7 9.11e-20
C47 top via23_4_712/m2_1_40# 0.347f
C48 m2_800_1156# via23_4_96/m2_1_40# 0.251f
C49 via23_4_598/m2_1_40# n5 0.452f
C50 via23_4_455/m2_1_40# n4 2.21e-19
C51 m3_6100_1156# via23_4_245/m2_1_40# 0.247f
C52 m2_35000_1156# m3_34700_1156# 0.181f
C53 m2_800_1156# via23_4_198/m2_1_40# 0.251f
C54 m2_41500_1156# n6 1.13f
C55 via23_4_459/m2_1_40# m3_23200_1156# 0.247f
C56 top via23_4_381/m2_1_40# 0.14f
C57 top via23_4_419/m2_1_40# 0.216f
C58 via23_4_250/m2_1_40# m3_7600_1156# 0.247f
C59 m2_2100_1156# via23_4_103/m2_1_40# 0.251f
C60 m3_8700_1156# m3_8900_1156# 3.35f
C61 top via23_4_379/m2_1_40# 0.14f
C62 top m3_38600_1156# 0.187f
C63 m2_9900_1156# n6 1.43e-19
C64 m2_35000_1156# n7 3.52f
C65 m2_7300_1156# via23_4_249/m2_1_40# 0.251f
C66 top m3_19300_1156# 0.187f
C67 m3_16700_1156# m3_17800_1156# 0.354f
C68 via23_4_711/m2_1_40# m2_40200_1156# 0.251f
C69 via23_4_675/m2_1_40# m3_33400_1156# 0.247f
C70 m2_17700_1156# m3_16700_1156# 0.023f
C71 via23_4_1/m2_1_40# m3_19300_1156# 0.247f
C72 via23_4_366/m2_1_40# m3_42500_1156# 0.247f
C73 m3_24500_1156# n7 1.98f
C74 top m3_30800_1156# 0.221f
C75 m3_31000_1156# via23_4_601/m2_1_40# 0.247f
C76 m2_2100_1156# n6 1.13f
C77 top m3_7400_1156# 0.187f
C78 via23_4_251/m2_1_40# n7 0.452f
C79 m3_24500_1156# n4 0.181f
C80 m3_27100_1156# n6 0.181f
C81 m2_7300_1156# n2 0.00855f
C82 m2_19000_1156# n1 8.05e-20
C83 via23_4_448/m2_1_40# n6 1.52e-19
C84 n3 m2_9900_1156# 5.59e-19
C85 m2_8600_1156# n1 8.05e-20
C86 via23_4_599/m2_1_40# m3_28400_1156# 0.247f
C87 top via23_4_590/m2_1_40# 0.347f
C88 m2_9900_1156# m3_8900_1156# 0.0061f
C89 via23_4_345/m2_1_40# n6 0.452f
C90 m3_42700_1156# via23_4_414/m2_1_40# 0.247f
C91 m3_12600_1156# n7 0.181f
C92 via23_4_198/m2_1_40# via23_4_213/m2_1_40# 0.199f
C93 via23_4_331/m2_1_40# m3_11500_1156# 0.247f
C94 top m3_36200_1156# 0.187f
C95 via23_4_90/m2_1_40# n1 9.38e-20
C96 via23_4_200/m2_1_40# via23_4_198/m2_1_40# 0.199f
C97 top via23_4_702/m2_1_40# 0.341f
C98 via23_4_89/m2_1_40# m3_11300_1156# 0.123f
C99 via23_4_369/m2_1_40# m2_40200_1156# 0.251f
C100 m2_2100_1156# n3 5.59e-19
C101 m2_800_1156# n1 8.05e-20
C102 via23_4_20/m2_1_40# n7 1.18e-19
C103 n5 via23_4_96/m2_1_40# 2.03e-19
C104 m2_33700_1156# n5 1.13f
C105 via23_4_20/m2_1_40# n4 2.85e-19
C106 via23_4_446/m2_1_40# n6 0.452f
C107 via23_4_95/m2_1_40# n6 1.52e-19
C108 m2_16400_1156# n7 1.05e-19
C109 via23_4_94/m2_1_40# n1 9.38e-20
C110 m3_41200_1156# n6 4.08f
C111 n6 via23_4_103/m2_1_40# 1.52e-19
C112 n0 m2_9900_1156# 6.36e-20
C113 via23_4_704/m2_1_40# m3_42700_1156# 0.247f
C114 m3_33600_1156# m3_34700_1156# 0.148f
C115 m3_41400_1156# m3_42500_1156# 0.148f
C116 m2_16400_1156# n4 3.19e-19
C117 via23_4_89/m2_1_40# n1 9.38e-20
C118 top via23_4_117/m2_1_40# 0.216f
C119 top m3_25800_1156# 0.187f
C120 top via23_4_447/m2_1_40# 0.14f
C121 top m2_31100_1156# 0.267f
C122 m3_11300_1156# n5 0.993f
C123 via23_4_95/m2_1_40# n3 4.28e-19
C124 m3_33400_1156# n6 0.00746f
C125 m2_13800_1156# n7 3.52f
C126 m2_2100_1156# n0 6.36e-20
C127 m2_4700_1156# m3_5000_1156# 0.181f
C128 via23_4_94/m2_1_40# m3_4800_1156# 0.247f
C129 m2_24600_1156# n2 1.36e-19
C130 via23_4_334/m2_1_40# m3_16500_1156# 0.247f
C131 m3_33600_1156# n7 1.98f
C132 m2_13800_1156# n4 3.19e-19
C133 n3 via23_4_103/m2_1_40# 4.28e-19
C134 via23_4_326/m2_1_40# n5 0.452f
C135 via23_4_3/m2_1_40# n6 0.452f
C136 via23_4_21/m2_1_40# n1 9.38e-20
C137 top via23_4_641/m2_1_40# 0.216f
C138 m2_2100_1156# m3_2400_1156# 0.181f
C139 m2_36300_1156# m3_36200_1156# 2.11f
C140 n6 via23_4_380/m2_1_40# 0.512f
C141 m2_35000_1156# m3_36000_1156# 0.0061f
C142 n5 n1 0.0771f
C143 via23_4_368/m2_1_40# m3_38800_1156# 0.247f
C144 m2_6000_1156# n1 8.05e-20
C145 n3 n6 0.313f
C146 m2_25900_1156# n6 2.39f
C147 top m3_39900_1156# 0.187f
C148 n3 via23_4_3/m2_1_40# 4.28e-19
C149 m2_4700_1156# n7 3.52f
C150 via23_4_9/m2_1_40# n6 1.52e-19
C151 m2_11200_1156# n6 1.13f
C152 m3_17800_1156# m3_18000_1156# 3.35f
C153 m2_12500_1156# n5 2.05e-19
C154 m3_15400_1156# n5 4.08f
C155 m2_28500_1156# n7 2.42f
C156 m2_4700_1156# n4 3.19e-19
C157 via23_4_460/m2_1_40# n5 0.0714f
C158 via23_4_429/m2_1_40# m2_42800_1156# 0.251f
C159 m2_17700_1156# m3_18000_1156# 0.181f
C160 top m3_32100_1156# 0.187f
C161 via23_4_368/m2_1_40# m2_38900_1156# 0.251f
C162 m2_3400_1156# n6 2.39f
C163 top m3_8700_1156# 0.187f
C164 via23_4_455/m2_1_40# n5 1.57e-19
C165 m2_40200_1156# n7 1.13f
C166 n2 m3_12800_1156# 0.021f
C167 via23_4_635/m2_1_40# m2_42800_1156# 0.251f
C168 n3 m2_11200_1156# 5.59e-19
C169 n3 via23_4_9/m2_1_40# 4.28e-19
C170 n2 m3_2200_1156# 0.021f
C171 m3_42500_1156# n7 4.08f
C172 top via23_4_599/m2_1_40# 0.347f
C173 m2_9900_1156# m3_10200_1156# 0.181f
C174 m3_5000_1156# m3_6100_1156# 0.148f
C175 via23_4_710/m2_1_40# n7 0.452f
C176 via23_4_378/m2_1_40# m3_33600_1156# 0.247f
C177 top via23_4_347/m2_1_40# 0.347f
C178 n0 n6 0.0802f
C179 top m2_41500_1156# 0.267f
C180 m2_3400_1156# n3 5.59e-19
C181 via23_4_2/m2_1_40# n1 0.251f
C182 m2_27200_1156# m3_27100_1156# 2.11f
C183 m2_27200_1156# via23_4_448/m2_1_40# 0.251f
C184 top m2_9900_1156# 0.267f
C185 m3_18000_1156# n7 3.1f
C186 m2_33700_1156# via23_4_676/m2_1_40# 0.251f
C187 m3_24500_1156# n5 0.00889f
C188 m3_2400_1156# n6 4.08f
C189 n3 n0 1.36f
C190 m3_7400_1156# via23_4_87/m2_1_40# 0.247f
C191 n0 m2_11200_1156# 6.36e-20
C192 top m2_2100_1156# 0.267f
C193 m3_6100_1156# n7 1.98f
C194 m3_42500_1156# m3_42700_1156# 3.35f
C195 m3_34700_1156# m3_34900_1156# 3.35f
C196 via23_4_675/m2_1_40# top 0.347f
C197 ndum m2_9900_1156# 3.15e-20
C198 top m3_27100_1156# 0.187f
C199 m3_41400_1156# via23_4_712/m2_1_40# 0.247f
C200 top via23_4_448/m2_1_40# 0.14f
C201 via23_4_678/m2_1_40# m3_36200_1156# 0.123f
C202 via23_4_598/m2_1_40# m3_28200_1156# 0.247f
C203 m3_900_1156# n2 0.021f
C204 n2 via23_4_91/m2_1_40# 0.169f
C205 m2_15100_1156# n7 2.39f
C206 m2_3400_1156# n0 6.36e-20
C207 top via23_4_345/m2_1_40# 0.347f
C208 ndum m2_2100_1156# 3.15e-20
C209 via23_4_20/m2_1_40# n5 2.03e-19
C210 m3_34900_1156# n7 1.19f
C211 m2_15100_1156# n4 3.19e-19
C212 n2 m3_10000_1156# 0.021f
C213 via23_4_23/m2_1_40# n6 1.52e-19
C214 m2_3400_1156# m3_2400_1156# 0.0061f
C215 top via23_4_446/m2_1_40# 0.14f
C216 top via23_4_95/m2_1_40# 0.14f
C217 m2_16400_1156# n5 2.39f
C218 m3_8700_1156# via23_4_88/m2_1_40# 0.247f
C219 via23_4_22/m2_1_40# n6 1.52e-19
C220 m2_7300_1156# n1 8.05e-20
C221 m2_20300_1156# m3_19300_1156# 0.0061f
C222 m2_27200_1156# n6 1.13f
C223 top m3_41200_1156# 0.187f
C224 top via23_4_103/m2_1_40# 0.14f
C225 m2_13800_1156# via23_4_21/m2_1_40# 0.251f
C226 via23_4_94/m2_1_40# m2_4700_1156# 0.251f
C227 via23_4_23/m2_1_40# n3 4.28e-19
C228 m3_18000_1156# m3_19100_1156# 0.148f
C229 m2_13800_1156# n5 2.05e-19
C230 via23_4_449/m2_1_40# m3_29500_1156# 0.123f
C231 m2_29800_1156# n7 3.52f
C232 via23_4_677/m2_1_40# m2_35000_1156# 0.251f
C233 m3_33600_1156# n5 0.181f
C234 m2_19000_1156# m3_18000_1156# 0.0061f
C235 top m3_33400_1156# 0.187f
C236 n3 via23_4_22/m2_1_40# 4.28e-19
C237 via23_4_346/m2_1_40# n7 0.227f
C238 via23_4_589/m2_1_40# m2_24600_1156# 0.251f
C239 n2 m3_14100_1156# 0.021f
C240 top n6 16.4f
C241 n2 m3_3500_1156# 0.021f
C242 top via23_4_3/m2_1_40# 0.14f
C243 m3_25800_1156# m3_25600_1156# 3.35f
C244 m3_6100_1156# m3_6300_1156# 3.35f
C245 m2_11200_1156# m3_10200_1156# 0.0061f
C246 via23_4_712/m2_1_40# n7 0.452f
C247 via23_4_1/m2_1_40# n6 1.52e-19
C248 top via23_4_380/m2_1_40# 0.14f
C249 m3_42700_1156# via23_4_705/m2_1_40# 0.247f
C250 top via23_4_218/m2_1_40# 0.347f
C251 via23_4_381/m2_1_40# n7 0.452f
C252 top m2_42800_1156# 0.267f
C253 ndum n6 0.0782f
C254 m2_4700_1156# n5 2.05e-19
C255 top via23_4_429/m2_1_40# 0.216f
C256 top m2_25900_1156# 0.267f
C257 via23_4_379/m2_1_40# n7 0.452f
C258 m3_38600_1156# n7 4.08f
C259 top n3 2.35f
C260 m2_28500_1156# n5 1.14f
C261 top m2_11200_1156# 0.316f
C262 top via23_4_9/m2_1_40# 0.14f
C263 m2_42800_1156# via23_4_367/m2_1_40# 0.251f
C264 top m3_8900_1156# 0.187f
C265 n3 via23_4_1/m2_1_40# 4.28e-19
C266 via23_4_429/m2_1_40# via23_4_367/m2_1_40# 0.199f
C267 via23_4_635/m2_1_40# top 0.216f
C268 via23_4_229/m2_1_40# m3_2200_1156# 0.247f
C269 n2 via23_4_96/m2_1_40# 0.169f
C270 m3_19300_1156# n4 4.08f
C271 m3_30800_1156# n7 3.14f
C272 n2 via23_4_354/m2_1_40# 0.247f
C273 ndum n3 1.36f
C274 m3_7400_1156# n7 0.181f
C275 top m2_3400_1156# 0.267f
C276 m3_34900_1156# m3_36000_1156# 0.354f
C277 ndum m2_11200_1156# 3.15e-20
C278 via23_4_218/m2_1_40# m3_3700_1156# 0.247f
C279 top m3_28400_1156# 0.187f
C280 m3_3500_1156# via23_4_91/m2_1_40# 0.247f
C281 n2 m3_23200_1156# 3.4f
C282 m2_24600_1156# via23_4_460/m2_1_40# 0.251f
C283 via23_4_366/m2_1_40# m2_41500_1156# 0.251f
C284 top via23_4_128/m2_1_40# 0.216f
C285 m3_42700_1156# via23_4_419/m2_1_40# 0.247f
C286 ndum m2_3400_1156# 3.15e-20
C287 m3_36200_1156# n7 0.181f
C288 via23_4_346/m2_1_40# m3_19100_1156# 0.247f
C289 m3_29700_1156# m2_29800_1156# 2.11f
C290 top via23_4_111/m2_1_40# 0.216f
C291 top n0 0.418f
C292 m2_36300_1156# n6 0.637f
C293 n2 m3_11300_1156# 0.021f
C294 via23_4_710/m2_1_40# m3_38800_1156# 0.247f
C295 m2_19000_1156# via23_4_346/m2_1_40# 0.251f
C296 m2_36300_1156# via23_4_380/m2_1_40# 0.0256f
C297 m2_3400_1156# m3_3700_1156# 0.181f
C298 m3_37500_1156# via23_4_381/m2_1_40# 0.247f
C299 via23_4_588/m2_1_40# m3_23200_1156# 0.247f
C300 top via23_4_333/m2_1_40# 0.347f
C301 top m3_13900_1156# 0.187f
C302 ndum n0 13.4f
C303 top m3_2400_1156# 0.187f
C304 m3_900_1156# via23_4_96/m2_1_40# 0.247f
C305 m3_37500_1156# m3_38600_1156# 0.148f
C306 m3_900_1156# via23_4_198/m2_1_40# 0.247f
C307 via23_4_88/m2_1_40# n6 1.52e-19
C308 via23_4_710/m2_1_40# m2_38900_1156# 0.251f
C309 m2_6000_1156# m3_6100_1156# 2.11f
C310 m3_25800_1156# n7 0.181f
C311 m3_11500_1156# n6 4.08f
C312 m3_19100_1156# m3_19300_1156# 3.35f
C313 n2 n1 2.02f
C314 m2_15100_1156# n5 1.13f
C315 via23_4_447/m2_1_40# n7 0.452f
C316 via23_4_381/m2_1_40# m2_37600_1156# 0.251f
C317 m2_31100_1156# n7 1.13f
C318 m2_24600_1156# m3_24500_1156# 2.11f
C319 m2_12500_1156# m3_12800_1156# 0.181f
C320 m2_19000_1156# m3_19300_1156# 0.181f
C321 via23_4_333/m2_1_40# m3_15200_1156# 0.247f
C322 m3_41400_1156# m2_41500_1156# 2.11f
C323 m3_42700_1156# via23_4_702/m2_1_40# 0.247f
C324 m3_38600_1156# m2_37600_1156# 0.0061f
C325 m3_38600_1156# via23_4_709/m2_1_40# 0.247f
C326 n3 via23_4_88/m2_1_40# 4.28e-19
C327 m3_33600_1156# via23_4_676/m2_1_40# 0.247f
C328 m2_12500_1156# n2 0.00855f
C329 n2 m3_15400_1156# 0.021f
C330 via23_4_439/m2_1_40# m3_33400_1156# 0.247f
C331 m3_29700_1156# m3_30800_1156# 0.354f
C332 n2 m3_4800_1156# 0.021f
C333 m3_36000_1156# via23_4_379/m2_1_40# 0.247f
C334 m2_20300_1156# via23_4_347/m2_1_40# 0.251f
C335 top via23_4_23/m2_1_40# 0.14f
C336 m2_11200_1156# m3_11500_1156# 0.181f
C337 m3_6300_1156# m3_7400_1156# 0.148f
C338 via23_4_439/m2_1_40# n6 1.52e-19
C339 via23_4_334/m2_1_40# n5 0.452f
C340 via23_4_711/m2_1_40# m3_41200_1156# 0.247f
C341 n2 via23_4_455/m2_1_40# 0.352f
C342 top via23_4_22/m2_1_40# 0.14f
C343 top m2_27200_1156# 0.267f
C344 m3_39900_1156# n7 4.08f
C345 via23_4_91/m2_1_40# n1 9.38e-20
C346 m2_29800_1156# n5 0.002f
C347 m3_16500_1156# n6 0.181f
C348 top m3_10200_1156# 0.187f
C349 via23_4_678/m2_1_40# n6 0.452f
C350 via23_4_711/m2_1_40# n6 0.452f
C351 via23_4_369/m2_1_40# m3_41200_1156# 0.247f
C352 m3_8700_1156# n7 2.16f
C353 m3_36000_1156# m3_36200_1156# 3.35f
C354 via23_4_22/m2_1_40# m3_15200_1156# 0.247f
C355 via23_4_87/m2_1_40# n6 0.452f
C356 n2 m3_24500_1156# 3.16e-19
C357 m3_42700_1156# via23_4_641/m2_1_40# 0.247f
C358 via23_4_332/m2_1_40# m3_13900_1156# 0.247f
C359 m3_40100_1156# m2_40200_1156# 2.11f
C360 via23_4_599/m2_1_40# n7 0.227f
C361 m3_12800_1156# m3_12600_1156# 3.35f
C362 top via23_4_1/m2_1_40# 0.14f
C363 via23_4_447/m2_1_40# m3_29700_1156# 0.247f
C364 via23_4_345/m2_1_40# m3_17800_1156# 0.247f
C365 top via23_4_367/m2_1_40# 0.136f
C366 m3_41400_1156# m3_41200_1156# 3.35f
C367 via23_4_677/m2_1_40# m3_34900_1156# 0.123f
C368 m2_41500_1156# n7 2.39f
C369 n2 m3_12600_1156# 0.021f
C370 via23_4_345/m2_1_40# m2_17700_1156# 0.251f
C371 top ndum 0.414f
C372 via23_4_369/m2_1_40# n6 0.512f
C373 via23_4_347/m2_1_40# n4 0.452f
C374 n3 via23_4_87/m2_1_40# 4.28e-19
C375 m2_800_1156# via23_4_117/m2_1_40# 0.251f
C376 n2 via23_4_20/m2_1_40# 0.169f
C377 m2_9900_1156# n7 2.39f
C378 top m3_15200_1156# 0.187f
C379 m3_30800_1156# n5 0.00889f
C380 top m3_3700_1156# 0.187f
C381 m2_9900_1156# n4 3.19e-19
C382 m3_38600_1156# m3_38800_1156# 3.35f
C383 n2 m3_16700_1156# 0.021f
C384 m3_41400_1156# n6 0.181f
C385 m2_2100_1156# n7 2.39f
C386 via23_4_95/m2_1_40# m3_5000_1156# 0.247f
C387 m2_16400_1156# n2 0.00855f
C388 m3_19300_1156# m3_20400_1156# 0.148f
C389 m2_25900_1156# m3_25600_1156# 0.181f
C390 via23_4_448/m2_1_40# n7 1.18e-19
C391 m2_2100_1156# n4 3.19e-19
C392 m2_13800_1156# m3_12800_1156# 0.0061f
C393 m2_20300_1156# n6 1.43e-19
C394 m3_38600_1156# m2_38900_1156# 0.181f
C395 via23_4_251/m2_1_40# m3_10000_1156# 0.247f
C396 top m2_36300_1156# 0.316f
C397 m2_13800_1156# n2 0.00855f
C398 m3_30800_1156# m3_31000_1156# 3.35f
C399 m3_28200_1156# m2_28500_1156# 0.181f
C400 n6 m3_17800_1156# 1.98f
C401 via23_4_3/m2_1_40# m3_17800_1156# 0.247f
C402 m3_7400_1156# m3_7600_1156# 3.35f
C403 m3_8700_1156# m2_8600_1156# 2.11f
C404 m2_17700_1156# n6 2.39f
C405 n1 via23_4_96/m2_1_40# 9.38e-20
C406 top m3_24300_1156# 0.187f
C407 via23_4_446/m2_1_40# n7 1.18e-19
C408 m2_17700_1156# via23_4_3/m2_1_40# 0.251f
C409 via23_4_354/m2_1_40# n1 0.251f
C410 via23_4_95/m2_1_40# n7 0.452f
C411 m2_20300_1156# n3 1.09f
C412 top via23_4_245/m2_1_40# 0.347f
C413 via23_4_95/m2_1_40# n4 2.85e-19
C414 m3_41200_1156# n7 0.00642f
C415 m3_25800_1156# n5 0.00889f
C416 top via23_4_88/m2_1_40# 0.14f
C417 via23_4_458/m2_1_40# m3_25800_1156# 0.247f
C418 via23_4_326/m2_1_40# m3_11300_1156# 0.123f
C419 via23_4_103/m2_1_40# n7 0.452f
C420 via23_4_447/m2_1_40# n5 0.0714f
C421 top via23_4_332/m2_1_40# 0.347f
C422 m2_31100_1156# n5 0.002f
C423 top m3_11500_1156# 0.187f
C424 m3_34700_1156# n6 0.00746f
C425 m2_17700_1156# n3 5.59e-19
C426 via23_4_103/m2_1_40# n4 2.85e-19
C427 m2_4700_1156# n2 0.00855f
C428 via23_4_23/m2_1_40# m3_16500_1156# 0.247f
C429 m2_2100_1156# m3_1100_1156# 0.0061f
C430 m3_36200_1156# m3_37300_1156# 0.148f
C431 n6 n7 20.9f
C432 m2_9900_1156# via23_4_90/m2_1_40# 0.251f
C433 via23_4_3/m2_1_40# n7 1.18e-19
C434 m2_20300_1156# n0 1.98e-19
C435 n6 n4 0.318f
C436 via23_4_449/m2_1_40# m2_28500_1156# 0.251f
C437 top via23_4_439/m2_1_40# 0.14f
C438 via23_4_3/m2_1_40# n4 2.85e-19
C439 n7 via23_4_380/m2_1_40# 1.18e-19
C440 m3_31000_1156# m2_31100_1156# 2.11f
C441 via23_4_218/m2_1_40# n7 0.452f
C442 m2_42800_1156# n7 1.13f
C443 m2_25900_1156# n7 1.13f
C444 via23_4_590/m2_1_40# m3_26900_1156# 0.247f
C445 m2_17700_1156# n0 6.36e-20
C446 n3 n7 0.623f
C447 m2_11200_1156# n7 1.05e-19
C448 via23_4_9/m2_1_40# n7 0.227f
C449 top m3_16500_1156# 0.187f
C450 m3_8900_1156# n7 4.08f
C451 m3_32100_1156# n5 0.00889f
C452 n3 n4 10.8f
C453 m2_11200_1156# n4 3.19e-19
C454 via23_4_9/m2_1_40# n4 2.85e-19
C455 m3_38800_1156# m3_39900_1156# 0.148f
C456 via23_4_366/m2_1_40# top 0.14f
C457 top via23_4_678/m2_1_40# 0.347f
C458 top via23_4_711/m2_1_40# 0.347f
C459 m2_12500_1156# n1 8.05e-20
C460 n2 m3_18000_1156# 0.021f
C461 m2_23300_1156# n6 1.43e-19
C462 m3_1100_1156# via23_4_103/m2_1_40# 0.247f
C463 via23_4_584/m2_1_40# n2 0.247f
C464 m2_3400_1156# n7 1.13f
C465 m2_7300_1156# m3_7400_1156# 2.11f
C466 m3_28400_1156# n7 1.98f
C467 top via23_4_87/m2_1_40# 0.14f
C468 via23_4_589/m2_1_40# m3_24500_1156# 0.247f
C469 m2_3400_1156# n4 3.19e-19
C470 via23_4_455/m2_1_40# n1 0.251f
C471 m3_6100_1156# n2 0.021f
C472 via23_4_642/m2_1_40# via23_4_641/m2_1_40# 0.199f
C473 m2_13800_1156# m3_14100_1156# 0.181f
C474 m3_42700_1156# m2_42800_1156# 2.11f
C475 m3_39900_1156# m2_38900_1156# 0.0061f
C476 m3_37500_1156# n6 0.188f
C477 via23_4_429/m2_1_40# m3_42700_1156# 0.247f
C478 n0 n7 0.0951f
C479 m2_23300_1156# n3 1.09f
C480 m2_15100_1156# n2 0.00855f
C481 via23_4_378/m2_1_40# n6 0.0598f
C482 m3_25800_1156# m3_26900_1156# 0.148f
C483 m3_29500_1156# m2_28500_1156# 0.0061f
C484 m3_31000_1156# m3_32100_1156# 0.148f
C485 top via23_4_369/m2_1_40# 0.14f
C486 m2_9900_1156# n5 1.13f
C487 n0 n4 0.0773f
C488 m3_7600_1156# m3_8700_1156# 0.148f
C489 m2_19000_1156# n6 1.43e-19
C490 via23_4_635/m2_1_40# m3_42700_1156# 0.247f
C491 via23_4_333/m2_1_40# n7 0.452f
C492 top m3_25600_1156# 0.187f
C493 m3_13900_1156# n7 2.16f
C494 m2_8600_1156# n6 1.43e-19
C495 m3_6300_1156# n6 4.08f
C496 m3_20400_1156# via23_4_347/m2_1_40# 0.247f
C497 m2_37600_1156# n6 1.13f
C498 m2_2100_1156# n5 2.05e-19
C499 via23_4_675/m2_1_40# n5 0.452f
C500 n6 via23_4_90/m2_1_40# 1.52e-19
C501 m3_27100_1156# n5 1.99f
C502 via23_4_448/m2_1_40# n5 0.523f
C503 top m3_41400_1156# 0.187f
C504 via23_4_459/m2_1_40# n6 1.52e-19
C505 m2_800_1156# n6 1.43e-19
C506 via23_4_9/m2_1_40# m3_19100_1156# 0.247f
C507 m3_36000_1156# n6 0.00746f
C508 m2_19000_1156# n3 5.59e-19
C509 m2_33700_1156# m3_33600_1156# 2.11f
C510 m2_36300_1156# via23_4_678/m2_1_40# 0.0256f
C511 n3 m2_8600_1156# 5.59e-19
C512 m2_19000_1156# via23_4_9/m2_1_40# 0.251f
C513 m2_23300_1156# n0 6.79e-20
C514 m3_24500_1156# via23_4_460/m2_1_40# 0.247f
C515 top m2_20300_1156# 0.267f
C516 via23_4_199/m2_1_40# via23_4_111/m2_1_40# 0.199f
C517 m2_8600_1156# m3_8900_1156# 0.181f
C518 n3 via23_4_90/m2_1_40# 4.28e-19
C519 via23_4_94/m2_1_40# n6 1.52e-19
C520 via23_4_20/m2_1_40# n1 9.38e-20
C521 m2_20300_1156# via23_4_1/m2_1_40# 0.251f
C522 top m3_17800_1156# 0.187f
C523 m2_800_1156# n3 5.59e-19
C524 m3_8900_1156# via23_4_90/m2_1_40# 0.247f
C525 via23_4_446/m2_1_40# n5 0.0714f
C526 m2_12500_1156# m3_12600_1156# 2.11f
C527 m2_32400_1156# m3_32100_1156# 0.181f
C528 via23_4_95/m2_1_40# n5 2.03e-19
C529 via23_4_89/m2_1_40# n6 1.52e-19
C530 via23_4_23/m2_1_40# n7 1.18e-19
C531 ndum m2_20300_1156# 9.94e-20
C532 top m2_17700_1156# 0.267f
C533 via23_4_95/m2_1_40# m2_6000_1156# 0.251f
C534 top m3_5000_1156# 0.187f
C535 via23_4_23/m2_1_40# n4 2.85e-19
C536 via23_4_103/m2_1_40# n5 2.03e-19
C537 m2_12500_1156# via23_4_20/m2_1_40# 0.251f
C538 via23_4_22/m2_1_40# n7 0.452f
C539 m2_16400_1156# n1 8.05e-20
C540 m2_27200_1156# n7 1.05e-19
C541 via23_4_94/m2_1_40# n3 4.28e-19
C542 m2_19000_1156# n0 6.36e-20
C543 via23_4_22/m2_1_40# n4 2.85e-19
C544 ndum m2_17700_1156# 3.15e-20
C545 n0 m2_8600_1156# 6.36e-20
C546 via23_4_89/m2_1_40# n3 4.28e-19
C547 m3_7400_1156# via23_4_249/m2_1_40# 0.247f
C548 m3_33400_1156# n5 4.08f
C549 top m3_34700_1156# 0.187f
C550 m3_39900_1156# m3_40100_1156# 3.35f
C551 via23_4_89/m2_1_40# m2_11200_1156# 0.0256f
C552 m2_800_1156# via23_4_128/m2_1_40# 0.251f
C553 via23_4_21/m2_1_40# n6 1.52e-19
C554 m2_13800_1156# n1 8.05e-20
C555 m3_31000_1156# via23_4_446/m2_1_40# 0.247f
C556 m2_16400_1156# m3_15400_1156# 0.0061f
C557 n2 m3_19300_1156# 0.0214f
C558 via23_4_600/m2_1_40# m2_29800_1156# 0.251f
C559 n6 n5 16.1f
C560 m2_800_1156# n0 6.36e-20
C561 via23_4_458/m2_1_40# n6 0.452f
C562 m2_800_1156# via23_4_111/m2_1_40# 0.251f
C563 via23_4_3/m2_1_40# n5 2.03e-19
C564 m2_6000_1156# n6 1.13f
C565 top via23_4_228/m2_1_40# 0.276f
C566 top n7 32.8f
C567 m3_7400_1156# n2 0.021f
C568 m2_15100_1156# m3_14100_1156# 0.0061f
C569 top n4 4.11f
C570 n3 via23_4_21/m2_1_40# 4.28e-19
C571 via23_4_1/m2_1_40# n7 1.18e-19
C572 m3_38800_1156# n6 0.00746f
C573 via23_4_675/m2_1_40# m2_32400_1156# 0.251f
C574 m3_26900_1156# m3_27100_1156# 3.35f
C575 n3 n5 0.161f
C576 m2_25900_1156# n5 0.002f
C577 m3_32100_1156# m3_32300_1156# 3.35f
C578 m3_29500_1156# m2_29800_1156# 0.181f
C579 via23_4_1/m2_1_40# n4 0.453f
C580 ndum n7 0.177f
C581 via23_4_458/m2_1_40# m2_25900_1156# 0.251f
C582 via23_4_9/m2_1_40# n5 2.03e-19
C583 m2_11200_1156# n5 0.636f
C584 m2_6000_1156# n3 5.59e-19
C585 m2_4700_1156# n1 8.05e-20
C586 ndum n4 0.0771f
C587 m3_31000_1156# n6 1.98f
C588 m3_15200_1156# n7 1.98f
C589 m3_3700_1156# n7 4.08f
C590 m2_38900_1156# n6 0.00135f
C591 m2_3400_1156# n5 2.05e-19
C592 via23_4_20/m2_1_40# m3_12600_1156# 0.123f
C593 m3_28400_1156# n5 0.19f
C594 top m2_23300_1156# 0.267f
C595 n3 m3_20400_1156# 0.174f
C596 via23_4_230/m2_1_40# m3_3500_1156# 0.247f
C597 top m3_42700_1156# 0.187f
C598 via23_4_2/m2_1_40# n6 1.17e-19
C599 top via23_4_199/m2_1_40# 0.216f
C600 m2_4700_1156# m3_4800_1156# 2.11f
C601 via23_4_600/m2_1_40# m3_30800_1156# 0.123f
C602 m3_5000_1156# via23_4_245/m2_1_40# 0.247f
C603 m3_37300_1156# n6 4.09f
C604 m3_42700_1156# via23_4_367/m2_1_40# 0.247f
C605 n0 n5 0.0772f
C606 ndum m2_23300_1156# 1.34e-19
C607 m3_37300_1156# via23_4_380/m2_1_40# 0.247f
C608 via23_4_642/m2_1_40# m2_42800_1156# 0.251f
C609 top m3_37500_1156# 0.187f
C610 m2_6000_1156# n0 6.36e-20
C611 m2_36300_1156# n7 1.13f
C612 m3_13900_1156# via23_4_21/m2_1_40# 0.247f
C613 top m3_1100_1156# 0.187f
C614 top via23_4_378/m2_1_40# 0.14f
C615 top m3_19100_1156# 0.187f
C616 n3 via23_4_2/m2_1_40# 0.453f
C617 via23_4_675/m2_1_40# m3_32300_1156# 0.247f
C618 m2_32400_1156# m3_33400_1156# 0.0061f
C619 top m2_19000_1156# 0.267f
C620 via23_4_366/m2_1_40# m3_41400_1156# 0.247f
C621 m2_16400_1156# m3_16700_1156# 0.181f
C622 top m3_29700_1156# 0.187f
C623 via23_4_635/m2_1_40# via23_4_642/m2_1_40# 0.199f
C624 top m3_6300_1156# 0.187f
C625 top m2_8600_1156# 0.267f
C626 via23_4_584/m2_1_40# n1 0.251f
C627 n0 m3_20400_1156# 3.12e-19
C628 m2_32400_1156# n6 1.13f
C629 via23_4_245/m2_1_40# n7 0.452f
C630 m3_24300_1156# n4 4.08f
C631 m3_26900_1156# n6 4.08f
C632 top m2_37600_1156# 0.267f
C633 top via23_4_709/m2_1_40# 0.347f
C634 via23_4_88/m2_1_40# n7 0.452f
C635 top via23_4_90/m2_1_40# 0.14f
C636 top via23_4_459/m2_1_40# 0.14f
C637 via23_4_332/m2_1_40# n7 0.452f
C638 ndum m2_19000_1156# 3.15e-20
C639 top m2_800_1156# 0.267f
C640 ndum m2_8600_1156# 3.15e-20
C641 via23_4_88/m2_1_40# n4 2.85e-19
C642 top m3_36000_1156# 0.187f
C643 m3_900_1156# via23_4_117/m2_1_40# 0.247f
C644 m3_40100_1156# m3_41200_1156# 0.148f
C645 via23_4_89/m2_1_40# m3_10200_1156# 0.247f
C646 m2_15100_1156# n1 8.05e-20
C647 m2_25900_1156# m3_26900_1156# 0.0061f
C648 n0 via23_4_2/m2_1_40# 0.381f
C649 ndum m2_800_1156# 3.15e-20
C650 top via23_4_94/m2_1_40# 0.14f
C651 m2_7300_1156# n6 2.39f
C652 m3_8700_1156# n2 0.021f
C653 via23_4_23/m2_1_40# n5 0.452f
C654 m2_23300_1156# m3_24300_1156# 0.0061f
C655 m2_15100_1156# m3_15400_1156# 0.181f
C656 top via23_4_89/m2_1_40# 0.14f
C657 via23_4_439/m2_1_40# n7 1.18e-19
C658 via23_4_22/m2_1_40# n5 2.03e-19
C659 m3_40100_1156# n6 1.99f
C660 m3_27100_1156# m3_28200_1156# 0.148f
C661 m2_27200_1156# n5 2.39f
C662 via23_4_448/m2_1_40# m3_28200_1156# 0.247f
C663 m3_32300_1156# m3_33400_1156# 0.148f
C664 m3_10200_1156# n5 4.08f
C665 m2_31100_1156# via23_4_601/m2_1_40# 0.251f
C666 m2_7300_1156# n3 5.59e-19
C667 m3_32300_1156# n6 0.181f
C668 top via23_4_213/m2_1_40# 0.216f
C669 top via23_4_200/m2_1_40# 0.216f
C670 via23_4_331/m2_1_40# m2_12500_1156# 0.251f
C671 via23_4_94/m2_1_40# m3_3700_1156# 0.247f
C672 via23_4_334/m2_1_40# m3_15400_1156# 0.247f
C673 top via23_4_220/m2_1_40# 0.219f
C674 top via23_4_21/m2_1_40# 0.14f
C675 m2_9900_1156# n2 0.00855f
C676 via23_4_366/m2_1_40# n7 0.503f
C677 top via23_4_458/m2_1_40# 0.14f
C678 top n5 8.2f
C679 m2_36300_1156# m3_36000_1156# 0.181f
C680 m2_2100_1156# m3_2200_1156# 2.11f
C681 m2_35000_1156# m3_34900_1156# 2.11f
C682 via23_4_87/m2_1_40# n7 1.18e-19
C683 top m2_6000_1156# 0.267f
C684 m2_2100_1156# n2 0.00855f
C685 via23_4_1/m2_1_40# n5 2.03e-19
C686 via23_4_459/m2_1_40# m3_24300_1156# 0.247f
C687 via23_4_250/m2_1_40# m3_8700_1156# 0.247f
C688 m2_8600_1156# via23_4_88/m2_1_40# 0.251f
C689 via23_4_87/m2_1_40# n4 2.85e-19
C690 m2_24600_1156# n6 1.43e-19
C691 ndum n5 0.0767f
C692 top m3_38800_1156# 0.187f
C693 m2_7300_1156# n0 6.36e-20
C694 ndum m2_6000_1156# 3.15e-20
C695 top m3_20400_1156# 0.187f
C696 via23_4_369/m2_1_40# n7 1.18e-19
C697 m3_15200_1156# n5 0.181f
C698 via23_4_1/m2_1_40# m3_20400_1156# 0.247f
C699 m2_17700_1156# m3_17800_1156# 2.11f
C700 m3_25600_1156# n7 4.08f
C701 top m3_31000_1156# 0.187f
C702 m3_32100_1156# via23_4_601/m2_1_40# 0.247f
C703 top m3_7600_1156# 0.187f
C704 top m2_38900_1156# 0.267f
C705 ndum m3_20400_1156# 1.58e-19
C706 via23_4_95/m2_1_40# n2 0.169f
C707 via23_4_599/m2_1_40# m3_29500_1156# 0.123f
C708 m3_41400_1156# n7 1.99f
C709 m3_2200_1156# via23_4_103/m2_1_40# 0.247f
C710 top via23_4_2/m2_1_40# 0.14f
C711 top via23_4_642/m2_1_40# 0.216f
C712 m2_9900_1156# m3_10000_1156# 2.11f
C713 via23_4_331/m2_1_40# m3_12600_1156# 0.123f
C714 top m3_37300_1156# 0.187f
C715 n2 via23_4_103/m2_1_40# 0.169f
C716 via23_4_704/m2_1_40# via23_4_705/m2_1_40# 0.199f
C717 via23_4_249/m2_1_40# n6 0.452f
C718 m2_20300_1156# n7 1.05e-19
C719 m2_27200_1156# m3_26900_1156# 0.181f
C720 via23_4_414/m2_1_40# via23_4_419/m2_1_40# 0.199f
C721 m2_20300_1156# n4 2.39f
C722 m3_17800_1156# n7 0.181f
C723 m3_24300_1156# n5 0.00889f
C724 m3_2200_1156# n6 0.181f
C725 top via23_4_677/m2_1_40# 0.347f
C726 n2 n6 0.39f
C727 m2_17700_1156# n7 1.13f
C728 m2_35000_1156# via23_4_379/m2_1_40# 0.251f
C729 m3_6300_1156# via23_4_87/m2_1_40# 0.247f
C730 n2 via23_4_3/m2_1_40# 0.169f
C731 m3_28200_1156# m3_28400_1156# 3.35f
C732 m3_5000_1156# n7 4.08f
C733 via23_4_334/m2_1_40# m2_16400_1156# 0.251f
C734 via23_4_88/m2_1_40# n5 2.03e-19
C735 m2_17700_1156# n4 3.19e-19
C736 m2_6000_1156# via23_4_245/m2_1_40# 0.251f
C737 top m3_26900_1156# 0.187f
C738 top m2_32400_1156# 0.267f
C739 via23_4_598/m2_1_40# m3_27100_1156# 0.247f
C740 via23_4_449/m2_1_40# n6 1.52e-19
C741 n3 n2 19.4f
C742 m3_34700_1156# n7 4.08f
C743 m2_11200_1156# n2 0.00855f
C744 via23_4_9/m2_1_40# n2 0.169f
C745 n2 m3_8900_1156# 0.021f
C746 m2_36300_1156# m3_37300_1156# 0.0061f
C747 top m2_7300_1156# 0.267f
C748 m2_3400_1156# n2 0.00855f
C749 via23_4_439/m2_1_40# n5 0.523f
C750 top via23_4_676/m2_1_40# 0.347f
C751 via23_4_91/m2_1_40# n6 0.452f
C752 m3_7600_1156# via23_4_88/m2_1_40# 0.247f
C753 via23_4_368/m2_1_40# m3_39900_1156# 0.247f
C754 n7 n4 0.678f
C755 top m3_40100_1156# 0.187f
C756 ndum m2_7300_1156# 3.15e-20
C757 via23_4_449/m2_1_40# m3_28400_1156# 0.247f
C758 m3_16500_1156# n5 1.98f
C759 n0 n2 1.42f
C760 via23_4_704/m2_1_40# via23_4_702/m2_1_40# 0.199f
C761 n3 via23_4_91/m2_1_40# 4.28e-19
C762 top m3_32300_1156# 0.187f
C763 m3_12800_1156# m3_13900_1156# 0.148f
C764 via23_4_229/m2_1_40# m2_2100_1156# 0.251f
C765 m3_2200_1156# m3_2400_1156# 3.35f
C766 n2 m3_13900_1156# 0.021f
C767 n6 via23_4_601/m2_1_40# 0.452f
C768 m2_23300_1156# n7 1.05e-19
C769 n2 m3_2400_1156# 0.021f
C770 via23_4_87/m2_1_40# n5 2.03e-19
C771 m3_42700_1156# n7 0.181f
C772 m2_3400_1156# via23_4_91/m2_1_40# 0.251f
C773 via23_4_378/m2_1_40# m3_34700_1156# 0.247f
C774 m3_8900_1156# m3_10000_1156# 0.148f
C775 m2_23300_1156# n4 2.39f
C776 m2_27200_1156# m3_28200_1156# 0.0061f
C777 via23_4_128/m2_1_40# m3_900_1156# 0.247f
C778 top m2_24600_1156# 0.267f
C779 m3_37500_1156# n7 1.98f
C780 m3_1100_1156# n7 4.08f
C781 via23_4_378/m2_1_40# n7 0.452f
C782 m3_900_1156# via23_4_111/m2_1_40# 0.247f
C783 m3_19100_1156# n7 1.98f
C784 m3_3500_1156# n6 1.98f
C785 m3_25600_1156# n5 0.00889f
C786 m2_9900_1156# n1 8.05e-20
C787 m3_19100_1156# n4 0.181f
C788 m2_19000_1156# n7 2.42f
C789 m3_29700_1156# n7 2.16f
C790 m2_8600_1156# n7 3.52f
C791 m3_28400_1156# m3_29500_1156# 0.148f
C792 via23_4_23/m2_1_40# n2 0.169f
C793 m2_19000_1156# n4 1.13f
C794 top m3_28200_1156# 0.187f
C795 m2_37600_1156# n7 2.39f
C796 m3_42500_1156# via23_4_712/m2_1_40# 0.247f
C797 m3_2400_1156# via23_4_91/m2_1_40# 0.247f
C798 via23_4_678/m2_1_40# m3_37300_1156# 0.247f
C799 via23_4_709/m2_1_40# n7 0.452f
C800 m2_8600_1156# n4 3.19e-19
C801 via23_4_90/m2_1_40# n7 0.452f
C802 m2_2100_1156# n1 8.05e-20
C803 via23_4_459/m2_1_40# n7 1.18e-19
C804 m2_33700_1156# m3_33400_1156# 0.181f
C805 n2 via23_4_22/m2_1_40# 0.169f
C806 via23_4_439/m2_1_40# m2_32400_1156# 0.251f
C807 via23_4_228/m2_1_40# m2_800_1156# 0.251f
C808 m2_800_1156# n7 1.13f
C809 via23_4_90/m2_1_40# n4 2.85e-19
C810 via23_4_346/m2_1_40# m3_18000_1156# 0.123f
C811 m3_36000_1156# n7 4.08f
C812 via23_4_459/m2_1_40# n4 0.541f
C813 m2_20300_1156# n5 2.05e-19
C814 m2_800_1156# n4 3.19e-19
C815 m2_33700_1156# n6 0.00135f
C816 n2 m3_10200_1156# 0.021f
C817 n6 via23_4_96/m2_1_40# 1.52e-19
C818 top via23_4_249/m2_1_40# 0.347f
C819 m2_3400_1156# m3_3500_1156# 2.11f
C820 via23_4_94/m2_1_40# n7 0.452f
C821 top m3_12800_1156# 0.187f
C822 m2_17700_1156# n5 2.05e-19
C823 top m3_2200_1156# 0.187f
C824 via23_4_94/m2_1_40# n4 2.85e-19
C825 via23_4_89/m2_1_40# n7 1.18e-19
C826 m2_20300_1156# m3_20400_1156# 2.11f
C827 top n2 1.32f
C828 n3 via23_4_96/m2_1_40# 4.28e-19
C829 via23_4_95/m2_1_40# n1 9.38e-20
C830 via23_4_89/m2_1_40# n4 2.85e-19
C831 m2_6000_1156# m3_5000_1156# 0.0061f
C832 n3 via23_4_354/m2_1_40# 0.452f
C833 m2_23300_1156# via23_4_459/m2_1_40# 0.251f
C834 n2 via23_4_1/m2_1_40# 0.169f
C835 m3_11300_1156# n6 0.181f
C836 m2_24600_1156# m3_24300_1156# 0.181f
C837 via23_4_103/m2_1_40# n1 9.38e-20
C838 n3 m3_23200_1156# 0.174f
C839 top via23_4_449/m2_1_40# 0.14f
C840 m2_800_1156# via23_4_199/m2_1_40# 0.251f
C841 via23_4_333/m2_1_40# m3_14100_1156# 0.247f
C842 m2_19000_1156# m3_19100_1156# 2.11f
C843 ndum n2 1.42f
C844 m3_13900_1156# m3_14100_1156# 3.35f
C845 m3_37500_1156# m2_37600_1156# 2.11f
C846 via23_4_251/m2_1_40# m2_9900_1156# 0.251f
C847 m3_37500_1156# via23_4_709/m2_1_40# 0.247f
C848 via23_4_368/m2_1_40# n6 0.0598f
C849 via23_4_228/m2_1_40# via23_4_220/m2_1_40# 0.199f
C850 via23_4_21/m2_1_40# n7 0.452f
C851 m3_2400_1156# m3_3500_1156# 0.148f
C852 n2 m3_15200_1156# 0.021f
C853 via23_4_439/m2_1_40# m3_32300_1156# 0.247f
C854 top via23_4_588/m2_1_40# 0.347f
C855 n2 m3_3700_1156# 0.021f
C856 n7 n5 1.06f
C857 via23_4_21/m2_1_40# n4 2.85e-19
C858 via23_4_458/m2_1_40# n7 1.18e-19
C859 m3_34900_1156# via23_4_379/m2_1_40# 0.123f
C860 via23_4_128/m2_1_40# via23_4_96/m2_1_40# 0.199f
C861 m2_800_1156# m3_1100_1156# 0.181f
C862 m2_11200_1156# m3_11300_1156# 2.11f
C863 m3_10000_1156# m3_10200_1156# 3.35f
C864 n6 n1 0.0843f
C865 m2_7300_1156# via23_4_87/m2_1_40# 0.251f
C866 via23_4_711/m2_1_40# m3_40100_1156# 0.247f
C867 n4 n5 11.4f
C868 m2_6000_1156# n7 2.39f
C869 via23_4_3/m2_1_40# n1 9.38e-20
C870 top m3_900_1156# 0.187f
C871 top via23_4_91/m2_1_40# 0.14f
C872 m2_37600_1156# via23_4_709/m2_1_40# 0.251f
C873 n0 via23_4_354/m2_1_40# 0.247f
C874 top via23_4_600/m2_1_40# 0.347f
C875 m2_6000_1156# n4 3.19e-19
C876 via23_4_326/m2_1_40# m2_11200_1156# 0.0256f
C877 top via23_4_250/m2_1_40# 0.347f
C878 m3_38800_1156# n7 2.16f
C879 n0 m3_23200_1156# 1.58e-19
C880 m2_27200_1156# via23_4_598/m2_1_40# 0.251f
C881 m2_12500_1156# n6 2.39f
C882 via23_4_460/m2_1_40# n6 1.52e-19
C883 top m3_10000_1156# 0.187f
C884 n3 n1 3.36f
C885 via23_4_200/m2_1_40# via23_4_199/m2_1_40# 0.199f
C886 m2_11200_1156# n1 8.05e-20
C887 via23_4_9/m2_1_40# n1 9.38e-20
C888 m3_20400_1156# n4 1.98f
C889 m3_31000_1156# n7 0.181f
C890 via23_4_455/m2_1_40# n6 1.17e-19
C891 via23_4_369/m2_1_40# m3_40100_1156# 0.247f
C892 m3_7600_1156# n7 4.08f
C893 m2_23300_1156# n5 2.05e-19
C894 via23_4_22/m2_1_40# m3_14100_1156# 0.247f
C895 via23_4_218/m2_1_40# m3_4800_1156# 0.247f
C896 top m3_29500_1156# 0.187f
C897 m2_38900_1156# n7 3.52f
C898 n2 m3_24300_1156# 4.18e-19
C899 m2_12500_1156# n3 5.59e-19
C900 top via23_4_601/m2_1_40# 0.347f
C901 m2_3400_1156# n1 8.05e-20
C902 via23_4_332/m2_1_40# m3_12800_1156# 0.247f
C903 top via23_4_598/m2_1_40# 0.347f
C904 m3_39900_1156# m2_40200_1156# 0.181f
C905 via23_4_2/m2_1_40# n7 9.11e-20
C906 via23_4_345/m2_1_40# m3_16700_1156# 0.123f
C907 m3_30800_1156# m2_29800_1156# 0.023f
C908 n2 via23_4_88/m2_1_40# 0.169f
C909 n3 via23_4_455/m2_1_40# 0.453f
C910 m2_35000_1156# n6 0.00135f
C911 via23_4_2/m2_1_40# n4 2.21e-19
C912 n2 m3_11500_1156# 0.021f
C913 via23_4_710/m2_1_40# m3_39900_1156# 0.247f
C914 m2_42800_1156# via23_4_414/m2_1_40# 0.251f
C915 via23_4_429/m2_1_40# via23_4_414/m2_1_40# 0.199f
C916 n0 n1 13.4f
C917 m3_38600_1156# via23_4_381/m2_1_40# 0.247f
C918 via23_4_588/m2_1_40# m3_24300_1156# 0.247f
C919 top m3_14100_1156# 0.187f
C920 via23_4_599/m2_1_40# m2_28500_1156# 0.251f
C921 m2_19000_1156# n5 2.05e-19
C922 top m3_3500_1156# 0.187f
C923 m3_29700_1156# n5 0.00889f
C924 via23_4_677/m2_1_40# n7 0.452f
C925 m2_8600_1156# n5 2.05e-19
C926 m2_800_1156# via23_4_213/m2_1_40# 0.251f
C927 m2_800_1156# via23_4_200/m2_1_40# 0.251f
C928 m2_12500_1156# n0 6.36e-20
C929 m2_800_1156# via23_4_220/m2_1_40# 0.251f
C930 m2_6000_1156# m3_6300_1156# 0.181f
C931 via23_4_90/m2_1_40# n5 2.03e-19
C932 m2_32400_1156# n7 1.05e-19
C933 m3_12600_1156# n6 1.01f
C934 via23_4_459/m2_1_40# n5 2.03e-19
C935 via23_4_642/m2_1_40# m3_42700_1156# 0.247f
C936 m2_24600_1156# m3_25600_1156# 0.0061f
C937 m2_800_1156# n5 2.05e-19
C938 via23_4_704/m2_1_40# m2_42800_1156# 0.251f
C939 via23_4_20/m2_1_40# n6 0.452f
C940 m3_42500_1156# m2_41500_1156# 0.0061f
C941 m3_14100_1156# m3_15200_1156# 0.148f
C942 via23_4_251/m2_1_40# m3_8900_1156# 0.247f
C943 m3_3500_1156# m3_3700_1156# 3.35f
C944 m3_34700_1156# via23_4_676/m2_1_40# 0.247f
C945 n2 m3_16500_1156# 0.021f
C946 top m2_33700_1156# 0.267f
C947 top via23_4_96/m2_1_40# 0.136f
C948 n6 m3_16700_1156# 3.14f
C949 top via23_4_229/m2_1_40# 0.347f
C950 top via23_4_354/m2_1_40# 0.347f
C951 via23_4_94/m2_1_40# n5 2.03e-19
C952 via23_4_447/m2_1_40# m2_29800_1156# 0.251f
C953 top via23_4_198/m2_1_40# 0.216f
C954 m3_37500_1156# m3_37300_1156# 3.35f
C955 via23_4_3/m2_1_40# m3_16700_1156# 0.123f
C956 m3_7600_1156# m2_8600_1156# 0.0061f
C957 m3_10200_1156# m3_11300_1156# 0.148f
C958 m2_16400_1156# n6 1.13f
C959 top m3_23200_1156# 0.187f
C960 via23_4_89/m2_1_40# n5 0.452f
C961 n3 via23_4_20/m2_1_40# 4.28e-19
C962 m2_7300_1156# n7 1.13f
C963 via23_4_676/m2_1_40# n7 0.452f
C964 via23_4_23/m2_1_40# n1 9.38e-20
C965 m2_7300_1156# n4 3.19e-19
C966 n2 via23_4_87/m2_1_40# 0.169f
C967 m3_33600_1156# m3_33400_1156# 3.35f
C968 via23_4_220/m2_1_40# via23_4_213/m2_1_40# 0.199f
C969 top via23_4_589/m2_1_40# 0.347f
C970 m3_40100_1156# n7 0.181f
C971 via23_4_326/m2_1_40# m3_10200_1156# 0.247f
C972 m2_13800_1156# n6 1.43e-19
C973 via23_4_22/m2_1_40# n1 9.38e-20
C974 ndum m3_23200_1156# 3.12e-19
C975 m2_37600_1156# m3_37300_1156# 0.181f
C976 top m3_11300_1156# 0.187f
C977 m3_33600_1156# n6 0.00746f
C978 m2_16400_1156# n3 5.59e-19
C979 via23_4_23/m2_1_40# m3_15400_1156# 0.247f
C980 via23_4_21/m2_1_40# n5 2.03e-19
C981 top via23_4_326/m2_1_40# 0.347f
C982 top via23_4_368/m2_1_40# 0.14f
C983 via23_4_458/m2_1_40# n5 0.0714f
C984 m2_13800_1156# n3 5.59e-19
C985 m2_6000_1156# n5 2.05e-19
C986 m3_41200_1156# m2_40200_1156# 0.0061f
C987 via23_4_447/m2_1_40# m3_30800_1156# 0.123f
C988 m3_30800_1156# m2_31100_1156# 0.181f
C989 top n1 0.983f
C990 via23_4_641/m2_1_40# via23_4_419/m2_1_40# 0.199f
C991 m2_4700_1156# n6 1.43e-19
C992 via23_4_677/m2_1_40# m3_36000_1156# 0.247f
C993 via23_4_1/m2_1_40# n1 9.38e-20
C994 n6 m2_28500_1156# 1.43e-19
C995 via23_4_590/m2_1_40# m3_25800_1156# 0.247f
C996 m2_16400_1156# n0 6.36e-20
C997 m2_24600_1156# n7 2.39f
C998 top m2_12500_1156# 0.267f
C999 m2_4700_1156# via23_4_218/m2_1_40# 0.251f
C1000 top m3_15400_1156# 0.187f
C1001 ndum n1 3.54f
C1002 m2_24600_1156# n4 1.13f
C1003 top via23_4_460/m2_1_40# 0.14f
C1004 m2_20300_1156# n2 0.256f
C1005 m3_31000_1156# n5 0.00889f
C1006 top m3_4800_1156# 0.187f
C1007 m2_40200_1156# n6 2.39f
C1008 m2_4700_1156# n3 5.59e-19
C1009 m3_23200_1156# m3_24300_1156# 0.148f
C1010 n2 m3_17800_1156# 0.021f
C1011 top via23_4_455/m2_1_40# 0.14f
C1012 m2_13800_1156# n0 6.36e-20
C1013 m2_7300_1156# m3_6300_1156# 0.0061f
C1014 ndum m2_12500_1156# 3.15e-20
C1015 via23_4_95/m2_1_40# m3_6100_1156# 0.247f
C1016 m2_17700_1156# n2 0.00855f
C1017 via23_4_2/m2_1_40# n5 1.57e-19
C1018 m3_5000_1156# n2 0.021f
C1019 top via23_4_414/m2_1_40# 0.216f
C1020 m3_42500_1156# m2_42800_1156# 0.181f
C1021 m2_13800_1156# m3_13900_1156# 2.11f
C1022 m3_15200_1156# m3_15400_1156# 3.35f
C1023 m3_38800_1156# m2_38900_1156# 2.11f
C1024 ndum via23_4_455/m2_1_40# 0.381f
C1025 m2_41500_1156# via23_4_712/m2_1_40# 0.251f
C1026 m3_3700_1156# m3_4800_1156# 0.148f
C1027 top m2_35000_1156# 0.267f
C1028 m3_28400_1156# m2_28500_1156# 2.11f
C1029 m3_11300_1156# m3_11500_1156# 3.35f
C1030 top m3_24500_1156# 0.187f
C1031 m2_4700_1156# n0 6.36e-20
C1032 m3_12800_1156# n7 4.08f
C1033 m3_6100_1156# n6 0.181f
C1034 m3_2200_1156# n7 1.98f
C1035 m3_19300_1156# via23_4_347/m2_1_40# 0.247f
C1036 via23_4_23/m2_1_40# m2_16400_1156# 0.251f
C1037 top via23_4_251/m2_1_40# 0.347f
C1038 n2 n7 0.78f
C1039 m2_32400_1156# n5 2.39f
C1040 m3_26900_1156# n5 0.00889f
C1041 via23_4_458/m2_1_40# m3_26900_1156# 0.247f
C1042 top via23_4_704/m2_1_40# 0.222f
C1043 m2_15100_1156# n6 1.43e-19
C1044 via23_4_584/m2_1_40# n3 0.452f
C1045 n2 n4 0.144f
C1046 via23_4_9/m2_1_40# m3_18000_1156# 0.123f
C1047 top m3_12600_1156# 0.221f
C1048 m3_34900_1156# n6 0.00746f
C1049 via23_4_88/m2_1_40# n1 9.38e-20
C1050 via23_4_449/m2_1_40# n7 0.227f
C1051 top via23_4_20/m2_1_40# 0.14f
C1052 m2_15100_1156# n3 5.59e-19
C1053 top m3_16700_1156# 0.221f
C1054 via23_4_331/m2_1_40# n6 0.452f
C1055 m2_7300_1156# n5 2.05e-19
C1056 via23_4_588/m2_1_40# n4 0.452f
C1057 m2_12500_1156# m3_11500_1156# 0.0061f
C1058 top m2_16400_1156# 0.267f
C1059 m2_23300_1156# n2 0.247f
C1060 via23_4_230/m2_1_40# n6 0.452f
C1061 m3_32100_1156# m2_31100_1156# 0.0061f
C1062 m3_900_1156# n7 0.181f
C1063 via23_4_228/m2_1_40# m3_900_1156# 0.247f
C1064 via23_4_91/m2_1_40# n7 1.18e-19
C1065 via23_4_600/m2_1_40# n7 0.452f
C1066 n6 m2_29800_1156# 1.43e-19
C1067 via23_4_250/m2_1_40# n7 0.452f
C1068 via23_4_91/m2_1_40# n4 2.85e-19
C1069 m2_42800_1156# via23_4_705/m2_1_40# 0.251f
C1070 ndum m2_16400_1156# 3.15e-20
C1071 top m2_13800_1156# 0.267f
C1072 m3_1100_1156# m3_2200_1156# 0.148f
C1073 m3_10000_1156# n7 1.98f
C1074 m3_6300_1156# via23_4_249/m2_1_40# 0.247f
C1075 m3_32300_1156# n5 1.99f
C1076 top m3_33600_1156# 0.187f
C1077 n2 m3_1100_1156# 0.021f
C1078 m3_24300_1156# m3_24500_1156# 3.35f
C1079 n2 m3_19100_1156# 0.0213f
C1080 via23_4_588/m2_1_40# m2_23300_1156# 0.251f
C1081 m2_15100_1156# n0 6.36e-20
C1082 m2_7300_1156# m3_7600_1156# 0.181f
C1083 ndum m2_13800_1156# 3.15e-20
C1084 via23_4_635/m2_1_40# via23_4_705/m2_1_40# 0.199f
C1085 m2_19000_1156# n2 0.00869f
C1086 m3_29500_1156# n7 3.1f
C1087 via23_4_589/m2_1_40# m3_25600_1156# 0.247f
C1088 m2_8600_1156# n2 0.00855f
C1089 m3_6300_1156# n2 0.021f
C1090 via23_4_381/m2_1_40# n6 0.0598f
C1091 via23_4_230/m2_1_40# m2_3400_1156# 0.251f
C1092 via23_4_333/m2_1_40# m2_15100_1156# 0.251f
C1093 m3_15400_1156# m3_16500_1156# 0.148f
C1094 via23_4_87/m2_1_40# n1 9.38e-20
C1095 m3_38600_1156# n6 0.00746f
C1096 n2 via23_4_90/m2_1_40# 0.169f
C1097 via23_4_379/m2_1_40# n6 0.0598f
C1098 m3_900_1156# via23_4_199/m2_1_40# 0.247f
C1099 top m2_4700_1156# 0.267f
C1100 m2_24600_1156# n5 0.002f
C1101 m2_800_1156# n2 0.00855f
C1102 m2_42800_1156# via23_4_419/m2_1_40# 0.251f
C1103 top m2_28500_1156# 0.267f
C1104 m3_11500_1156# m3_12600_1156# 0.354f
C1105 m3_14100_1156# n7 4.08f
C1106 m3_900_1156# m3_1100_1156# 3.35f
C1107 m3_7400_1156# n6 1.98f
C1108 ndum m2_4700_1156# 3.15e-20
C1109 m3_3500_1156# n7 0.181f
C1110 top m2_40200_1156# 0.267f
C1111 via23_4_20/m2_1_40# m3_11500_1156# 0.247f
C1112 via23_4_94/m2_1_40# n2 0.169f
C1113 m3_28200_1156# n5 4.09f
C1114 via23_4_230/m2_1_40# m3_2400_1156# 0.247f
C1115 via23_4_590/m2_1_40# n6 0.452f
C1116 top m3_42500_1156# 0.187f
C1117 via23_4_89/m2_1_40# n2 0.169f
C1118 top via23_4_710/m2_1_40# 0.347f
C1119 m2_4700_1156# m3_3700_1156# 0.0061f
C1120 via23_4_600/m2_1_40# m3_29700_1156# 0.247f
C1121 via23_4_446/m2_1_40# m2_31100_1156# 0.251f
C1122 m2_33700_1156# m3_34700_1156# 0.0061f
C1123 m3_36200_1156# n6 1f
C1124 via23_4_250/m2_1_40# m2_8600_1156# 0.251f
C1125 m3_25600_1156# via23_4_460/m2_1_40# 0.247f
C1126 m3_36200_1156# via23_4_380/m2_1_40# 0.123f
C1127 m2_15100_1156# via23_4_22/m2_1_40# 0.251f
C1128 m2_800_1156# m3_900_1156# 2.11f
C1129 m3_12800_1156# via23_4_21/m2_1_40# 0.247f
C1130 via23_4_590/m2_1_40# m2_25900_1156# 0.251f
C1131 m2_33700_1156# n7 2.39f
C1132 n7 via23_4_96/m2_1_40# 1.18e-19
C1133 top m3_18000_1156# 0.187f
C1134 m2_42800_1156# via23_4_702/m2_1_40# 0.251f
C1135 m2_20300_1156# n1 8.05e-20
C1136 m2_13800_1156# via23_4_332/m2_1_40# 0.251f
C1137 m3_10000_1156# via23_4_90/m2_1_40# 0.247f
C1138 via23_4_229/m2_1_40# n7 0.452f
C1139 top via23_4_584/m2_1_40# 0.347f
C1140 m3_29700_1156# m3_29500_1156# 3.35f
C1141 n2 via23_4_21/m2_1_40# 0.169f
C1142 m2_32400_1156# m3_32300_1156# 2.11f
C1143 n4 via23_4_96/m2_1_40# 2.85e-19
C1144 n2 n5 0.196f
C1145 top m3_6100_1156# 0.187f
C1146 m3_23200_1156# n4 1.99f
C1147 m3_25800_1156# n6 1.98f
C1148 m2_6000_1156# n2 0.00855f
C1149 m2_17700_1156# n1 8.05e-20
C1150 via23_4_447/m2_1_40# n6 1.52e-19
C1151 n1 VSUBS 3.76f
C1152 n5 VSUBS 16.9f
C1153 n4 VSUBS 8.19f
C1154 n3 VSUBS 5.86f
C1155 via23_4_200/m2_1_40# VSUBS 0.372f
C1156 via23_4_414/m2_1_40# VSUBS 0.372f
C1157 via23_4_447/m2_1_40# VSUBS 0.291f
C1158 via23_4_458/m2_1_40# VSUBS 0.291f
C1159 via23_4_446/m2_1_40# VSUBS 0.291f
C1160 via23_4_460/m2_1_40# VSUBS 0.291f
C1161 via23_4_220/m2_1_40# VSUBS 0.372f
C1162 via23_4_9/m2_1_40# VSUBS 0.364f
C1163 via23_4_459/m2_1_40# VSUBS 0.28f
C1164 via23_4_641/m2_1_40# VSUBS 0.372f
C1165 via23_4_455/m2_1_40# VSUBS 0.243f
C1166 via23_4_635/m2_1_40# VSUBS 0.372f
C1167 via23_4_601/m2_1_40# VSUBS 0.373f
C1168 via23_4_676/m2_1_40# VSUBS 0.373f
C1169 n0 VSUBS 2.8f
C1170 via23_4_3/m2_1_40# VSUBS 0.253f
C1171 via23_4_642/m2_1_40# VSUBS 0.372f
C1172 via23_4_709/m2_1_40# VSUBS 0.373f
C1173 via23_4_678/m2_1_40# VSUBS 0.485f
C1174 via23_4_117/m2_1_40# VSUBS 0.372f
C1175 via23_4_128/m2_1_40# VSUBS 0.372f
C1176 via23_4_677/m2_1_40# VSUBS 0.373f
C1177 via23_4_21/m2_1_40# VSUBS 0.253f
C1178 via23_4_103/m2_1_40# VSUBS 0.253f
C1179 via23_4_20/m2_1_40# VSUBS 0.253f
C1180 via23_4_91/m2_1_40# VSUBS 0.253f
C1181 via23_4_326/m2_1_40# VSUBS 0.485f
C1182 via23_4_111/m2_1_40# VSUBS 0.372f
C1183 via23_4_198/m2_1_40# VSUBS 0.372f
C1184 via23_4_379/m2_1_40# VSUBS 0.3f
C1185 via23_4_346/m2_1_40# VSUBS 0.485f
C1186 via23_4_1/m2_1_40# VSUBS 0.253f
C1187 via23_4_712/m2_1_40# VSUBS 0.373f
C1188 via23_4_199/m2_1_40# VSUBS 0.372f
C1189 via23_4_378/m2_1_40# VSUBS 0.3f
C1190 via23_4_334/m2_1_40# VSUBS 0.373f
C1191 via23_4_345/m2_1_40# VSUBS 0.373f
C1192 via23_4_89/m2_1_40# VSUBS 0.364f
C1193 via23_4_23/m2_1_40# VSUBS 0.253f
C1194 via23_4_711/m2_1_40# VSUBS 0.373f
C1195 via23_4_250/m2_1_40# VSUBS 0.373f
C1196 via23_4_333/m2_1_40# VSUBS 0.373f
C1197 n7 VSUBS 65.9f
C1198 via23_4_22/m2_1_40# VSUBS 0.253f
C1199 via23_4_710/m2_1_40# VSUBS 0.373f
C1200 via23_4_249/m2_1_40# VSUBS 0.373f
C1201 via23_4_367/m2_1_40# VSUBS 0.509f
C1202 via23_4_332/m2_1_40# VSUBS 0.373f
C1203 via23_4_2/m2_1_40# VSUBS 0.243f
C1204 via23_4_87/m2_1_40# VSUBS 0.253f
C1205 via23_4_705/m2_1_40# VSUBS 0.372f
C1206 via23_4_366/m2_1_40# VSUBS 0.308f
C1207 via23_4_331/m2_1_40# VSUBS 0.373f
C1208 via23_4_354/m2_1_40# VSUBS 0.373f
C1209 n6 VSUBS 31.9f
C1210 via23_4_88/m2_1_40# VSUBS 0.253f
C1211 via23_4_704/m2_1_40# VSUBS 0.372f
C1212 via23_4_369/m2_1_40# VSUBS 0.3f
C1213 via23_4_96/m2_1_40# VSUBS 0.388f
C1214 via23_4_368/m2_1_40# VSUBS 0.3f
C1215 via23_4_598/m2_1_40# VSUBS 0.373f
C1216 via23_4_95/m2_1_40# VSUBS 0.253f
C1217 via23_4_702/m2_1_40# VSUBS 0.509f
C1218 via23_4_347/m2_1_40# VSUBS 0.373f
C1219 via23_4_94/m2_1_40# VSUBS 0.253f
C1220 n2 VSUBS 7.31f
C1221 via23_4_675/m2_1_40# VSUBS 0.373f
C1222 via23_4_588/m2_1_40# VSUBS 0.373f
C1223 top VSUBS 30.9f
C1224 via23_4_381/m2_1_40# VSUBS 0.3f
C1225 via23_4_600/m2_1_40# VSUBS 0.373f
C1226 via23_4_380/m2_1_40# VSUBS 0.411f
C1227 via23_4_584/m2_1_40# VSUBS 0.373f
C1228 via23_4_599/m2_1_40# VSUBS 0.485f
C1229 via23_4_245/m2_1_40# VSUBS 0.373f
C1230 via23_4_90/m2_1_40# VSUBS 0.253f
C1231 via23_4_218/m2_1_40# VSUBS 0.373f
C1232 via23_4_251/m2_1_40# VSUBS 0.373f
C1233 via23_4_590/m2_1_40# VSUBS 0.373f
C1234 via23_4_230/m2_1_40# VSUBS 0.373f
C1235 via23_4_589/m2_1_40# VSUBS 0.373f
C1236 ndum VSUBS 6.68f
C1237 via23_4_228/m2_1_40# VSUBS 0.509f
C1238 via23_4_229/m2_1_40# VSUBS 0.373f
C1239 via23_4_419/m2_1_40# VSUBS 0.372f
C1240 via23_4_439/m2_1_40# VSUBS 0.291f
C1241 via23_4_429/m2_1_40# VSUBS 0.372f
C1242 via23_4_449/m2_1_40# VSUBS 0.402f
C1243 via23_4_213/m2_1_40# VSUBS 0.372f
C1244 via23_4_448/m2_1_40# VSUBS 0.291f
.ends

.subckt DAC enb en_buf ctl1 ctl0 dum ctl3 ctl4 ctl5 ctl6 ctl7 ctl2 vdd vss sample
+ out vin
Xinv2_0 vdd vdd ctl7 carray_0/n7 vss vss inv2
Xinv2_1 vdd vdd ctl6 carray_0/n6 vss vss inv2
Xinv2_2 vdd vdd dum carray_0/ndum vss vss inv2
Xinv2_3 vdd vdd ctl0 carray_0/n0 vss vss inv2
Xinv2_4 vdd vdd ctl1 carray_0/n1 vss vss inv2
Xinv2_5 vdd vdd ctl5 carray_0/n5 vss vss inv2
Xinv2_6 vdd vdd ctl4 carray_0/n4 vss vss inv2
Xinv2_7 vdd vdd ctl2 carray_0/n2 vss vss inv2
Xinv2_8 vdd vdd ctl3 carray_0/n3 vss vss inv2
Xsw_top_0 sample sw_top_0/m2_1158_361# vdd out vdd vin sw_top_0/m2_990_200# vss sw_top
Xcarray_0 carray_0/n2 carray_0/n3 carray_0/n0 carray_0/via23_4_702/m2_1_40# carray_0/m2_800_1156#
+ carray_0/via23_4_459/m2_1_40# carray_0/m2_27200_1156# carray_0/m2_23300_1156# carray_0/m2_28500_1156#
+ carray_0/via23_4_447/m2_1_40# carray_0/m2_24600_1156# carray_0/m2_29800_1156# carray_0/m2_35000_1156#
+ carray_0/m2_31100_1156# carray_0/m2_25900_1156# carray_0/via23_4_369/m2_1_40# carray_0/m2_36300_1156#
+ carray_0/via23_4_379/m2_1_40# carray_0/m2_32400_1156# carray_0/m2_37600_1156# carray_0/m3_42700_1156#
+ carray_0/m2_33700_1156# carray_0/m2_38900_1156# carray_0/m3_900_1156# carray_0/via23_4_635/m2_1_40#
+ carray_0/via23_4_455/m2_1_40# carray_0/via23_4_414/m2_1_40# carray_0/via23_4_439/m2_1_40#
+ carray_0/m2_40200_1156# carray_0/via23_4_460/m2_1_40# carray_0/via23_4_704/m2_1_40#
+ carray_0/m2_41500_1156# carray_0/via23_4_366/m2_1_40# carray_0/via23_4_429/m2_1_40#
+ carray_0/m2_42800_1156# carray_0/n4 carray_0/via23_4_128/m2_1_40# carray_0/via23_4_458/m2_1_40#
+ carray_0/ndum carray_0/via23_4_381/m2_1_40# carray_0/via23_4_419/m2_1_40# carray_0/via23_4_449/m2_1_40#
+ carray_0/via23_4_641/m2_1_40# carray_0/via23_4_378/m2_1_40# carray_0/n1 carray_0/n6
+ carray_0/via23_4_642/m2_1_40# carray_0/via23_4_368/m2_1_40# carray_0/via23_4_705/m2_1_40#
+ carray_0/via23_4_446/m2_1_40# carray_0/via23_4_96/m2_1_40# out carray_0/n5 carray_0/via23_4_448/m2_1_40#
+ carray_0/m3_42500_1156# vss carray_0/via23_4_380/m2_1_40# carray_0/n7 carray_0/via23_4_367/m2_1_40#
+ carray
Xsw_top_1 sample enb vdd out vdd vin en_buf vss sw_top
Xsw_top_2 sample enb vdd out vdd vin en_buf vss sw_top
Xsw_top_3 sample sw_top_3/m2_1158_361# vdd out vdd vin sw_top_3/m2_990_200# vss sw_top
* X0 vdd sample.t5 sw_top_0/m2_1158_361# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X1 vdd vss.t7 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=14.6 ps=142 w=0 l=0
* X2 out.t98 carray_0/via23_4_600/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X3 vdd vss.t1 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X4 out.t33 carray_0/via23_4_676/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X5 out.t10 carray_0/via23_4_709/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X6 out.t17 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X7 out.t277 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X8 carray_0/n1 ctl1.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X9 vdd sample.t17 enb vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X10 vss sample.t14 enb vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X11 out.t11 carray_0/via23_4_642/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X12 out.t314 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X13 out.t212 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X14 out.t168 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X15 carray_0/n4 ctl4.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X16 sw_top_3/m2_1158_361# sample.t31 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X17 sw_top_0/m2_1158_361# sample.t7 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X18 en_buf enb.t12 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X19 out.t177 carray_0/via23_4_635/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X20 out.t318 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X21 out.t237 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X22 out.t149 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X23 out.t339 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X24 out.t243 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X25 out.t113 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X26 out.t131 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X27 out.t120 carray_0/via23_4_705/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X28 out.t291 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X29 out.t255 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X30 out.t182 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X31 out.t39 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X32 out.t9 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X33 out.t153 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X34 out.t115 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X35 out en_buf vin vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X36 out.t29 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X37 out.t285 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X38 out.t194 carray_0/via23_4_87/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X39 out.t162 carray_0/via23_4_91/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X40 vin enb out vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X41 vdd enb.t15 en_buf vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X42 out.t172 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X43 out.t141 carray_0/via23_4_369/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X44 out.t70 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X45 carray_0/n2 ctl2.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X46 out.t13 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X47 out.t299 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X48 out.t152 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X49 en_buf enb vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X50 out.t90 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X51 out.t112 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X52 out.t27 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X53 carray_0/n5 ctl5.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X54 out.t108 carray_0/via23_4_2/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X55 out.t192 carray_0/via23_4_460/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X56 out.t84 carray_0/via23_4_449/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X57 out.t71 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X58 enb sample.t12 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X59 out.t82 carray_0/via23_4_704/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X60 out.t297 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X61 out.t265 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X62 out.t213 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X63 out.t165 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X64 out.t147 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X65 out.t295 carray_0/n3 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X66 out.t248 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X67 out.t214 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X68 out.t92 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X69 vss enb en_buf vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X70 out.t97 carray_0/via23_4_702/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X71 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=9.44 ps=103 w=0 l=0
* X72 out.t238 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X73 out.t49 carray_0/via23_4_326/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X74 out.t256 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X75 out.t205 carray_0/via23_4_346/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X76 out.t139 carray_0/via23_4_333/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X77 out.t290 carray_0/n3 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X78 out.t264 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X79 out.t188 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X80 out.t130 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X81 out.t110 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X82 vss ctl5.t0 carray_0/n5 vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X83 out.t268 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X84 vss sample.t16 enb vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X85 out.t246 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X86 vss sample.t8 enb vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X87 out.t196 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X88 out.t158 carray_0/via23_4_347/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X89 out.t287 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X90 out.t233 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X91 out en_buf vin vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X92 enb sample.t20 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X93 out.t171 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X94 out.t132 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X95 vin en_buf.t0 out vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X96 carray_0/ndum dum.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X97 carray_0/n1 ctl1.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X98 out.t292 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X99 out.t244 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X100 out enb.t7 vin vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=0 l=0
* X101 out.t55 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X102 vin enb.t2 out vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X103 out.t312 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X104 out.t86 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X105 out.t54 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X106 vin enb out vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X107 carray_0/n4 ctl4.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X108 out.t260 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X109 out.t331 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X110 out.t26 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X111 out.t307 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X112 out.t116 carray_0/n2 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X113 carray_0/n0 ctl0.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X114 out.t251 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X115 vdd sample.t9 enb vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X116 out.t170 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X117 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X118 vss dum.t0 carray_0/ndum vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X119 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X120 out.t286 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X121 out.t254 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X122 out.t236 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X123 out en_buf vin vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X124 out.t306 carray_0/n1 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X125 out.t166 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X126 out.t183 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X127 out.t129 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X128 vin en_buf out vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=0 l=0
* X129 en_buf enb vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X130 vin en_buf.t8 out vss sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=0 l=0
* X131 en_buf enb.t13 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X132 out.t159 carray_0/via23_4_229/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X133 out.t81 carray_0/via23_4_245/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X134 out enb vin vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X135 out enb.t1 vin vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X136 out.t64 carray_0/via23_4_251/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X137 out.t122 carray_0/via23_4_447/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X138 out.t160 carray_0/via23_4_378/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X139 out.t65 carray_0/via23_4_381/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X140 out.t296 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X141 out.t253 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X142 out.t199 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X143 out.t242 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X144 out.t215 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X145 out en_buf.t1 vin vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X146 out.t35 carray_0/via23_4_588/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X147 out.t157 carray_0/via23_4_598/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X148 out.t187 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X149 out.t259 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X150 out.t231 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X151 vin enb.t0 out vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X152 out.t283 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X153 vdd ctl0.t2 carray_0/n0 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X154 vin enb out vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X155 en_buf enb vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X156 out.t34 carray_0/via23_4_675/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X157 out.t87 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X158 enb sample.t10 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X159 out.t51 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X160 out.t77 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X161 vdd enb en_buf vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X162 out.t25 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X163 vin en_buf.t2 out vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X164 out.t227 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X165 out.t326 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X166 out.t59 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X167 vin enb out vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X168 out.t247 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X169 out.t52 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X170 out.t151 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X171 out enb.t9 vin vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X172 out.t252 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X173 vdd sample.t13 enb vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X174 vdd sample.t21 enb vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X175 out.t218 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X176 carray_0/n7 ctl7.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X177 out.t134 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X178 out.t263 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X179 vdd ctl1.t2 carray_0/n1 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X180 out.t5 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X181 enb sample.t18 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X182 out.t109 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X183 out.t20 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X184 out.t78 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X185 carray_0/n3 ctl3.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X186 out en_buf vin vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=0 l=0
* X187 vdd ctl4.t2 carray_0/n4 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X188 vss sample.t6 sw_top_0/m2_1158_361# vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X189 out.t101 carray_0/via23_4_367/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X190 vdd vss.t6 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X191 out.t66 carray_0/via23_4_89/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X192 out.t164 carray_0/via23_4_22/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X193 out.t72 carray_0/via23_4_9/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X194 vdd ctl7.t2 carray_0/n7 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X195 out.t329 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X196 out.t36 carray_0/via23_4_429/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X197 out.t313 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X198 out.t288 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X199 out.t280 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X200 out.t89 carray_0/via23_4_1/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X201 out.t62 carray_0/via23_4_678/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X202 out.t50 carray_0/via23_4_414/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X203 out.t0 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X204 en_buf enb.t17 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X205 out.t308 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X206 out.t261 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X207 en_buf enb vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X208 out.t293 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X209 out.t249 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X210 out.t128 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X211 out.t338 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X212 out.t257 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X213 out.t58 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X214 out.t2 carray_0/via23_4_712/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X215 out.t225 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X216 out.t189 carray_0/via23_4_345/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X217 out.t118 carray_0/via23_4_332/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X218 out.t269 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X219 out.t75 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X220 out enb.t4 vin vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X221 out.t273 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X222 out.t211 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X223 out.t311 carray_0/n1 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X224 out.t88 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X225 sw_top_3/m2_1158_361# sample.t28 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X226 out.t173 carray_0/n2 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X227 out.t67 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X228 out.t208 carray_0/via23_4_419/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X229 vss sample.t30 sw_top_3/m2_1158_361# vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X230 out.t303 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X231 out.t298 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X232 out.t272 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X233 out.t235 carray_0/via23_4_95/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X234 out.t143 carray_0/via23_4_103/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X235 out.t103 carray_0/via23_4_90/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X236 out.t330 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X237 out.t322 carray_0/n3 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X238 out.t21 carray_0/via23_4_641/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X239 enb sample.t11 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X240 enb sample.t19 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X241 out.t316 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X242 out.t245 carray_0/via23_4_200/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X243 out.t240 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X244 out.t270 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X245 out.t241 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X246 out.t184 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X247 out.t275 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X248 out.t94 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X249 carray_0/n7 ctl7.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X250 out.t230 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X251 out.t100 carray_0/via23_4_198/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X252 vss ctl1.t0 carray_0/n1 vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X253 out.t217 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X254 out.t282 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X255 out.t262 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X256 out.t181 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X257 out.t133 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X258 carray_0/n3 ctl3.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X259 out.t23 carray_0/via23_4_448/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X260 out.t179 carray_0/via23_4_459/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X261 out.t140 carray_0/via23_4_213/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X262 vss ctl4.t0 carray_0/n4 vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X263 out.t206 carray_0/via23_4_218/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X264 out.t234 carray_0/via23_4_250/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X265 out.t325 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X266 out.t220 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X267 out.t22 carray_0/via23_4_439/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X268 vss ctl7.t0 carray_0/n7 vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X269 vss ctl0.t0 carray_0/n0 vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X270 out.t203 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X271 out.t320 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X272 out.t319 carray_0/n3 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X273 out.t332 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X274 out.t327 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X275 vdd sample.t1 sw_top_0/m2_1158_361# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X276 vin en_buf out vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X277 out.t80 carray_0/via23_4_584/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X278 out.t63 carray_0/via23_4_590/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X279 vdd vss.t0 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X280 out.t321 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X281 out.t250 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X282 out.t232 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X283 out.t266 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X284 out enb vin vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X285 out.t119 carray_0/via23_4_220/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X286 out.t228 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X287 out.t198 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X288 out.t53 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X289 out.t32 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X290 out.t274 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X291 out.t135 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X292 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X293 out.t175 carray_0/via23_4_228/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X294 out.t24 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X295 out.t154 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X296 out.t44 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X297 out.t204 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X298 out.t328 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X299 out.t85 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X300 carray_0/n6 ctl6.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X301 out.t309 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X302 out.t4 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X303 out.t76 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X304 out.t335 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X305 out.t301 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X306 out.t219 carray_0/n4 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X307 out.t304 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X308 out.t104 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X309 out.t317 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X310 vdd vss.t5 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X311 vdd vss.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X312 out.t294 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X313 out.t145 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X314 out.t324 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X315 sw_top_3/m2_1158_361# sample.t26 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X316 out.t191 carray_0/via23_4_380/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X317 out en_buf.t3 vin vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=0 l=0
* X318 vdd sample.t25 sw_top_3/m2_1158_361# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X319 out.t15 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X320 vin en_buf out vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X321 vin en_buf.t7 out vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X322 out.t83 carray_0/via23_4_366/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X323 out enb vin vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X324 enb sample.t23 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X325 out.t146 carray_0/via23_4_21/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X326 enb sample.t15 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X327 out.t56 carray_0/via23_4_3/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X328 vin enb.t5 out vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X329 out.t41 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X330 out.t337 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X331 out.t7 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X332 out.t114 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X333 out.t186 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X334 out.t284 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X335 out.t57 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X336 vdd ctl3.t2 carray_0/n3 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X337 out.t117 carray_0/via23_4_601/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X338 out.t47 carray_0/via23_4_677/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X339 out.t137 carray_0/via23_4_710/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X340 out.t150 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X341 sw_top_0/m2_1158_361# sample.t4 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X342 out.t267 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X343 out.t74 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X344 out.t124 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X345 out.t289 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X346 out.t125 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X347 out.t68 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X348 vdd ctl6.t2 carray_0/n6 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X349 out en_buf.t6 vin vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X350 out en_buf vin vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X351 out.t14 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X352 out.t105 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X353 out.t99 carray_0/via23_4_331/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X354 vdd ctl2.t2 carray_0/n2 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X355 out.t38 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X356 out.t221 carray_0/via23_4_334/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X357 vdd vss.t4 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X358 out enb vin vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X359 vin enb.t3 out vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=0 l=0
* X360 out.t37 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X361 vin enb out vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=0 l=0
* X362 out.t163 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X363 out.t12 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X364 out.t28 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X365 out.t323 carray_0/n0 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X366 vss enb.t16 en_buf vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X367 out.t239 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X368 out.t167 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X369 vss enb en_buf vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X370 out.t333 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X371 vin en_buf out vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X372 vin en_buf.t5 out vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X373 out.t136 carray_0/n2 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X374 out.t69 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X375 out.t148 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X376 out.t91 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X377 out.t111 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X378 carray_0/n6 ctl6.t1 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X379 out.t276 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X380 out.t176 carray_0/via23_4_94/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X381 out.t209 carray_0/via23_4_88/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X382 out.t93 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X383 out.t300 carray_0/n3 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X384 out.t210 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X385 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X386 out.t31 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X387 out enb.t6 vin vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X388 out.t96 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X389 out.t258 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X390 out.t197 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X391 out.t40 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X392 out.t279 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X393 vss sample.t0 sw_top_0/m2_1158_361# vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X394 vss sample.t24 sw_top_3/m2_1158_361# vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X395 out.t216 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X396 out.t200 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X397 out.t3 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X398 out.t144 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X399 out.t161 carray_0/via23_4_455/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X400 out.t142 carray_0/via23_4_458/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X401 out.t336 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X402 vin en_buf out vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X403 out.t222 carray_0/via23_4_249/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X404 out.t190 carray_0/via23_4_230/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X405 out en_buf.t4 vin vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X406 vss sample.t22 enb vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X407 out.t310 carray_0/n3 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X408 out.t126 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X409 vin enb.t8 out vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X410 out.t156 carray_0/via23_4_711/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X411 sw_top_0/m2_1158_361# sample.t3 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X412 sw_top_3/m2_1158_361# sample.t27 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0 l=0
* X413 out.t334 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X414 out.t315 carray_0/n3 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X415 out.t305 carray_0/n3 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X416 en_buf enb.t14 vss vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X417 out.t195 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X418 out.t8 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X419 out.t123 carray_0/via23_4_96/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X420 vss ctl3.t0 carray_0/n3 vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X421 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X422 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X423 out.t174 carray_0/via23_4_354/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X424 out.t138 carray_0/via23_4_599/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X425 out.t48 carray_0/via23_4_589/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X426 out.t223 carray_0/via23_4_128/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X427 vss ctl6.t0 carray_0/n6 vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X428 out.t302 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X429 out.t271 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X430 out enb vin vdd sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=0 l=0
* X431 out.t193 carray_0/via23_4_117/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X432 vss ctl2.t0 carray_0/n2 vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0 l=0
* X433 out.t226 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X434 out.t185 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X435 out.t45 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X436 out.t46 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X437 vss enb.t10 en_buf vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0 l=0
* X438 out.t278 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X439 sw_top_0/m2_1158_361# sample.t2 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X440 out.t73 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X441 out.t1 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X442 out.t61 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X443 out.t155 carray_0/n2 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X444 carray_0/ndum dum.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X445 out.t107 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X446 out.t19 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X447 out.t30 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X448 out.t95 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X449 vdd vss.t2 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
* X450 out en_buf.t9 vin vss sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=0 l=0
* X451 out.t43 carray_0/ndum sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X452 out.t106 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X453 carray_0/n2 ctl2.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X454 vdd enb en_buf vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X455 vdd enb.t11 en_buf vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X456 carray_0/n0 ctl0.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X457 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
* X458 out.t207 carray_0/via23_4_111/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X459 carray_0/n5 ctl5.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=0 l=0
* X460 out.t102 carray_0/via23_4_446/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X461 vdd dum.t2 carray_0/ndum vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X462 out.t178 carray_0/via23_4_379/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X463 out.t121 carray_0/via23_4_368/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X464 out.t79 carray_0/via23_4_199/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X465 out.t6 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X466 out.t229 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X467 out.t169 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X468 out.t127 carray_0/via23_4_20/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X469 out.t180 carray_0/via23_4_23/m2_1_40# sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X470 out.t16 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X471 out.t201 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X472 out.t224 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X473 out.t202 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X474 out.t60 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X475 out.t18 carray_0/n7 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X476 vdd ctl5.t2 carray_0/n5 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=0 l=0
* X477 out.t42 carray_0/n6 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
* X478 vdd sample.t29 sw_top_3/m2_1158_361# vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=0 l=0
* X479 out.t281 carray_0/n5 sky130_fd_pr__cap_mim_m3_1 l=0 w=0
R0 ctl7.n0 ctl7.t2 212.081
R1 ctl7.n1 ctl7.t3 212.081
R2 ctl7.n0 ctl7.t0 139.78
R3 ctl7.n1 ctl7.t1 139.78
R4 ctl7.n1 ctl7.n0 61.346
R5 ctl7 ctl7.n1 44.6884
R6 vss.n134 vss.n133 17788.9
R7 vss.n135 vss.n134 4406.54
R8 vss.n124 vss.n123 3471.83
R9 vss.n675 vss.n674 1717.31
R10 vss.n457 vss.n456 1717.31
R11 vss.n296 vss.n295 1717.31
R12 vss.n675 vss.n673 611.246
R13 vss.n457 vss.n455 611.246
R14 vss.n296 vss.n294 611.246
R15 vss.n135 vss.n45 611.246
R16 vss.n123 vss.n48 511.757
R17 vss.n125 vss.n124 481.067
R18 vss.n56 vss.n55 294.462
R19 vss.n834 vss.n833 292.5
R20 vss.n833 vss.n832 292.5
R21 vss.n830 vss.n829 292.5
R22 vss.n829 vss.n828 292.5
R23 vss.n781 vss.n780 292.5
R24 vss.n780 vss.n779 292.5
R25 vss.n777 vss.n776 292.5
R26 vss.n776 vss.n775 292.5
R27 vss.n668 vss.n667 292.5
R28 vss.n666 vss.n665 292.5
R29 vss.n664 vss.n663 292.5
R30 vss.n662 vss.n661 292.5
R31 vss.n660 vss.n659 292.5
R32 vss.n658 vss.n657 292.5
R33 vss.n656 vss.n655 292.5
R34 vss.n654 vss.n653 292.5
R35 vss.n652 vss.n651 292.5
R36 vss.n650 vss.n649 292.5
R37 vss.n648 vss.n647 292.5
R38 vss.n646 vss.n645 292.5
R39 vss.n644 vss.n643 292.5
R40 vss.n642 vss.n641 292.5
R41 vss.n640 vss.n639 292.5
R42 vss.n638 vss.n637 292.5
R43 vss.n636 vss.n635 292.5
R44 vss.n634 vss.n633 292.5
R45 vss.n632 vss.n631 292.5
R46 vss.n629 vss.n628 292.5
R47 vss.n569 vss.n568 292.5
R48 vss.n573 vss.n572 292.5
R49 vss.n576 vss.n575 292.5
R50 vss.n575 vss.n574 292.5
R51 vss.n579 vss.n578 292.5
R52 vss.n578 vss.n577 292.5
R53 vss.n582 vss.n581 292.5
R54 vss.n581 vss.n580 292.5
R55 vss.n585 vss.n584 292.5
R56 vss.n584 vss.n583 292.5
R57 vss.n588 vss.n587 292.5
R58 vss.n587 vss.n586 292.5
R59 vss.n591 vss.n590 292.5
R60 vss.n590 vss.n589 292.5
R61 vss.n594 vss.n593 292.5
R62 vss.n593 vss.n592 292.5
R63 vss.n597 vss.n596 292.5
R64 vss.n596 vss.n595 292.5
R65 vss.n600 vss.n599 292.5
R66 vss.n599 vss.n598 292.5
R67 vss.n603 vss.n602 292.5
R68 vss.n602 vss.n601 292.5
R69 vss.n606 vss.n605 292.5
R70 vss.n605 vss.n604 292.5
R71 vss.n609 vss.n608 292.5
R72 vss.n608 vss.n607 292.5
R73 vss.n612 vss.n611 292.5
R74 vss.n611 vss.n610 292.5
R75 vss.n615 vss.n614 292.5
R76 vss.n614 vss.n613 292.5
R77 vss.n618 vss.n617 292.5
R78 vss.n617 vss.n616 292.5
R79 vss.n621 vss.n620 292.5
R80 vss.n620 vss.n619 292.5
R81 vss.n624 vss.n623 292.5
R82 vss.n623 vss.n622 292.5
R83 vss.n626 vss.n625 292.5
R84 vss.n450 vss.n449 292.5
R85 vss.n448 vss.n447 292.5
R86 vss.n446 vss.n445 292.5
R87 vss.n444 vss.n443 292.5
R88 vss.n442 vss.n441 292.5
R89 vss.n440 vss.n439 292.5
R90 vss.n438 vss.n437 292.5
R91 vss.n436 vss.n435 292.5
R92 vss.n434 vss.n433 292.5
R93 vss.n432 vss.n431 292.5
R94 vss.n430 vss.n429 292.5
R95 vss.n428 vss.n427 292.5
R96 vss.n426 vss.n425 292.5
R97 vss.n424 vss.n423 292.5
R98 vss.n422 vss.n421 292.5
R99 vss.n420 vss.n419 292.5
R100 vss.n418 vss.n417 292.5
R101 vss.n416 vss.n415 292.5
R102 vss.n414 vss.n413 292.5
R103 vss.n411 vss.n410 292.5
R104 vss.n499 vss.n498 292.5
R105 vss.n503 vss.n502 292.5
R106 vss.n506 vss.n505 292.5
R107 vss.n505 vss.n504 292.5
R108 vss.n509 vss.n508 292.5
R109 vss.n508 vss.n507 292.5
R110 vss.n512 vss.n511 292.5
R111 vss.n511 vss.n510 292.5
R112 vss.n515 vss.n514 292.5
R113 vss.n514 vss.n513 292.5
R114 vss.n518 vss.n517 292.5
R115 vss.n517 vss.n516 292.5
R116 vss.n521 vss.n520 292.5
R117 vss.n520 vss.n519 292.5
R118 vss.n524 vss.n523 292.5
R119 vss.n523 vss.n522 292.5
R120 vss.n527 vss.n526 292.5
R121 vss.n526 vss.n525 292.5
R122 vss.n530 vss.n529 292.5
R123 vss.n529 vss.n528 292.5
R124 vss.n533 vss.n532 292.5
R125 vss.n532 vss.n531 292.5
R126 vss.n536 vss.n535 292.5
R127 vss.n535 vss.n534 292.5
R128 vss.n539 vss.n538 292.5
R129 vss.n538 vss.n537 292.5
R130 vss.n542 vss.n541 292.5
R131 vss.n541 vss.n540 292.5
R132 vss.n545 vss.n544 292.5
R133 vss.n544 vss.n543 292.5
R134 vss.n548 vss.n547 292.5
R135 vss.n547 vss.n546 292.5
R136 vss.n551 vss.n550 292.5
R137 vss.n550 vss.n549 292.5
R138 vss.n554 vss.n553 292.5
R139 vss.n553 vss.n552 292.5
R140 vss.n556 vss.n555 292.5
R141 vss.n289 vss.n288 292.5
R142 vss.n287 vss.n286 292.5
R143 vss.n285 vss.n284 292.5
R144 vss.n283 vss.n282 292.5
R145 vss.n281 vss.n280 292.5
R146 vss.n279 vss.n278 292.5
R147 vss.n277 vss.n276 292.5
R148 vss.n275 vss.n274 292.5
R149 vss.n273 vss.n272 292.5
R150 vss.n271 vss.n270 292.5
R151 vss.n269 vss.n268 292.5
R152 vss.n267 vss.n266 292.5
R153 vss.n265 vss.n264 292.5
R154 vss.n263 vss.n262 292.5
R155 vss.n261 vss.n260 292.5
R156 vss.n259 vss.n258 292.5
R157 vss.n257 vss.n256 292.5
R158 vss.n255 vss.n254 292.5
R159 vss.n253 vss.n252 292.5
R160 vss.n250 vss.n249 292.5
R161 vss.n338 vss.n337 292.5
R162 vss.n342 vss.n341 292.5
R163 vss.n345 vss.n344 292.5
R164 vss.n344 vss.n343 292.5
R165 vss.n348 vss.n347 292.5
R166 vss.n347 vss.n346 292.5
R167 vss.n351 vss.n350 292.5
R168 vss.n350 vss.n349 292.5
R169 vss.n354 vss.n353 292.5
R170 vss.n353 vss.n352 292.5
R171 vss.n357 vss.n356 292.5
R172 vss.n356 vss.n355 292.5
R173 vss.n360 vss.n359 292.5
R174 vss.n359 vss.n358 292.5
R175 vss.n363 vss.n362 292.5
R176 vss.n362 vss.n361 292.5
R177 vss.n366 vss.n365 292.5
R178 vss.n365 vss.n364 292.5
R179 vss.n369 vss.n368 292.5
R180 vss.n368 vss.n367 292.5
R181 vss.n372 vss.n371 292.5
R182 vss.n371 vss.n370 292.5
R183 vss.n375 vss.n374 292.5
R184 vss.n374 vss.n373 292.5
R185 vss.n378 vss.n377 292.5
R186 vss.n377 vss.n376 292.5
R187 vss.n381 vss.n380 292.5
R188 vss.n380 vss.n379 292.5
R189 vss.n384 vss.n383 292.5
R190 vss.n383 vss.n382 292.5
R191 vss.n387 vss.n386 292.5
R192 vss.n386 vss.n385 292.5
R193 vss.n390 vss.n389 292.5
R194 vss.n389 vss.n388 292.5
R195 vss.n393 vss.n392 292.5
R196 vss.n392 vss.n391 292.5
R197 vss.n395 vss.n394 292.5
R198 vss.n40 vss.n39 292.5
R199 vss.n38 vss.n37 292.5
R200 vss.n36 vss.n35 292.5
R201 vss.n34 vss.n33 292.5
R202 vss.n32 vss.n31 292.5
R203 vss.n30 vss.n29 292.5
R204 vss.n28 vss.n27 292.5
R205 vss.n26 vss.n25 292.5
R206 vss.n24 vss.n23 292.5
R207 vss.n22 vss.n21 292.5
R208 vss.n20 vss.n19 292.5
R209 vss.n18 vss.n17 292.5
R210 vss.n16 vss.n15 292.5
R211 vss.n14 vss.n13 292.5
R212 vss.n12 vss.n11 292.5
R213 vss.n10 vss.n9 292.5
R214 vss.n8 vss.n7 292.5
R215 vss.n6 vss.n5 292.5
R216 vss.n4 vss.n3 292.5
R217 vss.n1 vss.n0 292.5
R218 vss.n177 vss.n176 292.5
R219 vss.n181 vss.n180 292.5
R220 vss.n184 vss.n183 292.5
R221 vss.n183 vss.n182 292.5
R222 vss.n187 vss.n186 292.5
R223 vss.n186 vss.n185 292.5
R224 vss.n190 vss.n189 292.5
R225 vss.n189 vss.n188 292.5
R226 vss.n193 vss.n192 292.5
R227 vss.n192 vss.n191 292.5
R228 vss.n196 vss.n195 292.5
R229 vss.n195 vss.n194 292.5
R230 vss.n199 vss.n198 292.5
R231 vss.n198 vss.n197 292.5
R232 vss.n202 vss.n201 292.5
R233 vss.n201 vss.n200 292.5
R234 vss.n205 vss.n204 292.5
R235 vss.n204 vss.n203 292.5
R236 vss.n208 vss.n207 292.5
R237 vss.n207 vss.n206 292.5
R238 vss.n211 vss.n210 292.5
R239 vss.n210 vss.n209 292.5
R240 vss.n214 vss.n213 292.5
R241 vss.n213 vss.n212 292.5
R242 vss.n217 vss.n216 292.5
R243 vss.n216 vss.n215 292.5
R244 vss.n220 vss.n219 292.5
R245 vss.n219 vss.n218 292.5
R246 vss.n223 vss.n222 292.5
R247 vss.n222 vss.n221 292.5
R248 vss.n226 vss.n225 292.5
R249 vss.n225 vss.n224 292.5
R250 vss.n229 vss.n228 292.5
R251 vss.n228 vss.n227 292.5
R252 vss.n232 vss.n231 292.5
R253 vss.n231 vss.n230 292.5
R254 vss.n234 vss.n233 292.5
R255 vss.n122 vss.n121 292.5
R256 vss.n123 vss.n122 292.5
R257 vss.n53 vss.n52 292.5
R258 vss.n52 vss.n51 292.5
R259 vss.n55 vss.n54 292.5
R260 vss.n717 vss.t5 188.089
R261 vss.n734 vss.t7 183.082
R262 vss.n787 vss.t3 183.082
R263 vss.n840 vss.t1 183.082
R264 vss.n122 vss.n49 172.611
R265 vss.n568 vss.n567 147.374
R266 vss.n498 vss.n497 147.374
R267 vss.n337 vss.n336 147.374
R268 vss.n176 vss.n175 147.374
R269 vss.n571 vss.n570 134.577
R270 vss.n501 vss.n500 134.577
R271 vss.n340 vss.n339 134.577
R272 vss.n179 vss.n178 134.577
R273 vss.n572 vss.n571 90.6382
R274 vss.n502 vss.n501 90.6382
R275 vss.n341 vss.n340 90.6382
R276 vss.n180 vss.n179 90.6382
R277 vss.n3 vss.n2 90.6381
R278 vss.n252 vss.n251 90.6381
R279 vss.n413 vss.n412 90.6381
R280 vss.n631 vss.n630 90.6381
R281 vss.n184 vss.n181 87.7181
R282 vss.n6 vss.n4 87.7181
R283 vss.n345 vss.n342 87.7181
R284 vss.n255 vss.n253 87.7181
R285 vss.n506 vss.n503 87.7181
R286 vss.n416 vss.n414 87.7181
R287 vss.n576 vss.n573 87.7181
R288 vss.n634 vss.n632 87.7181
R289 vss.n44 vss.n43 86.9123
R290 vss.n293 vss.n292 86.9123
R291 vss.n454 vss.n453 86.9123
R292 vss.n672 vss.n671 86.9123
R293 vss.n41 vss.n40 82.0711
R294 vss.n290 vss.n289 82.0711
R295 vss.n451 vss.n450 82.0711
R296 vss.n669 vss.n668 82.0711
R297 vss.n235 vss.n234 78.3064
R298 vss.n396 vss.n395 78.3064
R299 vss.n557 vss.n556 78.3064
R300 vss.n627 vss.n626 78.3064
R301 vss.n887 vss.n886 76.0005
R302 vss.n246 vss.n245 76.0005
R303 vss.n407 vss.n406 76.0005
R304 vss.n564 vss.n563 76.0005
R305 vss.n156 vss.n155 63.7358
R306 vss.n317 vss.n316 63.7358
R307 vss.n478 vss.n477 63.7358
R308 vss.n696 vss.n695 63.7358
R309 vss.n133 vss.n132 47.743
R310 vss.n130 vss.n129 47.743
R311 vss.n129 vss.n128 47.743
R312 vss.n128 vss.n127 47.743
R313 vss.n127 vss.n126 47.743
R314 vss.n126 vss.n125 47.743
R315 vss.n170 vss.n169 46.3534
R316 vss.n331 vss.n330 46.3534
R317 vss.n492 vss.n491 46.3534
R318 vss.n710 vss.n709 46.3534
R319 vss.n145 vss.n144 35.3848
R320 vss.n306 vss.n305 35.3848
R321 vss.n467 vss.n466 35.3848
R322 vss.n685 vss.n684 35.3848
R323 vss.n684 vss.n683 35.3848
R324 vss.n466 vss.n465 35.3848
R325 vss.n305 vss.n304 35.3848
R326 vss.n144 vss.n143 35.3848
R327 vss.n562 vss.t4 34.2973
R328 vss.n405 vss.t6 34.2973
R329 vss.n244 vss.t2 34.2973
R330 vss.n885 vss.t0 34.2973
R331 vss.n697 vss.n696 32.3305
R332 vss.n479 vss.n478 32.3305
R333 vss.n318 vss.n317 32.3305
R334 vss.n157 vss.n156 32.3305
R335 vss.n131 vss.n130 31.9637
R336 vss.n187 vss.n184 25.6005
R337 vss.n190 vss.n187 25.6005
R338 vss.n193 vss.n190 25.6005
R339 vss.n196 vss.n193 25.6005
R340 vss.n199 vss.n196 25.6005
R341 vss.n202 vss.n199 25.6005
R342 vss.n205 vss.n202 25.6005
R343 vss.n208 vss.n205 25.6005
R344 vss.n211 vss.n208 25.6005
R345 vss.n214 vss.n211 25.6005
R346 vss.n217 vss.n214 25.6005
R347 vss.n220 vss.n217 25.6005
R348 vss.n223 vss.n220 25.6005
R349 vss.n226 vss.n223 25.6005
R350 vss.n229 vss.n226 25.6005
R351 vss.n232 vss.n229 25.6005
R352 vss.n234 vss.n232 25.6005
R353 vss.n181 vss.n177 25.6005
R354 vss.n4 vss.n1 25.6005
R355 vss.n8 vss.n6 25.6005
R356 vss.n10 vss.n8 25.6005
R357 vss.n12 vss.n10 25.6005
R358 vss.n14 vss.n12 25.6005
R359 vss.n16 vss.n14 25.6005
R360 vss.n18 vss.n16 25.6005
R361 vss.n20 vss.n18 25.6005
R362 vss.n22 vss.n20 25.6005
R363 vss.n24 vss.n22 25.6005
R364 vss.n26 vss.n24 25.6005
R365 vss.n28 vss.n26 25.6005
R366 vss.n30 vss.n28 25.6005
R367 vss.n32 vss.n30 25.6005
R368 vss.n34 vss.n32 25.6005
R369 vss.n36 vss.n34 25.6005
R370 vss.n38 vss.n36 25.6005
R371 vss.n40 vss.n38 25.6005
R372 vss.n348 vss.n345 25.6005
R373 vss.n351 vss.n348 25.6005
R374 vss.n354 vss.n351 25.6005
R375 vss.n357 vss.n354 25.6005
R376 vss.n360 vss.n357 25.6005
R377 vss.n363 vss.n360 25.6005
R378 vss.n366 vss.n363 25.6005
R379 vss.n369 vss.n366 25.6005
R380 vss.n372 vss.n369 25.6005
R381 vss.n375 vss.n372 25.6005
R382 vss.n378 vss.n375 25.6005
R383 vss.n381 vss.n378 25.6005
R384 vss.n384 vss.n381 25.6005
R385 vss.n387 vss.n384 25.6005
R386 vss.n390 vss.n387 25.6005
R387 vss.n393 vss.n390 25.6005
R388 vss.n395 vss.n393 25.6005
R389 vss.n342 vss.n338 25.6005
R390 vss.n253 vss.n250 25.6005
R391 vss.n257 vss.n255 25.6005
R392 vss.n259 vss.n257 25.6005
R393 vss.n261 vss.n259 25.6005
R394 vss.n263 vss.n261 25.6005
R395 vss.n265 vss.n263 25.6005
R396 vss.n267 vss.n265 25.6005
R397 vss.n269 vss.n267 25.6005
R398 vss.n271 vss.n269 25.6005
R399 vss.n273 vss.n271 25.6005
R400 vss.n275 vss.n273 25.6005
R401 vss.n277 vss.n275 25.6005
R402 vss.n279 vss.n277 25.6005
R403 vss.n281 vss.n279 25.6005
R404 vss.n283 vss.n281 25.6005
R405 vss.n285 vss.n283 25.6005
R406 vss.n287 vss.n285 25.6005
R407 vss.n289 vss.n287 25.6005
R408 vss.n509 vss.n506 25.6005
R409 vss.n512 vss.n509 25.6005
R410 vss.n515 vss.n512 25.6005
R411 vss.n518 vss.n515 25.6005
R412 vss.n521 vss.n518 25.6005
R413 vss.n524 vss.n521 25.6005
R414 vss.n527 vss.n524 25.6005
R415 vss.n530 vss.n527 25.6005
R416 vss.n533 vss.n530 25.6005
R417 vss.n536 vss.n533 25.6005
R418 vss.n539 vss.n536 25.6005
R419 vss.n542 vss.n539 25.6005
R420 vss.n545 vss.n542 25.6005
R421 vss.n548 vss.n545 25.6005
R422 vss.n551 vss.n548 25.6005
R423 vss.n554 vss.n551 25.6005
R424 vss.n556 vss.n554 25.6005
R425 vss.n503 vss.n499 25.6005
R426 vss.n414 vss.n411 25.6005
R427 vss.n418 vss.n416 25.6005
R428 vss.n420 vss.n418 25.6005
R429 vss.n422 vss.n420 25.6005
R430 vss.n424 vss.n422 25.6005
R431 vss.n426 vss.n424 25.6005
R432 vss.n428 vss.n426 25.6005
R433 vss.n430 vss.n428 25.6005
R434 vss.n432 vss.n430 25.6005
R435 vss.n434 vss.n432 25.6005
R436 vss.n436 vss.n434 25.6005
R437 vss.n438 vss.n436 25.6005
R438 vss.n440 vss.n438 25.6005
R439 vss.n442 vss.n440 25.6005
R440 vss.n444 vss.n442 25.6005
R441 vss.n446 vss.n444 25.6005
R442 vss.n448 vss.n446 25.6005
R443 vss.n450 vss.n448 25.6005
R444 vss.n579 vss.n576 25.6005
R445 vss.n582 vss.n579 25.6005
R446 vss.n585 vss.n582 25.6005
R447 vss.n588 vss.n585 25.6005
R448 vss.n591 vss.n588 25.6005
R449 vss.n594 vss.n591 25.6005
R450 vss.n597 vss.n594 25.6005
R451 vss.n600 vss.n597 25.6005
R452 vss.n603 vss.n600 25.6005
R453 vss.n606 vss.n603 25.6005
R454 vss.n609 vss.n606 25.6005
R455 vss.n612 vss.n609 25.6005
R456 vss.n615 vss.n612 25.6005
R457 vss.n618 vss.n615 25.6005
R458 vss.n621 vss.n618 25.6005
R459 vss.n624 vss.n621 25.6005
R460 vss.n626 vss.n624 25.6005
R461 vss.n573 vss.n569 25.6005
R462 vss.n632 vss.n629 25.6005
R463 vss.n636 vss.n634 25.6005
R464 vss.n638 vss.n636 25.6005
R465 vss.n640 vss.n638 25.6005
R466 vss.n642 vss.n640 25.6005
R467 vss.n644 vss.n642 25.6005
R468 vss.n646 vss.n644 25.6005
R469 vss.n648 vss.n646 25.6005
R470 vss.n650 vss.n648 25.6005
R471 vss.n652 vss.n650 25.6005
R472 vss.n654 vss.n652 25.6005
R473 vss.n656 vss.n654 25.6005
R474 vss.n658 vss.n656 25.6005
R475 vss.n660 vss.n658 25.6005
R476 vss.n662 vss.n660 25.6005
R477 vss.n664 vss.n662 25.6005
R478 vss.n666 vss.n664 25.6005
R479 vss.n668 vss.n666 25.6005
R480 vss.n168 vss.n167 24.962
R481 vss.n329 vss.n328 24.962
R482 vss.n490 vss.n489 24.962
R483 vss.n708 vss.n707 24.962
R484 vss.n709 vss.n708 24.962
R485 vss.n491 vss.n490 24.962
R486 vss.n330 vss.n329 24.962
R487 vss.n169 vss.n168 24.962
R488 vss.n146 vss.n145 23.177
R489 vss.n307 vss.n306 23.177
R490 vss.n468 vss.n467 23.177
R491 vss.n686 vss.n685 23.177
R492 vss.n830 vss.n827 16.1455
R493 vss.n777 vss.n774 16.1455
R494 vss.n725 vss.n724 16.1455
R495 vss.n676 vss.n672 11.1897
R496 vss.n458 vss.n454 11.1897
R497 vss.n297 vss.n293 11.1897
R498 vss.n136 vss.n44 11.1897
R499 vss.n150 vss.n149 9.3005
R500 vss.n162 vss.n161 9.3005
R501 vss.n152 vss.n151 9.3005
R502 vss.n164 vss.n163 9.3005
R503 vss.n174 vss.n173 9.3005
R504 vss.n236 vss.n235 9.3005
R505 vss.n311 vss.n310 9.3005
R506 vss.n323 vss.n322 9.3005
R507 vss.n313 vss.n312 9.3005
R508 vss.n325 vss.n324 9.3005
R509 vss.n335 vss.n334 9.3005
R510 vss.n397 vss.n396 9.3005
R511 vss.n472 vss.n471 9.3005
R512 vss.n484 vss.n483 9.3005
R513 vss.n474 vss.n473 9.3005
R514 vss.n486 vss.n485 9.3005
R515 vss.n496 vss.n495 9.3005
R516 vss.n558 vss.n557 9.3005
R517 vss.n872 vss.n871 9.3005
R518 vss.n690 vss.n689 9.3005
R519 vss.n702 vss.n701 9.3005
R520 vss.n715 vss.n627 9.3005
R521 vss.n692 vss.n691 9.3005
R522 vss.n704 vss.n703 9.3005
R523 vss.n714 vss.n713 9.3005
R524 vss.n688 vss.n687 9.3005
R525 vss.n687 vss.n686 9.3005
R526 vss.n700 vss.n699 9.3005
R527 vss.n699 vss.n698 9.3005
R528 vss.n678 vss.n677 9.3005
R529 vss.n712 vss.n711 9.3005
R530 vss.n711 vss.n710 9.3005
R531 vss.n470 vss.n469 9.3005
R532 vss.n469 vss.n468 9.3005
R533 vss.n482 vss.n481 9.3005
R534 vss.n481 vss.n480 9.3005
R535 vss.n460 vss.n459 9.3005
R536 vss.n494 vss.n493 9.3005
R537 vss.n493 vss.n492 9.3005
R538 vss.n309 vss.n308 9.3005
R539 vss.n308 vss.n307 9.3005
R540 vss.n321 vss.n320 9.3005
R541 vss.n320 vss.n319 9.3005
R542 vss.n299 vss.n298 9.3005
R543 vss.n333 vss.n332 9.3005
R544 vss.n332 vss.n331 9.3005
R545 vss.n148 vss.n147 9.3005
R546 vss.n147 vss.n146 9.3005
R547 vss.n160 vss.n159 9.3005
R548 vss.n159 vss.n158 9.3005
R549 vss.n138 vss.n137 9.3005
R550 vss.n172 vss.n171 9.3005
R551 vss.n171 vss.n170 9.3005
R552 vss.n877 vss.n876 9.0005
R553 vss.n676 vss.n675 8.98038
R554 vss.n458 vss.n457 8.98038
R555 vss.n297 vss.n296 8.98038
R556 vss.n136 vss.n135 8.98038
R557 vss.n131 vss.n47 8.4537
R558 vss.n121 vss.n50 6.57927
R559 vss.n42 vss.n41 5.64756
R560 vss.n291 vss.n290 5.64756
R561 vss.n452 vss.n451 5.64756
R562 vss.n670 vss.n669 5.64756
R563 vss.n131 vss.n46 5.03498
R564 vss.n141 vss.n140 4.89462
R565 vss.n302 vss.n301 4.89462
R566 vss.n463 vss.n462 4.89462
R567 vss.n681 vss.n680 4.89462
R568 vss.n563 vss.n562 4.85762
R569 vss.n406 vss.n405 4.85762
R570 vss.n245 vss.n244 4.85762
R571 vss.n886 vss.n885 4.85762
R572 vss.n738 vss.n737 4.6505
R573 vss.n742 vss.n741 4.6505
R574 vss.n746 vss.n745 4.6505
R575 vss.n748 vss.n747 4.6505
R576 vss.n752 vss.n751 4.6505
R577 vss.n756 vss.n755 4.6505
R578 vss.n791 vss.n790 4.6505
R579 vss.n795 vss.n794 4.6505
R580 vss.n799 vss.n798 4.6505
R581 vss.n801 vss.n800 4.6505
R582 vss.n805 vss.n804 4.6505
R583 vss.n809 vss.n808 4.6505
R584 vss.n844 vss.n843 4.6505
R585 vss.n848 vss.n847 4.6505
R586 vss.n852 vss.n851 4.6505
R587 vss.n854 vss.n853 4.6505
R588 vss.n858 vss.n857 4.6505
R589 vss.n862 vss.n861 4.6505
R590 vss.n890 vss.n889 4.6505
R591 vss.n870 vss.n869 4.6505
R592 vss.n868 vss.n867 4.6505
R593 vss.n866 vss.n865 4.6505
R594 vss.n842 vss.n841 4.6505
R595 vss.n839 vss.n838 4.6505
R596 vss.n835 vss.n834 4.6505
R597 vss.n831 vss.n830 4.6505
R598 vss.n827 vss.n826 4.6505
R599 vss.n817 vss.n816 4.6505
R600 vss.n815 vss.n814 4.6505
R601 vss.n813 vss.n812 4.6505
R602 vss.n789 vss.n788 4.6505
R603 vss.n786 vss.n785 4.6505
R604 vss.n782 vss.n781 4.6505
R605 vss.n778 vss.n777 4.6505
R606 vss.n774 vss.n773 4.6505
R607 vss.n764 vss.n763 4.6505
R608 vss.n762 vss.n761 4.6505
R609 vss.n760 vss.n759 4.6505
R610 vss.n736 vss.n735 4.6505
R611 vss.n733 vss.n732 4.6505
R612 vss.n729 vss.n728 4.6505
R613 vss.n726 vss.n725 4.6505
R614 vss.n724 vss.n723 4.6505
R615 vss.n731 vss.n730 4.6505
R616 vss.n740 vss.n739 4.6505
R617 vss.n744 vss.n743 4.6505
R618 vss.n750 vss.n749 4.6505
R619 vss.n754 vss.n753 4.6505
R620 vss.n758 vss.n757 4.6505
R621 vss.n784 vss.n783 4.6505
R622 vss.n793 vss.n792 4.6505
R623 vss.n797 vss.n796 4.6505
R624 vss.n803 vss.n802 4.6505
R625 vss.n807 vss.n806 4.6505
R626 vss.n811 vss.n810 4.6505
R627 vss.n837 vss.n836 4.6505
R628 vss.n846 vss.n845 4.6505
R629 vss.n850 vss.n849 4.6505
R630 vss.n856 vss.n855 4.6505
R631 vss.n860 vss.n859 4.6505
R632 vss.n864 vss.n863 4.6505
R633 vss.n58 vss.n57 4.6505
R634 vss.n62 vss.n61 4.6505
R635 vss.n64 vss.n63 4.6505
R636 vss.n68 vss.n67 4.6505
R637 vss.n70 vss.n69 4.6505
R638 vss.n74 vss.n73 4.6505
R639 vss.n76 vss.n75 4.6505
R640 vss.n80 vss.n79 4.6505
R641 vss.n82 vss.n81 4.6505
R642 vss.n86 vss.n85 4.6505
R643 vss.n88 vss.n87 4.6505
R644 vss.n92 vss.n91 4.6505
R645 vss.n94 vss.n93 4.6505
R646 vss.n98 vss.n97 4.6505
R647 vss.n100 vss.n99 4.6505
R648 vss.n104 vss.n103 4.6505
R649 vss.n106 vss.n105 4.6505
R650 vss.n110 vss.n109 4.6505
R651 vss.n66 vss.n65 4.6505
R652 vss.n72 vss.n71 4.6505
R653 vss.n78 vss.n77 4.6505
R654 vss.n84 vss.n83 4.6505
R655 vss.n90 vss.n89 4.6505
R656 vss.n96 vss.n95 4.6505
R657 vss.n102 vss.n101 4.6505
R658 vss.n108 vss.n107 4.6505
R659 vss.n121 vss.n120 4.6505
R660 vss.n60 vss.n59 4.6505
R661 vss.n718 vss.n715 4.3758
R662 vss.n768 vss.n558 4.37575
R663 vss.n821 vss.n397 4.37575
R664 vss.n878 vss.n236 4.37575
R665 vss.n154 vss.n153 4.14168
R666 vss.n315 vss.n314 4.14168
R667 vss.n476 vss.n475 4.14168
R668 vss.n694 vss.n693 4.14168
R669 vss.n166 vss.n165 3.38874
R670 vss.n327 vss.n326 3.38874
R671 vss.n488 vss.n487 3.38874
R672 vss.n706 vss.n705 3.38874
R673 vss.n241 vss.n240 3.37584
R674 vss.n402 vss.n401 3.37584
R675 vss.n889 vss.n887 3.2005
R676 vss.n247 vss.n246 3.2005
R677 vss.n408 vss.n407 3.2005
R678 vss.n565 vss.n564 3.2005
R679 vss.n146 vss.n142 3.16936
R680 vss.n307 vss.n303 3.16936
R681 vss.n468 vss.n464 3.16936
R682 vss.n686 vss.n682 3.16936
R683 vss.n171 vss.n166 3.01226
R684 vss.n332 vss.n327 3.01226
R685 vss.n493 vss.n488 3.01226
R686 vss.n711 vss.n706 3.01226
R687 vss.n728 vss.n727 2.9544
R688 vss.n827 vss.n248 2.89365
R689 vss.n774 vss.n409 2.89365
R690 vss.n724 vss.n566 2.89365
R691 vss.n717 vss.n716 2.83522
R692 vss.n132 vss.n131 2.83268
R693 vss vss.n899 2.60076
R694 vss.n148 vss.n139 2.26191
R695 vss.n309 vss.n300 2.26191
R696 vss.n470 vss.n461 2.26191
R697 vss.n688 vss.n679 2.26191
R698 vss.n159 vss.n154 2.25932
R699 vss.n320 vss.n315 2.25932
R700 vss.n481 vss.n476 2.25932
R701 vss.n699 vss.n694 2.25932
R702 vss.n56 vss.n53 1.91313
R703 vss.n139 vss.n138 1.73128
R704 vss.n300 vss.n299 1.73128
R705 vss.n461 vss.n460 1.73128
R706 vss.n679 vss.n678 1.73128
R707 vss.n841 vss.n840 1.6005
R708 vss.n788 vss.n787 1.6005
R709 vss.n735 vss.n734 1.6005
R710 vss.n58 vss.n56 1.50714
R711 vss.n147 vss.n141 1.50638
R712 vss.n308 vss.n302 1.50638
R713 vss.n469 vss.n463 1.50638
R714 vss.n687 vss.n681 1.50638
R715 vss.n889 vss.n888 1.14023
R716 vss.n248 vss.n247 1.14023
R717 vss.n409 vss.n408 1.14023
R718 vss.n566 vss.n565 1.14023
R719 vss.n138 vss.n42 0.753441
R720 vss.n299 vss.n291 0.753441
R721 vss.n460 vss.n452 0.753441
R722 vss.n678 vss.n670 0.753441
R723 vss.n120 vss.n119 0.747896
R724 vss.n119 vss.n117 0.69215
R725 vss.n899 vss.n898 0.690998
R726 vss.n238 vss.n237 0.658034
R727 vss.n399 vss.n398 0.658034
R728 vss.n884 vss.n883 0.614199
R729 vss.n243 vss.n242 0.614199
R730 vss.n404 vss.n403 0.614199
R731 vss.n561 vss.n560 0.614199
R732 vss.n158 vss.n157 0.514956
R733 vss.n319 vss.n318 0.514956
R734 vss.n480 vss.n479 0.514956
R735 vss.n698 vss.n697 0.514956
R736 vss.n876 vss.n875 0.438856
R737 vss.n240 vss.n239 0.438856
R738 vss.n401 vss.n400 0.438856
R739 vss.n887 vss.n884 0.219678
R740 vss.n246 vss.n243 0.219678
R741 vss.n407 vss.n404 0.219678
R742 vss.n564 vss.n561 0.219678
R743 vss.n137 vss.n136 0.178872
R744 vss.n298 vss.n297 0.178872
R745 vss.n459 vss.n458 0.178872
R746 vss.n677 vss.n676 0.178872
R747 vss.n172 vss.n164 0.144522
R748 vss.n160 vss.n152 0.144522
R749 vss.n333 vss.n325 0.144522
R750 vss.n321 vss.n313 0.144522
R751 vss.n494 vss.n486 0.144522
R752 vss.n482 vss.n474 0.144522
R753 vss.n712 vss.n704 0.144522
R754 vss.n700 vss.n692 0.144522
R755 vss.n883 vss.n882 0.132007
R756 vss.n242 vss.n241 0.132007
R757 vss.n403 vss.n402 0.132007
R758 vss.n560 vss.n559 0.132007
R759 vss.n723 vss.n722 0.120292
R760 vss.n729 vss.n726 0.120292
R761 vss.n731 vss.n729 0.120292
R762 vss.n733 vss.n731 0.120292
R763 vss.n736 vss.n733 0.120292
R764 vss.n738 vss.n736 0.120292
R765 vss.n740 vss.n738 0.120292
R766 vss.n742 vss.n740 0.120292
R767 vss.n744 vss.n742 0.120292
R768 vss.n746 vss.n744 0.120292
R769 vss.n748 vss.n746 0.120292
R770 vss.n750 vss.n748 0.120292
R771 vss.n752 vss.n750 0.120292
R772 vss.n754 vss.n752 0.120292
R773 vss.n756 vss.n754 0.120292
R774 vss.n758 vss.n756 0.120292
R775 vss.n760 vss.n758 0.120292
R776 vss.n762 vss.n760 0.120292
R777 vss.n764 vss.n762 0.120292
R778 vss.n773 vss.n772 0.120292
R779 vss.n782 vss.n778 0.120292
R780 vss.n784 vss.n782 0.120292
R781 vss.n786 vss.n784 0.120292
R782 vss.n789 vss.n786 0.120292
R783 vss.n791 vss.n789 0.120292
R784 vss.n793 vss.n791 0.120292
R785 vss.n795 vss.n793 0.120292
R786 vss.n797 vss.n795 0.120292
R787 vss.n799 vss.n797 0.120292
R788 vss.n801 vss.n799 0.120292
R789 vss.n803 vss.n801 0.120292
R790 vss.n805 vss.n803 0.120292
R791 vss.n807 vss.n805 0.120292
R792 vss.n809 vss.n807 0.120292
R793 vss.n811 vss.n809 0.120292
R794 vss.n813 vss.n811 0.120292
R795 vss.n815 vss.n813 0.120292
R796 vss.n817 vss.n815 0.120292
R797 vss.n826 vss.n825 0.120292
R798 vss.n835 vss.n831 0.120292
R799 vss.n837 vss.n835 0.120292
R800 vss.n839 vss.n837 0.120292
R801 vss.n842 vss.n839 0.120292
R802 vss.n844 vss.n842 0.120292
R803 vss.n846 vss.n844 0.120292
R804 vss.n848 vss.n846 0.120292
R805 vss.n850 vss.n848 0.120292
R806 vss.n852 vss.n850 0.120292
R807 vss.n854 vss.n852 0.120292
R808 vss.n856 vss.n854 0.120292
R809 vss.n858 vss.n856 0.120292
R810 vss.n860 vss.n858 0.120292
R811 vss.n862 vss.n860 0.120292
R812 vss.n864 vss.n862 0.120292
R813 vss.n866 vss.n864 0.120292
R814 vss.n868 vss.n866 0.120292
R815 vss.n870 vss.n868 0.120292
R816 vss.n891 vss.n890 0.120292
R817 vss.n60 vss.n58 0.120292
R818 vss.n62 vss.n60 0.120292
R819 vss.n64 vss.n62 0.120292
R820 vss.n66 vss.n64 0.120292
R821 vss.n68 vss.n66 0.120292
R822 vss.n70 vss.n68 0.120292
R823 vss.n72 vss.n70 0.120292
R824 vss.n74 vss.n72 0.120292
R825 vss.n76 vss.n74 0.120292
R826 vss.n78 vss.n76 0.120292
R827 vss.n80 vss.n78 0.120292
R828 vss.n82 vss.n80 0.120292
R829 vss.n84 vss.n82 0.120292
R830 vss.n86 vss.n84 0.120292
R831 vss.n88 vss.n86 0.120292
R832 vss.n90 vss.n88 0.120292
R833 vss.n92 vss.n90 0.120292
R834 vss.n94 vss.n92 0.120292
R835 vss.n96 vss.n94 0.120292
R836 vss.n98 vss.n96 0.120292
R837 vss.n100 vss.n98 0.120292
R838 vss.n102 vss.n100 0.120292
R839 vss.n104 vss.n102 0.120292
R840 vss.n106 vss.n104 0.120292
R841 vss.n108 vss.n106 0.120292
R842 vss.n110 vss.n108 0.120292
R843 vss.n111 vss.n110 0.120292
R844 vss.n120 vss.n111 0.120292
R845 vss.n718 vss.n717 0.109392
R846 vss.n722 vss.n721 0.102062
R847 vss.n772 vss.n771 0.102062
R848 vss.n825 vss.n824 0.102062
R849 vss.n890 vss.n881 0.102062
R850 vss.n765 vss.n764 0.10076
R851 vss.n818 vss.n817 0.10076
R852 vss.n872 vss.n870 0.10076
R853 vss.n112 vss 0.0887192
R854 vss.n876 vss.n874 0.0881712
R855 vss.n239 vss.n238 0.0881712
R856 vss.n400 vss.n399 0.0881712
R857 vss.n893 vss 0.075897
R858 vss.n723 vss 0.0603958
R859 vss.n726 vss 0.0603958
R860 vss.n773 vss 0.0603958
R861 vss.n778 vss 0.0603958
R862 vss.n826 vss 0.0603958
R863 vss.n831 vss 0.0603958
R864 vss vss.n891 0.0603958
R865 vss.n719 vss.n718 0.0590102
R866 vss.n769 vss.n768 0.0588433
R867 vss.n822 vss.n821 0.0588433
R868 vss.n879 vss.n878 0.0588433
R869 vss.n878 vss.n877 0.0577417
R870 vss.n821 vss.n820 0.0577417
R871 vss.n768 vss.n767 0.0577417
R872 vss.n152 vss.n150 0.0358261
R873 vss.n313 vss.n311 0.0358261
R874 vss.n474 vss.n472 0.0358261
R875 vss.n692 vss.n690 0.0358261
R876 vss.n119 vss.n118 0.0308571
R877 vss.n164 vss.n162 0.0303913
R878 vss.n325 vss.n323 0.0303913
R879 vss.n486 vss.n484 0.0303913
R880 vss.n704 vss.n702 0.0303913
R881 vss.n899 vss.n892 0.0272857
R882 vss.n236 vss.n174 0.0249565
R883 vss.n397 vss.n335 0.0249565
R884 vss.n558 vss.n496 0.0249565
R885 vss.n715 vss.n714 0.0249565
R886 vss.n898 vss.n897 0.0240572
R887 vss.n174 vss.n172 0.0222391
R888 vss.n335 vss.n333 0.0222391
R889 vss.n496 vss.n494 0.0222391
R890 vss.n714 vss.n712 0.0222391
R891 vss.n896 vss.n895 0.0205
R892 vss.n897 vss.n896 0.0205
R893 vss.n116 vss.n115 0.0205
R894 vss.n115 vss.n114 0.0205
R895 vss.n766 vss.n765 0.0200312
R896 vss.n819 vss.n818 0.0200312
R897 vss.n873 vss.n872 0.0200312
R898 vss.n117 vss.n116 0.0187452
R899 vss.n721 vss.n720 0.0187292
R900 vss.n771 vss.n770 0.0187292
R901 vss.n824 vss.n823 0.0187292
R902 vss.n881 vss.n880 0.0187292
R903 vss.n162 vss.n160 0.0168043
R904 vss.n323 vss.n321 0.0168043
R905 vss.n484 vss.n482 0.0168043
R906 vss.n702 vss.n700 0.0168043
R907 vss.n898 vss.n894 0.0163636
R908 vss.n117 vss.n113 0.0142271
R909 vss.n113 vss.n112 0.0121722
R910 vss.n894 vss.n893 0.011753
R911 vss.n150 vss.n148 0.0113696
R912 vss.n311 vss.n309 0.0113696
R913 vss.n472 vss.n470 0.0113696
R914 vss.n690 vss.n688 0.0113696
R915 vss.n720 vss.n719 0.00440625
R916 vss.n770 vss.n769 0.00440625
R917 vss.n823 vss.n822 0.00440625
R918 vss.n880 vss.n879 0.00440625
R919 vss.n767 vss.n766 0.00310417
R920 vss.n820 vss.n819 0.00310417
R921 vss.n877 vss.n873 0.00310417
R922 ctl6.n0 ctl6.t2 212.081
R923 ctl6.n1 ctl6.t3 212.081
R924 ctl6.n0 ctl6.t0 139.78
R925 ctl6.n1 ctl6.t1 139.78
R926 ctl6.n1 ctl6.n0 61.346
R927 ctl6 ctl6.n1 44.6884
R928 dum.n0 dum.t2 212.081
R929 dum.n1 dum.t3 212.081
R930 dum.n0 dum.t0 139.78
R931 dum.n1 dum.t1 139.78
R932 dum.n1 dum.n0 61.346
R933 dum dum.n1 44.6494
R934 ctl0.n0 ctl0.t2 212.081
R935 ctl0.n1 ctl0.t3 212.081
R936 ctl0.n0 ctl0.t0 139.78
R937 ctl0.n1 ctl0.t1 139.78
R938 ctl0.n1 ctl0.n0 61.346
R939 ctl0 ctl0.n1 44.6884
R940 ctl1.n0 ctl1.t2 212.081
R941 ctl1.n1 ctl1.t3 212.081
R942 ctl1.n0 ctl1.t0 139.78
R943 ctl1.n1 ctl1.t1 139.78
R944 ctl1.n1 ctl1.n0 61.346
R945 ctl1 ctl1.n1 44.6884
R946 ctl5.n0 ctl5.t2 212.081
R947 ctl5.n1 ctl5.t3 212.081
R948 ctl5.n0 ctl5.t0 139.78
R949 ctl5.n1 ctl5.t1 139.78
R950 ctl5.n1 ctl5.n0 61.346
R951 ctl5 ctl5.n1 44.6884
R952 ctl4.n0 ctl4.t2 212.081
R953 ctl4.n1 ctl4.t3 212.081
R954 ctl4.n0 ctl4.t0 139.78
R955 ctl4.n1 ctl4.t1 139.78
R956 ctl4.n1 ctl4.n0 61.346
R957 ctl4 ctl4.n1 44.6884
R958 ctl2.n0 ctl2.t2 212.081
R959 ctl2.n1 ctl2.t3 212.081
R960 ctl2.n0 ctl2.t0 139.78
R961 ctl2.n1 ctl2.t1 139.78
R962 ctl2.n1 ctl2.n0 61.346
R963 ctl2 ctl2.n1 44.6884
R964 ctl3.n0 ctl3.t2 212.081
R965 ctl3.n1 ctl3.t3 212.081
R966 ctl3.n0 ctl3.t0 139.78
R967 ctl3.n1 ctl3.t1 139.78
R968 ctl3.n1 ctl3.n0 61.346
R969 ctl3 ctl3.n1 44.6884
R970 out.n23 out.n13 1.72892
R971 out.n18 out.n17 1.7055
R972 out.n48 out.n47 1.7055
R973 out.n71 out.n70 1.7055
R974 out.n6 out.n5 1.7055
R975 out.n9 out.n0 1.7055
R976 out.n67 out.n63 1.7055
R977 out.n44 out.n40 1.7055
R978 out.n22 out.n21 1.7055
R979 out.n76 out.n75 1.09861
R980 out.n53 out.n52 1.09651
R981 out.n30 out.n29 1.09651
R982 out.n52 out.n51 0.680902
R983 out.n75 out.n74 0.680902
R984 out.n85 out.n12 0.680902
R985 out.n425 out.n424 0.6115
R986 out.n424 out.n423 0.6115
R987 out.n423 out.n422 0.6115
R988 out.n422 out.n421 0.6115
R989 out.n421 out.n420 0.6115
R990 out.n420 out.n419 0.6115
R991 out.n419 out.n418 0.6115
R992 out.n418 out.n417 0.6115
R993 out.n417 out.n416 0.6115
R994 out.n416 out.n415 0.6115
R995 out.n415 out.n414 0.6115
R996 out.n414 out.n413 0.6115
R997 out.n413 out.n412 0.6115
R998 out.n412 out.n411 0.6115
R999 out.n411 out.n410 0.6115
R1000 out.n410 out.n409 0.6115
R1001 out.n409 out.n408 0.6115
R1002 out.n408 out.n407 0.6115
R1003 out.n407 out.n406 0.6115
R1004 out.n406 out.n405 0.6115
R1005 out.n405 out.n404 0.6115
R1006 out.n404 out.n403 0.6115
R1007 out.n403 out.n402 0.6115
R1008 out.n402 out.n401 0.6115
R1009 out.n401 out.n400 0.6115
R1010 out.n400 out.n399 0.6115
R1011 out.n399 out.n398 0.6115
R1012 out.n398 out.n397 0.6115
R1013 out.n397 out.n396 0.6115
R1014 out.n396 out.n395 0.6115
R1015 out.n395 out.n394 0.6115
R1016 out.n394 out.n393 0.6115
R1017 out.n393 out.n392 0.6115
R1018 out out.n85 0.512552
R1019 out.n24 out.n23 0.331771
R1020 out.n383 out.t123 0.301104
R1021 out.n374 out.t143 0.301104
R1022 out.n365 out.t162 0.301104
R1023 out.n356 out.t176 0.301104
R1024 out.n347 out.t235 0.301104
R1025 out.n338 out.t194 0.301104
R1026 out.n329 out.t209 0.301104
R1027 out.n320 out.t103 0.301104
R1028 out.n311 out.t66 0.301104
R1029 out.n302 out.t127 0.301104
R1030 out.n293 out.t146 0.301104
R1031 out.n284 out.t164 0.301104
R1032 out.n275 out.t180 0.301104
R1033 out.n266 out.t56 0.301104
R1034 out.n257 out.t72 0.301104
R1035 out.n248 out.t89 0.301104
R1036 out.n239 out.t108 0.301104
R1037 out.n230 out.t161 0.301104
R1038 out.n221 out.t179 0.301104
R1039 out.n212 out.t192 0.301104
R1040 out.n203 out.t142 0.301104
R1041 out.n194 out.t23 0.301104
R1042 out.n185 out.t84 0.301104
R1043 out.n176 out.t122 0.301104
R1044 out.n167 out.t102 0.301104
R1045 out.n158 out.t22 0.301104
R1046 out.n149 out.t160 0.301104
R1047 out.n140 out.t178 0.301104
R1048 out.n131 out.t191 0.301104
R1049 out.n122 out.t65 0.301104
R1050 out.n113 out.t121 0.301104
R1051 out.n104 out.t141 0.301104
R1052 out.n95 out.t83 0.301104
R1053 out.n86 out.t101 0.301104
R1054 out.n384 out.n383 0.301104
R1055 out.n385 out.n384 0.301104
R1056 out.n386 out.n385 0.301104
R1057 out.n387 out.n386 0.301104
R1058 out.n388 out.n387 0.301104
R1059 out.n389 out.n388 0.301104
R1060 out.n390 out.n389 0.301104
R1061 out.n391 out.n390 0.301104
R1062 out.n375 out.n374 0.301104
R1063 out.n376 out.n375 0.301104
R1064 out.n377 out.n376 0.301104
R1065 out.n378 out.n377 0.301104
R1066 out.n379 out.n378 0.301104
R1067 out.n380 out.n379 0.301104
R1068 out.n381 out.n380 0.301104
R1069 out.n382 out.n381 0.301104
R1070 out.n366 out.n365 0.301104
R1071 out.n367 out.n366 0.301104
R1072 out.n368 out.n367 0.301104
R1073 out.n369 out.n368 0.301104
R1074 out.n370 out.n369 0.301104
R1075 out.n371 out.n370 0.301104
R1076 out.n372 out.n371 0.301104
R1077 out.n373 out.n372 0.301104
R1078 out.n357 out.n356 0.301104
R1079 out.n358 out.n357 0.301104
R1080 out.n359 out.n358 0.301104
R1081 out.n360 out.n359 0.301104
R1082 out.n361 out.n360 0.301104
R1083 out.n362 out.n361 0.301104
R1084 out.n363 out.n362 0.301104
R1085 out.n364 out.n363 0.301104
R1086 out.n348 out.n347 0.301104
R1087 out.n349 out.n348 0.301104
R1088 out.n350 out.n349 0.301104
R1089 out.n351 out.n350 0.301104
R1090 out.n352 out.n351 0.301104
R1091 out.n353 out.n352 0.301104
R1092 out.n354 out.n353 0.301104
R1093 out.n355 out.n354 0.301104
R1094 out.n339 out.n338 0.301104
R1095 out.n340 out.n339 0.301104
R1096 out.n341 out.n340 0.301104
R1097 out.n342 out.n341 0.301104
R1098 out.n343 out.n342 0.301104
R1099 out.n344 out.n343 0.301104
R1100 out.n345 out.n344 0.301104
R1101 out.n346 out.n345 0.301104
R1102 out.n330 out.n329 0.301104
R1103 out.n331 out.n330 0.301104
R1104 out.n332 out.n331 0.301104
R1105 out.n333 out.n332 0.301104
R1106 out.n334 out.n333 0.301104
R1107 out.n335 out.n334 0.301104
R1108 out.n336 out.n335 0.301104
R1109 out.n337 out.n336 0.301104
R1110 out.n321 out.n320 0.301104
R1111 out.n322 out.n321 0.301104
R1112 out.n323 out.n322 0.301104
R1113 out.n324 out.n323 0.301104
R1114 out.n325 out.n324 0.301104
R1115 out.n326 out.n325 0.301104
R1116 out.n327 out.n326 0.301104
R1117 out.n328 out.n327 0.301104
R1118 out.n312 out.n311 0.301104
R1119 out.n313 out.n312 0.301104
R1120 out.n314 out.n313 0.301104
R1121 out.n315 out.n314 0.301104
R1122 out.n316 out.n315 0.301104
R1123 out.n317 out.n316 0.301104
R1124 out.n318 out.n317 0.301104
R1125 out.n319 out.n318 0.301104
R1126 out.n303 out.n302 0.301104
R1127 out.n304 out.n303 0.301104
R1128 out.n305 out.n304 0.301104
R1129 out.n306 out.n305 0.301104
R1130 out.n307 out.n306 0.301104
R1131 out.n308 out.n307 0.301104
R1132 out.n309 out.n308 0.301104
R1133 out.n310 out.n309 0.301104
R1134 out.n294 out.n293 0.301104
R1135 out.n295 out.n294 0.301104
R1136 out.n296 out.n295 0.301104
R1137 out.n297 out.n296 0.301104
R1138 out.n298 out.n297 0.301104
R1139 out.n299 out.n298 0.301104
R1140 out.n300 out.n299 0.301104
R1141 out.n301 out.n300 0.301104
R1142 out.n285 out.n284 0.301104
R1143 out.n286 out.n285 0.301104
R1144 out.n287 out.n286 0.301104
R1145 out.n288 out.n287 0.301104
R1146 out.n289 out.n288 0.301104
R1147 out.n290 out.n289 0.301104
R1148 out.n291 out.n290 0.301104
R1149 out.n292 out.n291 0.301104
R1150 out.n276 out.n275 0.301104
R1151 out.n277 out.n276 0.301104
R1152 out.n278 out.n277 0.301104
R1153 out.n279 out.n278 0.301104
R1154 out.n280 out.n279 0.301104
R1155 out.n281 out.n280 0.301104
R1156 out.n282 out.n281 0.301104
R1157 out.n283 out.n282 0.301104
R1158 out.n267 out.n266 0.301104
R1159 out.n268 out.n267 0.301104
R1160 out.n269 out.n268 0.301104
R1161 out.n270 out.n269 0.301104
R1162 out.n271 out.n270 0.301104
R1163 out.n272 out.n271 0.301104
R1164 out.n273 out.n272 0.301104
R1165 out.n274 out.n273 0.301104
R1166 out.n258 out.n257 0.301104
R1167 out.n259 out.n258 0.301104
R1168 out.n260 out.n259 0.301104
R1169 out.n261 out.n260 0.301104
R1170 out.n262 out.n261 0.301104
R1171 out.n263 out.n262 0.301104
R1172 out.n264 out.n263 0.301104
R1173 out.n265 out.n264 0.301104
R1174 out.n249 out.n248 0.301104
R1175 out.n250 out.n249 0.301104
R1176 out.n251 out.n250 0.301104
R1177 out.n252 out.n251 0.301104
R1178 out.n253 out.n252 0.301104
R1179 out.n254 out.n253 0.301104
R1180 out.n255 out.n254 0.301104
R1181 out.n256 out.n255 0.301104
R1182 out.n240 out.n239 0.301104
R1183 out.n241 out.n240 0.301104
R1184 out.n242 out.n241 0.301104
R1185 out.n243 out.n242 0.301104
R1186 out.n244 out.n243 0.301104
R1187 out.n245 out.n244 0.301104
R1188 out.n246 out.n245 0.301104
R1189 out.n247 out.n246 0.301104
R1190 out.n231 out.n230 0.301104
R1191 out.n232 out.n231 0.301104
R1192 out.n233 out.n232 0.301104
R1193 out.n234 out.n233 0.301104
R1194 out.n235 out.n234 0.301104
R1195 out.n236 out.n235 0.301104
R1196 out.n237 out.n236 0.301104
R1197 out.n238 out.n237 0.301104
R1198 out.n222 out.n221 0.301104
R1199 out.n223 out.n222 0.301104
R1200 out.n224 out.n223 0.301104
R1201 out.n225 out.n224 0.301104
R1202 out.n226 out.n225 0.301104
R1203 out.n227 out.n226 0.301104
R1204 out.n228 out.n227 0.301104
R1205 out.n229 out.n228 0.301104
R1206 out.n213 out.n212 0.301104
R1207 out.n214 out.n213 0.301104
R1208 out.n215 out.n214 0.301104
R1209 out.n216 out.n215 0.301104
R1210 out.n217 out.n216 0.301104
R1211 out.n218 out.n217 0.301104
R1212 out.n219 out.n218 0.301104
R1213 out.n220 out.n219 0.301104
R1214 out.n204 out.n203 0.301104
R1215 out.n205 out.n204 0.301104
R1216 out.n206 out.n205 0.301104
R1217 out.n207 out.n206 0.301104
R1218 out.n208 out.n207 0.301104
R1219 out.n209 out.n208 0.301104
R1220 out.n210 out.n209 0.301104
R1221 out.n211 out.n210 0.301104
R1222 out.n195 out.n194 0.301104
R1223 out.n196 out.n195 0.301104
R1224 out.n197 out.n196 0.301104
R1225 out.n198 out.n197 0.301104
R1226 out.n199 out.n198 0.301104
R1227 out.n200 out.n199 0.301104
R1228 out.n201 out.n200 0.301104
R1229 out.n202 out.n201 0.301104
R1230 out.n186 out.n185 0.301104
R1231 out.n187 out.n186 0.301104
R1232 out.n188 out.n187 0.301104
R1233 out.n189 out.n188 0.301104
R1234 out.n190 out.n189 0.301104
R1235 out.n191 out.n190 0.301104
R1236 out.n192 out.n191 0.301104
R1237 out.n193 out.n192 0.301104
R1238 out.n177 out.n176 0.301104
R1239 out.n178 out.n177 0.301104
R1240 out.n179 out.n178 0.301104
R1241 out.n180 out.n179 0.301104
R1242 out.n181 out.n180 0.301104
R1243 out.n182 out.n181 0.301104
R1244 out.n183 out.n182 0.301104
R1245 out.n184 out.n183 0.301104
R1246 out.n168 out.n167 0.301104
R1247 out.n169 out.n168 0.301104
R1248 out.n170 out.n169 0.301104
R1249 out.n171 out.n170 0.301104
R1250 out.n172 out.n171 0.301104
R1251 out.n173 out.n172 0.301104
R1252 out.n174 out.n173 0.301104
R1253 out.n175 out.n174 0.301104
R1254 out.n159 out.n158 0.301104
R1255 out.n160 out.n159 0.301104
R1256 out.n161 out.n160 0.301104
R1257 out.n162 out.n161 0.301104
R1258 out.n163 out.n162 0.301104
R1259 out.n164 out.n163 0.301104
R1260 out.n165 out.n164 0.301104
R1261 out.n166 out.n165 0.301104
R1262 out.n150 out.n149 0.301104
R1263 out.n151 out.n150 0.301104
R1264 out.n152 out.n151 0.301104
R1265 out.n153 out.n152 0.301104
R1266 out.n154 out.n153 0.301104
R1267 out.n155 out.n154 0.301104
R1268 out.n156 out.n155 0.301104
R1269 out.n157 out.n156 0.301104
R1270 out.n141 out.n140 0.301104
R1271 out.n142 out.n141 0.301104
R1272 out.n143 out.n142 0.301104
R1273 out.n144 out.n143 0.301104
R1274 out.n145 out.n144 0.301104
R1275 out.n146 out.n145 0.301104
R1276 out.n147 out.n146 0.301104
R1277 out.n148 out.n147 0.301104
R1278 out.n132 out.n131 0.301104
R1279 out.n133 out.n132 0.301104
R1280 out.n134 out.n133 0.301104
R1281 out.n135 out.n134 0.301104
R1282 out.n136 out.n135 0.301104
R1283 out.n137 out.n136 0.301104
R1284 out.n138 out.n137 0.301104
R1285 out.n139 out.n138 0.301104
R1286 out.n123 out.n122 0.301104
R1287 out.n124 out.n123 0.301104
R1288 out.n125 out.n124 0.301104
R1289 out.n126 out.n125 0.301104
R1290 out.n127 out.n126 0.301104
R1291 out.n128 out.n127 0.301104
R1292 out.n129 out.n128 0.301104
R1293 out.n130 out.n129 0.301104
R1294 out.n114 out.n113 0.301104
R1295 out.n115 out.n114 0.301104
R1296 out.n116 out.n115 0.301104
R1297 out.n117 out.n116 0.301104
R1298 out.n118 out.n117 0.301104
R1299 out.n119 out.n118 0.301104
R1300 out.n120 out.n119 0.301104
R1301 out.n121 out.n120 0.301104
R1302 out.n105 out.n104 0.301104
R1303 out.n106 out.n105 0.301104
R1304 out.n107 out.n106 0.301104
R1305 out.n108 out.n107 0.301104
R1306 out.n109 out.n108 0.301104
R1307 out.n110 out.n109 0.301104
R1308 out.n111 out.n110 0.301104
R1309 out.n112 out.n111 0.301104
R1310 out.n96 out.n95 0.301104
R1311 out.n97 out.n96 0.301104
R1312 out.n98 out.n97 0.301104
R1313 out.n99 out.n98 0.301104
R1314 out.n100 out.n99 0.301104
R1315 out.n101 out.n100 0.301104
R1316 out.n102 out.n101 0.301104
R1317 out.n103 out.n102 0.301104
R1318 out.n87 out.n86 0.301104
R1319 out.n88 out.n87 0.301104
R1320 out.n89 out.n88 0.301104
R1321 out.n90 out.n89 0.301104
R1322 out.n91 out.n90 0.301104
R1323 out.n92 out.n91 0.301104
R1324 out.n93 out.n92 0.301104
R1325 out.n94 out.n93 0.301104
R1326 out out.n425 0.165
R1327 out.n392 out.n391 0.14101
R1328 out.n393 out.n382 0.14101
R1329 out.n394 out.n373 0.14101
R1330 out.n395 out.n364 0.14101
R1331 out.n396 out.n355 0.14101
R1332 out.n397 out.n346 0.14101
R1333 out.n398 out.n337 0.14101
R1334 out.n399 out.n328 0.14101
R1335 out.n400 out.n319 0.14101
R1336 out.n401 out.n310 0.14101
R1337 out.n402 out.n301 0.14101
R1338 out.n403 out.n292 0.14101
R1339 out.n404 out.n283 0.14101
R1340 out.n405 out.n274 0.14101
R1341 out.n406 out.n265 0.14101
R1342 out.n407 out.n256 0.14101
R1343 out.n408 out.n247 0.14101
R1344 out.n409 out.n238 0.14101
R1345 out.n410 out.n229 0.14101
R1346 out.n411 out.n220 0.14101
R1347 out.n412 out.n211 0.14101
R1348 out.n413 out.n202 0.14101
R1349 out.n414 out.n193 0.14101
R1350 out.n415 out.n184 0.14101
R1351 out.n416 out.n175 0.14101
R1352 out.n417 out.n166 0.14101
R1353 out.n418 out.n157 0.14101
R1354 out.n419 out.n148 0.14101
R1355 out.n420 out.n139 0.14101
R1356 out.n421 out.n130 0.14101
R1357 out.n422 out.n121 0.14101
R1358 out.n423 out.n112 0.14101
R1359 out.n424 out.n103 0.14101
R1360 out.n425 out.n94 0.14101
R1361 out.n13 out 0.0505
R1362 out.n39 out 0.0505
R1363 out.n62 out 0.0505
R1364 out.n4 out 0.0505
R1365 out.n40 out.n39 0.03175
R1366 out.n63 out.n62 0.03175
R1367 out.n5 out.n4 0.03175
R1368 out.n23 out.n22 0.025645
R1369 out.n392 out 0.02306
R1370 out.n77 out.n76 0.023016
R1371 out.n85 out.n84 0.0221211
R1372 out.n54 out.n53 0.0221211
R1373 out.n31 out.n30 0.0221211
R1374 out.n75 out.n61 0.0221211
R1375 out.n52 out.n38 0.0221211
R1376 out.n29 out.n28 0.0221211
R1377 out.n15 out.n14 0.018125
R1378 out.n18 out.n16 0.018125
R1379 out.n19 out.n18 0.018125
R1380 out.n22 out.n20 0.018125
R1381 out.n51 out.n50 0.018125
R1382 out.n49 out.n48 0.018125
R1383 out.n48 out.n46 0.018125
R1384 out.n45 out.n44 0.018125
R1385 out.n44 out.n43 0.018125
R1386 out.n42 out.n41 0.018125
R1387 out.n74 out.n73 0.018125
R1388 out.n72 out.n71 0.018125
R1389 out.n71 out.n69 0.018125
R1390 out.n68 out.n67 0.018125
R1391 out.n67 out.n66 0.018125
R1392 out.n65 out.n64 0.018125
R1393 out.n12 out.n11 0.018125
R1394 out.n10 out.n9 0.018125
R1395 out.n9 out.n8 0.018125
R1396 out.n7 out.n6 0.018125
R1397 out.n6 out.n3 0.018125
R1398 out.n2 out.n1 0.018125
R1399 out.n83 out.n82 0.018125
R1400 out.n82 out.n81 0.018125
R1401 out.n80 out.n79 0.018125
R1402 out.n79 out.n78 0.018125
R1403 out.n60 out.n59 0.018125
R1404 out.n59 out.n58 0.018125
R1405 out.n57 out.n56 0.018125
R1406 out.n56 out.n55 0.018125
R1407 out.n37 out.n36 0.018125
R1408 out.n36 out.n35 0.018125
R1409 out.n34 out.n33 0.018125
R1410 out.n33 out.n32 0.018125
R1411 out.n27 out.n26 0.018125
R1412 out.n26 out.n25 0.018125
R1413 out.n16 out.n15 0.01225
R1414 out.n20 out.n19 0.01225
R1415 out.n50 out.n49 0.01225
R1416 out.n46 out.n45 0.01225
R1417 out.n43 out.n42 0.01225
R1418 out.n73 out.n72 0.01225
R1419 out.n69 out.n68 0.01225
R1420 out.n66 out.n65 0.01225
R1421 out.n11 out.n10 0.01225
R1422 out.n8 out.n7 0.01225
R1423 out.n3 out.n2 0.01225
R1424 out.n84 out.n83 0.01225
R1425 out.n81 out.n80 0.01225
R1426 out.n78 out.n77 0.01225
R1427 out.n61 out.n60 0.01225
R1428 out.n58 out.n57 0.01225
R1429 out.n55 out.n54 0.01225
R1430 out.n38 out.n37 0.01225
R1431 out.n35 out.n34 0.01225
R1432 out.n32 out.n31 0.01225
R1433 out.n28 out.n27 0.01225
R1434 out.n25 out.n24 0.01225
R1435 out.n383 out.t223 0.00050016
R1436 out.n384 out.t193 0.00050016
R1437 out.n385 out.t207 0.00050016
R1438 out.n386 out.t79 0.00050016
R1439 out.n387 out.t245 0.00050016
R1440 out.n388 out.t100 0.00050016
R1441 out.n389 out.t140 0.00050016
R1442 out.n390 out.t119 0.00050016
R1443 out.n391 out.t175 0.00050016
R1444 out.n374 out.t240 0.00050016
R1445 out.n375 out.t230 0.00050016
R1446 out.n376 out.t250 0.00050016
R1447 out.n377 out.t198 0.00050016
R1448 out.n378 out.t213 0.00050016
R1449 out.n379 out.t238 0.00050016
R1450 out.n380 out.t268 0.00050016
R1451 out.n381 out.t254 0.00050016
R1452 out.n382 out.t159 0.00050016
R1453 out.n365 out.t152 0.00050016
R1454 out.n366 out.t112 0.00050016
R1455 out.n367 out.t132 0.00050016
R1456 out.n368 out.t86 0.00050016
R1457 out.n369 out.t125 0.00050016
R1458 out.n370 out.t105 0.00050016
R1459 out.n371 out.t163 0.00050016
R1460 out.n372 out.t144 0.00050016
R1461 out.n373 out.t190 0.00050016
R1462 out.n356 out.t258 0.00050016
R1463 out.n357 out.t216 0.00050016
R1464 out.n358 out.t302 0.00050016
R1465 out.n359 out.t185 0.00050016
R1466 out.n360 out.t249 0.00050016
R1467 out.n361 out.t225 0.00050016
R1468 out.n362 out.t273 0.00050016
R1469 out.n363 out.t262 0.00050016
R1470 out.n364 out.t206 0.00050016
R1471 out.n347 out.t241 0.00050016
R1472 out.n348 out.t217 0.00050016
R1473 out.n349 out.t232 0.00050016
R1474 out.n350 out.t228 0.00050016
R1475 out.n351 out.t265 0.00050016
R1476 out.n352 out.t256 0.00050016
R1477 out.n353 out.t246 0.00050016
R1478 out.n354 out.t236 0.00050016
R1479 out.n355 out.t81 0.00050016
R1480 out.n338 out.t13 0.00050016
R1481 out.n339 out.t27 0.00050016
R1482 out.n340 out.t171 0.00050016
R1483 out.n341 out.t54 0.00050016
R1484 out.n342 out.t68 0.00050016
R1485 out.n343 out.t38 0.00050016
R1486 out.n344 out.t12 0.00050016
R1487 out.n345 out.t3 0.00050016
R1488 out.n346 out.t222 0.00050016
R1489 out.n329 out.t279 0.00050016
R1490 out.n330 out.t200 0.00050016
R1491 out.n331 out.t271 0.00050016
R1492 out.n332 out.t278 0.00050016
R1493 out.n333 out.t257 0.00050016
R1494 out.n334 out.t269 0.00050016
R1495 out.n335 out.t211 0.00050016
R1496 out.n336 out.t181 0.00050016
R1497 out.n337 out.t234 0.00050016
R1498 out.n320 out.t275 0.00050016
R1499 out.n321 out.t282 0.00050016
R1500 out.n322 out.t266 0.00050016
R1501 out.n323 out.t274 0.00050016
R1502 out.n324 out.t248 0.00050016
R1503 out.n325 out.t264 0.00050016
R1504 out.n326 out.t196 0.00050016
R1505 out.n327 out.t166 0.00050016
R1506 out.n328 out.t64 0.00050016
R1507 out.n311 out.t313 0.00050016
R1508 out.n312 out.t308 0.00050016
R1509 out.n313 out.t303 0.00050016
R1510 out.n314 out.t316 0.00050016
R1511 out.n315 out.t314 0.00050016
R1512 out.n316 out.t318 0.00050016
R1513 out.n317 out.t291 0.00050016
R1514 out.n318 out.t297 0.00050016
R1515 out.n319 out.t49 0.00050016
R1516 out.n302 out.t42 0.00050016
R1517 out.n303 out.t17 0.00050016
R1518 out.n304 out.t29 0.00050016
R1519 out.n305 out.t70 0.00050016
R1520 out.n306 out.t85 0.00050016
R1521 out.n307 out.t104 0.00050016
R1522 out.n308 out.t145 0.00050016
R1523 out.n309 out.t124 0.00050016
R1524 out.n310 out.t99 0.00050016
R1525 out.n293 out.t284 0.00050016
R1526 out.n294 out.t267 0.00050016
R1527 out.n295 out.t276 0.00050016
R1528 out.n296 out.t197 0.00050016
R1529 out.n297 out.t227 0.00050016
R1530 out.n298 out.t247 0.00050016
R1531 out.n299 out.t263 0.00050016
R1532 out.n300 out.t128 0.00050016
R1533 out.n301 out.t118 0.00050016
R1534 out.n284 out.t280 0.00050016
R1535 out.n285 out.t261 0.00050016
R1536 out.n286 out.t272 0.00050016
R1537 out.n287 out.t184 0.00050016
R1538 out.n288 out.t212 0.00050016
R1539 out.n289 out.t237 0.00050016
R1540 out.n290 out.t255 0.00050016
R1541 out.n291 out.t147 0.00050016
R1542 out.n292 out.t139 0.00050016
R1543 out.n275 out.t281 0.00050016
R1544 out.n276 out.t277 0.00050016
R1545 out.n277 out.t285 0.00050016
R1546 out.n278 out.t299 0.00050016
R1547 out.n279 out.t309 0.00050016
R1548 out.n280 out.t304 0.00050016
R1549 out.n281 out.t294 0.00050016
R1550 out.n282 out.t289 0.00050016
R1551 out.n283 out.t221 0.00050016
R1552 out.n266 out.t57 0.00050016
R1553 out.n267 out.t74 0.00050016
R1554 out.n268 out.t93 0.00050016
R1555 out.n269 out.t40 0.00050016
R1556 out.n270 out.t25 0.00050016
R1557 out.n271 out.t52 0.00050016
R1558 out.n272 out.t5 0.00050016
R1559 out.n273 out.t338 0.00050016
R1560 out.n274 out.t189 0.00050016
R1561 out.n257 out.t288 0.00050016
R1562 out.n258 out.t293 0.00050016
R1563 out.n259 out.t298 0.00050016
R1564 out.n260 out.t270 0.00050016
R1565 out.n261 out.t168 0.00050016
R1566 out.n262 out.t149 0.00050016
R1567 out.n263 out.t182 0.00050016
R1568 out.n264 out.t165 0.00050016
R1569 out.n265 out.t205 0.00050016
R1570 out.n248 out.t58 0.00050016
R1571 out.n249 out.t75 0.00050016
R1572 out.n250 out.t94 0.00050016
R1573 out.n251 out.t133 0.00050016
R1574 out.n252 out.t113 0.00050016
R1575 out.n253 out.t153 0.00050016
R1576 out.n254 out.t172 0.00050016
R1577 out.n255 out.t188 0.00050016
R1578 out.n256 out.t158 0.00050016
R1579 out.n239 out.t295 0.00050016
R1580 out.n240 out.t290 0.00050016
R1581 out.n241 out.t116 0.00050016
R1582 out.n242 out.t306 0.00050016
R1583 out.n243 out.t323 0.00050016
R1584 out.n244 out.t136 0.00050016
R1585 out.n245 out.t300 0.00050016
R1586 out.n246 out.t305 0.00050016
R1587 out.n247 out.t174 0.00050016
R1588 out.n230 out.t310 0.00050016
R1589 out.n231 out.t315 0.00050016
R1590 out.n232 out.t155 0.00050016
R1591 out.n233 out.t43 0.00050016
R1592 out.n234 out.t311 0.00050016
R1593 out.n235 out.t173 0.00050016
R1594 out.n236 out.t322 0.00050016
R1595 out.n237 out.t319 0.00050016
R1596 out.n238 out.t80 0.00050016
R1597 out.n221 out.t220 0.00050016
R1598 out.n222 out.t203 0.00050016
R1599 out.n223 out.t204 0.00050016
R1600 out.n224 out.t219 0.00050016
R1601 out.n225 out.t233 0.00050016
R1602 out.n226 out.t244 0.00050016
R1603 out.n227 out.t260 0.00050016
R1604 out.n228 out.t253 0.00050016
R1605 out.n229 out.t35 0.00050016
R1606 out.n212 out.t92 0.00050016
R1607 out.n213 out.t110 0.00050016
R1608 out.n214 out.t251 0.00050016
R1609 out.n215 out.t183 0.00050016
R1610 out.n216 out.t167 0.00050016
R1611 out.n217 out.t148 0.00050016
R1612 out.n218 out.t210 0.00050016
R1613 out.n219 out.t195 0.00050016
R1614 out.n220 out.t48 0.00050016
R1615 out.n203 out.t126 0.00050016
R1616 out.n204 out.t334 0.00050016
R1617 out.n205 out.t107 0.00050016
R1618 out.n206 out.t106 0.00050016
R1619 out.n207 out.t88 0.00050016
R1620 out.n208 out.t67 0.00050016
R1621 out.n209 out.t330 0.00050016
R1622 out.n210 out.t332 0.00050016
R1623 out.n211 out.t63 0.00050016
R1624 out.n194 out.t325 0.00050016
R1625 out.n195 out.t320 0.00050016
R1626 out.n196 out.t328 0.00050016
R1627 out.n197 out.t301 0.00050016
R1628 out.n198 out.t287 0.00050016
R1629 out.n199 out.t292 0.00050016
R1630 out.n200 out.t331 0.00050016
R1631 out.n201 out.t296 0.00050016
R1632 out.n202 out.t157 0.00050016
R1633 out.n185 out.t214 0.00050016
R1634 out.n186 out.t130 0.00050016
R1635 out.n187 out.t170 0.00050016
R1636 out.n188 out.t129 0.00050016
R1637 out.n189 out.t239 0.00050016
R1638 out.n190 out.t91 0.00050016
R1639 out.n191 out.t31 0.00050016
R1640 out.n192 out.t8 0.00050016
R1641 out.n193 out.t138 0.00050016
R1642 out.n176 out.t199 0.00050016
R1643 out.n177 out.t187 0.00050016
R1644 out.n178 out.t151 0.00050016
R1645 out.n179 out.t109 0.00050016
R1646 out.n180 out.t226 0.00050016
R1647 out.n181 out.t73 0.00050016
R1648 out.n182 out.t19 0.00050016
R1649 out.n183 out.t224 0.00050016
R1650 out.n184 out.t98 0.00050016
R1651 out.n167 out.t6 0.00050016
R1652 out.n168 out.t16 0.00050016
R1653 out.n169 out.t339 0.00050016
R1654 out.n170 out.t39 0.00050016
R1655 out.n171 out.t53 0.00050016
R1656 out.n172 out.t24 0.00050016
R1657 out.n173 out.t4 0.00050016
R1658 out.n174 out.t337 0.00050016
R1659 out.n175 out.t117 0.00050016
R1660 out.n158 out.t327 0.00050016
R1661 out.n159 out.t321 0.00050016
R1662 out.n160 out.t317 0.00050016
R1663 out.n161 out.t324 0.00050016
R1664 out.n162 out.t312 0.00050016
R1665 out.n163 out.t307 0.00050016
R1666 out.n164 out.t286 0.00050016
R1667 out.n165 out.t283 0.00050016
R1668 out.n166 out.t34 0.00050016
R1669 out.n149 out.t215 0.00050016
R1670 out.n150 out.t259 0.00050016
R1671 out.n151 out.t252 0.00050016
R1672 out.n152 out.t20 0.00050016
R1673 out.n153 out.t46 0.00050016
R1674 out.n154 out.t1 0.00050016
R1675 out.n155 out.t95 0.00050016
R1676 out.n156 out.t60 0.00050016
R1677 out.n157 out.t33 0.00050016
R1678 out.n140 out.t229 0.00050016
R1679 out.n141 out.t201 0.00050016
R1680 out.n142 out.t243 0.00050016
R1681 out.n143 out.t9 0.00050016
R1682 out.n144 out.t32 0.00050016
R1683 out.n145 out.t154 0.00050016
R1684 out.n146 out.t76 0.00050016
R1685 out.n147 out.t114 0.00050016
R1686 out.n148 out.t47 0.00050016
R1687 out.n131 out.t15 0.00050016
R1688 out.n132 out.t41 0.00050016
R1689 out.n133 out.t28 0.00050016
R1690 out.n134 out.t69 0.00050016
R1691 out.n135 out.t87 0.00050016
R1692 out.n136 out.t51 0.00050016
R1693 out.n137 out.t326 0.00050016
R1694 out.n138 out.t329 0.00050016
R1695 out.n139 out.t62 0.00050016
R1696 out.n122 out.t242 0.00050016
R1697 out.n123 out.t231 0.00050016
R1698 out.n124 out.t218 0.00050016
R1699 out.n125 out.t78 0.00050016
R1700 out.n126 out.t45 0.00050016
R1701 out.n127 out.t61 0.00050016
R1702 out.n128 out.t30 0.00050016
R1703 out.n129 out.t18 0.00050016
R1704 out.n130 out.t10 0.00050016
R1705 out.n113 out.t169 0.00050016
R1706 out.n114 out.t202 0.00050016
R1707 out.n115 out.t131 0.00050016
R1708 out.n116 out.t115 0.00050016
R1709 out.n117 out.t135 0.00050016
R1710 out.n118 out.t44 0.00050016
R1711 out.n119 out.t335 0.00050016
R1712 out.n120 out.t7 0.00050016
R1713 out.n121 out.t137 0.00050016
R1714 out.n104 out.t90 0.00050016
R1715 out.n105 out.t71 0.00050016
R1716 out.n106 out.t55 0.00050016
R1717 out.n107 out.t26 0.00050016
R1718 out.n108 out.t14 0.00050016
R1719 out.n109 out.t37 0.00050016
R1720 out.n110 out.t333 0.00050016
R1721 out.n111 out.t336 0.00050016
R1722 out.n112 out.t156 0.00050016
R1723 out.n95 out.t186 0.00050016
R1724 out.n96 out.t150 0.00050016
R1725 out.n97 out.t111 0.00050016
R1726 out.n98 out.t96 0.00050016
R1727 out.n99 out.t77 0.00050016
R1728 out.n100 out.t59 0.00050016
R1729 out.n101 out.t134 0.00050016
R1730 out.n102 out.t0 0.00050016
R1731 out.n103 out.t2 0.00050016
R1732 out.n86 out.t36 0.00050016
R1733 out.n87 out.t50 0.00050016
R1734 out.n88 out.t208 0.00050016
R1735 out.n89 out.t21 0.00050016
R1736 out.n90 out.t11 0.00050016
R1737 out.n91 out.t177 0.00050016
R1738 out.n92 out.t120 0.00050016
R1739 out.n93 out.t82 0.00050016
R1740 out.n94 out.t97 0.00050016
R1741 vin.n0 vin 1.62229
R1742 vin.n5 vin.n4 1.13247
R1743 vin.n3 vin.n0 1.13247
R1744 vin.n1 vin 0.592032
R1745 vin.n7 vin.n6 0.399502
R1746 vin.n6 vin.n5 0.286623
R1747 vin.n2 vin.n1 0.271427
R1748 vin vin.n7 0.203188
R1749 vin.n5 vin.n3 0.016595
R1750 vin.n1 vin 0.0114968
R1751 vin.n6 vin 0.0114968
R1752 vin.n3 vin.n2 0.00879751
R1753 sample.n20 sample.t7 212.081
R1754 sample.n26 sample.t5 212.081
R1755 sample.n24 sample.t2 212.081
R1756 sample.n22 sample.t1 212.081
R1757 sample.n10 sample.t15 212.081
R1758 sample.n16 sample.t13 212.081
R1759 sample.n14 sample.t10 212.081
R1760 sample.n12 sample.t9 212.081
R1761 sample.n0 sample.t31 212.081
R1762 sample.n6 sample.t29 212.081
R1763 sample.n4 sample.t26 212.081
R1764 sample.n2 sample.t25 212.081
R1765 sample.n35 sample.t23 212.081
R1766 sample.n33 sample.t21 212.081
R1767 sample.n38 sample.t18 212.081
R1768 sample.n36 sample.t17 212.081
R1769 sample.n20 sample.t3 139.78
R1770 sample.n26 sample.t0 139.78
R1771 sample.n24 sample.t4 139.78
R1772 sample.n22 sample.t6 139.78
R1773 sample.n10 sample.t11 139.78
R1774 sample.n16 sample.t8 139.78
R1775 sample.n14 sample.t12 139.78
R1776 sample.n12 sample.t14 139.78
R1777 sample.n0 sample.t27 139.78
R1778 sample.n6 sample.t24 139.78
R1779 sample.n4 sample.t28 139.78
R1780 sample.n2 sample.t30 139.78
R1781 sample.n35 sample.t19 139.78
R1782 sample.n33 sample.t16 139.78
R1783 sample.n38 sample.t20 139.78
R1784 sample.n36 sample.t22 139.78
R1785 sample.n23 sample.n21 97.5045
R1786 sample.n13 sample.n11 97.5045
R1787 sample.n3 sample.n1 97.5045
R1788 sample.n40 sample.n37 97.5045
R1789 sample.n28 sample.n27 76.0005
R1790 sample.n25 sample.n21 76.0005
R1791 sample.n18 sample.n17 76.0005
R1792 sample.n15 sample.n11 76.0005
R1793 sample.n8 sample.n7 76.0005
R1794 sample.n5 sample.n1 76.0005
R1795 sample.n40 sample.n39 76.0005
R1796 sample.n29 sample.n20 44.4802
R1797 sample.n19 sample.n10 44.4802
R1798 sample.n9 sample.n0 44.4802
R1799 sample.n42 sample.n35 44.4802
R1800 sample.n30 sample 33.6245
R1801 sample.n23 sample.n22 30.6732
R1802 sample.n24 sample.n23 30.6732
R1803 sample.n25 sample.n24 30.6732
R1804 sample.n26 sample.n25 30.6732
R1805 sample.n27 sample.n26 30.6732
R1806 sample.n27 sample.n20 30.6732
R1807 sample.n13 sample.n12 30.6732
R1808 sample.n14 sample.n13 30.6732
R1809 sample.n15 sample.n14 30.6732
R1810 sample.n16 sample.n15 30.6732
R1811 sample.n17 sample.n16 30.6732
R1812 sample.n17 sample.n10 30.6732
R1813 sample.n3 sample.n2 30.6732
R1814 sample.n4 sample.n3 30.6732
R1815 sample.n5 sample.n4 30.6732
R1816 sample.n6 sample.n5 30.6732
R1817 sample.n7 sample.n6 30.6732
R1818 sample.n7 sample.n0 30.6732
R1819 sample.n37 sample.n36 30.6732
R1820 sample.n39 sample.n38 30.6732
R1821 sample.n34 sample.n33 30.6732
R1822 sample.n35 sample.n34 30.6732
R1823 sample.n29 sample.n28 23.9042
R1824 sample.n19 sample.n18 23.9042
R1825 sample.n9 sample.n8 23.9042
R1826 sample.n42 sample.n41 23.9042
R1827 sample.n28 sample.n21 21.5045
R1828 sample.n18 sample.n11 21.5045
R1829 sample.n8 sample.n1 21.5045
R1830 sample.n41 sample.n40 21.5045
R1831 sample sample.n29 5.38578
R1832 sample sample.n19 5.38578
R1833 sample sample.n9 5.38578
R1834 sample sample.n42 5.38445
R1835 sample sample.n32 3.3673
R1836 sample.n32 sample.n31 3.30675
R1837 sample.n31 sample.n30 3.30675
R1838 sample.n30 sample 0.0610469
R1839 sample.n31 sample 0.0610469
R1840 sample.n32 sample 0.0610469
R1841 enb.n17 enb.t17 212.081
R1842 enb.n15 enb.t15 212.081
R1843 enb.n11 enb.t12 212.081
R1844 enb.n9 enb.t11 212.081
R1845 enb.n0 enb.t7 143.071
R1846 enb.n8 enb.t3 142.75
R1847 enb.n0 enb.t0 142.75
R1848 enb.n1 enb.t4 142.75
R1849 enb.n2 enb.t8 142.75
R1850 enb.n3 enb.t1 142.75
R1851 enb.n4 enb.t5 142.75
R1852 enb.n5 enb.t6 142.75
R1853 enb.n6 enb.t2 142.75
R1854 enb.n7 enb.t9 142.75
R1855 enb.n17 enb.t13 139.78
R1856 enb.n15 enb.t10 139.78
R1857 enb.n11 enb.t14 139.78
R1858 enb.n9 enb.t16 139.78
R1859 enb.n13 enb.n10 97.5045
R1860 enb.n13 enb.n12 76.0005
R1861 enb.n18 enb.n17 39.8685
R1862 enb.n10 enb.n9 30.6732
R1863 enb.n12 enb.n11 30.6732
R1864 enb.n16 enb.n15 30.6732
R1865 enb.n17 enb.n16 30.6732
R1866 enb.n14 enb.n13 21.5045
R1867 enb.n18 enb.n14 19.201
R1868 enb.n19 enb.n8 6.80862
R1869 enb.n19 enb.n18 4.11918
R1870 enb.n8 enb.n7 0.321152
R1871 enb.n7 enb.n6 0.321152
R1872 enb.n6 enb.n5 0.321152
R1873 enb.n5 enb.n4 0.321152
R1874 enb.n4 enb.n3 0.321152
R1875 enb.n3 enb.n2 0.321152
R1876 enb.n2 enb.n1 0.321152
R1877 enb.n1 enb.n0 0.321152
R1878 enb enb.n19 0.063
R1879 en_buf.n0 en_buf.t8 135.841
R1880 en_buf.n4 en_buf.t3 135.841
R1881 en_buf.n2 en_buf.t1 135.52
R1882 en_buf.n1 en_buf.t7 135.52
R1883 en_buf.n0 en_buf.t4 135.52
R1884 en_buf.n4 en_buf.t5 135.52
R1885 en_buf.n5 en_buf.t9 135.52
R1886 en_buf.n6 en_buf.t2 135.52
R1887 en_buf.n7 en_buf.t6 134.576
R1888 en_buf.n3 en_buf.t0 134.576
R1889 en_buf en_buf.n8 1.05289
R1890 en_buf.n1 en_buf.n0 0.321152
R1891 en_buf.n2 en_buf.n1 0.321152
R1892 en_buf.n6 en_buf.n5 0.321152
R1893 en_buf.n5 en_buf.n4 0.321152
R1894 en_buf.n3 en_buf.n2 0.315896
R1895 en_buf.n7 en_buf.n6 0.315896
R1896 en_buf.n8 en_buf.n3 0.121984
R1897 en_buf.n8 en_buf.n7 0.121984
C0 vin sw_top_3/m2_990_200# 0.0472f
C1 carray_0/n4 ctl7 1.72e-20
C2 ctl5 ctl4 0.193f
C3 vdd carray_0/via23_4_429/m2_1_40# 0.0108f
C4 carray_0/m2_24600_1156# sample 6.55e-20
C5 carray_0/m2_40200_1156# sample 6.55e-20
C6 ctl7 vdd 0.021f
C7 carray_0/m2_29800_1156# sample 6.55e-20
C8 carray_0/n4 sample 5.55e-19
C9 vin carray_0/via23_4_635/m2_1_40# 0.0175f
C10 ctl2 vdd 0.025f
C11 sw_top_0/m2_1158_361# en_buf 0.00725f
C12 carray_0/m2_42800_1156# carray_0/via23_4_641/m2_1_40# 2.84e-32
C13 vdd sample 0.303f
C14 sample carray_0/via23_4_369/m2_1_40# 9.23e-21
C15 vdd enb 0.0379f
C16 carray_0/n5 ctl7 3.35e-20
C17 ctl7 carray_0/n6 0.0169f
C18 en_buf out 0.0185f
C19 carray_0/n1 ctl1 0.0173f
C20 sample sw_top_3/m2_1158_361# 0.0218f
C21 enb sw_top_3/m2_1158_361# 0.0127f
C22 carray_0/m2_31100_1156# sample 6.55e-20
C23 en_buf sw_top_0/m2_990_200# 0.00185f
C24 vdd dum 0.0273f
C25 ctl2 ctl3 0.193f
C26 carray_0/m3_42700_1156# vdd 0.00943f
C27 carray_0/n4 carray_0/n2 4.38e-20
C28 sample carray_0/m2_41500_1156# 6.55e-20
C29 carray_0/n5 sample 0.0017f
C30 carray_0/n4 carray_0/via23_4_96/m2_1_40# 5.45e-19
C31 carray_0/via23_4_702/m2_1_40# enb 0.0244f
C32 sample carray_0/n6 0.0059f
C33 vdd carray_0/n0 0.0911f
C34 vdd carray_0/n2 0.0953f
C35 carray_0/m3_42700_1156# sw_top_3/m2_1158_361# 0.00278f
C36 sw_top_0/m2_1158_361# out 0.071f
C37 carray_0/n1 carray_0/n3 8.82e-20
C38 dum carray_0/n6 6.25e-20
C39 vdd sw_top_3/m2_990_200# 0.00684f
C40 out carray_0/via23_4_419/m2_1_40# 0.0569f
C41 carray_0/n4 carray_0/n7 3.37e-19
C42 sample carray_0/m2_42800_1156# 3.33e-19
C43 sw_top_0/m2_1158_361# sw_top_0/m2_990_200# -1.14e-31
C44 enb carray_0/m2_42800_1156# 0.00743f
C45 ctl3 carray_0/n2 0.0164f
C46 carray_0/n5 carray_0/n0 3.34e-19
C47 sw_top_0/m2_990_200# out 0.00532f
C48 vdd vin 0.572f
C49 sw_top_3/m2_1158_361# sw_top_3/m2_990_200# -1.14e-31
C50 carray_0/n6 carray_0/n0 1.07e-19
C51 carray_0/n5 carray_0/n2 4.38e-20
C52 carray_0/n6 carray_0/n2 4.38e-20
C53 carray_0/n3 out 0.00516f
C54 sw_top_0/m2_1158_361# carray_0/via23_4_367/m2_1_40# 0.00501f
C55 ctl0 sample 0.00375f
C56 carray_0/n5 carray_0/via23_4_96/m2_1_40# 0.00116f
C57 vdd carray_0/n7 0.0901f
C58 sample carray_0/via23_4_448/m2_1_40# 9.23e-21
C59 carray_0/m2_800_1156# carray_0/n2 0.00165f
C60 carray_0/via23_4_367/m2_1_40# out 8.98e-19
C61 carray_0/m3_42500_1156# sample 0.0051f
C62 out carray_0/via23_4_704/m2_1_40# 0.0569f
C63 sample carray_0/via23_4_439/m2_1_40# 9.23e-21
C64 vin sw_top_3/m2_1158_361# 0.141f
C65 ctl6 ctl7 0.193f
C66 carray_0/m3_42700_1156# carray_0/m2_42800_1156# 5.68e-32
C67 vdd carray_0/via23_4_635/m2_1_40# 0.0106f
C68 ctl0 dum 0.193f
C69 carray_0/via23_4_702/m2_1_40# vin 0.0292f
C70 sample carray_0/ndum 11.1f
C71 out carray_0/via23_4_642/m2_1_40# 0.045f
C72 carray_0/n3 ctl4 0.0164f
C73 carray_0/n5 carray_0/n7 3.54e-19
C74 sw_top_3/m2_1158_361# carray_0/via23_4_635/m2_1_40# 0.0215f
C75 carray_0/via23_4_446/m2_1_40# sample 9.23e-21
C76 carray_0/n6 carray_0/n7 1.2f
C77 vin carray_0/via23_4_705/m2_1_40# 0.0358f
C78 ctl0 carray_0/n0 0.0173f
C79 dum carray_0/ndum 0.0173f
C80 out carray_0/via23_4_641/m2_1_40# 0.0791f
C81 carray_0/m2_42800_1156# vin 0.00125f
C82 carray_0/n1 ctl7 0.00139f
C83 en_buf sample 0.124f
C84 ctl7 ctl1 0.193f
C85 sw_top_0/m2_1158_361# carray_0/via23_4_429/m2_1_40# 0.0214f
C86 carray_0/n0 carray_0/ndum 1.1f
C87 carray_0/via23_4_414/m2_1_40# vin 0.0351f
C88 out carray_0/via23_4_429/m2_1_40# 0.138f
C89 carray_0/via23_4_128/m2_1_40# carray_0/n2 0.0993f
C90 ctl0 carray_0/n7 1.64e-19
C91 carray_0/m2_42800_1156# carray_0/via23_4_635/m2_1_40# 2.84e-32
C92 carray_0/n4 vdd 0.0879f
C93 carray_0/via23_4_449/m2_1_40# sample 9.23e-21
C94 carray_0/n1 sample 0.00244f
C95 sample ctl1 0.00255f
C96 carray_0/m2_27200_1156# sample 6.55e-20
C97 carray_0/n7 carray_0/ndum 3.26e-19
C98 sw_top_0/m2_1158_361# sample 0.0218f
C99 sample carray_0/via23_4_455/m2_1_40# 4.62e-21
C100 sw_top_0/m2_1158_361# enb 0.00635f
C101 carray_0/n4 ctl3 0.00139f
C102 carray_0/n1 dum 1.97e-19
C103 sample out 0.00645f
C104 vdd sw_top_3/m2_1158_361# 0.0369f
C105 enb out 0.133f
C106 carray_0/n4 carray_0/n5 1.27f
C107 enb carray_0/via23_4_419/m2_1_40# 0.0258f
C108 carray_0/n4 carray_0/n6 6.52e-20
C109 ctl6 carray_0/n7 0.00139f
C110 en_buf sw_top_3/m2_990_200# 0.00369f
C111 carray_0/n4 carray_0/m2_800_1156# 5.11e-19
C112 vdd ctl3 0.021f
C113 sample carray_0/via23_4_447/m2_1_40# 9.23e-21
C114 carray_0/n3 ctl2 0.00139f
C115 sw_top_0/m2_990_200# sample 0.121f
C116 sw_top_0/m2_990_200# enb 1e-20
C117 carray_0/n5 vdd 0.0888f
C118 carray_0/n1 carray_0/n0 1.14f
C119 carray_0/via23_4_702/m2_1_40# vdd 0.0203f
C120 vdd carray_0/n6 0.0895f
C121 carray_0/n3 sample 3.92e-19
C122 ctl1 carray_0/n0 0.00139f
C123 sw_top_0/m2_1158_361# carray_0/m3_42700_1156# 0.00277f
C124 carray_0/via23_4_460/m2_1_40# sample 9.23e-21
C125 en_buf vin 0.0668f
C126 carray_0/m3_42700_1156# out 0.0285f
C127 carray_0/via23_4_367/m2_1_40# sample 0.0408f
C128 vdd carray_0/via23_4_705/m2_1_40# 0.00874f
C129 enb carray_0/via23_4_704/m2_1_40# 0.0236f
C130 carray_0/n4 ctl5 0.0164f
C131 carray_0/m2_25900_1156# sample 6.55e-20
C132 out carray_0/n2 0.0119f
C133 vdd ctl5 0.021f
C134 carray_0/via23_4_705/m2_1_40# sw_top_3/m2_1158_361# 0.0136f
C135 sample carray_0/via23_4_366/m2_1_40# 9.23e-21
C136 carray_0/m2_32400_1156# sample 6.55e-20
C137 vdd carray_0/m2_42800_1156# 0.0238f
C138 carray_0/n5 carray_0/n6 1.24f
C139 carray_0/n5 carray_0/m2_800_1156# 1.36e-19
C140 carray_0/n1 carray_0/n7 1.17f
C141 out sw_top_3/m2_990_200# 0.00924f
C142 carray_0/n6 carray_0/m2_800_1156# 2.66e-20
C143 vdd carray_0/via23_4_414/m2_1_40# 0.00801f
C144 ctl1 carray_0/n7 0.0172f
C145 carray_0/n3 carray_0/n2 1.34f
C146 ctl0 vdd 0.021f
C147 sample carray_0/via23_4_368/m2_1_40# 9.23e-21
C148 carray_0/m2_42800_1156# sw_top_3/m2_1158_361# 0.0031f
C149 carray_0/n3 carray_0/via23_4_96/m2_1_40# 8.98e-19
C150 sw_top_0/m2_1158_361# vin 0.116f
C151 enb carray_0/via23_4_641/m2_1_40# 0.0247f
C152 out vin 0.25f
C153 vin carray_0/via23_4_419/m2_1_40# 0.0402f
C154 carray_0/n5 ctl5 0.017f
C155 carray_0/n6 ctl5 0.00139f
C156 carray_0/m2_33700_1156# sample 6.55e-20
C157 sw_top_0/m2_990_200# vin 1.53e-20
C158 carray_0/n4 ctl6 1.72e-20
C159 vdd carray_0/ndum 0.124f
C160 sample carray_0/via23_4_378/m2_1_40# 9.23e-21
C161 sample carray_0/via23_4_458/m2_1_40# 9.23e-21
C162 carray_0/n5 ctl0 4.89e-20
C163 out carray_0/via23_4_635/m2_1_40# 0.152f
C164 ctl0 carray_0/n6 1.31e-19
C165 carray_0/n3 carray_0/n7 5.65e-19
C166 carray_0/via23_4_367/m2_1_40# vin 0.017f
C167 sample carray_0/via23_4_379/m2_1_40# 9.23e-21
C168 carray_0/via23_4_704/m2_1_40# vin 0.04f
C169 ctl6 vdd 0.021f
C170 ctl7 sample 0.00169f
C171 carray_0/m2_35000_1156# sample 6.55e-20
C172 vin carray_0/via23_4_642/m2_1_40# 0.0375f
C173 en_buf vdd 0.00684f
C174 carray_0/n5 ctl6 0.0166f
C175 enb sample 0.0218f
C176 ctl6 carray_0/n6 0.0171f
C177 carray_0/n4 carray_0/n1 6.52e-20
C178 en_buf sw_top_3/m2_1158_361# 0.00726f
C179 vin carray_0/via23_4_641/m2_1_40# 0.0325f
C180 carray_0/n4 ctl1 1.72e-20
C181 carray_0/n1 vdd 0.0908f
C182 carray_0/m2_36300_1156# sample 6.55e-20
C183 dum sample 0.00816f
C184 vdd ctl1 0.021f
C185 carray_0/m3_42700_1156# sample 0.0051f
C186 carray_0/n4 out 0.00281f
C187 carray_0/m3_42700_1156# enb 0.00364f
C188 ctl6 ctl5 0.193f
C189 carray_0/via23_4_429/m2_1_40# vin 0.0183f
C190 ctl0 carray_0/ndum 0.00139f
C191 ctl2 carray_0/n2 0.0168f
C192 sw_top_0/m2_1158_361# vdd 0.036f
C193 sample carray_0/n0 0.00854f
C194 vdd out 0.213f
C195 vdd carray_0/via23_4_419/m2_1_40# 0.0212f
C196 carray_0/n4 carray_0/n3 1.31f
C197 ctl7 carray_0/n7 0.0173f
C198 carray_0/m3_900_1156# carray_0/n2 0.0151f
C199 carray_0/n5 carray_0/n1 8.23e-20
C200 carray_0/n5 ctl1 3.35e-20
C201 carray_0/n1 carray_0/n6 1.07e-19
C202 ctl1 carray_0/n6 1.31e-19
C203 vdd sw_top_0/m2_990_200# 0.00684f
C204 sample sw_top_3/m2_990_200# 0.121f
C205 out sw_top_3/m2_1158_361# 0.0778f
C206 enb sw_top_3/m2_990_200# 0.00726f
C207 carray_0/n4 ctl4 0.0169f
C208 dum carray_0/n0 0.0178f
C209 carray_0/n3 vdd 0.086f
C210 sample carray_0/via23_4_381/m2_1_40# 9.23e-21
C211 vdd carray_0/via23_4_367/m2_1_40# 0.0196f
C212 vdd carray_0/via23_4_704/m2_1_40# 0.0226f
C213 sample vin 0.302f
C214 carray_0/m2_37600_1156# sample 6.55e-20
C215 carray_0/n5 out 0.00162f
C216 carray_0/via23_4_702/m2_1_40# out 0.0879f
C217 enb vin 0.172f
C218 vdd ctl4 0.021f
C219 sample carray_0/n7 4.96f
C220 sample carray_0/via23_4_459/m2_1_40# 9.23e-21
C221 out carray_0/via23_4_705/m2_1_40# 0.0454f
C222 carray_0/n3 ctl3 0.0168f
C223 carray_0/via23_4_96/m2_1_40# carray_0/n2 0.163f
C224 vdd carray_0/via23_4_642/m2_1_40# 0.0178f
C225 carray_0/n5 carray_0/n3 5.3e-20
C226 carray_0/via23_4_380/m2_1_40# sample 9.23e-21
C227 carray_0/n3 carray_0/n6 5.3e-20
C228 carray_0/n1 ctl0 0.0175f
C229 carray_0/m3_42700_1156# vin 9.27e-20
C230 carray_0/n3 carray_0/m2_800_1156# 9.73e-19
C231 dum carray_0/n7 2.59e-19
C232 ctl0 ctl1 0.193f
C233 sw_top_0/m2_1158_361# carray_0/m2_42800_1156# 0.00392f
C234 ctl3 ctl4 0.193f
C235 carray_0/m2_23300_1156# sample 6.55e-20
C236 carray_0/n5 ctl4 0.00139f
C237 out carray_0/m2_42800_1156# 0.0555f
C238 sw_top_3/m2_1158_361# carray_0/via23_4_642/m2_1_40# 0.00397f
C239 sw_top_0/m2_1158_361# carray_0/via23_4_414/m2_1_40# 0.0116f
C240 carray_0/m2_38900_1156# sample 6.55e-20
C241 vdd carray_0/via23_4_641/m2_1_40# 0.0208f
C242 out carray_0/via23_4_414/m2_1_40# 0.0451f
C243 carray_0/n7 carray_0/n0 1.45e-19
C244 carray_0/n7 carray_0/n2 7.53e-19
C245 carray_0/n1 carray_0/ndum 2.07e-19
C246 carray_0/m2_28500_1156# sample 6.55e-20
C247 enb.t3 vss 0.0729f
C248 enb.t9 vss 0.0729f
C249 enb.t2 vss 0.0729f
C250 enb.t6 vss 0.0729f
C251 enb.t5 vss 0.0729f
C252 enb.t1 vss 0.0729f
C253 enb.t8 vss 0.0729f
C254 enb.t4 vss 0.0729f
C255 enb.t0 vss 0.0729f
C256 enb.t7 vss 0.0731f
C257 enb.n0 vss 0.196f
C258 enb.n1 vss 0.103f
C259 enb.n2 vss 0.103f
C260 enb.n3 vss 0.103f
C261 enb.n4 vss 0.103f
C262 enb.n5 vss 0.103f
C263 enb.n6 vss 0.103f
C264 enb.n7 vss 0.103f
C265 enb.n8 vss 0.471f
C266 enb.t11 vss 0.0304f
C267 enb.t16 vss 0.0179f
C268 enb.n9 vss 0.041f
C269 enb.n10 vss 0.026f
C270 enb.t12 vss 0.0304f
C271 enb.t14 vss 0.0179f
C272 enb.n11 vss 0.0438f
C273 enb.n12 vss 0.0201f
C274 enb.n13 vss 0.0516f
C275 enb.n14 vss 0.0289f
C276 enb.t17 vss 0.0304f
C277 enb.t13 vss 0.0179f
C278 enb.t15 vss 0.0304f
C279 enb.t10 vss 0.0179f
C280 enb.n15 vss 0.0438f
C281 enb.n16 vss 0.0201f
C282 enb.n17 vss 0.051f
C283 enb.n18 vss 0.512f
C284 enb.n19 vss 1.14f
C285 sample.t31 vss 0.0132f
C286 sample.t27 vss 0.00777f
C287 sample.n0 vss 0.0219f
C288 sample.n1 vss 0.0224f
C289 sample.t29 vss 0.0132f
C290 sample.t24 vss 0.00777f
C291 sample.t26 vss 0.0132f
C292 sample.t28 vss 0.00777f
C293 sample.t25 vss 0.0132f
C294 sample.t30 vss 0.00777f
C295 sample.n2 vss 0.0178f
C296 sample.n3 vss 0.0113f
C297 sample.n4 vss 0.019f
C298 sample.n5 vss 0.0087f
C299 sample.n6 vss 0.019f
C300 sample.n7 vss 0.0087f
C301 sample.n8 vss 0.0139f
C302 sample.n9 vss 0.0295f
C303 sample.t15 vss 0.0132f
C304 sample.t11 vss 0.00777f
C305 sample.n10 vss 0.0219f
C306 sample.n11 vss 0.0224f
C307 sample.t13 vss 0.0132f
C308 sample.t8 vss 0.00777f
C309 sample.t10 vss 0.0132f
C310 sample.t12 vss 0.00777f
C311 sample.t9 vss 0.0132f
C312 sample.t14 vss 0.00777f
C313 sample.n12 vss 0.0178f
C314 sample.n13 vss 0.0113f
C315 sample.n14 vss 0.019f
C316 sample.n15 vss 0.0087f
C317 sample.n16 vss 0.019f
C318 sample.n17 vss 0.0087f
C319 sample.n18 vss 0.0139f
C320 sample.n19 vss 0.0295f
C321 sample.t7 vss 0.0132f
C322 sample.t3 vss 0.00777f
C323 sample.n20 vss 0.0219f
C324 sample.n21 vss 0.0224f
C325 sample.t5 vss 0.0132f
C326 sample.t0 vss 0.00777f
C327 sample.t2 vss 0.0132f
C328 sample.t4 vss 0.00777f
C329 sample.t1 vss 0.0132f
C330 sample.t6 vss 0.00777f
C331 sample.n22 vss 0.0178f
C332 sample.n23 vss 0.0113f
C333 sample.n24 vss 0.019f
C334 sample.n25 vss 0.0087f
C335 sample.n26 vss 0.019f
C336 sample.n27 vss 0.0087f
C337 sample.n28 vss 0.0139f
C338 sample.n29 vss 0.0295f
C339 sample.n30 vss 6.3f
C340 sample.n31 vss 0.534f
C341 sample.n32 vss 0.539f
C342 sample.t23 vss 0.0132f
C343 sample.t19 vss 0.00777f
C344 sample.t21 vss 0.0132f
C345 sample.t16 vss 0.00777f
C346 sample.n33 vss 0.019f
C347 sample.n34 vss 0.0087f
C348 sample.n35 vss 0.0219f
C349 sample.t17 vss 0.0132f
C350 sample.t22 vss 0.00777f
C351 sample.n36 vss 0.0178f
C352 sample.n37 vss 0.0113f
C353 sample.t18 vss 0.0132f
C354 sample.t20 vss 0.00777f
C355 sample.n38 vss 0.019f
C356 sample.n39 vss 0.0087f
C357 sample.n40 vss 0.0224f
C358 sample.n41 vss 0.0139f
C359 sample.n42 vss 0.0295f
C360 vin.n0 vss 2.41f
C361 vin.n1 vss 3.1f
C362 vin.n2 vss 1.5f
C363 vin.n4 vss 0.067f
C364 vin.n5 vss 1.53f
C365 vin.n6 vss 2.07f
C366 vin.n7 vss 3.38f
C367 out.n0 vss 0.0234f
C368 out.n1 vss 0.00829f
C369 out.n2 vss 0.00378f
C370 out.n3 vss 0.00378f
C371 out.n4 vss 0.0128f
C372 out.n5 vss 0.00756f
C373 out.n6 vss 0.00454f
C374 out.n7 vss 0.00378f
C375 out.n8 vss 0.00378f
C376 out.n9 vss 0.00454f
C377 out.n10 vss 0.00378f
C378 out.n11 vss 0.00378f
C379 out.n12 vss 0.00912f
C380 out.n13 vss 0.013f
C381 out.n14 vss 0.00912f
C382 out.n15 vss 0.00378f
C383 out.n16 vss 0.00378f
C384 out.n17 vss 0.0234f
C385 out.n18 vss 0.00454f
C386 out.n19 vss 0.00378f
C387 out.n20 vss 0.00378f
C388 out.n21 vss 0.00756f
C389 out.n22 vss 0.00789f
C390 out.n23 vss 0.0144f
C391 out.n24 vss 0.0222f
C392 out.n25 vss 0.00378f
C393 out.n26 vss 0.00454f
C394 out.n27 vss 0.00378f
C395 out.n28 vss 0.00462f
C396 out.n29 vss 0.143f
C397 out.n30 vss 0.143f
C398 out.n31 vss 0.00462f
C399 out.n32 vss 0.00378f
C400 out.n33 vss 0.00454f
C401 out.n34 vss 0.00378f
C402 out.n35 vss 0.00378f
C403 out.n36 vss 0.00454f
C404 out.n37 vss 0.00378f
C405 out.n38 vss 0.00462f
C406 out.n39 vss 0.0128f
C407 out.n40 vss 0.00756f
C408 out.n41 vss 0.00829f
C409 out.n42 vss 0.00378f
C410 out.n43 vss 0.00378f
C411 out.n44 vss 0.00454f
C412 out.n45 vss 0.00378f
C413 out.n46 vss 0.00378f
C414 out.n47 vss 0.0234f
C415 out.n48 vss 0.00454f
C416 out.n49 vss 0.00378f
C417 out.n50 vss 0.00378f
C418 out.n51 vss 0.00912f
C419 out.n52 vss 0.143f
C420 out.n53 vss 0.143f
C421 out.n54 vss 0.00462f
C422 out.n55 vss 0.00378f
C423 out.n56 vss 0.00454f
C424 out.n57 vss 0.00378f
C425 out.n58 vss 0.00378f
C426 out.n59 vss 0.00454f
C427 out.n60 vss 0.00378f
C428 out.n61 vss 0.00462f
C429 out.n62 vss 0.0128f
C430 out.n63 vss 0.00756f
C431 out.n64 vss 0.00829f
C432 out.n65 vss 0.00378f
C433 out.n66 vss 0.00378f
C434 out.n67 vss 0.00454f
C435 out.n68 vss 0.00378f
C436 out.n69 vss 0.00378f
C437 out.n70 vss 0.0234f
C438 out.n71 vss 0.00454f
C439 out.n72 vss 0.00378f
C440 out.n73 vss 0.00378f
C441 out.n74 vss 0.00912f
C442 out.n75 vss 0.144f
C443 out.n76 vss 0.143f
C444 out.n77 vss 0.00476f
C445 out.n78 vss 0.00378f
C446 out.n79 vss 0.00454f
C447 out.n80 vss 0.00378f
C448 out.n81 vss 0.00378f
C449 out.n82 vss 0.00454f
C450 out.n83 vss 0.00378f
C451 out.n84 vss 0.00462f
C452 out.n85 vss 0.0714f
C453 out.t97 vss 0.302f
C454 out.t82 vss 0.302f
C455 out.t120 vss 0.302f
C456 out.t177 vss 0.302f
C457 out.t11 vss 0.302f
C458 out.t21 vss 0.302f
C459 out.t208 vss 0.302f
C460 out.t50 vss 0.302f
C461 out.t36 vss 0.302f
C462 out.t101 vss 0.538f
C463 out.n86 vss 0.29f
C464 out.n87 vss 0.29f
C465 out.n88 vss 0.29f
C466 out.n89 vss 0.29f
C467 out.n90 vss 0.29f
C468 out.n91 vss 0.29f
C469 out.n92 vss 0.29f
C470 out.n93 vss 0.29f
C471 out.n94 vss 0.253f
C472 out.t2 vss 0.302f
C473 out.t0 vss 0.302f
C474 out.t134 vss 0.302f
C475 out.t59 vss 0.302f
C476 out.t77 vss 0.302f
C477 out.t96 vss 0.302f
C478 out.t111 vss 0.302f
C479 out.t150 vss 0.302f
C480 out.t186 vss 0.302f
C481 out.t83 vss 0.538f
C482 out.n95 vss 0.29f
C483 out.n96 vss 0.29f
C484 out.n97 vss 0.29f
C485 out.n98 vss 0.29f
C486 out.n99 vss 0.29f
C487 out.n100 vss 0.29f
C488 out.n101 vss 0.29f
C489 out.n102 vss 0.29f
C490 out.n103 vss 0.253f
C491 out.t156 vss 0.302f
C492 out.t336 vss 0.302f
C493 out.t333 vss 0.302f
C494 out.t37 vss 0.302f
C495 out.t14 vss 0.302f
C496 out.t26 vss 0.302f
C497 out.t55 vss 0.302f
C498 out.t71 vss 0.302f
C499 out.t90 vss 0.302f
C500 out.t141 vss 0.538f
C501 out.n104 vss 0.29f
C502 out.n105 vss 0.29f
C503 out.n106 vss 0.29f
C504 out.n107 vss 0.29f
C505 out.n108 vss 0.29f
C506 out.n109 vss 0.29f
C507 out.n110 vss 0.29f
C508 out.n111 vss 0.29f
C509 out.n112 vss 0.253f
C510 out.t137 vss 0.302f
C511 out.t7 vss 0.302f
C512 out.t335 vss 0.302f
C513 out.t44 vss 0.302f
C514 out.t135 vss 0.302f
C515 out.t115 vss 0.302f
C516 out.t131 vss 0.302f
C517 out.t202 vss 0.302f
C518 out.t169 vss 0.302f
C519 out.t121 vss 0.538f
C520 out.n113 vss 0.29f
C521 out.n114 vss 0.29f
C522 out.n115 vss 0.29f
C523 out.n116 vss 0.29f
C524 out.n117 vss 0.29f
C525 out.n118 vss 0.29f
C526 out.n119 vss 0.29f
C527 out.n120 vss 0.29f
C528 out.n121 vss 0.253f
C529 out.t10 vss 0.302f
C530 out.t18 vss 0.302f
C531 out.t30 vss 0.302f
C532 out.t61 vss 0.302f
C533 out.t45 vss 0.302f
C534 out.t78 vss 0.302f
C535 out.t218 vss 0.302f
C536 out.t231 vss 0.302f
C537 out.t242 vss 0.302f
C538 out.t65 vss 0.538f
C539 out.n122 vss 0.29f
C540 out.n123 vss 0.29f
C541 out.n124 vss 0.29f
C542 out.n125 vss 0.29f
C543 out.n126 vss 0.29f
C544 out.n127 vss 0.29f
C545 out.n128 vss 0.29f
C546 out.n129 vss 0.29f
C547 out.n130 vss 0.253f
C548 out.t62 vss 0.302f
C549 out.t329 vss 0.302f
C550 out.t326 vss 0.302f
C551 out.t51 vss 0.302f
C552 out.t87 vss 0.302f
C553 out.t69 vss 0.302f
C554 out.t28 vss 0.302f
C555 out.t41 vss 0.302f
C556 out.t15 vss 0.302f
C557 out.t191 vss 0.538f
C558 out.n131 vss 0.29f
C559 out.n132 vss 0.29f
C560 out.n133 vss 0.29f
C561 out.n134 vss 0.29f
C562 out.n135 vss 0.29f
C563 out.n136 vss 0.29f
C564 out.n137 vss 0.29f
C565 out.n138 vss 0.29f
C566 out.n139 vss 0.253f
C567 out.t47 vss 0.302f
C568 out.t114 vss 0.302f
C569 out.t76 vss 0.302f
C570 out.t154 vss 0.302f
C571 out.t32 vss 0.302f
C572 out.t9 vss 0.302f
C573 out.t243 vss 0.302f
C574 out.t201 vss 0.302f
C575 out.t229 vss 0.302f
C576 out.t178 vss 0.538f
C577 out.n140 vss 0.29f
C578 out.n141 vss 0.29f
C579 out.n142 vss 0.29f
C580 out.n143 vss 0.29f
C581 out.n144 vss 0.29f
C582 out.n145 vss 0.29f
C583 out.n146 vss 0.29f
C584 out.n147 vss 0.29f
C585 out.n148 vss 0.253f
C586 out.t33 vss 0.302f
C587 out.t60 vss 0.302f
C588 out.t95 vss 0.302f
C589 out.t1 vss 0.302f
C590 out.t46 vss 0.302f
C591 out.t20 vss 0.302f
C592 out.t252 vss 0.302f
C593 out.t259 vss 0.302f
C594 out.t215 vss 0.302f
C595 out.t160 vss 0.538f
C596 out.n149 vss 0.29f
C597 out.n150 vss 0.29f
C598 out.n151 vss 0.29f
C599 out.n152 vss 0.29f
C600 out.n153 vss 0.29f
C601 out.n154 vss 0.29f
C602 out.n155 vss 0.29f
C603 out.n156 vss 0.29f
C604 out.n157 vss 0.253f
C605 out.t34 vss 0.302f
C606 out.t283 vss 0.302f
C607 out.t286 vss 0.302f
C608 out.t307 vss 0.302f
C609 out.t312 vss 0.302f
C610 out.t324 vss 0.302f
C611 out.t317 vss 0.302f
C612 out.t321 vss 0.302f
C613 out.t327 vss 0.302f
C614 out.t22 vss 0.538f
C615 out.n158 vss 0.29f
C616 out.n159 vss 0.29f
C617 out.n160 vss 0.29f
C618 out.n161 vss 0.29f
C619 out.n162 vss 0.29f
C620 out.n163 vss 0.29f
C621 out.n164 vss 0.29f
C622 out.n165 vss 0.29f
C623 out.n166 vss 0.253f
C624 out.t117 vss 0.302f
C625 out.t337 vss 0.302f
C626 out.t4 vss 0.302f
C627 out.t24 vss 0.302f
C628 out.t53 vss 0.302f
C629 out.t39 vss 0.302f
C630 out.t339 vss 0.302f
C631 out.t16 vss 0.302f
C632 out.t6 vss 0.302f
C633 out.t102 vss 0.538f
C634 out.n167 vss 0.29f
C635 out.n168 vss 0.29f
C636 out.n169 vss 0.29f
C637 out.n170 vss 0.29f
C638 out.n171 vss 0.29f
C639 out.n172 vss 0.29f
C640 out.n173 vss 0.29f
C641 out.n174 vss 0.29f
C642 out.n175 vss 0.253f
C643 out.t98 vss 0.302f
C644 out.t224 vss 0.302f
C645 out.t19 vss 0.302f
C646 out.t73 vss 0.302f
C647 out.t226 vss 0.302f
C648 out.t109 vss 0.302f
C649 out.t151 vss 0.302f
C650 out.t187 vss 0.302f
C651 out.t199 vss 0.302f
C652 out.t122 vss 0.538f
C653 out.n176 vss 0.29f
C654 out.n177 vss 0.29f
C655 out.n178 vss 0.29f
C656 out.n179 vss 0.29f
C657 out.n180 vss 0.29f
C658 out.n181 vss 0.29f
C659 out.n182 vss 0.29f
C660 out.n183 vss 0.29f
C661 out.n184 vss 0.253f
C662 out.t138 vss 0.302f
C663 out.t8 vss 0.302f
C664 out.t31 vss 0.302f
C665 out.t91 vss 0.302f
C666 out.t239 vss 0.302f
C667 out.t129 vss 0.302f
C668 out.t170 vss 0.302f
C669 out.t130 vss 0.302f
C670 out.t214 vss 0.302f
C671 out.t84 vss 0.538f
C672 out.n185 vss 0.29f
C673 out.n186 vss 0.29f
C674 out.n187 vss 0.29f
C675 out.n188 vss 0.29f
C676 out.n189 vss 0.29f
C677 out.n190 vss 0.29f
C678 out.n191 vss 0.29f
C679 out.n192 vss 0.29f
C680 out.n193 vss 0.253f
C681 out.t157 vss 0.302f
C682 out.t296 vss 0.302f
C683 out.t331 vss 0.302f
C684 out.t292 vss 0.302f
C685 out.t287 vss 0.302f
C686 out.t301 vss 0.302f
C687 out.t328 vss 0.302f
C688 out.t320 vss 0.302f
C689 out.t325 vss 0.302f
C690 out.t23 vss 0.538f
C691 out.n194 vss 0.29f
C692 out.n195 vss 0.29f
C693 out.n196 vss 0.29f
C694 out.n197 vss 0.29f
C695 out.n198 vss 0.29f
C696 out.n199 vss 0.29f
C697 out.n200 vss 0.29f
C698 out.n201 vss 0.29f
C699 out.n202 vss 0.253f
C700 out.t63 vss 0.302f
C701 out.t332 vss 0.302f
C702 out.t330 vss 0.302f
C703 out.t67 vss 0.302f
C704 out.t88 vss 0.302f
C705 out.t106 vss 0.302f
C706 out.t107 vss 0.302f
C707 out.t334 vss 0.302f
C708 out.t126 vss 0.302f
C709 out.t142 vss 0.538f
C710 out.n203 vss 0.29f
C711 out.n204 vss 0.29f
C712 out.n205 vss 0.29f
C713 out.n206 vss 0.29f
C714 out.n207 vss 0.29f
C715 out.n208 vss 0.29f
C716 out.n209 vss 0.29f
C717 out.n210 vss 0.29f
C718 out.n211 vss 0.253f
C719 out.t48 vss 0.302f
C720 out.t195 vss 0.302f
C721 out.t210 vss 0.302f
C722 out.t148 vss 0.302f
C723 out.t167 vss 0.302f
C724 out.t183 vss 0.302f
C725 out.t251 vss 0.302f
C726 out.t110 vss 0.302f
C727 out.t92 vss 0.302f
C728 out.t192 vss 0.538f
C729 out.n212 vss 0.29f
C730 out.n213 vss 0.29f
C731 out.n214 vss 0.29f
C732 out.n215 vss 0.29f
C733 out.n216 vss 0.29f
C734 out.n217 vss 0.29f
C735 out.n218 vss 0.29f
C736 out.n219 vss 0.29f
C737 out.n220 vss 0.253f
C738 out.t35 vss 0.302f
C739 out.t253 vss 0.302f
C740 out.t260 vss 0.302f
C741 out.t244 vss 0.302f
C742 out.t233 vss 0.302f
C743 out.t219 vss 0.302f
C744 out.t204 vss 0.302f
C745 out.t203 vss 0.302f
C746 out.t220 vss 0.302f
C747 out.t179 vss 0.538f
C748 out.n221 vss 0.29f
C749 out.n222 vss 0.29f
C750 out.n223 vss 0.29f
C751 out.n224 vss 0.29f
C752 out.n225 vss 0.29f
C753 out.n226 vss 0.29f
C754 out.n227 vss 0.29f
C755 out.n228 vss 0.29f
C756 out.n229 vss 0.253f
C757 out.t80 vss 0.302f
C758 out.t319 vss 0.302f
C759 out.t322 vss 0.302f
C760 out.t173 vss 0.302f
C761 out.t311 vss 0.302f
C762 out.t43 vss 0.302f
C763 out.t155 vss 0.302f
C764 out.t315 vss 0.302f
C765 out.t310 vss 0.302f
C766 out.t161 vss 0.538f
C767 out.n230 vss 0.29f
C768 out.n231 vss 0.29f
C769 out.n232 vss 0.29f
C770 out.n233 vss 0.29f
C771 out.n234 vss 0.29f
C772 out.n235 vss 0.29f
C773 out.n236 vss 0.29f
C774 out.n237 vss 0.29f
C775 out.n238 vss 0.253f
C776 out.t174 vss 0.302f
C777 out.t305 vss 0.302f
C778 out.t300 vss 0.302f
C779 out.t136 vss 0.302f
C780 out.t323 vss 0.302f
C781 out.t306 vss 0.302f
C782 out.t116 vss 0.302f
C783 out.t290 vss 0.302f
C784 out.t295 vss 0.302f
C785 out.t108 vss 0.538f
C786 out.n239 vss 0.29f
C787 out.n240 vss 0.29f
C788 out.n241 vss 0.29f
C789 out.n242 vss 0.29f
C790 out.n243 vss 0.29f
C791 out.n244 vss 0.29f
C792 out.n245 vss 0.29f
C793 out.n246 vss 0.29f
C794 out.n247 vss 0.253f
C795 out.t158 vss 0.302f
C796 out.t188 vss 0.302f
C797 out.t172 vss 0.302f
C798 out.t153 vss 0.302f
C799 out.t113 vss 0.302f
C800 out.t133 vss 0.302f
C801 out.t94 vss 0.302f
C802 out.t75 vss 0.302f
C803 out.t58 vss 0.302f
C804 out.t89 vss 0.538f
C805 out.n248 vss 0.29f
C806 out.n249 vss 0.29f
C807 out.n250 vss 0.29f
C808 out.n251 vss 0.29f
C809 out.n252 vss 0.29f
C810 out.n253 vss 0.29f
C811 out.n254 vss 0.29f
C812 out.n255 vss 0.29f
C813 out.n256 vss 0.253f
C814 out.t205 vss 0.302f
C815 out.t165 vss 0.302f
C816 out.t182 vss 0.302f
C817 out.t149 vss 0.302f
C818 out.t168 vss 0.302f
C819 out.t270 vss 0.302f
C820 out.t298 vss 0.302f
C821 out.t293 vss 0.302f
C822 out.t288 vss 0.302f
C823 out.t72 vss 0.538f
C824 out.n257 vss 0.29f
C825 out.n258 vss 0.29f
C826 out.n259 vss 0.29f
C827 out.n260 vss 0.29f
C828 out.n261 vss 0.29f
C829 out.n262 vss 0.29f
C830 out.n263 vss 0.29f
C831 out.n264 vss 0.29f
C832 out.n265 vss 0.253f
C833 out.t189 vss 0.302f
C834 out.t338 vss 0.302f
C835 out.t5 vss 0.302f
C836 out.t52 vss 0.302f
C837 out.t25 vss 0.302f
C838 out.t40 vss 0.302f
C839 out.t93 vss 0.302f
C840 out.t74 vss 0.302f
C841 out.t57 vss 0.302f
C842 out.t56 vss 0.538f
C843 out.n266 vss 0.29f
C844 out.n267 vss 0.29f
C845 out.n268 vss 0.29f
C846 out.n269 vss 0.29f
C847 out.n270 vss 0.29f
C848 out.n271 vss 0.29f
C849 out.n272 vss 0.29f
C850 out.n273 vss 0.29f
C851 out.n274 vss 0.253f
C852 out.t221 vss 0.302f
C853 out.t289 vss 0.302f
C854 out.t294 vss 0.302f
C855 out.t304 vss 0.302f
C856 out.t309 vss 0.302f
C857 out.t299 vss 0.302f
C858 out.t285 vss 0.302f
C859 out.t277 vss 0.302f
C860 out.t281 vss 0.302f
C861 out.t180 vss 0.538f
C862 out.n275 vss 0.29f
C863 out.n276 vss 0.29f
C864 out.n277 vss 0.29f
C865 out.n278 vss 0.29f
C866 out.n279 vss 0.29f
C867 out.n280 vss 0.29f
C868 out.n281 vss 0.29f
C869 out.n282 vss 0.29f
C870 out.n283 vss 0.253f
C871 out.t139 vss 0.302f
C872 out.t147 vss 0.302f
C873 out.t255 vss 0.302f
C874 out.t237 vss 0.302f
C875 out.t212 vss 0.302f
C876 out.t184 vss 0.302f
C877 out.t272 vss 0.302f
C878 out.t261 vss 0.302f
C879 out.t280 vss 0.302f
C880 out.t164 vss 0.538f
C881 out.n284 vss 0.29f
C882 out.n285 vss 0.29f
C883 out.n286 vss 0.29f
C884 out.n287 vss 0.29f
C885 out.n288 vss 0.29f
C886 out.n289 vss 0.29f
C887 out.n290 vss 0.29f
C888 out.n291 vss 0.29f
C889 out.n292 vss 0.253f
C890 out.t118 vss 0.302f
C891 out.t128 vss 0.302f
C892 out.t263 vss 0.302f
C893 out.t247 vss 0.302f
C894 out.t227 vss 0.302f
C895 out.t197 vss 0.302f
C896 out.t276 vss 0.302f
C897 out.t267 vss 0.302f
C898 out.t284 vss 0.302f
C899 out.t146 vss 0.538f
C900 out.n293 vss 0.29f
C901 out.n294 vss 0.29f
C902 out.n295 vss 0.29f
C903 out.n296 vss 0.29f
C904 out.n297 vss 0.29f
C905 out.n298 vss 0.29f
C906 out.n299 vss 0.29f
C907 out.n300 vss 0.29f
C908 out.n301 vss 0.253f
C909 out.t99 vss 0.302f
C910 out.t124 vss 0.302f
C911 out.t145 vss 0.302f
C912 out.t104 vss 0.302f
C913 out.t85 vss 0.302f
C914 out.t70 vss 0.302f
C915 out.t29 vss 0.302f
C916 out.t17 vss 0.302f
C917 out.t42 vss 0.302f
C918 out.t127 vss 0.538f
C919 out.n302 vss 0.29f
C920 out.n303 vss 0.29f
C921 out.n304 vss 0.29f
C922 out.n305 vss 0.29f
C923 out.n306 vss 0.29f
C924 out.n307 vss 0.29f
C925 out.n308 vss 0.29f
C926 out.n309 vss 0.29f
C927 out.n310 vss 0.253f
C928 out.t49 vss 0.302f
C929 out.t297 vss 0.302f
C930 out.t291 vss 0.302f
C931 out.t318 vss 0.302f
C932 out.t314 vss 0.302f
C933 out.t316 vss 0.302f
C934 out.t303 vss 0.302f
C935 out.t308 vss 0.302f
C936 out.t313 vss 0.302f
C937 out.t66 vss 0.538f
C938 out.n311 vss 0.29f
C939 out.n312 vss 0.29f
C940 out.n313 vss 0.29f
C941 out.n314 vss 0.29f
C942 out.n315 vss 0.29f
C943 out.n316 vss 0.29f
C944 out.n317 vss 0.29f
C945 out.n318 vss 0.29f
C946 out.n319 vss 0.253f
C947 out.t64 vss 0.302f
C948 out.t166 vss 0.302f
C949 out.t196 vss 0.302f
C950 out.t264 vss 0.302f
C951 out.t248 vss 0.302f
C952 out.t274 vss 0.302f
C953 out.t266 vss 0.302f
C954 out.t282 vss 0.302f
C955 out.t275 vss 0.302f
C956 out.t103 vss 0.538f
C957 out.n320 vss 0.29f
C958 out.n321 vss 0.29f
C959 out.n322 vss 0.29f
C960 out.n323 vss 0.29f
C961 out.n324 vss 0.29f
C962 out.n325 vss 0.29f
C963 out.n326 vss 0.29f
C964 out.n327 vss 0.29f
C965 out.n328 vss 0.253f
C966 out.t234 vss 0.302f
C967 out.t181 vss 0.302f
C968 out.t211 vss 0.302f
C969 out.t269 vss 0.302f
C970 out.t257 vss 0.302f
C971 out.t278 vss 0.302f
C972 out.t271 vss 0.302f
C973 out.t200 vss 0.302f
C974 out.t279 vss 0.302f
C975 out.t209 vss 0.538f
C976 out.n329 vss 0.29f
C977 out.n330 vss 0.29f
C978 out.n331 vss 0.29f
C979 out.n332 vss 0.29f
C980 out.n333 vss 0.29f
C981 out.n334 vss 0.29f
C982 out.n335 vss 0.29f
C983 out.n336 vss 0.29f
C984 out.n337 vss 0.253f
C985 out.t222 vss 0.302f
C986 out.t3 vss 0.302f
C987 out.t12 vss 0.302f
C988 out.t38 vss 0.302f
C989 out.t68 vss 0.302f
C990 out.t54 vss 0.302f
C991 out.t171 vss 0.302f
C992 out.t27 vss 0.302f
C993 out.t13 vss 0.302f
C994 out.t194 vss 0.538f
C995 out.n338 vss 0.29f
C996 out.n339 vss 0.29f
C997 out.n340 vss 0.29f
C998 out.n341 vss 0.29f
C999 out.n342 vss 0.29f
C1000 out.n343 vss 0.29f
C1001 out.n344 vss 0.29f
C1002 out.n345 vss 0.29f
C1003 out.n346 vss 0.253f
C1004 out.t81 vss 0.302f
C1005 out.t236 vss 0.302f
C1006 out.t246 vss 0.302f
C1007 out.t256 vss 0.302f
C1008 out.t265 vss 0.302f
C1009 out.t228 vss 0.302f
C1010 out.t232 vss 0.302f
C1011 out.t217 vss 0.302f
C1012 out.t241 vss 0.302f
C1013 out.t235 vss 0.538f
C1014 out.n347 vss 0.29f
C1015 out.n348 vss 0.29f
C1016 out.n349 vss 0.29f
C1017 out.n350 vss 0.29f
C1018 out.n351 vss 0.29f
C1019 out.n352 vss 0.29f
C1020 out.n353 vss 0.29f
C1021 out.n354 vss 0.29f
C1022 out.n355 vss 0.253f
C1023 out.t206 vss 0.302f
C1024 out.t262 vss 0.302f
C1025 out.t273 vss 0.302f
C1026 out.t225 vss 0.302f
C1027 out.t249 vss 0.302f
C1028 out.t185 vss 0.302f
C1029 out.t302 vss 0.302f
C1030 out.t216 vss 0.302f
C1031 out.t258 vss 0.302f
C1032 out.t176 vss 0.538f
C1033 out.n356 vss 0.29f
C1034 out.n357 vss 0.29f
C1035 out.n358 vss 0.29f
C1036 out.n359 vss 0.29f
C1037 out.n360 vss 0.29f
C1038 out.n361 vss 0.29f
C1039 out.n362 vss 0.29f
C1040 out.n363 vss 0.29f
C1041 out.n364 vss 0.253f
C1042 out.t190 vss 0.302f
C1043 out.t144 vss 0.302f
C1044 out.t163 vss 0.302f
C1045 out.t105 vss 0.302f
C1046 out.t125 vss 0.302f
C1047 out.t86 vss 0.302f
C1048 out.t132 vss 0.302f
C1049 out.t112 vss 0.302f
C1050 out.t152 vss 0.302f
C1051 out.t162 vss 0.538f
C1052 out.n365 vss 0.29f
C1053 out.n366 vss 0.29f
C1054 out.n367 vss 0.29f
C1055 out.n368 vss 0.29f
C1056 out.n369 vss 0.29f
C1057 out.n370 vss 0.29f
C1058 out.n371 vss 0.29f
C1059 out.n372 vss 0.29f
C1060 out.n373 vss 0.253f
C1061 out.t159 vss 0.302f
C1062 out.t254 vss 0.302f
C1063 out.t268 vss 0.302f
C1064 out.t238 vss 0.302f
C1065 out.t213 vss 0.302f
C1066 out.t198 vss 0.302f
C1067 out.t250 vss 0.302f
C1068 out.t230 vss 0.302f
C1069 out.t240 vss 0.302f
C1070 out.t143 vss 0.538f
C1071 out.n374 vss 0.29f
C1072 out.n375 vss 0.29f
C1073 out.n376 vss 0.29f
C1074 out.n377 vss 0.29f
C1075 out.n378 vss 0.29f
C1076 out.n379 vss 0.29f
C1077 out.n380 vss 0.29f
C1078 out.n381 vss 0.29f
C1079 out.n382 vss 0.253f
C1080 out.t175 vss 0.302f
C1081 out.t119 vss 0.302f
C1082 out.t140 vss 0.302f
C1083 out.t100 vss 0.302f
C1084 out.t245 vss 0.302f
C1085 out.t79 vss 0.302f
C1086 out.t207 vss 0.302f
C1087 out.t193 vss 0.302f
C1088 out.t223 vss 0.302f
C1089 out.t123 vss 0.538f
C1090 out.n383 vss 0.29f
C1091 out.n384 vss 0.29f
C1092 out.n385 vss 0.29f
C1093 out.n386 vss 0.29f
C1094 out.n387 vss 0.29f
C1095 out.n388 vss 0.29f
C1096 out.n389 vss 0.29f
C1097 out.n390 vss 0.29f
C1098 out.n391 vss 0.253f
C1099 out.n392 vss 0.161f
C1100 out.n393 vss 0.279f
C1101 out.n394 vss 0.279f
C1102 out.n395 vss 0.279f
C1103 out.n396 vss 0.279f
C1104 out.n397 vss 0.279f
C1105 out.n398 vss 0.279f
C1106 out.n399 vss 0.279f
C1107 out.n400 vss 0.279f
C1108 out.n401 vss 0.279f
C1109 out.n402 vss 0.279f
C1110 out.n403 vss 0.279f
C1111 out.n404 vss 0.279f
C1112 out.n405 vss 0.279f
C1113 out.n406 vss 0.279f
C1114 out.n407 vss 0.279f
C1115 out.n408 vss 0.279f
C1116 out.n409 vss 0.279f
C1117 out.n410 vss 0.279f
C1118 out.n411 vss 0.279f
C1119 out.n412 vss 0.279f
C1120 out.n413 vss 0.279f
C1121 out.n414 vss 0.279f
C1122 out.n415 vss 0.279f
C1123 out.n416 vss 0.279f
C1124 out.n417 vss 0.279f
C1125 out.n418 vss 0.279f
C1126 out.n419 vss 0.279f
C1127 out.n420 vss 0.279f
C1128 out.n421 vss 0.279f
C1129 out.n422 vss 0.279f
C1130 out.n423 vss 0.279f
C1131 out.n424 vss 0.279f
C1132 out.n425 vss 0.189f
C1133 ctl7 vss 0.362f
C1134 ctl2 vss 0.509f
C1135 sw_top_3/m2_990_200# vss 1.81f
C1136 sw_top_3/m2_1158_361# vss 1.69f
C1137 dum vss 0.493f
C1138 ctl3 vss 0.362f
C1139 en_buf vss 3.48f
C1140 enb vss 3.17f
C1141 carray_0/n1 vss 4.01f
C1142 carray_0/n5 vss 17.2f
C1143 carray_0/n4 vss 8.48f
C1144 carray_0/n3 vss 6.16f
C1145 carray_0/m3_42700_1156# vss 1.78f
C1146 carray_0/m3_42500_1156# vss 1.02f
C1147 carray_0/m3_900_1156# vss 1.76f
C1148 carray_0/m2_42800_1156# vss 2.03f
C1149 carray_0/m2_41500_1156# vss 1.43f
C1150 carray_0/m2_40200_1156# vss 1.43f
C1151 carray_0/m2_38900_1156# vss 1.43f
C1152 carray_0/m2_37600_1156# vss 1.43f
C1153 carray_0/m2_36300_1156# vss 1.43f
C1154 carray_0/m2_35000_1156# vss 1.43f
C1155 carray_0/m2_33700_1156# vss 1.43f
C1156 carray_0/m2_32400_1156# vss 1.43f
C1157 carray_0/m2_31100_1156# vss 1.43f
C1158 carray_0/m2_29800_1156# vss 1.43f
C1159 carray_0/m2_28500_1156# vss 1.43f
C1160 carray_0/m2_27200_1156# vss 1.43f
C1161 carray_0/m2_25900_1156# vss 1.43f
C1162 carray_0/m2_24600_1156# vss 1.43f
C1163 carray_0/m2_23300_1156# vss 1.42f
C1164 carray_0/m2_800_1156# vss 2.03f
C1165 carray_0/via23_4_200/m2_1_40# vss 0.372f
C1166 carray_0/via23_4_414/m2_1_40# vss 0.372f
C1167 carray_0/via23_4_447/m2_1_40# vss 0.291f
C1168 carray_0/via23_4_458/m2_1_40# vss 0.291f
C1169 carray_0/via23_4_446/m2_1_40# vss 0.291f
C1170 carray_0/via23_4_460/m2_1_40# vss 0.291f
C1171 carray_0/via23_4_220/m2_1_40# vss 0.372f
C1172 carray_0/via23_4_9/m2_1_40# vss 0.364f
C1173 carray_0/via23_4_459/m2_1_40# vss 0.28f
C1174 carray_0/via23_4_641/m2_1_40# vss 0.372f
C1175 carray_0/via23_4_455/m2_1_40# vss 0.243f
C1176 carray_0/via23_4_635/m2_1_40# vss 0.372f
C1177 carray_0/via23_4_601/m2_1_40# vss 0.373f
C1178 carray_0/via23_4_676/m2_1_40# vss 0.373f
C1179 carray_0/n0 vss 3.04f
C1180 carray_0/via23_4_3/m2_1_40# vss 0.253f
C1181 carray_0/via23_4_642/m2_1_40# vss 0.372f
C1182 carray_0/via23_4_709/m2_1_40# vss 0.373f
C1183 carray_0/via23_4_678/m2_1_40# vss 0.485f
C1184 carray_0/via23_4_117/m2_1_40# vss 0.372f
C1185 carray_0/via23_4_128/m2_1_40# vss 0.372f
C1186 carray_0/via23_4_677/m2_1_40# vss 0.373f
C1187 carray_0/via23_4_21/m2_1_40# vss 0.253f
C1188 carray_0/via23_4_103/m2_1_40# vss 0.253f
C1189 carray_0/via23_4_20/m2_1_40# vss 0.253f
C1190 carray_0/via23_4_91/m2_1_40# vss 0.253f
C1191 carray_0/via23_4_326/m2_1_40# vss 0.485f
C1192 carray_0/via23_4_111/m2_1_40# vss 0.372f
C1193 carray_0/via23_4_198/m2_1_40# vss 0.372f
C1194 carray_0/via23_4_379/m2_1_40# vss 0.3f
C1195 carray_0/via23_4_346/m2_1_40# vss 0.485f
C1196 carray_0/via23_4_1/m2_1_40# vss 0.253f
C1197 carray_0/via23_4_712/m2_1_40# vss 0.373f
C1198 carray_0/via23_4_199/m2_1_40# vss 0.372f
C1199 carray_0/via23_4_378/m2_1_40# vss 0.3f
C1200 carray_0/via23_4_334/m2_1_40# vss 0.373f
C1201 carray_0/via23_4_345/m2_1_40# vss 0.373f
C1202 carray_0/via23_4_89/m2_1_40# vss 0.364f
C1203 carray_0/via23_4_23/m2_1_40# vss 0.253f
C1204 carray_0/via23_4_711/m2_1_40# vss 0.373f
C1205 carray_0/via23_4_250/m2_1_40# vss 0.373f
C1206 carray_0/via23_4_333/m2_1_40# vss 0.373f
C1207 carray_0/n7 vss 65.5f
C1208 carray_0/via23_4_22/m2_1_40# vss 0.253f
C1209 carray_0/via23_4_710/m2_1_40# vss 0.373f
C1210 carray_0/via23_4_249/m2_1_40# vss 0.373f
C1211 carray_0/via23_4_367/m2_1_40# vss 0.509f
C1212 carray_0/via23_4_332/m2_1_40# vss 0.373f
C1213 carray_0/via23_4_2/m2_1_40# vss 0.243f
C1214 carray_0/via23_4_87/m2_1_40# vss 0.253f
C1215 carray_0/via23_4_705/m2_1_40# vss 0.372f
C1216 carray_0/via23_4_366/m2_1_40# vss 0.308f
C1217 carray_0/via23_4_331/m2_1_40# vss 0.373f
C1218 carray_0/via23_4_354/m2_1_40# vss 0.373f
C1219 carray_0/n6 vss 32.2f
C1220 carray_0/via23_4_88/m2_1_40# vss 0.253f
C1221 carray_0/via23_4_704/m2_1_40# vss 0.372f
C1222 carray_0/via23_4_369/m2_1_40# vss 0.3f
C1223 carray_0/via23_4_96/m2_1_40# vss 0.388f
C1224 carray_0/via23_4_368/m2_1_40# vss 0.3f
C1225 carray_0/via23_4_598/m2_1_40# vss 0.373f
C1226 carray_0/via23_4_95/m2_1_40# vss 0.253f
C1227 carray_0/via23_4_702/m2_1_40# vss 0.509f
C1228 carray_0/via23_4_347/m2_1_40# vss 0.373f
C1229 carray_0/via23_4_94/m2_1_40# vss 0.253f
C1230 carray_0/n2 vss 8.06f
C1231 carray_0/via23_4_675/m2_1_40# vss 0.373f
C1232 carray_0/via23_4_588/m2_1_40# vss 0.373f
C1233 out vss 39f
C1234 carray_0/via23_4_381/m2_1_40# vss 0.3f
C1235 carray_0/via23_4_600/m2_1_40# vss 0.373f
C1236 carray_0/via23_4_380/m2_1_40# vss 0.411f
C1237 carray_0/via23_4_584/m2_1_40# vss 0.373f
C1238 carray_0/via23_4_599/m2_1_40# vss 0.485f
C1239 carray_0/via23_4_245/m2_1_40# vss 0.373f
C1240 carray_0/via23_4_90/m2_1_40# vss 0.253f
C1241 carray_0/via23_4_218/m2_1_40# vss 0.373f
C1242 carray_0/via23_4_251/m2_1_40# vss 0.373f
C1243 carray_0/via23_4_590/m2_1_40# vss 0.373f
C1244 carray_0/via23_4_230/m2_1_40# vss 0.373f
C1245 carray_0/via23_4_589/m2_1_40# vss 0.373f
C1246 carray_0/ndum vss 6.61f
C1247 carray_0/via23_4_228/m2_1_40# vss 0.509f
C1248 carray_0/via23_4_229/m2_1_40# vss 0.373f
C1249 carray_0/via23_4_419/m2_1_40# vss 0.372f
C1250 carray_0/via23_4_439/m2_1_40# vss 0.291f
C1251 carray_0/via23_4_429/m2_1_40# vss 0.372f
C1252 carray_0/via23_4_449/m2_1_40# vss 0.402f
C1253 carray_0/via23_4_213/m2_1_40# vss 0.372f
C1254 carray_0/via23_4_448/m2_1_40# vss 0.291f
C1255 ctl4 vss 0.362f
C1256 sample vss 32.3f
C1257 sw_top_0/m2_990_200# vss 1.81f
C1258 vin vss 17.2f
C1259 sw_top_0/m2_1158_361# vss 1.69f
C1260 ctl5 vss 0.362f
C1261 vdd vss 46.8f
C1262 ctl1 vss 0.363f
C1263 ctl0 vss 0.363f
C1264 ctl6 vss 0.362f
.ends
