magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 314 542
<< pwell >>
rect 1 -19 271 163
rect 30 -57 64 -19
<< scnmos >>
rect 79 7 109 137
rect 163 7 193 137
<< scpmoshvt >>
rect 79 257 109 457
rect 151 257 181 457
<< ndiff >>
rect 27 123 79 137
rect 27 89 35 123
rect 69 89 79 123
rect 27 55 79 89
rect 27 21 35 55
rect 69 21 79 55
rect 27 7 79 21
rect 109 123 163 137
rect 109 89 119 123
rect 153 89 163 123
rect 109 55 163 89
rect 109 21 119 55
rect 153 21 163 55
rect 109 7 163 21
rect 193 123 245 137
rect 193 89 203 123
rect 237 89 245 123
rect 193 55 245 89
rect 193 21 203 55
rect 237 21 245 55
rect 193 7 245 21
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 377 79 411
rect 27 343 35 377
rect 69 343 79 377
rect 27 309 79 343
rect 27 275 35 309
rect 69 275 79 309
rect 27 257 79 275
rect 109 257 151 457
rect 181 445 233 457
rect 181 411 191 445
rect 225 411 233 445
rect 181 377 233 411
rect 181 343 191 377
rect 225 343 233 377
rect 181 309 233 343
rect 181 275 191 309
rect 225 275 233 309
rect 181 257 233 275
<< ndiffc >>
rect 35 89 69 123
rect 35 21 69 55
rect 119 89 153 123
rect 119 21 153 55
rect 203 89 237 123
rect 203 21 237 55
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 35 275 69 309
rect 191 411 225 445
rect 191 343 225 377
rect 191 275 225 309
<< poly >>
rect 79 457 109 483
rect 151 457 181 483
rect 79 225 109 257
rect 22 209 109 225
rect 22 175 37 209
rect 71 175 109 209
rect 151 225 181 257
rect 151 209 255 225
rect 151 195 205 209
rect 22 159 109 175
rect 79 137 109 159
rect 163 175 205 195
rect 239 175 255 209
rect 163 159 255 175
rect 163 137 193 159
rect 79 -19 109 7
rect 163 -19 193 7
<< polycont >>
rect 37 175 71 209
rect 205 175 239 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 276 521
rect 19 445 85 450
rect 19 411 35 445
rect 69 411 85 445
rect 19 377 85 411
rect 19 343 35 377
rect 69 343 85 377
rect 19 309 85 343
rect 19 275 35 309
rect 69 293 85 309
rect 191 445 257 487
rect 225 411 257 445
rect 191 377 257 411
rect 225 343 257 377
rect 191 309 257 343
rect 69 275 155 293
rect 19 259 155 275
rect 225 275 257 309
rect 191 259 257 275
rect 17 209 87 225
rect 17 175 37 209
rect 71 175 87 209
rect 121 139 155 259
rect 189 209 259 225
rect 189 175 205 209
rect 239 175 259 209
rect 21 123 69 139
rect 21 89 35 123
rect 21 55 69 89
rect 21 21 35 55
rect 21 -23 69 21
rect 103 123 169 139
rect 103 89 119 123
rect 153 89 169 123
rect 103 55 169 89
rect 103 21 119 55
rect 153 21 169 55
rect 103 11 169 21
rect 203 123 257 139
rect 237 89 257 123
rect 203 55 257 89
rect 237 21 257 55
rect 203 -23 257 21
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 276 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
<< metal1 >>
rect 0 521 276 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 276 521
rect 0 456 276 487
rect 0 -23 276 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 276 -23
rect 0 -88 276 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 nor2_1
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 29 181 63 215 0 FreeSans 200 0 0 0 B
port 8 nsew
flabel locali s 30 385 64 419 0 FreeSans 200 0 0 0 Y
port 9 nsew
flabel locali s 213 181 247 215 0 FreeSans 200 0 0 0 A
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 276 504
string path 0.000 -1.000 6.900 -1.000 
<< end >>
