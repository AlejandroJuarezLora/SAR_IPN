* SPICE3 file created from sarlogic.ext - technology: sky130B

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X a_150_297# a_68_297#
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_68_297# a_150_297# 0.00477f
C1 X a_150_297# 4.96e-19
C2 VPB a_68_297# 0.0611f
C3 B A 0.0751f
C4 VPWR A 0.00846f
C5 VPB X 0.0209f
C6 B VGND 0.0437f
C7 VPWR VGND 0.0464f
C8 a_150_297# VGND 4.62e-19
C9 VPB A 0.031f
C10 VPWR B 0.00855f
C11 X a_68_297# 0.105f
C12 VPB VGND 0.0112f
C13 VPWR a_150_297# 0.00193f
C14 VPB B 0.0462f
C15 A a_68_297# 0.158f
C16 VPB VPWR 0.0805f
C17 A X 0.0131f
C18 a_68_297# VGND 0.118f
C19 X VGND 0.114f
C20 B a_68_297# 0.0984f
C21 VPWR a_68_297# 0.089f
C22 B X 1.65e-19
C23 VPWR X 0.129f
C24 A VGND 0.0347f
C25 VGND VNB 0.32f
C26 X VNB 0.101f
C27 A VNB 0.111f
C28 B VNB 0.183f
C29 VPWR VNB 0.269f
C30 VPB VNB 0.516f
C31 a_68_297# VNB 0.154f
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
C0 VGND VPWR 0.353f
C1 VPB VPWR 0.0625f
C2 VPB VGND 0.0797f
C3 VPWR VNB 0.47f
C4 VGND VNB 0.427f
C5 VPB VNB 0.339f
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
C0 VGND VPWR 1.57f
C1 VPB VPWR 0.137f
C2 VPB VGND 0.35f
C3 VPWR VNB 1.67f
C4 VGND VNB 1.47f
C5 VPB VNB 1.14f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X a_75_212#
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 VPB A 0.0525f
C1 a_75_212# X 0.107f
C2 X VGND 0.0545f
C3 VPB VPWR 0.0355f
C4 a_75_212# A 0.178f
C5 A VGND 0.0184f
C6 a_75_212# VPWR 0.134f
C7 VGND VPWR 0.0289f
C8 a_75_212# VPB 0.0571f
C9 VPB VGND 0.00507f
C10 A X 8.48e-19
C11 X VPWR 0.0896f
C12 VPB X 0.0128f
C13 a_75_212# VGND 0.105f
C14 A VPWR 0.0217f
C15 VGND VNB 0.207f
C16 VPWR VNB 0.176f
C17 X VNB 0.0942f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_75_212# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X a_80_21# a_209_297#
+ a_209_47# a_303_47#
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
C0 A2 X 3.42e-19
C1 A1 B1 0.101f
C2 a_209_297# a_303_47# 1.26e-19
C3 VGND X 0.0572f
C4 a_209_297# B1 0.00622f
C5 a_80_21# X 0.0765f
C6 A3 X 0.00625f
C7 VPB X 0.0108f
C8 X VPWR 0.117f
C9 a_303_47# A2 3.38e-19
C10 a_209_297# A1 0.0378f
C11 a_303_47# VGND 0.00661f
C12 a_209_297# a_209_47# 6.96e-20
C13 a_80_21# a_303_47# 0.0115f
C14 VGND B1 0.0172f
C15 a_80_21# B1 0.111f
C16 VPB B1 0.0342f
C17 a_303_47# VPWR 0.00105f
C18 B1 VPWR 0.0177f
C19 A2 A1 0.104f
C20 VGND A1 0.0135f
C21 a_80_21# A1 0.0367f
C22 a_209_297# A2 0.0366f
C23 VPB A1 0.0287f
C24 a_209_47# VGND 0.00696f
C25 a_209_297# VGND 0.0043f
C26 a_80_21# a_209_47# 0.0101f
C27 A3 a_209_47# 3.56e-19
C28 a_80_21# a_209_297# 0.0626f
C29 A1 VPWR 0.018f
C30 A3 a_209_297# 0.0268f
C31 a_209_297# VPB 0.00284f
C32 a_303_47# X 6.01e-19
C33 a_209_47# VPWR 0.00102f
C34 a_209_297# VPWR 0.205f
C35 VGND A2 0.0148f
C36 a_80_21# A2 0.0357f
C37 A3 A2 0.109f
C38 VPB A2 0.0285f
C39 a_80_21# VGND 0.216f
C40 A3 VGND 0.0169f
C41 VPB VGND 0.00769f
C42 A2 VPWR 0.0227f
C43 A1 X 1.56e-19
C44 A3 a_80_21# 0.117f
C45 a_80_21# VPB 0.051f
C46 A3 VPB 0.0297f
C47 VGND VPWR 0.0662f
C48 a_209_47# X 9.76e-19
C49 a_80_21# VPWR 0.0992f
C50 A3 VPWR 0.0403f
C51 VPB VPWR 0.0715f
C52 VGND VNB 0.41f
C53 VPWR VNB 0.332f
C54 X VNB 0.0895f
C55 B1 VNB 0.115f
C56 A1 VNB 0.0897f
C57 A2 VNB 0.0896f
C58 A3 VNB 0.0899f
C59 VPB VNB 0.693f
C60 a_209_297# VNB 0.00621f
C61 a_80_21# VNB 0.211f
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q a_1462_47# a_543_47#
+ a_651_413# a_193_47# a_805_47# a_448_47# a_639_47# a_1283_21# a_761_289# a_1108_47#
+ a_1217_47# a_1270_413# a_27_47#
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
C0 RESET_B a_1283_21# 0.278f
C1 a_1217_47# a_761_289# 4.2e-19
C2 VGND Q 0.0616f
C3 Q a_1108_47# 9.8e-19
C4 a_761_289# a_543_47# 0.21f
C5 a_193_47# a_1283_21# 0.0424f
C6 VPWR a_1283_21# 0.209f
C7 a_805_47# a_543_47# 0.00171f
C8 a_639_47# a_543_47# 0.0138f
C9 VPB a_761_289# 0.0994f
C10 VPB CLK 0.0693f
C11 a_27_47# a_1283_21# 0.0436f
C12 a_1462_47# VGND 0.00221f
C13 D a_543_47# 7.35e-20
C14 VGND a_1283_21# 0.24f
C15 a_1283_21# a_1108_47# 0.234f
C16 a_1217_47# RESET_B 6.03e-19
C17 VPB D 0.138f
C18 RESET_B a_543_47# 0.153f
C19 a_805_47# a_761_289# 3.69e-19
C20 a_1217_47# a_193_47# 2.36e-20
C21 a_639_47# a_761_289# 3.16e-19
C22 Q a_1283_21# 0.0598f
C23 a_193_47# a_543_47# 0.23f
C24 VPB RESET_B 0.138f
C25 a_27_47# a_1217_47# 2.56e-19
C26 a_448_47# a_543_47# 0.0498f
C27 VPWR a_543_47# 0.1f
C28 VPB a_193_47# 0.171f
C29 a_27_47# a_543_47# 0.115f
C30 a_651_413# a_543_47# 0.0572f
C31 a_1217_47# VGND 9.68e-19
C32 a_1462_47# a_1283_21# 0.0074f
C33 a_1217_47# a_1108_47# 0.00742f
C34 RESET_B a_761_289# 0.166f
C35 VPB VPWR 0.216f
C36 CLK RESET_B 1.09e-19
C37 a_448_47# VPB 0.0141f
C38 VGND a_543_47# 0.123f
C39 a_543_47# a_1108_47# 7.99e-20
C40 a_27_47# VPB 0.262f
C41 a_805_47# RESET_B 0.00316f
C42 a_651_413# VPB 0.0135f
C43 CLK a_193_47# 7.94e-19
C44 a_193_47# a_761_289# 0.186f
C45 a_639_47# RESET_B 9.54e-19
C46 CLK VPWR 0.0174f
C47 D RESET_B 4.72e-19
C48 VPB VGND 0.00999f
C49 VPWR a_761_289# 0.105f
C50 VPB a_1108_47# 0.113f
C51 a_1270_413# a_761_289# 2.6e-19
C52 a_639_47# a_193_47# 2.28e-19
C53 a_27_47# CLK 0.234f
C54 a_27_47# a_761_289# 0.0701f
C55 a_651_413# a_761_289# 0.0977f
C56 D a_193_47# 0.218f
C57 a_639_47# a_448_47# 4.61e-19
C58 a_448_47# D 0.156f
C59 D VPWR 0.0812f
C60 VGND a_761_289# 0.0734f
C61 VPB Q 0.011f
C62 CLK VGND 0.0172f
C63 a_761_289# a_1108_47# 0.0512f
C64 a_27_47# a_639_47# 0.00188f
C65 a_27_47# D 0.133f
C66 a_805_47# VGND 0.00579f
C67 RESET_B a_193_47# 0.0269f
C68 a_639_47# VGND 0.00863f
C69 RESET_B VPWR 0.0652f
C70 D VGND 0.0516f
C71 a_448_47# RESET_B 2.45e-19
C72 a_1270_413# RESET_B 2.06e-19
C73 a_27_47# RESET_B 0.296f
C74 a_651_413# RESET_B 0.0122f
C75 VPWR a_193_47# 0.396f
C76 a_448_47# a_193_47# 0.0642f
C77 VPB a_1283_21# 0.137f
C78 a_1270_413# a_193_47# 1.46e-19
C79 RESET_B VGND 0.288f
C80 a_448_47# VPWR 0.0681f
C81 RESET_B a_1108_47# 0.237f
C82 a_27_47# a_193_47# 0.906f
C83 a_651_413# a_193_47# 0.0346f
C84 a_1270_413# VPWR 7.19e-19
C85 a_27_47# a_448_47# 0.0931f
C86 a_27_47# VPWR 0.152f
C87 a_651_413# VPWR 0.129f
C88 VGND a_193_47# 0.0631f
C89 a_193_47# a_1108_47# 0.125f
C90 a_27_47# a_651_413# 9.73e-19
C91 a_448_47# VGND 0.0661f
C92 VPWR VGND 0.0502f
C93 RESET_B Q 9.12e-19
C94 VPWR a_1108_47# 0.173f
C95 a_1270_413# a_1108_47# 0.00645f
C96 a_27_47# VGND 0.254f
C97 a_27_47# a_1108_47# 0.102f
C98 Q a_193_47# 1.81e-19
C99 VPWR Q 0.0997f
C100 VGND a_1108_47# 0.148f
C101 a_1462_47# RESET_B 0.00288f
C102 VPB a_543_47# 0.0958f
C103 a_27_47# Q 2.63e-20
C104 Q VNB 0.0899f
C105 VGND VNB 1.02f
C106 VPWR VNB 0.831f
C107 RESET_B VNB 0.264f
C108 D VNB 0.16f
C109 CLK VNB 0.195f
C110 VPB VNB 1.85f
C111 a_651_413# VNB 0.00469f
C112 a_448_47# VNB 0.0139f
C113 a_1108_47# VNB 0.139f
C114 a_1283_21# VNB 0.299f
C115 a_543_47# VNB 0.158f
C116 a_761_289# VNB 0.121f
C117 a_193_47# VNB 0.274f
C118 a_27_47# VNB 0.496f
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
C0 VPB VGND 0.22f
C1 VPB VPWR 0.105f
C2 VGND VPWR 1.27f
C3 VPWR VNB 1.14f
C4 VGND VNB 0.992f
C5 VPB VNB 0.782f
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
C0 VPWR X 0.317f
C1 VGND a_27_47# 0.148f
C2 a_27_47# VPB 0.139f
C3 a_27_47# A 0.195f
C4 a_27_47# VPWR 0.219f
C5 VGND VPB 0.00583f
C6 a_27_47# X 0.328f
C7 VGND A 0.0431f
C8 VPB A 0.0321f
C9 VGND VPWR 0.057f
C10 VPB VPWR 0.0632f
C11 VGND X 0.216f
C12 VPB X 0.0122f
C13 A VPWR 0.022f
C14 A X 0.014f
C15 VGND VNB 0.358f
C16 X VNB 0.067f
C17 VPWR VNB 0.308f
C18 A VNB 0.148f
C19 VPB VNB 0.605f
C20 a_27_47# VNB 0.543f
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPWR VGND 0.0518f
C1 VPB A 0.0697f
C2 VPB a_27_47# 0.075f
C3 VPB X 0.00443f
C4 A VGND 0.0199f
C5 VGND a_27_47# 0.127f
C6 VGND X 0.111f
C7 VPB VGND 0.00642f
C8 A VPWR 0.0221f
C9 VPWR a_27_47# 0.153f
C10 VPWR X 0.169f
C11 VPB VPWR 0.0528f
C12 A a_27_47# 0.158f
C13 A X 0.00306f
C14 X a_27_47# 0.149f
C15 VGND VNB 0.284f
C16 X VNB 0.0215f
C17 VPWR VNB 0.25f
C18 A VNB 0.187f
C19 VPB VNB 0.428f
C20 a_27_47# VNB 0.284f
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_384_47# a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
C0 X VGND 0.0512f
C1 A1 a_81_21# 0.0568f
C2 VPWR a_81_21# 0.146f
C3 A1 A2 0.0921f
C4 VPWR A2 0.0201f
C5 A1 a_384_47# 0.00884f
C6 VPWR a_384_47# 4.08e-19
C7 a_81_21# B1 0.148f
C8 A1 VPB 0.0264f
C9 VPWR VPB 0.068f
C10 a_299_297# VGND 0.00772f
C11 B1 VPB 0.0387f
C12 VPWR A1 0.0209f
C13 a_81_21# X 0.112f
C14 A1 B1 0.0817f
C15 VPWR B1 0.0196f
C16 X VPB 0.0108f
C17 a_81_21# VGND 0.173f
C18 A2 VGND 0.0495f
C19 a_384_47# VGND 0.00366f
C20 a_81_21# a_299_297# 0.0821f
C21 VPWR X 0.0847f
C22 VPB VGND 0.00713f
C23 a_299_297# A2 0.0468f
C24 a_299_297# a_384_47# 1.48e-19
C25 X B1 3.04e-20
C26 a_299_297# VPB 0.0111f
C27 A1 VGND 0.0786f
C28 VPWR VGND 0.0579f
C29 A1 a_299_297# 0.0585f
C30 VPWR a_299_297# 0.202f
C31 B1 VGND 0.0181f
C32 a_81_21# A2 7.47e-19
C33 a_81_21# a_384_47# 0.00138f
C34 a_299_297# B1 0.00863f
C35 a_81_21# VPB 0.0593f
C36 VPB A2 0.0373f
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
C0 VPB VGND 0.116f
C1 VPWR VGND 0.546f
C2 VPB VPWR 0.0787f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
C0 VPB A 0.0806f
C1 VPWR VGND 0.0461f
C2 VGND a_145_75# 0.00468f
C3 VPWR a_59_75# 0.15f
C4 VGND B 0.0115f
C5 a_145_75# a_59_75# 0.00658f
C6 VGND X 0.0993f
C7 VGND VPB 0.008f
C8 a_59_75# B 0.143f
C9 X a_59_75# 0.109f
C10 VPWR a_145_75# 6.31e-19
C11 VPB a_59_75# 0.0563f
C12 VGND A 0.0147f
C13 VPWR B 0.0117f
C14 VPWR X 0.111f
C15 VPWR VPB 0.0729f
C16 a_59_75# A 0.0809f
C17 X a_145_75# 5.76e-19
C18 X B 0.00276f
C19 VPWR A 0.0362f
C20 VPB B 0.0629f
C21 VPB X 0.0127f
C22 VGND a_59_75# 0.116f
C23 B A 0.0971f
C24 X A 1.68e-19
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X a_27_297# a_109_47#
+ a_109_297# a_373_47#
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VGND a_109_297# 0.00426f
C1 B2 a_109_297# 0.0015f
C2 A2 VPWR 0.0178f
C3 a_27_297# VPWR 0.13f
C4 A2 VPB 0.0284f
C5 A2 X 0.0011f
C6 a_27_297# VPB 0.0591f
C7 a_27_297# X 0.108f
C8 A2 B1 1.81e-19
C9 a_27_297# B1 0.0838f
C10 A1 VPWR 0.0168f
C11 A1 VPB 0.0387f
C12 A1 X 2.98e-19
C13 A1 B1 0.0657f
C14 a_109_47# VPWR 0.00104f
C15 a_27_297# A2 0.161f
C16 a_373_47# VPWR 7.36e-19
C17 a_373_47# X 1.97e-19
C18 B1 a_109_47# 0.00145f
C19 VGND VPWR 0.0641f
C20 B2 VPWR 0.0126f
C21 VGND VPB 0.00746f
C22 VGND X 0.0543f
C23 B2 VPB 0.0299f
C24 B2 X 3.26e-20
C25 A2 A1 0.0738f
C26 a_27_297# A1 0.0839f
C27 VGND B1 0.0267f
C28 B2 B1 0.0739f
C29 a_27_297# a_109_47# 0.00393f
C30 A2 a_373_47# 6.81e-19
C31 VPWR a_109_297# 0.187f
C32 a_27_297# a_373_47# 0.0134f
C33 VPB a_109_297# 0.00882f
C34 X a_109_297# 0.00169f
C35 VGND A2 0.0162f
C36 A2 B2 8.94e-20
C37 VGND a_27_297# 0.257f
C38 a_27_297# B2 0.0567f
C39 B1 a_109_297# 0.0106f
C40 a_373_47# A1 0.00122f
C41 VGND A1 0.0137f
C42 A2 a_109_297# 0.00625f
C43 a_27_297# a_109_297# 0.171f
C44 VGND a_109_47# 0.00792f
C45 B2 a_109_47# 4.58e-19
C46 VGND a_373_47# 0.00344f
C47 A1 a_109_297# 0.0105f
C48 VGND B2 0.0538f
C49 VPB VPWR 0.0714f
C50 X VPWR 0.0914f
C51 X VPB 0.011f
C52 B1 VPWR 0.0139f
C53 B1 VPB 0.0317f
C54 B1 X 8.38e-20
C55 VGND VNB 0.421f
C56 X VNB 0.0917f
C57 VPWR VNB 0.328f
C58 A2 VNB 0.0927f
C59 A1 VNB 0.112f
C60 B1 VNB 0.112f
C61 B2 VNB 0.126f
C62 VPB VNB 0.693f
C63 a_109_297# VNB 0.00274f
C64 a_27_297# VNB 0.19f
.ends

.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X a_78_199# a_493_297#
+ a_215_47# a_292_297#
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPB VGND 0.00596f
C1 a_78_199# VGND 0.0684f
C2 VPWR A1 0.057f
C3 VPWR B2 0.0104f
C4 a_215_47# X 0.00228f
C5 VPB VPWR 0.0744f
C6 VPWR a_78_199# 0.211f
C7 a_215_47# B1 0.00758f
C8 A2 B1 3.91e-19
C9 A2 a_292_297# 4.41e-20
C10 VPWR VGND 0.0668f
C11 X B2 1.65e-19
C12 A2 a_215_47# 0.0439f
C13 VPB X 0.0107f
C14 X a_78_199# 0.105f
C15 B2 B1 0.0815f
C16 VPB B1 0.0388f
C17 B2 a_292_297# 4.98e-20
C18 a_78_199# B1 0.148f
C19 a_215_47# a_493_297# 3.25e-19
C20 A2 a_493_297# 0.0105f
C21 a_78_199# a_292_297# 0.013f
C22 a_215_47# A1 0.0498f
C23 X VGND 0.0472f
C24 A2 A1 0.0879f
C25 a_215_47# B2 0.0207f
C26 A2 B2 0.0676f
C27 B1 VGND 0.0119f
C28 VPB a_215_47# 9.85e-19
C29 a_215_47# a_78_199# 0.0907f
C30 VPB A2 0.0341f
C31 X VPWR 0.0911f
C32 A2 a_78_199# 0.0707f
C33 a_493_297# A1 9.88e-20
C34 a_292_297# VGND 0.00136f
C35 VPWR B1 0.0227f
C36 a_78_199# a_493_297# 3.15e-19
C37 VPWR a_292_297# 0.00854f
C38 a_215_47# VGND 0.258f
C39 A2 VGND 0.0153f
C40 VPB A1 0.0319f
C41 a_78_199# A1 4.58e-19
C42 VPB B2 0.0281f
C43 a_78_199# B2 0.0816f
C44 a_215_47# VPWR 0.00435f
C45 A2 VPWR 0.12f
C46 a_493_297# VGND 3.15e-19
C47 VPB a_78_199# 0.0517f
C48 X B1 6.11e-19
C49 X a_292_297# 4.46e-19
C50 VPWR a_493_297# 0.00283f
C51 A1 VGND 0.0146f
C52 B2 VGND 0.0103f
C53 VGND VNB 0.403f
C54 VPWR VNB 0.359f
C55 X VNB 0.0884f
C56 A1 VNB 0.132f
C57 A2 VNB 0.0971f
C58 B2 VNB 0.0913f
C59 B1 VNB 0.11f
C60 VPB VNB 0.693f
C61 a_215_47# VNB 0.0357f
C62 a_78_199# VNB 0.154f
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
C0 VPB VPWR 0.0858f
C1 VPWR VGND 0.903f
C2 VPB VGND 0.161f
C3 VPWR VNB 0.867f
C4 VGND VNB 0.761f
C5 VPB VNB 0.605f
.ends

.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y a_408_47# a_218_47#
+ a_27_47#
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176 pd=1.39 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.12 ps=1.04 w=0.65 l=0.15
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.176 ps=1.39 w=1 l=0.15
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.04 as=0.109 ps=1.36 w=0.42 l=0.15
C0 C A_N 0.0603f
C1 VPB a_218_47# 1.44e-19
C2 C VPB 0.0536f
C3 VPB B 0.082f
C4 VGND a_27_47# 0.119f
C5 a_408_47# a_27_47# 0.0212f
C6 VGND VPWR 0.0834f
C7 a_408_47# VPWR 0.00288f
C8 Y a_27_47# 0.35f
C9 VPB A_N 0.0913f
C10 Y VPWR 0.457f
C11 a_408_47# VGND 0.243f
C12 a_218_47# a_27_47# 0.00788f
C13 C a_27_47# 0.0792f
C14 a_218_47# VPWR 0.00305f
C15 B a_27_47# 0.176f
C16 VGND Y 0.0176f
C17 a_408_47# Y 0.0985f
C18 C VPWR 0.032f
C19 B VPWR 0.0305f
C20 VGND a_218_47# 0.173f
C21 a_408_47# a_218_47# 0.097f
C22 a_27_47# A_N 0.0854f
C23 C VGND 0.0348f
C24 VGND B 0.0223f
C25 C a_408_47# 7.76e-20
C26 a_408_47# B 0.0409f
C27 VPWR A_N 0.023f
C28 VPB a_27_47# 0.098f
C29 C Y 0.0232f
C30 B Y 0.031f
C31 VPB VPWR 0.0961f
C32 VGND A_N 0.0459f
C33 a_408_47# A_N 5.25e-20
C34 C a_218_47# 0.0806f
C35 B a_218_47# 0.0867f
C36 VGND VPB 0.00877f
C37 Y A_N 0.00302f
C38 C B 0.0583f
C39 VPB Y 0.0201f
C40 a_218_47# A_N 0.00187f
C41 VPWR a_27_47# 0.174f
C42 VGND VNB 0.483f
C43 Y VNB 0.0685f
C44 VPWR VNB 0.41f
C45 B VNB 0.227f
C46 C VNB 0.176f
C47 A_N VNB 0.171f
C48 VPB VNB 0.871f
C49 a_408_47# VNB 0.0232f
C50 a_218_47# VNB 0.0113f
C51 a_27_47# VNB 0.296f
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q a_1462_47# a_543_47#
+ a_651_413# a_193_47# a_805_47# a_448_47# a_639_47# a_1283_21# a_761_289# a_1108_47#
+ a_1217_47# a_1270_413# a_27_47#
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
C0 a_1108_47# VGND 0.148f
C1 RESET_B Q 8.96e-19
C2 VPWR VGND 0.0719f
C3 a_27_47# a_651_413# 9.73e-19
C4 a_27_47# VPB 0.262f
C5 a_193_47# a_651_413# 0.0346f
C6 a_1283_21# RESET_B 0.279f
C7 a_193_47# VPB 0.171f
C8 a_639_47# VGND 0.00863f
C9 a_448_47# VGND 0.0661f
C10 a_543_47# D 7.35e-20
C11 a_805_47# RESET_B 0.00316f
C12 a_761_289# VGND 0.0734f
C13 a_1283_21# a_1462_47# 0.0074f
C14 a_1108_47# Q 9.64e-19
C15 VPWR Q 0.169f
C16 a_27_47# CLK 0.234f
C17 a_1283_21# a_1108_47# 0.234f
C18 a_193_47# CLK 7.94e-19
C19 a_1283_21# VPWR 0.23f
C20 a_543_47# RESET_B 0.153f
C21 a_651_413# VPB 0.0135f
C22 a_805_47# a_761_289# 3.69e-19
C23 VGND Q 0.11f
C24 a_27_47# D 0.133f
C25 a_1283_21# VGND 0.259f
C26 a_193_47# D 0.218f
C27 a_543_47# a_1108_47# 7.99e-20
C28 a_543_47# VPWR 0.1f
C29 a_1217_47# RESET_B 6.03e-19
C30 a_805_47# VGND 0.00579f
C31 a_543_47# a_639_47# 0.0138f
C32 a_543_47# a_448_47# 0.0498f
C33 a_1270_413# RESET_B 2.06e-19
C34 a_543_47# a_761_289# 0.21f
C35 VPB CLK 0.0693f
C36 a_27_47# RESET_B 0.296f
C37 a_193_47# RESET_B 0.0269f
C38 a_1283_21# Q 0.0963f
C39 a_1217_47# a_1108_47# 0.00742f
C40 a_543_47# VGND 0.123f
C41 a_1270_413# a_1108_47# 0.00645f
C42 a_1270_413# VPWR 7.19e-19
C43 a_761_289# a_1217_47# 4.2e-19
C44 VPB D 0.138f
C45 a_27_47# a_1108_47# 0.102f
C46 a_27_47# VPWR 0.152f
C47 a_193_47# a_1108_47# 0.125f
C48 a_193_47# VPWR 0.396f
C49 a_27_47# a_639_47# 0.00188f
C50 a_1217_47# VGND 9.68e-19
C51 a_1270_413# a_761_289# 2.6e-19
C52 a_193_47# a_639_47# 2.28e-19
C53 a_27_47# a_448_47# 0.0931f
C54 a_193_47# a_448_47# 0.0642f
C55 a_805_47# a_543_47# 0.00171f
C56 a_27_47# a_761_289# 0.0701f
C57 a_193_47# a_761_289# 0.186f
C58 a_651_413# RESET_B 0.0122f
C59 VPB RESET_B 0.138f
C60 a_27_47# VGND 0.254f
C61 a_193_47# VGND 0.0631f
C62 a_651_413# VPWR 0.129f
C63 a_1108_47# VPB 0.115f
C64 VPB VPWR 0.234f
C65 CLK RESET_B 1.09e-19
C66 a_27_47# Q 2.57e-20
C67 a_193_47# Q 1.79e-19
C68 a_448_47# VPB 0.0141f
C69 a_27_47# a_1283_21# 0.0436f
C70 a_1283_21# a_193_47# 0.0425f
C71 a_761_289# a_651_413# 0.0977f
C72 a_761_289# VPB 0.0994f
C73 D RESET_B 4.72e-19
C74 VPB VGND 0.0122f
C75 CLK VPWR 0.0174f
C76 a_27_47# a_543_47# 0.115f
C77 a_193_47# a_543_47# 0.23f
C78 VPB Q 0.00555f
C79 CLK VGND 0.0172f
C80 D VPWR 0.0812f
C81 a_1283_21# VPB 0.168f
C82 a_448_47# D 0.156f
C83 a_27_47# a_1217_47# 2.56e-19
C84 a_193_47# a_1217_47# 2.36e-20
C85 a_1462_47# RESET_B 0.00288f
C86 a_193_47# a_1270_413# 1.46e-19
C87 a_1108_47# RESET_B 0.237f
C88 RESET_B VPWR 0.0652f
C89 D VGND 0.0516f
C90 a_639_47# RESET_B 9.54e-19
C91 a_543_47# a_651_413# 0.0572f
C92 a_448_47# RESET_B 2.45e-19
C93 a_543_47# VPB 0.0958f
C94 a_27_47# a_193_47# 0.906f
C95 a_761_289# RESET_B 0.166f
C96 a_1108_47# VPWR 0.174f
C97 RESET_B VGND 0.288f
C98 a_448_47# VPWR 0.0681f
C99 a_448_47# a_639_47# 4.61e-19
C100 a_1462_47# VGND 0.00221f
C101 a_761_289# a_1108_47# 0.0512f
C102 a_761_289# VPWR 0.105f
C103 a_761_289# a_639_47# 3.16e-19
C104 Q VNB 0.0296f
C105 VGND VNB 1.1f
C106 VPWR VNB 0.902f
C107 RESET_B VNB 0.263f
C108 D VNB 0.16f
C109 CLK VNB 0.195f
C110 VPB VNB 1.93f
C111 a_651_413# VNB 0.00469f
C112 a_448_47# VNB 0.0139f
C113 a_1108_47# VNB 0.137f
C114 a_1283_21# VNB 0.389f
C115 a_543_47# VNB 0.158f
C116 a_761_289# VNB 0.121f
C117 a_193_47# VNB 0.273f
C118 a_27_47# VNB 0.496f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VGND a_285_47# 0.00552f
C1 X VPB 0.0154f
C2 A VPB 0.051f
C3 VGND X 0.173f
C4 VGND A 0.0325f
C5 VPWR a_35_297# 0.096f
C6 VPWR a_117_297# 0.00852f
C7 a_35_297# a_117_297# 0.00641f
C8 VGND VPB 0.00696f
C9 VPWR a_285_297# 0.246f
C10 a_35_297# a_285_297# 0.025f
C11 VPWR B 0.0703f
C12 B a_35_297# 0.203f
C13 VPWR a_285_47# 8.6e-19
C14 a_35_297# a_285_47# 0.00723f
C15 B a_117_297# 0.00777f
C16 X VPWR 0.0537f
C17 X a_35_297# 0.166f
C18 A VPWR 0.0348f
C19 A a_35_297# 0.0633f
C20 B a_285_297# 0.0553f
C21 X a_117_297# 2.25e-19
C22 B a_285_47# 3.98e-19
C23 VPWR VPB 0.0689f
C24 a_35_297# VPB 0.0699f
C25 X a_285_297# 0.0712f
C26 VGND VPWR 0.0643f
C27 A a_285_297# 0.00749f
C28 VGND a_35_297# 0.177f
C29 X B 0.0149f
C30 A B 0.221f
C31 X a_285_47# 0.00206f
C32 VGND a_117_297# 0.00177f
C33 a_285_297# VPB 0.0133f
C34 VGND a_285_297# 0.00394f
C35 A X 0.00166f
C36 B VPB 0.0697f
C37 VGND B 0.0304f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
C0 X A 8.48e-19
C1 VPB VPWR 0.0355f
C2 VPB VGND 0.00505f
C3 VPB a_27_47# 0.0592f
C4 VPWR A 0.0215f
C5 A VGND 0.0184f
C6 a_27_47# A 0.181f
C7 VPB A 0.0524f
C8 VPWR X 0.0897f
C9 X VGND 0.0546f
C10 X a_27_47# 0.107f
C11 VPB X 0.0128f
C12 VPWR VGND 0.029f
C13 VPWR a_27_47# 0.135f
C14 a_27_47# VGND 0.105f
C15 VGND VNB 0.207f
C16 X VNB 0.0941f
C17 VPWR VNB 0.175f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_27_47# VNB 0.208f
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X a_27_413# a_297_47# a_207_413#
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_297_47# X 8.17e-20
C1 VPB a_207_413# 0.0478f
C2 A_N VGND 0.0473f
C3 A_N VPWR 0.0182f
C4 VPB B 0.111f
C5 VPB VGND 0.00763f
C6 VPB VPWR 0.0634f
C7 a_297_47# a_207_413# 0.00476f
C8 a_27_413# a_207_413# 0.185f
C9 a_297_47# VGND 0.00504f
C10 a_297_47# VPWR 6.35e-19
C11 A_N VPB 0.0801f
C12 X a_207_413# 0.0716f
C13 a_27_413# B 0.0926f
C14 VGND a_27_413# 0.0863f
C15 VPWR a_27_413# 0.108f
C16 B X 0.0303f
C17 VGND X 0.0652f
C18 VPWR X 0.0552f
C19 A_N a_27_413# 0.198f
C20 VPB a_27_413# 0.0834f
C21 B a_207_413# 0.182f
C22 VGND a_207_413# 0.115f
C23 VPWR a_207_413# 0.111f
C24 VPB X 0.0122f
C25 VGND B 0.0187f
C26 VPWR B 0.0867f
C27 VPWR VGND 0.0564f
C28 A_N a_207_413# 8.2e-19
C29 VGND VNB 0.368f
C30 X VNB 0.0892f
C31 VPWR VNB 0.292f
C32 B VNB 0.132f
C33 A_N VNB 0.201f
C34 VPB VNB 0.605f
C35 a_207_413# VNB 0.137f
C36 a_27_413# VNB 0.197f
.ends

.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X a_212_413# a_27_413# a_297_47#
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.229 ps=1.75 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.75 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VGND a_212_413# 0.137f
C1 VPWR a_212_413# 0.132f
C2 VGND A_N 0.0469f
C3 A_N VPWR 0.0181f
C4 VGND X 0.103f
C5 A_N a_212_413# 7.63e-19
C6 VPWR X 0.112f
C7 VGND VPB 0.00913f
C8 VGND B 0.0188f
C9 VPB VPWR 0.0784f
C10 VGND a_297_47# 0.00553f
C11 VGND a_27_413# 0.0862f
C12 a_212_413# X 0.109f
C13 VPWR B 0.0871f
C14 a_297_47# VPWR 6.75e-19
C15 a_27_413# VPWR 0.109f
C16 VPB a_212_413# 0.0794f
C17 B a_212_413# 0.182f
C18 a_297_47# a_212_413# 0.00539f
C19 a_27_413# a_212_413# 0.183f
C20 VPB A_N 0.0808f
C21 A_N a_27_413# 0.194f
C22 VPB X 0.00781f
C23 B X 0.0303f
C24 a_297_47# X 8.32e-20
C25 VPB B 0.113f
C26 VGND VPWR 0.0772f
C27 VPB a_27_413# 0.0853f
C28 a_27_413# B 0.0875f
C29 VGND VNB 0.437f
C30 X VNB 0.0366f
C31 VPWR VNB 0.358f
C32 B VNB 0.133f
C33 A_N VNB 0.202f
C34 VPB VNB 0.693f
C35 a_212_413# VNB 0.228f
C36 a_27_413# VNB 0.196f
.ends

.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y a_277_297# a_27_297#
+ a_694_21# a_474_297#
X0 VPWR D_N a_694_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_27_297# B a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_474_297# a_694_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_277_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y a_694_21# a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND D_N a_694_21# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_474_297# C a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 Y a_694_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_277_297# C a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND a_694_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_277_297# C 0.0172f
C1 a_474_297# C 0.0918f
C2 a_694_21# C 0.0591f
C3 VPB VGND 0.0139f
C4 VPWR VGND 0.107f
C5 VPB A 0.0568f
C6 VPWR A 0.0387f
C7 VPB D_N 0.115f
C8 VPB B 0.0615f
C9 VPWR D_N 0.04f
C10 VPWR B 0.0233f
C11 Y a_27_297# 0.00665f
C12 a_277_297# a_27_297# 0.145f
C13 a_474_297# a_27_297# 0.0551f
C14 VGND Y 0.597f
C15 Y A 0.0854f
C16 Y D_N 0.00144f
C17 VPWR VPB 0.12f
C18 B Y 0.135f
C19 a_277_297# VGND 0.00337f
C20 VGND a_474_297# 0.0139f
C21 VGND a_694_21# 0.154f
C22 a_277_297# D_N 1.67e-19
C23 a_474_297# D_N 0.00185f
C24 a_277_297# B 0.021f
C25 a_474_297# B 0.0297f
C26 C a_27_297# 1.05e-19
C27 D_N a_694_21# 0.0977f
C28 VPB Y 0.00707f
C29 VGND C 0.0304f
C30 VPWR Y 0.0138f
C31 B C 0.0392f
C32 a_277_297# VPB 0.0101f
C33 VPB a_474_297# 0.0135f
C34 a_277_297# VPWR 0.183f
C35 VPWR a_474_297# 0.142f
C36 VPB a_694_21# 0.107f
C37 VPWR a_694_21# 0.0917f
C38 VPB C 0.0577f
C39 VGND a_27_297# 0.00756f
C40 VPWR C 0.021f
C41 a_474_297# Y 0.126f
C42 A a_27_297# 0.132f
C43 D_N a_27_297# 4.51e-19
C44 B a_27_297# 0.0932f
C45 Y a_694_21# 0.122f
C46 a_277_297# a_474_297# 0.149f
C47 VGND A 0.0583f
C48 VGND D_N 0.0436f
C49 VGND B 0.0316f
C50 a_474_297# a_694_21# 0.0922f
C51 Y C 0.113f
C52 B A 0.0717f
C53 VPB a_27_297# 0.0177f
C54 VPWR a_27_297# 0.237f
C55 VGND VNB 0.698f
C56 Y VNB 0.0244f
C57 VPWR VNB 0.536f
C58 D_N VNB 0.176f
C59 C VNB 0.181f
C60 B VNB 0.187f
C61 A VNB 0.21f
C62 VPB VNB 1.14f
C63 a_474_297# VNB 7.04e-19
C64 a_277_297# VNB 0.0042f
C65 a_27_297# VNB 0.0363f
C66 a_694_21# VNB 0.257f
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y a_109_297#
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 Y B 0.0877f
C1 VPB A 0.0415f
C2 VPB VPWR 0.0449f
C3 Y VGND 0.154f
C4 A B 0.0584f
C5 B VPWR 0.0148f
C6 A VGND 0.0486f
C7 VGND VPWR 0.0314f
C8 a_109_297# VGND 0.00128f
C9 VPB B 0.0367f
C10 A Y 0.0471f
C11 Y VPWR 0.0995f
C12 VPB VGND 0.00456f
C13 Y a_109_297# 0.0113f
C14 B VGND 0.0451f
C15 VPB Y 0.0139f
C16 A VPWR 0.0528f
C17 a_109_297# VPWR 0.00638f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y a_27_47#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPWR Y 0.398f
C1 VPWR VGND 0.0476f
C2 VPWR B 0.06f
C3 A Y 0.178f
C4 A VGND 0.018f
C5 A B 0.0748f
C6 VPB Y 0.0159f
C7 VPWR A 0.0315f
C8 VPB VGND 0.00576f
C9 a_27_47# Y 0.0956f
C10 VPB B 0.0568f
C11 VGND a_27_47# 0.259f
C12 B a_27_47# 0.0896f
C13 VPWR VPB 0.0664f
C14 VPWR a_27_47# 0.00338f
C15 VPB A 0.0571f
C16 A a_27_47# 0.0374f
C17 VPB a_27_47# 1.51e-19
C18 VGND Y 0.0208f
C19 B Y 0.062f
C20 B VGND 0.029f
C21 VGND VNB 0.296f
C22 Y VNB 0.063f
C23 VPWR VNB 0.309f
C24 A VNB 0.198f
C25 B VNB 0.209f
C26 VPB VNB 0.516f
C27 a_27_47# VNB 0.0484f
.ends

.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X a_373_53# a_215_311#
+ a_301_53# a_109_53#
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.1 w=0.65 l=0.15
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.1 as=0.0536 ps=0.675 w=0.42 l=0.15
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPWR a_109_53# 0.0609f
C1 C VPB 0.0346f
C2 VPB X 0.00646f
C3 VPB VPWR 0.144f
C4 a_373_53# a_215_311# 0.0026f
C5 a_373_53# VGND 0.00282f
C6 VPB a_109_53# 0.0621f
C7 VPWR A_N 0.0362f
C8 C B 0.0684f
C9 X B 8.71e-19
C10 C a_215_311# 0.19f
C11 X a_215_311# 0.125f
C12 a_109_53# A_N 0.0949f
C13 VPWR B 0.132f
C14 C VGND 0.0706f
C15 a_301_53# VPWR 1.15e-19
C16 X VGND 0.139f
C17 a_215_311# VPWR 0.179f
C18 VGND VPWR 0.0802f
C19 VPB A_N 0.0535f
C20 B a_109_53# 0.0797f
C21 a_301_53# a_109_53# 1.81e-19
C22 a_215_311# a_109_53# 0.179f
C23 C a_373_53# 0.00415f
C24 VGND a_109_53# 0.0717f
C25 VPB B 0.0926f
C26 a_373_53# VPWR 4.26e-19
C27 VPB a_215_311# 0.0818f
C28 VPB VGND 0.0111f
C29 a_215_311# A_N 6.83e-19
C30 VGND A_N 0.044f
C31 C X 0.0161f
C32 C VPWR 0.00933f
C33 X VPWR 0.193f
C34 a_215_311# B 0.0583f
C35 a_215_311# a_301_53# 0.0049f
C36 VGND B 0.00805f
C37 VGND a_301_53# 5.98e-19
C38 VGND a_215_311# 0.144f
C39 VGND VNB 0.485f
C40 X VNB 0.0401f
C41 C VNB 0.114f
C42 A_N VNB 0.188f
C43 VPWR VNB 0.428f
C44 B VNB 0.0998f
C45 VPB VNB 0.782f
C46 a_109_53# VNB 0.154f
C47 a_215_311# VNB 0.233f
.ends

.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q a_1140_413# a_1296_47#
+ a_1182_261# a_586_47# a_1602_47# a_956_413# a_1224_47# a_193_47# a_796_47# a_381_47#
+ a_1056_47# a_1032_413# a_562_413# a_652_21# a_476_47# a_27_47#
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
C0 a_1602_47# SET_B 0.00213f
C1 a_652_21# a_956_413# 3.11e-19
C2 CLK VGND 0.0194f
C3 a_652_21# VPWR 0.144f
C4 a_27_47# VPB 0.226f
C5 a_476_47# VPWR 0.12f
C6 D a_381_47# 0.14f
C7 a_796_47# VGND 0.00583f
C8 a_27_47# a_956_413# 0.00294f
C9 a_27_47# VPWR 0.438f
C10 a_1032_413# a_193_47# 0.0573f
C11 a_652_21# a_1224_47# 1.57e-19
C12 a_1032_413# SET_B 0.215f
C13 a_652_21# VGND 0.0761f
C14 a_586_47# a_381_47# 3.7e-19
C15 a_476_47# VGND 0.178f
C16 a_1224_47# a_27_47# 1.63e-19
C17 CLK a_193_47# 0.00156f
C18 a_27_47# VGND 0.164f
C19 a_1602_47# a_1182_261# 0.144f
C20 a_1056_47# a_1032_413# 0.0016f
C21 VPB VPWR 0.218f
C22 a_796_47# SET_B 0.00149f
C23 VPWR a_956_413# 0.00457f
C24 a_1032_413# a_1140_413# 0.00523f
C25 a_1602_47# Q 0.0715f
C26 a_652_21# a_193_47# 0.0849f
C27 a_476_47# a_193_47# 0.215f
C28 VPB VGND 0.0173f
C29 a_652_21# SET_B 0.157f
C30 a_1032_413# a_1182_261# 0.344f
C31 a_476_47# SET_B 0.203f
C32 VGND a_956_413# 3.4e-19
C33 a_27_47# a_193_47# 0.797f
C34 VPWR VGND 0.0687f
C35 a_27_47# SET_B 0.0407f
C36 a_652_21# a_1056_47# 3.94e-19
C37 a_1032_413# Q 0.00365f
C38 a_652_21# a_381_47# 7.79e-20
C39 a_1224_47# VGND 0.00169f
C40 a_476_47# a_381_47# 0.0356f
C41 a_1056_47# a_27_47# 0.00248f
C42 VPB a_193_47# 0.179f
C43 a_652_21# a_562_413# 9.35e-20
C44 VGND a_1296_47# 0.00523f
C45 a_1602_47# a_1032_413# 0.111f
C46 a_476_47# a_562_413# 0.00972f
C47 VPB SET_B 0.143f
C48 a_27_47# a_381_47# 0.0729f
C49 VPWR a_193_47# 0.101f
C50 a_562_413# a_27_47# 0.0018f
C51 SET_B VPWR 0.0807f
C52 a_1182_261# a_27_47# 0.0608f
C53 a_476_47# D 1.36e-19
C54 VPB a_381_47# 0.0101f
C55 a_1224_47# SET_B 8.75e-19
C56 VGND a_193_47# 0.219f
C57 SET_B VGND 0.338f
C58 SET_B a_1296_47# 0.00167f
C59 a_27_47# D 0.103f
C60 Q a_27_47# 1.08e-19
C61 VPWR a_381_47# 0.0942f
C62 a_1182_261# VPB 0.112f
C63 a_1140_413# VPWR 0.00334f
C64 a_562_413# VPWR 0.0041f
C65 a_586_47# a_476_47# 0.00807f
C66 a_1056_47# VGND 0.00386f
C67 a_1602_47# a_27_47# 2.39e-19
C68 a_1182_261# VPWR 0.123f
C69 VGND a_381_47# 0.0787f
C70 VPB D 0.0485f
C71 Q VPB 0.0174f
C72 a_652_21# a_1032_413# 0.00971f
C73 SET_B a_193_47# 0.202f
C74 a_476_47# a_1032_413# 0.00329f
C75 D VPWR 0.0158f
C76 Q VPWR 0.0704f
C77 a_1182_261# VGND 0.0628f
C78 a_1182_261# a_1296_47# 1.84e-19
C79 a_1602_47# VPB 0.0453f
C80 a_1032_413# a_27_47# 0.183f
C81 a_1602_47# VPWR 0.135f
C82 a_1056_47# SET_B 0.00152f
C83 a_652_21# a_796_47# 0.00196f
C84 a_476_47# a_796_47# 0.00184f
C85 a_381_47# a_193_47# 0.157f
C86 D VGND 0.014f
C87 Q VGND 0.0595f
C88 a_27_47# CLK 0.214f
C89 a_562_413# a_193_47# 4.45e-20
C90 a_1140_413# SET_B 6.31e-19
C91 a_1032_413# VPB 0.177f
C92 a_1032_413# a_956_413# 0.00212f
C93 a_1182_261# a_193_47# 0.0728f
C94 a_652_21# a_476_47# 0.26f
C95 a_1602_47# VGND 0.0942f
C96 a_1032_413# VPWR 0.257f
C97 a_1182_261# SET_B 0.12f
C98 a_586_47# VGND 0.00172f
C99 a_652_21# a_27_47# 0.19f
C100 VPB CLK 0.0702f
C101 a_476_47# a_27_47# 0.223f
C102 D a_193_47# 0.0606f
C103 Q a_193_47# 6.4e-20
C104 a_1224_47# a_1032_413# 0.00536f
C105 a_562_413# a_381_47# 8.75e-19
C106 CLK VPWR 0.0194f
C107 Q SET_B 4.58e-19
C108 a_1032_413# VGND 0.157f
C109 a_1032_413# a_1296_47# 0.00384f
C110 a_1602_47# a_193_47# 4.3e-19
C111 a_652_21# VPB 0.0992f
C112 a_476_47# VPB 0.146f
C113 a_586_47# a_193_47# 0.00206f
C114 Q VNB 0.0834f
C115 VGND VNB 1.08f
C116 VPWR VNB 0.875f
C117 SET_B VNB 0.247f
C118 D VNB 0.107f
C119 CLK VNB 0.196f
C120 VPB VNB 1.93f
C121 a_381_47# VNB 0.0203f
C122 a_1602_47# VNB 0.126f
C123 a_1032_413# VNB 0.305f
C124 a_1182_261# VNB 0.128f
C125 a_476_47# VNB 0.286f
C126 a_652_21# VNB 0.119f
C127 a_193_47# VNB 0.322f
C128 a_27_47# VNB 0.437f
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X a_505_21# a_535_374# a_439_47#
+ a_218_47# a_76_199# a_218_374#
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPWR a_218_47# 4.95e-19
C1 A1 S 0.0872f
C2 a_218_374# VGND 7.29e-19
C3 S VGND 0.033f
C4 VPWR A0 0.00732f
C5 a_76_199# a_218_374# 0.00557f
C6 VPWR X 0.128f
C7 S a_76_199# 0.318f
C8 a_505_21# VPB 0.0781f
C9 A1 a_505_21# 0.0993f
C10 VPWR a_535_374# 8.63e-19
C11 A0 S 0.0341f
C12 A1 VPB 0.0721f
C13 a_505_21# VGND 0.124f
C14 A1 a_439_47# 0.00498f
C15 VPB VGND 0.0134f
C16 a_439_47# VGND 0.00354f
C17 S X 0.00823f
C18 A1 VGND 0.0752f
C19 a_76_199# VPB 0.0481f
C20 S a_535_374# 0.00526f
C21 A1 a_76_199# 0.187f
C22 A0 a_505_21# 0.0383f
C23 VPWR a_218_374# 0.00177f
C24 A0 VPB 0.107f
C25 a_76_199# VGND 0.16f
C26 VPWR S 0.392f
C27 A0 a_439_47# 0.00369f
C28 a_218_47# VGND 0.00328f
C29 X VPB 0.012f
C30 A0 A1 0.267f
C31 A0 VGND 0.0432f
C32 a_76_199# a_218_47# 0.00783f
C33 S a_218_374# 0.00688f
C34 X VGND 0.0586f
C35 A0 a_76_199# 0.0544f
C36 VPWR a_505_21# 0.0818f
C37 VPWR VPB 0.11f
C38 VPWR a_439_47# 4.69e-19
C39 X a_76_199# 0.0776f
C40 a_535_374# VGND 6.38e-19
C41 X a_218_47# 2.88e-19
C42 VPWR A1 0.0114f
C43 VPWR VGND 0.0804f
C44 a_76_199# a_535_374# 6.64e-19
C45 S a_505_21# 0.198f
C46 S VPB 0.168f
C47 VPWR a_76_199# 0.0542f
C48 VGND VNB 0.499f
C49 A1 VNB 0.14f
C50 A0 VNB 0.134f
C51 S VNB 0.268f
C52 VPWR VNB 0.419f
C53 X VNB 0.0924f
C54 VPB VNB 0.871f
C55 a_505_21# VNB 0.247f
C56 a_76_199# VNB 0.139f
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 Y A 0.0894f
C1 A VGND 0.0638f
C2 VPB VPWR 0.0521f
C3 VPWR A 0.0631f
C4 Y VGND 0.155f
C5 VPB A 0.0742f
C6 VPWR Y 0.209f
C7 VPWR VGND 0.0423f
C8 VPB Y 0.0061f
C9 VPB VGND 0.00649f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X a_161_47#
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
C0 VPWR VPB 0.102f
C1 VPB X 0.013f
C2 A VPB 0.0756f
C3 VPWR a_161_47# 0.338f
C4 a_161_47# X 0.301f
C5 VGND VPB 0.01f
C6 VPWR X 0.508f
C7 A a_161_47# 0.202f
C8 VGND a_161_47# 0.234f
C9 A VPWR 0.0505f
C10 A X 3.93e-19
C11 VPWR VGND 0.102f
C12 VGND X 0.364f
C13 A VGND 0.0417f
C14 VPB a_161_47# 0.187f
C15 VGND VNB 0.533f
C16 X VNB 0.0506f
C17 VPWR VNB 0.48f
C18 A VNB 0.24f
C19 VPB VNB 0.871f
C20 a_161_47# VNB 0.593f
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X a_110_47#
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
C0 A a_110_47# 0.307f
C1 VPWR X 1.36f
C2 VPWR VPB 0.184f
C3 A X 0.00292f
C4 A VPB 0.133f
C5 VGND a_110_47# 0.512f
C6 VPWR A 0.112f
C7 VGND X 0.977f
C8 VPB VGND 0.0114f
C9 VPWR VGND 0.187f
C10 A VGND 0.115f
C11 X a_110_47# 1.62f
C12 VPB a_110_47# 0.528f
C13 VPB X 0.0315f
C14 VPWR a_110_47# 0.67f
C15 VGND VNB 1.01f
C16 X VNB 0.111f
C17 VPWR VNB 0.835f
C18 A VNB 0.495f
C19 VPB VNB 1.85f
C20 a_110_47# VNB 1.73f
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X a_382_297# a_297_47#
+ a_79_21#
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPWR B1 0.0213f
C1 a_79_21# B1 0.134f
C2 A1 a_297_47# 0.0492f
C3 VGND VPWR 0.0588f
C4 VPWR VPB 0.0624f
C5 VGND a_79_21# 0.129f
C6 a_79_21# VPB 0.0489f
C7 A1 A2 0.102f
C8 VGND B1 0.0182f
C9 VPB B1 0.0328f
C10 a_297_47# A2 0.048f
C11 A1 a_382_297# 2.25e-19
C12 VGND VPB 0.0049f
C13 a_382_297# a_297_47# 8.13e-19
C14 VPWR A1 0.0449f
C15 a_79_21# A1 7.71e-19
C16 a_382_297# A2 0.0145f
C17 VPWR a_297_47# 0.0056f
C18 a_79_21# a_297_47# 0.0326f
C19 VPWR X 0.0958f
C20 a_79_21# X 0.104f
C21 a_297_47# B1 0.00637f
C22 X B1 3.56e-19
C23 VGND A1 0.0157f
C24 A1 VPB 0.0412f
C25 VPWR A2 0.0835f
C26 a_79_21# A2 0.0889f
C27 VGND a_297_47# 0.125f
C28 a_297_47# VPB 7.6e-19
C29 A2 B1 0.0665f
C30 VGND X 0.0736f
C31 X VPB 0.011f
C32 VPWR a_382_297# 0.00566f
C33 a_79_21# a_382_297# 0.00145f
C34 VGND A2 0.0171f
C35 A2 VPB 0.0334f
C36 a_79_21# VPWR 0.201f
C37 VGND a_382_297# 8.23e-19
C38 VGND VNB 0.352f
C39 VPWR VNB 0.304f
C40 X VNB 0.0935f
C41 A1 VNB 0.152f
C42 A2 VNB 0.0981f
C43 B1 VNB 0.101f
C44 VPB VNB 0.605f
C45 a_297_47# VNB 0.0348f
C46 a_79_21# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y a_199_47# a_113_297#
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
C0 VGND a_199_47# 0.00428f
C1 A1 VPB 0.0264f
C2 VPB Y 0.0146f
C3 a_113_297# a_199_47# 2.42e-19
C4 VGND A1 0.078f
C5 VGND Y 0.0654f
C6 A1 a_113_297# 0.05f
C7 a_113_297# Y 0.0909f
C8 VPB VPWR 0.0424f
C9 VGND VPWR 0.037f
C10 A1 a_199_47# 0.00917f
C11 B1 VPB 0.0389f
C12 a_199_47# Y 0.00151f
C13 VPB A2 0.0373f
C14 a_113_297# VPWR 0.177f
C15 VGND B1 0.0436f
C16 VGND A2 0.0495f
C17 A1 Y 0.0813f
C18 B1 a_113_297# 0.00758f
C19 a_199_47# VPWR 4.76e-19
C20 a_113_297# A2 0.0476f
C21 A1 VPWR 0.0154f
C22 VPWR Y 0.0447f
C23 B1 A1 0.0518f
C24 B1 Y 0.113f
C25 A1 A2 0.0912f
C26 A2 Y 0.00122f
C27 B1 VPWR 0.0134f
C28 VGND VPB 0.00548f
C29 A2 VPWR 0.0147f
C30 VPB a_113_297# 0.0108f
C31 VGND a_113_297# 0.00882f
C32 VGND VNB 0.286f
C33 VPWR VNB 0.211f
C34 Y VNB 0.0544f
C35 A2 VNB 0.144f
C36 A1 VNB 0.0981f
C37 B1 VNB 0.162f
C38 VPB VNB 0.428f
C39 a_113_297# VNB 0.034f
.ends

.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X a_114_297# a_304_297# a_220_297#
+ a_32_297#
X0 VPWR A a_304_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X1 a_304_297# B a_220_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND C a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X3 a_220_297# C a_114_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X4 a_32_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_32_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X7 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A a_32_297# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_32_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X11 X a_32_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_32_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X13 a_114_297# D a_32_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X14 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VGND a_32_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 X a_32_297# 0.366f
C1 VGND C 0.0169f
C2 B VGND 0.0177f
C3 VPB C 0.0291f
C4 a_220_297# a_32_297# 0.00132f
C5 VGND D 0.0469f
C6 a_304_297# a_32_297# 0.00167f
C7 A X 0.0157f
C8 VPB B 0.0282f
C9 VPB D 0.0392f
C10 a_304_297# A 7.1e-19
C11 VPB VGND 0.00682f
C12 VPWR a_32_297# 0.153f
C13 B X 0.0046f
C14 A VPWR 0.0525f
C15 a_220_297# C 0.0108f
C16 VPWR a_114_297# 0.00839f
C17 a_220_297# B 0.00641f
C18 a_304_297# B 0.0126f
C19 X VGND 0.245f
C20 VPB X 0.0126f
C21 a_220_297# VGND 0.00137f
C22 A a_32_297# 0.111f
C23 a_304_297# VGND 1e-18
C24 VPWR C 0.044f
C25 a_114_297# a_32_297# 0.0144f
C26 B VPWR 0.0827f
C27 VPWR D 0.0136f
C28 VPWR VGND 0.0835f
C29 C a_32_297# 0.122f
C30 B a_32_297# 0.0415f
C31 VPB VPWR 0.0864f
C32 a_32_297# D 0.106f
C33 a_304_297# X 5.61e-19
C34 C a_114_297# 0.0112f
C35 B A 0.108f
C36 VGND a_32_297# 0.292f
C37 VPB a_32_297# 0.135f
C38 VPWR X 0.358f
C39 A VGND 0.0184f
C40 VGND a_114_297# 0.00223f
C41 B C 0.163f
C42 VPB A 0.031f
C43 a_220_297# VPWR 0.00615f
C44 a_304_297# VPWR 0.00556f
C45 C D 0.0464f
C46 VGND VNB 0.509f
C47 X VNB 0.0584f
C48 VPWR VNB 0.423f
C49 A VNB 0.0911f
C50 B VNB 0.0892f
C51 C VNB 0.0907f
C52 D VNB 0.158f
C53 VPB VNB 0.871f
C54 a_32_297# VNB 0.454f
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y a_129_47# a_47_47# a_285_47#
+ a_377_297#
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 a_377_297# B 0.00254f
C1 a_47_47# VPB 0.0444f
C2 Y A 0.00181f
C3 VGND A 0.0635f
C4 VPB B 0.0643f
C5 VGND a_129_47# 0.00547f
C6 Y VPWR 0.107f
C7 VGND VPWR 0.0665f
C8 a_285_47# A 0.0353f
C9 Y a_47_47# 0.143f
C10 VGND a_47_47# 0.104f
C11 a_285_47# VPWR 0.00255f
C12 Y a_377_297# 0.00188f
C13 VGND a_377_297# 0.00125f
C14 Y B 0.00334f
C15 VGND B 0.0389f
C16 a_285_47# a_47_47# 0.0175f
C17 VPWR A 0.0349f
C18 Y VPB 0.00878f
C19 VGND VPB 0.00568f
C20 a_285_47# B 0.067f
C21 a_129_47# VPWR 9.47e-19
C22 a_47_47# A 0.0307f
C23 a_285_47# VPB 5.53e-19
C24 A B 0.236f
C25 a_129_47# a_47_47# 0.00369f
C26 a_47_47# VPWR 0.273f
C27 a_377_297# VPWR 0.00559f
C28 a_129_47# B 0.00236f
C29 Y VGND 0.0381f
C30 VPWR B 0.0408f
C31 A VPB 0.0822f
C32 a_377_297# a_47_47# 0.00899f
C33 Y a_285_47# 0.0439f
C34 a_47_47# B 0.356f
C35 VGND a_285_47# 0.211f
C36 VPWR VPB 0.0718f
C37 VGND VNB 0.4f
C38 Y VNB 0.0783f
C39 VPWR VNB 0.352f
C40 A VNB 0.217f
C41 B VNB 0.212f
C42 VPB VNB 0.693f
C43 a_285_47# VNB 0.0174f
C44 a_47_47# VNB 0.199f
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 X VGND 0.115f
C1 VPB a_27_47# 0.0686f
C2 VGND VPWR 0.0381f
C3 X A 0.0123f
C4 VPWR A 0.022f
C5 VGND VPB 0.00461f
C6 X VPWR 0.139f
C7 VPB A 0.0335f
C8 X VPB 0.00837f
C9 VGND a_27_47# 0.105f
C10 VPB VPWR 0.0438f
C11 A a_27_47# 0.209f
C12 X a_27_47# 0.165f
C13 VGND A 0.0453f
C14 VPWR a_27_47# 0.167f
C15 VGND VNB 0.263f
C16 X VNB 0.0731f
C17 VPWR VNB 0.221f
C18 A VNB 0.148f
C19 VPB VNB 0.428f
C20 a_27_47# VNB 0.32f
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y a_113_47#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
C0 a_113_47# VPWR 1.78e-19
C1 B Y 0.0481f
C2 Y A 0.0855f
C3 B VPWR 0.0478f
C4 A VPWR 0.0444f
C5 B A 0.051f
C6 VPB Y 0.00618f
C7 VPB VPWR 0.0509f
C8 VGND Y 0.139f
C9 VGND a_113_47# 0.0019f
C10 VPB B 0.0391f
C11 VGND VPWR 0.0322f
C12 VPB A 0.0379f
C13 VGND B 0.0544f
C14 VGND A 0.00949f
C15 VGND VPB 0.0044f
C16 a_113_47# Y 0.00937f
C17 Y VPWR 0.211f
C18 VGND VNB 0.232f
C19 Y VNB 0.0557f
C20 VPWR VNB 0.245f
C21 A VNB 0.143f
C22 B VNB 0.146f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y a_193_297# a_109_297#
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 C VGND 0.0167f
C1 VPB C 0.0369f
C2 B C 0.0936f
C3 VPWR A 0.0477f
C4 VPB VGND 0.00466f
C5 C VPWR 0.0094f
C6 B VGND 0.0192f
C7 B VPB 0.0286f
C8 Y A 0.111f
C9 VPWR VGND 0.0406f
C10 VPB VPWR 0.0471f
C11 C Y 0.0919f
C12 B VPWR 0.013f
C13 a_109_297# VGND 8.05e-19
C14 a_193_297# VGND 6.78e-19
C15 a_109_297# B 0.00897f
C16 B a_193_297# 7.73e-19
C17 Y VGND 0.132f
C18 VPB Y 0.0139f
C19 B Y 0.202f
C20 a_109_297# VPWR 0.00216f
C21 a_193_297# VPWR 0.00239f
C22 Y VPWR 0.171f
C23 VGND A 0.0483f
C24 VPB A 0.0436f
C25 a_109_297# Y 0.0112f
C26 a_193_297# Y 0.0153f
C27 B A 0.0566f
C28 VGND VNB 0.266f
C29 VPWR VNB 0.237f
C30 Y VNB 0.0806f
C31 A VNB 0.177f
C32 B VNB 0.0934f
C33 C VNB 0.144f
C34 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_181_47# a_109_47# a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VGND VPWR 0.0475f
C1 A B 0.0869f
C2 C B 0.0746f
C3 a_109_47# VPWR 3.29e-19
C4 VGND VPB 0.00604f
C5 A VPWR 0.0185f
C6 C VPWR 0.00464f
C7 VGND X 0.0708f
C8 a_27_47# B 0.0625f
C9 VGND a_181_47# 0.00261f
C10 A VPB 0.0426f
C11 C VPB 0.0347f
C12 a_27_47# VPWR 0.145f
C13 C X 0.0149f
C14 C a_181_47# 0.00151f
C15 a_27_47# VPB 0.0501f
C16 VPWR B 0.128f
C17 VGND a_109_47# 0.00123f
C18 X a_27_47# 0.087f
C19 a_27_47# a_181_47# 0.00401f
C20 VPB B 0.0836f
C21 A VGND 0.0154f
C22 C VGND 0.0703f
C23 X B 0.00111f
C24 A a_109_47# 6.45e-19
C25 VPB VPWR 0.0795f
C26 VGND a_27_47# 0.134f
C27 X VPWR 0.0766f
C28 a_27_47# a_109_47# 0.00517f
C29 a_181_47# VPWR 3.97e-19
C30 VGND B 0.00714f
C31 X VPB 0.0121f
C32 A a_27_47# 0.157f
C33 C a_27_47# 0.186f
C34 VGND VNB 0.3f
C35 X VNB 0.0923f
C36 C VNB 0.12f
C37 A VNB 0.174f
C38 VPWR VNB 0.274f
C39 B VNB 0.102f
C40 VPB VNB 0.516f
C41 a_27_47# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X a_103_199# a_253_47#
+ a_337_297# a_253_297#
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.201 pd=1.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.213 ps=1.42 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 B1 VGND 0.0154f
C1 a_337_297# VPWR 0.00348f
C2 a_253_47# A1 0.00334f
C3 VPB VGND 0.00633f
C4 VGND X 0.109f
C5 B1 VPWR 0.019f
C6 a_253_47# VGND 0.2f
C7 VPB VPWR 0.0727f
C8 X VPWR 0.12f
C9 a_103_199# A1 0.123f
C10 VPB B1 0.0344f
C11 B1 X 8.93e-20
C12 a_253_47# a_337_297# 0.00219f
C13 A3 VGND 0.0139f
C14 a_253_47# VPWR 0.00261f
C15 VPB X 0.0155f
C16 a_253_47# B1 0.013f
C17 a_337_297# A3 0.00758f
C18 A3 VPWR 0.011f
C19 a_103_199# VGND 0.102f
C20 a_253_297# VGND 0.00119f
C21 A2 A1 0.0802f
C22 A3 B1 0.0736f
C23 VPB a_253_47# 0.00165f
C24 a_253_47# X 3.38e-19
C25 a_103_199# a_337_297# 0.0101f
C26 a_103_199# VPWR 0.377f
C27 a_253_297# VPWR 0.00267f
C28 VPB A3 0.031f
C29 A3 X 1.42e-19
C30 a_103_199# B1 0.102f
C31 A2 VGND 0.0133f
C32 a_337_297# A2 0.00555f
C33 a_253_47# A3 0.03f
C34 a_103_199# VPB 0.0492f
C35 a_103_199# X 0.0762f
C36 A2 VPWR 0.00974f
C37 a_103_199# a_253_47# 0.0606f
C38 a_253_297# a_253_47# 0.00137f
C39 VPB A2 0.0284f
C40 A2 X 2.55e-19
C41 a_103_199# A3 0.0854f
C42 VGND A1 0.0432f
C43 a_253_47# A2 0.0303f
C44 a_103_199# a_253_297# 0.0148f
C45 A1 VPWR 0.0115f
C46 A2 A3 0.137f
C47 a_337_297# VGND 0.00153f
C48 a_103_199# A2 0.0856f
C49 VGND VPWR 0.0651f
C50 a_253_297# A2 0.00458f
C51 VPB A1 0.0271f
C52 A1 X 7.36e-19
C53 VGND VNB 0.391f
C54 VPWR VNB 0.349f
C55 X VNB 0.0972f
C56 B1 VNB 0.121f
C57 A3 VNB 0.0896f
C58 A2 VNB 0.0885f
C59 A1 VNB 0.0902f
C60 VPB VNB 0.693f
C61 a_253_47# VNB 0.011f
C62 a_103_199# VNB 0.196f
.ends

.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y a_27_297#
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
C0 B VPB 0.121f
C1 VGND VPWR 0.0816f
C2 VPB A 0.12f
C3 VGND Y 0.564f
C4 a_27_297# VPWR 0.6f
C5 VGND B 0.0485f
C6 a_27_297# Y 0.253f
C7 VGND A 0.0864f
C8 a_27_297# B 0.0595f
C9 Y VPWR 0.0299f
C10 VGND VPB 0.00743f
C11 a_27_297# A 0.199f
C12 B VPWR 0.0294f
C13 a_27_297# VPB 0.0259f
C14 VPWR A 0.0795f
C15 B Y 0.354f
C16 Y A 0.165f
C17 VPWR VPB 0.0815f
C18 VGND a_27_297# 0.0127f
C19 B A 0.0625f
C20 Y VPB 0.019f
C21 VGND VNB 0.531f
C22 Y VNB 0.0831f
C23 VPWR VNB 0.401f
C24 B VNB 0.379f
C25 A VNB 0.392f
C26 VPB VNB 0.871f
C27 a_27_297# VNB 0.062f
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y a_27_297#
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 A B 0.0712f
C1 VPWR B 0.0174f
C2 VPB Y 0.00961f
C3 B VPB 0.0566f
C4 a_27_297# Y 0.152f
C5 VPWR A 0.0418f
C6 a_27_297# B 0.0451f
C7 VGND Y 0.289f
C8 A VPB 0.0563f
C9 VPWR VPB 0.05f
C10 B VGND 0.0294f
C11 a_27_297# A 0.0889f
C12 a_27_297# VPWR 0.321f
C13 a_27_297# VPB 0.0203f
C14 A VGND 0.0597f
C15 VPWR VGND 0.0467f
C16 B Y 0.179f
C17 VPB VGND 0.00613f
C18 A Y 0.0523f
C19 a_27_297# VGND 0.00726f
C20 VPWR Y 0.0127f
C21 VGND VNB 0.343f
C22 Y VNB 0.0641f
C23 VPWR VNB 0.249f
C24 B VNB 0.198f
C25 A VNB 0.207f
C26 VPB VNB 0.516f
C27 a_27_297# VNB 0.0647f
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X a_193_297# a_465_47#
+ a_205_47# a_109_297# a_27_47#
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
C0 VPWR a_193_297# 0.169f
C1 VGND a_27_47# 0.395f
C2 A2 VPWR 0.0209f
C3 X VPWR 0.0897f
C4 VPWR a_205_47# 1.62e-19
C5 A1 VPB 0.0343f
C6 B1 a_193_297# 0.00869f
C7 a_109_297# VPB 0.00421f
C8 VPWR A1 0.0161f
C9 X B1 9.58e-20
C10 X a_465_47# 1.56e-19
C11 A2 a_193_297# 0.00683f
C12 VPWR a_109_297# 0.15f
C13 C1 VPB 0.0367f
C14 X a_193_297# 0.00367f
C15 B2 VPB 0.0256f
C16 A1 B1 0.0609f
C17 VGND VPB 0.00844f
C18 A1 a_465_47# 7.06e-19
C19 X A2 0.00157f
C20 C1 VPWR 0.0139f
C21 VPWR B2 0.00842f
C22 B1 a_109_297# 0.00736f
C23 A1 a_193_297# 0.0109f
C24 VPWR VGND 0.0722f
C25 a_27_47# VPB 0.0512f
C26 A2 A1 0.0692f
C27 a_109_297# a_193_297# 0.0927f
C28 X A1 2.77e-19
C29 C1 B1 6.46e-19
C30 B2 B1 0.0784f
C31 B1 VGND 0.0133f
C32 VPWR a_27_47# 0.099f
C33 X a_109_297# 3.99e-19
C34 VGND a_465_47# 0.00257f
C35 B2 a_193_297# 0.00126f
C36 VGND a_193_297# 0.00438f
C37 C1 A2 9.03e-21
C38 A1 a_109_297# 1.05e-19
C39 B1 a_27_47# 0.112f
C40 C1 X 5.03e-20
C41 X B2 6.77e-20
C42 a_27_47# a_465_47# 0.013f
C43 A2 VGND 0.0168f
C44 X VGND 0.061f
C45 VGND a_205_47# 0.00156f
C46 a_27_47# a_193_297# 0.144f
C47 C1 A1 1.77e-20
C48 A1 VGND 0.0126f
C49 A2 a_27_47# 0.153f
C50 X a_27_47# 0.0921f
C51 a_27_47# a_205_47# 0.00762f
C52 VPWR VPB 0.0799f
C53 C1 a_109_297# 0.00739f
C54 B2 a_109_297# 0.0133f
C55 VGND a_109_297# 0.00284f
C56 A1 a_27_47# 0.0984f
C57 B1 VPB 0.0321f
C58 C1 B2 0.0726f
C59 C1 VGND 0.0196f
C60 B2 VGND 0.0174f
C61 a_27_47# a_109_297# 0.0961f
C62 a_193_297# VPB 0.00774f
C63 VPWR B1 0.00982f
C64 VPWR a_465_47# 5.05e-19
C65 A2 VPB 0.027f
C66 C1 a_27_47# 0.0792f
C67 B2 a_27_47# 0.0959f
C68 X VPB 0.0113f
C69 VGND VNB 0.437f
C70 X VNB 0.0919f
C71 VPWR VNB 0.364f
C72 A2 VNB 0.0896f
C73 A1 VNB 0.106f
C74 B1 VNB 0.108f
C75 B2 VNB 0.0887f
C76 C1 VNB 0.139f
C77 VPB VNB 0.782f
C78 a_193_297# VNB 0.0011f
C79 a_109_297# VNB 7.11e-19
C80 a_27_47# VNB 0.216f
.ends

.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X a_548_47# a_639_47#
+ a_476_47# a_174_21# a_505_280# a_27_47#
X0 a_174_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.331 ps=1.71 w=0.42 l=0.15
X2 a_476_47# a_27_47# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.331 pd=1.71 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.141 ps=1.33 w=1 l=0.15
X5 a_548_47# a_505_280# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.109 ps=1.36 w=0.42 l=0.15
X7 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X8 VPWR D a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND D a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VPWR a_505_280# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X11 a_505_280# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X12 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_505_280# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0924 ps=0.86 w=0.42 l=0.15
X14 a_639_47# C a_548_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.064 ps=0.725 w=0.42 l=0.15
X15 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPB VPWR 0.098f
C1 a_548_47# C 0.00375f
C2 a_27_47# A_N 0.134f
C3 a_174_21# VPWR 0.217f
C4 VPB X 0.00317f
C5 a_548_47# a_505_280# 8.83e-19
C6 a_27_47# C 8.75e-19
C7 a_505_280# B_N 0.0891f
C8 a_639_47# D 0.00323f
C9 C D 0.177f
C10 a_174_21# X 0.106f
C11 a_505_280# a_27_47# 0.103f
C12 VGND VPWR 0.0933f
C13 VPB B_N 0.0745f
C14 a_505_280# D 0.0541f
C15 a_476_47# C 0.00125f
C16 a_639_47# C 0.00114f
C17 a_548_47# a_174_21# 0.00101f
C18 a_27_47# VPB 0.106f
C19 VPB D 0.0656f
C20 a_174_21# B_N 4.33e-19
C21 VGND X 0.0746f
C22 a_476_47# a_505_280# 9.37e-20
C23 VPB A_N 0.0969f
C24 a_639_47# a_505_280# 8e-19
C25 a_505_280# C 0.136f
C26 a_174_21# a_27_47# 0.267f
C27 a_174_21# D 0.00723f
C28 a_548_47# VGND 0.00415f
C29 VPB C 0.0541f
C30 a_174_21# A_N 0.0431f
C31 VGND B_N 0.045f
C32 X VPWR 0.0141f
C33 a_476_47# a_174_21# 0.00228f
C34 a_27_47# VGND 0.0942f
C35 a_505_280# VPB 0.105f
C36 a_639_47# a_174_21# 2.58e-19
C37 a_174_21# C 0.0449f
C38 VGND D 0.0513f
C39 a_548_47# VPWR 6.01e-19
C40 VGND A_N 0.0173f
C41 B_N VPWR 0.0156f
C42 a_174_21# a_505_280# 0.145f
C43 a_27_47# VPWR 0.206f
C44 a_476_47# VGND 0.00259f
C45 a_639_47# VGND 0.0041f
C46 VGND C 0.0328f
C47 VPWR D 0.0148f
C48 a_174_21# VPB 0.0845f
C49 A_N VPWR 0.0167f
C50 a_505_280# VGND 0.0924f
C51 a_27_47# X 0.117f
C52 a_476_47# VPWR 5.59e-19
C53 a_639_47# VPWR 5.43e-19
C54 VPWR C 0.0151f
C55 VGND VPB 0.0142f
C56 A_N X 0.00242f
C57 a_505_280# VPWR 0.129f
C58 B_N D 0.117f
C59 a_174_21# VGND 0.143f
C60 VGND VNB 0.548f
C61 X VNB 0.00543f
C62 VPWR VNB 0.446f
C63 B_N VNB 0.162f
C64 D VNB 0.11f
C65 C VNB 0.109f
C66 A_N VNB 0.199f
C67 VPB VNB 0.959f
C68 a_505_280# VNB 0.198f
C69 a_27_47# VNB 0.212f
C70 a_174_21# VNB 0.219f
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X a_109_93# a_368_53# a_209_311#
+ a_296_53#
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0536 ps=0.675 w=0.42 l=0.15
C0 VPWR a_296_53# 1.15e-19
C1 C X 0.0176f
C2 VGND X 0.0647f
C3 X a_209_311# 0.0877f
C4 VPWR a_109_93# 0.0984f
C5 C a_368_53# 0.00415f
C6 VGND a_368_53# 0.0031f
C7 a_368_53# a_209_311# 0.0026f
C8 a_109_93# a_296_53# 1.84e-19
C9 X B 0.00119f
C10 C VPWR 0.005f
C11 VGND VPWR 0.0657f
C12 VPWR a_209_311# 0.155f
C13 VGND a_296_53# 6.07e-19
C14 a_209_311# a_296_53# 0.0049f
C15 X A_N 1.44e-19
C16 C a_109_93# 3.91e-20
C17 VGND a_109_93# 0.0784f
C18 a_109_93# a_209_311# 0.168f
C19 B VPWR 0.131f
C20 VGND C 0.0678f
C21 C a_209_311# 0.19f
C22 VGND a_209_311# 0.131f
C23 B a_109_93# 0.0802f
C24 VPWR A_N 0.0513f
C25 C B 0.0671f
C26 A_N a_109_93# 0.117f
C27 VGND B 0.00796f
C28 B a_209_311# 0.0609f
C29 X VPB 0.0119f
C30 C A_N 7.6e-19
C31 VGND A_N 0.045f
C32 A_N a_209_311# 0.00515f
C33 VPWR VPB 0.104f
C34 B A_N 2.03e-19
C35 VPB a_109_93# 0.0652f
C36 C VPB 0.0339f
C37 VGND VPB 0.00909f
C38 VPB a_209_311# 0.0515f
C39 B VPB 0.0914f
C40 VPB A_N 0.111f
C41 X VPWR 0.0732f
C42 VPWR a_368_53# 4.26e-19
C43 VGND VNB 0.44f
C44 X VNB 0.0925f
C45 C VNB 0.114f
C46 B VNB 0.101f
C47 VPWR VNB 0.342f
C48 A_N VNB 0.197f
C49 VPB VNB 0.693f
C50 a_209_311# VNB 0.143f
C51 a_109_93# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X a_256_47# a_584_47#
+ a_93_21# a_250_297# a_346_47#
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
C0 a_346_47# VGND 0.00514f
C1 VPWR B1 0.01f
C2 VGND A1 0.0133f
C3 a_93_21# A2 0.0747f
C4 a_250_297# B2 0.0344f
C5 a_93_21# VGND 0.251f
C6 VGND A2 0.0114f
C7 VPB B1 0.0276f
C8 VPWR B2 0.0108f
C9 a_256_47# a_93_21# 0.0114f
C10 a_584_47# a_93_21# 0.00278f
C11 a_93_21# A3 0.124f
C12 a_256_47# A2 0.00256f
C13 a_250_297# A1 0.0129f
C14 A3 A2 0.0788f
C15 a_346_47# VPWR 0.00109f
C16 a_256_47# VGND 0.00394f
C17 a_584_47# VGND 0.00683f
C18 VGND A3 0.00974f
C19 VPB B2 0.0355f
C20 a_250_297# a_93_21# 0.188f
C21 X B1 3.83e-20
C22 VPWR A1 0.016f
C23 a_250_297# A2 0.0129f
C24 a_256_47# A3 4.42e-19
C25 a_250_297# VGND 0.0072f
C26 a_93_21# VPWR 0.0907f
C27 VPWR A2 0.0133f
C28 VPB A1 0.0296f
C29 VPWR VGND 0.076f
C30 a_584_47# a_250_297# 2.43e-19
C31 a_250_297# A3 0.00602f
C32 VPB a_93_21# 0.0485f
C33 VPB A2 0.0287f
C34 a_256_47# VPWR 9.47e-19
C35 a_584_47# VPWR 9.47e-19
C36 VPWR A3 0.0158f
C37 VPB VGND 0.00788f
C38 X A1 6.03e-20
C39 B2 B1 0.0823f
C40 a_250_297# VPWR 0.313f
C41 a_93_21# X 0.0841f
C42 VPB A3 0.0291f
C43 X A2 1.19e-19
C44 a_346_47# B1 5.39e-20
C45 X VGND 0.06f
C46 A1 B1 0.0965f
C47 VPB a_250_297# 0.00616f
C48 a_93_21# B1 0.0774f
C49 X A3 2.45e-19
C50 B1 A2 1.44e-20
C51 VPB VPWR 0.0756f
C52 A1 B2 3.14e-19
C53 VGND B1 0.0344f
C54 a_250_297# X 5.42e-19
C55 a_93_21# B2 0.0147f
C56 a_256_47# B1 2.07e-20
C57 a_346_47# A1 0.00465f
C58 a_584_47# B1 0.00143f
C59 B1 A3 7.88e-22
C60 B2 A2 1.46e-19
C61 X VPWR 0.0849f
C62 VGND B2 0.0469f
C63 a_346_47# a_93_21# 0.0119f
C64 a_346_47# A2 0.00252f
C65 a_250_297# B1 0.0125f
C66 a_93_21# A1 0.0641f
C67 VPB X 0.0108f
C68 A1 A2 0.0971f
C69 B2 A3 9.12e-20
C70 VGND VNB 0.465f
C71 VPWR VNB 0.365f
C72 X VNB 0.0937f
C73 B2 VNB 0.14f
C74 B1 VNB 0.101f
C75 A1 VNB 0.0951f
C76 A2 VNB 0.0921f
C77 A3 VNB 0.0929f
C78 VPB VNB 0.782f
C79 a_250_297# VNB 0.0278f
C80 a_93_21# VNB 0.151f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPWR a_303_47# 4.83e-19
C1 B C 0.161f
C2 D C 0.18f
C3 B a_27_47# 0.13f
C4 D a_27_47# 0.107f
C5 VGND a_109_47# 0.00223f
C6 X VPB 0.0111f
C7 VGND VPB 0.00852f
C8 VPWR a_109_47# 4.66e-19
C9 VPB VPWR 0.077f
C10 B A 0.0839f
C11 VGND a_197_47# 0.00387f
C12 VPWR a_197_47# 5.24e-19
C13 C VGND 0.0408f
C14 C VPWR 0.021f
C15 X a_27_47# 0.0754f
C16 VGND a_27_47# 0.132f
C17 VPWR a_27_47# 0.326f
C18 VGND A 0.0151f
C19 C a_303_47# 0.00527f
C20 VPWR A 0.044f
C21 a_303_47# a_27_47# 0.00119f
C22 B VGND 0.0453f
C23 X D 0.00746f
C24 D VGND 0.0898f
C25 B VPWR 0.0231f
C26 C a_109_47# 1.72e-20
C27 D VPWR 0.0207f
C28 C VPB 0.0609f
C29 a_27_47# a_109_47# 0.00578f
C30 VPB a_27_47# 0.082f
C31 D a_303_47# 0.00119f
C32 C a_197_47# 0.00123f
C33 VPB A 0.0907f
C34 a_27_47# a_197_47# 0.00167f
C35 X VGND 0.0903f
C36 B a_109_47# 0.00153f
C37 C a_27_47# 0.0516f
C38 X VPWR 0.0945f
C39 VGND VPWR 0.0662f
C40 B VPB 0.0643f
C41 D VPB 0.0782f
C42 B a_197_47# 0.00623f
C43 a_27_47# A 0.153f
C44 VGND a_303_47# 0.00381f
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X a_27_47#
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_27_47# VGND 0.163f
C1 X VGND 0.23f
C2 a_27_47# X 0.207f
C3 A VGND 0.0194f
C4 VPWR VGND 0.072f
C5 VPB VGND 0.00796f
C6 A a_27_47# 0.17f
C7 a_27_47# VPWR 0.218f
C8 A X 4.66e-19
C9 VPWR X 0.333f
C10 a_27_47# VPB 0.132f
C11 VPB X 0.00899f
C12 A VPWR 0.016f
C13 A VPB 0.0361f
C14 VPWR VPB 0.0711f
C15 VGND VNB 0.378f
C16 X VNB 0.039f
C17 VPWR VNB 0.325f
C18 A VNB 0.14f
C19 VPB VNB 0.605f
C20 a_27_47# VNB 0.461f
.ends

.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y a_655_47# a_465_47#
+ a_215_47# a_27_47#
X0 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_465_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VGND D a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X3 a_215_47# B a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_655_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_655_47# C a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.37 pd=1.74 as=0.135 ps=1.27 w=1 l=0.15
X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_465_47# C a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=2.8 as=0.135 ps=1.27 w=1 l=0.15
X13 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X14 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.37 ps=1.74 w=1 l=0.15
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
C0 D a_655_47# 0.0973f
C1 C B 0.0362f
C2 B VGND 0.0218f
C3 a_27_47# VGND 0.109f
C4 VPWR a_215_47# 0.00471f
C5 Y a_215_47# 0.0832f
C6 VPWR VPB 0.132f
C7 Y VPB 0.0192f
C8 VPB D 0.0786f
C9 A_N a_27_47# 0.155f
C10 VPWR a_465_47# 0.00194f
C11 Y a_465_47# 0.00307f
C12 a_655_47# a_215_47# 0.0234f
C13 VPB a_655_47# 4.11e-19
C14 VPWR B 0.035f
C15 C VGND 0.0214f
C16 B Y 0.152f
C17 VPWR a_27_47# 0.186f
C18 Y a_27_47# 0.0941f
C19 a_655_47# a_465_47# 0.0905f
C20 A_N VGND 0.0171f
C21 VPB a_215_47# 2.32e-19
C22 B a_655_47# 3.69e-19
C23 a_465_47# a_215_47# 0.089f
C24 VPB a_465_47# 2.49e-19
C25 VPWR C 0.035f
C26 VPWR VGND 0.112f
C27 C Y 0.133f
C28 Y VGND 0.018f
C29 B a_215_47# 0.109f
C30 C D 0.0696f
C31 D VGND 0.0336f
C32 B VPB 0.071f
C33 a_27_47# a_215_47# 0.0716f
C34 VPWR A_N 0.0201f
C35 Y A_N 0.00283f
C36 VPB a_27_47# 0.0973f
C37 C a_655_47# 0.115f
C38 a_655_47# VGND 0.178f
C39 B a_465_47# 0.0119f
C40 A_N a_655_47# 2.96e-19
C41 VPWR Y 0.82f
C42 B a_27_47# 0.0532f
C43 C a_215_47# 7.48e-20
C44 a_215_47# VGND 0.16f
C45 VPWR D 0.0768f
C46 Y D 0.0577f
C47 C VPB 0.0658f
C48 VPB VGND 0.0109f
C49 A_N a_215_47# 0.00211f
C50 A_N VPB 0.106f
C51 VPWR a_655_47# 0.00433f
C52 Y a_655_47# 0.0111f
C53 C a_465_47# 0.00942f
C54 a_465_47# VGND 0.182f
C55 VGND VNB 0.63f
C56 Y VNB 0.0153f
C57 VPWR VNB 0.547f
C58 D VNB 0.246f
C59 C VNB 0.195f
C60 B VNB 0.208f
C61 A_N VNB 0.209f
C62 VPB VNB 1.14f
C63 a_655_47# VNB 0.0373f
C64 a_465_47# VNB 0.01f
C65 a_215_47# VNB 0.0194f
C66 a_27_47# VNB 0.283f
.ends

.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y a_388_297# a_297_47#
+ a_105_352#
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
C0 a_297_47# VGND 0.163f
C1 A2 Y 0.0526f
C2 a_105_352# VPB 0.0584f
C3 A1 VPB 0.034f
C4 a_297_47# VPWR 0.00498f
C5 a_105_352# A2 0.0533f
C6 A2 A1 0.0751f
C7 VPB B1_N 0.144f
C8 VGND VPWR 0.0578f
C9 a_297_47# Y 0.0476f
C10 a_105_352# a_297_47# 0.00424f
C11 VGND Y 0.0397f
C12 a_297_47# A1 0.055f
C13 a_388_297# A2 0.00169f
C14 A2 VPB 0.0263f
C15 a_105_352# VGND 0.0687f
C16 a_297_47# B1_N 5.28e-19
C17 VGND A1 0.0148f
C18 Y VPWR 0.154f
C19 VGND B1_N 0.0552f
C20 a_105_352# VPWR 0.085f
C21 a_388_297# a_297_47# 0.0023f
C22 a_297_47# VPB 7.84e-19
C23 A1 VPWR 0.0533f
C24 A2 a_297_47# 0.0544f
C25 a_388_297# VGND 0.00201f
C26 VGND VPB 0.00719f
C27 a_105_352# Y 0.137f
C28 VPWR B1_N 0.0709f
C29 A1 Y 0.00408f
C30 A2 VGND 0.0152f
C31 a_388_297# VPWR 0.0132f
C32 VPWR VPB 0.0754f
C33 Y B1_N 0.0049f
C34 A2 VPWR 0.0247f
C35 a_105_352# B1_N 0.172f
C36 a_388_297# Y 0.00711f
C37 Y VPB 0.00665f
C38 VGND VNB 0.384f
C39 Y VNB 0.0183f
C40 VPWR VNB 0.327f
C41 A1 VNB 0.134f
C42 A2 VNB 0.0904f
C43 B1_N VNB 0.232f
C44 VPB VNB 0.605f
C45 a_297_47# VNB 0.0343f
C46 a_105_352# VNB 0.149f
.ends

.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y a_27_93# a_206_47#
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
C0 B a_27_93# 0.177f
C1 VPWR VPB 0.0788f
C2 A_N a_27_93# 0.0854f
C3 Y a_27_93# 0.144f
C4 VGND a_206_47# 0.00612f
C5 VPWR VGND 0.0468f
C6 A_N B 0.0602f
C7 Y B 0.00954f
C8 VPB a_27_93# 0.0511f
C9 Y A_N 0.00194f
C10 VGND a_27_93# 0.1f
C11 VPB B 0.0322f
C12 VPWR a_206_47# 8.87e-19
C13 A_N VPB 0.0445f
C14 Y VPB 0.0264f
C15 VGND B 0.0181f
C16 A_N VGND 0.0118f
C17 Y VGND 0.109f
C18 a_27_93# a_206_47# 0.00698f
C19 VPWR a_27_93# 0.0714f
C20 VGND VPB 0.00942f
C21 VPWR B 0.0176f
C22 Y a_206_47# 0.00332f
C23 A_N VPWR 0.00835f
C24 Y VPWR 0.184f
C25 VGND VNB 0.312f
C26 Y VNB 0.0943f
C27 A_N VNB 0.145f
C28 VPWR VNB 0.279f
C29 B VNB 0.102f
C30 VPB VNB 0.516f
C31 a_27_93# VNB 0.168f
.ends

.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X a_215_297# a_27_413#
+ a_298_297# a_382_47#
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.136 ps=1.1 w=0.65 l=0.15
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.258 ps=1.45 w=0.65 l=0.15
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.1 as=0.111 ps=1.37 w=0.42 l=0.15
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.258 pd=1.45 as=0.091 ps=0.93 w=0.65 l=0.15
C0 B1_N VGND 0.0492f
C1 a_215_297# VPWR 0.13f
C2 X A1 1.5e-19
C3 VPB A2 0.0417f
C4 a_27_413# B1_N 0.237f
C5 a_298_297# A1 0.0494f
C6 a_382_47# A1 5.63e-19
C7 X A2 0.00569f
C8 a_215_297# A1 0.093f
C9 B1_N VPB 0.103f
C10 B1_N X 2.01e-19
C11 a_298_297# A2 0.0357f
C12 a_27_413# VGND 0.0982f
C13 VPWR A1 0.0215f
C14 a_215_297# A2 0.0949f
C15 VPB VGND 0.0117f
C16 a_298_297# B1_N 8.44e-19
C17 B1_N a_215_297# 0.00479f
C18 VPWR A2 0.0307f
C19 a_27_413# VPB 0.0987f
C20 X VGND 0.0573f
C21 B1_N VPWR 0.019f
C22 a_27_413# X 4.11e-20
C23 a_298_297# VGND 0.00393f
C24 a_382_47# VGND 0.0053f
C25 A2 A1 0.112f
C26 a_215_297# VGND 0.272f
C27 VPB X 0.0117f
C28 a_298_297# a_27_413# 0.00498f
C29 B1_N A1 1.31e-20
C30 a_27_413# a_215_297# 0.141f
C31 VPWR VGND 0.0789f
C32 a_298_297# VPB 0.00345f
C33 VPB a_215_297# 0.0546f
C34 a_27_413# VPWR 0.107f
C35 B1_N A2 4.62e-21
C36 a_382_47# X 5.12e-19
C37 a_215_297# X 0.0802f
C38 VGND A1 0.0144f
C39 VPB VPWR 0.0976f
C40 a_298_297# a_382_47# 1.58e-20
C41 a_27_413# A1 0.0573f
C42 a_298_297# a_215_297# 0.0718f
C43 a_382_47# a_215_297# 0.0105f
C44 VPWR X 0.115f
C45 VGND A2 0.0197f
C46 VPB A1 0.0277f
C47 a_298_297# VPWR 0.196f
C48 a_382_47# VPWR 8.53e-19
C49 a_27_413# A2 8.92e-20
C50 VGND VNB 0.44f
C51 X VNB 0.089f
C52 VPWR VNB 0.366f
C53 A2 VNB 0.108f
C54 A1 VNB 0.0893f
C55 B1_N VNB 0.29f
C56 VPB VNB 0.782f
C57 a_298_297# VNB 0.0039f
C58 a_215_297# VNB 0.153f
C59 a_27_413# VNB 0.172f
.ends

.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X a_396_47# a_206_47# a_490_47#
+ a_314_297# a_204_297# a_27_47#
X0 a_204_297# A1 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.16 ps=1.32 w=1 l=0.15
X1 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR S a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 a_204_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.162 ps=1.33 w=1 l=0.15
X5 a_396_47# A0 a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.26 ps=2.52 w=1 l=0.15
X6 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.109 ps=0.985 w=0.65 l=0.15
X7 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 a_490_47# A1 a_396_47# VNB sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.104 ps=0.97 w=0.65 l=0.15
X11 VGND S a_490_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.275 ps=1.5 w=0.65 l=0.15
X12 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 a_396_47# A0 a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.26 ps=1.45 w=0.65 l=0.15
X14 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X15 VPWR S a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X16 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND S a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
C0 S a_204_297# 0.0097f
C1 a_314_297# a_27_47# 7.66e-19
C2 VGND a_396_47# 0.257f
C3 A0 a_27_47# 0.0551f
C4 A1 a_27_47# 9.52e-20
C5 a_314_297# a_396_47# 0.12f
C6 S a_27_47# 0.208f
C7 a_490_47# S 0.0127f
C8 VPB X 0.0118f
C9 VPWR X 0.299f
C10 A0 a_396_47# 0.00958f
C11 a_206_47# VPWR 0.00256f
C12 A1 a_396_47# 0.0444f
C13 a_204_297# a_27_47# 0.0153f
C14 S a_396_47# 0.297f
C15 VGND X 0.222f
C16 VGND a_206_47# 0.0161f
C17 VPB VPWR 0.119f
C18 a_314_297# X 0.0111f
C19 a_204_297# a_396_47# 0.0127f
C20 VPB VGND 0.0113f
C21 a_314_297# a_206_47# 5.08e-20
C22 VGND VPWR 0.108f
C23 a_490_47# a_27_47# 2.12e-19
C24 A0 X 5.48e-20
C25 A1 X 8.93e-20
C26 VPB a_314_297# 0.00854f
C27 a_314_297# VPWR 0.0706f
C28 S X 0.00188f
C29 A0 a_206_47# 6.55e-19
C30 a_396_47# a_27_47# 0.00537f
C31 S a_206_47# 0.0209f
C32 a_490_47# a_396_47# 0.0245f
C33 VGND a_314_297# 0.00385f
C34 A0 VPB 0.0475f
C35 A0 VPWR 0.0115f
C36 VPB A1 0.0325f
C37 A1 VPWR 0.00928f
C38 a_204_297# X 3.48e-19
C39 VPB S 0.0837f
C40 S VPWR 0.0403f
C41 a_204_297# a_206_47# 1.91e-19
C42 A0 VGND 0.0151f
C43 A1 VGND 0.0108f
C44 VGND S 0.133f
C45 VPB a_204_297# 0.0121f
C46 a_204_297# VPWR 0.227f
C47 a_27_47# X 3.79e-19
C48 A0 a_314_297# 0.0263f
C49 A1 a_314_297# 0.00665f
C50 a_490_47# X 2e-19
C51 S a_314_297# 0.00998f
C52 a_206_47# a_27_47# 0.00106f
C53 VGND a_204_297# 0.00392f
C54 A0 A1 0.0812f
C55 VPB a_27_47# 0.0485f
C56 a_27_47# VPWR 0.152f
C57 a_396_47# X 0.305f
C58 A0 S 0.0358f
C59 A1 S 0.0942f
C60 a_204_297# a_314_297# 0.14f
C61 a_490_47# VPWR 0.00182f
C62 a_206_47# a_396_47# 0.00414f
C63 VGND a_27_47# 0.0676f
C64 VGND a_490_47# 0.00792f
C65 A0 a_204_297# 0.00948f
C66 A1 a_204_297# 0.00593f
C67 VPB a_396_47# 0.135f
C68 a_396_47# VPWR 0.121f
C69 VGND VNB 0.632f
C70 X VNB 0.075f
C71 VPWR VNB 0.536f
C72 A1 VNB 0.098f
C73 A0 VNB 0.115f
C74 S VNB 0.265f
C75 VPB VNB 1.14f
C76 a_314_297# VNB 0.00495f
C77 a_204_297# VNB 0.00597f
C78 a_396_47# VNB 0.407f
C79 a_27_47# VNB 0.191f
.ends

.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y a_109_297# a_27_47#
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_27_47# VGND 0.142f
C1 A2 Y 0.124f
C2 B1 VPB 0.0741f
C3 a_27_47# VPWR 0.00663f
C4 B1 A2 0.0472f
C5 VPB A1 0.0327f
C6 VGND VPWR 0.0381f
C7 a_27_47# Y 0.0517f
C8 A2 A1 0.0986f
C9 B1 a_27_47# 0.00471f
C10 VGND Y 0.0289f
C11 a_109_297# A2 0.00993f
C12 A2 VPB 0.0305f
C13 B1 VGND 0.016f
C14 a_27_47# A1 0.037f
C15 Y VPWR 0.105f
C16 VGND A1 0.0163f
C17 B1 VPWR 0.0433f
C18 a_109_297# a_27_47# 5.37e-19
C19 a_27_47# VPB 8.4e-19
C20 A2 a_27_47# 0.0388f
C21 a_109_297# VGND 4.56e-19
C22 VGND VPB 0.00462f
C23 VPWR A1 0.0497f
C24 B1 Y 0.0811f
C25 A2 VGND 0.0183f
C26 a_109_297# VPWR 0.00401f
C27 VPWR VPB 0.056f
C28 Y A1 8.9e-19
C29 A2 VPWR 0.109f
C30 a_109_297# Y 5.24e-19
C31 Y VPB 0.00672f
C32 VGND VNB 0.254f
C33 Y VNB 0.0545f
C34 VPWR VNB 0.271f
C35 B1 VNB 0.152f
C36 A2 VNB 0.0962f
C37 A1 VNB 0.138f
C38 VPB VNB 0.428f
C39 a_27_47# VNB 0.0311f
.ends

.subckt sarlogic VGND VPWR cal clk clkc comp ctln[0] ctln[1] ctln[2] ctln[3] ctln[4]
+ ctln[5] ctln[6] ctln[7] ctlp[0] ctlp[1] ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6]
+ ctlp[7] en result[0] result[1] result[2] result[3] result[4] result[5] result[6]
+ result[7] rstn sample trim[0] trim[1] trim[2] trim[3] trim[4] trimb[0] trimb[1]
+ trimb[2] trimb[3] trimb[4] valid
X_294_ net2 cal_count\[2\] VGND VGND VPWR VPWR _130_ _294_/a_150_297# _294_/a_68_297#
+ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_0_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_277_ _117_ VGND VGND VPWR VPWR _032_ _277_/a_75_212# sky130_fd_sc_hd__clkbuf_1
X_200_ cal_itt\[1\] cal_itt\[0\] cal_itt\[2\] _062_ VGND VGND VPWR VPWR _071_ _200_/a_80_21#
+ _200_/a_209_297# _200_/a_209_47# _200_/a_303_47# sky130_fd_sc_hd__a31o_1
X_329_ clknet_2_2__leaf_clk _026_ net46 VGND VGND VPWR VPWR trim_mask\[2\] _329_/a_1462_47#
+ _329_/a_543_47# _329_/a_651_413# _329_/a_193_47# _329_/a_805_47# _329_/a_448_47#
+ _329_/a_639_47# _329_/a_1283_21# _329_/a_761_289# _329_/a_1108_47# _329_/a_1217_47#
+ _329_/a_1270_413# _329_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput31 net31 VGND VGND VPWR VPWR trim[0] output31/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput20 net20 VGND VGND VPWR VPWR ctlp[6] output20/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput7 net7 VGND VGND VPWR VPWR ctln[1] output7/a_27_47# sky130_fd_sc_hd__buf_2
X_293_ cal_count\[0\] _126_ _125_ VGND VGND VPWR VPWR _129_ _293_/a_384_47# _293_/a_81_21#
+ _293_/a_299_297# sky130_fd_sc_hd__a21o_1
XFILLER_0_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_276_ _110_ _116_ VGND VGND VPWR VPWR _117_ _276_/a_145_75# _276_/a_59_75# sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_259_ trim_mask\[3\] _104_ _064_ trim_mask\[4\] VGND VGND VPWR VPWR _027_ _259_/a_27_297#
+ _259_/a_109_47# _259_/a_109_297# _259_/a_373_47# sky130_fd_sc_hd__a22o_1
X_328_ clknet_2_2__leaf_clk _025_ net46 VGND VGND VPWR VPWR trim_mask\[1\] _328_/a_1462_47#
+ _328_/a_543_47# _328_/a_651_413# _328_/a_193_47# _328_/a_805_47# _328_/a_448_47#
+ _328_/a_639_47# _328_/a_1283_21# _328_/a_761_289# _328_/a_1108_47# _328_/a_1217_47#
+ _328_/a_1270_413# _328_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput32 net32 VGND VGND VPWR VPWR trim[1] output32/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput21 net21 VGND VGND VPWR VPWR ctlp[7] output21/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput10 net10 VGND VGND VPWR VPWR ctln[4] output10/a_27_47# sky130_fd_sc_hd__buf_2
Xoutput8 net8 VGND VGND VPWR VPWR ctln[2] output8/a_27_47# sky130_fd_sc_hd__buf_2
X_292_ cal_count\[1\] _122_ _128_ _123_ VGND VGND VPWR VPWR _036_ _292_/a_78_199#
+ _292_/a_493_297# _292_/a_215_47# _292_/a_292_297# sky130_fd_sc_hd__o22a_1
XFILLER_0_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_275_ trim_mask\[3\] net50 trim_val\[3\] VGND VGND VPWR VPWR _116_ _275_/a_384_47#
+ _275_/a_81_21# _275_/a_299_297# sky130_fd_sc_hd__a21o_1
X_189_ _051_ _050_ _048_ VGND VGND VPWR VPWR _062_ _189_/a_408_47# _189_/a_218_47#
+ _189_/a_27_47# sky130_fd_sc_hd__nand3b_2
X_258_ trim_mask\[2\] _104_ _064_ trim_mask\[3\] VGND VGND VPWR VPWR _026_ _258_/a_27_297#
+ _258_/a_109_47# _258_/a_109_297# _258_/a_373_47# sky130_fd_sc_hd__a22o_1
X_327_ clknet_2_2__leaf_clk _024_ net46 VGND VGND VPWR VPWR trim_mask\[0\] _327_/a_1462_47#
+ _327_/a_543_47# _327_/a_651_413# _327_/a_193_47# _327_/a_805_47# _327_/a_448_47#
+ _327_/a_639_47# _327_/a_1283_21# _327_/a_761_289# _327_/a_1108_47# _327_/a_1217_47#
+ _327_/a_1270_413# _327_/a_27_47# sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput33 net33 VGND VGND VPWR VPWR trim[2] output33/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput22 net22 VGND VGND VPWR VPWR result[0] output22/a_27_47# sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR ctln[5] output11/a_27_47# sky130_fd_sc_hd__buf_2
Xoutput9 net9 VGND VGND VPWR VPWR ctln[3] output9/a_27_47# sky130_fd_sc_hd__buf_2
XFILLER_0_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_291_ cal_count\[0\] _127_ VGND VGND VPWR VPWR _128_ _291_/a_117_297# _291_/a_285_297#
+ _291_/a_285_47# _291_/a_35_297# sky130_fd_sc_hd__xor2_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_19_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_274_ _115_ VGND VGND VPWR VPWR _031_ _274_/a_75_212# sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_188_ _061_ VGND VGND VPWR VPWR net5 _188_/a_27_47# sky130_fd_sc_hd__buf_1
X_257_ trim_mask\[1\] _104_ _064_ trim_mask\[2\] VGND VGND VPWR VPWR _025_ _257_/a_27_297#
+ _257_/a_109_47# _257_/a_109_297# _257_/a_373_47# sky130_fd_sc_hd__a22o_1
X_326_ clknet_2_1__leaf_clk _023_ net43 VGND VGND VPWR VPWR mask\[7\] _326_/a_1462_47#
+ _326_/a_543_47# _326_/a_651_413# _326_/a_193_47# _326_/a_805_47# _326_/a_448_47#
+ _326_/a_639_47# _326_/a_1283_21# _326_/a_761_289# _326_/a_1108_47# _326_/a_1217_47#
+ _326_/a_1270_413# _326_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_309_ clknet_2_1__leaf_clk _006_ net43 VGND VGND VPWR VPWR net24 _309_/a_1462_47#
+ _309_/a_543_47# _309_/a_651_413# _309_/a_193_47# _309_/a_805_47# _309_/a_448_47#
+ _309_/a_639_47# _309_/a_1283_21# _309_/a_761_289# _309_/a_1108_47# _309_/a_1217_47#
+ _309_/a_1270_413# _309_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_7_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput34 net34 VGND VGND VPWR VPWR trim[3] output34/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput23 net23 VGND VGND VPWR VPWR result[1] output23/a_27_47# sky130_fd_sc_hd__buf_2
Xoutput12 net12 VGND VGND VPWR VPWR ctln[6] output12/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_290_ _125_ _126_ VGND VGND VPWR VPWR _127_ _290_/a_27_413# _290_/a_297_47# _290_/a_207_413#
+ sky130_fd_sc_hd__and2b_1
X_273_ _110_ _114_ VGND VGND VPWR VPWR _115_ _273_/a_145_75# _273_/a_59_75# sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_20_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_187_ clknet_2_3__leaf_clk en_co_clk VGND VGND VPWR VPWR _061_ _187_/a_212_413# _187_/a_27_413#
+ _187_/a_297_47# sky130_fd_sc_hd__and2b_2
X_256_ trim_mask\[0\] _104_ _064_ trim_mask\[1\] VGND VGND VPWR VPWR _024_ _256_/a_27_297#
+ _256_/a_109_47# _256_/a_109_297# _256_/a_373_47# sky130_fd_sc_hd__a22o_1
X_325_ clknet_2_1__leaf_clk _022_ net43 VGND VGND VPWR VPWR mask\[6\] _325_/a_1462_47#
+ _325_/a_543_47# _325_/a_651_413# _325_/a_193_47# _325_/a_805_47# _325_/a_448_47#
+ _325_/a_639_47# _325_/a_1283_21# _325_/a_761_289# _325_/a_1108_47# _325_/a_1217_47#
+ _325_/a_1270_413# _325_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_239_ _050_ calibrate _048_ _051_ VGND VGND VPWR VPWR _098_ _239_/a_277_297# _239_/a_27_297#
+ _239_/a_694_21# _239_/a_474_297# sky130_fd_sc_hd__nor4b_2
X_308_ clknet_2_0__leaf_clk _005_ net43 VGND VGND VPWR VPWR net23 _308_/a_1462_47#
+ _308_/a_543_47# _308_/a_651_413# _308_/a_193_47# _308_/a_805_47# _308_/a_448_47#
+ _308_/a_639_47# _308_/a_1283_21# _308_/a_761_289# _308_/a_1108_47# _308_/a_1217_47#
+ _308_/a_1270_413# _308_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput35 net35 VGND VGND VPWR VPWR trim[4] output35/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput24 net24 VGND VGND VPWR VPWR result[2] output24/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput13 net13 VGND VGND VPWR VPWR ctln[7] output13/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_272_ trim_mask\[2\] net48 trim_val\[2\] VGND VGND VPWR VPWR _114_ _272_/a_384_47#
+ _272_/a_81_21# _272_/a_299_297# sky130_fd_sc_hd__a21o_1
X_341_ clknet_2_3__leaf_clk _038_ net46 VGND VGND VPWR VPWR cal_count\[3\] _341_/a_1462_47#
+ _341_/a_543_47# _341_/a_651_413# _341_/a_193_47# _341_/a_805_47# _341_/a_448_47#
+ _341_/a_639_47# _341_/a_1283_21# _341_/a_761_289# _341_/a_1108_47# _341_/a_1217_47#
+ _341_/a_1270_413# _341_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_186_ _059_ _060_ VGND VGND VPWR VPWR net41 _186_/a_109_297# sky130_fd_sc_hd__nor2_1
X_255_ net30 _103_ VGND VGND VPWR VPWR _104_ _255_/a_27_47# sky130_fd_sc_hd__nand2_2
X_324_ clknet_2_1__leaf_clk _021_ net44 VGND VGND VPWR VPWR mask\[5\] _324_/a_1462_47#
+ _324_/a_543_47# _324_/a_651_413# _324_/a_193_47# _324_/a_805_47# _324_/a_448_47#
+ _324_/a_639_47# _324_/a_1283_21# _324_/a_761_289# _324_/a_1108_47# _324_/a_1217_47#
+ _324_/a_1270_413# _324_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_169_ state\[1\] state\[2\] state\[0\] VGND VGND VPWR VPWR _053_ _169_/a_373_53#
+ _169_/a_215_311# _169_/a_301_53# _169_/a_109_53# sky130_fd_sc_hd__and3b_2
X_238_ _097_ VGND VGND VPWR VPWR _013_ _238_/a_75_212# sky130_fd_sc_hd__clkbuf_1
X_307_ clknet_2_0__leaf_clk _004_ net45 VGND VGND VPWR VPWR net22 _307_/a_1462_47#
+ _307_/a_543_47# _307_/a_651_413# _307_/a_193_47# _307_/a_805_47# _307_/a_448_47#
+ _307_/a_639_47# _307_/a_1283_21# _307_/a_761_289# _307_/a_1108_47# _307_/a_1217_47#
+ _307_/a_1270_413# _307_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput36 net36 VGND VGND VPWR VPWR trimb[0] output36/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput25 net25 VGND VGND VPWR VPWR result[3] output25/a_27_47# sky130_fd_sc_hd__buf_2
Xoutput14 net14 VGND VGND VPWR VPWR ctlp[0] output14/a_27_47# sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_271_ _113_ VGND VGND VPWR VPWR _030_ _271_/a_75_212# sky130_fd_sc_hd__clkbuf_1
X_340_ clknet_2_3__leaf_clk _037_ net47 VGND VGND VPWR VPWR cal_count\[2\] _340_/a_1140_413#
+ _340_/a_1296_47# _340_/a_1182_261# _340_/a_586_47# _340_/a_1602_47# _340_/a_956_413#
+ _340_/a_1224_47# _340_/a_193_47# _340_/a_796_47# _340_/a_381_47# _340_/a_1056_47#
+ _340_/a_1032_413# _340_/a_562_413# _340_/a_652_21# _340_/a_476_47# _340_/a_27_47#
+ sky130_fd_sc_hd__dfstp_1
X_185_ net54 state\[0\] VGND VGND VPWR VPWR _060_ _185_/a_150_297# _185_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_254_ _092_ net42 VGND VGND VPWR VPWR _103_ _254_/a_109_297# sky130_fd_sc_hd__nor2_1
X_323_ clknet_2_1__leaf_clk _020_ net47 VGND VGND VPWR VPWR mask\[4\] _323_/a_1462_47#
+ _323_/a_543_47# _323_/a_651_413# _323_/a_193_47# _323_/a_805_47# _323_/a_448_47#
+ _323_/a_639_47# _323_/a_1283_21# _323_/a_761_289# _323_/a_1108_47# _323_/a_1217_47#
+ _323_/a_1270_413# _323_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_168_ _050_ _051_ VGND VGND VPWR VPWR _052_ _168_/a_27_413# _168_/a_297_47# _168_/a_207_413#
+ sky130_fd_sc_hd__and2b_1
X_237_ _048_ _090_ _096_ VGND VGND VPWR VPWR _097_ _237_/a_505_21# _237_/a_535_374#
+ _237_/a_439_47# _237_/a_218_47# _237_/a_76_199# _237_/a_218_374# sky130_fd_sc_hd__mux2_1
X_306_ clknet_2_0__leaf_clk _003_ net44 VGND VGND VPWR VPWR cal_itt\[3\] _306_/a_1462_47#
+ _306_/a_543_47# _306_/a_651_413# _306_/a_193_47# _306_/a_805_47# _306_/a_448_47#
+ _306_/a_639_47# _306_/a_1283_21# _306_/a_761_289# _306_/a_1108_47# _306_/a_1217_47#
+ _306_/a_1270_413# _306_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_34 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput37 net37 VGND VGND VPWR VPWR trimb[1] output37/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput26 net26 VGND VGND VPWR VPWR result[4] output26/a_27_47# sky130_fd_sc_hd__buf_2
Xoutput15 net15 VGND VGND VPWR VPWR ctlp[1] output15/a_27_47# sky130_fd_sc_hd__buf_2
XFILLER_0_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_270_ _110_ _112_ VGND VGND VPWR VPWR _113_ _270_/a_145_75# _270_/a_59_75# sky130_fd_sc_hd__and2_1
X_322_ clknet_2_1__leaf_clk _019_ net44 VGND VGND VPWR VPWR mask\[3\] _322_/a_1462_47#
+ _322_/a_543_47# _322_/a_651_413# _322_/a_193_47# _322_/a_805_47# _322_/a_448_47#
+ _322_/a_639_47# _322_/a_1283_21# _322_/a_761_289# _322_/a_1108_47# _322_/a_1217_47#
+ _322_/a_1270_413# _322_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_184_ net55 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__inv_2
X_253_ mask\[7\] _102_ _074_ VGND VGND VPWR VPWR _023_ _253_/a_384_47# _253_/a_81_21#
+ _253_/a_299_297# sky130_fd_sc_hd__a21o_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_167_ state\[1\] VGND VGND VPWR VPWR _051_ _167_/a_161_47# sky130_fd_sc_hd__buf_6
X_236_ _092_ _095_ VGND VGND VPWR VPWR _096_ _236_/a_109_297# sky130_fd_sc_hd__nor2_1
X_305_ clknet_2_1__leaf_clk _002_ net43 VGND VGND VPWR VPWR cal_itt\[2\] _305_/a_1462_47#
+ _305_/a_543_47# _305_/a_651_413# _305_/a_193_47# _305_/a_805_47# _305_/a_448_47#
+ _305_/a_639_47# _305_/a_1283_21# _305_/a_761_289# _305_/a_1108_47# _305_/a_1217_47#
+ _305_/a_1270_413# _305_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_219_ _074_ _083_ VGND VGND VPWR VPWR _008_ _219_/a_109_297# sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_11_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput38 net38 VGND VGND VPWR VPWR trimb[2] output38/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput27 net27 VGND VGND VPWR VPWR result[5] output27/a_27_47# sky130_fd_sc_hd__buf_2
Xoutput16 net16 VGND VGND VPWR VPWR ctlp[2] output16/a_27_47# sky130_fd_sc_hd__buf_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk clkbuf_0_clk/a_110_47# sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_183_ net35 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__inv_2
X_252_ net52 VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__inv_2
X_321_ clknet_2_1__leaf_clk _018_ net43 VGND VGND VPWR VPWR mask\[2\] _321_/a_1462_47#
+ _321_/a_543_47# _321_/a_651_413# _321_/a_193_47# _321_/a_805_47# _321_/a_448_47#
+ _321_/a_639_47# _321_/a_1283_21# _321_/a_761_289# _321_/a_1108_47# _321_/a_1217_47#
+ _321_/a_1270_413# _321_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_235_ net55 _094_ net54 VGND VGND VPWR VPWR _095_ _235_/a_382_297# _235_/a_297_47#
+ _235_/a_79_21# sky130_fd_sc_hd__o21a_1
X_304_ clknet_2_3__leaf_clk _001_ net47 VGND VGND VPWR VPWR cal_itt\[1\] _304_/a_1462_47#
+ _304_/a_543_47# _304_/a_651_413# _304_/a_193_47# _304_/a_805_47# _304_/a_448_47#
+ _304_/a_639_47# _304_/a_1283_21# _304_/a_761_289# _304_/a_1108_47# _304_/a_1217_47#
+ _304_/a_1270_413# _304_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_166_ state\[2\] VGND VGND VPWR VPWR _050_ _166_/a_161_47# sky130_fd_sc_hd__buf_6
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_149_ mask\[4\] net26 VGND VGND VPWR VPWR _043_ _149_/a_150_297# _149_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_218_ mask\[4\] _078_ net26 VGND VGND VPWR VPWR _083_ _218_/a_199_47# _218_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
Xoutput39 net39 VGND VGND VPWR VPWR trimb[3] output39/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput28 net28 VGND VGND VPWR VPWR result[6] output28/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput17 net17 VGND VGND VPWR VPWR ctlp[3] output17/a_27_47# sky130_fd_sc_hd__buf_2
XFILLER_0_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk clkbuf_2_0__f_clk/a_110_47#
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_182_ _058_ VGND VGND VPWR VPWR net35 _182_/a_27_47# sky130_fd_sc_hd__buf_1
X_251_ mask\[7\] net52 _101_ mask\[6\] VGND VGND VPWR VPWR _022_ _251_/a_27_297# _251_/a_109_47#
+ _251_/a_109_297# _251_/a_373_47# sky130_fd_sc_hd__a22o_1
X_320_ clknet_2_0__leaf_clk _017_ net44 VGND VGND VPWR VPWR mask\[1\] _320_/a_1462_47#
+ _320_/a_543_47# _320_/a_651_413# _320_/a_193_47# _320_/a_805_47# _320_/a_448_47#
+ _320_/a_639_47# _320_/a_1283_21# _320_/a_761_289# _320_/a_1108_47# _320_/a_1217_47#
+ _320_/a_1270_413# _320_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_165_ _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__inv_2
X_234_ mask\[0\] _049_ VGND VGND VPWR VPWR _094_ _234_/a_109_297# sky130_fd_sc_hd__nor2_1
X_303_ clknet_2_3__leaf_clk _000_ net47 VGND VGND VPWR VPWR cal_itt\[0\] _303_/a_1462_47#
+ _303_/a_543_47# _303_/a_651_413# _303_/a_193_47# _303_/a_805_47# _303_/a_448_47#
+ _303_/a_639_47# _303_/a_1283_21# _303_/a_761_289# _303_/a_1108_47# _303_/a_1217_47#
+ _303_/a_1270_413# _303_/a_27_47# sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_148_ net17 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__inv_2
X_217_ _074_ _082_ VGND VGND VPWR VPWR _007_ _217_/a_109_297# sky130_fd_sc_hd__nor2_1
Xoutput29 net29 VGND VGND VPWR VPWR result[7] output29/a_27_47# sky130_fd_sc_hd__buf_2
Xoutput18 net18 VGND VGND VPWR VPWR ctlp[4] output18/a_27_47# sky130_fd_sc_hd__buf_2
XFILLER_0_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_181_ trim_val\[4\] trim_mask\[4\] VGND VGND VPWR VPWR _058_ _181_/a_150_297# _181_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_250_ mask\[6\] net53 _101_ mask\[5\] VGND VGND VPWR VPWR _021_ _250_/a_27_297# _250_/a_109_47#
+ _250_/a_109_297# _250_/a_373_47# sky130_fd_sc_hd__a22o_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_164_ state\[0\] VGND VGND VPWR VPWR _048_ _164_/a_161_47# sky130_fd_sc_hd__buf_6
X_233_ calibrate _093_ _074_ net1 VGND VGND VPWR VPWR _012_ _233_/a_27_297# _233_/a_109_47#
+ _233_/a_109_297# _233_/a_373_47# sky130_fd_sc_hd__a22o_1
X_302_ cal_count\[3\] _066_ _136_ _092_ VGND VGND VPWR VPWR _038_ _302_/a_27_297#
+ _302_/a_109_47# _302_/a_109_297# _302_/a_373_47# sky130_fd_sc_hd__a22o_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_147_ _042_ VGND VGND VPWR VPWR net17 _147_/a_27_47# sky130_fd_sc_hd__buf_1
X_216_ mask\[3\] _078_ net25 VGND VGND VPWR VPWR _082_ _216_/a_199_47# _216_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput19 net19 VGND VGND VPWR VPWR ctlp[5] output19/a_27_47# sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_180_ net34 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__inv_2
Xfanout43 net45 VGND VGND VPWR VPWR net43 fanout43/a_27_47# sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_18_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_163_ net31 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__inv_2
X_232_ net54 _049_ _090_ _092_ VGND VGND VPWR VPWR _093_ _232_/a_114_297# _232_/a_304_297#
+ _232_/a_220_297# _232_/a_32_297# sky130_fd_sc_hd__or4_4
X_301_ _134_ _135_ VGND VGND VPWR VPWR _136_ _301_/a_129_47# _301_/a_47_47# _301_/a_285_47#
+ _301_/a_377_297# sky130_fd_sc_hd__xnor2_1
X_146_ mask\[3\] net25 VGND VGND VPWR VPWR _042_ _146_/a_150_297# _146_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_215_ _074_ _081_ VGND VGND VPWR VPWR _006_ _215_/a_109_297# sky130_fd_sc_hd__nor2_1
XFILLER_0_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout44 net45 VGND VGND VPWR VPWR net44 fanout44/a_27_47# sky130_fd_sc_hd__buf_2
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_162_ _047_ VGND VGND VPWR VPWR net31 _162_/a_27_47# sky130_fd_sc_hd__buf_1
X_231_ _091_ VGND VGND VPWR VPWR _092_ _231_/a_161_47# sky130_fd_sc_hd__buf_6
X_300_ cal_count\[3\] net2 VGND VGND VPWR VPWR _135_ _300_/a_129_47# _300_/a_47_47#
+ _300_/a_285_47# _300_/a_377_297# sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 cal VGND VGND VPWR VPWR net1 input1/a_75_212# sky130_fd_sc_hd__clkbuf_1
X_145_ net16 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__inv_2
X_214_ mask\[2\] _078_ net24 VGND VGND VPWR VPWR _081_ _214_/a_199_47# _214_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout45 net4 VGND VGND VPWR VPWR net45 fanout45/a_27_47# sky130_fd_sc_hd__buf_2
X_161_ trim_val\[0\] trim_mask\[0\] VGND VGND VPWR VPWR _047_ _161_/a_150_297# _161_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_230_ _053_ _063_ VGND VGND VPWR VPWR _091_ _230_/a_145_75# _230_/a_59_75# sky130_fd_sc_hd__and2_1
Xinput2 comp VGND VGND VPWR VPWR net2 input2/a_27_47# sky130_fd_sc_hd__clkbuf_2
X_144_ _041_ VGND VGND VPWR VPWR net16 _144_/a_27_47# sky130_fd_sc_hd__buf_1
X_213_ _074_ _080_ VGND VGND VPWR VPWR _005_ _213_/a_109_297# sky130_fd_sc_hd__nor2_1
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout46 net4 VGND VGND VPWR VPWR net46 fanout46/a_27_47# sky130_fd_sc_hd__clkbuf_4
X_160_ net21 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__inv_2
X_289_ net2 cal_count\[1\] VGND VGND VPWR VPWR _126_ _289_/a_150_297# _289_/a_68_297#
+ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 en VGND VGND VPWR VPWR net3 input3/a_75_212# sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_143_ mask\[2\] net24 VGND VGND VPWR VPWR _041_ _143_/a_150_297# _143_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_212_ mask\[1\] _078_ net23 VGND VGND VPWR VPWR _080_ _212_/a_199_47# _212_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout47 net4 VGND VGND VPWR VPWR net47 fanout47/a_27_47# sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_288_ net2 cal_count\[1\] VGND VGND VPWR VPWR _125_ _288_/a_145_75# _288_/a_59_75#
+ sky130_fd_sc_hd__and2_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk clkbuf_2_1__f_clk/a_110_47#
+ sky130_fd_sc_hd__clkbuf_16
Xinput4 rstn VGND VGND VPWR VPWR net4 input4/a_27_47# sky130_fd_sc_hd__buf_1
X_142_ net15 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__inv_2
X_211_ _074_ _079_ VGND VGND VPWR VPWR _004_ _211_/a_109_297# sky130_fd_sc_hd__nor2_1
XFILLER_0_22_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_287_ _124_ VGND VGND VPWR VPWR _035_ _287_/a_75_212# sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_141_ _040_ VGND VGND VPWR VPWR net15 _141_/a_27_47# sky130_fd_sc_hd__buf_1
X_210_ mask\[0\] _078_ net22 VGND VGND VPWR VPWR _079_ _210_/a_199_47# _210_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
X_339_ clknet_2_3__leaf_clk _036_ net47 VGND VGND VPWR VPWR cal_count\[1\] _339_/a_1140_413#
+ _339_/a_1296_47# _339_/a_1182_261# _339_/a_586_47# _339_/a_1602_47# _339_/a_956_413#
+ _339_/a_1224_47# _339_/a_193_47# _339_/a_796_47# _339_/a_381_47# _339_/a_1056_47#
+ _339_/a_1032_413# _339_/a_562_413# _339_/a_652_21# _339_/a_476_47# _339_/a_27_47#
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_147 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_286_ _122_ _123_ cal_count\[0\] VGND VGND VPWR VPWR _124_ _286_/a_505_21# _286_/a_535_374#
+ _286_/a_439_47# _286_/a_218_47# _286_/a_76_199# _286_/a_218_374# sky130_fd_sc_hd__mux2_1
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_140_ net23 mask\[1\] VGND VGND VPWR VPWR _040_ _140_/a_150_297# _140_/a_68_297#
+ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_269_ trim_mask\[1\] net49 trim_val\[1\] VGND VGND VPWR VPWR _112_ _269_/a_384_47#
+ _269_/a_81_21# _269_/a_299_297# sky130_fd_sc_hd__a21o_1
X_338_ clknet_2_3__leaf_clk _035_ net47 VGND VGND VPWR VPWR cal_count\[0\] _338_/a_1140_413#
+ _338_/a_1296_47# _338_/a_1182_261# _338_/a_586_47# _338_/a_1602_47# _338_/a_956_413#
+ _338_/a_1224_47# _338_/a_193_47# _338_/a_796_47# _338_/a_381_47# _338_/a_1056_47#
+ _338_/a_1032_413# _338_/a_562_413# _338_/a_652_21# _338_/a_476_47# _338_/a_27_47#
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_285_ _053_ _063_ VGND VGND VPWR VPWR _123_ _285_/a_113_47# sky130_fd_sc_hd__nand2_1
XFILLER_0_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_199_ _065_ _069_ _070_ VGND VGND VPWR VPWR _001_ _199_/a_193_297# _199_/a_109_297#
+ sky130_fd_sc_hd__nor3_1
X_268_ _111_ VGND VGND VPWR VPWR _029_ _268_/a_75_212# sky130_fd_sc_hd__clkbuf_1
X_337_ clknet_2_0__leaf_clk _034_ net44 VGND VGND VPWR VPWR en_co_clk _337_/a_1462_47#
+ _337_/a_543_47# _337_/a_651_413# _337_/a_193_47# _337_/a_805_47# _337_/a_448_47#
+ _337_/a_639_47# _337_/a_1283_21# _337_/a_761_289# _337_/a_1108_47# _337_/a_1217_47#
+ _337_/a_1270_413# _337_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_284_ _053_ _065_ VGND VGND VPWR VPWR _122_ _284_/a_150_297# _284_/a_68_297# sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_17_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_198_ cal_itt\[1\] cal_itt\[0\] _067_ VGND VGND VPWR VPWR _070_ _198_/a_181_47# _198_/a_109_47#
+ _198_/a_27_47# sky130_fd_sc_hd__and3_1
X_267_ _109_ _110_ VGND VGND VPWR VPWR _111_ _267_/a_145_75# _267_/a_59_75# sky130_fd_sc_hd__and2_1
X_336_ clknet_2_2__leaf_clk _033_ net46 VGND VGND VPWR VPWR trim_val\[4\] _336_/a_1462_47#
+ _336_/a_543_47# _336_/a_651_413# _336_/a_193_47# _336_/a_805_47# _336_/a_448_47#
+ _336_/a_639_47# _336_/a_1283_21# _336_/a_761_289# _336_/a_1108_47# _336_/a_1217_47#
+ _336_/a_1270_413# _336_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_319_ clknet_2_0__leaf_clk _016_ net43 VGND VGND VPWR VPWR mask\[0\] _319_/a_1462_47#
+ _319_/a_543_47# _319_/a_651_413# _319_/a_193_47# _319_/a_805_47# _319_/a_448_47#
+ _319_/a_639_47# _319_/a_1283_21# _319_/a_761_289# _319_/a_1108_47# _319_/a_1217_47#
+ _319_/a_1270_413# _319_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_283_ _121_ VGND VGND VPWR VPWR _034_ _283_/a_75_212# sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_197_ cal_itt\[0\] _067_ cal_itt\[1\] VGND VGND VPWR VPWR _069_ _197_/a_199_47# _197_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
X_266_ _048_ _106_ VGND VGND VPWR VPWR _110_ _266_/a_150_297# _266_/a_68_297# sky130_fd_sc_hd__or2_1
X_335_ clknet_2_2__leaf_clk _032_ net46 VGND VGND VPWR VPWR trim_val\[3\] _335_/a_1462_47#
+ _335_/a_543_47# _335_/a_651_413# _335_/a_193_47# _335_/a_805_47# _335_/a_448_47#
+ _335_/a_639_47# _335_/a_1283_21# _335_/a_761_289# _335_/a_1108_47# _335_/a_1217_47#
+ _335_/a_1270_413# _335_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_249_ mask\[5\] net53 _101_ mask\[4\] VGND VGND VPWR VPWR _020_ _249_/a_27_297# _249_/a_109_47#
+ _249_/a_109_297# _249_/a_373_47# sky130_fd_sc_hd__a22o_1
X_318_ clknet_2_0__leaf_clk _015_ net45 VGND VGND VPWR VPWR state\[2\] _318_/a_1462_47#
+ _318_/a_543_47# _318_/a_651_413# _318_/a_193_47# _318_/a_805_47# _318_/a_448_47#
+ _318_/a_639_47# _318_/a_1283_21# _318_/a_761_289# _318_/a_1108_47# _318_/a_1217_47#
+ _318_/a_1270_413# _318_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_282_ _065_ _120_ VGND VGND VPWR VPWR _121_ _282_/a_150_297# _282_/a_68_297# sky130_fd_sc_hd__or2_1
X_334_ clknet_2_2__leaf_clk _031_ net46 VGND VGND VPWR VPWR trim_val\[2\] _334_/a_1462_47#
+ _334_/a_543_47# _334_/a_651_413# _334_/a_193_47# _334_/a_805_47# _334_/a_448_47#
+ _334_/a_639_47# _334_/a_1283_21# _334_/a_761_289# _334_/a_1108_47# _334_/a_1217_47#
+ _334_/a_1270_413# _334_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_196_ _068_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
X_265_ trim_mask\[0\] _108_ trim_val\[0\] VGND VGND VPWR VPWR _109_ _265_/a_384_47#
+ _265_/a_81_21# _265_/a_299_297# sky130_fd_sc_hd__a21o_1
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_179_ _057_ VGND VGND VPWR VPWR net34 _179_/a_27_47# sky130_fd_sc_hd__buf_1
X_248_ mask\[4\] net53 _101_ mask\[3\] VGND VGND VPWR VPWR _019_ _248_/a_27_297# _248_/a_109_47#
+ _248_/a_109_297# _248_/a_373_47# sky130_fd_sc_hd__a22o_1
X_317_ clknet_2_0__leaf_clk _014_ net45 VGND VGND VPWR VPWR state\[1\] _317_/a_1462_47#
+ _317_/a_543_47# _317_/a_651_413# _317_/a_193_47# _317_/a_805_47# _317_/a_448_47#
+ _317_/a_639_47# _317_/a_1283_21# _317_/a_761_289# _317_/a_1108_47# _317_/a_1217_47#
+ _317_/a_1270_413# _317_/a_27_47# sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk clkbuf_2_2__f_clk/a_110_47#
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_281_ _090_ _092_ _095_ en_co_clk VGND VGND VPWR VPWR _120_ _281_/a_103_199# _281_/a_253_47#
+ _281_/a_337_297# _281_/a_253_297# sky130_fd_sc_hd__o31a_1
XFILLER_0_11_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ _062_ _067_ cal_itt\[0\] VGND VGND VPWR VPWR _068_ _195_/a_505_21# _195_/a_535_374#
+ _195_/a_439_47# _195_/a_218_47# _195_/a_76_199# _195_/a_218_374# sky130_fd_sc_hd__mux2_1
X_264_ _106_ _107_ VGND VGND VPWR VPWR _108_ _264_/a_27_297# sky130_fd_sc_hd__nor2_4
X_333_ clknet_2_2__leaf_clk _030_ net46 VGND VGND VPWR VPWR trim_val\[1\] _333_/a_1462_47#
+ _333_/a_543_47# _333_/a_651_413# _333_/a_193_47# _333_/a_805_47# _333_/a_448_47#
+ _333_/a_639_47# _333_/a_1283_21# _333_/a_761_289# _333_/a_1108_47# _333_/a_1217_47#
+ _333_/a_1270_413# _333_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_247_ mask\[3\] net52 _101_ mask\[2\] VGND VGND VPWR VPWR _018_ _247_/a_27_297# _247_/a_109_47#
+ _247_/a_109_297# _247_/a_373_47# sky130_fd_sc_hd__a22o_1
X_316_ clknet_2_0__leaf_clk _013_ net45 VGND VGND VPWR VPWR state\[0\] _316_/a_1462_47#
+ _316_/a_543_47# _316_/a_651_413# _316_/a_193_47# _316_/a_805_47# _316_/a_448_47#
+ _316_/a_639_47# _316_/a_1283_21# _316_/a_761_289# _316_/a_1108_47# _316_/a_1217_47#
+ _316_/a_1270_413# _316_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_178_ trim_val\[3\] trim_mask\[3\] VGND VGND VPWR VPWR _057_ _178_/a_150_297# _178_/a_68_297#
+ sky130_fd_sc_hd__or2_1
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_280_ _119_ VGND VGND VPWR VPWR _033_ _280_/a_75_212# sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ trim_mask\[0\] _064_ _066_ VGND VGND VPWR VPWR _067_ _194_/a_199_47# _194_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
X_263_ net54 _059_ _048_ VGND VGND VPWR VPWR _107_ _263_/a_382_297# _263_/a_297_47#
+ _263_/a_79_21# sky130_fd_sc_hd__o21a_1
X_332_ clknet_2_2__leaf_clk _029_ net46 VGND VGND VPWR VPWR trim_val\[0\] _332_/a_1462_47#
+ _332_/a_543_47# _332_/a_651_413# _332_/a_193_47# _332_/a_805_47# _332_/a_448_47#
+ _332_/a_639_47# _332_/a_1283_21# _332_/a_761_289# _332_/a_1108_47# _332_/a_1217_47#
+ _332_/a_1270_413# _332_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_22_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_177_ net33 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__inv_2
X_246_ mask\[2\] net52 _101_ mask\[1\] VGND VGND VPWR VPWR _017_ _246_/a_27_297# _246_/a_109_47#
+ _246_/a_109_297# _246_/a_373_47# sky130_fd_sc_hd__a22o_1
X_315_ clknet_2_0__leaf_clk _012_ net45 VGND VGND VPWR VPWR calibrate _315_/a_1462_47#
+ _315_/a_543_47# _315_/a_651_413# _315_/a_193_47# _315_/a_805_47# _315_/a_448_47#
+ _315_/a_639_47# _315_/a_1283_21# _315_/a_761_289# _315_/a_1108_47# _315_/a_1217_47#
+ _315_/a_1270_413# _315_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_229_ _087_ _089_ VGND VGND VPWR VPWR _090_ _229_/a_27_297# sky130_fd_sc_hd__nor2_2
XFILLER_0_18_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_193_ _053_ _065_ VGND VGND VPWR VPWR _066_ _193_/a_109_297# sky130_fd_sc_hd__nor2_1
X_262_ _053_ _063_ _105_ net55 net42 VGND VGND VPWR VPWR _106_ _262_/a_193_297# _262_/a_465_47#
+ _262_/a_205_47# _262_/a_109_297# _262_/a_27_47# sky130_fd_sc_hd__a221o_1
X_331_ clknet_2_2__leaf_clk _028_ net45 VGND VGND VPWR VPWR trim_mask\[4\] _331_/a_1462_47#
+ _331_/a_543_47# _331_/a_651_413# _331_/a_193_47# _331_/a_805_47# _331_/a_448_47#
+ _331_/a_639_47# _331_/a_1283_21# _331_/a_761_289# _331_/a_1108_47# _331_/a_1217_47#
+ _331_/a_1270_413# _331_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_176_ _056_ VGND VGND VPWR VPWR net33 _176_/a_27_47# sky130_fd_sc_hd__buf_1
X_245_ mask\[1\] net52 _101_ mask\[0\] VGND VGND VPWR VPWR _016_ _245_/a_27_297# _245_/a_109_47#
+ _245_/a_109_297# _245_/a_373_47# sky130_fd_sc_hd__a22o_1
X_314_ clknet_2_1__leaf_clk _011_ net43 VGND VGND VPWR VPWR net29 _314_/a_1462_47#
+ _314_/a_543_47# _314_/a_651_413# _314_/a_193_47# _314_/a_805_47# _314_/a_448_47#
+ _314_/a_639_47# _314_/a_1283_21# _314_/a_761_289# _314_/a_1108_47# _314_/a_1217_47#
+ _314_/a_1270_413# _314_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_159_ _046_ VGND VGND VPWR VPWR net21 _159_/a_27_47# sky130_fd_sc_hd__buf_1
X_228_ _052_ _088_ _048_ VGND VGND VPWR VPWR _089_ _228_/a_382_297# _228_/a_297_47#
+ _228_/a_79_21# sky130_fd_sc_hd__o21a_1
Xclone1 state\[2\] VGND VGND VPWR VPWR net55 clone1/a_27_47# sky130_fd_sc_hd__buf_2
XFILLER_0_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_192_ net54 _050_ _048_ net3 VGND VGND VPWR VPWR _065_ _192_/a_548_47# _192_/a_639_47#
+ _192_/a_476_47# _192_/a_174_21# _192_/a_505_280# _192_/a_27_47# sky130_fd_sc_hd__and4bb_2
X_261_ _048_ cal_count\[3\] VGND VGND VPWR VPWR _105_ _261_/a_113_47# sky130_fd_sc_hd__nand2_1
X_330_ clknet_2_2__leaf_clk _027_ net46 VGND VGND VPWR VPWR trim_mask\[3\] _330_/a_1462_47#
+ _330_/a_543_47# _330_/a_651_413# _330_/a_193_47# _330_/a_805_47# _330_/a_448_47#
+ _330_/a_639_47# _330_/a_1283_21# _330_/a_761_289# _330_/a_1108_47# _330_/a_1217_47#
+ _330_/a_1270_413# _330_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_175_ trim_val\[2\] trim_mask\[2\] VGND VGND VPWR VPWR _056_ _175_/a_150_297# _175_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_244_ _065_ net51 VGND VGND VPWR VPWR _101_ _244_/a_27_297# sky130_fd_sc_hd__nor2_2
X_313_ clknet_2_1__leaf_clk _010_ net43 VGND VGND VPWR VPWR net28 _313_/a_1462_47#
+ _313_/a_543_47# _313_/a_651_413# _313_/a_193_47# _313_/a_805_47# _313_/a_448_47#
+ _313_/a_639_47# _313_/a_1283_21# _313_/a_761_289# _313_/a_1108_47# _313_/a_1217_47#
+ _313_/a_1270_413# _313_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_158_ mask\[7\] net29 VGND VGND VPWR VPWR _046_ _158_/a_150_297# _158_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_227_ _051_ net55 trim_mask\[0\] VGND VGND VPWR VPWR _088_ _227_/a_109_93# _227_/a_368_53#
+ _227_/a_209_311# _227_/a_296_53# sky130_fd_sc_hd__and3b_1
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_75 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_260_ calibrate _049_ _052_ _104_ trim_mask\[4\] VGND VGND VPWR VPWR _028_ _260_/a_256_47#
+ _260_/a_584_47# _260_/a_93_21# _260_/a_250_297# _260_/a_346_47# sky130_fd_sc_hd__a32o_1
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_191_ _062_ _063_ VGND VGND VPWR VPWR _064_ _191_/a_27_297# sky130_fd_sc_hd__nor2_2
X_174_ net32 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__inv_2
X_243_ net55 _060_ _096_ _100_ VGND VGND VPWR VPWR _015_ _243_/a_27_297# _243_/a_109_47#
+ _243_/a_109_297# _243_/a_373_47# sky130_fd_sc_hd__a22o_1
X_312_ clknet_2_1__leaf_clk _009_ net44 VGND VGND VPWR VPWR net27 _312_/a_1462_47#
+ _312_/a_543_47# _312_/a_651_413# _312_/a_193_47# _312_/a_805_47# _312_/a_448_47#
+ _312_/a_639_47# _312_/a_1283_21# _312_/a_761_289# _312_/a_1108_47# _312_/a_1217_47#
+ _312_/a_1270_413# _312_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire42 _098_ VGND VGND VPWR VPWR net42 wire42/a_75_212# sky130_fd_sc_hd__clkbuf_1
X_157_ net20 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__inv_2
X_226_ net3 _062_ _075_ _060_ VGND VGND VPWR VPWR _087_ _226_/a_109_47# _226_/a_197_47#
+ _226_/a_303_47# _226_/a_27_47# sky130_fd_sc_hd__and4_1
XFILLER_0_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_209_ _077_ VGND VGND VPWR VPWR _078_ _209_/a_27_47# sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_13_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_190_ cal_itt\[3\] cal_itt\[2\] cal_itt\[1\] cal_itt\[0\] VGND VGND VPWR VPWR _063_
+ _190_/a_655_47# _190_/a_465_47# _190_/a_215_47# _190_/a_27_47# sky130_fd_sc_hd__nand4b_2
X_173_ _055_ VGND VGND VPWR VPWR net32 _173_/a_27_47# sky130_fd_sc_hd__buf_1
X_242_ calibrate _048_ _052_ VGND VGND VPWR VPWR _100_ _242_/a_382_297# _242_/a_297_47#
+ _242_/a_79_21# sky130_fd_sc_hd__o21a_1
X_311_ clknet_2_1__leaf_clk _008_ net44 VGND VGND VPWR VPWR net26 _311_/a_1462_47#
+ _311_/a_543_47# _311_/a_651_413# _311_/a_193_47# _311_/a_805_47# _311_/a_448_47#
+ _311_/a_639_47# _311_/a_1283_21# _311_/a_761_289# _311_/a_1108_47# _311_/a_1217_47#
+ _311_/a_1270_413# _311_/a_27_47# sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_1_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_156_ _045_ VGND VGND VPWR VPWR net20 _156_/a_27_47# sky130_fd_sc_hd__buf_1
X_225_ _074_ _086_ VGND VGND VPWR VPWR _011_ _225_/a_109_297# sky130_fd_sc_hd__nor2_1
X_139_ net14 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__inv_2
X_208_ _065_ net2 _076_ VGND VGND VPWR VPWR _077_ _208_/a_505_21# _208_/a_535_374#
+ _208_/a_439_47# _208_/a_218_47# _208_/a_76_199# _208_/a_218_374# sky130_fd_sc_hd__mux2_1
XFILLER_0_0_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk clkbuf_2_3__f_clk/a_110_47#
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_310_ clknet_2_1__leaf_clk _007_ net43 VGND VGND VPWR VPWR net25 _310_/a_1462_47#
+ _310_/a_543_47# _310_/a_651_413# _310_/a_193_47# _310_/a_805_47# _310_/a_448_47#
+ _310_/a_639_47# _310_/a_1283_21# _310_/a_761_289# _310_/a_1108_47# _310_/a_1217_47#
+ _310_/a_1270_413# _310_/a_27_47# sky130_fd_sc_hd__dfrtp_1
X_172_ trim_val\[1\] trim_mask\[1\] VGND VGND VPWR VPWR _055_ _172_/a_150_297# _172_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_241_ _092_ _099_ _095_ VGND VGND VPWR VPWR _014_ _241_/a_388_297# _241_/a_297_47#
+ _241_/a_105_352# sky130_fd_sc_hd__o21bai_1
XFILLER_0_2_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_155_ mask\[6\] net28 VGND VGND VPWR VPWR _045_ _155_/a_150_297# _155_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_224_ mask\[7\] _078_ net29 VGND VGND VPWR VPWR _086_ _224_/a_199_47# _224_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
X_138_ _039_ VGND VGND VPWR VPWR net14 _138_/a_27_47# sky130_fd_sc_hd__buf_1
X_207_ _075_ _049_ VGND VGND VPWR VPWR _076_ _207_/a_109_297# sky130_fd_sc_hd__nor2_1
XFILLER_0_20_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_171_ _054_ VGND VGND VPWR VPWR net30 _171_/a_27_47# sky130_fd_sc_hd__clkbuf_2
X_240_ _087_ _098_ VGND VGND VPWR VPWR _099_ _240_/a_109_297# sky130_fd_sc_hd__nor2_1
XFILLER_0_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer1 _108_ VGND VGND VPWR VPWR net48 rebuffer1/a_75_212# sky130_fd_sc_hd__clkbuf_1
X_223_ _074_ _085_ VGND VGND VPWR VPWR _010_ _223_/a_109_297# sky130_fd_sc_hd__nor2_1
X_154_ net19 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__inv_2
X_137_ net22 mask\[0\] VGND VGND VPWR VPWR _039_ _137_/a_150_297# _137_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_206_ _050_ _051_ VGND VGND VPWR VPWR _075_ _206_/a_27_93# _206_/a_206_47# sky130_fd_sc_hd__nand2b_1
X_170_ _049_ _052_ _053_ VGND VGND VPWR VPWR _054_ _170_/a_384_47# _170_/a_81_21#
+ _170_/a_299_297# sky130_fd_sc_hd__a21o_1
X_299_ _129_ _130_ _131_ VGND VGND VPWR VPWR _134_ _299_/a_215_297# _299_/a_27_413#
+ _299_/a_298_297# _299_/a_382_47# sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer2 _108_ VGND VGND VPWR VPWR net49 rebuffer2/a_75_212# sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_5_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_153_ _044_ VGND VGND VPWR VPWR net19 _153_/a_27_47# sky130_fd_sc_hd__buf_1
X_222_ mask\[6\] _078_ net28 VGND VGND VPWR VPWR _085_ _222_/a_199_47# _222_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
Xclone7 state\[1\] VGND VGND VPWR VPWR net54 clone7/a_27_47# sky130_fd_sc_hd__clkbuf_2
X_205_ _065_ VGND VGND VPWR VPWR _074_ _205_/a_27_47# sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_298_ cal_count\[2\] _122_ _133_ _123_ VGND VGND VPWR VPWR _037_ _298_/a_78_199#
+ _298_/a_493_297# _298_/a_215_47# _298_/a_292_297# sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_21_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer3 _108_ VGND VGND VPWR VPWR net50 rebuffer3/a_75_212# sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_152_ mask\[5\] net27 VGND VGND VPWR VPWR _044_ _152_/a_150_297# _152_/a_68_297#
+ sky130_fd_sc_hd__or2_1
X_221_ _074_ _084_ VGND VGND VPWR VPWR _009_ _221_/a_109_297# sky130_fd_sc_hd__nor2_1
X_204_ _073_ VGND VGND VPWR VPWR _003_ _204_/a_75_212# sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_297_ _129_ _132_ VGND VGND VPWR VPWR _133_ _297_/a_129_47# _297_/a_47_47# _297_/a_285_47#
+ _297_/a_377_297# sky130_fd_sc_hd__xnor2_1
Xrebuffer4 _076_ VGND VGND VPWR VPWR net51 rebuffer4/a_27_47# sky130_fd_sc_hd__buf_1
X_151_ net18 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__inv_2
X_220_ mask\[5\] _078_ net27 VGND VGND VPWR VPWR _084_ _220_/a_199_47# _220_/a_113_297#
+ sky130_fd_sc_hd__a21oi_1
X_203_ cal_itt\[3\] _072_ VGND VGND VPWR VPWR _073_ _203_/a_145_75# _203_/a_59_75#
+ sky130_fd_sc_hd__and2_1
XFILLER_0_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_296_ _130_ _131_ VGND VGND VPWR VPWR _132_ _296_/a_113_47# sky130_fd_sc_hd__nand2_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer5 net51 VGND VGND VPWR VPWR net52 rebuffer5/a_161_47# sky130_fd_sc_hd__buf_6
X_150_ _043_ VGND VGND VPWR VPWR net18 _150_/a_27_47# sky130_fd_sc_hd__buf_1
X_279_ trim_val\[4\] _118_ _108_ VGND VGND VPWR VPWR _119_ _279_/a_396_47# _279_/a_206_47#
+ _279_/a_490_47# _279_/a_314_297# _279_/a_204_297# _279_/a_27_47# sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_202_ cal_itt\[2\] _070_ _072_ VGND VGND VPWR VPWR _002_ _202_/a_382_297# _202_/a_297_47#
+ _202_/a_79_21# sky130_fd_sc_hd__o21a_1
XFILLER_0_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput40 net40 VGND VGND VPWR VPWR trimb[4] output40/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput5 net5 VGND VGND VPWR VPWR clkc output5/a_27_47# sky130_fd_sc_hd__buf_1
X_295_ net2 cal_count\[2\] VGND VGND VPWR VPWR _131_ _295_/a_113_47# sky130_fd_sc_hd__nand2_1
Xrebuffer6 _076_ VGND VGND VPWR VPWR net53 rebuffer6/a_27_47# sky130_fd_sc_hd__buf_1
X_278_ _062_ net40 net30 VGND VGND VPWR VPWR _118_ _278_/a_109_297# _278_/a_27_47#
+ sky130_fd_sc_hd__o21ai_1
X_201_ _067_ _071_ VGND VGND VPWR VPWR _072_ _201_/a_113_47# sky130_fd_sc_hd__nand2_1
XFILLER_0_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput41 net41 VGND VGND VPWR VPWR valid output41/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput30 net30 VGND VGND VPWR VPWR sample output30/a_27_47# sky130_fd_sc_hd__clkbuf_4
Xoutput6 net6 VGND VGND VPWR VPWR ctln[0] output6/a_27_47# sky130_fd_sc_hd__buf_2
C0 _074_ _011_ 0.0529f
C1 VPWR _231_/a_161_47# 0.0566f
C2 _302_/a_27_297# net40 1.71e-19
C3 net50 _280_/a_75_212# 6.72e-19
C4 _290_/a_27_413# _127_ 6.21e-19
C5 ctlp[1] net29 5.91e-19
C6 net16 _112_ 0.0667f
C7 _272_/a_299_297# net16 0.00392f
C8 _089_ _090_ 0.0252f
C9 _313_/a_27_47# _085_ 0.00843f
C10 _026_ trim_mask\[3\] 0.00642f
C11 VPWR trim_mask\[3\] 0.219f
C12 net43 _019_ 6.48e-19
C13 net21 _312_/a_27_47# 2.25e-21
C14 _170_/a_384_47# _049_ 0.0013f
C15 _170_/a_81_21# _054_ 0.00672f
C16 _323_/a_543_47# mask\[4\] 8.93e-19
C17 _024_ _053_ 5.87e-20
C18 net12 _208_/a_76_199# 0.0113f
C19 net30 _170_/a_81_21# 2.4e-19
C20 _187_/a_27_413# clkc 3.36e-19
C21 _239_/a_27_297# _049_ 0.012f
C22 net50 _257_/a_373_47# 1.65e-19
C23 _303_/a_805_47# net19 6.71e-19
C24 _337_/a_1217_47# en_co_clk 3.92e-19
C25 calibrate state\[1\] 0.00217f
C26 _012_ net45 1.38e-19
C27 cal_count\[1\] _036_ 2.79e-20
C28 VPWR _107_ 0.786f
C29 _312_/a_27_47# _312_/a_1283_21# -9.15e-20
C30 _033_ _330_/a_448_47# 6.61e-19
C31 _336_/a_1108_47# net46 -0.0141f
C32 _328_/a_1283_21# trim_mask\[1\] 0.0273f
C33 _341_/a_1283_21# _058_ 1.27e-20
C34 _051_ en_co_clk 0.00346f
C35 VPWR _001_ 1.42f
C36 _320_/a_27_47# _246_/a_27_297# 2.32e-20
C37 _188_/a_27_47# _061_ 0.0308f
C38 net1 _316_/a_448_47# 1.29e-20
C39 VPWR _333_/a_1108_47# 0.00663f
C40 VPWR _166_/a_161_47# 0.104f
C41 _149_/a_68_297# _311_/a_27_47# 1.72e-21
C42 _092_ net18 4.21e-19
C43 _290_/a_27_413# _126_ 0.00183f
C44 _128_ _291_/a_117_297# 7.95e-21
C45 _309_/a_193_47# _216_/a_113_297# 4.52e-20
C46 _200_/a_209_297# cal_itt\[1\] 0.00592f
C47 net44 _208_/a_76_199# 2.12e-20
C48 _168_/a_207_413# _227_/a_209_311# 3.67e-21
C49 _325_/a_1270_413# net13 1.29e-19
C50 cal_count\[0\] net33 0.00507f
C51 _063_ net19 0.824f
C52 _231_/a_161_47# _063_ 0.00133f
C53 mask\[6\] _021_ 0.017f
C54 _049_ _203_/a_59_75# 7.54e-22
C55 trim_mask\[0\] net40 0.00625f
C56 _022_ net26 8.91e-20
C57 result[1] clknet_2_0__leaf_clk 0.0172f
C58 _237_/a_505_21# _099_ 0.0337f
C59 _237_/a_76_199# _092_ 0.0622f
C60 _323_/a_543_47# _020_ 1.98e-19
C61 _192_/a_27_47# _049_ 0.00826f
C62 _048_ _089_ 0.164f
C63 VPWR _155_/a_68_297# 0.0185f
C64 _322_/a_193_47# _205_/a_27_47# 0.0108f
C65 _208_/a_76_199# _003_ 4.11e-20
C66 _104_ trim_mask\[2\] 0.479f
C67 mask\[1\] net14 0.00984f
C68 VPWR _279_/a_27_47# 0.0371f
C69 _331_/a_1462_47# _028_ 2.52e-19
C70 _061_ net33 0.0164f
C71 en_co_clk _316_/a_1283_21# 3.25e-21
C72 _028_ _260_/a_93_21# 0.00127f
C73 clknet_2_2__leaf_clk _260_/a_250_297# 1.54e-21
C74 _327_/a_761_289# clknet_2_3__leaf_clk 3e-20
C75 _256_/a_27_297# net46 7.71e-19
C76 _101_ _209_/a_27_47# 0.0126f
C77 VPWR _325_/a_1108_47# 0.0223f
C78 net13 _095_ 0.00928f
C79 net12 _059_ 4.92e-20
C80 net4 _330_/a_1283_21# 4.47e-19
C81 _255_/a_27_47# _227_/a_109_93# 2.21e-19
C82 result[2] clknet_2_1__leaf_clk 2.89e-20
C83 _107_ _063_ 0.019f
C84 trim_mask\[0\] _267_/a_145_75# 0.0029f
C85 _040_ _248_/a_109_297# 4.45e-20
C86 _002_ cal_itt\[3\] 1.29e-19
C87 fanout46/a_27_47# _336_/a_1283_21# 0.0114f
C88 _325_/a_27_47# _046_ 7.78e-20
C89 net15 _282_/a_68_297# 0.00169f
C90 _104_ _329_/a_27_47# 1.59e-19
C91 _340_/a_1032_413# net37 9.31e-37
C92 _064_ clkbuf_2_3__f_clk/a_110_47# 0.0533f
C93 _094_ _337_/a_448_47# 0.025f
C94 _327_/a_639_47# net18 6.77e-19
C95 VPWR _181_/a_68_297# 0.00971f
C96 _214_/a_199_47# mask\[2\] 0.00137f
C97 mask\[1\] _040_ 0.41f
C98 _051_ _235_/a_297_47# 1.85e-20
C99 _036_ _001_ 0.00281f
C100 net10 trim_val\[3\] 5.28e-22
C101 VPWR _248_/a_109_297# 0.00318f
C102 _306_/a_448_47# clk 7.3e-22
C103 _185_/a_68_297# net41 0.0201f
C104 _121_ _120_ 0.00162f
C105 net12 _306_/a_1108_47# 0.00227f
C106 _059_ net44 0.00165f
C107 trim_val\[3\] clknet_2_2__leaf_clk 0.00266f
C108 _080_ _016_ 8.64e-21
C109 _033_ _027_ 2.18e-19
C110 _103_ _254_/a_109_297# 9.83e-19
C111 _255_/a_27_47# net42 5.16e-19
C112 _320_/a_761_289# mask\[2\] 1.96e-19
C113 net1 _013_ 0.00186f
C114 VPWR mask\[1\] 2.13f
C115 _068_ _067_ 0.0116f
C116 cal_itt\[2\] cal_itt\[3\] 0.00647f
C117 _068_ _070_ 0.0108f
C118 _253_/a_81_21# _310_/a_193_47# 0.00844f
C119 _053_ clkbuf_2_3__f_clk/a_110_47# 0.133f
C120 _107_ _260_/a_346_47# 2.81e-19
C121 VPWR _185_/a_68_297# 0.0255f
C122 result[7] _078_ 2.78e-20
C123 _309_/a_651_413# net25 1.1e-19
C124 net12 _075_ 0.057f
C125 _303_/a_761_289# mask\[4\] 5.88e-19
C126 _078_ net30 0.0868f
C127 clkbuf_2_1__f_clk/a_110_47# _319_/a_651_413# 9.92e-19
C128 clknet_2_1__leaf_clk _319_/a_193_47# 8.29e-19
C129 comp _129_ 0.00337f
C130 clknet_2_0__leaf_clk _049_ 0.221f
C131 _063_ _279_/a_27_47# 3.67e-19
C132 _318_/a_27_47# net45 2.94e-19
C133 _325_/a_651_413# _101_ 2.38e-19
C134 _325_/a_1108_47# net52 2.36e-21
C135 _216_/a_199_47# _101_ 1.55e-20
C136 mask\[3\] _245_/a_373_47# 7.06e-20
C137 _306_/a_1108_47# net44 0.0124f
C138 input3/a_75_212# en 0.0154f
C139 _326_/a_193_47# _023_ 0.0414f
C140 _326_/a_761_289# _102_ 1.46e-19
C141 _326_/a_543_47# mask\[7\] 0.00755f
C142 cal_itt\[2\] _262_/a_205_47# 3.12e-20
C143 trim_mask\[3\] net50 0.0656f
C144 clkbuf_2_0__f_clk/a_110_47# net55 6.68e-20
C145 _293_/a_81_21# net2 5.27e-19
C146 clkbuf_2_2__f_clk/a_110_47# _330_/a_1108_47# 0.00167f
C147 _286_/a_76_199# _338_/a_193_47# 0.00114f
C148 _324_/a_27_47# mask\[5\] 2.42e-19
C149 _255_/a_27_47# net30 0.00224f
C150 _340_/a_476_47# cal_count\[0\] 7.26e-21
C151 net23 mask\[1\] 0.831f
C152 net22 _078_ 0.0116f
C153 net50 _107_ 4.2e-20
C154 net44 _075_ 0.0155f
C155 clk _088_ 8.97e-20
C156 _187_/a_27_413# _136_ 1.29e-19
C157 _210_/a_199_47# net45 1.19e-19
C158 _248_/a_373_47# _101_ 2.72e-19
C159 _340_/a_27_47# net2 1.21e-19
C160 VPWR _118_ 0.138f
C161 _088_ clone7/a_27_47# 6.68e-21
C162 VPWR _327_/a_1283_21# 0.0136f
C163 _306_/a_1108_47# _003_ 5.47e-21
C164 _317_/a_639_47# _014_ 9.32e-19
C165 _317_/a_1108_47# state\[1\] 9.14e-19
C166 _317_/a_1270_413# net45 -3.58e-20
C167 _136_ _332_/a_27_47# 0.00475f
C168 trim_mask\[2\] _267_/a_59_75# 3.93e-21
C169 _136_ _268_/a_75_212# 0.0029f
C170 _074_ _313_/a_761_289# 2.01e-20
C171 _232_/a_32_297# _100_ 1.42e-20
C172 _315_/a_27_47# _315_/a_1108_47# -2.98e-20
C173 net4 _195_/a_218_374# 7.36e-19
C174 output27/a_27_47# output28/a_27_47# 0.00249f
C175 output16/a_27_47# output39/a_27_47# 8.52e-19
C176 _167_/a_161_47# calibrate 1.95e-20
C177 _322_/a_1270_413# mask\[3\] 3.62e-19
C178 mask\[1\] net52 0.0404f
C179 _058_ _119_ 4.32e-19
C180 _259_/a_109_297# _119_ 1.16e-20
C181 net2 _144_/a_27_47# 6.55e-20
C182 _064_ cal_count\[3\] 0.297f
C183 _110_ _336_/a_1108_47# 0.0126f
C184 net13 state\[0\] 0.143f
C185 _097_ net45 0.235f
C186 _312_/a_27_47# _045_ 6.75e-19
C187 _249_/a_27_297# _312_/a_193_47# 2.91e-21
C188 _064_ _257_/a_27_297# 0.025f
C189 net19 _279_/a_396_47# 0.0147f
C190 _320_/a_1108_47# _077_ 2.9e-19
C191 _265_/a_81_21# _109_ 0.0132f
C192 ctlp[3] ctlp[4] 0.00165f
C193 _074_ _143_/a_68_297# 2.68e-20
C194 _309_/a_27_47# mask\[2\] 7.45e-21
C195 clk _108_ 2.39e-21
C196 net48 _056_ 0.0137f
C197 trim_val\[2\] net33 0.00704f
C198 _334_/a_1283_21# net34 0.0166f
C199 trim_mask\[1\] _066_ 1.32e-21
C200 mask\[7\] _310_/a_1108_47# 1.79e-19
C201 _102_ _310_/a_1283_21# 4.63e-19
C202 _023_ _310_/a_543_47# 7.13e-19
C203 _149_/a_150_297# net26 1.05e-19
C204 _053_ cal_count\[3\] 0.0162f
C205 VPWR _281_/a_337_297# -4.67e-19
C206 _192_/a_548_47# _065_ 1.74e-20
C207 net45 _315_/a_543_47# 6.61e-20
C208 clknet_2_0__leaf_clk _315_/a_1108_47# 0.016f
C209 _014_ _315_/a_1283_21# 6.06e-19
C210 _071_ _065_ 6.44e-20
C211 _090_ _092_ 0.0602f
C212 _218_/a_113_297# mask\[4\] 0.00258f
C213 VPWR _288_/a_145_75# -1.44e-19
C214 _103_ _262_/a_27_47# 2.31e-19
C215 net16 net33 0.11f
C216 _063_ _118_ 0.00299f
C217 net8 _114_ 3.77e-19
C218 _107_ _279_/a_396_47# 0.0111f
C219 _058_ _266_/a_150_297# 4.73e-20
C220 _321_/a_543_47# clknet_2_1__leaf_clk 0.0142f
C221 output32/a_27_47# net34 0.0191f
C222 _336_/a_27_47# net30 6.14e-21
C223 net4 _108_ 0.0253f
C224 _004_ net30 0.125f
C225 ctln[1] clk 0.00132f
C226 _286_/a_439_47# _122_ 5.37e-22
C227 _340_/a_27_47# _123_ 0.519f
C228 clone1/a_27_47# _049_ 0.0108f
C229 net54 _089_ 4.07e-20
C230 _253_/a_81_21# _224_/a_113_297# 1.29e-21
C231 _060_ _087_ 6.92e-19
C232 cal_count\[0\] _338_/a_193_47# 8.11e-20
C233 _124_ _338_/a_476_47# 0.00285f
C234 _242_/a_297_47# _099_ 4.21e-19
C235 _324_/a_1217_47# mask\[5\] 1.52e-19
C236 VPWR output19/a_27_47# 0.0697f
C237 _262_/a_27_47# _105_ 0.0527f
C238 _168_/a_27_413# _336_/a_27_47# 4.62e-21
C239 _110_ _162_/a_27_47# 9.22e-20
C240 _033_ _032_ 5.83e-21
C241 _322_/a_761_289# mask\[2\] 1.89e-19
C242 _055_ _108_ 0.00609f
C243 _004_ net22 0.00877f
C244 _079_ _078_ 0.0126f
C245 ctln[1] net4 0.0343f
C246 clknet_2_0__leaf_clk state\[1\] 0.027f
C247 net9 _304_/a_193_47# 0.0014f
C248 output14/a_27_47# net14 0.00571f
C249 trim[0] _055_ 0.0624f
C250 net31 net34 0.966f
C251 comp _297_/a_47_47# 1.17e-19
C252 _122_ _108_ 4.53e-21
C253 _301_/a_47_47# _332_/a_761_289# 2.67e-19
C254 ctln[2] ctln[3] 0.00303f
C255 trim_mask\[4\] _279_/a_490_47# 9.91e-21
C256 clknet_2_2__leaf_clk trim_val\[4\] 1.6e-19
C257 _327_/a_543_47# clknet_2_2__leaf_clk 0.00175f
C258 _060_ _263_/a_297_47# 0.00436f
C259 state\[2\] _090_ 3.14e-19
C260 _329_/a_193_47# net46 0.00137f
C261 VPWR _330_/a_761_289# 0.00452f
C262 _339_/a_193_47# _286_/a_505_21# 1.07e-19
C263 _048_ _092_ 0.273f
C264 _275_/a_299_297# _178_/a_68_297# 0.00615f
C265 _103_ wire42/a_75_212# 0.0649f
C266 _096_ net30 1.8e-20
C267 _323_/a_761_289# _068_ 1.5e-21
C268 output5/a_27_47# _131_ 0.00106f
C269 net3 _095_ 0.193f
C270 _337_/a_27_47# _049_ 0.0504f
C271 _259_/a_373_47# clknet_2_2__leaf_clk 3.54e-21
C272 cal_itt\[1\] _304_/a_1283_21# 0.00297f
C273 _331_/a_27_47# _330_/a_448_47# 3.88e-21
C274 _331_/a_448_47# _330_/a_27_47# 3.88e-21
C275 _189_/a_408_47# net12 4.34e-22
C276 trim_mask\[4\] _092_ 2.7e-22
C277 _181_/a_150_297# _279_/a_27_47# 1.25e-19
C278 net46 net18 0.0539f
C279 mask\[2\] _101_ 0.13f
C280 net50 _118_ 0.00284f
C281 state\[2\] _242_/a_382_297# 2.81e-19
C282 cal_count\[0\] output40/a_27_47# 3.06e-19
C283 mask\[0\] _319_/a_448_47# 0.0264f
C284 _105_ wire42/a_75_212# 8.03e-20
C285 _293_/a_299_297# _127_ 2.03e-20
C286 VPWR output14/a_27_47# 0.0741f
C287 _076_ net53 0.0273f
C288 _319_/a_543_47# clknet_2_0__leaf_clk 0.0375f
C289 _319_/a_193_47# net45 2.36e-19
C290 calibrate _240_/a_109_297# 1.7e-21
C291 _321_/a_805_47# _042_ 2.51e-19
C292 _307_/a_1108_47# _137_/a_68_297# 3.43e-19
C293 _286_/a_505_21# clknet_2_3__leaf_clk 0.0797f
C294 _305_/a_1108_47# net44 9.86e-21
C295 mask\[6\] _313_/a_27_47# 4.14e-19
C296 _200_/a_80_21# clkbuf_0_clk/a_110_47# 1.35e-20
C297 net5 output5/a_27_47# 0.0154f
C298 output11/a_27_47# net11 0.0201f
C299 net44 _311_/a_639_47# -3.61e-19
C300 net21 _084_ 1.92e-20
C301 net27 _312_/a_193_47# 1.15e-19
C302 _300_/a_47_47# _298_/a_215_47# 1.54e-20
C303 _273_/a_145_75# _031_ 6.16e-19
C304 trim_mask\[2\] fanout46/a_27_47# 0.00289f
C305 net2 net34 0.0237f
C306 _189_/a_408_47# net44 1.14e-20
C307 en_co_clk _087_ 1.01e-24
C308 cal_count\[0\] _338_/a_796_47# 2.06e-20
C309 VPWR _306_/a_1283_21# 0.0317f
C310 _327_/a_27_47# _109_ 2.68e-21
C311 _312_/a_1283_21# _084_ 1.03e-21
C312 _319_/a_193_47# _065_ 5.84e-19
C313 clkbuf_2_0__f_clk/a_110_47# _121_ 0.00357f
C314 _134_ _300_/a_47_47# 7.21e-19
C315 _301_/a_377_297# net2 7.35e-19
C316 _322_/a_1108_47# _077_ 5.29e-19
C317 cal_itt\[1\] _091_ 0.00111f
C318 rebuffer4/a_27_47# rebuffer6/a_27_47# 1.62e-19
C319 _176_/a_27_47# net33 0.00261f
C320 _241_/a_105_352# _099_ 0.00617f
C321 _341_/a_193_47# net2 9.68e-20
C322 _341_/a_1108_47# _300_/a_285_47# 8.66e-20
C323 state\[2\] _048_ 0.0104f
C324 _293_/a_299_297# _126_ 0.00805f
C325 _058_ _333_/a_639_47# 4.87e-19
C326 net31 _133_ 1.06e-20
C327 output33/a_27_47# _047_ 4.2e-22
C328 net2 _299_/a_298_297# 3.72e-20
C329 net35 trim_val\[0\] 0.138f
C330 VPWR _062_ 2.77f
C331 _262_/a_205_47# net55 3.16e-19
C332 _102_ _251_/a_109_297# 6.74e-19
C333 mask\[7\] _251_/a_109_47# 0.00419f
C334 net9 _340_/a_1182_261# 9.58e-19
C335 _041_ clknet_2_1__leaf_clk 0.0101f
C336 _319_/a_27_47# _319_/a_193_47# -0.325f
C337 state\[2\] trim_mask\[4\] 0.168f
C338 _079_ _004_ 0.0613f
C339 _102_ _042_ 1.59e-20
C340 _307_/a_543_47# _074_ 0.0152f
C341 _307_/a_761_289# calibrate 3.2e-20
C342 en_co_clk _263_/a_297_47# 8.37e-19
C343 _326_/a_543_47# net28 7.67e-20
C344 _325_/a_193_47# mask\[5\] 3.3e-20
C345 _002_ clk 5.38e-20
C346 _279_/a_396_47# _118_ 0.00755f
C347 _279_/a_204_297# trim_val\[4\] 3.12e-19
C348 _329_/a_1462_47# net46 5.11e-19
C349 _189_/a_27_47# _098_ 1.09e-19
C350 _339_/a_652_21# cal_count\[0\] 0.0264f
C351 _065_ _202_/a_79_21# 0.0512f
C352 ctlp[7] _078_ 5.41e-19
C353 _234_/a_109_297# _337_/a_193_47# 9.28e-20
C354 _304_/a_543_47# _065_ 0.00211f
C355 _337_/a_1217_47# _049_ 1.93e-19
C356 _317_/a_193_47# _316_/a_761_289# 1.78e-20
C357 _317_/a_27_47# _316_/a_543_47# 1.37e-20
C358 net43 _314_/a_761_289# 0.0102f
C359 _068_ clknet_2_3__leaf_clk 1.16e-19
C360 clk _317_/a_1283_21# 0.00588f
C361 VPWR _195_/a_76_199# 3.42e-19
C362 _331_/a_27_47# _027_ 4.98e-19
C363 clknet_2_2__leaf_clk _330_/a_193_47# 0.0438f
C364 _028_ _330_/a_27_47# 5.1e-19
C365 _190_/a_27_47# _092_ 3.77e-20
C366 _051_ _049_ 0.0328f
C367 trim_val\[1\] net34 0.00267f
C368 net49 _055_ 1.29e-20
C369 VPWR _326_/a_1283_21# 0.0848f
C370 _314_/a_805_47# net14 6.71e-19
C371 _051_ _318_/a_761_289# 4.03e-21
C372 _329_/a_1283_21# _031_ 0.00166f
C373 VPWR _334_/a_1283_21# 0.0334f
C374 _189_/a_27_47# clknet_0_clk 0.0512f
C375 _181_/a_150_297# _118_ 8.55e-19
C376 _306_/a_448_47# _101_ 8.21e-21
C377 clkbuf_2_1__f_clk/a_110_47# clknet_0_clk 0.0385f
C378 output25/a_27_47# _310_/a_27_47# 0.0112f
C379 _002_ net4 7.04e-21
C380 net21 _085_ 8.48e-20
C381 net15 _046_ 0.135f
C382 state\[0\] net3 0.135f
C383 net17 _042_ 0.0282f
C384 trimb[0] net33 0.00141f
C385 net9 trim_mask\[0\] 0.0947f
C386 _307_/a_1270_413# _039_ 3.69e-19
C387 VPWR _286_/a_535_374# -7.62e-19
C388 _340_/a_1182_261# _132_ 5.78e-20
C389 _330_/a_193_47# net11 3.59e-19
C390 _330_/a_543_47# net19 0.0116f
C391 cal_itt\[2\] clk 0.0131f
C392 _071_ clkbuf_0_clk/a_110_47# 0.0217f
C393 _256_/a_27_297# rebuffer3/a_75_212# 4.76e-21
C394 net4 _317_/a_1283_21# 0.0129f
C395 VPWR _137_/a_68_297# 0.0358f
C396 _303_/a_193_47# _068_ 0.00885f
C397 _274_/a_75_212# trim_mask\[1\] 1.93e-19
C398 output32/a_27_47# VPWR 0.141f
C399 _078_ _313_/a_543_47# 0.0015f
C400 net2 _133_ 0.00134f
C401 _300_/a_47_47# cal_count\[3\] 0.041f
C402 _012_ _013_ 1.91e-19
C403 _182_/a_27_47# _058_ 0.0149f
C404 _337_/a_543_47# net45 3.42e-20
C405 _063_ _062_ 0.251f
C406 _337_/a_1108_47# clknet_2_0__leaf_clk 7.25e-20
C407 VPWR _335_/a_761_289# 0.0079f
C408 net28 _314_/a_639_47# 0.00177f
C409 _323_/a_761_289# _042_ 0.0184f
C410 _309_/a_543_47# _310_/a_1108_47# 2.66e-20
C411 _237_/a_505_21# _093_ 4.38e-19
C412 _035_ _065_ 5.27e-20
C413 trim_mask\[3\] _330_/a_543_47# 5.37e-21
C414 _167_/a_161_47# clknet_2_0__leaf_clk 1.92e-20
C415 _309_/a_27_47# _074_ 0.0189f
C416 _015_ _185_/a_68_297# 0.00565f
C417 _326_/a_651_413# net43 0.00166f
C418 _319_/a_1462_47# _065_ 1.27e-19
C419 _257_/a_109_297# _335_/a_1108_47# 1.11e-20
C420 _323_/a_448_47# clknet_2_1__leaf_clk 1.99e-19
C421 VPWR _187_/a_212_413# -0.00205f
C422 net13 calibrate 0.00629f
C423 cal_itt\[2\] net4 1.64e-21
C424 VPWR _314_/a_805_47# 2.69e-19
C425 VPWR _332_/a_193_47# -0.292f
C426 _289_/a_68_297# _122_ 1.55e-19
C427 _228_/a_79_21# _242_/a_79_21# 0.0132f
C428 fanout43/a_27_47# _212_/a_113_297# 7.26e-19
C429 clk _318_/a_651_413# 0.0263f
C430 _104_ _050_ 0.0258f
C431 _337_/a_543_47# _065_ 1.69e-19
C432 _048_ _226_/a_197_47# 0.00231f
C433 _110_ _329_/a_193_47# 2.48e-19
C434 _143_/a_150_297# _078_ 0.00132f
C435 _195_/a_76_199# _063_ 5.74e-19
C436 net31 VPWR 1.09f
C437 _326_/a_1283_21# net52 0.0128f
C438 net9 _338_/a_652_21# 5.31e-20
C439 net23 _137_/a_68_297# 2.59e-19
C440 fanout45/a_27_47# net45 0.0324f
C441 net3 _226_/a_27_47# 0.00183f
C442 _336_/a_27_47# _336_/a_639_47# -0.0015f
C443 _102_ _022_ 1.9e-20
C444 _314_/a_1108_47# _046_ 3.69e-20
C445 result[1] _308_/a_761_289# 0.00102f
C446 _281_/a_103_199# _095_ 0.0669f
C447 _060_ _099_ 0.00621f
C448 net54 _092_ 0.204f
C449 _289_/a_68_297# _299_/a_27_413# 6.12e-19
C450 _249_/a_27_297# mask\[5\] 0.0277f
C451 _059_ _107_ 9.45e-19
C452 VPWR _310_/a_448_47# -0.00224f
C453 _306_/a_1108_47# net19 2.19e-21
C454 _110_ net18 0.0157f
C455 mask\[3\] mask\[5\] 7.12e-22
C456 _340_/a_1032_413# cal_count\[2\] 0.00921f
C457 clknet_0_clk _227_/a_109_93# 2.5e-19
C458 _322_/a_761_289# _074_ 0.0107f
C459 net12 _078_ 0.111f
C460 calibrate _331_/a_193_47# 1.61e-19
C461 _329_/a_1108_47# trim_mask\[1\] 2.78e-20
C462 _169_/a_215_311# _060_ 5.66e-19
C463 _169_/a_109_53# net54 3.91e-19
C464 net27 _152_/a_68_297# 0.00901f
C465 net34 _296_/a_113_47# 1.59e-19
C466 _209_/a_27_47# _077_ 0.156f
C467 clknet_2_2__leaf_clk _330_/a_1462_47# 4.64e-19
C468 output12/a_27_47# net45 5.09e-20
C469 _040_ _247_/a_27_297# 4.86e-21
C470 VPWR _113_ 0.157f
C471 _248_/a_27_297# mask\[2\] 0.00222f
C472 _123_ _133_ 0.0618f
C473 _081_ mask\[0\] 1.69e-19
C474 net42 _098_ 0.173f
C475 net2 _040_ 1.61e-21
C476 _328_/a_27_47# trim_mask\[2\] 3.93e-19
C477 _327_/a_1270_413# _058_ 1.09e-19
C478 mask\[1\] _208_/a_76_199# 3.42e-19
C479 _328_/a_1462_47# trim_mask\[0\] 8.3e-20
C480 _292_/a_78_199# net2 0.0528f
C481 _334_/a_543_47# clknet_2_2__leaf_clk 7.44e-19
C482 clkbuf_2_1__f_clk/a_110_47# _245_/a_27_297# 0.0172f
C483 _331_/a_1462_47# _052_ 5.97e-20
C484 net50 _062_ 1.8e-19
C485 _052_ _260_/a_93_21# 0.0953f
C486 net43 _310_/a_639_47# 7.29e-19
C487 _311_/a_448_47# net53 0.00818f
C488 _022_ _010_ 5.28e-19
C489 VPWR _247_/a_27_297# 0.0708f
C490 _078_ net44 0.0366f
C491 _325_/a_27_47# net15 8.47e-19
C492 net42 clknet_0_clk 0.104f
C493 _101_ _244_/a_27_297# 0.0181f
C494 _045_ _084_ 0.0144f
C495 VPWR net2 1.44f
C496 mask\[5\] _220_/a_113_297# 0.032f
C497 _249_/a_109_297# _084_ 5e-20
C498 _064_ _058_ 0.12f
C499 _259_/a_109_297# _064_ 9.79e-19
C500 VPWR _305_/a_1283_21# 0.00312f
C501 _307_/a_27_47# _210_/a_113_297# 7.96e-20
C502 _107_ _075_ 5.06e-19
C503 _328_/a_27_47# _329_/a_27_47# 2.08e-20
C504 _341_/a_1283_21# net16 2.94e-20
C505 _231_/a_161_47# _195_/a_505_21# 0.0015f
C506 _051_ state\[1\] 0.354f
C507 VPWR _311_/a_1270_413# -2.28e-19
C508 output10/a_27_47# _335_/a_1108_47# 2.48e-20
C509 state\[2\] _169_/a_373_53# 1.35e-19
C510 net9 _298_/a_78_199# 0.00188f
C511 _042_ clknet_2_3__leaf_clk 1.61e-20
C512 state\[2\] net54 0.00408f
C513 _324_/a_27_47# clknet_2_1__leaf_clk 0.0144f
C514 net47 fanout47/a_27_47# 0.0251f
C515 _076_ _205_/a_27_47# 3.4e-20
C516 _074_ _101_ 0.969f
C517 _335_/a_193_47# clknet_2_2__leaf_clk 0.0017f
C518 VPWR _189_/a_218_47# -6.73e-19
C519 net30 _098_ 8.93e-20
C520 net14 net29 0.0335f
C521 _282_/a_150_297# _065_ 2.58e-19
C522 _182_/a_27_47# en_co_clk 6.91e-20
C523 net13 _232_/a_304_297# 9e-19
C524 _276_/a_145_75# VPWR 0.00165f
C525 _333_/a_193_47# net46 0.0284f
C526 clknet_0_clk _054_ 3.05e-19
C527 _053_ _058_ 0.00145f
C528 _323_/a_27_47# _150_/a_27_47# 1.06e-20
C529 net9 _341_/a_1108_47# 0.00738f
C530 _041_ net45 1.44e-20
C531 _336_/a_543_47# _033_ 4.03e-19
C532 clknet_0_clk net30 0.237f
C533 mask\[4\] _084_ 3.07e-20
C534 _265_/a_81_21# net46 0.00127f
C535 _232_/a_32_297# net41 4.77e-21
C536 _332_/a_27_47# clknet_2_2__leaf_clk 0.0281f
C537 _120_ _095_ 0.0354f
C538 en_co_clk _099_ 0.00304f
C539 _303_/a_193_47# _042_ 2.78e-21
C540 _235_/a_79_21# _050_ 2.2e-19
C541 _050_ net15 3.54e-20
C542 _339_/a_1140_413# _123_ 0.00177f
C543 cal_itt\[1\] clkbuf_2_3__f_clk/a_110_47# 0.0102f
C544 _268_/a_75_212# clknet_2_2__leaf_clk 0.0215f
C545 net43 _305_/a_651_413# 0.00129f
C546 _308_/a_27_47# net22 1.73e-19
C547 output25/a_27_47# clknet_2_1__leaf_clk 0.0196f
C548 _321_/a_27_47# _321_/a_1108_47# -2.98e-20
C549 _319_/a_193_47# _282_/a_68_297# 4.88e-19
C550 trim_mask\[3\] _335_/a_543_47# 4.03e-20
C551 net50 _335_/a_761_289# 0.00471f
C552 trim_val\[3\] _335_/a_1283_21# 0.00206f
C553 _168_/a_27_413# clknet_0_clk 0.00165f
C554 _214_/a_113_297# clknet_2_0__leaf_clk 1.88e-20
C555 _247_/a_27_297# net52 0.0162f
C556 _293_/a_81_21# _144_/a_27_47# 0.0184f
C557 _247_/a_109_47# _101_ 2.72e-19
C558 VPWR _232_/a_32_297# 0.0782f
C559 _008_ _311_/a_448_47# 0.00199f
C560 VPWR _221_/a_109_297# -6.61e-19
C561 _292_/a_78_199# _123_ 0.0152f
C562 _062_ _279_/a_396_47# 1.82e-19
C563 _041_ _065_ 0.204f
C564 _317_/a_761_289# net14 6.77e-20
C565 _014_ _316_/a_1270_413# 5.82e-20
C566 net45 _316_/a_651_413# 0.00164f
C567 _307_/a_193_47# _315_/a_193_47# 2.34e-19
C568 _309_/a_27_47# net26 4.53e-21
C569 trim_val\[4\] _278_/a_27_47# 3.3e-19
C570 calibrate _260_/a_93_21# 0.007f
C571 net2 _063_ 1.05e-19
C572 VPWR trim_val\[1\] 0.607f
C573 trim_mask\[4\] net46 0.468f
C574 _320_/a_543_47# _078_ 7.94e-20
C575 _305_/a_1283_21# _063_ 3.38e-19
C576 _337_/a_193_47# _337_/a_1283_21# -6.53e-19
C577 _337_/a_27_47# _337_/a_1108_47# -2.98e-20
C578 _307_/a_448_47# net30 4.57e-19
C579 net24 _320_/a_27_47# 1.18e-19
C580 VPWR net29 0.807f
C581 _126_ _339_/a_27_47# 1.75e-20
C582 _320_/a_193_47# clknet_2_0__leaf_clk 0.00228f
C583 VPWR _123_ 2.87f
C584 net9 _339_/a_476_47# 0.0108f
C585 _257_/a_373_47# trim_mask\[1\] 0.00244f
C586 _256_/a_109_297# _302_/a_27_297# 4.61e-21
C587 net27 mask\[5\] 0.689f
C588 _036_ net2 0.152f
C589 _074_ _312_/a_448_47# 2.76e-20
C590 net13 _317_/a_1108_47# 2.3e-20
C591 net47 _287_/a_75_212# 0.0126f
C592 _097_ _013_ 8.57e-19
C593 _250_/a_373_47# net53 0.00125f
C594 _042_ net20 1.83e-22
C595 _291_/a_117_297# cal_count\[0\] 0.00146f
C596 clknet_0_clk _072_ 0.00187f
C597 _042_ net53 0.369f
C598 _331_/a_27_47# _171_/a_27_47# 3.56e-21
C599 net25 net15 4.23e-21
C600 net4 _336_/a_193_47# 0.0115f
C601 _324_/a_193_47# mask\[6\] 6.26e-20
C602 _333_/a_543_47# rebuffer2/a_75_212# 0.00125f
C603 _110_ _191_/a_27_297# 4.33e-20
C604 _237_/a_505_21# _192_/a_505_280# 9.76e-19
C605 _092_ net40 1.05e-19
C606 VPWR _227_/a_209_311# -0.0067f
C607 _333_/a_1283_21# _108_ 0.0051f
C608 _187_/a_27_413# trim_val\[0\] 9.02e-21
C609 _307_/a_1108_47# mask\[0\] 8.21e-19
C610 _307_/a_1283_21# _078_ 0.0109f
C611 _307_/a_448_47# net22 1.88e-19
C612 VPWR _251_/a_373_47# -4.3e-19
C613 trim[4] net35 0.00211f
C614 trim_val\[0\] _332_/a_27_47# 1.07e-19
C615 _051_ _336_/a_651_413# 7.37e-21
C616 _307_/a_27_47# net45 0.00153f
C617 _307_/a_761_289# clknet_2_0__leaf_clk 2.62e-19
C618 _329_/a_805_47# net9 4.44e-19
C619 trim[3] _334_/a_193_47# 1.78e-19
C620 VPWR _317_/a_761_289# 0.0113f
C621 output35/a_27_47# comp 3.98e-20
C622 _060_ _226_/a_109_47# 8.38e-19
C623 _136_ _066_ 0.0389f
C624 output27/a_27_47# result[5] 0.00955f
C625 _322_/a_448_47# _042_ 2.87e-20
C626 _298_/a_292_297# cal_count\[2\] 7.38e-20
C627 _235_/a_382_297# _092_ 0.00169f
C628 _304_/a_651_413# _136_ 3.08e-19
C629 _304_/a_543_47# _038_ 2.52e-20
C630 clk net55 0.00591f
C631 _293_/a_299_297# net47 2.46e-20
C632 _064_ en_co_clk 3.22e-20
C633 net8 net34 0.0332f
C634 net55 clone7/a_27_47# 0.0294f
C635 _304_/a_651_413# _284_/a_68_297# 3e-20
C636 ctlp[7] _313_/a_1108_47# 1.83e-19
C637 _033_ _106_ 6.82e-20
C638 rebuffer3/a_75_212# net18 0.0112f
C639 _269_/a_81_21# _333_/a_193_47# 0.00164f
C640 cal_itt\[1\] cal_count\[3\] 7.38e-21
C641 _276_/a_59_75# clknet_2_2__leaf_clk 8.39e-22
C642 _123_ _063_ 0.00752f
C643 trim_mask\[0\] _091_ 7.39e-20
C644 _113_ _333_/a_448_47# 1.68e-20
C645 _030_ _333_/a_1108_47# 1.61e-19
C646 _256_/a_109_297# trim_mask\[0\] 0.0723f
C647 _315_/a_193_47# output41/a_27_47# 5.23e-20
C648 _340_/a_193_47# net47 9.57e-19
C649 ctln[7] _318_/a_448_47# 5.95e-20
C650 net13 _318_/a_1270_413# 5.91e-20
C651 cal_itt\[0\] _198_/a_27_47# 0.00901f
C652 calibrate net3 0.00995f
C653 _319_/a_1283_21# _121_ 0.00141f
C654 net4 net55 1.05e-20
C655 clknet_2_1__leaf_clk _312_/a_543_47# 2.56e-19
C656 net44 _319_/a_651_413# 2.61e-20
C657 _308_/a_448_47# net24 9.84e-21
C658 _301_/a_47_47# clkc 7.43e-20
C659 mask\[0\] net14 0.00272f
C660 _308_/a_1108_47# net45 0.012f
C661 net28 result[7] 0.11f
C662 _007_ _310_/a_27_47# 0.0361f
C663 _036_ _123_ 0.0118f
C664 _008_ _042_ 6.43e-21
C665 VPWR _296_/a_113_47# -1.33e-19
C666 _053_ en_co_clk 0.014f
C667 _065_ net18 0.661f
C668 _341_/a_651_413# _065_ 9.16e-19
C669 VPWR _114_ 0.104f
C670 _309_/a_193_47# _078_ 0.0278f
C671 _276_/a_59_75# net11 9.67e-20
C672 _292_/a_215_47# net16 0.00111f
C673 _119_ _049_ 1.08e-19
C674 _251_/a_373_47# net52 6.65e-19
C675 _237_/a_76_199# net45 3.57e-21
C676 _237_/a_505_21# _014_ 2.65e-20
C677 VPWR ctlp[1] 0.175f
C678 _101_ net26 0.261f
C679 _336_/a_761_289# clkbuf_2_2__f_clk/a_110_47# 0.00792f
C680 net43 _203_/a_59_75# 1.14e-20
C681 net25 _310_/a_193_47# 0.00792f
C682 net15 _246_/a_109_47# 5.78e-20
C683 _051_ _337_/a_1108_47# 1.6e-19
C684 VPWR _318_/a_1108_47# 0.0217f
C685 output36/a_27_47# output38/a_27_47# 0.00249f
C686 _325_/a_1283_21# _074_ 0.00417f
C687 _117_ _275_/a_299_297# 2.22e-19
C688 _276_/a_145_75# net50 1.8e-20
C689 _327_/a_27_47# net46 0.00414f
C690 _167_/a_161_47# _051_ 0.00947f
C691 _189_/a_408_47# _107_ 0.00102f
C692 _035_ _338_/a_476_47# 0.0101f
C693 net13 clknet_2_0__leaf_clk 0.164f
C694 net4 _067_ 0.0556f
C695 _289_/a_68_297# _297_/a_285_47# 2.98e-19
C696 trim_mask\[2\] _336_/a_1108_47# 1.12e-19
C697 net4 _070_ 0.138f
C698 trim_mask\[0\] _033_ 0.00407f
C699 _024_ _106_ 7.33e-22
C700 _324_/a_639_47# _021_ 1.9e-19
C701 comp net40 2.43e-19
C702 VPWR _168_/a_207_413# 0.00658f
C703 ctlp[6] output21/a_27_47# 4.08e-19
C704 state\[2\] _228_/a_382_297# 1.95e-19
C705 _087_ _049_ 8.72e-19
C706 _259_/a_109_297# _027_ 0.00307f
C707 _259_/a_27_297# net46 0.00358f
C708 _328_/a_1108_47# VPWR 0.00673f
C709 _208_/a_218_374# _076_ 4.55e-19
C710 _208_/a_505_21# _077_ 4.91e-20
C711 trim_val\[0\] _332_/a_1217_47# 3.85e-20
C712 VPWR mask\[0\] 1.1f
C713 _207_/a_109_297# _076_ 0.00288f
C714 _074_ _248_/a_27_297# 0.00126f
C715 _307_/a_1217_47# net45 8.84e-20
C716 calibrate _241_/a_388_297# 9.09e-20
C717 _308_/a_1283_21# _319_/a_193_47# 1.03e-19
C718 _308_/a_1108_47# _319_/a_27_47# 1.09e-19
C719 _311_/a_1283_21# _152_/a_68_297# 6.2e-22
C720 VPWR output24/a_27_47# 0.0801f
C721 _110_ _265_/a_81_21# 0.00533f
C722 _307_/a_1283_21# _004_ 1.29e-20
C723 en_co_clk _226_/a_109_47# 1.05e-19
C724 _321_/a_27_47# _214_/a_113_297# 8.73e-21
C725 _315_/a_1270_413# net14 1.25e-19
C726 trim_mask\[3\] trim_mask\[1\] 1.44e-19
C727 _322_/a_543_47# _078_ 7.59e-21
C728 _019_ _042_ 7.08e-19
C729 mask\[6\] net21 0.00186f
C730 _104_ _228_/a_79_21# 0.0025f
C731 _110_ _048_ 0.0039f
C732 _319_/a_1108_47# clknet_0_clk 0.0083f
C733 net47 _136_ 0.00242f
C734 _122_ _067_ 1.5e-19
C735 net47 _284_/a_68_297# 0.00446f
C736 _304_/a_805_47# _122_ 6.43e-19
C737 net14 ctln[0] 0.00137f
C738 VPWR _150_/a_27_47# 0.0513f
C739 _021_ _312_/a_193_47# 1.23e-20
C740 _340_/a_652_21# _122_ 0.00191f
C741 _112_ _333_/a_543_47# 0.00315f
C742 net49 _333_/a_1283_21# 1.09e-19
C743 trim_val\[1\] _333_/a_448_47# 9.97e-20
C744 trim_mask\[1\] _333_/a_1108_47# 4.23e-19
C745 _293_/a_81_21# _299_/a_298_297# 2.3e-21
C746 _304_/a_761_289# net18 0.01f
C747 _110_ trim_mask\[4\] 0.0431f
C748 trim_mask\[2\] _256_/a_27_297# 5.93e-21
C749 _258_/a_27_297# trim_mask\[0\] 6.41e-20
C750 _107_ _170_/a_81_21# 0.00403f
C751 _340_/a_1032_413# _041_ 9.24e-22
C752 trim_mask\[0\] _024_ 0.122f
C753 _340_/a_796_47# net47 3.82e-19
C754 _315_/a_448_47# valid 0.00102f
C755 _325_/a_193_47# clknet_2_1__leaf_clk 0.00679f
C756 _144_/a_27_47# net34 3.57e-21
C757 net23 mask\[0\] 0.241f
C758 _108_ trim_val\[4\] 0.263f
C759 _327_/a_543_47# _108_ 5.7e-19
C760 _340_/a_652_21# _037_ 7.99e-19
C761 _005_ net24 0.00456f
C762 net23 output24/a_27_47# 0.0138f
C763 net5 clknet_2_3__leaf_clk 7.24e-20
C764 net43 clknet_2_0__leaf_clk 0.373f
C765 _327_/a_761_289# _111_ 2.55e-19
C766 result[4] _310_/a_27_47# 0.0131f
C767 _309_/a_1462_47# _078_ 0.00213f
C768 mask\[4\] _311_/a_193_47# 0.0256f
C769 _107_ _227_/a_296_53# 9.57e-20
C770 _323_/a_448_47# _043_ 7.3e-22
C771 mask\[1\] _247_/a_109_297# 1.12e-20
C772 clkbuf_0_clk/a_110_47# _041_ 6.5e-21
C773 VPWR _315_/a_1270_413# -1.45e-19
C774 _053_ _286_/a_76_199# 1.01e-19
C775 _337_/a_639_47# net44 -7.75e-19
C776 _329_/a_27_47# _256_/a_27_297# 1.23e-19
C777 _313_/a_761_289# _010_ 4.31e-19
C778 net35 _108_ 0.00122f
C779 _062_ _278_/a_109_297# 2.94e-21
C780 mask\[0\] net52 5.84e-19
C781 _058_ _332_/a_1108_47# 0.00185f
C782 _334_/a_193_47# _057_ 5.45e-20
C783 _233_/a_109_47# cal 1.54e-19
C784 _233_/a_109_297# net1 0.00361f
C785 net48 clknet_2_2__leaf_clk 2.26e-20
C786 _058_ _029_ 0.00671f
C787 _239_/a_474_297# _048_ 0.00726f
C788 _328_/a_27_47# _333_/a_27_47# 1.45e-19
C789 _327_/a_1217_47# net46 2.16e-19
C790 _291_/a_117_297# net16 7.79e-19
C791 _146_/a_68_297# mask\[1\] 1.08e-21
C792 clkbuf_2_0__f_clk/a_110_47# _095_ 0.117f
C793 VPWR ctln[0] 0.0202f
C794 net31 input2/a_27_47# 0.00901f
C795 clknet_2_2__leaf_clk net30 0.00237f
C796 _043_ net18 0.0203f
C797 clk _316_/a_543_47# 4.67e-19
C798 _149_/a_68_297# _303_/a_761_289# 5.23e-19
C799 net39 net33 1.61e-20
C800 _302_/a_27_297# clkbuf_2_3__f_clk/a_110_47# 2.93e-20
C801 net12 ctln[6] 0.00602f
C802 output14/a_27_47# _314_/a_27_47# 0.0023f
C803 _293_/a_81_21# _133_ 1.84e-20
C804 _168_/a_27_413# clknet_2_2__leaf_clk 6.96e-20
C805 _059_ _062_ 0.102f
C806 net3 _317_/a_1108_47# 1.46e-20
C807 _254_/a_109_297# _050_ 1.84e-20
C808 _323_/a_193_47# net47 -0.00111f
C809 _328_/a_1283_21# clknet_2_2__leaf_clk 0.0763f
C810 _106_ clkbuf_2_3__f_clk/a_110_47# 0.00664f
C811 _304_/a_448_47# clknet_2_3__leaf_clk 0.0162f
C812 _136_ _301_/a_47_47# 0.00153f
C813 _340_/a_27_47# _133_ 2.33e-22
C814 VPWR net8 0.25f
C815 _341_/a_27_47# _136_ 0.0151f
C816 _302_/a_109_297# net18 0.0044f
C817 mask\[5\] _311_/a_1283_21# 5.66e-20
C818 _060_ _093_ 0.00231f
C819 _007_ clknet_2_1__leaf_clk 0.233f
C820 _325_/a_761_289# mask\[6\] 0.0219f
C821 _338_/a_27_47# _122_ 0.00155f
C822 _341_/a_27_47# _284_/a_68_297# 3.15e-19
C823 _048_ _192_/a_476_47# 0.00151f
C824 net45 _090_ 1.49e-20
C825 net48 _333_/a_651_413# 6.72e-21
C826 _041_ _338_/a_476_47# 3.12e-19
C827 net47 _338_/a_1140_413# -6.31e-19
C828 net3 _192_/a_27_47# 0.0394f
C829 clknet_2_1__leaf_clk _249_/a_27_297# 0.058f
C830 _338_/a_27_47# _338_/a_381_47# -0.00438f
C831 _306_/a_193_47# rebuffer4/a_27_47# 3.29e-21
C832 net13 _321_/a_27_47# 4.31e-21
C833 _051_ clkbuf_2_2__f_clk/a_110_47# 6.84e-19
C834 mask\[3\] clknet_2_1__leaf_clk 0.737f
C835 net13 _337_/a_27_47# 0.0153f
C836 _335_/a_27_47# _330_/a_1108_47# 8.91e-19
C837 _335_/a_193_47# _330_/a_1283_21# 0.00203f
C838 _100_ net41 0.0383f
C839 net16 _333_/a_639_47# 0.0015f
C840 net2 input2/a_27_47# 0.0135f
C841 _110_ _327_/a_27_47# 1.76e-20
C842 _277_/a_75_212# trim_val\[3\] 4.8e-19
C843 _340_/a_1032_413# _129_ 4.17e-19
C844 _232_/a_32_297# _034_ 1.16e-19
C845 result[4] _310_/a_1217_47# 6.14e-21
C846 mask\[4\] _311_/a_1462_47# 0.00185f
C847 _090_ _065_ 1.37e-19
C848 _168_/a_297_47# _107_ 2.5e-19
C849 VPWR _319_/a_448_47# 0.0023f
C850 _062_ _075_ 0.281f
C851 VPWR _230_/a_145_75# -4.39e-19
C852 trim_mask\[0\] clkbuf_2_3__f_clk/a_110_47# 0.127f
C853 net47 clknet_0_clk 5.33e-19
C854 _012_ net1 0.0346f
C855 _104_ fanout46/a_27_47# 0.0101f
C856 _300_/a_47_47# en_co_clk 1.4e-19
C857 VPWR _100_ 0.248f
C858 _323_/a_193_47# net44 0.00488f
C859 _320_/a_448_47# _143_/a_68_297# 9.86e-19
C860 _328_/a_1108_47# _333_/a_448_47# 6.86e-21
C861 trim[4] _332_/a_27_47# 6.64e-20
C862 net15 _314_/a_1108_47# 1.64e-20
C863 _074_ _156_/a_27_47# 2.4e-19
C864 net47 _339_/a_27_47# 0.012f
C865 output20/a_27_47# VPWR 0.0522f
C866 trim_mask\[0\] _134_ 1.05e-19
C867 net12 _098_ 0.0253f
C868 _326_/a_761_289# _314_/a_761_289# 0.00117f
C869 _326_/a_193_47# _314_/a_543_47# 2.28e-19
C870 _326_/a_543_47# _314_/a_193_47# 1.97e-20
C871 trim_mask\[1\] _118_ 4.41e-20
C872 _340_/a_1032_413# _339_/a_1032_413# 7.46e-19
C873 net46 net40 0.33f
C874 _303_/a_1283_21# _035_ 0.00101f
C875 _327_/a_1283_21# trim_mask\[1\] 5.11e-23
C876 _198_/a_27_47# _069_ 0.044f
C877 clknet_2_1__leaf_clk _220_/a_113_297# 0.00345f
C878 _195_/a_505_21# _062_ 1.26e-20
C879 net2 _208_/a_76_199# 9.76e-19
C880 _255_/a_27_47# _107_ 0.00512f
C881 _302_/a_27_297# cal_count\[3\] 0.013f
C882 trim[3] trim_val\[2\] 8.5e-19
C883 net30 _279_/a_204_297# 1.45e-19
C884 _330_/a_639_47# net46 -7.75e-19
C885 net12 clknet_0_clk 0.0103f
C886 _048_ net45 4.74e-19
C887 _293_/a_81_21# VPWR 0.00604f
C888 net43 _319_/a_639_47# -5.18e-19
C889 net12 _320_/a_1108_47# 7.6e-22
C890 _323_/a_1462_47# net47 -6.49e-19
C891 net3 clknet_2_0__leaf_clk 0.0115f
C892 _326_/a_27_47# _310_/a_27_47# 9.43e-22
C893 net43 _321_/a_27_47# 0.149f
C894 _106_ cal_count\[3\] 0.00111f
C895 VPWR _336_/a_805_47# 2.92e-19
C896 _198_/a_109_47# _067_ 0.00165f
C897 VPWR _264_/a_27_297# 0.0252f
C898 VPWR _304_/a_1270_413# 4.74e-20
C899 _334_/a_27_47# net46 0.206f
C900 mask\[6\] _045_ 0.00847f
C901 VPWR _340_/a_27_47# -0.227f
C902 net43 _337_/a_27_47# 5.87e-20
C903 mask\[6\] _249_/a_109_297# 1.44e-19
C904 _341_/a_1217_47# _136_ 1.18e-19
C905 _038_ net18 0.0268f
C906 _103_ _048_ 0.481f
C907 net45 trim_mask\[4\] 0.103f
C908 _250_/a_109_297# mask\[5\] 0.0121f
C909 _078_ _155_/a_68_297# 0.00101f
C910 fanout47/a_27_47# net19 0.00323f
C911 _093_ en_co_clk 0.00338f
C912 trim_mask\[4\] rebuffer3/a_75_212# 1.36e-21
C913 ctlp[7] net28 0.00152f
C914 net43 _069_ 7.84e-21
C915 _182_/a_27_47# net16 7.97e-19
C916 clkbuf_2_1__f_clk/a_110_47# mask\[2\] 0.014f
C917 net51 _208_/a_218_47# 1.68e-19
C918 _110_ _178_/a_68_297# 0.0586f
C919 result[4] clknet_2_1__leaf_clk 0.0505f
C920 _319_/a_1283_21# _016_ 6.74e-20
C921 _048_ _065_ 0.0175f
C922 _099_ _049_ 0.0156f
C923 _230_/a_145_75# _063_ 6.66e-19
C924 net44 clknet_0_clk 0.00545f
C925 _334_/a_27_47# _334_/a_639_47# -0.00188f
C926 _338_/a_476_47# net18 0.00994f
C927 _341_/a_27_47# _341_/a_761_289# -0.017f
C928 clone1/a_27_47# _260_/a_93_21# 2.25e-20
C929 _320_/a_1108_47# net44 -0.00283f
C930 VPWR _144_/a_27_47# 0.0478f
C931 net47 _303_/a_27_47# 0.00738f
C932 cal_itt\[2\] _190_/a_655_47# 7.83e-20
C933 _048_ _105_ 0.152f
C934 _336_/a_27_47# net19 0.0145f
C935 _169_/a_215_311# _049_ 6.23e-21
C936 _169_/a_215_311# _318_/a_761_289# 0.00109f
C937 net13 _051_ 0.0111f
C938 _290_/a_207_413# _288_/a_59_75# 1.16e-19
C939 _332_/a_448_47# net40 6.16e-19
C940 mask\[6\] mask\[4\] 5.62e-20
C941 net28 _313_/a_543_47# 0.0358f
C942 output18/a_27_47# ctlp[4] 0.0188f
C943 output21/a_27_47# net21 0.00609f
C944 _329_/a_193_47# trim_mask\[2\] 2.65e-19
C945 trim_mask\[0\] cal_count\[3\] 2.78e-19
C946 clknet_0_clk _003_ 1.8e-20
C947 ctln[4] _335_/a_1108_47# 2.83e-19
C948 net4 clknet_2_3__leaf_clk 0.0256f
C949 _014_ _241_/a_105_352# 0.0343f
C950 VPWR _321_/a_1270_413# 3.1e-20
C951 _339_/a_193_47# _122_ 6.01e-21
C952 _116_ _104_ 1.8e-20
C953 net27 clknet_2_1__leaf_clk 0.0557f
C954 _276_/a_59_75# _330_/a_1283_21# 7.73e-20
C955 _041_ _339_/a_1182_261# 0.0204f
C956 mask\[1\] _078_ 0.884f
C957 _257_/a_27_297# trim_mask\[0\] 6.95e-19
C958 _333_/a_1108_47# _056_ 1.92e-19
C959 clknet_2_1__leaf_clk _222_/a_113_297# 0.0129f
C960 VPWR _313_/a_1283_21# 0.0288f
C961 net47 _339_/a_586_47# 1.16e-19
C962 VPWR _337_/a_1270_413# 6.54e-20
C963 _264_/a_27_297# _063_ 3.05e-19
C964 _336_/a_27_47# _107_ 0.00341f
C965 _309_/a_27_47# _102_ 4.1e-21
C966 _037_ _339_/a_193_47# 2.07e-20
C967 trim_mask\[2\] net18 0.00588f
C968 output22/a_27_47# _307_/a_27_47# 0.0112f
C969 _316_/a_193_47# net14 3.78e-20
C970 _289_/a_68_297# _288_/a_59_75# 0.00852f
C971 _050_ wire42/a_75_212# 3.15e-19
C972 net34 _133_ 2.23e-20
C973 clknet_2_1__leaf_clk rebuffer5/a_161_47# 0.011f
C974 _159_/a_27_47# _313_/a_543_47# 9.58e-20
C975 _051_ _331_/a_193_47# 0.00143f
C976 _292_/a_292_297# net47 4.05e-19
C977 _340_/a_1032_413# _297_/a_47_47# 6.74e-20
C978 _015_ _318_/a_1108_47# 1.26e-19
C979 state\[2\] _318_/a_193_47# 0.00398f
C980 fanout44/a_27_47# clknet_2_0__leaf_clk 0.0446f
C981 _036_ _340_/a_27_47# 0.00113f
C982 _128_ _340_/a_1182_261# 3.45e-20
C983 mask\[0\] _034_ 8.14e-22
C984 _134_ _298_/a_78_199# 2.16e-19
C985 _122_ clknet_2_3__leaf_clk 0.15f
C986 _081_ net14 0.0112f
C987 net36 _126_ 6.86e-20
C988 _303_/a_27_47# net44 0.00597f
C989 _323_/a_1108_47# net18 2.68e-19
C990 _320_/a_543_47# clknet_0_clk 0.00449f
C991 _262_/a_109_297# _092_ 1.19e-19
C992 net43 _321_/a_1217_47# 7.34e-19
C993 trim[1] net37 0.0301f
C994 _326_/a_543_47# _074_ 0.0147f
C995 _338_/a_381_47# clknet_2_3__leaf_clk 0.0159f
C996 ctln[6] ctln[7] 0.00465f
C997 _320_/a_193_47# _320_/a_651_413# -0.00701f
C998 _309_/a_761_289# _081_ 1.59e-19
C999 _309_/a_27_47# _006_ 0.0365f
C1000 _334_/a_1217_47# net46 1.06e-20
C1001 _271_/a_75_212# net46 0.0424f
C1002 _066_ clknet_2_2__leaf_clk 6.69e-19
C1003 _194_/a_113_297# trim_mask\[4\] 1.81e-20
C1004 clk valid 5.35e-20
C1005 _316_/a_193_47# net41 0.0258f
C1006 VPWR _340_/a_586_47# 2.04e-19
C1007 _037_ clknet_2_3__leaf_clk 0.0387f
C1008 net43 _313_/a_651_413# 0.0032f
C1009 _329_/a_193_47# _115_ 7.12e-20
C1010 _021_ mask\[5\] 5.92e-20
C1011 _315_/a_1108_47# _099_ 1.31e-19
C1012 _129_ _298_/a_292_297# 2.17e-20
C1013 _299_/a_298_297# _133_ 1.4e-21
C1014 _336_/a_1283_21# trim_mask\[4\] 0.052f
C1015 _036_ _144_/a_27_47# 6.61e-21
C1016 _306_/a_27_47# clknet_2_1__leaf_clk 5.04e-20
C1017 _061_ _161_/a_68_297# 2.27e-20
C1018 _234_/a_109_297# _092_ 3.9e-19
C1019 _308_/a_193_47# _307_/a_543_47# 1.91e-19
C1020 _059_ _232_/a_32_297# 4.28e-19
C1021 _338_/a_1224_47# net18 1.57e-19
C1022 _336_/a_27_47# _279_/a_27_47# 1.13e-20
C1023 _081_ _040_ 0.165f
C1024 _283_/a_75_212# _065_ 0.0287f
C1025 rebuffer1/a_75_212# rebuffer2/a_75_212# 5.35e-19
C1026 mask\[3\] net45 4.53e-21
C1027 _327_/a_27_47# rebuffer3/a_75_212# 3.91e-19
C1028 _050_ _319_/a_193_47# 5.42e-21
C1029 _107_ _096_ 3.94e-19
C1030 VPWR _316_/a_193_47# 0.0464f
C1031 _332_/a_27_47# _108_ 0.445f
C1032 _332_/a_193_47# _332_/a_761_289# -0.0113f
C1033 _332_/a_27_47# _332_/a_543_47# -0.00297f
C1034 net47 _303_/a_1217_47# 2.63e-19
C1035 output34/a_27_47# net33 0.00131f
C1036 _189_/a_218_47# _075_ 4.95e-20
C1037 _268_/a_75_212# _108_ 0.0365f
C1038 _328_/a_639_47# _058_ 5.31e-19
C1039 _335_/a_639_47# net46 0.00387f
C1040 _104_ _328_/a_27_47# 0.0099f
C1041 _053_ _049_ 0.32f
C1042 _053_ _318_/a_761_289# 8.36e-20
C1043 state\[0\] _318_/a_543_47# 4.69e-20
C1044 clk _331_/a_448_47# 0.00869f
C1045 _097_ net1 3.15e-20
C1046 net12 _322_/a_1108_47# 0.00241f
C1047 _105_ _190_/a_27_47# 9.22e-20
C1048 net12 _331_/a_1108_47# 0.00143f
C1049 VPWR _081_ 0.565f
C1050 _110_ net40 1.8e-20
C1051 trim_val\[2\] _057_ 5.23e-20
C1052 _251_/a_27_297# _085_ 1.1e-19
C1053 mask\[6\] _222_/a_199_47# 4.87e-19
C1054 _327_/a_27_47# _065_ 2.04e-20
C1055 _333_/a_1108_47# _173_/a_27_47# 4.54e-19
C1056 _329_/a_1462_47# trim_mask\[2\] 5.43e-19
C1057 mask\[3\] _065_ 2.22e-20
C1058 net43 _023_ 0.00497f
C1059 state\[1\] _099_ 6.04e-22
C1060 _324_/a_448_47# net44 0.00173f
C1061 net2 _295_/a_113_47# 1.11e-19
C1062 _332_/a_1270_413# net46 5.88e-19
C1063 _324_/a_1108_47# _323_/a_27_47# 2.06e-19
C1064 _324_/a_1283_21# _323_/a_193_47# 0.00889f
C1065 _041_ _339_/a_1296_47# 0.00205f
C1066 _094_ clkbuf_2_1__f_clk/a_110_47# 2.84e-21
C1067 net3 _337_/a_27_47# 6.19e-19
C1068 net16 _057_ 1.4e-20
C1069 _326_/a_27_47# clknet_2_1__leaf_clk 0.138f
C1070 _308_/a_193_47# _138_/a_27_47# 7.99e-20
C1071 _189_/a_27_47# _088_ 8.22e-20
C1072 _110_ _267_/a_145_75# 5.4e-19
C1073 VPWR _323_/a_27_47# 0.0702f
C1074 result[0] _307_/a_1108_47# 3.43e-19
C1075 _030_ _332_/a_193_47# 6.47e-22
C1076 clknet_2_0__leaf_clk _281_/a_103_199# 1.79e-19
C1077 _309_/a_1108_47# _214_/a_113_297# 6.28e-19
C1078 net1 _315_/a_543_47# 0.00105f
C1079 _102_ _101_ 0.00317f
C1080 _322_/a_1108_47# net44 0.0188f
C1081 _169_/a_215_311# state\[1\] 0.0644f
C1082 _074_ _310_/a_1108_47# 5.17e-19
C1083 _314_/a_27_47# net29 0.00203f
C1084 _292_/a_493_297# _122_ 2.52e-19
C1085 net54 net45 0.00148f
C1086 _309_/a_193_47# _308_/a_27_47# 4.17e-21
C1087 _309_/a_27_47# _308_/a_193_47# 1.51e-19
C1088 _233_/a_373_47# _093_ 0.00125f
C1089 _340_/a_193_47# _001_ 5.65e-20
C1090 _233_/a_109_297# _012_ 0.051f
C1091 _110_ _334_/a_27_47# 0.00314f
C1092 net31 _030_ 1.25e-20
C1093 VPWR net34 0.923f
C1094 net21 _313_/a_1270_413# 5.17e-20
C1095 _051_ _260_/a_93_21# 0.00143f
C1096 net23 _081_ 0.0986f
C1097 _104_ _262_/a_27_47# 8.47e-20
C1098 _282_/a_68_297# _090_ 3.1e-19
C1099 _062_ _170_/a_81_21# 6.81e-21
C1100 _311_/a_27_47# _311_/a_448_47# -0.00346f
C1101 _311_/a_193_47# _311_/a_1108_47# -0.00656f
C1102 VPWR _301_/a_377_297# 0.00365f
C1103 _061_ _300_/a_47_47# 2.52e-20
C1104 _302_/a_109_297# trim_mask\[4\] 2.67e-20
C1105 net30 _278_/a_27_47# 0.0016f
C1106 _341_/a_1108_47# cal_count\[3\] 0.0541f
C1107 VPWR _338_/a_956_413# 2.06e-20
C1108 comp _132_ 0.00448f
C1109 _341_/a_805_47# clknet_2_3__leaf_clk 8.08e-19
C1110 VPWR _341_/a_193_47# -0.305f
C1111 en_co_clk _192_/a_505_280# 0.0534f
C1112 cal_itt\[1\] en_co_clk 0.133f
C1113 net4 _266_/a_68_297# 0.00574f
C1114 _323_/a_543_47# _303_/a_651_413# 4.92e-20
C1115 _323_/a_1108_47# _303_/a_1108_47# 1.46e-20
C1116 net2 _332_/a_761_289# 1.86e-20
C1117 _050_ _206_/a_27_93# 0.0521f
C1118 trim_mask\[0\] _242_/a_297_47# 2.27e-21
C1119 net54 _065_ 0.0141f
C1120 _316_/a_1462_47# net41 0.00184f
C1121 _339_/a_27_47# _339_/a_956_413# -0.00135f
C1122 _319_/a_761_289# _092_ 2.39e-20
C1123 net13 _320_/a_651_413# 0.00125f
C1124 _081_ net52 1.28e-19
C1125 VPWR _299_/a_298_297# -0.00451f
C1126 _272_/a_81_21# _334_/a_543_47# 6.99e-19
C1127 _320_/a_1283_21# _040_ 0.00251f
C1128 _053_ _262_/a_193_297# 0.00716f
C1129 _113_ _030_ 0.018f
C1130 clknet_2_1__leaf_clk _314_/a_448_47# 0.00142f
C1131 _307_/a_1108_47# net14 0.00335f
C1132 net15 _318_/a_27_47# 7.97e-21
C1133 mask\[0\] output30/a_27_47# 2.42e-21
C1134 _210_/a_113_297# sample 3.8e-19
C1135 _336_/a_27_47# _118_ 1.22e-19
C1136 _336_/a_193_47# trim_val\[4\] 0.0126f
C1137 clkbuf_2_2__f_clk/a_110_47# _119_ 0.151f
C1138 result[0] net14 0.00258f
C1139 VPWR _316_/a_1462_47# 6.13e-20
C1140 net4 _199_/a_109_297# 7.7e-19
C1141 _303_/a_1283_21# net18 6.47e-19
C1142 output27/a_27_47# _011_ 0.00178f
C1143 net44 _263_/a_79_21# 9.65e-21
C1144 _029_ _332_/a_639_47# 2.29e-19
C1145 trim_mask\[0\] _265_/a_299_297# 9.81e-19
C1146 VPWR _320_/a_1283_21# 0.0209f
C1147 _060_ _243_/a_27_297# 0.0719f
C1148 _185_/a_68_297# _096_ 0.00131f
C1149 clk _028_ 0.0679f
C1150 _050_ _337_/a_543_47# 5.57e-20
C1151 _087_ _240_/a_109_297# 0.00257f
C1152 _229_/a_27_297# _098_ 4.93e-19
C1153 net54 _243_/a_109_297# 4.43e-19
C1154 fanout43/a_27_47# net45 0.08f
C1155 clknet_2_1__leaf_clk _310_/a_761_289# 0.0198f
C1156 _047_ trim_val\[0\] 0.0259f
C1157 _333_/a_805_47# net32 6.64e-20
C1158 output21/a_27_47# _045_ 0.0124f
C1159 _088_ _227_/a_109_93# 4e-20
C1160 _326_/a_193_47# mask\[6\] 4.14e-20
C1161 _326_/a_543_47# net26 2.32e-20
C1162 fanout44/a_27_47# _337_/a_27_47# 8.93e-21
C1163 _136_ _001_ 0.00119f
C1164 clkbuf_2_0__f_clk/a_110_47# calibrate 7e-21
C1165 _333_/a_1108_47# _172_/a_68_297# 1.43e-19
C1166 _292_/a_78_199# _133_ 1.09e-20
C1167 _128_ _298_/a_78_199# 1.32e-20
C1168 _304_/a_1283_21# _092_ 4.48e-20
C1169 _308_/a_761_289# net43 0.00883f
C1170 _308_/a_543_47# _005_ 0.00354f
C1171 _117_ net46 5.03e-19
C1172 ctlp[6] _312_/a_193_47# 1.31e-19
C1173 _258_/a_373_47# clknet_2_2__leaf_clk 0.00199f
C1174 _308_/a_805_47# net14 5.85e-19
C1175 _341_/a_193_47# _063_ 1.35e-20
C1176 net12 net11 0.00123f
C1177 net4 _028_ 0.0109f
C1178 net49 _332_/a_27_47# 5.23e-20
C1179 _051_ net3 0.0124f
C1180 VPWR _307_/a_1108_47# 0.0112f
C1181 VPWR _323_/a_1217_47# 1.75e-19
C1182 clknet_2_0__leaf_clk _120_ 0.0431f
C1183 net31 trim_mask\[1\] 4.83e-19
C1184 VPWR _133_ 0.932f
C1185 _053_ state\[1\] 0.0276f
C1186 _314_/a_1217_47# net29 1.37e-19
C1187 net45 rebuffer5/a_161_47# 3.93e-19
C1188 _329_/a_448_47# _026_ 0.00413f
C1189 _329_/a_448_47# VPWR 0.00307f
C1190 result[7] _314_/a_193_47# 0.0012f
C1191 VPWR result[0] 0.162f
C1192 _110_ _271_/a_75_212# 0.00989f
C1193 _305_/a_1108_47# net2 1.43e-20
C1194 net43 _320_/a_651_413# 2.97e-20
C1195 _097_ net15 0.211f
C1196 _335_/a_805_47# _032_ 1.01e-19
C1197 net31 _290_/a_27_413# 0.00589f
C1198 _309_/a_761_289# net14 6.88e-19
C1199 _321_/a_761_289# mask\[3\] 5.12e-21
C1200 _321_/a_543_47# net25 2.89e-20
C1201 _313_/a_1108_47# _155_/a_68_297# 2.65e-19
C1202 _305_/a_27_47# _305_/a_639_47# -0.0015f
C1203 net42 _088_ 0.00164f
C1204 _309_/a_193_47# _309_/a_543_47# -0.0129f
C1205 net12 _209_/a_27_47# 0.0021f
C1206 _042_ _311_/a_27_47# 3.4e-21
C1207 _038_ trim_mask\[4\] 1.02e-19
C1208 net43 _140_/a_68_297# 3.96e-19
C1209 clknet_2_0__leaf_clk _076_ 0.00551f
C1210 _067_ _190_/a_655_47# 6.58e-21
C1211 VPWR _341_/a_1462_47# 6.25e-20
C1212 _065_ rebuffer5/a_161_47# 6.42e-19
C1213 _305_/a_27_47# clknet_2_1__leaf_clk 0.0266f
C1214 net14 net41 0.0116f
C1215 _306_/a_761_289# clknet_2_0__leaf_clk 2.53e-19
C1216 _320_/a_1283_21# net52 2.4e-19
C1217 _306_/a_27_47# net45 1.56e-20
C1218 clknet_2_1__leaf_clk _311_/a_1283_21# 0.00123f
C1219 _313_/a_193_47# _158_/a_68_297# 2.04e-19
C1220 _303_/a_1270_413# clknet_2_3__leaf_clk 3.05e-19
C1221 _269_/a_81_21# _269_/a_384_47# 5.55e-35
C1222 _091_ _092_ 0.115f
C1223 _323_/a_193_47# net19 0.0188f
C1224 _117_ _335_/a_651_413# 1.39e-19
C1225 _305_/a_639_47# net51 3.68e-19
C1226 _327_/a_193_47# _302_/a_27_297# 5.93e-20
C1227 _341_/a_27_47# clknet_2_2__leaf_clk 1.33e-19
C1228 _113_ trim_mask\[1\] 0.0392f
C1229 _030_ trim_val\[1\] 1.15e-19
C1230 _321_/a_193_47# mask\[4\] 2.97e-20
C1231 _067_ trim_val\[4\] 0.00182f
C1232 _274_/a_75_212# clknet_2_2__leaf_clk 3.4e-20
C1233 VPWR _308_/a_805_47# 4.2e-19
C1234 _195_/a_218_374# net30 8.83e-21
C1235 _306_/a_448_47# _072_ 1.94e-20
C1236 _094_ net30 2.27e-19
C1237 trim_mask\[2\] _175_/a_68_297# 0.00261f
C1238 _337_/a_1283_21# _092_ 7.91e-20
C1239 _337_/a_1108_47# _099_ 2.94e-21
C1240 VPWR net14 1.08f
C1241 net3 _316_/a_1283_21# 0.00391f
C1242 trim_mask\[2\] _333_/a_193_47# 2.63e-20
C1243 cal_count\[1\] _339_/a_27_47# 9.04e-22
C1244 net44 _209_/a_27_47# 0.00315f
C1245 net45 sample 4.04e-20
C1246 clknet_2_1__leaf_clk net51 0.331f
C1247 _088_ _054_ 0.0123f
C1248 _167_/a_161_47# _099_ 4.06e-21
C1249 _306_/a_27_47# _065_ 9.37e-21
C1250 net16 _334_/a_1270_413# 1.15e-20
C1251 _088_ net30 2.51e-19
C1252 net26 _310_/a_1108_47# 1.19e-19
C1253 clkbuf_0_clk/a_110_47# _190_/a_27_47# 0.012f
C1254 rebuffer3/a_75_212# net40 0.0347f
C1255 VPWR _237_/a_439_47# -2.74e-19
C1256 _058_ _302_/a_27_297# 0.00216f
C1257 VPWR _309_/a_761_289# -4.42e-20
C1258 _116_ fanout46/a_27_47# 9.48e-21
C1259 en_co_clk _243_/a_27_297# 0.00177f
C1260 _328_/a_193_47# net46 -2.55e-20
C1261 _253_/a_299_297# net25 5.91e-19
C1262 output28/a_27_47# result[6] 0.00425f
C1263 calibrate _317_/a_27_47# 4.43e-22
C1264 VPWR _339_/a_1140_413# -3.83e-19
C1265 net9 net46 1.8f
C1266 _104_ _336_/a_1108_47# 0.0578f
C1267 net54 _337_/a_761_289# 1.02e-19
C1268 _058_ _106_ 5.05e-19
C1269 _324_/a_543_47# net53 8.7e-19
C1270 _290_/a_27_413# net2 5.47e-21
C1271 _019_ _320_/a_761_289# 1.17e-19
C1272 _094_ net22 0.00156f
C1273 _169_/a_215_311# _167_/a_161_47# 7.46e-19
C1274 net31 output33/a_27_47# 0.00225f
C1275 VPWR _040_ 0.121f
C1276 VPWR net41 0.334f
C1277 _065_ net40 1.05e-19
C1278 net13 _322_/a_651_413# 0.00105f
C1279 _300_/a_47_47# net16 2.14e-19
C1280 _247_/a_27_297# _018_ 0.00761f
C1281 VPWR _292_/a_78_199# 0.0154f
C1282 trim_mask\[2\] trim_mask\[4\] 0.014f
C1283 _146_/a_68_297# net29 1.71e-20
C1284 _337_/a_1270_413# _034_ 1.66e-20
C1285 net23 net14 0.00709f
C1286 net48 _108_ 0.00159f
C1287 net49 _332_/a_1217_47# 3.38e-20
C1288 VPWR _324_/a_1108_47# 0.0164f
C1289 clknet_0_clk net19 0.0411f
C1290 _322_/a_761_289# net53 4.45e-21
C1291 _110_ _269_/a_384_47# 1.12e-19
C1292 _301_/a_47_47# trim_val\[0\] 2.33e-21
C1293 _026_ VPWR 0.0678f
C1294 _309_/a_1108_47# net43 -0.0159f
C1295 _304_/a_193_47# en_co_clk 2.08e-20
C1296 _108_ _054_ 1.4e-20
C1297 mask\[0\] _137_/a_150_297# 0.00141f
C1298 _327_/a_193_47# trim_mask\[0\] 0.0048f
C1299 _053_ _304_/a_1108_47# 7.74e-19
C1300 net4 _279_/a_314_297# 0.00558f
C1301 _257_/a_109_297# _119_ 1.08e-19
C1302 net30 _108_ 0.0409f
C1303 _107_ _098_ 0.0442f
C1304 cal_itt\[0\] _068_ 0.0453f
C1305 _305_/a_543_47# _002_ 0.0363f
C1306 net16 _332_/a_1108_47# 0.0106f
C1307 _277_/a_75_212# _335_/a_193_47# 0.00452f
C1308 VPWR _322_/a_1283_21# 0.0587f
C1309 net9 _300_/a_377_297# 5.89e-20
C1310 net16 _029_ 4.6e-19
C1311 VPWR _331_/a_1283_21# 0.0453f
C1312 _329_/a_27_47# trim_mask\[4\] 4.49e-19
C1313 _329_/a_1108_47# clknet_2_2__leaf_clk 0.00393f
C1314 _314_/a_761_289# _011_ 7.65e-19
C1315 net52 net14 2.19e-20
C1316 _311_/a_651_413# net26 0.0265f
C1317 _232_/a_32_297# _232_/a_114_297# -5.24e-19
C1318 net23 _040_ 0.0416f
C1319 net43 result[6] 7.22e-20
C1320 _309_/a_1283_21# _101_ 8.96e-19
C1321 _322_/a_193_47# _322_/a_651_413# -0.00399f
C1322 trim_mask\[0\] _058_ 0.142f
C1323 _064_ _256_/a_109_47# 0.00199f
C1324 _104_ _256_/a_27_297# 0.0651f
C1325 clknet_0_clk _107_ 0.039f
C1326 _324_/a_193_47# _312_/a_193_47# 7.32e-21
C1327 _250_/a_109_297# clknet_2_1__leaf_clk 9.25e-19
C1328 result[7] _074_ 1.76e-20
C1329 _093_ _049_ 0.0933f
C1330 VPWR _303_/a_805_47# 2.3e-19
C1331 trim_val\[1\] trim_mask\[1\] 0.163f
C1332 _074_ net30 0.0754f
C1333 _185_/a_150_297# _316_/a_193_47# 1.56e-20
C1334 _328_/a_1283_21# _108_ 5.16e-21
C1335 _245_/a_109_297# _101_ 9.95e-19
C1336 _327_/a_1283_21# _136_ 0.00212f
C1337 _327_/a_27_47# _038_ 2.98e-20
C1338 net15 _319_/a_193_47# 0.0179f
C1339 net48 _031_ 0.00259f
C1340 net9 _332_/a_448_47# 7.31e-20
C1341 _305_/a_761_289# _203_/a_59_75# 1.9e-20
C1342 _086_ _310_/a_27_47# 3.93e-22
C1343 VPWR net23 0.425f
C1344 _040_ net52 0.153f
C1345 _308_/a_761_289# _080_ 4.22e-19
C1346 result[4] _253_/a_81_21# 9.76e-20
C1347 _101_ net53 0.0928f
C1348 cal_itt\[2\] _305_/a_543_47# 9.12e-20
C1349 net37 cal_count\[2\] 1.17e-19
C1350 _128_ _339_/a_1224_47# 1.82e-19
C1351 _329_/a_651_413# trim_mask\[3\] 6.01e-19
C1352 _066_ _278_/a_27_47# 3.47e-20
C1353 _194_/a_113_297# net40 6.94e-19
C1354 _336_/a_1283_21# net40 3.24e-21
C1355 _059_ _100_ 0.0368f
C1356 net12 _044_ 4.19e-20
C1357 _074_ net22 0.191f
C1358 _303_/a_543_47# _000_ 0.00206f
C1359 _328_/a_1462_47# net46 0.00138f
C1360 _110_ _117_ 0.0388f
C1361 _313_/a_193_47# _084_ 3.03e-21
C1362 VPWR net52 0.583f
C1363 _337_/a_27_47# _120_ 6.92e-19
C1364 _337_/a_193_47# en_co_clk 0.0291f
C1365 _303_/a_27_47# net19 0.015f
C1366 VPWR _063_ 1.06f
C1367 _292_/a_78_199# _036_ 0.00115f
C1368 clkbuf_2_0__f_clk/a_110_47# _192_/a_27_47# 4.09e-20
C1369 _164_/a_161_47# net41 1.53e-19
C1370 input1/a_75_212# _316_/a_193_47# 1.11e-19
C1371 _015_ _316_/a_193_47# 7.75e-21
C1372 _328_/a_1108_47# _030_ 0.00135f
C1373 _270_/a_59_75# _332_/a_193_47# 1.72e-20
C1374 output8/a_27_47# net46 8.79e-19
C1375 VPWR _036_ 0.808f
C1376 net31 _270_/a_59_75# 2.36e-20
C1377 _097_ _012_ 7.01e-20
C1378 _321_/a_651_413# mask\[2\] 1.94e-19
C1379 _337_/a_27_47# _076_ 8.74e-20
C1380 net44 _044_ 9.19e-19
C1381 VPWR _164_/a_161_47# 0.0878f
C1382 _303_/a_805_47# _063_ 6.23e-21
C1383 net8 _334_/a_1108_47# 0.0184f
C1384 _078_ _247_/a_27_297# 0.0114f
C1385 _327_/a_1462_47# trim_mask\[0\] 5.41e-21
C1386 _280_/a_75_212# clknet_2_2__leaf_clk 0.0284f
C1387 output23/a_27_47# net22 6.71e-20
C1388 net23 net52 0.00459f
C1389 net2 _078_ 6.06e-20
C1390 _251_/a_27_297# mask\[6\] 0.0749f
C1391 mask\[6\] _250_/a_109_47# 0.00348f
C1392 _312_/a_448_47# net20 0.0146f
C1393 VPWR _260_/a_346_47# -9.01e-19
C1394 _100_ _075_ 1.35e-20
C1395 _008_ _101_ 0.00877f
C1396 _312_/a_448_47# net53 7.79e-20
C1397 _308_/a_27_47# mask\[1\] 3.15e-20
C1398 _074_ _315_/a_651_413# 0.00346f
C1399 _012_ _315_/a_543_47# 0.00477f
C1400 calibrate _315_/a_448_47# 8.06e-19
C1401 _064_ _258_/a_109_297# 1.38e-21
C1402 _259_/a_27_297# trim_mask\[2\] 9.79e-20
C1403 _239_/a_694_21# net42 1.79e-19
C1404 _331_/a_761_289# _028_ 0.0322f
C1405 _331_/a_543_47# clknet_2_2__leaf_clk 3.85e-19
C1406 _113_ _270_/a_59_75# 0.00141f
C1407 _021_ clknet_2_1__leaf_clk 0.143f
C1408 _281_/a_103_199# _316_/a_1283_21# 4.66e-21
C1409 _331_/a_651_413# _260_/a_93_21# 9.66e-21
C1410 VPWR _083_ 0.0607f
C1411 state\[0\] clk 2.86e-19
C1412 _317_/a_27_47# _317_/a_1108_47# -2.98e-20
C1413 _317_/a_193_47# _317_/a_1283_21# -5.93e-19
C1414 _060_ _316_/a_1108_47# 1.92e-20
C1415 net48 net49 0.00261f
C1416 mask\[1\] clknet_0_clk 1.17e-19
C1417 _101_ _016_ 0.0161f
C1418 _272_/a_384_47# trim_val\[2\] 3.41e-19
C1419 _272_/a_81_21# net48 0.00492f
C1420 _143_/a_150_297# mask\[2\] 3.43e-19
C1421 net33 rebuffer1/a_75_212# 5.32e-20
C1422 net15 _319_/a_1462_47# 6.83e-20
C1423 _110_ _328_/a_193_47# 4.66e-20
C1424 _320_/a_1108_47# mask\[1\] 0.0533f
C1425 output32/a_27_47# clkc 4.89e-21
C1426 _276_/a_59_75# _277_/a_75_212# 0.0157f
C1427 _305_/a_448_47# _072_ 2.59e-19
C1428 _322_/a_1283_21# _083_ 4.82e-19
C1429 net31 _056_ 9.97e-20
C1430 _321_/a_543_47# net15 0.00541f
C1431 _110_ net9 0.138f
C1432 clkbuf_2_0__f_clk/a_110_47# clknet_2_0__leaf_clk 0.208f
C1433 trim[4] _047_ 0.0025f
C1434 net45 net51 1.03e-19
C1435 _005_ _213_/a_109_297# 0.00125f
C1436 _290_/a_207_413# _127_ 0.0186f
C1437 _305_/a_27_47# _065_ 8.53e-20
C1438 _259_/a_27_297# _329_/a_27_47# 7.3e-21
C1439 _065_ _311_/a_1283_21# 2.03e-21
C1440 _235_/a_297_47# _337_/a_193_47# 6.67e-21
C1441 _235_/a_79_21# _337_/a_543_47# 1.39e-19
C1442 _313_/a_193_47# _085_ 0.0013f
C1443 net21 _312_/a_193_47# 2.49e-21
C1444 VPWR net50 0.269f
C1445 trim_mask\[0\] en_co_clk 4.6e-20
C1446 cal_itt\[0\] _042_ 1.18e-20
C1447 _323_/a_1283_21# mask\[4\] 0.0627f
C1448 net30 _170_/a_299_297# 8.72e-20
C1449 _171_/a_27_47# _049_ 0.00707f
C1450 state\[0\] net4 0.0129f
C1451 output10/a_27_47# _275_/a_81_21# 8.07e-20
C1452 _306_/a_27_47# clkbuf_0_clk/a_110_47# 1.17e-20
C1453 _187_/a_212_413# clkc 7.77e-19
C1454 clkbuf_2_3__f_clk/a_110_47# _092_ 0.00248f
C1455 _239_/a_277_297# _049_ 0.0076f
C1456 input2/a_27_47# net34 0.00866f
C1457 _093_ state\[1\] 3.64e-20
C1458 _340_/a_1032_413# net40 8.48e-21
C1459 _337_/a_1462_47# en_co_clk 5.11e-19
C1460 _303_/a_1217_47# net19 1.84e-19
C1461 _312_/a_27_47# _312_/a_1108_47# -2.98e-20
C1462 _074_ _079_ 0.0205f
C1463 _328_/a_1108_47# trim_mask\[1\] 0.048f
C1464 _336_/a_448_47# net46 1.09e-21
C1465 _065_ net51 0.0819f
C1466 net31 clkc 0.146f
C1467 trim_mask\[2\] _178_/a_68_297# 4.08e-20
C1468 VPWR _333_/a_448_47# 0.018f
C1469 _090_ _242_/a_79_21# 1.33e-20
C1470 _019_ _101_ 0.0724f
C1471 clknet_0_clk _118_ 2.72e-21
C1472 _002_ net30 0.00184f
C1473 fanout45/a_27_47# net15 0.00307f
C1474 _128_ _291_/a_285_297# 7.1e-19
C1475 _078_ net29 0.109f
C1476 _290_/a_207_413# _126_ 0.0121f
C1477 _200_/a_80_21# _071_ 0.00109f
C1478 net44 _208_/a_505_21# 2.17e-19
C1479 output32/a_27_47# _173_/a_27_47# 5.36e-21
C1480 net2 fanout47/a_27_47# 5.94e-20
C1481 _023_ result[5] 8.38e-19
C1482 _051_ _076_ 8.68e-19
C1483 net44 mask\[2\] 0.00622f
C1484 _326_/a_27_47# _253_/a_81_21# 1.02e-19
C1485 _319_/a_1108_47# _244_/a_27_297# 4.17e-20
C1486 net28 _155_/a_68_297# 0.00694f
C1487 _064_ clkbuf_2_2__f_clk/a_110_47# 2.53e-20
C1488 _304_/a_193_47# cal_count\[0\] 7.48e-20
C1489 _304_/a_543_47# _124_ 8.48e-20
C1490 _162_/a_27_47# net37 0.0246f
C1491 clknet_2_1__leaf_clk _086_ 0.00107f
C1492 VPWR _217_/a_109_297# -0.00161f
C1493 _237_/a_505_21# _092_ 3.2e-21
C1494 _237_/a_218_374# _099_ 2.1e-19
C1495 _005_ _212_/a_113_297# 6.78e-19
C1496 _192_/a_505_280# _049_ 9.03e-19
C1497 net50 _063_ 2.42e-20
C1498 VPWR _155_/a_150_297# -5.53e-19
C1499 _322_/a_761_289# _205_/a_27_47# 0.00152f
C1500 _289_/a_68_297# _126_ 6.69e-19
C1501 cal_itt\[2\] net30 0.00218f
C1502 _321_/a_27_47# _310_/a_1283_21# 5.37e-21
C1503 output9/a_27_47# ctln[3] 0.00992f
C1504 _042_ clknet_2_0__leaf_clk 1.44e-20
C1505 _331_/a_639_47# trim_mask\[4\] 2.12e-19
C1506 net31 _173_/a_27_47# 0.00232f
C1507 VPWR _279_/a_396_47# 0.0215f
C1508 _256_/a_109_297# net46 2.51e-20
C1509 _028_ _260_/a_250_297# 4.5e-19
C1510 _306_/a_27_47# _204_/a_75_212# 0.00414f
C1511 _327_/a_543_47# clknet_2_3__leaf_clk 1.94e-19
C1512 VPWR _325_/a_448_47# 0.00338f
C1513 net13 _099_ 0.00749f
C1514 net4 _330_/a_1108_47# 9.85e-20
C1515 VPWR _216_/a_113_297# 0.0761f
C1516 _317_/a_27_47# clknet_2_0__leaf_clk 0.0895f
C1517 _002_ _072_ 0.0995f
C1518 _066_ _108_ 0.0118f
C1519 _263_/a_79_21# _107_ 0.00791f
C1520 _053_ clkbuf_2_2__f_clk/a_110_47# 4.79e-19
C1521 net26 _072_ 1.07e-20
C1522 _248_/a_27_297# net53 0.06f
C1523 mask\[1\] _245_/a_27_297# 0.0144f
C1524 net2 clkc 3.18e-19
C1525 _038_ net40 2.03e-19
C1526 fanout46/a_27_47# _336_/a_1108_47# 0.00191f
C1527 _048_ _242_/a_79_21# 0.0352f
C1528 _325_/a_193_47# _046_ 6.44e-20
C1529 net15 _282_/a_150_297# 1.95e-19
C1530 _104_ _329_/a_193_47# 5.06e-20
C1531 net46 net32 2.32e-19
C1532 VPWR _181_/a_150_297# -4.93e-19
C1533 clknet_2_2__leaf_clk net19 0.125f
C1534 _327_/a_805_47# net18 2.75e-19
C1535 _094_ _337_/a_651_413# 8.78e-22
C1536 net13 _169_/a_215_311# 0.0132f
C1537 _333_/a_27_47# _333_/a_193_47# -0.0618f
C1538 _035_ _124_ 0.003f
C1539 _069_ _068_ 1.84e-20
C1540 net5 _135_ 1.05e-19
C1541 input2/a_27_47# _133_ 1.69e-19
C1542 cal_count\[3\] _092_ 0.0602f
C1543 net10 trim_mask\[3\] 0.00217f
C1544 VPWR _248_/a_109_47# -6.03e-19
C1545 _265_/a_81_21# _333_/a_27_47# 8.6e-21
C1546 output25/a_27_47# net25 0.0216f
C1547 _254_/a_109_297# wire42/a_75_212# 6.01e-20
C1548 net12 _306_/a_448_47# 0.00883f
C1549 trim_mask\[3\] clknet_2_2__leaf_clk 0.0111f
C1550 _203_/a_59_75# cal_itt\[3\] 0.0588f
C1551 net3 _263_/a_297_47# 2.03e-19
C1552 _325_/a_639_47# net43 2.23e-19
C1553 _033_ net46 0.175f
C1554 _104_ net18 0.0279f
C1555 net19 net11 0.00896f
C1556 input1/a_75_212# net14 0.00531f
C1557 trim_val\[1\] _056_ 5.31e-19
C1558 _101_ _205_/a_27_47# 0.0103f
C1559 _320_/a_543_47# mask\[2\] 3.55e-19
C1560 _320_/a_27_47# _017_ 0.25f
C1561 _134_ comp 1.07e-19
C1562 cal_itt\[2\] _072_ 0.145f
C1563 cal_itt\[0\] cal_itt\[3\] 0.00179f
C1564 trim[1] _162_/a_27_47# 6.46e-19
C1565 VPWR _185_/a_150_297# 2.07e-19
C1566 net13 _246_/a_27_297# 1.03e-19
C1567 _107_ clknet_2_2__leaf_clk 0.00487f
C1568 _107_ _260_/a_584_47# 7.02e-20
C1569 net43 _158_/a_68_297# 3.83e-20
C1570 _288_/a_59_75# trimb[4] 2.54e-20
C1571 _303_/a_543_47# mask\[4\] 0.0017f
C1572 _333_/a_1108_47# clknet_2_2__leaf_clk 2.36e-21
C1573 clknet_2_1__leaf_clk _319_/a_761_289# 1.4e-19
C1574 _014_ _049_ 1.21e-21
C1575 comp _130_ 9.2e-19
C1576 _308_/a_1283_21# fanout43/a_27_47# 0.00444f
C1577 _063_ _279_/a_396_47# 2.43e-20
C1578 _318_/a_193_47# net45 -9.53e-19
C1579 _325_/a_448_47# net52 1.96e-20
C1580 _325_/a_1270_413# _101_ 1.05e-20
C1581 _324_/a_1283_21# _044_ 5.4e-19
C1582 _189_/a_27_47# net55 8.85e-21
C1583 _306_/a_448_47# net44 3.68e-19
C1584 input3/a_75_212# net3 0.00197f
C1585 _326_/a_761_289# _023_ 8.7e-19
C1586 _326_/a_543_47# _102_ 1.05e-19
C1587 _326_/a_1283_21# mask\[7\] 0.019f
C1588 ctlp[7] _074_ 0.0518f
C1589 _341_/a_1108_47# en_co_clk 1.08e-19
C1590 _050_ _090_ 0.0666f
C1591 VPWR _034_ 0.275f
C1592 _249_/a_373_47# net53 0.00136f
C1593 _015_ net41 0.00932f
C1594 cal output41/a_27_47# 0.0251f
C1595 input1/a_75_212# net41 0.0639f
C1596 output39/a_27_47# net16 0.00133f
C1597 clkbuf_2_2__f_clk/a_110_47# _330_/a_448_47# 8.5e-19
C1598 _286_/a_76_199# _338_/a_652_21# 1.79e-19
C1599 _047_ _108_ 0.00591f
C1600 _324_/a_193_47# mask\[5\] 4.16e-19
C1601 VPWR output26/a_27_47# 0.094f
C1602 _340_/a_1182_261# cal_count\[0\] 1.02e-20
C1603 net12 _094_ 1.21e-20
C1604 mask\[0\] _078_ 0.0857f
C1605 trim[0] _047_ 5.54e-19
C1606 clk _052_ 0.0283f
C1607 _187_/a_212_413# _136_ 1.66e-19
C1608 _340_/a_193_47# net2 1.9e-19
C1609 _052_ clone7/a_27_47# 2.83e-37
C1610 net12 _088_ 3.71e-19
C1611 _024_ net46 0.0198f
C1612 _015_ VPWR 0.242f
C1613 VPWR input1/a_75_212# 0.0681f
C1614 _306_/a_448_47# _003_ 0.00243f
C1615 VPWR _327_/a_1108_47# 0.0204f
C1616 _141_/a_27_47# _040_ 0.0116f
C1617 _136_ _332_/a_193_47# 0.00381f
C1618 _317_/a_805_47# _014_ 3.81e-19
C1619 _317_/a_448_47# state\[1\] 7.84e-20
C1620 net31 _172_/a_68_297# 0.0148f
C1621 output22/a_27_47# sample 4.4e-21
C1622 result[0] output30/a_27_47# 0.00176f
C1623 _074_ _313_/a_543_47# 2.34e-20
C1624 _232_/a_32_297# _096_ 0.0796f
C1625 _315_/a_193_47# _315_/a_1108_47# -0.00656f
C1626 state\[2\] _331_/a_27_47# 1.55e-21
C1627 _312_/a_1283_21# _152_/a_68_297# 3.24e-19
C1628 net4 _195_/a_535_374# 2.01e-19
C1629 _167_/a_161_47# _093_ 2.98e-20
C1630 _325_/a_1283_21# _019_ 9.46e-20
C1631 _322_/a_639_47# mask\[3\] 2.74e-19
C1632 _287_/a_75_212# _123_ 2.48e-19
C1633 trim_mask\[2\] _334_/a_27_47# 0.00247f
C1634 _125_ net38 1.01e-19
C1635 net13 _084_ 5.3e-20
C1636 net4 _052_ 8.16e-20
C1637 _094_ net44 0.14f
C1638 net13 _053_ 5.12e-19
C1639 _305_/a_27_47# clkbuf_0_clk/a_110_47# 7.19e-20
C1640 VPWR _141_/a_27_47# 0.0633f
C1641 _125_ _339_/a_1182_261# 9.71e-21
C1642 net9 _065_ 3.57e-20
C1643 _312_/a_193_47# _045_ 3.32e-19
C1644 _243_/a_27_297# _049_ 6.11e-19
C1645 _325_/a_27_47# _325_/a_193_47# -0.0524f
C1646 trim_val\[0\] _333_/a_1108_47# 2.64e-21
C1647 VPWR input2/a_27_47# 0.171f
C1648 trim_val\[1\] _173_/a_27_47# 0.1f
C1649 net19 _279_/a_204_297# 3.29e-19
C1650 _064_ _257_/a_109_297# 0.00587f
C1651 _265_/a_299_297# _109_ 0.00133f
C1652 _050_ _048_ 0.117f
C1653 _019_ _248_/a_27_297# 0.00879f
C1654 _062_ _098_ 3.97e-19
C1655 _334_/a_1108_47# net34 0.00409f
C1656 _114_ _056_ 1.67e-19
C1657 _227_/a_109_93# net55 0.0174f
C1658 _102_ _310_/a_1108_47# 0.00168f
C1659 VPWR _281_/a_253_47# -6.1e-19
C1660 _040_ _208_/a_76_199# 1.12e-19
C1661 _262_/a_27_47# wire42/a_75_212# 3.51e-19
C1662 _225_/a_109_297# _011_ 0.00438f
C1663 net45 _315_/a_1283_21# 0.0662f
C1664 _014_ _315_/a_1108_47# 3.11e-19
C1665 clknet_2_0__leaf_clk _315_/a_448_47# 0.00154f
C1666 output36/a_27_47# _126_ 2.66e-19
C1667 _321_/a_27_47# _042_ 0.106f
C1668 _218_/a_199_47# mask\[4\] 0.00145f
C1669 _053_ _198_/a_27_47# 3.78e-20
C1670 clknet_0_clk _062_ 0.142f
C1671 _061_ trim_mask\[0\] 5.78e-19
C1672 _050_ trim_mask\[4\] 0.228f
C1673 _103_ _262_/a_109_297# 1.2e-19
C1674 _107_ _279_/a_204_297# 0.00129f
C1675 _053_ _331_/a_193_47# 1.48e-22
C1676 _321_/a_1283_21# clknet_2_1__leaf_clk 0.0101f
C1677 clk calibrate 6.08e-20
C1678 _336_/a_193_47# net30 5.93e-22
C1679 trim_mask\[0\] _332_/a_639_47# 0.00131f
C1680 _115_ _334_/a_27_47# 0.00138f
C1681 VPWR _193_/a_109_297# -7.56e-19
C1682 calibrate clone7/a_27_47# 0.0232f
C1683 net12 _074_ 4.02e-19
C1684 _339_/a_1182_261# net40 4.04e-20
C1685 VPWR _208_/a_76_199# 0.0151f
C1686 _340_/a_193_47# _123_ 0.0182f
C1687 _136_ net2 0.0141f
C1688 clknet_2_1__leaf_clk _313_/a_27_47# 0.617f
C1689 _060_ _089_ 3.49e-19
C1690 clkbuf_2_2__f_clk/a_110_47# _027_ 0.0137f
C1691 _041_ _124_ 0.112f
C1692 cal_count\[0\] _338_/a_652_21# 2.2e-20
C1693 _242_/a_297_47# _092_ 2.32e-20
C1694 _324_/a_1462_47# mask\[5\] 6.42e-19
C1695 net20 _156_/a_27_47# 0.00307f
C1696 net44 _244_/a_27_297# 0.0642f
C1697 _234_/a_109_297# _065_ 2.4e-19
C1698 _168_/a_207_413# _336_/a_27_47# 3.37e-21
C1699 net42 net55 0.0904f
C1700 _141_/a_27_47# net52 0.0406f
C1701 clknet_0_clk _195_/a_76_199# 1.29e-19
C1702 _237_/a_76_199# net15 0.00477f
C1703 _015_ _164_/a_161_47# 0.0142f
C1704 _328_/a_27_47# _336_/a_1108_47# 3.63e-20
C1705 _322_/a_543_47# mask\[2\] 7.1e-19
C1706 _110_ net32 4.19e-20
C1707 calibrate net4 2.6e-19
C1708 _004_ mask\[0\] 8.96e-20
C1709 _014_ state\[1\] 1.65e-20
C1710 net13 _085_ 6.8e-21
C1711 VPWR output30/a_27_47# 0.0452f
C1712 net54 _242_/a_79_21# 1.39e-19
C1713 _074_ net44 0.137f
C1714 VPWR _278_/a_109_297# -1.67e-19
C1715 mask\[1\] _209_/a_27_47# 0.00518f
C1716 _301_/a_47_47# _108_ 1.67e-20
C1717 _301_/a_47_47# _332_/a_543_47# 1.61e-20
C1718 clknet_2_2__leaf_clk _118_ 2.09e-19
C1719 result[5] result[6] 0.035f
C1720 net19 _044_ 0.00728f
C1721 ctlp[2] trimb[3] 0.00996f
C1722 _327_/a_1283_21# clknet_2_2__leaf_clk 0.00475f
C1723 trim_mask\[2\] _271_/a_75_212# 8.82e-19
C1724 _119_ _330_/a_27_47# 8.06e-19
C1725 _341_/a_27_47# _108_ 5.19e-20
C1726 _319_/a_805_47# _049_ 2.4e-20
C1727 _244_/a_27_297# _003_ 9.28e-20
C1728 _110_ _033_ 0.00853f
C1729 _047_ net49 4.23e-21
C1730 _000_ mask\[5\] 1.37e-19
C1731 VPWR _330_/a_543_47# 0.0134f
C1732 _329_/a_543_47# _027_ 1.42e-20
C1733 _329_/a_761_289# net46 1.16e-19
C1734 _125_ _339_/a_1296_47# 7.89e-21
C1735 _339_/a_27_47# _286_/a_535_374# 7e-20
C1736 net37 _129_ 1.3e-19
C1737 net55 _054_ 4.54e-20
C1738 _275_/a_299_297# _178_/a_150_297# 8.01e-20
C1739 _059_ net41 0.127f
C1740 mask\[5\] _312_/a_1283_21# 5.46e-20
C1741 net12 _305_/a_448_47# 2.34e-19
C1742 _323_/a_543_47# _068_ 6.22e-19
C1743 _307_/a_1283_21# _094_ 8.61e-21
C1744 net55 net30 0.0559f
C1745 net3 _099_ 0.0116f
C1746 _337_/a_193_47# _049_ 0.0219f
C1747 _064_ _025_ 6.73e-20
C1748 cal_itt\[1\] _304_/a_1108_47# 7.9e-19
C1749 _200_/a_209_47# _106_ 1.13e-19
C1750 output14/a_27_47# net28 0.0464f
C1751 _134_ net46 6.57e-20
C1752 trim_val\[1\] _172_/a_68_297# 0.0814f
C1753 _314_/a_27_47# net14 0.00552f
C1754 net52 _208_/a_76_199# 0.00104f
C1755 _341_/a_1270_413# net46 -3.58e-20
C1756 _168_/a_27_413# net55 2.98e-20
C1757 _146_/a_68_297# _081_ 1.07e-20
C1758 net27 _046_ 0.0365f
C1759 VPWR _059_ 0.389f
C1760 state\[2\] _242_/a_297_47# 0.00228f
C1761 _328_/a_27_47# _256_/a_27_297# 0.0111f
C1762 _321_/a_27_47# _022_ 7.92e-21
C1763 output34/a_27_47# trim[3] 0.00978f
C1764 _169_/a_215_311# net3 5.43e-20
C1765 _046_ _222_/a_113_297# 0.0555f
C1766 _188_/a_27_47# _131_ 7.53e-22
C1767 _136_ _123_ 5.71e-19
C1768 _319_/a_1283_21# clknet_2_0__leaf_clk 0.0582f
C1769 _319_/a_761_289# net45 7.31e-20
C1770 _321_/a_1217_47# _042_ 1.61e-19
C1771 _339_/a_1032_413# net37 4.63e-21
C1772 _305_/a_448_47# net44 0.00192f
C1773 mask\[6\] _313_/a_193_47# 1.19e-20
C1774 _200_/a_209_297# clkbuf_0_clk/a_110_47# 6.87e-20
C1775 net44 _311_/a_805_47# -0.001f
C1776 net27 _312_/a_761_289# 3.47e-19
C1777 state\[1\] _243_/a_27_297# 3.97e-19
C1778 _053_ _260_/a_93_21# 0.00615f
C1779 _106_ _049_ 2e-20
C1780 _274_/a_75_212# _031_ 0.00317f
C1781 clkbuf_2_1__f_clk/a_110_47# _121_ 5.11e-19
C1782 _110_ _024_ 1.51e-21
C1783 net43 _085_ 0.00429f
C1784 mask\[7\] net29 1.03f
C1785 _340_/a_1182_261# net16 7.99e-19
C1786 output10/a_27_47# _057_ 4.11e-19
C1787 _124_ net18 0.022f
C1788 cal_count\[0\] _338_/a_1056_47# 4.68e-20
C1789 VPWR _306_/a_1108_47# 0.0189f
C1790 _327_/a_1283_21# trim_val\[0\] 2.3e-20
C1791 _312_/a_1108_47# _084_ 1.83e-20
C1792 _135_ _122_ 2.59e-19
C1793 _188_/a_27_47# net5 0.00215f
C1794 _187_/a_27_413# clknet_2_3__leaf_clk 0.00665f
C1795 _241_/a_105_352# _092_ 9.7e-21
C1796 _241_/a_388_297# _099_ 0.00252f
C1797 _241_/a_297_47# _095_ 0.00293f
C1798 _341_/a_761_289# net2 1.57e-22
C1799 VPWR _314_/a_27_47# 0.0448f
C1800 _293_/a_384_47# _126_ 2.2e-20
C1801 _058_ _333_/a_805_47# 2.61e-19
C1802 cal en 0.0365f
C1803 net47 net26 0.00334f
C1804 _218_/a_113_297# _076_ 5.93e-20
C1805 _058_ _109_ 0.0221f
C1806 VPWR _075_ 0.187f
C1807 net33 _131_ 0.00541f
C1808 _262_/a_465_47# net55 2.93e-19
C1809 mask\[7\] _251_/a_373_47# -2.76e-19
C1810 net8 _056_ 0.00123f
C1811 net12 _239_/a_694_21# 0.0098f
C1812 net9 _340_/a_1032_413# 0.00332f
C1813 _319_/a_27_47# _319_/a_761_289# -0.0166f
C1814 _007_ net25 0.0825f
C1815 _104_ _048_ 0.0872f
C1816 _067_ _072_ 0.0109f
C1817 _072_ _070_ 0.00384f
C1818 trim_mask\[0\] _049_ 0.00997f
C1819 cal_count\[3\] net46 0.0785f
C1820 _279_/a_204_297# _118_ 0.00873f
C1821 _189_/a_218_47# _098_ 9.31e-21
C1822 _339_/a_476_47# cal_count\[0\] 0.0503f
C1823 net2 clknet_0_clk 1.8e-20
C1824 _008_ _077_ 1.23e-20
C1825 _065_ _202_/a_382_297# 0.00191f
C1826 net12 _002_ 4.08e-19
C1827 trim_mask\[0\] net16 0.0753f
C1828 _097_ fanout45/a_27_47# 2.22e-19
C1829 _032_ clkbuf_2_2__f_clk/a_110_47# 1.45e-19
C1830 net25 mask\[3\] 0.0723f
C1831 _305_/a_1283_21# clknet_0_clk 0.00155f
C1832 net54 _050_ 2.65e-19
C1833 net12 net26 0.102f
C1834 _294_/a_150_297# net33 3.68e-19
C1835 net43 _314_/a_543_47# 0.00373f
C1836 _304_/a_1283_21# _065_ 0.00232f
C1837 _337_/a_1462_47# _049_ 4.02e-19
C1838 clk _317_/a_1108_47# 0.00521f
C1839 _317_/a_27_47# _316_/a_1283_21# 4.57e-20
C1840 _317_/a_193_47# _316_/a_543_47# 2.29e-20
C1841 _104_ trim_mask\[4\] 0.215f
C1842 net2 _339_/a_27_47# 1.57e-19
C1843 VPWR _195_/a_505_21# 0.0498f
C1844 net5 net33 3.09e-19
C1845 _257_/a_27_297# net46 1.93e-20
C1846 _028_ _330_/a_193_47# 2e-19
C1847 clknet_2_2__leaf_clk _330_/a_761_289# 0.0325f
C1848 _331_/a_193_47# _027_ 1.93e-19
C1849 trim_mask\[1\] net34 5.19e-20
C1850 _314_/a_1217_47# net14 1.84e-19
C1851 VPWR _326_/a_1108_47# 0.0412f
C1852 _112_ _055_ -1.01e-24
C1853 _329_/a_1108_47# _031_ 8.91e-19
C1854 VPWR _334_/a_1108_47# 0.0162f
C1855 _189_/a_218_47# clknet_0_clk 0.0521f
C1856 _290_/a_27_413# net34 0.0108f
C1857 _306_/a_651_413# _101_ 7.37e-21
C1858 VPWR _295_/a_113_47# 3.07e-19
C1859 _306_/a_1108_47# _063_ 9.17e-21
C1860 output25/a_27_47# _310_/a_193_47# 2.18e-19
C1861 _231_/a_161_47# _278_/a_27_47# 3.92e-20
C1862 _320_/a_27_47# clknet_2_1__leaf_clk 0.00248f
C1863 clk _203_/a_59_75# 0.0113f
C1864 _320_/a_448_47# clkbuf_2_1__f_clk/a_110_47# 9.72e-19
C1865 _053_ net3 1.05e-20
C1866 _331_/a_543_47# _088_ 1.96e-21
C1867 _238_/a_75_212# _316_/a_27_47# 9.84e-19
C1868 VPWR _286_/a_218_47# -3.98e-19
C1869 _340_/a_1032_413# _132_ 6.76e-20
C1870 _325_/a_27_47# net27 1.97e-20
C1871 _002_ net44 0.0123f
C1872 _235_/a_79_21# _090_ 0.001f
C1873 net15 _090_ 7.61e-19
C1874 cal_itt\[0\] clk 7.41e-21
C1875 net4 _317_/a_1108_47# 0.0157f
C1876 _308_/a_639_47# _074_ 0.00194f
C1877 net44 net26 0.0738f
C1878 VPWR _137_/a_150_297# 3.84e-19
C1879 _335_/a_27_47# _119_ 1.68e-19
C1880 _325_/a_27_47# _222_/a_113_297# 1.15e-19
C1881 _078_ _313_/a_1283_21# 3.27e-20
C1882 _232_/a_32_297# _098_ 6.57e-21
C1883 net14 _310_/a_651_413# 0.00145f
C1884 _300_/a_377_297# cal_count\[3\] 3.69e-19
C1885 _090_ _228_/a_79_21# 1.96e-20
C1886 _229_/a_27_297# _088_ 1.01e-19
C1887 _337_/a_448_47# clknet_2_0__leaf_clk 0.00471f
C1888 VPWR _335_/a_543_47# 0.0157f
C1889 net28 _314_/a_805_47# 7.38e-19
C1890 ctlp[1] mask\[7\] 5.33e-20
C1891 _239_/a_694_21# _003_ 3.62e-21
C1892 _263_/a_79_21# _062_ 3.44e-19
C1893 _237_/a_218_374# _093_ 1.07e-19
C1894 trim_mask\[3\] _330_/a_1283_21# 0.00306f
C1895 _323_/a_543_47# _042_ 0.0296f
C1896 _309_/a_193_47# _074_ 0.0142f
C1897 _107_ _278_/a_27_47# 9.64e-19
C1898 _015_ _185_/a_150_297# 5.02e-19
C1899 _058_ _092_ 9.34e-19
C1900 _232_/a_32_297# clknet_0_clk 2.86e-21
C1901 VPWR _187_/a_297_47# -6.75e-19
C1902 net9 _038_ 1.21e-20
C1903 cal_itt\[0\] net4 0.122f
C1904 net13 _093_ 5.91e-20
C1905 VPWR _314_/a_1217_47# 1.22e-19
C1906 ctln[4] _275_/a_81_21# 8.88e-19
C1907 _253_/a_81_21# _086_ 3.17e-21
C1908 VPWR _332_/a_761_289# 0.0162f
C1909 _051_ cal_itt\[3\] 3.84e-20
C1910 clk _318_/a_1270_413# 3.55e-19
C1911 _020_ _152_/a_68_297# 0.00129f
C1912 _337_/a_1283_21# _065_ 5.5e-21
C1913 cal_itt\[2\] net44 4.51e-19
C1914 _048_ _226_/a_303_47# 0.00242f
C1915 _110_ _329_/a_761_289# 7.05e-19
C1916 _110_ clkbuf_2_3__f_clk/a_110_47# 1.11e-20
C1917 _195_/a_505_21# _063_ 1.54e-19
C1918 trim_mask\[0\] _262_/a_193_297# 3.38e-19
C1919 net9 _338_/a_476_47# 7.29e-20
C1920 _326_/a_1108_47# net52 9.47e-19
C1921 _227_/a_209_311# _098_ 7.16e-19
C1922 _336_/a_27_47# _264_/a_27_297# 1.96e-20
C1923 result[1] _308_/a_543_47# 2.56e-19
C1924 _281_/a_253_297# _095_ 0.00135f
C1925 _281_/a_103_199# _099_ 7.1e-21
C1926 _304_/a_27_47# _304_/a_448_47# -0.0105f
C1927 _325_/a_1108_47# mask\[2\] 4.31e-20
C1928 mask\[5\] _045_ 3.91e-21
C1929 _339_/a_27_47# _123_ 0.522f
C1930 _060_ _092_ 0.0391f
C1931 _289_/a_68_297# _299_/a_215_297# 6.49e-20
C1932 result[4] net25 1.25e-20
C1933 _249_/a_109_297# mask\[5\] 0.00411f
C1934 _267_/a_59_75# _265_/a_81_21# 0.00147f
C1935 output33/a_27_47# net34 0.0216f
C1936 VPWR _310_/a_651_413# -0.0083f
C1937 _116_ net18 0.0016f
C1938 _073_ _203_/a_59_75# 0.0023f
C1939 _340_/a_1602_47# cal_count\[2\] 0.0603f
C1940 _275_/a_81_21# _335_/a_27_47# 3.69e-19
C1941 _337_/a_27_47# _319_/a_1283_21# 1.4e-19
C1942 cal_itt\[0\] _122_ 6.25e-20
C1943 _234_/a_109_297# _282_/a_68_297# 6.46e-21
C1944 _100_ _096_ 0.017f
C1945 _235_/a_79_21# _048_ 0.0273f
C1946 _048_ net15 0.0177f
C1947 _322_/a_543_47# _074_ 0.00617f
C1948 _071_ _041_ 1.8e-20
C1949 clk clknet_2_0__leaf_clk 0.0705f
C1950 _121_ net30 0.0346f
C1951 _169_/a_109_53# _060_ 0.00124f
C1952 cal_itt\[0\] _338_/a_381_47# 4.41e-19
C1953 net27 _152_/a_150_297# 3.75e-19
C1954 rstn output6/a_27_47# 4.51e-19
C1955 input4/a_27_47# net6 0.00163f
C1956 _048_ _228_/a_79_21# 0.0501f
C1957 _167_/a_161_47# _243_/a_27_297# 0.0011f
C1958 VPWR _030_ 0.0841f
C1959 _101_ _311_/a_27_47# 6.71e-21
C1960 _033_ _105_ 1.58e-21
C1961 _081_ _078_ 0.0702f
C1962 _006_ net22 7.26e-21
C1963 _327_/a_639_47# _058_ 9.54e-19
C1964 _104_ _327_/a_27_47# 7.3e-20
C1965 mask\[1\] _208_/a_505_21# 5.76e-20
C1966 net16 _298_/a_78_199# 1.26e-20
C1967 mask\[5\] mask\[4\] 0.071f
C1968 _091_ _194_/a_113_297# 3.02e-20
C1969 _230_/a_59_75# _067_ 8.66e-19
C1970 _334_/a_1283_21# clknet_2_2__leaf_clk 1.24e-20
C1971 trim_mask\[2\] net9 0.0102f
C1972 _052_ _260_/a_250_297# 0.00202f
C1973 _146_/a_68_297# _040_ 1.18e-21
C1974 _306_/a_27_47# _050_ 3.23e-20
C1975 mask\[1\] mask\[2\] 0.014f
C1976 net43 _310_/a_805_47# 5.25e-19
C1977 _311_/a_651_413# net53 0.00167f
C1978 net4 clknet_2_0__leaf_clk 0.0188f
C1979 VPWR _247_/a_109_297# -0.0189f
C1980 net22 _121_ 7.52e-21
C1981 _324_/a_27_47# _250_/a_27_297# 1.46e-20
C1982 _259_/a_109_47# _064_ 8.36e-20
C1983 _259_/a_27_297# _104_ 0.0401f
C1984 mask\[5\] _220_/a_199_47# 0.00114f
C1985 clknet_2_1__leaf_clk rebuffer6/a_27_47# 0.0024f
C1986 _307_/a_193_47# _210_/a_113_297# 1.15e-19
C1987 VPWR _305_/a_1108_47# -0.00694f
C1988 _328_/a_193_47# _329_/a_27_47# 9.64e-20
C1989 VPWR _311_/a_639_47# 2.33e-19
C1990 state\[2\] _060_ 1.84e-19
C1991 VPWR _146_/a_68_297# 0.00871f
C1992 _324_/a_193_47# clknet_2_1__leaf_clk 0.00561f
C1993 _329_/a_27_47# net9 0.0128f
C1994 _335_/a_761_289# clknet_2_2__leaf_clk 2.9e-19
C1995 _024_ _065_ 3.21e-19
C1996 VPWR _189_/a_408_47# 4.54e-19
C1997 trim_mask\[2\] trim[2] 1.25e-19
C1998 _023_ _011_ 0.00513f
C1999 _066_ _067_ 0.0427f
C2000 _328_/a_27_47# net18 2.45e-21
C2001 _110_ cal_count\[3\] 4.11e-20
C2002 _333_/a_761_289# net46 4.86e-19
C2003 output8/a_27_47# _179_/a_27_47# 1.48e-19
C2004 _322_/a_27_47# clknet_2_1__leaf_clk 0.00946f
C2005 _104_ net54 0.00148f
C2006 _323_/a_193_47# _150_/a_27_47# 1.52e-19
C2007 _127_ trimb[1] 6.52e-19
C2008 _336_/a_1283_21# _033_ 2.48e-20
C2009 _332_/a_193_47# clknet_2_2__leaf_clk 0.00223f
C2010 _265_/a_299_297# net46 3.28e-19
C2011 _018_ net14 9.06e-21
C2012 en_co_clk _092_ 0.274f
C2013 net9 _115_ 2.05e-20
C2014 _107_ _088_ 0.0421f
C2015 mask\[5\] _020_ 0.00722f
C2016 net43 _305_/a_1270_413# 4.73e-20
C2017 _271_/a_75_212# _333_/a_27_47# 1.15e-19
C2018 _308_/a_27_47# mask\[0\] 6.38e-21
C2019 _308_/a_193_47# net22 8.85e-20
C2020 _324_/a_27_47# _009_ 5.42e-21
C2021 _321_/a_27_47# _321_/a_448_47# -0.00719f
C2022 net24 _214_/a_113_297# 0.00348f
C2023 _340_/a_27_47# _340_/a_193_47# -0.0176f
C2024 net50 _335_/a_543_47# 0.00214f
C2025 trim_val\[3\] _335_/a_1108_47# 6.12e-19
C2026 _170_/a_81_21# net41 1.75e-22
C2027 _168_/a_207_413# clknet_0_clk 2.23e-19
C2028 trim_mask\[3\] _335_/a_1283_21# 0.0277f
C2029 _308_/a_27_47# output24/a_27_47# 3.92e-20
C2030 net28 net29 0.0207f
C2031 _247_/a_109_297# net52 0.00428f
C2032 _293_/a_299_297# _144_/a_27_47# 3.09e-19
C2033 _247_/a_373_47# _101_ 0.00199f
C2034 VPWR _232_/a_114_297# -0.00259f
C2035 _008_ _311_/a_651_413# 2.01e-20
C2036 _108_ net19 8.39e-19
C2037 _292_/a_292_297# _123_ 0.00332f
C2038 _005_ clknet_2_1__leaf_clk 1.3e-21
C2039 _317_/a_543_47# net14 1.93e-19
C2040 _286_/a_439_47# _001_ 4.44e-20
C2041 _014_ _316_/a_639_47# 8.45e-19
C2042 net45 _316_/a_1270_413# 1.6e-19
C2043 _026_ trim_mask\[1\] 1.47e-19
C2044 calibrate _260_/a_250_297# 0.0028f
C2045 mask\[0\] clknet_0_clk 0.00866f
C2046 _337_/a_651_413# net55 4.2e-19
C2047 VPWR trim_mask\[1\] 1.67f
C2048 _118_ _278_/a_27_47# 0.0163f
C2049 net15 _283_/a_75_212# 5.67e-19
C2050 _231_/a_161_47# _108_ 2.1e-19
C2051 clkbuf_0_clk/a_110_47# _304_/a_1283_21# 1.75e-20
C2052 _320_/a_1283_21# _078_ 4.8e-19
C2053 trimb[1] _126_ 4.36e-19
C2054 _305_/a_1108_47# _063_ 2.71e-19
C2055 _337_/a_27_47# _337_/a_448_47# -0.00346f
C2056 _337_/a_193_47# _337_/a_1108_47# -0.00207f
C2057 VPWR _290_/a_27_413# 0.0276f
C2058 net13 mask\[6\] 0.015f
C2059 net24 _320_/a_193_47# 9.63e-20
C2060 _146_/a_68_297# net52 0.00178f
C2061 _320_/a_27_47# net45 1.04e-20
C2062 _320_/a_761_289# clknet_2_0__leaf_clk 4.81e-19
C2063 VPWR _170_/a_81_21# -3.11e-19
C2064 trim[1] _265_/a_81_21# 4.51e-20
C2065 output32/a_27_47# trim_val\[0\] 0.00905f
C2066 _330_/a_1283_21# _118_ 3.87e-22
C2067 clknet_2_3__leaf_clk net30 3.13e-21
C2068 _113_ clknet_2_2__leaf_clk 0.174f
C2069 clkbuf_2_1__f_clk/a_110_47# _016_ 0.0198f
C2070 trimb[2] net16 3.94e-19
C2071 _306_/a_1217_47# _050_ 3.14e-20
C2072 _291_/a_285_297# cal_count\[0\] 1.19e-20
C2073 _327_/a_27_47# _267_/a_59_75# 5.67e-21
C2074 VPWR _018_ 0.155f
C2075 _107_ _108_ 0.0581f
C2076 _331_/a_193_47# _171_/a_27_47# 1.18e-21
C2077 _097_ _237_/a_76_199# 0.00292f
C2078 net4 _336_/a_761_289# 0.0085f
C2079 mask\[3\] net15 0.00596f
C2080 _304_/a_27_47# net4 1.42e-21
C2081 _324_/a_1283_21# net26 1.34e-21
C2082 VPWR _227_/a_296_53# -6.7e-20
C2083 _326_/a_27_47# net25 2.09e-19
C2084 output8/a_27_47# trim_mask\[2\] 3e-19
C2085 _333_/a_1108_47# _108_ 0.0171f
C2086 _187_/a_212_413# trim_val\[0\] 1.02e-19
C2087 _320_/a_27_47# _065_ 1.76e-20
C2088 _307_/a_1108_47# _078_ 0.0138f
C2089 _307_/a_651_413# net22 0.00352f
C2090 _064_ _330_/a_27_47# 5.22e-21
C2091 trim_val\[0\] _332_/a_193_47# 1.25e-20
C2092 _265_/a_81_21# _332_/a_651_413# 2.18e-21
C2093 result[0] _078_ 4.11e-20
C2094 _126_ trimb[4] 0.00797f
C2095 _307_/a_193_47# net45 -5.4e-19
C2096 _307_/a_543_47# clknet_2_0__leaf_clk 6.3e-19
C2097 _239_/a_694_21# _229_/a_27_297# 8.56e-21
C2098 trim[3] _334_/a_761_289# 9.11e-20
C2099 _329_/a_1217_47# net9 4.37e-19
C2100 net34 _056_ 0.0887f
C2101 net33 _055_ 0.0246f
C2102 net31 trim_val\[0\] 1.55e-19
C2103 VPWR _317_/a_543_47# 0.009f
C2104 output40/a_27_47# _131_ 3.38e-21
C2105 _322_/a_193_47# mask\[6\] 5.57e-22
C2106 _060_ _226_/a_197_47# 1.78e-19
C2107 net43 output29/a_27_47# 4.29e-20
C2108 _322_/a_651_413# _042_ 2.18e-20
C2109 _122_ net33 9.06e-21
C2110 _298_/a_493_297# cal_count\[2\] 8.07e-20
C2111 _235_/a_297_47# _092_ 0.00256f
C2112 _304_/a_1270_413# _136_ 1.97e-21
C2113 _294_/a_68_297# comp 1.28e-19
C2114 net12 net55 0.00863f
C2115 net47 _067_ 0.0716f
C2116 _041_ _202_/a_79_21# 4.47e-20
C2117 net47 _070_ 0.00159f
C2118 _304_/a_27_47# _122_ 0.0101f
C2119 _053_ _330_/a_27_47# 9.79e-21
C2120 _083_ _311_/a_639_47# 2.45e-20
C2121 clknet_2_1__leaf_clk net21 0.00953f
C2122 fanout46/a_27_47# trim_mask\[4\] 0.00133f
C2123 net33 _299_/a_27_413# 1.21e-19
C2124 VPWR output33/a_27_47# 0.026f
C2125 net34 clkc 0.00407f
C2126 _030_ _333_/a_448_47# 0.00211f
C2127 net43 mask\[6\] 0.413f
C2128 _340_/a_652_21# net47 0.00132f
C2129 _037_ _304_/a_27_47# 0.00269f
C2130 net54 _235_/a_79_21# 0.0668f
C2131 ctln[7] _318_/a_651_413# 3.69e-20
C2132 net13 _318_/a_639_47# 0.00132f
C2133 cal_itt\[1\] _198_/a_27_47# 0.0581f
C2134 _093_ net3 0.0565f
C2135 _108_ _279_/a_27_47# 0.0267f
C2136 ctlp[1] net28 3.32e-19
C2137 _319_/a_1108_47# _121_ 1.8e-19
C2138 clknet_2_1__leaf_clk _312_/a_1283_21# 3.11e-20
C2139 net44 _319_/a_1270_413# 1.27e-20
C2140 _078_ net14 0.304f
C2141 _301_/a_377_297# clkc 7.52e-20
C2142 _105_ clkbuf_2_3__f_clk/a_110_47# 0.00233f
C2143 _018_ net52 0.189f
C2144 _129_ cal_count\[2\] 0.127f
C2145 _007_ _310_/a_193_47# 0.0339f
C2146 net2 _209_/a_27_47# 9.21e-20
C2147 net44 net55 0.00485f
C2148 _309_/a_761_289# _078_ 0.0257f
C2149 net4 _069_ 0.0991f
C2150 _323_/a_1283_21# _149_/a_68_297# 0.00781f
C2151 _074_ _155_/a_68_297# 0.0534f
C2152 _237_/a_218_374# _014_ 1.21e-19
C2153 _313_/a_27_47# _313_/a_639_47# -0.0015f
C2154 _336_/a_543_47# clkbuf_2_2__f_clk/a_110_47# 0.00882f
C2155 mask\[0\] _245_/a_27_297# 0.0172f
C2156 _181_/a_68_297# _108_ 0.0216f
C2157 net15 _246_/a_373_47# 4.75e-19
C2158 _038_ _091_ 1.84e-20
C2159 net25 _310_/a_761_289# 0.00128f
C2160 mask\[3\] _310_/a_193_47# 1.41e-20
C2161 VPWR _318_/a_448_47# 5.97e-19
C2162 trim_val\[1\] clknet_2_2__leaf_clk 2.5e-20
C2163 _325_/a_1108_47# _074_ 7.48e-19
C2164 _327_/a_193_47# net46 0.00521f
C2165 net24 net13 2.64e-19
C2166 _041_ _035_ 0.126f
C2167 cal_itt\[1\] net43 6.61e-21
C2168 _035_ _338_/a_1182_261# 1.83e-21
C2169 _078_ _040_ 0.00184f
C2170 _339_/a_1032_413# cal_count\[2\] 3.38e-21
C2171 _331_/a_448_47# net30 5.29e-20
C2172 _324_/a_805_47# _021_ 7.78e-20
C2173 _312_/a_543_47# _009_ 1.98e-19
C2174 cal_count\[1\] _289_/a_68_297# 0.0465f
C2175 net34 _173_/a_27_47# 0.0121f
C2176 VPWR _168_/a_297_47# -4.65e-19
C2177 net44 _070_ 0.00138f
C2178 state\[2\] _228_/a_297_47# 3.69e-19
C2179 _089_ _049_ 0.00246f
C2180 _259_/a_109_297# net46 0.00236f
C2181 _058_ net46 0.0779f
C2182 _328_/a_448_47# _026_ 2.79e-19
C2183 _328_/a_448_47# VPWR -0.00275f
C2184 _050_ net51 4.53e-21
C2185 _208_/a_218_374# _077_ 1.1e-19
C2186 _330_/a_27_47# _330_/a_448_47# -0.00642f
C2187 _208_/a_535_374# _076_ 2.47e-19
C2188 trim_val\[0\] _332_/a_1462_47# 1.25e-19
C2189 VPWR _078_ 3.79f
C2190 _307_/a_1462_47# net45 5.4e-19
C2191 _168_/a_27_413# _331_/a_448_47# 2.27e-21
C2192 _308_/a_1108_47# _319_/a_193_47# 9.39e-20
C2193 _308_/a_27_47# _319_/a_448_47# 6.41e-22
C2194 _194_/a_113_297# clkbuf_2_3__f_clk/a_110_47# 5.57e-19
C2195 _110_ _265_/a_299_297# 0.00182f
C2196 _307_/a_1108_47# _004_ 5.47e-21
C2197 _307_/a_651_413# _079_ 4.5e-20
C2198 cal_count\[3\] rebuffer3/a_75_212# 0.012f
C2199 _100_ _098_ 0.048f
C2200 net50 trim_mask\[1\] 0.191f
C2201 _315_/a_639_47# net14 7.18e-19
C2202 output39/a_27_47# net39 0.00827f
C2203 _322_/a_1283_21# _078_ 0.0128f
C2204 result[0] _004_ 0.00119f
C2205 _065_ rebuffer6/a_27_47# 3.73e-19
C2206 clk input4/a_27_47# 0.00296f
C2207 net27 net15 0.008f
C2208 _074_ mask\[1\] 0.0263f
C2209 _266_/a_68_297# net30 0.0328f
C2210 net45 _331_/a_27_47# 0.00209f
C2211 net15 _222_/a_113_297# 2.39e-19
C2212 _257_/a_27_297# rebuffer3/a_75_212# 9.43e-22
C2213 _254_/a_109_297# _048_ 0.0011f
C2214 net31 net36 0.0626f
C2215 _341_/a_27_47# _067_ 1.77e-19
C2216 VPWR _255_/a_27_47# -5.75e-19
C2217 _325_/a_193_47# _250_/a_27_297# 5.85e-20
C2218 _336_/a_1108_47# net18 1.3e-20
C2219 _051_ clk 0.357f
C2220 _065_ cal_count\[3\] 0.0151f
C2221 _002_ net19 1.69e-20
C2222 trim_mask\[1\] _333_/a_448_47# 4.06e-19
C2223 net49 _333_/a_1108_47# 0.00521f
C2224 trim_val\[1\] _333_/a_651_413# 4.79e-19
C2225 _340_/a_476_47# _122_ 0.00178f
C2226 net47 _338_/a_27_47# 0.0602f
C2227 _304_/a_543_47# net18 0.00332f
C2228 net26 net19 0.0105f
C2229 output24/a_27_47# result[3] 0.00182f
C2230 _051_ clone7/a_27_47# 1.21e-20
C2231 _107_ _170_/a_299_297# 0.00161f
C2232 _258_/a_109_297# trim_mask\[0\] 3.49e-20
C2233 _016_ net30 1.45e-19
C2234 _340_/a_1056_47# net47 6.27e-19
C2235 _315_/a_651_413# valid 7.82e-19
C2236 net13 _243_/a_27_297# 0.00819f
C2237 _325_/a_761_289# clknet_2_1__leaf_clk 6.93e-20
C2238 net23 _078_ 0.0113f
C2239 _108_ _118_ 0.351f
C2240 input4/a_27_47# net4 0.00198f
C2241 _064_ _335_/a_27_47# 4.61e-20
C2242 _327_/a_1283_21# _108_ 1.58e-19
C2243 _340_/a_476_47# _037_ 0.00251f
C2244 _239_/a_694_21# _107_ 0.00576f
C2245 net43 net24 0.069f
C2246 VPWR _270_/a_59_75# 0.0433f
C2247 _105_ cal_count\[3\] 0.0103f
C2248 _005_ net45 8.46e-20
C2249 _327_/a_543_47# _111_ 2.05e-19
C2250 result[4] _310_/a_193_47# 9.51e-19
C2251 _097_ _090_ 7.45e-19
C2252 _305_/a_193_47# _092_ 1.07e-20
C2253 mask\[4\] _311_/a_761_289# 0.0219f
C2254 _107_ _227_/a_368_53# 2.25e-19
C2255 _090_ _192_/a_548_47# 6.74e-20
C2256 _004_ net14 0.00343f
C2257 _051_ net4 0.324f
C2258 VPWR _315_/a_639_47# 8.62e-19
C2259 _230_/a_59_75# clknet_2_3__leaf_clk 0.00118f
C2260 _337_/a_805_47# net44 -0.00125f
C2261 result[6] _011_ 0.0016f
C2262 _313_/a_543_47# _010_ 0.00132f
C2263 _062_ _278_/a_27_47# 0.0153f
C2264 _291_/a_35_297# _127_ 0.167f
C2265 _078_ net52 0.0217f
C2266 net35 _332_/a_1283_21# 0.019f
C2267 _058_ _332_/a_448_47# 0.00217f
C2268 clkbuf_2_2__f_clk/a_110_47# _106_ 5.96e-21
C2269 _293_/a_81_21# _339_/a_27_47# 5.65e-20
C2270 ctln[4] _057_ 1.27e-19
C2271 _233_/a_109_47# net1 0.00476f
C2272 _002_ _001_ 2.75e-20
C2273 trimb[0] trimb[2] 0.0503f
C2274 _024_ _038_ 0.00259f
C2275 output35/a_27_47# net37 0.0127f
C2276 cal_itt\[2\] net19 9.46e-19
C2277 clknet_2_0__leaf_clk _101_ 0.137f
C2278 _328_/a_27_47# _333_/a_193_47# 2.74e-21
C2279 _327_/a_1462_47# net46 0.00119f
C2280 _291_/a_285_297# net16 0.00445f
C2281 _035_ net18 0.0212f
C2282 net9 _333_/a_27_47# 2.54e-21
C2283 clkbuf_2_0__f_clk/a_110_47# _099_ 0.00122f
C2284 trim_mask\[2\] _033_ 0.00893f
C2285 _340_/a_27_47# _339_/a_27_47# 3.88e-20
C2286 VPWR fanout47/a_27_47# 0.103f
C2287 _028_ net30 6.27e-21
C2288 net47 net17 1.8e-20
C2289 _256_/a_27_297# net18 0.0106f
C2290 clk _316_/a_1283_21# 5.68e-19
C2291 _316_/a_27_47# _316_/a_543_47# -0.00482f
C2292 _267_/a_59_75# net40 2.5e-20
C2293 _149_/a_68_297# _303_/a_543_47# 0.00374f
C2294 _297_/a_47_47# cal_count\[2\] 8.68e-19
C2295 _330_/a_27_47# _027_ 0.484f
C2296 output14/a_27_47# _314_/a_193_47# 0.00632f
C2297 _136_ net34 2.33e-20
C2298 VPWR _056_ 0.293f
C2299 _194_/a_113_297# cal_count\[3\] 1.5e-19
C2300 _125_ net37 0.00738f
C2301 _168_/a_27_413# _028_ 4.62e-19
C2302 _168_/a_207_413# clknet_2_2__leaf_clk 4.38e-20
C2303 _291_/a_35_297# _126_ 0.00393f
C2304 _144_/a_27_47# _339_/a_27_47# 1.08e-19
C2305 _066_ clknet_2_3__leaf_clk 0.29f
C2306 cal_itt\[2\] _107_ 5.64e-19
C2307 _059_ _075_ 2.71e-19
C2308 _323_/a_761_289# net47 1.56e-20
C2309 _058_ _269_/a_81_21# 3.09e-19
C2310 cal_itt\[2\] _001_ 2.07e-20
C2311 _304_/a_761_289# cal_count\[3\] 9.6e-21
C2312 VPWR _336_/a_27_47# 0.0988f
C2313 _328_/a_639_47# _025_ 2.82e-19
C2314 _328_/a_27_47# trim_mask\[4\] 9.71e-19
C2315 _328_/a_1108_47# clknet_2_2__leaf_clk 0.0568f
C2316 _304_/a_651_413# clknet_2_3__leaf_clk 6.03e-20
C2317 VPWR _004_ 0.0206f
C2318 _340_/a_1032_413# _298_/a_215_47# 1.11e-19
C2319 net4 _316_/a_1283_21# 0.00105f
C2320 _250_/a_27_297# _249_/a_27_297# 8.82e-20
C2321 _341_/a_193_47# _136_ 0.0113f
C2322 trim_mask\[0\] clkbuf_2_2__f_clk/a_110_47# 4.42e-20
C2323 _235_/a_79_21# _235_/a_382_297# 2.22e-34
C2324 _257_/a_27_297# _336_/a_1283_21# 1.8e-20
C2325 _097_ _048_ 0.0686f
C2326 _326_/a_27_47# net15 6.55e-22
C2327 _325_/a_543_47# mask\[6\] 0.0357f
C2328 _341_/a_193_47# _284_/a_68_297# 2.51e-20
C2329 _048_ _192_/a_548_47# 0.0016f
C2330 _325_/a_1108_47# net26 7.08e-20
C2331 _083_ _078_ 0.146f
C2332 _076_ rebuffer4/a_27_47# 0.0648f
C2333 state\[1\] _089_ 3.47e-20
C2334 _325_/a_639_47# _042_ 1.01e-19
C2335 clknet_2_1__leaf_clk _045_ 0.0454f
C2336 _041_ _338_/a_1182_261# 8.03e-20
C2337 _340_/a_1224_47# _122_ 7.52e-20
C2338 _338_/a_193_47# _338_/a_381_47# -0.00594f
C2339 net47 _338_/a_586_47# 0.00227f
C2340 VPWR clkc 0.265f
C2341 net3 _192_/a_505_280# 0.0117f
C2342 clknet_2_1__leaf_clk _249_/a_109_297# 0.00341f
C2343 _277_/a_75_212# net19 2.95e-21
C2344 _258_/a_27_297# trim_mask\[2\] 0.0884f
C2345 _306_/a_761_289# rebuffer4/a_27_47# 2.69e-21
C2346 trim_mask\[2\] _024_ 3e-21
C2347 net13 _321_/a_193_47# 1.73e-20
C2348 _053_ _068_ 0.00191f
C2349 _228_/a_79_21# _228_/a_382_297# 2.22e-34
C2350 clkbuf_0_clk/a_110_47# clkbuf_2_3__f_clk/a_110_47# 0.00246f
C2351 _048_ _262_/a_27_47# 0.101f
C2352 trim[1] output35/a_27_47# 9.24e-19
C2353 output32/a_27_47# trim[4] 0.00125f
C2354 _064_ _335_/a_1217_47# 3.56e-20
C2355 _104_ _335_/a_639_47# 7.42e-20
C2356 net13 _337_/a_193_47# 0.0177f
C2357 _335_/a_193_47# _330_/a_1108_47# 1.74e-20
C2358 _096_ net41 1.83e-20
C2359 _110_ _327_/a_193_47# 6.59e-21
C2360 net16 _333_/a_805_47# 0.00127f
C2361 _340_/a_1602_47# _129_ 4.04e-19
C2362 _277_/a_75_212# trim_mask\[3\] 3.63e-19
C2363 net37 net40 0.016f
C2364 result[4] _310_/a_1462_47# 2.78e-20
C2365 VPWR _287_/a_75_212# 0.0176f
C2366 net16 _109_ 0.0017f
C2367 net44 _121_ 2.33e-20
C2368 VPWR _319_/a_651_413# 0.00135f
C2369 _329_/a_27_47# _258_/a_27_297# 0.0111f
C2370 _000_ _065_ 6.57e-20
C2371 _329_/a_27_47# _024_ 1.74e-20
C2372 _237_/a_76_199# fanout45/a_27_47# 2.12e-21
C2373 _300_/a_377_297# en_co_clk 3.47e-21
C2374 VPWR _096_ 0.218f
C2375 _323_/a_761_289# net44 0.00124f
C2376 clknet_2_1__leaf_clk mask\[4\] 0.0601f
C2377 _110_ _058_ 0.0486f
C2378 trim[4] _332_/a_193_47# 1.01e-20
C2379 _249_/a_27_297# _009_ 4.03e-20
C2380 net47 _339_/a_193_47# 0.00452f
C2381 _336_/a_27_47# _063_ 9.79e-21
C2382 net31 trim[4] 0.109f
C2383 _323_/a_27_47# _323_/a_193_47# -0.00606f
C2384 _326_/a_761_289# _314_/a_543_47# 3.66e-20
C2385 _326_/a_543_47# _314_/a_761_289# 3.17e-20
C2386 _326_/a_1108_47# _314_/a_27_47# 2.25e-20
C2387 _326_/a_27_47# _314_/a_1108_47# 6.19e-20
C2388 _340_/a_1602_47# _339_/a_1032_413# 1.29e-19
C2389 _303_/a_1108_47# _035_ 7.31e-20
C2390 VPWR _173_/a_27_47# 0.0272f
C2391 _198_/a_109_47# _069_ 6.92e-19
C2392 clknet_2_1__leaf_clk _220_/a_199_47# 2.53e-20
C2393 _195_/a_218_374# _062_ 2.49e-20
C2394 net2 _208_/a_505_21# 0.0475f
C2395 _049_ _279_/a_490_47# 5.81e-20
C2396 _136_ _133_ 7.12e-19
C2397 _200_/a_209_47# _092_ 0.00314f
C2398 _302_/a_109_297# cal_count\[3\] 0.00669f
C2399 _229_/a_27_297# net55 6.38e-20
C2400 _247_/a_27_297# mask\[2\] 6.85e-19
C2401 _038_ clkbuf_2_3__f_clk/a_110_47# 7.24e-21
C2402 net30 _279_/a_314_297# 2.29e-19
C2403 _330_/a_805_47# net46 -0.00125f
C2404 ctlp[0] _314_/a_448_47# 5.04e-19
C2405 _088_ _062_ 1.38e-19
C2406 _293_/a_299_297# VPWR 0.0692f
C2407 net43 _319_/a_805_47# -0.0011f
C2408 net3 _014_ 0.0126f
C2409 _048_ wire42/a_75_212# 0.0537f
C2410 _326_/a_193_47# _310_/a_27_47# 1.33e-20
C2411 _326_/a_27_47# _310_/a_193_47# 2.81e-21
C2412 net24 _080_ 0.0117f
C2413 output7/a_27_47# net15 0.00137f
C2414 net43 _321_/a_193_47# 0.0192f
C2415 _198_/a_181_47# _067_ 0.00107f
C2416 VPWR _336_/a_1217_47# 5.34e-19
C2417 net47 clknet_2_3__leaf_clk 0.481f
C2418 VPWR _304_/a_639_47# 3.32e-19
C2419 _198_/a_181_47# _070_ 2.89e-20
C2420 _334_/a_193_47# net46 0.0151f
C2421 VPWR _340_/a_193_47# 0.0306f
C2422 net43 _337_/a_193_47# 3.14e-20
C2423 _250_/a_109_47# mask\[5\] 0.00168f
C2424 _341_/a_1462_47# _136_ 1.99e-19
C2425 ctlp[7] net20 4.56e-19
C2426 _315_/a_27_47# _241_/a_297_47# 1.52e-21
C2427 _110_ _178_/a_150_297# 0.00108f
C2428 _116_ _178_/a_68_297# 3.67e-20
C2429 net51 _208_/a_439_47# 4.69e-19
C2430 _319_/a_651_413# net52 3.39e-19
C2431 _319_/a_1108_47# _016_ 1.93e-19
C2432 output14/a_27_47# _074_ 1.54e-19
C2433 net27 _224_/a_113_297# 0.0472f
C2434 _092_ _049_ 0.291f
C2435 _216_/a_113_297# _078_ 0.0308f
C2436 _095_ net30 1.44e-19
C2437 net8 clknet_2_2__leaf_clk 0.0058f
C2438 _041_ net18 0.00946f
C2439 _321_/a_27_47# _101_ 0.457f
C2440 clknet_2_1__leaf_clk _020_ 0.349f
C2441 _338_/a_1182_261# net18 0.00254f
C2442 _341_/a_27_47# _341_/a_543_47# -0.00469f
C2443 _341_/a_193_47# _341_/a_761_289# -0.0177f
C2444 _320_/a_543_47# _121_ 5.22e-20
C2445 clone1/a_27_47# _260_/a_250_297# 7.24e-21
C2446 net13 _321_/a_1462_47# 2.3e-19
C2447 _320_/a_448_47# net44 -1.86e-19
C2448 _263_/a_79_21# _100_ 2.66e-19
C2449 _341_/a_1283_21# _037_ 9.46e-20
C2450 net47 _303_/a_193_47# 0.00512f
C2451 _071_ _190_/a_27_47# 0.00405f
C2452 cal_itt\[0\] _190_/a_655_47# 0.00446f
C2453 cal_itt\[1\] _190_/a_465_47# 0.00167f
C2454 _041_ _129_ 0.00225f
C2455 _336_/a_193_47# net19 0.014f
C2456 output31/a_27_47# net37 1.08e-19
C2457 _335_/a_27_47# _027_ 6.08e-20
C2458 _094_ _137_/a_68_297# 5.3e-20
C2459 _062_ _108_ 0.0054f
C2460 _169_/a_215_311# _318_/a_543_47# 4.71e-20
C2461 _332_/a_651_413# net40 6.24e-19
C2462 _262_/a_27_47# _190_/a_27_47# 2.9e-21
C2463 net27 _250_/a_27_297# 8.68e-19
C2464 net28 _313_/a_1283_21# 0.0902f
C2465 net50 _336_/a_27_47# 2.82e-21
C2466 _329_/a_761_289# trim_mask\[2\] 2.59e-19
C2467 _164_/a_161_47# _096_ 0.00593f
C2468 net4 _261_/a_113_47# 1.27e-19
C2469 _014_ _241_/a_388_297# 0.00143f
C2470 net45 _241_/a_105_352# 9.84e-19
C2471 VPWR _321_/a_639_47# 2.07e-19
C2472 _309_/a_1108_47# _143_/a_68_297# 1.04e-20
C2473 net3 _243_/a_27_297# 0.00209f
C2474 mask\[7\] net14 3.5e-19
C2475 _117_ _104_ 8.64e-20
C2476 _012_ sample 3.98e-19
C2477 _333_/a_1283_21# net33 0.00975f
C2478 clknet_2_1__leaf_clk _222_/a_199_47# 4.52e-19
C2479 _041_ _339_/a_1032_413# 0.044f
C2480 net47 _339_/a_796_47# -7.54e-19
C2481 net44 clknet_2_3__leaf_clk 0.00416f
C2482 VPWR _337_/a_639_47# 2.44e-19
C2483 VPWR _313_/a_1108_47# 0.0234f
C2484 _336_/a_193_47# _107_ 0.00241f
C2485 _309_/a_27_47# _023_ 1.73e-22
C2486 _042_ _084_ 6.34e-21
C2487 _340_/a_193_47# _063_ 3.52e-20
C2488 _310_/a_193_47# _310_/a_761_289# -0.00517f
C2489 output22/a_27_47# _307_/a_193_47# 2.18e-19
C2490 _334_/a_1283_21# _108_ 4.38e-19
C2491 _046_ _313_/a_27_47# 0.0294f
C2492 VPWR _172_/a_68_297# 0.00573f
C2493 _038_ cal_count\[3\] 0.0216f
C2494 state\[2\] _049_ 0.00628f
C2495 _015_ _318_/a_448_47# 0.00397f
C2496 state\[2\] _318_/a_761_289# 0.00114f
C2497 VPWR _136_ 0.481f
C2498 _308_/a_639_47# _006_ 1.56e-20
C2499 _337_/a_543_47# _090_ 8.11e-22
C2500 _128_ _340_/a_1032_413# 0.0117f
C2501 _036_ _340_/a_193_47# 1.63e-19
C2502 _134_ _298_/a_292_297# 6.3e-20
C2503 VPWR _284_/a_68_297# 0.0151f
C2504 _301_/a_47_47# clknet_2_3__leaf_clk 0.117f
C2505 _303_/a_193_47# net44 0.00334f
C2506 _306_/a_1283_21# _305_/a_448_47# 3.74e-19
C2507 net55 net19 1.79e-20
C2508 _262_/a_193_297# _092_ 9.77e-20
C2509 _326_/a_1283_21# _074_ 5.88e-20
C2510 _329_/a_193_47# net18 5.13e-20
C2511 net27 _009_ 3.17e-19
C2512 _341_/a_27_47# clknet_2_3__leaf_clk 0.567f
C2513 _281_/a_103_199# _192_/a_505_280# 0.00113f
C2514 _320_/a_27_47# _320_/a_639_47# -0.0015f
C2515 _309_/a_543_47# _081_ 6.06e-19
C2516 _309_/a_193_47# _006_ 0.0343f
C2517 _323_/a_27_47# _303_/a_27_47# 1.62e-20
C2518 _316_/a_761_289# net41 0.0219f
C2519 VPWR _340_/a_796_47# 3.86e-19
C2520 trim[1] output31/a_27_47# 0.00179f
C2521 output32/a_27_47# trim[0] 1.44e-19
C2522 result[2] _007_ 4.52e-19
C2523 net43 _313_/a_1270_413# -2.06e-19
C2524 _129_ _298_/a_493_297# 1.98e-20
C2525 _336_/a_1108_47# trim_mask\[4\] 0.0389f
C2526 VPWR mask\[7\] 0.441f
C2527 _306_/a_193_47# clknet_2_1__leaf_clk 1.45e-19
C2528 net12 net20 0.0134f
C2529 _081_ _245_/a_27_297# 1.53e-19
C2530 _264_/a_27_297# clknet_2_2__leaf_clk 7.38e-19
C2531 net12 net53 0.0178f
C2532 _308_/a_27_47# _307_/a_1108_47# 4.25e-21
C2533 _308_/a_543_47# _307_/a_761_289# 2.14e-20
C2534 _308_/a_1108_47# _307_/a_27_47# 3.02e-20
C2535 _308_/a_761_289# _307_/a_543_47# 7.82e-20
C2536 output27/a_27_47# result[7] 0.00234f
C2537 clk _119_ 2.39e-20
C2538 net16 comp 3e-20
C2539 result[0] _308_/a_27_47# 0.00211f
C2540 _187_/a_27_413# _332_/a_1283_21# 1.11e-19
C2541 _048_ _206_/a_27_93# 2.7e-20
C2542 _338_/a_1296_47# net18 2.78e-19
C2543 _336_/a_27_47# _279_/a_396_47# 0.00922f
C2544 _336_/a_193_47# _279_/a_27_47# 0.0013f
C2545 _326_/a_27_47# _224_/a_113_297# 2.65e-20
C2546 _107_ net55 0.116f
C2547 VPWR _316_/a_761_289# 0.00842f
C2548 _303_/a_1108_47# _041_ 4.03e-20
C2549 _067_ net19 0.0106f
C2550 _332_/a_193_47# _332_/a_543_47# -0.02f
C2551 _332_/a_193_47# _108_ 0.397f
C2552 _332_/a_27_47# _332_/a_1283_21# -8.77e-19
C2553 net47 _303_/a_1462_47# 0.00104f
C2554 net19 _070_ 0.0709f
C2555 _189_/a_408_47# _075_ 1.97e-19
C2556 VPWR ctln[6] 0.0347f
C2557 _111_ _332_/a_27_47# 2.22e-19
C2558 _231_/a_161_47# _067_ 0.0161f
C2559 _335_/a_805_47# net46 0.00132f
C2560 net31 _108_ 0.0162f
C2561 _328_/a_805_47# _058_ 2.61e-19
C2562 _104_ _328_/a_193_47# 2.53e-20
C2563 _268_/a_75_212# _111_ 0.0121f
C2564 clk _331_/a_651_413# 0.00269f
C2565 _104_ net9 3.84e-19
C2566 net31 trim[0] 0.00511f
C2567 net44 net20 0.0362f
C2568 ctln[6] _331_/a_1283_21# 1.83e-21
C2569 net44 net53 0.123f
C2570 _058_ rebuffer3/a_75_212# 0.0034f
C2571 net4 _119_ 0.648f
C2572 _327_/a_193_47# _065_ 1.61e-20
C2573 _333_/a_27_47# net32 7.72e-20
C2574 net42 _226_/a_27_47# 4.92e-20
C2575 _324_/a_651_413# net44 0.00317f
C2576 state\[1\] _092_ 0.00946f
C2577 _048_ _337_/a_543_47# 5.1e-21
C2578 trim_mask\[2\] _257_/a_27_297# 0.00807f
C2579 _324_/a_1108_47# _323_/a_193_47# 7.71e-20
C2580 net3 _337_/a_193_47# 6.11e-19
C2581 _256_/a_27_297# trim_mask\[4\] 0.0098f
C2582 _025_ trim_mask\[0\] 0.00129f
C2583 _001_ _067_ 9.01e-19
C2584 _001_ _070_ 0.013f
C2585 _326_/a_193_47# clknet_2_1__leaf_clk 0.0245f
C2586 _308_/a_27_47# net14 0.00787f
C2587 _189_/a_218_47# _088_ 1.17e-19
C2588 _058_ _065_ 8.88e-19
C2589 _050_ _336_/a_448_47# 8.9e-21
C2590 _113_ _108_ 9.94e-20
C2591 VPWR _323_/a_193_47# -0.293f
C2592 result[0] _307_/a_448_47# 6.73e-19
C2593 _169_/a_109_53# state\[1\] 0.0393f
C2594 _074_ _310_/a_448_47# 0.00248f
C2595 _314_/a_193_47# net29 0.00644f
C2596 mask\[7\] net52 0.121f
C2597 _339_/a_1032_413# _129_ 6.61e-20
C2598 _292_/a_215_47# _122_ 0.0632f
C2599 _322_/a_448_47# net44 5.15e-19
C2600 _060_ net45 1.14e-19
C2601 _309_/a_27_47# _308_/a_761_289# 3.48e-21
C2602 _309_/a_193_47# _308_/a_193_47# 1.43e-21
C2603 _233_/a_109_47# _012_ 3.65e-20
C2604 net4 _087_ 2.67e-20
C2605 _110_ _334_/a_193_47# 0.00154f
C2606 net21 _313_/a_639_47# 1.32e-19
C2607 _335_/a_27_47# _032_ 0.0366f
C2608 net12 _008_ 0.00728f
C2609 _051_ _260_/a_250_297# 2.34e-19
C2610 _325_/a_193_47# _321_/a_543_47# 8.89e-21
C2611 _188_/a_27_47# net35 1.73e-19
C2612 _104_ _262_/a_109_297# 4.63e-19
C2613 _282_/a_150_297# _090_ 2.4e-20
C2614 _226_/a_197_47# _049_ 7.09e-20
C2615 _078_ _208_/a_76_199# 9.44e-19
C2616 _311_/a_193_47# _311_/a_448_47# -0.00482f
C2617 VPWR _301_/a_129_47# -7.64e-19
C2618 _325_/a_27_47# _313_/a_27_47# 7.57e-19
C2619 _306_/a_1283_21# _002_ 2.36e-19
C2620 ctln[3] _057_ 0.0412f
C2621 _187_/a_27_413# _135_ 0.00107f
C2622 _103_ _060_ 8.17e-21
C2623 _341_/a_448_47# cal_count\[3\] 0.0163f
C2624 VPWR _338_/a_1140_413# 1.88e-20
C2625 _291_/a_35_297# net47 8.66e-20
C2626 mask\[0\] mask\[2\] 1.12e-19
C2627 _341_/a_1217_47# clknet_2_3__leaf_clk 0.00112f
C2628 VPWR _341_/a_761_289# 0.00858f
C2629 en_co_clk _192_/a_476_47# 1.07e-19
C2630 _120_ _192_/a_505_280# 0.183f
C2631 net2 _108_ 4.09e-20
C2632 net2 _332_/a_543_47# 1.14e-19
C2633 net4 _266_/a_150_297# 1.65e-19
C2634 _094_ _232_/a_32_297# 1.95e-21
C2635 _060_ _065_ 5.79e-21
C2636 _013_ output41/a_27_47# 2.01e-20
C2637 net13 _320_/a_1270_413# 1.5e-19
C2638 VPWR _299_/a_382_47# -4.75e-19
C2639 _040_ clknet_0_clk 0.0218f
C2640 _321_/a_27_47# _248_/a_27_297# 1.74e-20
C2641 trim_mask\[1\] _334_/a_1108_47# 9.68e-21
C2642 VPWR _098_ 0.0378f
C2643 _272_/a_299_297# _334_/a_543_47# 1.49e-19
C2644 _008_ net44 6.48e-19
C2645 _320_/a_1108_47# _040_ 0.0346f
C2646 output13/a_27_47# net13 0.0457f
C2647 _053_ _262_/a_205_47# 1.72e-19
C2648 VPWR _308_/a_27_47# 0.0953f
C2649 state\[2\] state\[1\] 0.204f
C2650 _113_ _031_ 0.00248f
C2651 output22/a_27_47# _005_ 1.31e-20
C2652 net15 _318_/a_193_47# 7.1e-21
C2653 _336_/a_193_47# _118_ 3.81e-21
C2654 mask\[1\] _319_/a_1270_413# 8.1e-21
C2655 clk input3/a_75_212# 0.00131f
C2656 trim_mask\[0\] _333_/a_543_47# 1.73e-19
C2657 net4 _199_/a_193_297# 4.24e-19
C2658 _303_/a_1108_47# net18 2.39e-19
C2659 _071_ _306_/a_27_47# 1.97e-21
C2660 _029_ _332_/a_805_47# 9.23e-20
C2661 VPWR clknet_0_clk 0.814f
C2662 trim_mask\[0\] _265_/a_384_47# 0.00132f
C2663 net35 net33 0.415f
C2664 net50 _136_ 0.00145f
C2665 _185_/a_68_297# net55 3.84e-19
C2666 net54 _243_/a_109_47# 1.14e-19
C2667 _060_ _243_/a_109_297# 0.00385f
C2668 VPWR _320_/a_1108_47# 0.00694f
C2669 _050_ _337_/a_1283_21# 0.00416f
C2670 _181_/a_68_297# _067_ 3.4e-20
C2671 VPWR _339_/a_27_47# -0.259f
C2672 net12 _028_ 0.00295f
C2673 _286_/a_439_47# _123_ 5.37e-20
C2674 clknet_2_1__leaf_clk _310_/a_543_47# 0.0364f
C2675 _022_ _085_ 0.00128f
C2676 _333_/a_1217_47# net32 7.32e-20
C2677 _088_ _227_/a_209_311# 0.00384f
C2678 _326_/a_761_289# mask\[6\] 2.18e-21
C2679 net9 _267_/a_59_75# 3.47e-19
C2680 _326_/a_1283_21# net26 2.13e-20
C2681 fanout44/a_27_47# _337_/a_193_47# 4.94e-20
C2682 cal_itt\[2\] _062_ 0.00126f
C2683 clkbuf_2_0__f_clk/a_110_47# _093_ 2.69e-21
C2684 net15 _317_/a_639_47# 0.00103f
C2685 _308_/a_543_47# net43 0.00229f
C2686 _308_/a_27_47# net23 2.61e-19
C2687 _308_/a_1283_21# _005_ 4.73e-20
C2688 ctlp[6] _312_/a_761_289# 0.00104f
C2689 _191_/a_27_297# net18 1.36e-19
C2690 net49 _332_/a_193_47# 1.04e-19
C2691 trim_val\[1\] _108_ 0.139f
C2692 _324_/a_1283_21# clknet_2_3__leaf_clk 5.51e-21
C2693 _112_ _332_/a_27_47# 6.36e-19
C2694 _050_ _033_ 9.69e-19
C2695 VPWR _323_/a_1462_47# 1.98e-19
C2696 VPWR _307_/a_448_47# 0.00114f
C2697 net45 en_co_clk 2.3e-20
C2698 trim[0] trim_val\[1\] 0.00247f
C2699 net31 net49 0.00371f
C2700 _314_/a_1462_47# net29 4.31e-19
C2701 _288_/a_59_75# net33 0.00892f
C2702 _019_ net44 8.34e-20
C2703 en_co_clk rebuffer3/a_75_212# 1.38e-21
C2704 trimb[2] net39 0.00735f
C2705 _329_/a_651_413# VPWR 0.0028f
C2706 input2/a_27_47# clkc 5.42e-19
C2707 _327_/a_27_47# _256_/a_27_297# 5.24e-19
C2708 net31 _290_/a_207_413# 7.34e-19
C2709 _309_/a_543_47# net14 0.0113f
C2710 _335_/a_1217_47# _032_ 1.04e-20
C2711 _015_ _096_ 1.64e-19
C2712 _321_/a_543_47# mask\[3\] 2.36e-20
C2713 cal_itt\[2\] _195_/a_76_199# 5.23e-21
C2714 _129_ _297_/a_47_47# 0.0425f
C2715 net42 _052_ 5.72e-21
C2716 _103_ en_co_clk 1.3e-20
C2717 _125_ cal_count\[2\] 2.52e-20
C2718 trim_val\[2\] net46 0.00456f
C2719 _324_/a_1108_47# _303_/a_27_47# 1.54e-20
C2720 clknet_2_0__leaf_clk _077_ -1.01e-24
C2721 clknet_0_clk net52 0.119f
C2722 en_co_clk _065_ 0.198f
C2723 clknet_0_clk _063_ 0.0459f
C2724 _305_/a_193_47# clknet_2_1__leaf_clk 1.36e-19
C2725 _074_ net29 3.58e-19
C2726 _320_/a_1108_47# net52 2.33e-20
C2727 _306_/a_543_47# clknet_2_0__leaf_clk 1.49e-19
C2728 _306_/a_193_47# net45 4.54e-22
C2729 clknet_2_1__leaf_clk _311_/a_1108_47# 0.00435f
C2730 _313_/a_193_47# _158_/a_150_297# 9.72e-20
C2731 net28 net14 0.398f
C2732 VPWR _303_/a_27_47# 0.0756f
C2733 _078_ _314_/a_27_47# 9.87e-19
C2734 _323_/a_761_289# net19 0.00947f
C2735 _043_ mask\[4\] 0.0669f
C2736 _305_/a_805_47# net51 1.55e-19
C2737 _030_ trim_mask\[1\] 0.104f
C2738 _113_ net49 0.0029f
C2739 _114_ _334_/a_448_47# 2.07e-19
C2740 trim_val\[2\] _334_/a_639_47# 1.48e-19
C2741 _234_/a_109_297# net15 0.00108f
C2742 net16 net46 0.0561f
C2743 VPWR _308_/a_1217_47# 5.6e-20
C2744 _140_/a_68_297# _101_ 0.00187f
C2745 _040_ _245_/a_27_297# 1.86e-19
C2746 _337_/a_1108_47# _092_ 2.64e-19
C2747 net3 _316_/a_1108_47# 9.66e-19
C2748 trim_mask\[2\] _333_/a_761_289# 4.36e-20
C2749 _128_ _339_/a_1182_261# 0.0153f
C2750 _036_ _339_/a_27_47# 0.042f
C2751 cal_count\[1\] _339_/a_193_47# -1.26e-21
C2752 calibrate _227_/a_109_93# 3.13e-20
C2753 _052_ _054_ 3.87e-19
C2754 _306_/a_193_47# _065_ 1.17e-20
C2755 _052_ net30 1.34e-20
C2756 net7 output6/a_27_47# 1.39e-19
C2757 clkbuf_0_clk/a_110_47# _190_/a_215_47# 0.00413f
C2758 _004_ output30/a_27_47# 0.0445f
C2759 _058_ _302_/a_109_297# 0.00122f
C2760 _211_/a_109_297# sample 3.96e-19
C2761 VPWR _309_/a_543_47# -0.00123f
C2762 _117_ fanout46/a_27_47# 5.57e-19
C2763 en_co_clk _243_/a_109_297# 7.06e-19
C2764 _281_/a_253_47# _096_ 2.32e-19
C2765 _328_/a_761_289# net46 0.00311f
C2766 mask\[7\] _216_/a_113_297# 1.54e-19
C2767 _325_/a_448_47# mask\[7\] 5.89e-20
C2768 _253_/a_299_297# mask\[3\] 1.23e-21
C2769 net12 _205_/a_27_47# 0.00291f
C2770 VPWR _339_/a_586_47# 5.47e-20
C2771 cal_count\[2\] net40 0.00976f
C2772 calibrate _317_/a_193_47# 4.8e-21
C2773 _093_ _317_/a_27_47# 6.21e-22
C2774 VPWR _245_/a_27_297# 0.024f
C2775 _292_/a_78_199# _292_/a_292_297# -1.09e-21
C2776 _104_ _336_/a_448_47# 2.61e-19
C2777 net54 _337_/a_543_47# 1.26e-21
C2778 ctln[1] _317_/a_761_289# 2.4e-20
C2779 _168_/a_27_413# _052_ 0.00112f
C2780 _324_/a_1283_21# net53 2.43e-21
C2781 _290_/a_207_413# net2 1.2e-19
C2782 _094_ mask\[0\] 0.0048f
C2783 _169_/a_109_53# _167_/a_161_47# 3.05e-19
C2784 _328_/a_27_47# _271_/a_75_212# 1.35e-20
C2785 _326_/a_1108_47# _078_ 0.00364f
C2786 result[3] net14 8.01e-20
C2787 ctlp[0] _086_ 1.04e-19
C2788 net7 net45 1.3e-20
C2789 VPWR net28 1.8f
C2790 _237_/a_76_199# _090_ 0.00486f
C2791 cal_count\[1\] trimb[4] 5.25e-20
C2792 VPWR _292_/a_292_297# 4.73e-19
C2793 _247_/a_109_297# _018_ 8.09e-19
C2794 net37 _132_ 0.00591f
C2795 trim_val\[0\] net34 8.77e-19
C2796 net42 calibrate 3.11e-19
C2797 VPWR _324_/a_448_47# 0.00366f
C2798 net44 _205_/a_27_47# 0.00463f
C2799 _043_ _020_ 2.16e-21
C2800 _341_/a_543_47# _001_ 2.66e-19
C2801 _303_/a_27_47# _063_ 4.53e-21
C2802 _309_/a_448_47# net43 3.46e-20
C2803 _210_/a_113_297# _039_ 6.7e-20
C2804 _327_/a_761_289# trim_mask\[0\] 7.95e-19
C2805 net4 _279_/a_206_47# 3.06e-19
C2806 _146_/a_68_297# _018_ 0.00373f
C2807 _002_ net2 0.0574f
C2808 _305_/a_1283_21# _002_ 0.00336f
C2809 net23 _245_/a_27_297# 0.0304f
C2810 cal_itt\[1\] _068_ 0.171f
C2811 net16 _332_/a_448_47# 4.27e-19
C2812 _316_/a_27_47# _095_ 1.61e-19
C2813 _277_/a_75_212# _335_/a_761_289# 7.23e-19
C2814 net2 _289_/a_68_297# 0.0256f
C2815 VPWR _322_/a_1108_47# 0.0234f
C2816 net9 _300_/a_129_47# 4.46e-19
C2817 _329_/a_448_47# clknet_2_2__leaf_clk 1.12e-19
C2818 _329_/a_193_47# trim_mask\[4\] 1.26e-19
C2819 _314_/a_543_47# _011_ 0.00283f
C2820 _099_ clone7/a_27_47# 7.04e-20
C2821 net12 _095_ 6.2e-21
C2822 VPWR _331_/a_1108_47# 0.0235f
C2823 _311_/a_1270_413# net26 4.38e-19
C2824 VPWR _159_/a_27_47# 0.0491f
C2825 state\[2\] _167_/a_161_47# 7.2e-19
C2826 ctlp[1] _074_ 5.89e-19
C2827 _309_/a_1108_47# _101_ 0.00106f
C2828 _064_ _256_/a_373_47# 2.84e-19
C2829 _104_ _256_/a_109_297# 0.00107f
C2830 _320_/a_1283_21# _209_/a_27_47# 0.0148f
C2831 _251_/a_27_297# clknet_2_1__leaf_clk 0.0348f
C2832 calibrate _054_ 6.74e-19
C2833 VPWR _303_/a_1217_47# 1.15e-19
C2834 _169_/a_215_311# clk 2.62e-20
C2835 trim_val\[1\] net49 0.115f
C2836 VPWR result[3] 0.0946f
C2837 _245_/a_27_297# net52 0.031f
C2838 calibrate net30 0.00261f
C2839 net15 _319_/a_761_289# 0.00236f
C2840 _327_/a_1108_47# _136_ 0.00119f
C2841 trim_mask\[4\] net18 0.366f
C2842 _169_/a_215_311# clone7/a_27_47# 6.11e-19
C2843 _328_/a_1283_21# _111_ 2.19e-19
C2844 clknet_2_3__leaf_clk net19 0.0276f
C2845 _114_ _031_ 0.00585f
C2846 _305_/a_543_47# _203_/a_59_75# 7.48e-19
C2847 trim[1] trim[2] 3.16e-20
C2848 _006_ mask\[1\] 3.35e-19
C2849 cal_itt\[2\] net2 0.0512f
C2850 _231_/a_161_47# clknet_2_3__leaf_clk 0.00105f
C2851 net19 _153_/a_27_47# 0.0105f
C2852 net28 net52 0.00395f
C2853 cal_itt\[2\] _305_/a_1283_21# 0.0316f
C2854 net16 _269_/a_81_21# 0.00875f
C2855 _128_ _339_/a_1296_47# 3.98e-19
C2856 _237_/a_76_199# _048_ 0.0131f
C2857 mask\[3\] _041_ 8.1e-20
C2858 _058_ _038_ 0.00111f
C2859 _059_ _096_ 0.0162f
C2860 calibrate net22 1.75e-20
C2861 _169_/a_215_311# net4 0.0528f
C2862 _303_/a_1283_21# _000_ 9.79e-21
C2863 _074_ mask\[0\] 1.13e-20
C2864 _116_ _117_ 0.221f
C2865 net24 _310_/a_1283_21# 3.61e-22
C2866 output24/a_27_47# _074_ 0.0126f
C2867 _303_/a_193_47# net19 0.0168f
C2868 net31 output5/a_27_47# 0.00676f
C2869 _337_/a_193_47# _120_ 9.35e-20
C2870 _337_/a_761_289# en_co_clk 0.00551f
C2871 _292_/a_493_297# cal_count\[1\] 0.00114f
C2872 _292_/a_292_297# _036_ 6.14e-19
C2873 _104_ _033_ 0.0252f
C2874 _107_ clknet_2_3__leaf_clk 0.00643f
C2875 VPWR _263_/a_79_21# 0.00206f
C2876 clkbuf_2_0__f_clk/a_110_47# _192_/a_505_280# 0.00268f
C2877 _001_ clknet_2_3__leaf_clk 0.381f
C2878 output15/a_27_47# _251_/a_27_297# 7.82e-21
C2879 clknet_0_clk _279_/a_396_47# 1.14e-20
C2880 net26 net29 2.24e-20
C2881 net31 _270_/a_145_75# 2.11e-20
C2882 _321_/a_1270_413# mask\[2\] 6e-20
C2883 _289_/a_68_297# _123_ 6.19e-21
C2884 _337_/a_193_47# _076_ 3.9e-20
C2885 _218_/a_113_297# _101_ 2.38e-19
C2886 _110_ trim_val\[2\] 2.39e-19
C2887 _227_/a_209_311# _227_/a_368_53# 8.88e-34
C2888 clknet_2_1__leaf_clk _049_ 5.62e-19
C2889 ctln[2] _334_/a_1283_21# 8.69e-19
C2890 net8 _334_/a_448_47# 0.00107f
C2891 _323_/a_27_47# _044_ 4.75e-20
C2892 _232_/a_32_297# _192_/a_174_21# 0.0237f
C2893 net31 output36/a_27_47# 0.00817f
C2894 net36 net34 0.206f
C2895 net10 VPWR 0.0521f
C2896 _136_ _193_/a_109_297# 4.88e-19
C2897 net45 _039_ 0.214f
C2898 _304_/a_761_289# _286_/a_76_199# 9.16e-22
C2899 _251_/a_109_297# mask\[6\] 0.00185f
C2900 mask\[6\] _250_/a_373_47# 4.1e-19
C2901 output23/a_27_47# output24/a_27_47# 0.0217f
C2902 _250_/a_27_297# _021_ 0.0107f
C2903 _026_ clknet_2_2__leaf_clk 0.0985f
C2904 _312_/a_651_413# net20 0.00219f
C2905 _096_ _075_ 5.91e-20
C2906 _110_ net16 0.0575f
C2907 VPWR clknet_2_2__leaf_clk 2.08f
C2908 net55 _062_ 0.00671f
C2909 VPWR _260_/a_584_47# -8.99e-19
C2910 mask\[6\] _042_ 1.95e-19
C2911 _308_/a_193_47# mask\[1\] 6.5e-20
C2912 calibrate _315_/a_651_413# 0.0256f
C2913 _012_ _315_/a_1283_21# 4.1e-20
C2914 _146_/a_68_297# _078_ 5.82e-19
C2915 trim_mask\[2\] _058_ 0.00127f
C2916 _259_/a_109_297# trim_mask\[2\] 8.17e-20
C2917 _104_ _258_/a_27_297# 0.0723f
C2918 _064_ _258_/a_109_47# 0.00199f
C2919 _322_/a_543_47# _019_ 2.8e-19
C2920 _104_ _024_ 0.00764f
C2921 _300_/a_285_47# cal_count\[2\] 1.85e-20
C2922 _239_/a_27_297# net42 0.00125f
C2923 _331_/a_1283_21# clknet_2_2__leaf_clk 5.33e-20
C2924 _331_/a_543_47# _028_ 0.0336f
C2925 _113_ _270_/a_145_75# 8.31e-19
C2926 _030_ _270_/a_59_75# 3.44e-19
C2927 _064_ net4 0.0666f
C2928 clkbuf_0_clk/a_110_47# en_co_clk 3.63e-19
C2929 _053_ clk 0.00574f
C2930 _317_/a_193_47# _317_/a_1108_47# -0.00677f
C2931 state\[0\] _316_/a_27_47# 2.39e-19
C2932 _272_/a_81_21# _114_ 0.00604f
C2933 _272_/a_299_297# net48 0.0443f
C2934 _237_/a_505_21# _050_ 0.00133f
C2935 net2 output5/a_27_47# 9.38e-19
C2936 _332_/a_27_47# net33 7.1e-21
C2937 net12 state\[0\] 1.7e-20
C2938 _053_ clone7/a_27_47# 8.25e-20
C2939 _046_ net21 0.0107f
C2940 clkbuf_2_1__f_clk/a_110_47# clknet_2_0__leaf_clk 0.0448f
C2941 VPWR net11 0.265f
C2942 _110_ _328_/a_761_289# 5.43e-20
C2943 _320_/a_448_47# mask\[1\] 0.0111f
C2944 _305_/a_651_413# _072_ 0.00299f
C2945 _040_ _209_/a_27_47# 3.17e-19
C2946 _322_/a_1108_47# _083_ 0.00198f
C2947 _305_/a_193_47# _065_ 7.67e-20
C2948 _067_ _062_ 0.035f
C2949 VPWR _236_/a_109_297# -0.00218f
C2950 _062_ _070_ 3.11e-20
C2951 _331_/a_448_47# net19 5.77e-19
C2952 _259_/a_27_297# _329_/a_193_47# 3.28e-19
C2953 _327_/a_27_47# net18 0.0237f
C2954 _181_/a_68_297# clknet_2_3__leaf_clk 3.62e-21
C2955 net15 _313_/a_27_47# 0.00107f
C2956 net8 _108_ 4.46e-19
C2957 _088_ _100_ 3.2e-19
C2958 _170_/a_384_47# _054_ 1.88e-20
C2959 _323_/a_1108_47# mask\[4\] 0.019f
C2960 net5 _300_/a_47_47# 7.07e-21
C2961 net12 _208_/a_218_374# 6.82e-19
C2962 _318_/a_27_47# _318_/a_193_47# -0.019f
C2963 _034_ clknet_0_clk 0.127f
C2964 net12 _207_/a_109_297# 4.37e-19
C2965 output10/a_27_47# _275_/a_299_297# 4.68e-19
C2966 _053_ net4 1.21f
C2967 _306_/a_193_47# clkbuf_0_clk/a_110_47# 2.77e-19
C2968 VPWR _209_/a_27_47# 0.0457f
C2969 _282_/a_68_297# en_co_clk 2.2e-21
C2970 _239_/a_474_297# _049_ 0.00562f
C2971 _021_ _009_ 2.08e-20
C2972 _086_ _224_/a_113_297# 0.00758f
C2973 _259_/a_27_297# net18 0.00703f
C2974 _328_/a_448_47# trim_mask\[1\] 0.0164f
C2975 _322_/a_1283_21# _209_/a_27_47# 9.72e-19
C2976 VPWR _333_/a_651_413# 0.00154f
C2977 _195_/a_76_199# _067_ 3.99e-20
C2978 _081_ mask\[2\] 3.52e-19
C2979 _015_ clknet_0_clk 2e-20
C2980 _266_/a_68_297# net19 0.00778f
C2981 VPWR trim_val\[0\] 0.146f
C2982 cal_count\[1\] _291_/a_35_297# 4.78e-21
C2983 _290_/a_297_47# _126_ 1.43e-19
C2984 _038_ en_co_clk 2.04e-19
C2985 _309_/a_543_47# _216_/a_113_297# 2.12e-19
C2986 _200_/a_209_297# _071_ 4.88e-19
C2987 net12 _226_/a_27_47# 2.37e-20
C2988 _050_ _331_/a_27_47# 7.37e-19
C2989 net44 _207_/a_109_297# 2.44e-19
C2990 _336_/a_639_47# _052_ 4.96e-21
C2991 _053_ _122_ 0.19f
C2992 net8 _031_ 0.00114f
C2993 net20 _155_/a_68_297# 2.23e-19
C2994 _325_/a_805_47# net13 1.81e-19
C2995 _326_/a_27_47# _253_/a_299_297# 9.57e-19
C2996 _326_/a_193_47# _253_/a_81_21# 2.09e-19
C2997 net28 _155_/a_150_297# 8.39e-21
C2998 _078_ _018_ 0.00646f
C2999 clk _330_/a_448_47# 7.28e-19
C3000 _041_ rebuffer5/a_161_47# 4.56e-21
C3001 _275_/a_81_21# trim_val\[3\] 0.0377f
C3002 _314_/a_1108_47# _313_/a_27_47# 1.43e-20
C3003 _041_ _125_ 0.0167f
C3004 _053_ _037_ 0.00216f
C3005 _141_/a_27_47# clknet_0_clk 0.0326f
C3006 mask\[6\] _022_ 0.0576f
C3007 _325_/a_1108_47# net53 2.71e-20
C3008 _328_/a_27_47# _328_/a_193_47# -0.328f
C3009 result[1] net45 3.22e-20
C3010 _320_/a_1108_47# _141_/a_27_47# 2e-19
C3011 net30 _203_/a_59_75# 0.0435f
C3012 _266_/a_68_297# _107_ 0.00884f
C3013 _237_/a_218_374# _092_ 5.89e-19
C3014 net43 _212_/a_113_297# 0.00838f
C3015 net37 net32 0.0391f
C3016 _328_/a_27_47# net9 0.00722f
C3017 output31/a_27_47# _162_/a_27_47# 8.1e-20
C3018 _048_ _090_ 0.282f
C3019 _192_/a_476_47# _049_ 1.44e-19
C3020 _322_/a_543_47# _205_/a_27_47# 0.00358f
C3021 net44 _226_/a_27_47# 4.7e-21
C3022 _311_/a_1283_21# _202_/a_79_21# 5.95e-21
C3023 cal_itt\[0\] net30 3.6e-20
C3024 _321_/a_193_47# _310_/a_1283_21# 3.21e-20
C3025 _321_/a_27_47# _310_/a_1108_47# 3.19e-20
C3026 net24 _042_ 1.88e-19
C3027 _178_/a_68_297# net18 0.00254f
C3028 VPWR _279_/a_204_297# -0.00176f
C3029 clknet_2_3__leaf_clk _118_ 5.75e-20
C3030 _331_/a_805_47# trim_mask\[4\] 1.36e-19
C3031 _306_/a_193_47# _204_/a_75_212# 5.35e-19
C3032 net52 _209_/a_27_47# 8.83e-19
C3033 VPWR _325_/a_651_413# 0.00142f
C3034 VPWR _216_/a_199_47# -3.48e-19
C3035 net13 _092_ 0.0585f
C3036 _317_/a_27_47# _014_ 0.0376f
C3037 _317_/a_193_47# clknet_2_0__leaf_clk 0.583f
C3038 _309_/a_1283_21# mask\[1\] 0.00327f
C3039 output25/a_27_47# _007_ 0.0163f
C3040 _264_/a_27_297# _108_ 0.00481f
C3041 _048_ _242_/a_382_297# 0.00132f
C3042 _189_/a_27_47# clone1/a_27_47# 4.91e-19
C3043 _325_/a_761_289# _046_ 0.00305f
C3044 _199_/a_109_297# _001_ 8.77e-19
C3045 _028_ net19 0.00127f
C3046 _333_/a_193_47# _175_/a_68_297# 8.23e-20
C3047 _104_ clkbuf_2_3__f_clk/a_110_47# 1.77e-19
C3048 _327_/a_1217_47# net18 5.39e-20
C3049 _315_/a_27_47# net30 8.1e-21
C3050 net13 _169_/a_109_53# 0.00396f
C3051 mask\[7\] _314_/a_27_47# 1.54e-19
C3052 _041_ net40 5.18e-22
C3053 net10 net50 0.0105f
C3054 _265_/a_81_21# _333_/a_193_47# 2.14e-21
C3055 VPWR _248_/a_373_47# -4.25e-19
C3056 trim[4] net34 0.0953f
C3057 ctlp[6] ctlp[5] 1.96e-20
C3058 _320_/a_1108_47# _208_/a_76_199# 6.13e-20
C3059 net12 _306_/a_651_413# 0.00178f
C3060 _030_ _173_/a_27_47# 1.16e-20
C3061 net50 clknet_2_2__leaf_clk 0.0136f
C3062 _203_/a_59_75# _072_ 0.00556f
C3063 _203_/a_145_75# cal_itt\[3\] 0.00121f
C3064 _325_/a_805_47# net43 -0.00123f
C3065 _320_/a_193_47# _017_ 0.0979f
C3066 _308_/a_27_47# output30/a_27_47# 3.05e-21
C3067 cal_itt\[0\] _072_ 0.00264f
C3068 cal_itt\[1\] cal_itt\[3\] 0.00338f
C3069 net22 _315_/a_27_47# 2.45e-20
C3070 net51 _206_/a_27_93# 8.31e-21
C3071 _043_ _311_/a_1108_47# 2.32e-20
C3072 _107_ _028_ 7.9e-19
C3073 trim_mask\[1\] _336_/a_27_47# 4.07e-20
C3074 _309_/a_448_47# _082_ 1.16e-19
C3075 _333_/a_448_47# clknet_2_2__leaf_clk 1.96e-20
C3076 trim[1] net32 0.146f
C3077 clknet_2_1__leaf_clk _319_/a_543_47# 6.88e-19
C3078 _083_ _209_/a_27_47# 1.29e-20
C3079 net45 _049_ 0.00196f
C3080 _308_/a_1108_47# fanout43/a_27_47# 0.00423f
C3081 net13 mask\[5\] 9.08e-20
C3082 _318_/a_761_289# net45 1.29e-19
C3083 net8 _272_/a_81_21# 0.00281f
C3084 clknet_2_0__leaf_clk net30 1.38f
C3085 state\[2\] net13 0.127f
C3086 _306_/a_651_413# net44 8.36e-19
C3087 _326_/a_543_47# _023_ 0.00108f
C3088 _326_/a_1283_21# _102_ 0.00375f
C3089 _326_/a_1108_47# mask\[7\] 0.0213f
C3090 net43 _092_ 2.25e-20
C3091 clk _027_ 0.00154f
C3092 VPWR net36 0.114f
C3093 VPWR _044_ 0.289f
C3094 net1 output41/a_27_47# 0.189f
C3095 _213_/a_109_297# _080_ 0.00379f
C3096 _048_ trim_mask\[4\] 2.84e-20
C3097 _097_ _315_/a_1283_21# 7.8e-21
C3098 clkbuf_2_2__f_clk/a_110_47# _330_/a_651_413# 2.2e-19
C3099 _286_/a_76_199# _338_/a_476_47# 0.00437f
C3100 _103_ _049_ 0.0125f
C3101 net2 _067_ 3.42e-19
C3102 _047_ _332_/a_1283_21# 1.23e-20
C3103 _324_/a_761_289# mask\[5\] 2.14e-19
C3104 net2 _070_ 0.38f
C3105 _059_ _098_ 1.04e-19
C3106 _340_/a_1032_413# cal_count\[0\] 2.03e-20
C3107 _305_/a_1283_21# _067_ 2.17e-19
C3108 _305_/a_1283_21# _070_ 0.00139f
C3109 _328_/a_1217_47# net9 1.84e-20
C3110 _065_ _049_ 0.339f
C3111 _125_ _129_ 0.00637f
C3112 _187_/a_297_47# _136_ 1.17e-19
C3113 net22 clknet_2_0__leaf_clk 0.0104f
C3114 _320_/a_27_47# net15 4.44e-21
C3115 net12 _052_ 0.00248f
C3116 VPWR _327_/a_448_47# 0.00283f
C3117 _307_/a_27_47# sample 0.00361f
C3118 net4 _027_ 2.02e-19
C3119 _136_ _332_/a_761_289# 2.34e-20
C3120 _059_ clknet_0_clk 0.0276f
C3121 _105_ _049_ 0.00221f
C3122 _074_ _313_/a_1283_21# 3.85e-19
C3123 _232_/a_32_297# net55 0.0307f
C3124 net9 cal_count\[2\] 1.69e-20
C3125 state\[2\] _331_/a_193_47# 1.43e-20
C3126 clknet_2_2__leaf_clk _279_/a_396_47# 5.22e-19
C3127 net4 _195_/a_218_47# 7.62e-19
C3128 _325_/a_1108_47# _019_ 2.67e-19
C3129 _322_/a_805_47# mask\[3\] 4.33e-20
C3130 mask\[1\] _016_ 0.00126f
C3131 trim_mask\[2\] _334_/a_193_47# 0.00989f
C3132 fanout46/a_27_47# _033_ 0.0622f
C3133 output25/a_27_47# result[4] 0.0022f
C3134 result[3] output26/a_27_47# 1.88e-20
C3135 _319_/a_27_47# _049_ 0.0011f
C3136 _104_ cal_count\[3\] 1.88e-20
C3137 _324_/a_27_47# net27 2.02e-19
C3138 _305_/a_193_47# clkbuf_0_clk/a_110_47# 0.00157f
C3139 mask\[7\] _314_/a_1217_47# 6.99e-20
C3140 _125_ _339_/a_1032_413# 1.43e-20
C3141 output33/a_27_47# _056_ 0.171f
C3142 _312_/a_761_289# _045_ 6.66e-20
C3143 _100_ _170_/a_299_297# 8.93e-20
C3144 _243_/a_109_297# _049_ 0.00162f
C3145 trim_val\[0\] _333_/a_448_47# 5.91e-20
C3146 net18 net40 0.0116f
C3147 net12 _311_/a_27_47# 7.12e-21
C3148 _064_ _257_/a_109_47# 0.00344f
C3149 _104_ _257_/a_27_297# 0.0807f
C3150 net19 _279_/a_314_297# 0.00139f
C3151 _104_ _331_/a_27_47# 1.07e-19
C3152 net43 mask\[5\] 2.36e-21
C3153 _239_/a_694_21# _100_ 0.0016f
C3154 _306_/a_1108_47# clknet_0_clk 3.47e-19
C3155 _019_ _248_/a_109_297# 0.00723f
C3156 _129_ net40 0.083f
C3157 net48 net33 1.38e-20
C3158 _260_/a_93_21# _092_ 1.12e-20
C3159 _227_/a_209_311# net55 0.0362f
C3160 _246_/a_27_297# _101_ 0.0635f
C3161 _080_ _212_/a_113_297# 0.00838f
C3162 output37/a_27_47# net37 0.0225f
C3163 _273_/a_59_75# net46 0.0121f
C3164 trim_mask\[1\] _336_/a_1217_47# 2.91e-21
C3165 _127_ net33 0.0235f
C3166 net13 _017_ 9.55e-19
C3167 net45 _315_/a_1108_47# 0.0084f
C3168 _014_ _315_/a_448_47# 1.1e-21
C3169 _321_/a_193_47# _042_ 0.00809f
C3170 _019_ mask\[1\] 2.67e-20
C3171 _132_ cal_count\[2\] 0.00622f
C3172 _079_ _315_/a_27_47# 1.26e-20
C3173 _040_ mask\[2\] 0.0363f
C3174 _123_ _067_ 5.69e-19
C3175 clknet_0_clk _075_ 0.261f
C3176 net44 _311_/a_27_47# 0.0073f
C3177 _107_ _279_/a_314_297# 0.00207f
C3178 _048_ _283_/a_75_212# 8.48e-21
C3179 _321_/a_1108_47# clknet_2_1__leaf_clk 0.00232f
C3180 calibrate _316_/a_27_47# 2.84e-20
C3181 trim_mask\[0\] _332_/a_805_47# 8.96e-19
C3182 _336_/a_761_289# net30 2.25e-21
C3183 _258_/a_27_297# fanout46/a_27_47# 2.53e-20
C3184 _115_ _334_/a_193_47# 0.00186f
C3185 _093_ clone7/a_27_47# 3.26e-20
C3186 _339_/a_1032_413# net40 2.31e-19
C3187 net12 calibrate 0.0079f
C3188 VPWR _208_/a_505_21# 0.00607f
C3189 _340_/a_652_21# _123_ 0.0316f
C3190 clknet_2_1__leaf_clk _313_/a_193_47# 0.596f
C3191 _189_/a_27_47# _051_ 0.0288f
C3192 net54 _090_ 0.259f
C3193 clkbuf_2_2__f_clk/a_110_47# net46 0.0262f
C3194 cal_count\[0\] _338_/a_476_47# 0.00994f
C3195 clone1/a_27_47# net30 5.12e-21
C3196 _327_/a_27_47# _265_/a_81_21# 1.9e-21
C3197 VPWR mask\[2\] 0.319f
C3198 _300_/a_47_47# _122_ 3.83e-19
C3199 cal_itt\[0\] _230_/a_59_75# 0.0479f
C3200 _074_ _081_ 0.0162f
C3201 _126_ net33 0.46f
C3202 _293_/a_81_21# _289_/a_68_297# 5.27e-19
C3203 _322_/a_1283_21# mask\[2\] 8.98e-21
C3204 _305_/a_27_47# _041_ 1.2e-20
C3205 _328_/a_193_47# _336_/a_1108_47# 2.05e-20
C3206 _093_ net4 2.32e-20
C3207 _058_ _333_/a_27_47# 0.00266f
C3208 net34 _108_ 0.00839f
C3209 _004_ _078_ 1.57e-20
C3210 net45 state\[1\] 0.104f
C3211 net54 _242_/a_382_297# 1.17e-20
C3212 trim[0] net34 0.105f
C3213 _062_ clknet_2_3__leaf_clk 0.177f
C3214 _079_ clknet_2_0__leaf_clk 0.0308f
C3215 _134_ net37 1.79e-20
C3216 VPWR output17/a_27_47# 0.0723f
C3217 VPWR _278_/a_27_47# 6.54e-19
C3218 mask\[7\] _146_/a_68_297# 2.69e-19
C3219 _327_/a_1108_47# clknet_2_2__leaf_clk 3.11e-19
C3220 _327_/a_27_47# trim_mask\[4\] 0.00152f
C3221 state\[2\] _260_/a_93_21# 0.00652f
C3222 _101_ _084_ 1.37e-19
C3223 _119_ _330_/a_193_47# 2.15e-19
C3224 _341_/a_193_47# _108_ 1.06e-19
C3225 _319_/a_1217_47# _049_ 5.28e-20
C3226 _313_/a_27_47# _009_ 1.71e-21
C3227 _041_ net51 4.43e-20
C3228 ctlp[1] _223_/a_109_297# 8.48e-19
C3229 _329_/a_543_47# net46 1.81e-19
C3230 VPWR _330_/a_1283_21# 0.0386f
C3231 net23 mask\[2\] 2.03e-20
C3232 net37 _130_ 0.0221f
C3233 mask\[5\] _312_/a_1108_47# 2.34e-20
C3234 net12 _305_/a_651_413# 3.15e-19
C3235 VPWR trim[4] 0.255f
C3236 _307_/a_1108_47# _094_ 3.31e-23
C3237 net3 _092_ 0.0901f
C3238 _229_/a_27_297# _226_/a_27_47# 1.02e-19
C3239 _313_/a_448_47# net29 1.76e-20
C3240 _337_/a_761_289# _049_ 0.00926f
C3241 _259_/a_27_297# trim_mask\[4\] 0.01f
C3242 cal_itt\[1\] _304_/a_448_47# 7.03e-20
C3243 _125_ _297_/a_47_47# 0.001f
C3244 _337_/a_27_47# net30 2.09e-19
C3245 trim_val\[1\] _172_/a_150_297# 0.00172f
C3246 trim_mask\[1\] _172_/a_68_297# 0.00653f
C3247 _314_/a_193_47# net14 0.0067f
C3248 _031_ net34 7.71e-23
C3249 _322_/a_27_47# net15 6.81e-20
C3250 _341_/a_639_47# net46 1.26e-19
C3251 net54 _048_ 0.0101f
C3252 _168_/a_207_413# net55 1.95e-21
C3253 mask\[2\] net52 0.333f
C3254 net4 _032_ 3.38e-21
C3255 _328_/a_193_47# _256_/a_27_297# 3.43e-19
C3256 _169_/a_109_53# net3 4.79e-20
C3257 _321_/a_193_47# _022_ 7.1e-19
C3258 mask\[1\] _205_/a_27_47# 9.85e-20
C3259 _319_/a_543_47# net45 6.88e-20
C3260 _319_/a_1108_47# clknet_2_0__leaf_clk 0.061f
C3261 _286_/a_535_374# clknet_2_3__leaf_clk 2.46e-19
C3262 _305_/a_651_413# net44 0.00382f
C3263 _051_ _227_/a_109_93# 0.00531f
C3264 net31 trimb[1] 0.109f
C3265 mask\[6\] _313_/a_761_289# 1.34e-21
C3266 net44 _311_/a_1217_47# -1.47e-19
C3267 state\[1\] _243_/a_109_297# 9.96e-21
C3268 net27 _312_/a_543_47# 2.14e-19
C3269 _053_ _260_/a_250_297# 0.00772f
C3270 _233_/a_373_47# _013_ 5.79e-20
C3271 _338_/a_27_47# _123_ 0.0015f
C3272 net28 _314_/a_27_47# 0.0118f
C3273 _064_ trim_val\[3\] 4.87e-20
C3274 _191_/a_27_297# net40 1.45e-19
C3275 _063_ _278_/a_27_47# 3.44e-19
C3276 _102_ net29 2.32e-20
C3277 _340_/a_1032_413# net16 8.39e-19
C3278 VPWR _306_/a_448_47# 0.00263f
C3279 _327_/a_1108_47# trim_val\[0\] 1.75e-21
C3280 _312_/a_448_47# _084_ 4.93e-20
C3281 _301_/a_47_47# _135_ 0.0423f
C3282 _301_/a_285_47# net2 3.31e-19
C3283 _297_/a_47_47# net40 0.015f
C3284 _187_/a_212_413# clknet_2_3__leaf_clk 8.26e-19
C3285 _178_/a_68_297# trim_mask\[4\] 2.49e-20
C3286 _241_/a_297_47# _099_ 0.0598f
C3287 VPWR _314_/a_193_47# 0.0233f
C3288 _341_/a_27_47# _135_ 1.04e-20
C3289 _069_ _072_ 4.94e-20
C3290 _058_ _333_/a_1217_47# 1.11e-19
C3291 cal net3 0.00534f
C3292 state\[2\] net3 6.86e-20
C3293 clk _171_/a_27_47# 0.0124f
C3294 net31 trimb[4] 0.109f
C3295 net42 _051_ 0.00681f
C3296 _308_/a_1283_21# _039_ 0.0101f
C3297 net12 _239_/a_27_297# 0.00146f
C3298 _319_/a_193_47# _319_/a_761_289# -0.0119f
C3299 _319_/a_27_47# _319_/a_543_47# -0.00936f
C3300 _185_/a_68_297# _095_ 5.79e-20
C3301 _007_ mask\[3\] 1.14e-19
C3302 _059_ _263_/a_79_21# 0.00233f
C3303 result[0] _074_ 0.0228f
C3304 _279_/a_206_47# trim_val\[4\] 0.0017f
C3305 _279_/a_314_297# _118_ 0.00906f
C3306 _088_ net41 1.32e-20
C3307 _339_/a_1182_261# cal_count\[0\] 0.065f
C3308 net8 ctln[2] 0.0038f
C3309 trim_val\[3\] _057_ 0.00755f
C3310 _065_ _202_/a_297_47# 2.28e-19
C3311 net4 _171_/a_27_47# 1.45e-20
C3312 fanout47/a_27_47# _287_/a_75_212# 1.92e-20
C3313 state\[0\] _166_/a_161_47# 2.4e-19
C3314 _214_/a_113_297# clknet_2_1__leaf_clk 2.91e-20
C3315 _305_/a_1108_47# clknet_0_clk 1.24e-19
C3316 _060_ _050_ 2.31e-19
C3317 _110_ _273_/a_59_75# 0.00312f
C3318 _282_/a_68_297# _049_ 0.0134f
C3319 _010_ net29 8.13e-20
C3320 _304_/a_1108_47# _065_ 0.00918f
C3321 net43 _314_/a_1283_21# 0.00325f
C3322 clk _317_/a_448_47# 0.00205f
C3323 _317_/a_193_47# _316_/a_1283_21# 1.12e-20
C3324 _317_/a_27_47# _316_/a_1108_47# 1.69e-20
C3325 net2 _339_/a_193_47# 4.56e-20
C3326 cal_itt\[0\] net47 0.279f
C3327 VPWR _195_/a_218_374# -0.00159f
C3328 VPWR _094_ 0.152f
C3329 _028_ _330_/a_761_289# 5.82e-23
C3330 clknet_2_2__leaf_clk _330_/a_543_47# 0.0413f
C3331 _257_/a_109_297# net46 5.48e-21
C3332 _209_/a_27_47# _208_/a_76_199# 5.06e-20
C3333 _051_ _054_ 0.0162f
C3334 _314_/a_1462_47# net14 2.52e-19
C3335 VPWR _326_/a_448_47# 0.00366f
C3336 _329_/a_448_47# _031_ 3.97e-20
C3337 VPWR _334_/a_448_47# 0.00341f
C3338 _051_ net30 0.705f
C3339 _189_/a_408_47# clknet_0_clk 0.0319f
C3340 VPWR _088_ 0.502f
C3341 _290_/a_207_413# net34 0.0122f
C3342 _106_ _262_/a_205_47# 6.6e-20
C3343 _328_/a_27_47# _258_/a_27_297# 1.75e-19
C3344 _328_/a_27_47# _024_ 0.00115f
C3345 _320_/a_193_47# clknet_2_1__leaf_clk 1.11e-20
C3346 _266_/a_68_297# _062_ 3.65e-20
C3347 net15 net21 1.66e-20
C3348 clk _203_/a_145_75# 9.6e-19
C3349 _238_/a_75_212# _316_/a_193_47# 2.94e-19
C3350 _110_ clkbuf_2_2__f_clk/a_110_47# 0.0083f
C3351 _331_/a_543_47# _052_ 2.78e-21
C3352 net12 _203_/a_59_75# 2.86e-19
C3353 net43 _310_/a_27_47# 0.0147f
C3354 VPWR _286_/a_439_47# -4.05e-19
C3355 _340_/a_1602_47# _132_ 6.93e-20
C3356 _330_/a_1108_47# net19 9.02e-20
C3357 _325_/a_193_47# net27 9.9e-20
C3358 net50 _278_/a_27_47# 1.62e-19
C3359 cal_itt\[1\] clk 1.25e-20
C3360 _308_/a_805_47# _074_ 6.63e-19
C3361 _168_/a_27_413# _051_ 0.0374f
C3362 _321_/a_651_413# clknet_2_0__leaf_clk 4.04e-20
C3363 _303_/a_543_47# _068_ 0.0027f
C3364 _274_/a_75_212# _112_ 4.98e-19
C3365 _335_/a_193_47# _119_ 1.36e-20
C3366 net2 trimb[4] 1.08e-19
C3367 _324_/a_27_47# _311_/a_1283_21# 2.45e-20
C3368 _074_ net14 0.926f
C3369 _229_/a_27_297# _052_ 3.29e-20
C3370 result[0] output23/a_27_47# 1.11e-20
C3371 output22/a_27_47# result[1] 0.00288f
C3372 _182_/a_27_47# net35 0.00288f
C3373 net2 clknet_2_3__leaf_clk 0.106f
C3374 _337_/a_651_413# clknet_2_0__leaf_clk 1.08e-20
C3375 VPWR _335_/a_1283_21# 0.0165f
C3376 _323_/a_27_47# net26 4.04e-19
C3377 result[6] _314_/a_639_47# 3.88e-19
C3378 net28 _314_/a_1217_47# 2.55e-20
C3379 _107_ _226_/a_27_47# 0.00327f
C3380 _263_/a_79_21# _075_ 0.00358f
C3381 _309_/a_1108_47# _310_/a_1108_47# 1.55e-20
C3382 _323_/a_1283_21# _042_ 0.0354f
C3383 _237_/a_535_374# _093_ 7.79e-20
C3384 trim_mask\[3\] _330_/a_1108_47# 6.69e-19
C3385 _167_/a_161_47# net45 0.00532f
C3386 ctlp[6] _009_ 2.05e-20
C3387 _098_ _170_/a_81_21# 1.2e-21
C3388 net44 _203_/a_59_75# 1.65e-19
C3389 cal_itt\[1\] net4 0.407f
C3390 VPWR _314_/a_1462_47# 0.00178f
C3391 _265_/a_81_21# net40 1.62e-20
C3392 ctln[4] _275_/a_299_297# 0.00151f
C3393 VPWR _332_/a_543_47# 0.0113f
C3394 VPWR _108_ 1.23f
C3395 _051_ _072_ 8.19e-19
C3396 _059_ _236_/a_109_297# 4.7e-21
C3397 _074_ _040_ 4.02e-21
C3398 _337_/a_1108_47# _065_ 9.33e-19
C3399 _074_ net41 2.02e-19
C3400 _012_ output41/a_27_47# 9.78e-19
C3401 _303_/a_193_47# net2 1.18e-20
C3402 _110_ _329_/a_543_47# 9.34e-19
C3403 result[4] _007_ 7.64e-20
C3404 VPWR _244_/a_27_297# 0.063f
C3405 trim[0] VPWR 0.225f
C3406 net9 _041_ 0.00973f
C3407 _304_/a_27_47# _066_ 2.59e-21
C3408 net9 _338_/a_1182_261# 0.0012f
C3409 net24 _143_/a_68_297# 0.00693f
C3410 trim_mask\[2\] trim_val\[2\] 0.162f
C3411 _336_/a_193_47# _264_/a_27_297# 1.49e-21
C3412 result[1] _308_/a_1283_21# 1.68e-19
C3413 mask\[7\] _078_ 0.271f
C3414 _281_/a_103_199# _092_ 0.0118f
C3415 _281_/a_337_297# _095_ 0.00157f
C3416 _304_/a_193_47# _304_/a_448_47# -0.00373f
C3417 _339_/a_193_47# _123_ 0.017f
C3418 _200_/a_80_21# clkbuf_2_3__f_clk/a_110_47# 0.00682f
C3419 _249_/a_109_47# mask\[5\] 9.26e-19
C3420 VPWR _310_/a_1270_413# -1.62e-19
C3421 VPWR _074_ 2.52f
C3422 _003_ _203_/a_59_75# 4.94e-20
C3423 trim_mask\[4\] net40 0.00108f
C3424 _117_ net18 8.86e-19
C3425 _340_/a_381_47# cal_count\[2\] 1.81e-20
C3426 ctln[1] VPWR 0.00266f
C3427 _275_/a_81_21# _335_/a_193_47# 0.00133f
C3428 _275_/a_299_297# _335_/a_27_47# 1.03e-19
C3429 trim_mask\[2\] net16 0.0178f
C3430 _337_/a_193_47# _319_/a_1283_21# 3.92e-20
C3431 _337_/a_27_47# _319_/a_1108_47# 3.29e-20
C3432 _050_ en_co_clk 0.112f
C3433 cal_itt\[1\] _122_ 1.33e-20
C3434 ctlp[1] _010_ 0.00232f
C3435 _100_ net55 0.253f
C3436 output10/a_27_47# net46 1.46e-20
C3437 _322_/a_1283_21# _074_ 0.00292f
C3438 cal_itt\[1\] _073_ 4.66e-20
C3439 clknet_2_0__leaf_clk _316_/a_27_47# 0.0349f
C3440 clk _014_ 0.0041f
C3441 state\[0\] _185_/a_68_297# 0.0685f
C3442 cal_itt\[0\] _341_/a_27_47# 1.88e-19
C3443 _025_ net46 0.0067f
C3444 net12 clknet_2_0__leaf_clk 1.37e-19
C3445 _026_ _031_ 1.79e-20
C3446 VPWR _031_ 0.104f
C3447 net27 _007_ 2.83e-20
C3448 _101_ _311_/a_193_47# 4.59e-21
C3449 calibrate _229_/a_27_297# 0.0647f
C3450 _064_ trim_val\[4\] 0.0378f
C3451 _123_ clknet_2_3__leaf_clk 0.156f
C3452 _327_/a_805_47# _058_ 4.69e-19
C3453 _104_ _327_/a_193_47# 1.35e-19
C3454 mask\[1\] _208_/a_218_374# 1.34e-19
C3455 _330_/a_1108_47# _279_/a_27_47# 5.98e-21
C3456 output24/a_27_47# _006_ 0.00974f
C3457 net27 _249_/a_27_297# 4e-20
C3458 _334_/a_1108_47# clknet_2_2__leaf_clk 8.02e-20
C3459 _304_/a_1283_21# _035_ 1.83e-21
C3460 _052_ _260_/a_256_47# 0.00327f
C3461 _306_/a_193_47# _050_ 1.23e-21
C3462 net43 _310_/a_1217_47# 9.72e-19
C3463 _311_/a_1270_413# net53 4.26e-20
C3464 net27 mask\[3\] 1.52e-20
C3465 net13 clknet_2_1__leaf_clk 7.95e-20
C3466 net23 _074_ 0.211f
C3467 _063_ _108_ 6.65e-19
C3468 net4 _014_ 5.39e-20
C3469 VPWR _247_/a_109_47# -0.00104f
C3470 mask\[0\] _121_ 0.00291f
C3471 _115_ trim_val\[2\] 0.0012f
C3472 _324_/a_193_47# _250_/a_27_297# 2.84e-19
C3473 _047_ net33 0.0023f
C3474 VPWR output23/a_27_47# 0.0236f
C3475 _104_ _058_ 0.00402f
C3476 _259_/a_373_47# _064_ 8.77e-19
C3477 _259_/a_109_297# _104_ 0.00431f
C3478 output28/a_27_47# clknet_2_1__leaf_clk 0.0131f
C3479 net44 clknet_2_0__leaf_clk 0.173f
C3480 _126_ output40/a_27_47# 0.0463f
C3481 VPWR _305_/a_448_47# 0.00286f
C3482 VPWR _311_/a_805_47# 1.18e-19
C3483 _052_ net19 2.02e-21
C3484 VPWR _146_/a_150_297# -6.23e-19
C3485 _324_/a_761_289# clknet_2_1__leaf_clk 4.73e-19
C3486 _329_/a_193_47# net9 0.0159f
C3487 _115_ net16 0.013f
C3488 mask\[3\] rebuffer5/a_161_47# 1.65e-21
C3489 _179_/a_27_47# _176_/a_27_47# 1.77e-20
C3490 _056_ _172_/a_68_297# 3.39e-19
C3491 _074_ net52 0.0103f
C3492 _335_/a_543_47# clknet_2_2__leaf_clk 1.7e-19
C3493 _276_/a_59_75# _119_ 6.99e-22
C3494 net15 _241_/a_105_352# 0.00353f
C3495 _333_/a_543_47# net46 0.0208f
C3496 _243_/a_27_297# clone7/a_27_47# 0.0806f
C3497 _322_/a_193_47# clknet_2_1__leaf_clk 9.42e-19
C3498 _304_/a_1270_413# _067_ 8.41e-20
C3499 clknet_2_0__leaf_clk _003_ 0.00196f
C3500 net9 net18 0.0456f
C3501 net9 _341_/a_651_413# 3.15e-19
C3502 _337_/a_1283_21# _206_/a_27_93# 0.00185f
C3503 _336_/a_1108_47# _033_ 1.94e-21
C3504 net34 output5/a_27_47# 0.00396f
C3505 net27 _220_/a_113_297# 0.0022f
C3506 _332_/a_761_289# clknet_2_2__leaf_clk 2.34e-19
C3507 output23/a_27_47# net23 0.023f
C3508 _120_ _092_ 0.076f
C3509 net16 net38 0.0476f
C3510 _304_/a_27_47# net47 0.00459f
C3511 _107_ _052_ 0.0314f
C3512 _071_ clkbuf_2_3__f_clk/a_110_47# 0.00225f
C3513 _311_/a_27_47# net19 7.96e-22
C3514 net43 _305_/a_639_47# -7.75e-19
C3515 output13/a_27_47# _318_/a_543_47# 1.95e-19
C3516 net16 _339_/a_1182_261# 8.18e-19
C3517 _136_ clkc 5.39e-20
C3518 _308_/a_193_47# mask\[0\] 3.45e-20
C3519 _308_/a_27_47# _078_ 0.00772f
C3520 _308_/a_761_289# net22 1.74e-19
C3521 _321_/a_193_47# _321_/a_448_47# -0.00373f
C3522 net24 _214_/a_199_47# 4.81e-19
C3523 _340_/a_27_47# _340_/a_652_21# -0.00438f
C3524 net50 _335_/a_1283_21# 0.00823f
C3525 trim_mask\[3\] _335_/a_1108_47# 0.00393f
C3526 net4 _243_/a_27_297# 3.76e-21
C3527 net26 net14 0.00702f
C3528 _308_/a_193_47# output24/a_27_47# 1.55e-19
C3529 _247_/a_109_47# net52 0.00475f
C3530 _262_/a_27_47# clkbuf_2_3__f_clk/a_110_47# 0.00344f
C3531 VPWR _232_/a_220_297# -4.59e-19
C3532 _186_/a_109_297# net54 1.18e-20
C3533 _292_/a_493_297# _123_ 4.54e-20
C3534 net43 clknet_2_1__leaf_clk 0.304f
C3535 clkbuf_0_clk/a_110_47# _202_/a_297_47# 6.77e-20
C3536 _014_ _316_/a_805_47# 3.89e-19
C3537 net45 _316_/a_639_47# -3.61e-19
C3538 _078_ clknet_0_clk 3.17e-20
C3539 _092_ _076_ 4.94e-20
C3540 VPWR net49 0.198f
C3541 VPWR _272_/a_81_21# 0.0334f
C3542 _327_/a_27_47# net40 8.8e-20
C3543 clkbuf_0_clk/a_110_47# _304_/a_1108_47# 4.44e-19
C3544 _320_/a_1108_47# _078_ 8.98e-19
C3545 VPWR _290_/a_207_413# 0.00668f
C3546 _320_/a_193_47# net45 4.53e-20
C3547 _320_/a_543_47# clknet_2_0__leaf_clk 0.0014f
C3548 net50 _108_ 0.13f
C3549 VPWR _170_/a_299_297# 0.0249f
C3550 net9 _339_/a_1032_413# 7.41e-19
C3551 _083_ _074_ 0.0151f
C3552 output36/a_27_47# net34 0.0153f
C3553 trim[1] _265_/a_299_297# 7.76e-20
C3554 _162_/a_27_47# net32 5.19e-19
C3555 _326_/a_27_47# _007_ 0.00105f
C3556 _030_ clknet_2_2__leaf_clk 0.179f
C3557 VPWR _239_/a_694_21# -0.00501f
C3558 _238_/a_75_212# net14 2.88e-21
C3559 _291_/a_285_47# cal_count\[0\] 0.00164f
C3560 _255_/a_27_47# clknet_0_clk 9.47e-19
C3561 _097_ _237_/a_505_21# 2.46e-19
C3562 net4 _336_/a_543_47# 0.0072f
C3563 output34/a_27_47# net46 8.6e-19
C3564 _324_/a_543_47# mask\[6\] 7.79e-22
C3565 _324_/a_27_47# _021_ 0.146f
C3566 _129_ _132_ 0.0828f
C3567 _062_ _095_ 4.99e-20
C3568 _324_/a_1108_47# net26 1.04e-19
C3569 _304_/a_193_47# net4 8.89e-21
C3570 VPWR _227_/a_368_53# -3.12e-19
C3571 _326_/a_193_47# net25 1.29e-19
C3572 _291_/a_35_297# net2 5.01e-19
C3573 _320_/a_193_47# _065_ 4.41e-20
C3574 _019_ _247_/a_27_297# 9.77e-21
C3575 _307_/a_1270_413# net22 2.15e-19
C3576 _307_/a_651_413# mask\[0\] 1.44e-20
C3577 _064_ _330_/a_193_47# 2.68e-21
C3578 VPWR _002_ 0.0886f
C3579 VPWR net26 2.11f
C3580 trim_val\[0\] _332_/a_761_289# 0.00308f
C3581 _307_/a_761_289# net45 1.39e-20
C3582 _307_/a_1283_21# clknet_2_0__leaf_clk 3.93e-19
C3583 VPWR _289_/a_68_297# 0.0258f
C3584 net47 _069_ 3.22e-19
C3585 _058_ _267_/a_59_75# 0.00906f
C3586 trim[3] _334_/a_543_47# 2.57e-20
C3587 _156_/a_27_47# _084_ 0.00229f
C3588 VPWR _317_/a_1283_21# 0.00805f
C3589 _238_/a_75_212# net41 1.43e-19
C3590 _060_ _226_/a_303_47# 1.78e-19
C3591 calibrate _107_ 0.0534f
C3592 _328_/a_27_47# _257_/a_27_297# 2.44e-19
C3593 _322_/a_1283_21# net26 0.00125f
C3594 _192_/a_174_21# net41 2.35e-21
C3595 _251_/a_27_297# _046_ 5.07e-19
C3596 _298_/a_78_199# _131_ 0.00179f
C3597 _298_/a_215_47# cal_count\[2\] 0.0222f
C3598 net27 _222_/a_113_297# 2.1e-19
C3599 _304_/a_639_47# _136_ 2.96e-19
C3600 output38/a_27_47# output39/a_27_47# 0.0523f
C3601 ctln[2] net34 0.00136f
C3602 _304_/a_193_47# _122_ 0.00922f
C3603 _053_ _330_/a_193_47# 1.33e-19
C3604 _083_ _311_/a_805_47# 1.62e-20
C3605 _110_ output10/a_27_47# 4.1e-20
C3606 _274_/a_75_212# net33 7.24e-21
C3607 clknet_2_3__leaf_clk _150_/a_27_47# 6.4e-22
C3608 net12 _337_/a_27_47# 1.79e-21
C3609 VPWR _238_/a_75_212# 0.0485f
C3610 _134_ cal_count\[2\] 0.0359f
C3611 _269_/a_299_297# _333_/a_761_289# 2.18e-19
C3612 _304_/a_1217_47# net47 1.99e-19
C3613 VPWR _192_/a_174_21# 0.00833f
C3614 _341_/a_27_47# _304_/a_27_47# 4.05e-20
C3615 cal_itt\[2\] VPWR 0.365f
C3616 _258_/a_27_297# _256_/a_27_297# 1.26e-20
C3617 _256_/a_373_47# trim_mask\[0\] 2.23e-19
C3618 _256_/a_27_297# _024_ 0.0129f
C3619 fanout47/a_27_47# clknet_0_clk 3.52e-21
C3620 _340_/a_476_47# net47 0.0015f
C3621 _037_ _304_/a_193_47# 8.53e-19
C3622 _060_ _235_/a_79_21# 7.13e-20
C3623 net13 _318_/a_805_47# 5.87e-19
C3624 cal_itt\[0\] _198_/a_181_47# 4.2e-20
C3625 cal_itt\[1\] _198_/a_109_47# 4.34e-19
C3626 _108_ _279_/a_396_47# 0.0356f
C3627 _308_/a_1462_47# mask\[0\] 4.24e-19
C3628 _308_/a_1217_47# _078_ 3.07e-19
C3629 net43 _210_/a_113_297# 1.58e-19
C3630 trim_val\[3\] _032_ 2.72e-19
C3631 _030_ trim_val\[0\] 0.00101f
C3632 clknet_2_1__leaf_clk _312_/a_1108_47# 1.32e-19
C3633 _262_/a_27_47# cal_count\[3\] 4.56e-19
C3634 _308_/a_639_47# clknet_2_0__leaf_clk 1.44e-19
C3635 result[6] result[7] 0.0507f
C3636 _130_ cal_count\[2\] 0.15f
C3637 _007_ _310_/a_761_289# 0.00229f
C3638 _308_/a_27_47# _004_ 2.88e-20
C3639 _217_/a_109_297# _074_ 0.00223f
C3640 net42 _087_ 2.68e-20
C3641 net35 _161_/a_68_297# 2.12e-19
C3642 _309_/a_543_47# _078_ 0.00886f
C3643 _309_/a_1283_21# mask\[0\] 1.94e-19
C3644 _094_ _034_ 0.0183f
C3645 clk _106_ 1.91e-20
C3646 _119_ _054_ 0.00224f
C3647 _002_ net52 2.54e-20
C3648 _237_/a_218_374# net45 8.89e-20
C3649 _074_ _155_/a_150_297# 5.4e-19
C3650 mask\[6\] _101_ 0.369f
C3651 _309_/a_27_47# net24 0.0466f
C3652 _237_/a_535_374# _014_ 1.51e-20
C3653 _337_/a_27_47# net44 0.00213f
C3654 _058_ net37 3.24e-19
C3655 cal_itt\[0\] _303_/a_639_47# 1.44e-19
C3656 _071_ _303_/a_448_47# 6.22e-20
C3657 _336_/a_27_47# clknet_0_clk 0.0028f
C3658 _336_/a_1283_21# clkbuf_2_2__f_clk/a_110_47# 0.0067f
C3659 net52 net26 0.0105f
C3660 _119_ net30 6.18e-19
C3661 mask\[0\] _245_/a_109_297# 0.00491f
C3662 _078_ _245_/a_27_297# 6.43e-20
C3663 _181_/a_150_297# _108_ 5.77e-19
C3664 VPWR _318_/a_651_413# -0.00632f
C3665 net25 _310_/a_543_47# 8.59e-19
C3666 _082_ _310_/a_27_47# 1.67e-19
C3667 trim_mask\[1\] clknet_2_2__leaf_clk 0.374f
C3668 net21 _009_ 5.24e-21
C3669 _327_/a_761_289# net46 0.004f
C3670 net13 net45 0.226f
C3671 _035_ _338_/a_1032_413# 4.03e-20
C3672 net28 _078_ 0.0029f
C3673 _339_/a_1602_47# cal_count\[2\] 8.14e-20
C3674 _306_/a_27_47# rebuffer5/a_161_47# 0.0041f
C3675 _324_/a_1217_47# _021_ 2.14e-20
C3676 cal_count\[1\] _289_/a_150_297# 0.00101f
C3677 _321_/a_1283_21# _041_ 9.15e-20
C3678 output35/a_27_47# net40 0.0147f
C3679 net4 _106_ 0.0182f
C3680 _328_/a_651_413# VPWR -0.00924f
C3681 _330_/a_193_47# _330_/a_448_47# -0.00297f
C3682 _277_/a_75_212# VPWR 0.0702f
C3683 _208_/a_535_374# _077_ 2.83e-20
C3684 _208_/a_218_47# _076_ 0.00129f
C3685 _164_/a_161_47# _317_/a_1283_21# 7.1e-20
C3686 _074_ _248_/a_109_47# 4.39e-19
C3687 cal_itt\[2\] _063_ 0.208f
C3688 net13 _065_ 0.058f
C3689 _028_ _227_/a_209_311# 6.9e-20
C3690 _307_/a_448_47# _004_ 0.00455f
C3691 _096_ _098_ 4.83e-19
C3692 VPWR ctlp[2] 0.101f
C3693 _315_/a_805_47# net14 5.85e-19
C3694 _136_ _284_/a_68_297# 0.00218f
C3695 _322_/a_1108_47# _078_ 0.0161f
C3696 cal_count\[3\] wire42/a_75_212# 2.12e-20
C3697 trim_mask\[0\] clk 0.00535f
C3698 _104_ _228_/a_297_47# 0.03f
C3699 _080_ clknet_2_1__leaf_clk 5.41e-19
C3700 _319_/a_651_413# clknet_0_clk 3.18e-19
C3701 _078_ _159_/a_27_47# 0.0319f
C3702 _125_ net40 0.227f
C3703 _322_/a_193_47# net45 5.96e-21
C3704 _266_/a_150_297# net30 0.00133f
C3705 net45 _331_/a_193_47# 0.00447f
C3706 _242_/a_79_21# _049_ 0.0147f
C3707 _326_/a_27_47# net27 0.00215f
C3708 _287_/a_75_212# _339_/a_27_47# 2.52e-21
C3709 trimb[0] net38 0.00705f
C3710 _185_/a_68_297# calibrate 5.21e-20
C3711 _325_/a_27_47# _251_/a_27_297# 0.00122f
C3712 VPWR output5/a_27_47# 0.0888f
C3713 _341_/a_193_47# _067_ 2.28e-20
C3714 clknet_0_clk _096_ 0.0288f
C3715 _325_/a_193_47# _250_/a_109_297# 6.47e-20
C3716 _164_/a_161_47# _192_/a_174_21# 1.47e-20
C3717 _083_ net26 0.143f
C3718 mask\[6\] _312_/a_448_47# 2.83e-21
C3719 result[3] _078_ 3.52e-19
C3720 _297_/a_47_47# _132_ 0.0162f
C3721 _021_ _312_/a_543_47# 2.75e-20
C3722 _340_/a_1182_261# _122_ 0.00579f
C3723 net13 _319_/a_27_47# 1.88e-21
C3724 trim_val\[1\] _333_/a_1270_413# 1.87e-19
C3725 trim_mask\[1\] _333_/a_651_413# 0.00123f
C3726 net47 _338_/a_193_47# 0.306f
C3727 trim[1] _058_ 0.00145f
C3728 _235_/a_79_21# en_co_clk 0.00618f
C3729 net15 en_co_clk 0.00947f
C3730 net12 _051_ 0.23f
C3731 _107_ _170_/a_384_47# 8.79e-20
C3732 _315_/a_1270_413# valid 2.99e-20
C3733 _340_/a_1224_47# net47 3.38e-21
C3734 _198_/a_27_47# _065_ 2.44e-19
C3735 net13 _243_/a_109_297# 0.00326f
C3736 _325_/a_543_47# clknet_2_1__leaf_clk 0.00214f
C3737 trim_mask\[0\] net4 0.0222f
C3738 _064_ _335_/a_193_47# 5e-19
C3739 _327_/a_1108_47# _108_ 1.55e-19
C3740 _340_/a_1182_261# _037_ 0.00151f
C3741 _239_/a_27_297# _107_ 0.00349f
C3742 _005_ result[2] 4.79e-21
C3743 VPWR _270_/a_145_75# 0.00144f
C3744 net43 net45 0.378f
C3745 _327_/a_1283_21# _111_ 0.0362f
C3746 net16 _333_/a_27_47# 0.0152f
C3747 mask\[3\] net51 4.53e-21
C3748 result[4] _310_/a_761_289# 2.56e-19
C3749 output26/a_27_47# _074_ 1.55e-19
C3750 mask\[4\] _311_/a_543_47# 0.0356f
C3751 _090_ _192_/a_639_47# 1.09e-19
C3752 VPWR _315_/a_805_47# 4.89e-19
C3753 _226_/a_27_47# _062_ 0.0104f
C3754 _071_ _000_ 1.61e-20
C3755 _313_/a_1283_21# _010_ 2.58e-19
C3756 _291_/a_117_297# _127_ 9.99e-20
C3757 net35 _332_/a_1108_47# 0.00429f
C3758 VPWR output36/a_27_47# 0.139f
C3759 mask\[0\] _016_ 0.0328f
C3760 _058_ _332_/a_651_413# 9.61e-19
C3761 _334_/a_543_47# _057_ 1.22e-19
C3762 _293_/a_299_297# _339_/a_27_47# 3.38e-20
C3763 _233_/a_373_47# net1 0.00105f
C3764 _074_ input1/a_75_212# 0.00827f
C3765 _058_ fanout46/a_27_47# 1.08e-19
C3766 _051_ net44 0.00365f
C3767 net24 _101_ 0.00937f
C3768 cal_itt\[0\] net19 0.0181f
C3769 _291_/a_285_47# net16 5.96e-19
C3770 net43 _065_ 0.0751f
C3771 cal_itt\[0\] _231_/a_161_47# 0.0693f
C3772 clkbuf_2_0__f_clk/a_110_47# _092_ 0.0808f
C3773 _340_/a_27_47# _339_/a_193_47# 0.00117f
C3774 _340_/a_193_47# _339_/a_27_47# 0.00126f
C3775 _294_/a_68_297# net37 8.7e-20
C3776 _256_/a_109_297# net18 0.00587f
C3777 clk _316_/a_1108_47# 5.5e-19
C3778 en_co_clk net37 1.95e-19
C3779 _297_/a_377_297# cal_count\[2\] 5.95e-20
C3780 _330_/a_27_47# net46 -2.05e-19
C3781 _330_/a_193_47# _027_ 0.522f
C3782 output14/a_27_47# _314_/a_761_289# 0.00321f
C3783 _293_/a_81_21# trimb[4] 9.37e-20
C3784 _128_ cal_count\[2\] 0.00309f
C3785 net43 _319_/a_27_47# 0.00142f
C3786 cal_itt\[0\] _107_ 3.22e-19
C3787 _168_/a_207_413# _028_ 0.00369f
C3788 _291_/a_117_297# _126_ 7.6e-19
C3789 _144_/a_27_47# _339_/a_193_47# 3.33e-21
C3790 _058_ _269_/a_299_297# 6.04e-19
C3791 _323_/a_543_47# net47 1.26e-20
C3792 _042_ _152_/a_68_297# 1.02e-20
C3793 cal_itt\[0\] _001_ 0.0135f
C3794 VPWR _336_/a_193_47# 0.0244f
C3795 _304_/a_543_47# cal_count\[3\] 3.03e-21
C3796 _232_/a_32_297# _095_ 4.99e-19
C3797 _328_/a_805_47# _025_ 1.11e-19
C3798 _328_/a_448_47# clknet_2_2__leaf_clk 0.0164f
C3799 _136_ _301_/a_129_47# 4.21e-19
C3800 _216_/a_199_47# _018_ 3.21e-20
C3801 _340_/a_1602_47# _298_/a_215_47# 3.17e-21
C3802 net4 _316_/a_1108_47# 0.00387f
C3803 net9 trim_mask\[4\] 2.61e-20
C3804 _340_/a_27_47# clknet_2_3__leaf_clk 0.0257f
C3805 VPWR ctln[2] 0.00906f
C3806 _341_/a_761_289# _136_ 0.00384f
C3807 _302_/a_373_47# net18 5.13e-19
C3808 net15 net7 0.0193f
C3809 _250_/a_27_297# _249_/a_109_297# 1.58e-19
C3810 net45 _260_/a_93_21# 2.59e-20
C3811 _257_/a_27_297# _336_/a_1108_47# 3.7e-19
C3812 _081_ _006_ 0.0291f
C3813 clkbuf_2_1__f_clk/a_110_47# _246_/a_27_297# 0.0105f
C3814 _325_/a_1283_21# mask\[6\] 0.0692f
C3815 _048_ _192_/a_639_47# 0.0024f
C3816 _077_ rebuffer4/a_27_47# 2.14e-20
C3817 _033_ net18 1.37e-20
C3818 _340_/a_1296_47# _122_ 6.42e-19
C3819 _041_ _338_/a_1032_413# 3.51e-19
C3820 net47 _338_/a_796_47# 0.00142f
C3821 net3 _192_/a_476_47# 9.36e-19
C3822 _314_/a_27_47# _314_/a_193_47# -0.0235f
C3823 _059_ _094_ 0.0451f
C3824 _258_/a_109_297# trim_mask\[2\] 0.00109f
C3825 _306_/a_543_47# rebuffer4/a_27_47# 1.06e-19
C3826 _144_/a_27_47# trimb[4] 4.07e-21
C3827 _255_/a_27_47# clknet_2_2__leaf_clk 4.21e-20
C3828 _103_ _260_/a_93_21# 1.08e-20
C3829 _082_ clknet_2_1__leaf_clk 0.00131f
C3830 _048_ _262_/a_109_297# 0.0145f
C3831 _059_ _088_ 7.29e-21
C3832 _104_ _335_/a_805_47# 1.17e-20
C3833 _050_ _049_ 0.4f
C3834 _326_/a_651_413# output14/a_27_47# 1.35e-20
C3835 net13 _337_/a_761_289# 0.00672f
C3836 _335_/a_543_47# _330_/a_1283_21# 4.14e-19
C3837 net55 net41 9.56e-19
C3838 _110_ _327_/a_761_289# 1.61e-20
C3839 _277_/a_75_212# net50 0.00108f
C3840 _108_ _278_/a_109_297# 1.2e-19
C3841 _250_/a_27_297# mask\[4\] 2.19e-19
C3842 output20/a_27_47# net20 0.043f
C3843 net27 _311_/a_1283_21# 2.42e-19
C3844 _270_/a_59_75# clknet_2_2__leaf_clk 0.0016f
C3845 VPWR _319_/a_1270_413# 4.74e-20
C3846 _329_/a_193_47# _258_/a_27_297# 3.43e-19
C3847 _323_/a_1283_21# net4 5.5e-20
C3848 _078_ _209_/a_27_47# 0.0167f
C3849 _256_/a_27_297# cal_count\[3\] 3.52e-20
C3850 _329_/a_1283_21# trim_mask\[0\] 5.88e-20
C3851 VPWR net55 1.07f
C3852 _323_/a_543_47# net44 0.00197f
C3853 VPWR _223_/a_109_297# 4.7e-20
C3854 _045_ _009_ 0.00719f
C3855 _320_/a_27_47# _041_ 7.84e-19
C3856 trim[4] _332_/a_761_289# 1.68e-19
C3857 _074_ output30/a_27_47# 0.0204f
C3858 _336_/a_193_47# _063_ 1.36e-19
C3859 net47 _339_/a_652_21# 7.51e-19
C3860 _305_/a_27_47# rebuffer5/a_161_47# 5.84e-21
C3861 _257_/a_27_297# _256_/a_27_297# 8.33e-19
C3862 _326_/a_193_47# _314_/a_1108_47# 3.21e-21
C3863 _326_/a_1108_47# _314_/a_193_47# 5.19e-20
C3864 _326_/a_543_47# _314_/a_543_47# 0.00139f
C3865 _340_/a_1602_47# _339_/a_1602_47# 1.04e-20
C3866 _258_/a_27_297# net18 0.00591f
C3867 cal_count\[1\] net33 0.0109f
C3868 _147_/a_27_47# net18 0.00164f
C3869 _024_ net18 0.029f
C3870 _198_/a_181_47# _069_ 2.15e-19
C3871 _189_/a_27_47# _053_ 2.5e-19
C3872 _097_ _241_/a_105_352# 8.1e-19
C3873 _094_ _075_ 1.22e-19
C3874 output8/a_27_47# _175_/a_68_297# 8.9e-21
C3875 trim_mask\[2\] _273_/a_59_75# 0.0537f
C3876 _200_/a_303_47# _092_ 0.00324f
C3877 _247_/a_109_297# mask\[2\] 1.54e-19
C3878 _330_/a_1217_47# net46 5.12e-20
C3879 _308_/a_193_47# _081_ 1.5e-21
C3880 _052_ _062_ 2.54e-20
C3881 _293_/a_384_47# VPWR -4.08e-19
C3882 _122_ _298_/a_78_199# 0.0191f
C3883 net43 _319_/a_1217_47# -1.9e-19
C3884 VPWR _067_ 0.513f
C3885 net51 rebuffer5/a_161_47# 0.0911f
C3886 VPWR _070_ 0.422f
C3887 net3 net45 0.264f
C3888 _326_/a_193_47# _310_/a_193_47# 3.85e-21
C3889 _326_/a_761_289# _310_/a_27_47# 3.13e-20
C3890 net43 _321_/a_761_289# 0.0155f
C3891 VPWR _336_/a_1462_47# 8.89e-19
C3892 _080_ net45 0.00397f
C3893 VPWR _304_/a_805_47# 1.82e-19
C3894 output26/a_27_47# net26 0.0218f
C3895 _037_ _298_/a_78_199# 0.00177f
C3896 ctln[4] net46 1.77e-19
C3897 _334_/a_761_289# net46 0.00139f
C3898 VPWR _340_/a_652_21# 0.0062f
C3899 trim_mask\[2\] clkbuf_2_2__f_clk/a_110_47# 1.07e-19
C3900 net43 _337_/a_761_289# 6.51e-20
C3901 _341_/a_639_47# _038_ 0.00196f
C3902 _021_ _249_/a_27_297# 7.91e-20
C3903 _250_/a_373_47# mask\[5\] 2.82e-19
C3904 _299_/a_27_413# _298_/a_78_199# 4.16e-20
C3905 _025_ _336_/a_1283_21# 6.6e-21
C3906 _336_/a_27_47# clknet_2_2__leaf_clk 0.0181f
C3907 _042_ mask\[5\] 0.00943f
C3908 _117_ _178_/a_68_297# 7.35e-20
C3909 _328_/a_193_47# _327_/a_27_47# 2.52e-20
C3910 _328_/a_27_47# _327_/a_193_47# 2.53e-20
C3911 _319_/a_448_47# _016_ 0.00175f
C3912 _341_/a_1108_47# _122_ 9.16e-20
C3913 output27/a_27_47# net29 5.41e-20
C3914 net27 _224_/a_199_47# 6.1e-21
C3915 _091_ _191_/a_27_297# 1.14e-19
C3916 _325_/a_651_413# _078_ 2.26e-19
C3917 _216_/a_199_47# _078_ 0.00136f
C3918 _270_/a_59_75# trim_val\[0\] 1.89e-21
C3919 _161_/a_68_297# _332_/a_27_47# 5.68e-21
C3920 _099_ net30 7.54e-20
C3921 _327_/a_27_47# net9 5.13e-22
C3922 state\[0\] _232_/a_32_297# 8.12e-19
C3923 _321_/a_193_47# _101_ 0.493f
C3924 _306_/a_27_47# net51 0.00529f
C3925 net3 _065_ 0.0566f
C3926 _015_ _317_/a_1283_21# 9.37e-19
C3927 _338_/a_1032_413# net18 0.00919f
C3928 _341_/a_193_47# _341_/a_543_47# -0.0233f
C3929 _034_ _192_/a_174_21# 6.52e-19
C3930 _063_ net55 5.98e-19
C3931 _263_/a_79_21# _096_ 5.63e-20
C3932 _341_/a_1108_47# _037_ 2.26e-19
C3933 net47 _303_/a_761_289# 0.00453f
C3934 _071_ _190_/a_215_47# 0.00714f
C3935 cal_itt\[1\] _190_/a_655_47# 0.019f
C3936 _336_/a_761_289# net19 6.83e-19
C3937 clkbuf_0_clk/a_110_47# _198_/a_27_47# 0.0095f
C3938 _328_/a_27_47# _058_ 0.00513f
C3939 _335_/a_193_47# _027_ 9.9e-20
C3940 _335_/a_27_47# net46 0.0483f
C3941 net15 _039_ 8.96e-21
C3942 _273_/a_59_75# _115_ 0.0101f
C3943 trimb[1] net34 0.0785f
C3944 _262_/a_109_297# _190_/a_27_47# 8.03e-21
C3945 net27 _250_/a_109_297# 6.97e-20
C3946 net28 _313_/a_1108_47# 0.043f
C3947 _266_/a_68_297# _264_/a_27_297# 7.02e-20
C3948 mask\[0\] _095_ 0.00186f
C3949 _015_ _192_/a_174_21# 1.97e-19
C3950 net50 _336_/a_193_47# 1.03e-20
C3951 cal_itt\[0\] _118_ 0.0023f
C3952 _329_/a_543_47# trim_mask\[2\] 2.01e-19
C3953 _074_ _314_/a_27_47# 0.00141f
C3954 _164_/a_161_47# net55 8.54e-19
C3955 net43 _253_/a_81_21# 0.0109f
C3956 net45 _241_/a_388_297# 0.00113f
C3957 VPWR _321_/a_805_47# 1.18e-19
C3958 _286_/a_76_199# _124_ 0.0223f
C3959 net46 rebuffer1/a_75_212# 3.52e-20
C3960 _102_ net14 1.21e-20
C3961 _067_ _063_ 0.54f
C3962 result[5] clknet_2_1__leaf_clk 0.0773f
C3963 _063_ _070_ 0.0225f
C3964 _053_ _227_/a_109_93# 8.89e-20
C3965 _020_ _009_ 1.89e-20
C3966 calibrate _062_ 3.45e-19
C3967 _110_ _330_/a_27_47# 0.00698f
C3968 _041_ _339_/a_1602_47# 0.0475f
C3969 _333_/a_1108_47# net33 0.00671f
C3970 VPWR _313_/a_448_47# 0.00137f
C3971 net47 _339_/a_1056_47# -7.95e-19
C3972 VPWR _337_/a_805_47# 1.5e-19
C3973 _336_/a_761_289# _107_ 0.00133f
C3974 _309_/a_543_47# mask\[7\] 8.38e-21
C3975 _307_/a_27_47# _307_/a_193_47# -0.1f
C3976 net43 clkbuf_0_clk/a_110_47# 4.46e-19
C3977 mask\[1\] clknet_2_0__leaf_clk 7.16e-19
C3978 clknet_0_clk _098_ 4.99e-20
C3979 _050_ state\[1\] 4.82e-20
C3980 _092_ cal_itt\[3\] 4.32e-20
C3981 _304_/a_27_47# _001_ 0.19f
C3982 _246_/a_27_297# net30 7.56e-21
C3983 _323_/a_27_47# clknet_2_3__leaf_clk 1.16e-20
C3984 _310_/a_193_47# _310_/a_543_47# -0.0129f
C3985 _107_ clone1/a_27_47# 0.00977f
C3986 clknet_2_1__leaf_clk _120_ 8.85e-21
C3987 net34 trimb[4] 0.0785f
C3988 _041_ rebuffer6/a_27_47# 0.0359f
C3989 VPWR _172_/a_150_297# -1.53e-20
C3990 _046_ _313_/a_193_47# 9.45e-19
C3991 _051_ _331_/a_543_47# 0.00194f
C3992 _018_ mask\[2\] 3.7e-19
C3993 _292_/a_215_47# net47 1.11e-19
C3994 state\[2\] _318_/a_543_47# 7.62e-19
C3995 fanout44/a_27_47# net45 0.00723f
C3996 net26 _208_/a_76_199# 1.14e-21
C3997 _293_/a_81_21# _291_/a_35_297# 6.66e-19
C3998 _128_ _340_/a_1602_47# 7.48e-19
C3999 cal_count\[0\] net37 2.9e-19
C4000 _134_ _298_/a_493_297# 8.56e-20
C4001 mask\[7\] net28 0.0586f
C4002 VPWR _284_/a_150_297# -5.76e-19
C4003 _303_/a_761_289# net44 2.45e-19
C4004 _006_ net14 0.0111f
C4005 _306_/a_1283_21# _305_/a_651_413# 8.82e-19
C4006 net9 _178_/a_68_297# 2.97e-19
C4007 _051_ _229_/a_27_297# 6.43e-21
C4008 VPWR _338_/a_27_47# 0.0341f
C4009 _053_ net42 0.0279f
C4010 _341_/a_193_47# clknet_2_3__leaf_clk 0.525f
C4011 _200_/a_80_21# en_co_clk 0.0268f
C4012 _323_/a_27_47# _303_/a_193_47# 9.08e-21
C4013 _323_/a_193_47# _303_/a_27_47# 4.37e-21
C4014 _309_/a_1283_21# _081_ 0.00119f
C4015 _309_/a_761_289# _006_ 6.55e-19
C4016 clknet_2_1__leaf_clk _076_ 0.0855f
C4017 net43 _282_/a_68_297# 6.96e-20
C4018 _069_ net19 2.78e-20
C4019 _316_/a_193_47# valid 8.33e-20
C4020 _316_/a_543_47# net41 0.0356f
C4021 _104_ _049_ 0.307f
C4022 VPWR _340_/a_1056_47# 4.86e-19
C4023 _236_/a_109_297# _096_ 7e-20
C4024 net43 _313_/a_639_47# -7.06e-19
C4025 _064_ net30 0.184f
C4026 _336_/a_448_47# trim_mask\[4\] 0.025f
C4027 VPWR _102_ 0.235f
C4028 _322_/a_27_47# _041_ 7.15e-20
C4029 _306_/a_761_289# clknet_2_1__leaf_clk 1.63e-19
C4030 fanout44/a_27_47# _065_ 0.024f
C4031 _308_/a_193_47# _307_/a_1108_47# 6.41e-22
C4032 _308_/a_543_47# _307_/a_543_47# 8.87e-19
C4033 _308_/a_1108_47# _307_/a_193_47# 5.24e-20
C4034 _269_/a_299_297# _334_/a_193_47# 2.19e-21
C4035 _061_ net37 0.00617f
C4036 mask\[6\] _156_/a_27_47# 7.31e-22
C4037 _187_/a_27_413# _332_/a_1108_47# 0.00112f
C4038 _187_/a_212_413# _332_/a_1283_21# 4.47e-19
C4039 _336_/a_27_47# _279_/a_204_297# 1.34e-19
C4040 _336_/a_193_47# _279_/a_396_47# 0.0116f
C4041 _006_ _040_ 1e-19
C4042 _326_/a_193_47# _224_/a_113_297# 4.52e-20
C4043 _134_ _129_ 0.0296f
C4044 VPWR _316_/a_543_47# 0.0132f
C4045 _332_/a_27_47# _332_/a_1108_47# -2.98e-20
C4046 _332_/a_761_289# _108_ 0.0315f
C4047 _332_/a_193_47# _332_/a_1283_21# -6.53e-19
C4048 net31 rebuffer2/a_75_212# 6.95e-19
C4049 _029_ _332_/a_27_47# 0.152f
C4050 _328_/a_1217_47# _058_ 1e-20
C4051 _335_/a_1217_47# net46 7.02e-19
C4052 _053_ _054_ 0.339f
C4053 _268_/a_75_212# _029_ 0.00964f
C4054 fanout44/a_27_47# _319_/a_27_47# 6.12e-21
C4055 _040_ _121_ 2.96e-20
C4056 clk _331_/a_1270_413# 5.04e-20
C4057 _053_ net30 0.173f
C4058 _001_ _069_ 0.0139f
C4059 _129_ _130_ 0.18f
C4060 ctln[6] _331_/a_1108_47# 3.54e-20
C4061 VPWR _006_ 0.357f
C4062 _251_/a_27_297# net15 0.0133f
C4063 _333_/a_193_47# net32 1.66e-19
C4064 VPWR net17 0.994f
C4065 _324_/a_1270_413# net44 1.27e-19
C4066 _323_/a_27_47# net53 0.00178f
C4067 _089_ clone7/a_27_47# 8.68e-20
C4068 _124_ cal_count\[0\] 0.00903f
C4069 net12 _087_ 0.00185f
C4070 _053_ _168_/a_27_413# 1.27e-19
C4071 net12 _218_/a_113_297# 0.00206f
C4072 VPWR _121_ 0.172f
C4073 _110_ _330_/a_1217_47# 4.53e-19
C4074 _276_/a_59_75# _027_ 1.64e-21
C4075 trim_mask\[2\] _257_/a_109_297# 5.32e-19
C4076 _324_/a_1283_21# _323_/a_543_47# 3.32e-19
C4077 VPWR _010_ 0.0401f
C4078 _256_/a_109_297# trim_mask\[4\] 0.00264f
C4079 net12 _312_/a_27_47# 1.3e-19
C4080 _326_/a_761_289# clknet_2_1__leaf_clk 4.07e-20
C4081 _308_/a_193_47# net14 0.0121f
C4082 _189_/a_408_47# _088_ 6.59e-20
C4083 _113_ rebuffer2/a_75_212# 3.36e-21
C4084 input2/a_27_47# output5/a_27_47# 4.01e-20
C4085 _030_ _108_ 1.99e-20
C4086 VPWR _323_/a_761_289# 0.0108f
C4087 result[0] _307_/a_651_413# 5.48e-19
C4088 net45 _281_/a_103_199# 4.61e-20
C4089 cal _315_/a_448_47# 0.00123f
C4090 _102_ net52 0.0806f
C4091 _322_/a_651_413# net44 2.81e-20
C4092 clknet_2_3__leaf_clk _133_ 0.00197f
C4093 _074_ _310_/a_651_413# 0.00464f
C4094 _314_/a_761_289# net29 0.00218f
C4095 _309_/a_27_47# _308_/a_543_47# 3.47e-19
C4096 _309_/a_193_47# _308_/a_761_289# 2.21e-21
C4097 _110_ ctln[4] 1.91e-19
C4098 _110_ _334_/a_761_289# 6.43e-21
C4099 net21 _313_/a_805_47# 7.65e-20
C4100 _128_ _041_ 0.012f
C4101 _335_/a_193_47# _032_ 0.00635f
C4102 _325_/a_27_47# _321_/a_1108_47# 8.37e-21
C4103 output38/a_27_47# trimb[2] 0.00959f
C4104 net23 _006_ 0.00178f
C4105 _048_ _033_ 3.33e-21
C4106 trim[1] _061_ 6.73e-21
C4107 _226_/a_303_47# _049_ 1.13e-19
C4108 _311_/a_193_47# _311_/a_651_413# -0.00701f
C4109 _306_/a_1108_47# _002_ 8.81e-19
C4110 VPWR _301_/a_285_47# 0.00869f
C4111 _325_/a_193_47# _313_/a_27_47# 7.04e-19
C4112 _187_/a_212_413# _135_ 4.37e-19
C4113 _097_ en_co_clk 0.00288f
C4114 _136_ clknet_2_2__leaf_clk 0.00225f
C4115 output35/a_27_47# _132_ 4.05e-20
C4116 _341_/a_651_413# cal_count\[3\] 0.0265f
C4117 cal_count\[3\] net18 0.423f
C4118 net44 _312_/a_27_47# 0.00291f
C4119 _078_ mask\[2\] 0.116f
C4120 _341_/a_1462_47# clknet_2_3__leaf_clk 0.00219f
C4121 VPWR _341_/a_543_47# 0.0077f
C4122 en_co_clk _192_/a_548_47# 9.46e-20
C4123 _071_ en_co_clk 0.125f
C4124 _051_ net19 7.23e-20
C4125 _339_/a_1032_413# _339_/a_1602_47# -1.42e-32
C4126 net31 _135_ 6.2e-21
C4127 _033_ trim_mask\[4\] 0.0193f
C4128 _276_/a_59_75# _335_/a_448_47# 4.67e-19
C4129 _110_ _335_/a_27_47# 0.0268f
C4130 _305_/a_27_47# net51 0.0281f
C4131 _257_/a_27_297# net18 0.00956f
C4132 _321_/a_193_47# _248_/a_27_297# 1.67e-19
C4133 _005_ _307_/a_27_47# 1.8e-20
C4134 _320_/a_448_47# _040_ 0.0214f
C4135 _053_ _262_/a_465_47# 4.5e-19
C4136 net15 _049_ 0.0163f
C4137 _235_/a_79_21# _049_ 0.00169f
C4138 _030_ _031_ 2.09e-19
C4139 VPWR _308_/a_193_47# 0.0386f
C4140 output22/a_27_47# net43 1.91e-19
C4141 _307_/a_651_413# net14 9.07e-20
C4142 result[7] _085_ 1.61e-21
C4143 _320_/a_1283_21# net53 4.06e-21
C4144 _336_/a_543_47# trim_val\[4\] 1.05e-19
C4145 _336_/a_761_289# _118_ 3.01e-19
C4146 _326_/a_651_413# net29 1.1e-19
C4147 _306_/a_1283_21# _203_/a_59_75# 0.00131f
C4148 _000_ _041_ 0.2f
C4149 _121_ net52 2.08e-20
C4150 trim_mask\[0\] _333_/a_1283_21# 2.4e-20
C4151 net9 net40 0.0692f
C4152 net39 net38 0.067f
C4153 _125_ _132_ 0.00249f
C4154 _088_ _170_/a_81_21# 0.0285f
C4155 _228_/a_79_21# _049_ 0.025f
C4156 net27 _086_ 0.193f
C4157 _321_/a_27_47# mask\[1\] 3.14e-21
C4158 _029_ _332_/a_1217_47# 2.47e-21
C4159 _110_ rebuffer1/a_75_212# 9.81e-20
C4160 _071_ _306_/a_193_47# 6.82e-21
C4161 cal_itt\[2\] _306_/a_1108_47# 1.91e-20
C4162 _036_ net17 0.00164f
C4163 _042_ _310_/a_27_47# 1.81e-20
C4164 VPWR trimb[1] 0.208f
C4165 _074_ _146_/a_68_297# 4.36e-21
C4166 VPWR _320_/a_448_47# 5.38e-19
C4167 _051_ _107_ 0.156f
C4168 _060_ _243_/a_109_47# 0.00527f
C4169 _050_ _337_/a_1108_47# 3.29e-20
C4170 VPWR _339_/a_193_47# 0.0137f
C4171 _191_/a_27_297# clkbuf_2_3__f_clk/a_110_47# 0.00122f
C4172 trim_mask\[1\] _335_/a_1283_21# 1.15e-20
C4173 clknet_2_1__leaf_clk _310_/a_1283_21# 0.0376f
C4174 _167_/a_161_47# _050_ 1.97e-20
C4175 _062_ _203_/a_59_75# 6.02e-20
C4176 _051_ _166_/a_161_47# 0.0551f
C4177 net45 _330_/a_27_47# 7.48e-21
C4178 _333_/a_1462_47# net32 2.91e-19
C4179 _088_ _227_/a_296_53# 1.25e-20
C4180 _052_ _227_/a_209_311# 2.19e-20
C4181 _322_/a_448_47# _320_/a_1283_21# 2.48e-20
C4182 _326_/a_543_47# mask\[6\] 1.16e-21
C4183 fanout44/a_27_47# _337_/a_761_289# 4.89e-20
C4184 cal_itt\[0\] _062_ 0.232f
C4185 net15 _317_/a_805_47# 5.85e-19
C4186 _308_/a_1283_21# net43 0.0163f
C4187 _308_/a_193_47# net23 2.34e-19
C4188 _308_/a_1108_47# _005_ 1.51e-19
C4189 net9 _334_/a_27_47# 0.00213f
C4190 trim_mask\[2\] _025_ 9.3e-20
C4191 ctlp[6] _312_/a_543_47# 9.17e-19
C4192 _258_/a_27_297# trim_mask\[4\] 0.0102f
C4193 trim_val\[1\] rebuffer2/a_75_212# 1.75e-20
C4194 comp _131_ 0.00527f
C4195 _024_ trim_mask\[4\] 4.44e-19
C4196 ctln[6] net11 6.71e-19
C4197 _324_/a_1108_47# clknet_2_3__leaf_clk 2.62e-19
C4198 _112_ _332_/a_193_47# 0.00101f
C4199 trim_mask\[1\] _108_ 0.0105f
C4200 VPWR _307_/a_651_413# 0.00101f
C4201 net45 _120_ 4.53e-21
C4202 net31 _112_ 1.19e-20
C4203 trim[0] trim_mask\[1\] 7.26e-19
C4204 VPWR trimb[4] 0.248f
C4205 _288_/a_145_75# net33 6.02e-19
C4206 _294_/a_68_297# cal_count\[2\] 0.0026f
C4207 net2 _135_ 0.036f
C4208 _329_/a_1270_413# VPWR 1.09e-19
C4209 result[7] _314_/a_543_47# 3.7e-20
C4210 _132_ net40 0.201f
C4211 VPWR clknet_2_3__leaf_clk 1.3f
C4212 _327_/a_27_47# _256_/a_109_297# 3.33e-19
C4213 _327_/a_193_47# _256_/a_27_297# 2.86e-20
C4214 net43 _320_/a_639_47# 5.05e-20
C4215 _263_/a_79_21# _098_ 4.91e-19
C4216 net16 net37 2.55e-20
C4217 en_co_clk cal_count\[2\] 1.66e-19
C4218 _015_ net55 0.00146f
C4219 _321_/a_1283_21# mask\[3\] 5.87e-20
C4220 cal_itt\[0\] _195_/a_76_199# 0.0611f
C4221 cal_itt\[2\] _195_/a_505_21# 3.68e-21
C4222 calibrate _232_/a_32_297# 2.97e-19
C4223 VPWR _153_/a_27_47# 0.0988f
C4224 _130_ _297_/a_47_47# 5.4e-20
C4225 _129_ _297_/a_377_297# 0.00335f
C4226 _329_/a_27_47# _025_ 1.44e-20
C4227 _309_/a_193_47# _309_/a_1108_47# -0.00656f
C4228 net5 comp 6.19e-20
C4229 _128_ _129_ 4.32e-20
C4230 net45 _076_ 1.28e-20
C4231 _064_ _230_/a_59_75# 0.00158f
C4232 _120_ _065_ 0.0481f
C4233 _256_/a_27_297# _058_ 0.0068f
C4234 _305_/a_761_289# clknet_2_1__leaf_clk 3.05e-20
C4235 clknet_0_clk _263_/a_79_21# 4.48e-22
C4236 net14 valid 0.00598f
C4237 _320_/a_448_47# net52 5.81e-19
C4238 _306_/a_1283_21# clknet_2_0__leaf_clk 1.09e-20
C4239 clknet_2_1__leaf_clk _311_/a_448_47# 1.68e-20
C4240 VPWR _303_/a_193_47# 0.0141f
C4241 _078_ _314_/a_193_47# 0.00266f
C4242 _323_/a_543_47# net19 0.00603f
C4243 _060_ _206_/a_27_93# 0.00643f
C4244 _276_/a_59_75# _032_ 0.0323f
C4245 _309_/a_1283_21# _040_ 3.64e-19
C4246 trim_mask\[1\] _031_ 2.04e-20
C4247 _030_ net49 4.69e-20
C4248 _113_ _112_ 0.108f
C4249 _182_/a_27_47# _047_ 4.27e-20
C4250 trim_val\[2\] _334_/a_805_47# 9.25e-20
C4251 VPWR _308_/a_1462_47# 4.04e-19
C4252 output34/a_27_47# _179_/a_27_47# 4.2e-19
C4253 _306_/a_639_47# cal_itt\[3\] 2.69e-19
C4254 _065_ _076_ 0.635f
C4255 _337_/a_448_47# _092_ 0.00126f
C4256 _106_ trim_val\[4\] 0.0101f
C4257 trim_mask\[2\] _333_/a_543_47# 2.97e-20
C4258 calibrate _227_/a_209_311# 2.51e-19
C4259 _036_ _339_/a_193_47# -0.00571f
C4260 _128_ _339_/a_1032_413# 0.0126f
C4261 _319_/a_27_47# _120_ 1.8e-20
C4262 _306_/a_761_289# _065_ 1.3e-21
C4263 _053_ _230_/a_59_75# 0.00252f
C4264 clkbuf_0_clk/a_110_47# _190_/a_465_47# 0.00282f
C4265 _058_ _302_/a_109_47# 6.13e-20
C4266 net41 valid 0.00746f
C4267 VPWR _309_/a_1283_21# 0.0468f
C4268 en_co_clk _243_/a_109_47# 4.69e-20
C4269 _328_/a_543_47# net46 0.00143f
C4270 _326_/a_27_47# _086_ 2.59e-20
C4271 _102_ _216_/a_113_297# 3.99e-20
C4272 _064_ _066_ 6.91e-19
C4273 _093_ _317_/a_193_47# 3.73e-21
C4274 VPWR _339_/a_796_47# 1.16e-19
C4275 VPWR _245_/a_109_297# -0.00187f
C4276 cal_count\[3\] _191_/a_27_297# 0.0689f
C4277 _063_ clknet_2_3__leaf_clk 0.0185f
C4278 ctln[3] net46 4.12e-20
C4279 rebuffer4/a_27_47# _072_ 8.44e-21
C4280 _259_/a_27_297# _033_ 4.61e-19
C4281 output33/a_27_47# _108_ 6.33e-19
C4282 clknet_0_clk clknet_2_2__leaf_clk 0.0807f
C4283 _104_ _336_/a_651_413# 5.97e-19
C4284 _324_/a_1108_47# net53 1.86e-21
C4285 _168_/a_207_413# _052_ 0.00851f
C4286 _185_/a_68_297# _051_ 1.82e-20
C4287 trim[0] output33/a_27_47# 9.86e-19
C4288 output31/a_27_47# trim[2] 0.00245f
C4289 _328_/a_193_47# _271_/a_75_212# 1.96e-19
C4290 trim[1] net16 5.53e-20
C4291 VPWR valid 0.261f
C4292 VPWR net20 0.288f
C4293 net15 state\[1\] 1.16e-19
C4294 _235_/a_79_21# state\[1\] 1.16e-21
C4295 _237_/a_505_21# _090_ 0.0476f
C4296 net13 _322_/a_639_47# 0.00121f
C4297 VPWR net53 0.388f
C4298 _300_/a_129_47# net16 4.35e-20
C4299 VPWR _292_/a_493_297# -3e-19
C4300 _036_ clknet_2_3__leaf_clk 0.0321f
C4301 _280_/a_75_212# _119_ 0.0291f
C4302 output21/a_27_47# _156_/a_27_47# 1.13e-19
C4303 net13 _046_ 7.78e-20
C4304 _322_/a_448_47# _040_ 2.36e-19
C4305 VPWR _324_/a_651_413# 0.00156f
C4306 _048_ clkbuf_2_3__f_clk/a_110_47# 0.00413f
C4307 _322_/a_1283_21# net53 3.23e-20
C4308 _053_ _066_ 0.0457f
C4309 _303_/a_193_47# _063_ 8.5e-21
C4310 net28 _159_/a_27_47# 1.04e-20
C4311 _309_/a_1283_21# net23 0.00142f
C4312 _309_/a_651_413# net43 0.00265f
C4313 _304_/a_543_47# en_co_clk 2.76e-20
C4314 trim[4] clkc 0.0371f
C4315 trim_mask\[0\] trim_val\[4\] 0.0422f
C4316 _258_/a_27_297# _327_/a_27_47# 2.01e-21
C4317 _327_/a_543_47# trim_mask\[0\] 5.05e-19
C4318 _327_/a_27_47# _024_ 0.0798f
C4319 net4 _279_/a_490_47# 0.00201f
C4320 _053_ _304_/a_651_413# 0.00352f
C4321 net23 _245_/a_109_297# 0.00553f
C4322 clk _092_ 0.034f
C4323 _305_/a_1108_47# _002_ 0.0343f
C4324 net16 _332_/a_651_413# 0.00193f
C4325 _255_/a_27_47# _088_ 2.94e-20
C4326 _316_/a_193_47# _095_ 1.18e-19
C4327 _277_/a_75_212# _335_/a_543_47# 6.3e-19
C4328 VPWR _322_/a_448_47# -0.00285f
C4329 net9 _300_/a_285_47# 8.04e-19
C4330 _016_ net14 1.04e-20
C4331 VPWR _331_/a_448_47# 0.00216f
C4332 _314_/a_1283_21# _011_ 4.1e-20
C4333 net12 _099_ 0.00188f
C4334 _092_ clone7/a_27_47# 2.66e-19
C4335 _067_ _193_/a_109_297# 4.22e-21
C4336 _100_ _226_/a_27_47# 1.35e-20
C4337 _051_ _118_ 2.39e-21
C4338 _146_/a_68_297# net26 8.47e-20
C4339 trim_mask\[0\] net35 0.012f
C4340 _104_ _256_/a_109_47# 0.00354f
C4341 _320_/a_1108_47# _209_/a_27_47# 2.12e-19
C4342 _251_/a_109_297# clknet_2_1__leaf_clk 1.3e-19
C4343 _324_/a_27_47# _312_/a_1283_21# 1.2e-19
C4344 _250_/a_373_47# clknet_2_1__leaf_clk 2.72e-19
C4345 en_co_clk _206_/a_27_93# 0.00658f
C4346 VPWR _303_/a_1462_47# 2.56e-19
C4347 _093_ net30 9.79e-21
C4348 trim_val\[1\] _112_ 0.00575f
C4349 trim_mask\[1\] net49 0.0777f
C4350 _042_ clknet_2_1__leaf_clk 0.665f
C4351 _245_/a_373_47# _101_ 8.5e-19
C4352 net2 _203_/a_59_75# 7.02e-22
C4353 _327_/a_448_47# _136_ 5.57e-19
C4354 _261_/a_113_47# net19 1.68e-19
C4355 net15 _319_/a_543_47# 0.00861f
C4356 _328_/a_1283_21# _029_ 5.83e-21
C4357 net4 _092_ 0.0098f
C4358 _086_ _310_/a_761_289# 1.59e-22
C4359 _078_ _244_/a_27_297# 4.42e-20
C4360 cal_itt\[0\] net2 0.00936f
C4361 net27 _313_/a_27_47# 3.51e-20
C4362 VPWR _266_/a_68_297# 0.0237f
C4363 result[4] _253_/a_384_47# 1.3e-20
C4364 cal_itt\[0\] _305_/a_1283_21# 1.59e-20
C4365 cal_itt\[2\] _305_/a_1108_47# 0.00671f
C4366 _071_ _305_/a_193_47# 1.05e-19
C4367 net3 _013_ 1.05e-19
C4368 net16 _269_/a_299_297# 0.00983f
C4369 _237_/a_505_21# _048_ 0.00334f
C4370 _229_/a_27_297# _087_ 0.0076f
C4371 _329_/a_639_47# trim_mask\[3\] 1.18e-19
C4372 _313_/a_27_47# _222_/a_113_297# 2.2e-19
C4373 output32/a_27_47# _188_/a_27_47# 2.58e-19
C4374 VPWR _008_ 0.202f
C4375 net50 clknet_2_3__leaf_clk 3.78e-21
C4376 net43 _322_/a_639_47# 1.83e-20
C4377 output35/a_27_47# net32 0.00105f
C4378 _078_ _310_/a_1270_413# 1.98e-19
C4379 _059_ net55 0.0964f
C4380 _169_/a_109_53# net4 0.0193f
C4381 net43 _046_ 0.0109f
C4382 _074_ _078_ 0.166f
C4383 _303_/a_1108_47# _000_ 5.47e-21
C4384 _128_ _297_/a_47_47# 1.51e-21
C4385 _322_/a_1283_21# _008_ 4.31e-20
C4386 VPWR _016_ 0.393f
C4387 _337_/a_543_47# en_co_clk 0.003f
C4388 clone1/a_27_47# _062_ 1.74e-19
C4389 _303_/a_761_289# net19 0.00894f
C4390 _107_ _261_/a_113_47# 1.17e-19
C4391 _292_/a_215_47# cal_count\[1\] 1.72e-19
C4392 VPWR _263_/a_382_297# -3.35e-19
C4393 VPWR _199_/a_109_297# 5.7e-19
C4394 _188_/a_27_47# _187_/a_212_413# 0.00133f
C4395 clk cal 2.95e-20
C4396 state\[2\] clk 0.0574f
C4397 _092_ _073_ 4.32e-20
C4398 _322_/a_1270_413# _101_ 1.37e-19
C4399 _041_ mask\[4\] 1.8e-20
C4400 state\[2\] clone7/a_27_47# 9.29e-19
C4401 _270_/a_59_75# _108_ 1.9e-19
C4402 _034_ _121_ 0.0156f
C4403 _019_ _040_ 8.42e-20
C4404 _337_/a_761_289# _076_ 1.76e-19
C4405 _048_ cal_count\[3\] 0.00449f
C4406 net44 _246_/a_27_297# 2.21e-20
C4407 ctln[2] _334_/a_1108_47# 1.72e-20
C4408 net8 _334_/a_651_413# 0.00203f
C4409 _325_/a_27_47# net13 0.00283f
C4410 _323_/a_193_47# _044_ 1.39e-21
C4411 VPWR _291_/a_35_297# 0.0126f
C4412 _232_/a_32_297# _192_/a_27_47# 8.26e-19
C4413 state\[2\] net4 0.325f
C4414 _053_ net47 0.0146f
C4415 output32/a_27_47# net33 0.00242f
C4416 _340_/a_1602_47# en_co_clk 5.5e-22
C4417 _068_ _065_ 0.00939f
C4418 net23 _016_ 0.0433f
C4419 _190_/a_27_47# clkbuf_2_3__f_clk/a_110_47# 0.00108f
C4420 _304_/a_543_47# _286_/a_76_199# 3.01e-20
C4421 _251_/a_109_47# mask\[6\] 0.00241f
C4422 trim_mask\[4\] cal_count\[3\] 1.55e-20
C4423 _083_ net53 0.0625f
C4424 _250_/a_109_297# _021_ 1.12e-19
C4425 VPWR _019_ 0.155f
C4426 _266_/a_68_297# _063_ 1.54e-20
C4427 VPWR _028_ 0.127f
C4428 _312_/a_1270_413# net20 4.33e-20
C4429 net55 _075_ 2.15e-19
C4430 _308_/a_761_289# mask\[1\] 5.96e-19
C4431 _074_ _315_/a_639_47# 0.00164f
C4432 calibrate _315_/a_1270_413# 4.47e-19
C4433 _093_ _315_/a_651_413# 8.82e-19
C4434 _012_ _315_/a_1108_47# 1.26e-19
C4435 _336_/a_1283_21# _335_/a_27_47# 6.38e-21
C4436 cal_itt\[0\] _123_ 0.00309f
C4437 _064_ _258_/a_373_47# 6.38e-21
C4438 _104_ _258_/a_109_297# 0.0539f
C4439 _239_/a_277_297# net42 2.29e-19
C4440 _022_ clknet_2_1__leaf_clk 0.144f
C4441 _331_/a_27_47# trim_mask\[4\] 2.44e-19
C4442 _331_/a_1283_21# _028_ 0.00204f
C4443 _331_/a_1108_47# clknet_2_2__leaf_clk 1.1e-19
C4444 _257_/a_27_297# trim_mask\[4\] 0.0106f
C4445 clknet_2_3__leaf_clk _279_/a_396_47# 4.93e-20
C4446 _324_/a_1270_413# net19 3.32e-20
C4447 _187_/a_212_413# net33 0.0027f
C4448 _119_ net19 0.442f
C4449 state\[0\] _316_/a_193_47# 3.53e-19
C4450 _317_/a_193_47# _317_/a_448_47# -0.00482f
C4451 net12 _084_ 0.00227f
C4452 net52 _016_ 0.0267f
C4453 _272_/a_299_297# _114_ 2.49e-19
C4454 _143_/a_68_297# _017_ 3.47e-19
C4455 _309_/a_27_47# _212_/a_113_297# 1.24e-20
C4456 _056_ _108_ 0.00425f
C4457 net24 clkbuf_2_1__f_clk/a_110_47# 0.00181f
C4458 net12 _053_ 0.00965f
C4459 _320_/a_651_413# mask\[1\] 0.0278f
C4460 _305_/a_1270_413# _072_ 5.67e-19
C4461 net31 net33 0.485f
C4462 _336_/a_27_47# _108_ 6.55e-19
C4463 _110_ ctln[3] 1.44e-20
C4464 _094_ _096_ 2.17e-19
C4465 trim_mask\[3\] _119_ 0.0315f
C4466 clkbuf_2_0__f_clk/a_110_47# net45 9.16e-19
C4467 net13 _050_ 0.00894f
C4468 _259_/a_109_297# _329_/a_193_47# 3.97e-19
C4469 net15 _313_/a_193_47# 1.11e-19
C4470 _327_/a_1283_21# _341_/a_1283_21# 1.03e-20
C4471 _235_/a_297_47# _337_/a_543_47# 1.22e-20
C4472 _327_/a_193_47# net18 0.00863f
C4473 _313_/a_543_47# _085_ 1.84e-19
C4474 _052_ _100_ 0.00158f
C4475 mask\[1\] _140_/a_68_297# 0.0335f
C4476 _323_/a_448_47# mask\[4\] 1.8e-19
C4477 _035_ _286_/a_76_199# 1.97e-19
C4478 _069_ _195_/a_76_199# 5.64e-21
C4479 output29/a_27_47# result[7] 0.01f
C4480 _167_/a_161_47# net15 1.04e-19
C4481 _188_/a_27_47# net2 0.00103f
C4482 _171_/a_27_47# _054_ 0.0217f
C4483 _119_ _107_ 0.0048f
C4484 _171_/a_27_47# net30 0.0196f
C4485 net44 _084_ 1.46e-19
C4486 trim[4] _136_ 7.1e-20
C4487 _282_/a_68_297# _120_ 0.0049f
C4488 _074_ _004_ 0.0892f
C4489 _058_ net18 0.0388f
C4490 _328_/a_1108_47# _112_ 1.1e-20
C4491 _328_/a_651_413# trim_mask\[1\] 0.0265f
C4492 _325_/a_27_47# net43 0.0112f
C4493 _312_/a_27_47# net19 6.86e-20
C4494 clkbuf_2_0__f_clk/a_110_47# _065_ 0.0331f
C4495 _259_/a_109_297# net18 5.32e-19
C4496 _336_/a_1270_413# net46 -1.07e-19
C4497 _322_/a_1108_47# _209_/a_27_47# 1.04e-19
C4498 net1 _316_/a_639_47# 7.19e-21
C4499 _195_/a_505_21# _067_ 0.0392f
C4500 _019_ net52 9.79e-21
C4501 _168_/a_27_413# _171_/a_27_47# 0.00107f
C4502 _113_ net33 4.06e-22
C4503 _008_ _083_ 0.0415f
C4504 mask\[4\] net18 0.00596f
C4505 _266_/a_150_297# net19 2.11e-19
C4506 _275_/a_81_21# net19 2.46e-21
C4507 _050_ _331_/a_193_47# 0.00139f
C4508 comp _299_/a_27_413# 4.35e-19
C4509 _107_ _087_ 0.0797f
C4510 _325_/a_1217_47# net13 1.36e-19
C4511 clkbuf_2_0__f_clk/a_110_47# _319_/a_27_47# 4.99e-19
C4512 _326_/a_761_289# _253_/a_81_21# 1.8e-19
C4513 _326_/a_193_47# _253_/a_299_297# 3.25e-19
C4514 _166_/a_161_47# _087_ 1.03e-19
C4515 _047_ _161_/a_68_297# 0.00495f
C4516 _275_/a_299_297# trim_val\[3\] 7.4e-19
C4517 _275_/a_81_21# trim_mask\[3\] 0.00518f
C4518 _341_/a_27_47# _053_ 0.017f
C4519 _104_ clkbuf_2_2__f_clk/a_110_47# 0.0012f
C4520 _314_/a_1108_47# _313_/a_193_47# 7.01e-21
C4521 net14 _095_ 1.78e-20
C4522 net2 net33 0.612f
C4523 VPWR _205_/a_27_47# 0.117f
C4524 _024_ net40 5.23e-20
C4525 result[1] result[2] 0.0367f
C4526 clknet_2_1__leaf_clk _011_ 0.185f
C4527 _328_/a_27_47# _328_/a_761_289# -0.0166f
C4528 _266_/a_150_297# _107_ 1.6e-19
C4529 _237_/a_218_47# _099_ 0.00187f
C4530 _078_ net26 0.062f
C4531 _323_/a_448_47# _020_ 0.00196f
C4532 output23/a_27_47# _004_ 9.22e-20
C4533 _305_/a_193_47# _202_/a_79_21# 2.48e-19
C4534 net43 _050_ 1.75e-20
C4535 _192_/a_548_47# _049_ 4.47e-20
C4536 _328_/a_193_47# net9 0.00793f
C4537 _270_/a_59_75# net49 3.31e-19
C4538 _322_/a_1283_21# _205_/a_27_47# 0.00472f
C4539 _076_ _204_/a_75_212# 7.8e-20
C4540 cal_itt\[1\] net30 0.00168f
C4541 _321_/a_448_47# _310_/a_27_47# 6.41e-22
C4542 _321_/a_193_47# _310_/a_1108_47# 2.49e-20
C4543 _261_/a_113_47# _118_ 1.73e-20
C4544 _178_/a_150_297# net18 3.05e-19
C4545 _331_/a_1217_47# trim_mask\[4\] 2.58e-19
C4546 VPWR _279_/a_314_297# -0.0145f
C4547 _256_/a_373_47# net46 5.19e-20
C4548 trim[0] _173_/a_27_47# 2.73e-19
C4549 output31/a_27_47# net32 0.00155f
C4550 _051_ _062_ 0.0911f
C4551 calibrate _100_ 0.631f
C4552 VPWR _325_/a_1270_413# 9.11e-20
C4553 _317_/a_193_47# _014_ -0.00111f
C4554 _317_/a_761_289# clknet_2_0__leaf_clk 0.0196f
C4555 _317_/a_27_47# net45 0.00289f
C4556 _309_/a_1108_47# mask\[1\] 1.15e-19
C4557 _262_/a_27_47# _049_ 0.00201f
C4558 _263_/a_297_47# _107_ 2.06e-19
C4559 net54 _237_/a_505_21# 1.53e-19
C4560 _095_ net41 4.84e-20
C4561 _322_/a_27_47# mask\[3\] 0.307f
C4562 _248_/a_109_47# net53 0.00321f
C4563 mask\[1\] _245_/a_109_47# 0.00256f
C4564 _327_/a_27_47# _257_/a_27_297# 0.00109f
C4565 _307_/a_193_47# fanout43/a_27_47# 1.71e-21
C4566 _048_ _242_/a_297_47# 1.57e-19
C4567 output37/a_27_47# _125_ 0.0117f
C4568 _325_/a_543_47# _046_ 1.31e-19
C4569 _325_/a_651_413# _159_/a_27_47# 1.26e-19
C4570 _199_/a_193_297# _001_ 4.91e-19
C4571 _324_/a_27_47# mask\[4\] 9.76e-21
C4572 _315_/a_193_47# net30 1.98e-21
C4573 clknet_2_2__leaf_clk net11 3.85e-20
C4574 _094_ _337_/a_639_47# 0.00511f
C4575 _327_/a_1462_47# net18 5.71e-20
C4576 net13 _169_/a_301_53# 2.46e-19
C4577 _333_/a_27_47# _333_/a_543_47# -0.00787f
C4578 mask\[7\] _314_/a_193_47# 5.51e-19
C4579 _035_ cal_count\[0\] 2.29e-19
C4580 _312_/a_27_47# _155_/a_68_297# 2.1e-21
C4581 input2/a_27_47# trimb[4] 0.00219f
C4582 result[3] _216_/a_199_47# 5.04e-20
C4583 VPWR _095_ 0.552f
C4584 trim_mask\[4\] _242_/a_297_47# 4.81e-21
C4585 net12 _306_/a_1270_413# 3.74e-20
C4586 _320_/a_1108_47# _208_/a_505_21# 5.98e-21
C4587 _203_/a_145_75# _072_ 6.42e-19
C4588 _321_/a_27_47# _247_/a_27_297# 0.00133f
C4589 clknet_0_clk mask\[2\] 1.5e-19
C4590 net43 net25 0.26f
C4591 _325_/a_1217_47# net43 -3.08e-19
C4592 _312_/a_1217_47# net19 3.38e-20
C4593 _266_/a_68_297# _279_/a_396_47# 0.00121f
C4594 trim_val\[1\] net33 0.127f
C4595 net52 _205_/a_27_47# 6.74e-22
C4596 _320_/a_761_289# _017_ 7.03e-19
C4597 _320_/a_1108_47# mask\[2\] 5.22e-21
C4598 _272_/a_81_21# _056_ 2.92e-20
C4599 _308_/a_193_47# output30/a_27_47# 1.86e-20
C4600 cal_itt\[1\] _072_ 2.1e-20
C4601 cal_itt\[2\] _255_/a_27_47# 8.54e-20
C4602 mask\[0\] _315_/a_27_47# 1.54e-19
C4603 net22 _315_/a_193_47# 0.00108f
C4604 _253_/a_81_21# _310_/a_1283_21# 6.89e-19
C4605 cal_itt\[0\] _150_/a_27_47# 4.47e-22
C4606 trim_mask\[1\] _336_/a_193_47# 0.00141f
C4607 _090_ _241_/a_105_352# 1.71e-19
C4608 _123_ net33 4.06e-22
C4609 net12 rebuffer4/a_27_47# -2.1e-36
C4610 net2 _069_ 0.0612f
C4611 output35/a_27_47# _130_ 0.00105f
C4612 clknet_2_1__leaf_clk _319_/a_1283_21# 0.0013f
C4613 _187_/a_27_413# trim_mask\[0\] 5.9e-21
C4614 _050_ _260_/a_93_21# 0.0243f
C4615 _318_/a_27_47# state\[1\] 4.72e-21
C4616 _318_/a_543_47# net45 8.06e-20
C4617 net8 _272_/a_299_297# 6.57e-19
C4618 _305_/a_1283_21# _069_ 5.34e-20
C4619 _014_ net30 1.8e-20
C4620 _306_/a_1270_413# net44 9.21e-20
C4621 trim_val\[0\] clknet_2_2__leaf_clk 2.4e-19
C4622 output37/a_27_47# net40 2.1e-20
C4623 _304_/a_27_47# _123_ 1.94e-19
C4624 trim_mask\[0\] _332_/a_27_47# 0.00555f
C4625 wire42/a_75_212# _049_ 0.00225f
C4626 _326_/a_1283_21# _023_ 4.1e-20
C4627 _326_/a_448_47# mask\[7\] 8.14e-20
C4628 _326_/a_1108_47# _102_ 0.00202f
C4629 en_co_clk net18 0.00801f
C4630 _214_/a_113_297# net15 1.13e-20
C4631 trim_mask\[0\] _268_/a_75_212# 6.85e-19
C4632 _294_/a_68_297# _129_ 4.36e-19
C4633 input1/a_75_212# valid 1.27e-19
C4634 _097_ _315_/a_1108_47# 2.42e-20
C4635 _041_ _286_/a_76_199# 0.0591f
C4636 net16 cal_count\[2\] 0.0127f
C4637 _286_/a_76_199# _338_/a_1182_261# 7.41e-21
C4638 _047_ _332_/a_1108_47# 1.66e-19
C4639 _324_/a_27_47# _020_ 6.39e-20
C4640 _324_/a_543_47# mask\[5\] 2.57e-19
C4641 clkbuf_0_clk/a_110_47# _068_ 0.0139f
C4642 en_co_clk _129_ 4.52e-19
C4643 _337_/a_1283_21# net51 9.5e-20
C4644 _305_/a_1108_47# _067_ 7.47e-19
C4645 _305_/a_1108_47# _070_ 0.00102f
C4646 _119_ _118_ 2.59e-19
C4647 _328_/a_1462_47# net9 2.57e-19
C4648 net44 rebuffer4/a_27_47# 0.00187f
C4649 net47 _300_/a_47_47# 1.31e-20
C4650 _125_ _130_ 4.49e-21
C4651 mask\[0\] clknet_2_0__leaf_clk 0.0635f
C4652 net22 _014_ 5.06e-20
C4653 _340_/a_476_47# net2 2.46e-19
C4654 _320_/a_193_47# net15 1.55e-19
C4655 _172_/a_68_297# _108_ 0.0102f
C4656 VPWR _327_/a_651_413# 0.00143f
C4657 clone1/a_27_47# _227_/a_209_311# 0.011f
C4658 net4 net46 0.0243f
C4659 _136_ _332_/a_543_47# 8.86e-19
C4660 _136_ _108_ 0.008f
C4661 _317_/a_1217_47# net45 8.84e-20
C4662 _237_/a_76_199# en_co_clk 4.52e-20
C4663 trim[0] _172_/a_68_297# 5.41e-20
C4664 _074_ _313_/a_1108_47# 6.62e-20
C4665 _232_/a_114_297# net55 0.00257f
C4666 _315_/a_193_47# _315_/a_651_413# -0.00355f
C4667 _284_/a_68_297# _108_ 1.4e-20
C4668 clknet_2_2__leaf_clk _279_/a_204_297# 5.17e-20
C4669 net8 output9/a_27_47# 3.66e-19
C4670 net4 _195_/a_439_47# 4.03e-19
C4671 _064_ _280_/a_75_212# 0.0176f
C4672 trim_mask\[2\] _334_/a_761_289# 1.47e-20
C4673 _232_/a_32_297# _337_/a_27_47# 5.83e-20
C4674 mask\[3\] net21 9.79e-21
C4675 _319_/a_193_47# _049_ 0.00111f
C4676 _110_ _336_/a_1270_413# 1.39e-19
C4677 _324_/a_193_47# net27 2.33e-19
C4678 _134_ net40 1.8e-19
C4679 _125_ _339_/a_1602_47# 1.71e-20
C4680 _164_/a_161_47# _095_ 5.12e-19
C4681 _312_/a_543_47# _045_ 1.35e-19
C4682 net55 _170_/a_81_21# 1.88e-19
C4683 net46 _055_ 0.00649f
C4684 state\[0\] net41 0.272f
C4685 net12 _311_/a_193_47# 1.11e-19
C4686 VPWR output27/a_27_47# 0.101f
C4687 _104_ _331_/a_193_47# 1.36e-22
C4688 _104_ _257_/a_109_297# 0.0259f
C4689 _064_ _257_/a_373_47# 1.56e-20
C4690 _122_ net46 1.07e-20
C4691 _123_ _069_ 5.86e-20
C4692 _130_ net40 0.0102f
C4693 trim_mask\[2\] _335_/a_27_47# 3.11e-19
C4694 _260_/a_250_297# _092_ 4.55e-21
C4695 _050_ net3 0.031f
C4696 _246_/a_109_297# _101_ 0.0195f
C4697 _023_ _310_/a_448_47# 4.05e-19
C4698 _080_ _212_/a_199_47# 2.22e-34
C4699 _037_ net46 1.3e-20
C4700 output6/a_27_47# net6 0.0531f
C4701 mask\[7\] _074_ 0.0747f
C4702 VPWR state\[0\] 0.792f
C4703 _273_/a_145_75# net46 3.61e-19
C4704 trim_mask\[1\] _336_/a_1462_47# 1.97e-21
C4705 _043_ _042_ 0.019f
C4706 net45 _315_/a_448_47# 1.84e-21
C4707 clknet_2_0__leaf_clk _315_/a_1270_413# 1.67e-19
C4708 _014_ _315_/a_651_413# 7.28e-21
C4709 _321_/a_761_289# _042_ 0.00526f
C4710 mask\[5\] _101_ 0.243f
C4711 _189_/a_27_47# trim_mask\[0\] 3.41e-19
C4712 _079_ _315_/a_193_47# 7.45e-20
C4713 _005_ fanout43/a_27_47# 4.32e-19
C4714 net44 _311_/a_193_47# 0.0065f
C4715 _306_/a_27_47# rebuffer6/a_27_47# 2.16e-21
C4716 _053_ _331_/a_543_47# 1.42e-21
C4717 trim_mask\[2\] rebuffer1/a_75_212# 0.053f
C4718 _321_/a_448_47# clknet_2_1__leaf_clk 1.61e-19
C4719 _093_ _316_/a_27_47# 2.78e-20
C4720 calibrate _316_/a_193_47# 4.87e-20
C4721 _336_/a_543_47# net30 3.34e-21
C4722 net47 _285_/a_113_47# 3.32e-19
C4723 trim_mask\[0\] _332_/a_1217_47# 0.00108f
C4724 _339_/a_1602_47# net40 1.88e-20
C4725 VPWR _208_/a_218_374# 3.86e-19
C4726 _340_/a_476_47# _123_ 0.0324f
C4727 VPWR _207_/a_109_297# -0.00199f
C4728 clknet_2_1__leaf_clk _313_/a_761_289# 0.0433f
C4729 _060_ _090_ 0.00512f
C4730 _189_/a_218_47# _051_ 4.44e-34
C4731 _041_ cal_count\[0\] 0.419f
C4732 _088_ _098_ 2.83e-19
C4733 cal_count\[0\] _338_/a_1182_261# 0.00246f
C4734 _286_/a_76_199# net18 0.0103f
C4735 clkbuf_2_0__f_clk/a_110_47# _282_/a_68_297# 0.0126f
C4736 _301_/a_47_47# _300_/a_47_47# 0.0163f
C4737 _006_ _310_/a_651_413# 1.1e-20
C4738 cal_itt\[1\] _230_/a_59_75# 9.72e-19
C4739 _262_/a_205_47# _105_ 1.74e-20
C4740 _106_ _227_/a_109_93# 3.64e-19
C4741 _237_/a_218_374# net15 1.97e-19
C4742 _094_ clknet_0_clk 0.0166f
C4743 _341_/a_27_47# _300_/a_47_47# 1.01e-20
C4744 _192_/a_174_21# _096_ 2.5e-20
C4745 net31 output40/a_27_47# 0.00659f
C4746 _293_/a_299_297# _289_/a_68_297# 0.00117f
C4747 _305_/a_193_47# _041_ 7.19e-21
C4748 _322_/a_1108_47# mask\[2\] 8.23e-21
C4749 _206_/a_27_93# _049_ 0.00282f
C4750 _058_ _333_/a_193_47# 0.00218f
C4751 _107_ _099_ 0.0643f
C4752 clknet_0_clk _088_ 5.9e-20
C4753 _058_ _265_/a_81_21# 0.0124f
C4754 net13 net15 0.00271f
C4755 VPWR _226_/a_27_47# 0.0133f
C4756 net13 _235_/a_79_21# 0.0118f
C4757 cal_count\[3\] net40 0.412f
C4758 _301_/a_285_47# _332_/a_761_289# 8.57e-20
C4759 _143_/a_68_297# clknet_2_1__leaf_clk 4.36e-21
C4760 _327_/a_193_47# trim_mask\[4\] 0.00205f
C4761 _327_/a_448_47# clknet_2_2__leaf_clk 0.00253f
C4762 state\[2\] _260_/a_250_297# 0.00858f
C4763 _102_ _146_/a_68_297# 1.65e-19
C4764 mask\[7\] _146_/a_150_297# 1.25e-20
C4765 _058_ _048_ 2.11e-19
C4766 _319_/a_1462_47# _049_ 9.02e-20
C4767 output39/a_27_47# trimb[3] 0.0122f
C4768 _051_ _232_/a_32_297# 1.22e-21
C4769 _257_/a_27_297# net40 5.9e-22
C4770 _115_ rebuffer1/a_75_212# 9.01e-19
C4771 VPWR _330_/a_1108_47# 0.0309f
C4772 _329_/a_1283_21# net46 0.0721f
C4773 ctlp[7] mask\[6\] 5.34e-19
C4774 cal_itt\[1\] _066_ 9.54e-25
C4775 en_co_clk _297_/a_47_47# 2.85e-20
C4776 net42 _106_ 1.56e-19
C4777 _337_/a_543_47# _049_ 0.0111f
C4778 _259_/a_109_297# trim_mask\[4\] 1.06e-20
C4779 _104_ _025_ 8.86e-19
C4780 _058_ trim_mask\[4\] 0.134f
C4781 _104_ _260_/a_93_21# 0.00152f
C4782 _019_ _141_/a_27_47# 4.93e-20
C4783 _337_/a_193_47# net30 7.21e-20
C4784 ctlp[0] output28/a_27_47# 0.0347f
C4785 output14/a_27_47# result[6] 6.17e-19
C4786 _050_ fanout44/a_27_47# 1.33e-21
C4787 trim_mask\[1\] _172_/a_150_297# 5.26e-20
C4788 net49 _172_/a_68_297# 0.00295f
C4789 _314_/a_761_289# net14 0.00489f
C4790 trim_mask\[0\] _227_/a_109_93# 0.0225f
C4791 _128_ _125_ 8.35e-19
C4792 _341_/a_805_47# net46 6.17e-20
C4793 state\[0\] _164_/a_161_47# 0.0325f
C4794 _322_/a_193_47# net15 1.58e-21
C4795 output5/a_27_47# clkc 0.00267f
C4796 _060_ _048_ 0.392f
C4797 net27 net21 0.448f
C4798 _017_ _101_ 1.05e-22
C4799 mask\[0\] _319_/a_639_47# 0.00449f
C4800 clknet_0_clk _108_ 1.25e-20
C4801 _321_/a_761_289# _022_ 7.48e-20
C4802 net21 _222_/a_113_297# 4.04e-19
C4803 fanout46/a_27_47# clkbuf_2_2__f_clk/a_110_47# 0.0029f
C4804 _319_/a_1283_21# net45 6.73e-19
C4805 _319_/a_448_47# clknet_2_0__leaf_clk 0.0139f
C4806 _307_/a_27_47# _039_ 7.99e-19
C4807 _064_ net19 4.18e-20
C4808 _286_/a_218_47# clknet_2_3__leaf_clk 2.48e-19
C4809 net2 output40/a_27_47# 0.0013f
C4810 _051_ _227_/a_209_311# 0.00186f
C4811 mask\[6\] _313_/a_543_47# 8.25e-21
C4812 _308_/a_27_47# _074_ 0.0183f
C4813 net44 _311_/a_1462_47# -6.57e-19
C4814 _064_ _231_/a_161_47# 7e-19
C4815 state\[1\] _243_/a_109_47# 1.67e-19
C4816 net27 _312_/a_1283_21# 0.0118f
C4817 mask\[0\] _337_/a_27_47# 7.17e-20
C4818 _053_ _260_/a_256_47# 0.00107f
C4819 _338_/a_193_47# _123_ 0.00678f
C4820 _106_ net30 0.084f
C4821 _135_ net34 1.32e-20
C4822 _064_ trim_mask\[3\] 0.254f
C4823 net28 _314_/a_193_47# 0.0133f
C4824 _309_/a_27_47# _310_/a_27_47# 2.63e-19
C4825 en_co_clk _090_ 0.00578f
C4826 net43 net15 0.0355f
C4827 _110_ net4 0.326f
C4828 _023_ net29 1.43e-21
C4829 _340_/a_1602_47# net16 0.00324f
C4830 cal_count\[0\] _338_/a_1296_47# 9.23e-20
C4831 cal_count\[0\] net18 0.00559f
C4832 VPWR _306_/a_651_413# 6.68e-19
C4833 _319_/a_1283_21# _065_ 8.51e-19
C4834 _255_/a_27_47# net55 0.00894f
C4835 trim_mask\[0\] net42 3.74e-20
C4836 _301_/a_377_297# _135_ 0.00351f
C4837 _326_/a_651_413# net14 0.00477f
C4838 _053_ net19 0.0347f
C4839 _064_ _107_ 0.00119f
C4840 _241_/a_297_47# _092_ 0.00534f
C4841 _341_/a_193_47# _135_ 0.00145f
C4842 _341_/a_1283_21# net2 0.00641f
C4843 VPWR _314_/a_761_289# 0.00786f
C4844 cal_count\[0\] _129_ 0.0507f
C4845 _128_ net40 2.4e-21
C4846 _332_/a_761_289# clknet_2_3__leaf_clk 1.75e-20
C4847 _053_ _231_/a_161_47# 8.17e-19
C4848 net1 net3 8.1e-20
C4849 _119_ _062_ 1.74e-19
C4850 net35 _109_ 3.95e-20
C4851 _308_/a_1108_47# _039_ 0.00137f
C4852 _336_/a_27_47# _336_/a_193_47# -0.172f
C4853 net8 net33 1.21e-19
C4854 output23/a_27_47# _308_/a_27_47# 0.0112f
C4855 net12 _239_/a_277_297# 0.00306f
C4856 trim[2] net32 6.26e-20
C4857 mask\[7\] net26 0.0661f
C4858 net9 _340_/a_381_47# 0.003f
C4859 _319_/a_193_47# _319_/a_543_47# -0.0102f
C4860 _185_/a_68_297# _099_ 7.19e-21
C4861 _307_/a_448_47# _074_ 0.00471f
C4862 _059_ _263_/a_382_297# 0.00146f
C4863 _053_ _107_ 0.0484f
C4864 trim_mask\[0\] _054_ 5.81e-20
C4865 _052_ net41 0.00169f
C4866 _279_/a_206_47# _118_ 3.03e-20
C4867 _339_/a_1032_413# cal_count\[0\] 0.0796f
C4868 trim_mask\[0\] net30 0.0433f
C4869 _053_ _001_ 5.28e-19
C4870 trim_mask\[3\] _057_ 0.00156f
C4871 _327_/a_27_47# _327_/a_193_47# -0.0436f
C4872 _050_ _281_/a_103_199# 0.018f
C4873 _053_ _166_/a_161_47# 0.0314f
C4874 net12 mask\[6\] 0.00824f
C4875 _282_/a_150_297# _049_ 2.91e-19
C4876 net25 _082_ 0.302f
C4877 _034_ _095_ 4.95e-20
C4878 clk _317_/a_651_413# 0.00154f
C4879 _317_/a_193_47# _316_/a_1108_47# 9.92e-21
C4880 _317_/a_543_47# _316_/a_543_47# 9.85e-20
C4881 net43 _314_/a_1108_47# 0.00566f
C4882 VPWR _195_/a_535_374# 3.56e-20
C4883 cal_itt\[1\] net47 6.69e-19
C4884 _169_/a_215_311# _185_/a_68_297# 3.85e-19
C4885 _257_/a_109_47# net46 1.94e-21
C4886 _028_ _330_/a_543_47# 1.48e-21
C4887 clknet_2_2__leaf_clk _330_/a_1283_21# 0.00182f
C4888 VPWR _326_/a_651_413# 0.00244f
C4889 _051_ _318_/a_1108_47# 2.53e-19
C4890 _329_/a_651_413# _031_ 1.38e-19
C4891 VPWR _334_/a_651_413# 0.013f
C4892 trim_mask\[0\] _168_/a_27_413# 1.5e-20
C4893 _048_ en_co_clk 0.0131f
C4894 VPWR _052_ 0.0475f
C4895 _290_/a_297_47# net34 1.65e-19
C4896 _064_ _279_/a_27_47# 1.42e-20
C4897 _327_/a_27_47# _058_ 0.033f
C4898 _106_ _262_/a_465_47# 3.9e-19
C4899 _328_/a_193_47# _258_/a_27_297# 8.11e-20
C4900 _328_/a_27_47# _258_/a_109_297# 3.66e-19
C4901 _328_/a_1283_21# trim_mask\[0\] 4.74e-19
C4902 _249_/a_27_297# mask\[4\] 0.00435f
C4903 clkbuf_0_clk/a_110_47# cal_itt\[3\] 0.01f
C4904 _258_/a_27_297# net9 6.46e-19
C4905 net9 _024_ 2.6e-20
C4906 _116_ clkbuf_2_2__f_clk/a_110_47# 3.83e-19
C4907 _305_/a_27_47# rebuffer6/a_27_47# 6.02e-20
C4908 _015_ _095_ 1.44e-20
C4909 _331_/a_1283_21# _052_ 2.16e-19
C4910 net9 _147_/a_27_47# 6.92e-19
C4911 mask\[1\] _246_/a_27_297# 0.00327f
C4912 _325_/a_761_289# net27 3.28e-20
C4913 mask\[3\] mask\[4\] 0.0432f
C4914 net43 _310_/a_193_47# 0.0135f
C4915 _330_/a_448_47# net19 0.00495f
C4916 _168_/a_207_413# _051_ 0.0276f
C4917 mask\[6\] net44 2.19e-21
C4918 _324_/a_27_47# _311_/a_1108_47# 2.8e-21
C4919 _155_/a_68_297# _084_ 8.19e-19
C4920 _324_/a_193_47# _311_/a_1283_21# 4.08e-19
C4921 calibrate net14 0.0958f
C4922 _259_/a_27_297# _058_ 1.34e-20
C4923 _064_ _181_/a_68_297# 0.00196f
C4924 VPWR _335_/a_1108_47# 0.0183f
C4925 _323_/a_193_47# net26 0.00549f
C4926 net28 _314_/a_1462_47# 7.77e-20
C4927 net16 _041_ 0.0106f
C4928 fanout47/a_27_47# _067_ 5.48e-19
C4929 _323_/a_1108_47# _042_ 0.0531f
C4930 net50 _330_/a_1108_47# 1.17e-20
C4931 fanout47/a_27_47# _070_ 1.46e-19
C4932 _309_/a_543_47# _074_ 0.00391f
C4933 VPWR _311_/a_27_47# 0.00882f
C4934 net51 rebuffer6/a_27_47# 3.53e-19
C4935 _101_ _310_/a_27_47# 5.73e-22
C4936 VPWR rebuffer2/a_75_212# 0.0884f
C4937 _239_/a_694_21# _098_ 0.00544f
C4938 VPWR _332_/a_1283_21# 0.0247f
C4939 _337_/a_448_47# _065_ 1.52e-19
C4940 calibrate net41 0.0278f
C4941 _110_ _329_/a_1283_21# 2.51e-19
C4942 VPWR _111_ 0.171f
C4943 net28 _074_ 0.0147f
C4944 trim_mask\[0\] _262_/a_465_47# 4.46e-19
C4945 net12 _318_/a_639_47# 2.31e-19
C4946 _053_ _181_/a_68_297# 5.41e-22
C4947 _290_/a_27_413# trimb[1] 0.00504f
C4948 net9 _338_/a_1032_413# 0.00191f
C4949 fanout45/a_27_47# state\[1\] 0.0119f
C4950 _326_/a_651_413# net52 1.99e-20
C4951 mask\[4\] _220_/a_113_297# 1.03e-20
C4952 clk output6/a_27_47# 0.00421f
C4953 result[1] _308_/a_1108_47# 3.76e-19
C4954 _281_/a_253_297# _092_ 0.00117f
C4955 _281_/a_253_47# _095_ 0.0243f
C4956 _102_ _078_ 0.00123f
C4957 trim[4] trim_val\[0\] 1.61e-19
C4958 _322_/a_27_47# net51 3.21e-20
C4959 _339_/a_652_21# _123_ 0.0317f
C4960 _200_/a_209_297# clkbuf_2_3__f_clk/a_110_47# 2.65e-19
C4961 _249_/a_373_47# mask\[5\] -3e-19
C4962 _249_/a_27_297# _020_ 0.0112f
C4963 VPWR _310_/a_639_47# 7.41e-19
C4964 _340_/a_27_47# _304_/a_27_47# 0.00162f
C4965 VPWR calibrate 4.16f
C4966 _204_/a_75_212# cal_itt\[3\] 5.57e-19
C4967 _003_ _203_/a_145_75# 5.24e-20
C4968 _340_/a_562_413# cal_count\[2\] 6.34e-21
C4969 _275_/a_81_21# _335_/a_761_289# 0.00132f
C4970 _275_/a_299_297# _335_/a_193_47# 6.67e-20
C4971 _050_ _120_ 0.0965f
C4972 _096_ net55 0.0642f
C4973 _235_/a_297_47# _048_ 0.0341f
C4974 _322_/a_1108_47# _074_ 6.87e-19
C4975 _143_/a_68_297# _065_ 8.62e-20
C4976 calibrate _331_/a_1283_21# 1.23e-19
C4977 clk net45 0.323f
C4978 _317_/a_27_47# _013_ 2.38e-19
C4979 clknet_2_0__leaf_clk _316_/a_193_47# 0.0036f
C4980 _014_ _316_/a_27_47# 0.0202f
C4981 net3 net15 0.0611f
C4982 state\[0\] _185_/a_150_297# 0.00186f
C4983 _235_/a_79_21# net3 0.0348f
C4984 cal_itt\[0\] _341_/a_193_47# 0.00165f
C4985 net54 _060_ 0.201f
C4986 input4/a_27_47# ctln[0] 3.49e-19
C4987 net4 output6/a_27_47# 0.0302f
C4988 cal_count\[0\] _297_/a_47_47# 4.49e-21
C4989 _074_ _159_/a_27_47# 1.62e-19
C4990 net45 clone7/a_27_47# 1.48e-20
C4991 _290_/a_27_413# trimb[4] 9.58e-19
C4992 output26/a_27_47# output27/a_27_47# 0.00269f
C4993 _006_ _078_ 3.87e-19
C4994 _064_ _118_ 0.0875f
C4995 _309_/a_27_47# clknet_2_1__leaf_clk 0.03f
C4996 _327_/a_1217_47# _058_ 1.84e-19
C4997 mask\[1\] _208_/a_535_374# 2.87e-20
C4998 net27 _045_ 6.13e-19
C4999 result[3] _074_ 6.03e-19
C5000 net16 _298_/a_493_297# 3.42e-20
C5001 _081_ clknet_2_0__leaf_clk 2.17e-20
C5002 _103_ clk 0.00537f
C5003 _292_/a_215_47# net2 0.0383f
C5004 _334_/a_448_47# clknet_2_2__leaf_clk 5.24e-19
C5005 _304_/a_1108_47# _035_ 3.54e-20
C5006 trim_mask\[4\] _228_/a_297_47# 1.96e-19
C5007 en_co_clk _190_/a_27_47# 1.15e-19
C5008 _052_ _260_/a_346_47# 0.00403f
C5009 net43 _310_/a_1462_47# 0.00125f
C5010 _311_/a_639_47# net53 6.89e-19
C5011 clk _065_ 2.07e-20
C5012 _027_ net19 0.0148f
C5013 net4 net45 0.176f
C5014 VPWR _247_/a_373_47# -7.36e-19
C5015 _078_ _010_ 8.71e-19
C5016 _324_/a_193_47# _250_/a_109_297# 4.14e-19
C5017 clknet_0_clk _192_/a_174_21# 0.013f
C5018 cal_itt\[2\] clknet_0_clk 0.186f
C5019 VPWR _135_ 0.173f
C5020 net24 net44 2.51e-21
C5021 _333_/a_27_47# rebuffer1/a_75_212# 6.92e-21
C5022 output21/a_27_47# ctlp[7] 0.0448f
C5023 VPWR _305_/a_651_413# 0.0015f
C5024 trim_mask\[3\] _027_ 0.0619f
C5025 trim_val\[3\] net46 0.0741f
C5026 VPWR _311_/a_1217_47# 4.26e-20
C5027 _053_ _118_ 1.98e-19
C5028 _015_ state\[0\] 0.268f
C5029 net9 _298_/a_215_47# 2.06e-20
C5030 _324_/a_543_47# clknet_2_1__leaf_clk 8.78e-19
C5031 _329_/a_761_289# net9 0.00805f
C5032 output11/a_27_47# ctln[5] 0.0111f
C5033 _335_/a_1283_21# clknet_2_2__leaf_clk 4.35e-20
C5034 net16 _129_ 0.791f
C5035 net43 _224_/a_113_297# 0.0107f
C5036 net4 _065_ 0.0126f
C5037 _302_/a_27_297# _066_ 0.117f
C5038 net27 mask\[4\] 9.99e-19
C5039 net15 _241_/a_388_297# 0.00192f
C5040 net9 _134_ 8.17e-20
C5041 _304_/a_651_413# _302_/a_27_297# 9.19e-21
C5042 output23/a_27_47# result[3] 0.00101f
C5043 _333_/a_1283_21# net46 -8.84e-19
C5044 _237_/a_76_199# _049_ 2.74e-19
C5045 net4 _105_ 0.00345f
C5046 net9 _341_/a_1270_413# 9.87e-20
C5047 _337_/a_1108_47# _206_/a_27_93# 0.00254f
C5048 _336_/a_448_47# _033_ 0.0023f
C5049 _083_ _311_/a_27_47# 0.0291f
C5050 _303_/a_27_47# net26 6.75e-20
C5051 net27 _220_/a_199_47# 0.00142f
C5052 _059_ _095_ 7.45e-19
C5053 clknet_2_2__leaf_clk _108_ 0.124f
C5054 _332_/a_543_47# clknet_2_2__leaf_clk 0.00121f
C5055 _304_/a_193_47# net47 0.00757f
C5056 _322_/a_1217_47# net51 1.93e-20
C5057 _110_ _257_/a_109_47# 2.49e-21
C5058 _164_/a_161_47# calibrate 0.0444f
C5059 net43 _305_/a_805_47# -0.00125f
C5060 net43 _250_/a_27_297# 4.17e-21
C5061 net16 _339_/a_1032_413# 0.00115f
C5062 net13 _318_/a_27_47# 0.0199f
C5063 _308_/a_193_47# _078_ 0.00934f
C5064 _308_/a_543_47# net22 5.67e-19
C5065 _340_/a_27_47# _340_/a_476_47# -0.0112f
C5066 _340_/a_193_47# _340_/a_652_21# 7.11e-33
C5067 net50 _335_/a_1108_47# 0.0118f
C5068 _170_/a_384_47# net41 4.96e-22
C5069 _122_ _065_ 0.079f
C5070 result[6] net29 5.77e-20
C5071 _262_/a_109_297# clkbuf_2_3__f_clk/a_110_47# 9e-20
C5072 _247_/a_373_47# net52 1.9e-20
C5073 mask\[5\] _156_/a_27_47# 2.11e-21
C5074 VPWR _232_/a_304_297# -0.00104f
C5075 _188_/a_27_47# net34 0.00426f
C5076 _065_ _073_ 3.23e-20
C5077 _186_/a_109_297# _060_ 0.00175f
C5078 _292_/a_215_47# _123_ 0.00424f
C5079 _307_/a_543_47# _315_/a_761_289# 5.13e-21
C5080 _307_/a_27_47# _315_/a_1108_47# 4.72e-21
C5081 net54 en_co_clk 0.012f
C5082 _307_/a_761_289# _315_/a_543_47# 5.13e-21
C5083 _307_/a_1108_47# _315_/a_27_47# 4.72e-21
C5084 _014_ _316_/a_1217_47# 7.1e-20
C5085 net45 _316_/a_805_47# -0.001f
C5086 calibrate _260_/a_346_47# 0.00138f
C5087 VPWR _112_ 0.539f
C5088 VPWR _272_/a_299_297# 0.0626f
C5089 _327_/a_193_47# net40 2.47e-20
C5090 _037_ _065_ 1.04e-20
C5091 _051_ _100_ 0.00624f
C5092 VPWR _290_/a_297_47# -6.35e-19
C5093 net2 _199_/a_193_297# 3.07e-19
C5094 _320_/a_1283_21# clknet_2_0__leaf_clk 2.89e-20
C5095 VPWR _170_/a_384_47# -3.54e-19
C5096 _326_/a_193_47# _007_ 1.42e-19
C5097 net27 _020_ 2.32e-20
C5098 _031_ clknet_2_2__leaf_clk 0.0711f
C5099 _074_ _312_/a_639_47# 5.75e-21
C5100 clknet_2_1__leaf_clk _101_ 1.01f
C5101 mask\[0\] _140_/a_68_297# 0.00105f
C5102 trim_mask\[0\] _066_ 0.0196f
C5103 VPWR _239_/a_27_297# 0.0189f
C5104 _058_ net40 0.00678f
C5105 net28 net26 1.3e-20
C5106 _244_/a_27_297# _209_/a_27_47# 7.42e-20
C5107 _317_/a_1108_47# net41 3.16e-21
C5108 _097_ _237_/a_218_374# 9.3e-19
C5109 net4 _336_/a_1283_21# 5.48e-19
C5110 _130_ _132_ 0.259f
C5111 _075_ _095_ 8.5e-20
C5112 _062_ _099_ 2.25e-21
C5113 _312_/a_27_47# _221_/a_109_297# 5.89e-20
C5114 _324_/a_193_47# _021_ 0.0164f
C5115 _326_/a_193_47# mask\[3\] 2.68e-20
C5116 _326_/a_761_289# net25 1.58e-19
C5117 _320_/a_761_289# _065_ 7.65e-21
C5118 _307_/a_1270_413# mask\[0\] 4.86e-21
C5119 _307_/a_639_47# net22 9.4e-19
C5120 _019_ _247_/a_109_297# 6.51e-21
C5121 _064_ _330_/a_761_289# 1.87e-21
C5122 _104_ _330_/a_27_47# 3.03e-20
C5123 trim_val\[0\] _108_ 0.37f
C5124 trim_val\[0\] _332_/a_543_47# 1.9e-19
C5125 _109_ _332_/a_27_47# 4.37e-19
C5126 mask\[1\] rebuffer4/a_27_47# 2.18e-20
C5127 _307_/a_543_47# net45 6.61e-20
C5128 _307_/a_1108_47# clknet_2_0__leaf_clk 3.1e-19
C5129 ctln[5] _330_/a_193_47# 1.07e-20
C5130 _167_/a_161_47# fanout45/a_27_47# 1.28e-19
C5131 net9 cal_count\[3\] 0.129f
C5132 VPWR _289_/a_150_297# 5.32e-19
C5133 _058_ _267_/a_145_75# 2.95e-19
C5134 _051_ _264_/a_27_297# 1.79e-20
C5135 trim[3] _334_/a_1283_21# 2.13e-19
C5136 VPWR output9/a_27_47# 0.0397f
C5137 _074_ _209_/a_27_47# 0.00126f
C5138 net34 net33 0.433f
C5139 VPWR _317_/a_1108_47# -0.00974f
C5140 result[0] clknet_2_0__leaf_clk 0.152f
C5141 _315_/a_27_47# net14 0.0117f
C5142 _136_ _067_ 8.31e-19
C5143 _093_ _107_ 1.73e-19
C5144 _192_/a_27_47# net41 2.68e-21
C5145 _251_/a_109_297# _046_ 1.51e-19
C5146 _237_/a_76_199# _315_/a_1108_47# 7.92e-21
C5147 net27 _222_/a_199_47# 0.00143f
C5148 net47 _302_/a_27_297# 4.88e-20
C5149 _304_/a_805_47# _136_ 1.62e-19
C5150 _284_/a_68_297# _067_ 4.38e-19
C5151 VPWR _203_/a_59_75# 0.0152f
C5152 _304_/a_761_289# _122_ 0.00631f
C5153 _032_ net19 1.11e-19
C5154 _225_/a_109_297# net14 5.22e-19
C5155 VPWR _192_/a_27_47# 0.0176f
C5156 cal_itt\[0\] VPWR 1.27f
C5157 _341_/a_193_47# _304_/a_27_47# 5.81e-21
C5158 _341_/a_27_47# _304_/a_193_47# 3.33e-21
C5159 _311_/a_1462_47# net19 5.5e-20
C5160 output32/a_27_47# _182_/a_27_47# 0.0126f
C5161 net15 _281_/a_103_199# 0.0132f
C5162 _256_/a_109_297# _024_ 0.00564f
C5163 _340_/a_1182_261# net47 -4.58e-19
C5164 _037_ _304_/a_761_289# 1.29e-19
C5165 net54 _235_/a_297_47# 9.56e-19
C5166 _315_/a_27_47# net41 1.9e-20
C5167 _043_ net4 1.61e-20
C5168 ctln[7] _318_/a_639_47# 6.41e-20
C5169 net13 _318_/a_1217_47# 1.14e-19
C5170 _071_ _198_/a_27_47# 1.22e-20
C5171 _012_ net3 2.04e-20
C5172 _108_ _279_/a_204_297# 0.00144f
C5173 trim_mask\[3\] _032_ 0.00318f
C5174 clknet_2_1__leaf_clk _312_/a_448_47# 4.56e-19
C5175 _262_/a_109_297# cal_count\[3\] 2.87e-19
C5176 _308_/a_1270_413# net45 1.41e-19
C5177 _186_/a_109_297# en_co_clk 9.86e-20
C5178 _294_/a_68_297# _125_ 6.58e-20
C5179 trim_mask\[0\] _047_ 1.32e-19
C5180 _007_ _310_/a_543_47# 4.36e-19
C5181 net16 _297_/a_47_47# 1.68e-20
C5182 _308_/a_193_47# _004_ 1.44e-20
C5183 clknet_2_0__leaf_clk net14 0.527f
C5184 net45 _138_/a_27_47# 0.0027f
C5185 _309_/a_1283_21# _078_ 0.0767f
C5186 _309_/a_1108_47# mask\[0\] 3.55e-19
C5187 VPWR _315_/a_27_47# 0.123f
C5188 _309_/a_193_47# net24 0.551f
C5189 _337_/a_193_47# net44 0.00133f
C5190 cal_itt\[0\] _303_/a_805_47# 8.9e-20
C5191 _309_/a_27_47# net45 2.73e-20
C5192 _336_/a_193_47# clknet_0_clk 7.24e-19
C5193 _336_/a_1108_47# clkbuf_2_2__f_clk/a_110_47# 0.00155f
C5194 mask\[0\] _245_/a_109_47# 6.4e-19
C5195 _078_ _245_/a_109_297# 1.34e-20
C5196 _082_ _310_/a_193_47# 0.00178f
C5197 net25 _310_/a_1283_21# 0.0691f
C5198 net49 clknet_2_2__leaf_clk 3.7e-21
C5199 VPWR _318_/a_1270_413# -7.21e-20
C5200 net46 trim_val\[4\] 0.00792f
C5201 output27/a_27_47# _314_/a_27_47# 3.9e-19
C5202 _327_/a_543_47# net46 0.0027f
C5203 _110_ trim_val\[3\] 0.211f
C5204 _071_ net43 0.00629f
C5205 _064_ _062_ 0.464f
C5206 _035_ _338_/a_1602_47# 6.62e-21
C5207 _078_ net20 1.54e-19
C5208 _258_/a_27_297# _033_ 9.34e-20
C5209 _078_ net53 0.229f
C5210 VPWR _225_/a_109_297# -0.0013f
C5211 fanout47/a_27_47# clknet_2_3__leaf_clk 1.9e-20
C5212 _040_ clknet_2_0__leaf_clk 0.0704f
C5213 clknet_2_0__leaf_clk net41 0.123f
C5214 _128_ net9 0.00665f
C5215 clkbuf_0_clk/a_110_47# clk 0.0082f
C5216 _063_ _203_/a_59_75# 3.84e-19
C5217 _089_ _054_ 6.64e-21
C5218 _090_ _049_ 0.222f
C5219 net35 net46 0.00522f
C5220 _259_/a_373_47# net46 1.02e-19
C5221 _050_ clkbuf_2_0__f_clk/a_110_47# 0.0678f
C5222 net33 _133_ 5.06e-20
C5223 _328_/a_1270_413# VPWR -2.21e-19
C5224 _208_/a_439_47# _076_ 6.37e-19
C5225 _164_/a_161_47# _317_/a_1108_47# 8.6e-20
C5226 _294_/a_68_297# net40 0.0078f
C5227 cal_itt\[0\] _063_ 0.299f
C5228 _059_ _226_/a_27_47# 0.00764f
C5229 _064_ _195_/a_76_199# 1.78e-19
C5230 net55 _098_ 0.0966f
C5231 VPWR clknet_2_0__leaf_clk 4.98f
C5232 _053_ _062_ 0.162f
C5233 _315_/a_1217_47# net14 2.37e-19
C5234 mask\[7\] _313_/a_448_47# 4.96e-21
C5235 _304_/a_27_47# _133_ 0.00172f
C5236 en_co_clk net40 0.084f
C5237 _328_/a_27_47# _025_ 0.256f
C5238 _136_ _284_/a_150_297# 1.5e-19
C5239 _271_/a_75_212# _058_ 0.00186f
C5240 _303_/a_193_47# fanout47/a_27_47# 2.48e-19
C5241 clkbuf_0_clk/a_110_47# net4 0.0159f
C5242 _319_/a_1270_413# clknet_0_clk 9.87e-20
C5243 net12 trim_mask\[0\] 5.52e-21
C5244 _341_/a_27_47# _302_/a_27_297# 4.17e-19
C5245 _242_/a_382_297# _049_ 3.21e-19
C5246 net45 _331_/a_761_289# 0.00291f
C5247 _326_/a_193_47# net27 3.19e-20
C5248 trimb[2] trimb[3] 0.0408f
C5249 _287_/a_75_212# _339_/a_193_47# 4.91e-21
C5250 _185_/a_68_297# _093_ 7.18e-20
C5251 clknet_0_clk net55 0.344f
C5252 _144_/a_27_47# output40/a_27_47# 2.19e-20
C5253 trim_val\[2\] _175_/a_68_297# 0.0438f
C5254 _325_/a_27_47# _042_ 1.4e-19
C5255 _297_/a_377_297# _132_ 0.00119f
C5256 net13 _319_/a_193_47# 1.73e-20
C5257 _112_ _333_/a_448_47# 0.00367f
C5258 trim_mask\[1\] _333_/a_1270_413# 1.17e-20
C5259 net49 _333_/a_651_413# 0.00301f
C5260 _340_/a_1032_413# _122_ 0.0353f
C5261 net47 _338_/a_652_21# 0.0163f
C5262 _304_/a_1108_47# net18 6.42e-19
C5263 clknet_2_3__leaf_clk clkc 1.48e-19
C5264 net15 _120_ 0.0591f
C5265 _235_/a_382_297# en_co_clk 3.21e-19
C5266 _053_ _195_/a_76_199# 0.00262f
C5267 _258_/a_27_297# _024_ 8.17e-20
C5268 _340_/a_1296_47# net47 6.52e-19
C5269 net49 trim_val\[0\] 4.74e-20
C5270 net13 _243_/a_109_47# 0.00167f
C5271 _107_ _171_/a_27_47# 0.00468f
C5272 _325_/a_1283_21# clknet_2_1__leaf_clk 5.54e-20
C5273 _104_ _335_/a_27_47# 1.78e-19
C5274 _327_/a_448_47# _108_ 9.48e-19
C5275 _340_/a_1032_413# _037_ 1.39e-19
C5276 _239_/a_277_297# _107_ 5.69e-19
C5277 net43 result[2] 5.53e-20
C5278 net16 _175_/a_68_297# 0.00422f
C5279 net23 clknet_2_0__leaf_clk 7.41e-19
C5280 VPWR _188_/a_27_47# 0.065f
C5281 _327_/a_1108_47# _111_ 0.00162f
C5282 net16 _333_/a_193_47# 0.0161f
C5283 _008_ _078_ 0.165f
C5284 result[4] _310_/a_543_47# 0.00118f
C5285 mask\[7\] _102_ 0.114f
C5286 _287_/a_75_212# clknet_2_3__leaf_clk 4.39e-22
C5287 clk _204_/a_75_212# 4.17e-19
C5288 net16 _265_/a_81_21# 0.0035f
C5289 mask\[4\] _311_/a_1283_21# 0.0672f
C5290 clknet_0_clk _067_ 0.00189f
C5291 VPWR _315_/a_1217_47# 2.13e-19
C5292 clknet_0_clk _070_ 0.00135f
C5293 _226_/a_27_47# _075_ 0.0121f
C5294 _091_ clkbuf_2_3__f_clk/a_110_47# 0.00418f
C5295 _048_ _049_ 0.509f
C5296 _337_/a_1462_47# net44 2.44e-19
C5297 _313_/a_1108_47# _010_ 3.47e-19
C5298 _291_/a_285_297# _127_ 4.1e-19
C5299 _078_ _016_ 3.68e-20
C5300 _058_ _332_/a_1270_413# 3.02e-20
C5301 _334_/a_1283_21# _057_ 1.12e-19
C5302 _189_/a_27_47# _092_ 0.018f
C5303 calibrate input1/a_75_212# 0.00115f
C5304 _015_ calibrate 0.0209f
C5305 clknet_2_1__leaf_clk _248_/a_27_297# 2.24e-20
C5306 cal_itt\[1\] net19 0.215f
C5307 clknet_2_0__leaf_clk net52 0.139f
C5308 net45 _101_ 0.349f
C5309 cal_itt\[1\] _231_/a_161_47# 3.16e-19
C5310 trim_mask\[0\] _301_/a_47_47# 3.95e-20
C5311 trim_mask\[4\] _049_ 0.16f
C5312 _340_/a_193_47# _339_/a_193_47# 4.41e-21
C5313 _256_/a_109_47# net18 4.58e-20
C5314 clk _316_/a_448_47# 2.08e-19
C5315 _101_ _065_ 0.669f
C5316 _330_/a_761_289# _027_ 0.0431f
C5317 _330_/a_193_47# net46 -0.00287f
C5318 net27 _310_/a_543_47# 1.76e-21
C5319 output14/a_27_47# _314_/a_543_47# 0.00343f
C5320 _293_/a_299_297# trimb[4] 1.92e-19
C5321 VPWR net33 0.731f
C5322 _164_/a_161_47# clknet_2_0__leaf_clk 4.38e-20
C5323 _291_/a_285_297# _126_ 0.00108f
C5324 net43 _319_/a_193_47# -0.00263f
C5325 cal_itt\[1\] _107_ 3.8e-19
C5326 _323_/a_1283_21# net47 0.0156f
C5327 cal_itt\[1\] _001_ 0.00103f
C5328 mask\[7\] _010_ 0.00329f
C5329 _158_/a_68_297# net29 0.00632f
C5330 net47 _298_/a_78_199# 8.16e-19
C5331 VPWR _336_/a_761_289# 0.00658f
C5332 _232_/a_32_297# _099_ 0.0651f
C5333 _328_/a_1217_47# _025_ 2.82e-21
C5334 _019_ _078_ 5.23e-20
C5335 _328_/a_651_413# clknet_2_2__leaf_clk 0.00165f
C5336 VPWR _304_/a_27_47# 0.0869f
C5337 _304_/a_639_47# clknet_2_3__leaf_clk 2.64e-19
C5338 _136_ _301_/a_285_47# 0.00565f
C5339 _038_ _122_ 0.00538f
C5340 mask\[6\] _155_/a_68_297# 0.0356f
C5341 _340_/a_193_47# clknet_2_3__leaf_clk 0.00909f
C5342 _341_/a_543_47# _136_ 0.0067f
C5343 _020_ _311_/a_1283_21# 6.17e-19
C5344 _035_ _339_/a_381_47# 9.09e-21
C5345 VPWR clone1/a_27_47# 0.0322f
C5346 _257_/a_109_297# _336_/a_1108_47# 1.54e-19
C5347 clkbuf_2_1__f_clk/a_110_47# _246_/a_109_297# 2.46e-19
C5348 _325_/a_27_47# _022_ 0.263f
C5349 _325_/a_1108_47# mask\[6\] 0.0407f
C5350 _204_/a_75_212# _073_ 0.0101f
C5351 _319_/a_27_47# _101_ 6.81e-20
C5352 _097_ net3 5.88e-20
C5353 _326_/a_27_47# _326_/a_193_47# -0.0178f
C5354 _169_/a_215_311# _232_/a_32_297# 1.86e-20
C5355 net25 _042_ 7.41e-19
C5356 _041_ _338_/a_1602_47# 2.1e-19
C5357 state\[1\] _090_ 5.04e-20
C5358 _334_/a_27_47# _334_/a_193_47# -0.00453f
C5359 net47 _338_/a_1056_47# 0.00112f
C5360 _303_/a_27_47# _067_ 1.31e-22
C5361 net3 _192_/a_548_47# 0.00123f
C5362 clknet_2_1__leaf_clk _249_/a_373_47# 0.00105f
C5363 fanout43/a_27_47# _039_ 2.5e-19
C5364 _277_/a_75_212# net11 4.84e-20
C5365 _303_/a_27_47# _070_ 8.05e-20
C5366 trim_mask\[2\] net4 9.27e-20
C5367 _048_ _262_/a_193_297# 0.0224f
C5368 _321_/a_27_47# _040_ 1.17e-21
C5369 net13 _337_/a_543_47# 0.014f
C5370 net43 _202_/a_79_21# 0.00122f
C5371 _110_ trim_val\[4\] 0.0123f
C5372 _227_/a_109_93# _092_ 4.21e-21
C5373 _110_ _327_/a_543_47# 1.92e-20
C5374 _074_ mask\[2\] 0.00154f
C5375 _040_ _337_/a_27_47# 4.82e-21
C5376 _108_ _278_/a_27_47# 3.51e-19
C5377 _336_/a_27_47# _266_/a_68_297# 5.87e-21
C5378 _250_/a_109_297# mask\[4\] 3.11e-19
C5379 _091_ cal_count\[3\] 2.04e-19
C5380 VPWR _319_/a_639_47# 2.37e-19
C5381 _061_ output35/a_27_47# 7.29e-19
C5382 VPWR _321_/a_27_47# 0.031f
C5383 _125_ cal_count\[0\] 0.422f
C5384 _330_/a_1283_21# _108_ 4.09e-21
C5385 _283_/a_75_212# _049_ 0.0032f
C5386 _053_ net2 8.1e-20
C5387 _320_/a_193_47# _041_ 0.00174f
C5388 trim[4] _332_/a_543_47# 7.31e-20
C5389 _305_/a_27_47# en_co_clk 3.78e-21
C5390 net47 _339_/a_476_47# 0.00316f
C5391 VPWR _337_/a_27_47# -0.00141f
C5392 _212_/a_113_297# net22 4.11e-19
C5393 _257_/a_27_297# _256_/a_109_297# 8.48e-20
C5394 _322_/a_27_47# _321_/a_1283_21# 1.92e-19
C5395 _323_/a_193_47# _323_/a_761_289# -0.00517f
C5396 VPWR _069_ 0.187f
C5397 net34 output40/a_27_47# 0.0147f
C5398 _258_/a_109_297# net18 0.00283f
C5399 clk _013_ 1.58e-19
C5400 _189_/a_218_47# _053_ 1.22e-19
C5401 _097_ _241_/a_388_297# 0.0012f
C5402 _195_/a_218_47# _062_ 0.00222f
C5403 net42 _092_ 0.0209f
C5404 trim_mask\[2\] _273_/a_145_75# 0.00278f
C5405 _302_/a_373_47# cal_count\[3\] 1.46e-19
C5406 _087_ _100_ 0.0124f
C5407 _247_/a_109_47# mask\[2\] 4.16e-19
C5408 _136_ clknet_2_3__leaf_clk 0.181f
C5409 _171_/a_27_47# _118_ 1.86e-20
C5410 _330_/a_1462_47# net46 4.31e-19
C5411 _308_/a_27_47# _006_ 1.37e-20
C5412 _308_/a_761_289# _081_ 9.1e-22
C5413 _048_ state\[1\] 6.16e-19
C5414 en_co_clk net51 1.77e-19
C5415 output32/a_27_47# _161_/a_68_297# 0.00593f
C5416 _122_ _298_/a_292_297# 4.28e-19
C5417 net43 _319_/a_1462_47# -6.49e-19
C5418 _284_/a_68_297# clknet_2_3__leaf_clk 0.002f
C5419 ctlp[1] _158_/a_68_297# 3.63e-19
C5420 _306_/a_193_47# _305_/a_27_47# 1.92e-19
C5421 _306_/a_27_47# _305_/a_193_47# 1.34e-19
C5422 _326_/a_27_47# _310_/a_543_47# 6.4e-21
C5423 _326_/a_761_289# _310_/a_193_47# 6.88e-21
C5424 _326_/a_543_47# _310_/a_27_47# 9.08e-19
C5425 net43 _321_/a_543_47# 0.0348f
C5426 _078_ _205_/a_27_47# 0.0386f
C5427 output7/a_27_47# net7 0.0154f
C5428 VPWR _304_/a_1217_47# 7.1e-20
C5429 output20/a_27_47# _312_/a_27_47# 4.41e-19
C5430 net12 output13/a_27_47# 0.00349f
C5431 _037_ _298_/a_292_297# 6.13e-19
C5432 _334_/a_543_47# net46 0.0233f
C5433 state\[2\] _227_/a_109_93# 8.42e-20
C5434 cal_count\[0\] net40 0.0315f
C5435 VPWR _340_/a_476_47# 0.0301f
C5436 net43 _337_/a_543_47# 3.35e-20
C5437 _341_/a_805_47# _038_ 7.31e-19
C5438 _059_ calibrate 0.0092f
C5439 _336_/a_27_47# _028_ 1.05e-19
C5440 _025_ _336_/a_1108_47# 6.48e-20
C5441 _336_/a_193_47# clknet_2_2__leaf_clk 0.00505f
C5442 clkbuf_2_1__f_clk/a_110_47# _017_ 0.0101f
C5443 _338_/a_1224_47# _122_ 1.73e-19
C5444 _328_/a_193_47# _327_/a_193_47# 4e-20
C5445 _319_/a_639_47# net52 6.3e-20
C5446 _319_/a_651_413# _016_ 6.95e-19
C5447 _341_/a_1108_47# _301_/a_47_47# 4.46e-20
C5448 _341_/a_448_47# _122_ 3.67e-19
C5449 _221_/a_109_297# _084_ 0.00265f
C5450 _121_ clknet_0_clk 0.0132f
C5451 _092_ net30 0.0074f
C5452 _306_/a_193_47# net51 0.00189f
C5453 _327_/a_193_47# net9 9.64e-20
C5454 _015_ _317_/a_1108_47# 5.52e-19
C5455 _321_/a_27_47# net52 0.0211f
C5456 _321_/a_761_289# _101_ 0.0432f
C5457 _338_/a_1602_47# net18 7.99e-19
C5458 _303_/a_1217_47# _070_ 6.83e-20
C5459 _081_ _140_/a_68_297# 0.0504f
C5460 _034_ _192_/a_27_47# 3.76e-21
C5461 _320_/a_1270_413# net44 -3.58e-20
C5462 net31 _161_/a_68_297# 4.7e-19
C5463 _263_/a_79_21# net55 0.0508f
C5464 net47 _303_/a_543_47# 0.00192f
C5465 _303_/a_27_47# _338_/a_27_47# 1.71e-19
C5466 _071_ _190_/a_465_47# 0.00198f
C5467 _336_/a_543_47# net19 0.00765f
C5468 output18/a_27_47# net18 0.0143f
C5469 _061_ net40 0.0224f
C5470 _335_/a_761_289# _027_ 1.21e-19
C5471 _335_/a_193_47# net46 0.0241f
C5472 clknet_2_1__leaf_clk _156_/a_27_47# 5.37e-20
C5473 _328_/a_193_47# _058_ 0.00399f
C5474 _069_ _063_ 0.0696f
C5475 _053_ _123_ 0.0956f
C5476 net54 _049_ 0.284f
C5477 _060_ _318_/a_193_47# 9.79e-21
C5478 net9 _058_ 0.0376f
C5479 _262_/a_193_297# _190_/a_27_47# 8.1e-21
C5480 net27 _251_/a_27_297# 2.01e-19
C5481 net28 _313_/a_448_47# 0.0249f
C5482 _015_ _192_/a_27_47# 3.58e-20
C5483 _051_ net41 0.116f
C5484 _329_/a_1283_21# trim_mask\[2\] 0.00891f
C5485 _074_ _314_/a_193_47# 0.00484f
C5486 _187_/a_27_413# net46 3.5e-19
C5487 net43 _253_/a_299_297# 6.99e-20
C5488 net45 _241_/a_297_47# 1.02e-19
C5489 VPWR input4/a_27_47# 0.0803f
C5490 VPWR _321_/a_1217_47# 4.26e-20
C5491 net3 _243_/a_109_47# 8.21e-21
C5492 _286_/a_505_21# _124_ 1.38e-20
C5493 _332_/a_27_47# net46 0.0347f
C5494 _023_ net14 0.0179f
C5495 _339_/a_1182_261# _122_ 2.09e-19
C5496 _053_ _227_/a_209_311# 6.7e-20
C5497 _308_/a_27_47# _308_/a_193_47# -0.0426f
C5498 _268_/a_75_212# net46 0.0145f
C5499 _110_ _330_/a_193_47# 0.00736f
C5500 _258_/a_27_297# _257_/a_27_297# 8.59e-20
C5501 _041_ _339_/a_381_47# 0.0194f
C5502 net47 _339_/a_1224_47# -3.85e-19
C5503 VPWR _337_/a_1217_47# 1.14e-19
C5504 calibrate _075_ 1.61e-20
C5505 _025_ _256_/a_27_297# 2.61e-20
C5506 VPWR _313_/a_651_413# 5.62e-19
C5507 _336_/a_543_47# _107_ 0.00213f
C5508 _307_/a_27_47# _307_/a_761_289# -0.00751f
C5509 net13 _041_ 0.0129f
C5510 net24 mask\[1\] 0.00304f
C5511 VPWR _051_ 0.884f
C5512 clkbuf_2_0__f_clk/a_110_47# net15 0.0194f
C5513 _304_/a_193_47# _001_ 0.0178f
C5514 _092_ _072_ 4.89e-20
C5515 input1/a_75_212# _315_/a_27_47# 1.03e-21
C5516 _310_/a_193_47# _310_/a_1283_21# -5.93e-19
C5517 _329_/a_27_47# _329_/a_1283_21# -0.0013f
C5518 state\[2\] _054_ 1.37e-20
C5519 _046_ _313_/a_761_289# 0.00279f
C5520 net21 _313_/a_27_47# 7.59e-19
C5521 _340_/a_1032_413# _297_/a_285_47# 4.99e-20
C5522 state\[2\] _318_/a_1283_21# 0.00403f
C5523 _303_/a_1283_21# net4 0.00105f
C5524 state\[2\] net30 9.58e-20
C5525 _293_/a_299_297# _291_/a_35_297# 6.34e-20
C5526 _036_ _340_/a_476_47# 6.1e-19
C5527 _134_ _298_/a_215_47# 0.00196f
C5528 _301_/a_129_47# clknet_2_3__leaf_clk 0.0029f
C5529 _303_/a_543_47# net44 5.09e-19
C5530 _306_/a_1108_47# _305_/a_651_413# 1.35e-19
C5531 net9 _178_/a_150_297# 6.58e-20
C5532 _167_/a_161_47# _090_ 8.23e-21
C5533 _034_ clknet_2_0__leaf_clk 0.0621f
C5534 _097_ _281_/a_103_199# 3.28e-19
C5535 _326_/a_448_47# _074_ 0.00612f
C5536 mask\[2\] net26 7.52e-20
C5537 VPWR _338_/a_193_47# -0.00666f
C5538 _338_/a_1140_413# clknet_2_3__leaf_clk 9.56e-19
C5539 _341_/a_761_289# clknet_2_3__leaf_clk 0.0701f
C5540 _309_/a_1108_47# _081_ 0.00126f
C5541 _309_/a_543_47# _006_ 4.36e-19
C5542 _200_/a_209_297# en_co_clk 0.0454f
C5543 clknet_2_1__leaf_clk _077_ 2.07e-20
C5544 _323_/a_193_47# _303_/a_193_47# 7.45e-21
C5545 _323_/a_27_47# _303_/a_761_289# 1.76e-20
C5546 _323_/a_761_289# _303_/a_27_47# 9.42e-21
C5547 _316_/a_1283_21# net41 0.0673f
C5548 VPWR _340_/a_1224_47# 9.06e-20
C5549 net43 _313_/a_805_47# -0.00124f
C5550 _339_/a_27_47# _339_/a_193_47# -0.248f
C5551 fanout46/a_27_47# _335_/a_27_47# 7.43e-20
C5552 VPWR _023_ 0.602f
C5553 _322_/a_193_47# _041_ 1.44e-20
C5554 _306_/a_543_47# clknet_2_1__leaf_clk 1.07e-19
C5555 net2 rebuffer4/a_27_47# 0.0326f
C5556 _269_/a_81_21# _334_/a_543_47# 1.89e-20
C5557 net29 _085_ 1.86e-19
C5558 _015_ clknet_2_0__leaf_clk 0.0843f
C5559 _334_/a_448_47# _031_ 1.37e-19
C5560 input1/a_75_212# clknet_2_0__leaf_clk 6.32e-20
C5561 _187_/a_212_413# _332_/a_1108_47# 4.77e-20
C5562 _336_/a_761_289# _279_/a_396_47# 1.09e-19
C5563 _336_/a_193_47# _279_/a_204_297# 7.53e-21
C5564 _134_ _130_ 5.7e-20
C5565 output22/a_27_47# _138_/a_27_47# 1.07e-20
C5566 VPWR _316_/a_1283_21# 0.0296f
C5567 _332_/a_543_47# _108_ 0.042f
C5568 _332_/a_193_47# _332_/a_1108_47# -0.00863f
C5569 _332_/a_27_47# _332_/a_448_47# -0.00297f
C5570 _029_ _332_/a_193_47# 2.73e-19
C5571 clknet_0_clk clknet_2_3__leaf_clk 0.00249f
C5572 trim[0] _108_ 9.39e-20
C5573 _335_/a_1462_47# net46 0.00126f
C5574 _328_/a_1462_47# _058_ 1.06e-19
C5575 _106_ net19 0.159f
C5576 _051_ _063_ 7.4e-20
C5577 _049_ rebuffer5/a_161_47# 4.88e-19
C5578 clk _331_/a_639_47# 0.00121f
C5579 _185_/a_68_297# _243_/a_27_297# 8.18e-19
C5580 net43 _041_ 5.66e-19
C5581 output38/a_27_47# net38 0.0202f
C5582 fanout44/a_27_47# _319_/a_193_47# 1.05e-19
C5583 output14/a_27_47# output29/a_27_47# 0.00355f
C5584 _339_/a_27_47# clknet_2_3__leaf_clk 0.00662f
C5585 net28 _010_ 0.0643f
C5586 _141_/a_27_47# clknet_2_0__leaf_clk 3.11e-19
C5587 net8 trim[3] 2.86e-19
C5588 _251_/a_109_297# net15 0.00109f
C5589 _333_/a_761_289# net32 1.34e-19
C5590 output21/a_27_47# _155_/a_68_297# 0.005f
C5591 net16 _125_ 0.0151f
C5592 _326_/a_27_47# _251_/a_27_297# 5.41e-21
C5593 _042_ net15 0.00595f
C5594 _324_/a_639_47# net44 0.00103f
C5595 _323_/a_193_47# net53 0.00126f
C5596 output36/a_27_47# net36 0.0227f
C5597 _339_/a_1296_47# _122_ 9.69e-20
C5598 _332_/a_1217_47# net46 -3.08e-19
C5599 net12 _089_ 0.0146f
C5600 _048_ _337_/a_1108_47# 2.81e-21
C5601 net15 _317_/a_27_47# 0.0147f
C5602 net12 _218_/a_199_47# 1.39e-19
C5603 _110_ _330_/a_1462_47# 4.63e-19
C5604 _276_/a_59_75# net46 3.42e-21
C5605 net3 _337_/a_543_47# 1.35e-21
C5606 _256_/a_109_47# trim_mask\[4\] 2.05e-19
C5607 net12 _312_/a_193_47# 8.37e-19
C5608 _306_/a_27_47# _049_ 8.61e-19
C5609 _106_ _107_ 0.123f
C5610 _326_/a_543_47# clknet_2_1__leaf_clk 6.62e-19
C5611 _308_/a_761_289# net14 0.0137f
C5612 VPWR output40/a_27_47# 0.141f
C5613 _308_/a_1283_21# _138_/a_27_47# 5.15e-19
C5614 net9 en_co_clk 0.0171f
C5615 VPWR _323_/a_543_47# 0.00119f
C5616 result[0] _307_/a_1270_413# 7.73e-21
C5617 cal _315_/a_651_413# 5.19e-19
C5618 _023_ net52 6.2e-21
C5619 _314_/a_543_47# net29 0.00118f
C5620 _322_/a_1270_413# net44 -1.89e-19
C5621 cal_count\[3\] clkbuf_2_3__f_clk/a_110_47# 0.0047f
C5622 _309_/a_27_47# _308_/a_1283_21# 6.42e-21
C5623 _309_/a_193_47# _308_/a_543_47# 8.5e-21
C5624 _300_/a_47_47# net2 0.0422f
C5625 net54 state\[1\] 0.189f
C5626 _113_ _029_ 5.19e-19
C5627 _110_ _334_/a_543_47# 3.4e-20
C5628 net21 _313_/a_1217_47# 5.32e-20
C5629 _335_/a_761_289# _032_ 2.11e-19
C5630 _128_ _338_/a_1032_413# 2.37e-20
C5631 _325_/a_193_47# _321_/a_1108_47# 3.1e-20
C5632 _305_/a_27_47# _305_/a_193_47# -0.329f
C5633 trim_mask\[0\] net19 0.287f
C5634 _078_ _208_/a_218_374# 4.08e-19
C5635 _134_ cal_count\[3\] 0.0058f
C5636 _311_/a_1283_21# _311_/a_1108_47# 5.68e-32
C5637 _311_/a_27_47# _311_/a_639_47# -0.0015f
C5638 _325_/a_193_47# _313_/a_193_47# 1.55e-20
C5639 _325_/a_27_47# _313_/a_761_289# 4.52e-22
C5640 _061_ _300_/a_285_47# 2.76e-20
C5641 trim_mask\[0\] _231_/a_161_47# 0.0047f
C5642 fanout45/a_27_47# net3 0.0249f
C5643 net44 _312_/a_193_47# 0.00527f
C5644 _341_/a_1270_413# cal_count\[3\] 4.21e-19
C5645 net16 net40 0.129f
C5646 en_co_clk _192_/a_639_47# 1.02e-19
C5647 VPWR _341_/a_1283_21# 0.0149f
C5648 _135_ _332_/a_761_289# 3.35e-21
C5649 trim_mask\[3\] trim_mask\[0\] 3.32e-21
C5650 net2 _029_ 1.01e-24
C5651 _339_/a_193_47# _339_/a_586_47# -7.91e-19
C5652 _303_/a_27_47# clknet_2_3__leaf_clk 0.617f
C5653 _230_/a_59_75# _092_ 0.0421f
C5654 _110_ _335_/a_193_47# 0.0115f
C5655 _116_ _335_/a_27_47# 4.14e-20
C5656 VPWR ctlp[4] 0.172f
C5657 _257_/a_109_297# net18 0.0056f
C5658 _294_/a_68_297# _132_ 0.0139f
C5659 _305_/a_193_47# net51 0.00359f
C5660 _321_/a_193_47# _248_/a_109_297# 2.5e-19
C5661 ctlp[1] _085_ 0.0037f
C5662 _005_ _307_/a_193_47# 4.58e-20
C5663 net43 _307_/a_27_47# 4.95e-19
C5664 trim_val\[2\] _334_/a_27_47# 2.19e-19
C5665 _096_ _095_ 0.0479f
C5666 _100_ _099_ 0.0406f
C5667 output13/a_27_47# ctln[7] 0.034f
C5668 en_co_clk _132_ 1.15e-19
C5669 VPWR _308_/a_761_289# 0.023f
C5670 trim_mask\[0\] _107_ 0.0667f
C5671 _336_/a_543_47# _118_ 0.0115f
C5672 _336_/a_1283_21# trim_val\[4\] 0.00319f
C5673 _106_ _279_/a_27_47# 0.00751f
C5674 output23/a_27_47# _074_ 0.00436f
C5675 trim_mask\[0\] _333_/a_1108_47# 3.4e-19
C5676 _052_ _170_/a_81_21# 0.00584f
C5677 clknet_2_0__leaf_clk output30/a_27_47# 0.0847f
C5678 _088_ _170_/a_299_297# 0.0463f
C5679 _228_/a_382_297# _049_ 2.38e-19
C5680 _321_/a_193_47# mask\[1\] 4.19e-21
C5681 _140_/a_68_297# _040_ 3.34e-19
C5682 _029_ _332_/a_1462_47# 6.53e-22
C5683 _110_ _332_/a_27_47# 0.00426f
C5684 _042_ _310_/a_193_47# 2.53e-20
C5685 _303_/a_27_47# _303_/a_193_47# -0.322f
C5686 _277_/a_75_212# _330_/a_1283_21# 1.37e-19
C5687 _060_ _243_/a_373_47# 0.00382f
C5688 _169_/a_215_311# _100_ 3.01e-21
C5689 VPWR _320_/a_651_413# -0.00822f
C5690 _090_ _240_/a_109_297# 3.4e-19
C5691 VPWR _339_/a_652_21# 0.00337f
C5692 trim_mask\[1\] _335_/a_1108_47# 3.39e-21
C5693 ctlp[6] net21 3.56e-20
C5694 clknet_2_1__leaf_clk _310_/a_1108_47# 0.0679f
C5695 _062_ _203_/a_145_75# 6.54e-20
C5696 net45 _330_/a_193_47# 5.82e-23
C5697 _022_ net15 0.00821f
C5698 _047_ _109_ 6.2e-21
C5699 _322_/a_651_413# _320_/a_1283_21# 2.66e-20
C5700 _066_ _092_ 0.0851f
C5701 _088_ _227_/a_368_53# 5.81e-20
C5702 _326_/a_1283_21# mask\[6\] 2.47e-19
C5703 _300_/a_47_47# _123_ 7.17e-20
C5704 fanout44/a_27_47# _337_/a_543_47# 0.00143f
C5705 VPWR _140_/a_68_297# 0.0459f
C5706 cal_itt\[1\] _062_ 0.262f
C5707 net15 _317_/a_1217_47# 2.97e-20
C5708 _333_/a_27_47# _055_ 3.54e-19
C5709 _292_/a_215_47# _133_ 1.3e-20
C5710 net9 _334_/a_193_47# 0.00121f
C5711 _308_/a_1108_47# net43 0.0274f
C5712 _308_/a_761_289# net23 2.72e-19
C5713 _308_/a_448_47# _005_ 0.0128f
C5714 _258_/a_109_297# trim_mask\[4\] 0.00592f
C5715 trim_mask\[1\] rebuffer2/a_75_212# 1.16e-20
C5716 _337_/a_27_47# _034_ 0.00634f
C5717 net49 _108_ 0.118f
C5718 trim[4] output5/a_27_47# 0.00118f
C5719 _059_ clknet_2_0__leaf_clk 2.05e-19
C5720 VPWR _307_/a_1270_413# -4.49e-20
C5721 trim[0] net49 1.66e-19
C5722 VPWR _261_/a_113_47# -4.57e-20
C5723 _329_/a_639_47# _026_ 7.96e-19
C5724 _329_/a_639_47# VPWR 2.96e-19
C5725 trim_mask\[0\] _279_/a_27_47# 0.028f
C5726 net43 _320_/a_805_47# 7.98e-21
C5727 _321_/a_1108_47# mask\[3\] 1.86e-21
C5728 _321_/a_448_47# net25 8.78e-21
C5729 _313_/a_27_47# _045_ 9.7e-21
C5730 _094_ _192_/a_174_21# 4.06e-19
C5731 cal_itt\[0\] _195_/a_505_21# 0.0676f
C5732 cal_itt\[1\] _195_/a_76_199# 0.0366f
C5733 _308_/a_27_47# _016_ 2.75e-21
C5734 _200_/a_80_21# _068_ 4.85e-19
C5735 _093_ _232_/a_32_297# 0.00394f
C5736 _129_ _297_/a_129_47# 2.57e-19
C5737 _303_/a_27_47# net53 1.37e-21
C5738 _329_/a_193_47# _025_ 9.52e-21
C5739 _309_/a_193_47# _309_/a_448_47# -0.00482f
C5740 net23 _140_/a_68_297# 0.0123f
C5741 net48 net46 9.52e-19
C5742 clknet_0_clk _016_ 7.76e-21
C5743 _309_/a_1283_21# _245_/a_27_297# 1.68e-20
C5744 trim_mask\[0\] _181_/a_68_297# 0.0193f
C5745 _256_/a_109_297# _058_ 0.00327f
C5746 trim_val\[3\] trim_mask\[2\] 3.18e-19
C5747 _305_/a_543_47# clknet_2_1__leaf_clk 6.69e-20
C5748 clk _050_ 0.0344f
C5749 _320_/a_651_413# net52 1.67e-19
C5750 _306_/a_1108_47# clknet_2_0__leaf_clk 6.95e-20
C5751 _306_/a_543_47# net45 1e-21
C5752 calibrate _170_/a_81_21# 0.0066f
C5753 result[6] net14 4.91e-20
C5754 output10/a_27_47# net18 0.00701f
C5755 VPWR _303_/a_761_289# 0.00879f
C5756 _050_ clone7/a_27_47# 5.91e-21
C5757 _078_ _314_/a_761_289# 0.00156f
C5758 _048_ _240_/a_109_297# 3.92e-19
C5759 _323_/a_1283_21# net19 0.00502f
C5760 net8 _057_ 0.159f
C5761 _276_/a_145_75# _032_ 0.00138f
C5762 net46 net30 3.76e-21
C5763 _025_ net18 0.00262f
C5764 _303_/a_1108_47# _198_/a_27_47# 5.29e-21
C5765 _030_ _112_ 0.0213f
C5766 trim_val\[2\] _334_/a_1217_47# 1.34e-19
C5767 clkbuf_2_1__f_clk/a_110_47# clknet_2_1__leaf_clk 0.00895f
C5768 _065_ _077_ 0.173f
C5769 _306_/a_805_47# cal_itt\[3\] 1.57e-19
C5770 _058_ net32 0.00353f
C5771 _106_ _118_ 0.00544f
C5772 _128_ _339_/a_1602_47# 0.00794f
C5773 _036_ _339_/a_652_21# 2.56e-19
C5774 _048_ clkbuf_2_2__f_clk/a_110_47# 3.38e-21
C5775 _028_ _098_ 1.39e-20
C5776 clknet_2_0__leaf_clk _075_ 0.00194f
C5777 _319_/a_193_47# _120_ 1.44e-20
C5778 _329_/a_27_47# trim_val\[3\] 8.78e-20
C5779 _050_ net4 0.773f
C5780 _306_/a_543_47# _065_ 2.85e-21
C5781 _053_ _230_/a_145_75# 4.01e-19
C5782 net16 _334_/a_1217_47# 6.83e-21
C5783 _285_/a_113_47# _123_ 2.29e-19
C5784 clkbuf_0_clk/a_110_47# _190_/a_655_47# 0.00389f
C5785 _058_ _302_/a_373_47# 3.46e-20
C5786 VPWR _309_/a_1108_47# 0.0332f
C5787 _074_ net26 1.16f
C5788 net12 _152_/a_68_297# 4.73e-20
C5789 en_co_clk _243_/a_373_47# 7.94e-20
C5790 _276_/a_59_75# _110_ 0.0527f
C5791 _328_/a_1283_21# net46 0.0688f
C5792 _326_/a_193_47# _086_ 0.00579f
C5793 state\[0\] _096_ 2.01e-19
C5794 VPWR _339_/a_1056_47# 1.63e-19
C5795 _261_/a_113_47# _063_ 5.07e-19
C5796 VPWR _245_/a_109_47# -4.32e-19
C5797 clknet_0_clk _028_ 8.37e-20
C5798 clkbuf_2_2__f_clk/a_110_47# trim_mask\[4\] 2.14e-19
C5799 _104_ _336_/a_1270_413# 3.05e-19
C5800 _060_ _337_/a_1283_21# 3.9e-20
C5801 net54 _337_/a_1108_47# 1.55e-20
C5802 _001_ _298_/a_78_199# 9.76e-20
C5803 _064_ _264_/a_27_297# 3.08e-19
C5804 _168_/a_297_47# _052_ 9.31e-19
C5805 _324_/a_448_47# net53 7.43e-19
C5806 _019_ _320_/a_1108_47# 5.18e-20
C5807 _326_/a_651_413# _078_ 9.07e-20
C5808 ctlp[0] _011_ 4.62e-19
C5809 net47 _092_ 0.0024f
C5810 VPWR result[6] 0.161f
C5811 _305_/a_27_47# _049_ 5.51e-20
C5812 _237_/a_218_374# _090_ 1.53e-19
C5813 net13 _322_/a_805_47# 5.18e-19
C5814 _300_/a_285_47# net16 2.73e-19
C5815 VPWR _292_/a_215_47# 0.00312f
C5816 _247_/a_373_47# _018_ 5.05e-20
C5817 _238_/a_75_212# _074_ 1.47e-21
C5818 VPWR _324_/a_1270_413# 5.39e-20
C5819 _026_ _119_ 2.56e-20
C5820 net44 _152_/a_68_297# 0.00258f
C5821 VPWR _119_ 0.109f
C5822 _322_/a_1108_47# net53 9.34e-20
C5823 _050_ _073_ 3.44e-20
C5824 net13 _090_ 0.0117f
C5825 _303_/a_761_289# _063_ 7.96e-20
C5826 mask\[6\] _247_/a_27_297# 1.11e-20
C5827 _134_ _265_/a_299_297# 7.39e-21
C5828 _309_/a_1270_413# net43 -3.58e-20
C5829 _309_/a_1108_47# net23 0.00161f
C5830 trim_mask\[0\] _118_ 0.202f
C5831 _304_/a_1283_21# en_co_clk 6.54e-20
C5832 _258_/a_27_297# _327_/a_193_47# 7.13e-19
C5833 _258_/a_109_297# _327_/a_27_47# 6.37e-21
C5834 net9 cal_count\[0\] 0.045f
C5835 _327_/a_1283_21# trim_mask\[0\] 0.0329f
C5836 _327_/a_193_47# _024_ 0.0853f
C5837 _087_ net41 1.99e-19
C5838 net51 _049_ 0.00338f
C5839 _071_ _068_ 0.319f
C5840 _305_/a_448_47# _002_ 0.0276f
C5841 net23 _245_/a_109_47# 0.00378f
C5842 net16 _332_/a_1270_413# 1.39e-19
C5843 _316_/a_761_289# _095_ 9.69e-20
C5844 _053_ _340_/a_27_47# 0.00282f
C5845 fanout44/a_27_47# _041_ 4.69e-21
C5846 VPWR _322_/a_651_413# -0.0037f
C5847 _000_ rebuffer6/a_27_47# 2.8e-20
C5848 net12 _092_ 0.00962f
C5849 VPWR _331_/a_651_413# 0.00222f
C5850 _314_/a_1108_47# _011_ 1.26e-19
C5851 clknet_2_2__leaf_clk clknet_2_3__leaf_clk 1.6e-20
C5852 _250_/a_27_297# _042_ 5.22e-20
C5853 _078_ _311_/a_27_47# 2.01e-19
C5854 _208_/a_505_21# _070_ 5.95e-22
C5855 _015_ _051_ 0.0399f
C5856 _076_ _202_/a_79_21# 9.14e-20
C5857 _258_/a_27_297# _058_ 7.2e-19
C5858 _309_/a_651_413# _101_ 1.95e-20
C5859 _104_ _256_/a_373_47# 0.00343f
C5860 _024_ _058_ 0.047f
C5861 _324_/a_193_47# _312_/a_1283_21# 1.08e-19
C5862 _324_/a_27_47# _312_/a_1108_47# 7.23e-19
C5863 VPWR _087_ 0.208f
C5864 VPWR _218_/a_113_297# -0.01f
C5865 en_co_clk _206_/a_206_47# 2.33e-19
C5866 _110_ _227_/a_109_93# 4.49e-21
C5867 trim_mask\[1\] _112_ 0.216f
C5868 _245_/a_109_47# net52 3.87e-21
C5869 _245_/a_27_297# _016_ 0.00193f
C5870 _185_/a_68_297# _316_/a_1108_47# 3.02e-20
C5871 _272_/a_299_297# trim_mask\[1\] 1.52e-20
C5872 VPWR _312_/a_27_47# 0.0156f
C5873 net15 _319_/a_1283_21# 8.76e-19
C5874 _086_ _310_/a_543_47# 2.06e-21
C5875 output31/a_27_47# _176_/a_27_47# 8.27e-21
C5876 _322_/a_1283_21# _218_/a_113_297# 1.4e-19
C5877 cal_itt\[1\] net2 5.03e-19
C5878 trim[3] net34 0.061f
C5879 net44 _092_ 7.09e-20
C5880 net27 _313_/a_193_47# 5.06e-22
C5881 VPWR _266_/a_150_297# -4.13e-19
C5882 input3/a_75_212# net14 0.00162f
C5883 output26/a_27_47# _023_ 0.00178f
C5884 cal_itt\[0\] _305_/a_1108_47# 7.11e-20
C5885 net37 _131_ 0.00604f
C5886 net16 _269_/a_384_47# 4.9e-19
C5887 _237_/a_218_374# _048_ 7.33e-19
C5888 _229_/a_27_297# _089_ 0.0679f
C5889 _067_ _278_/a_27_47# 6.89e-19
C5890 _329_/a_805_47# trim_mask\[3\] 4.63e-20
C5891 cal_count\[0\] _132_ 8.08e-21
C5892 _091_ en_co_clk 0.00219f
C5893 VPWR _275_/a_81_21# 0.00341f
C5894 _182_/a_27_47# net34 3.82e-22
C5895 output29/a_27_47# net29 0.0153f
C5896 _237_/a_76_199# net3 9.98e-19
C5897 calibrate _078_ 2.42e-20
C5898 _303_/a_448_47# _000_ 0.00455f
C5899 net24 _310_/a_448_47# 2.92e-21
C5900 net13 _048_ 0.00631f
C5901 _322_/a_1108_47# _008_ 0.00155f
C5902 _320_/a_193_47# _283_/a_75_212# 5.64e-21
C5903 _059_ _337_/a_27_47# 2.77e-19
C5904 _303_/a_543_47# net19 0.0109f
C5905 _337_/a_1283_21# en_co_clk 0.065f
C5906 _097_ clkbuf_2_0__f_clk/a_110_47# 2.21e-19
C5907 VPWR _263_/a_297_47# -0.00102f
C5908 ctlp[6] _045_ 6.87e-19
C5909 _042_ _009_ 5.83e-21
C5910 VPWR _199_/a_193_297# 1.72e-20
C5911 clk net1 2.9e-20
C5912 cal _316_/a_27_47# 8.2e-19
C5913 net12 mask\[5\] 0.318f
C5914 _270_/a_59_75# rebuffer2/a_75_212# 3.49e-20
C5915 _092_ _003_ 4.53e-21
C5916 en output41/a_27_47# 0.00805f
C5917 _081_ _246_/a_27_297# 2.76e-19
C5918 net5 net37 0.00267f
C5919 state\[2\] net12 0.261f
C5920 mask\[6\] net29 6.37e-19
C5921 _341_/a_27_47# _092_ 0.00324f
C5922 _101_ _046_ 0.00309f
C5923 trim_val\[0\] clknet_2_3__leaf_clk 3.62e-22
C5924 _337_/a_543_47# _076_ 1.22e-19
C5925 _336_/a_27_47# _052_ 3.51e-20
C5926 mask\[7\] output27/a_27_47# 1.11e-19
C5927 _320_/a_193_47# mask\[3\] 9.22e-21
C5928 _110_ net48 0.00265f
C5929 _095_ _098_ 2.5e-20
C5930 result[7] clknet_2_1__leaf_clk 0.00252f
C5931 _104_ clk 0.00692f
C5932 trim_mask\[2\] trim_val\[4\] 0.00455f
C5933 net8 _334_/a_1270_413# 1.46e-19
C5934 VPWR input3/a_75_212# 0.0914f
C5935 _325_/a_193_47# net13 0.00405f
C5936 VPWR _291_/a_117_297# -2.55e-20
C5937 _078_ _247_/a_373_47# 1.2e-20
C5938 clknet_2_1__leaf_clk net30 2.02e-20
C5939 _104_ clone7/a_27_47# 2.64e-21
C5940 net24 _247_/a_27_297# 5.06e-20
C5941 _190_/a_215_47# clkbuf_2_3__f_clk/a_110_47# 3.87e-20
C5942 net44 mask\[5\] 0.0319f
C5943 _251_/a_373_47# mask\[6\] 0.00286f
C5944 _110_ net30 0.214f
C5945 _002_ net26 4.53e-21
C5946 _250_/a_109_47# _021_ 6.05e-20
C5947 _312_/a_639_47# net20 0.00117f
C5948 clknet_0_clk _095_ 0.161f
C5949 _308_/a_543_47# mask\[1\] 1.21e-19
C5950 _012_ _315_/a_448_47# 0.00445f
C5951 calibrate _315_/a_639_47# 2.29e-19
C5952 _074_ _315_/a_805_47# 6.43e-19
C5953 net54 _240_/a_109_297# 1.28e-21
C5954 _336_/a_1108_47# _335_/a_27_47# 1.46e-19
C5955 cal_itt\[1\] _123_ 4.01e-20
C5956 _259_/a_373_47# trim_mask\[2\] 2.72e-20
C5957 _239_/a_474_297# net42 3.84e-19
C5958 _331_/a_1108_47# _028_ 0.00379f
C5959 _331_/a_193_47# trim_mask\[4\] 3.68e-19
C5960 _331_/a_448_47# clknet_2_2__leaf_clk 6.21e-19
C5961 _104_ net4 0.166f
C5962 _257_/a_109_297# trim_mask\[4\] 0.0018f
C5963 _281_/a_253_47# _316_/a_1283_21# 1.96e-20
C5964 _317_/a_193_47# _317_/a_651_413# -0.00701f
C5965 state\[0\] _316_/a_761_289# 2.3e-19
C5966 _309_/a_193_47# _212_/a_113_297# 2.38e-20
C5967 clkbuf_2_1__f_clk/a_110_47# net45 0.158f
C5968 _110_ _328_/a_1283_21# 5.34e-21
C5969 _320_/a_1270_413# mask\[1\] 4.37e-19
C5970 _321_/a_448_47# net15 0.00623f
C5971 _336_/a_193_47# _108_ 3.78e-19
C5972 _094_ net55 0.221f
C5973 net50 _119_ 0.00107f
C5974 _305_/a_543_47# _065_ 3.64e-20
C5975 cal_itt\[2\] _002_ 0.0339f
C5976 output15/a_27_47# result[7] 4.15e-20
C5977 ctlp[1] output29/a_27_47# 1.47e-19
C5978 _327_/a_761_289# net18 7.42e-19
C5979 _189_/a_27_47# _103_ 1.28e-19
C5980 ctln[2] _108_ 1.05e-19
C5981 _088_ net55 0.0428f
C5982 _097_ _317_/a_27_47# 4.22e-21
C5983 _035_ _286_/a_505_21# 2.02e-20
C5984 mask\[1\] _140_/a_150_297# 2.2e-19
C5985 clknet_2_1__leaf_clk _072_ 1.55e-20
C5986 _106_ _062_ 0.0208f
C5987 net12 _208_/a_218_47# 1.76e-19
C5988 _318_/a_193_47# _318_/a_761_289# -0.00517f
C5989 _218_/a_113_297# _083_ 2.39e-19
C5990 clkbuf_2_1__f_clk/a_110_47# _065_ 6.09e-19
C5991 _059_ _337_/a_1217_47# 1.23e-19
C5992 _058_ _134_ 4.45e-19
C5993 _066_ net46 2.54e-19
C5994 _059_ _051_ 0.0305f
C5995 calibrate _004_ 2.09e-19
C5996 _325_/a_193_47# net43 0.0113f
C5997 _336_/a_639_47# net46 -7.75e-19
C5998 _328_/a_1270_413# trim_mask\[1\] 4.1e-19
C5999 _312_/a_193_47# net19 4.79e-20
C6000 _259_/a_109_47# net18 3.1e-19
C6001 _232_/a_32_297# _014_ 1.2e-20
C6002 VPWR _333_/a_639_47# 8.68e-19
C6003 _068_ _202_/a_79_21# 0.00218f
C6004 _030_ net33 1.44e-20
C6005 _309_/a_27_47# net25 2.54e-19
C6006 _050_ _331_/a_761_289# 0.00234f
C6007 _210_/a_113_297# net30 0.0281f
C6008 clkbuf_2_1__f_clk/a_110_47# _319_/a_27_47# 0.0219f
C6009 comp _299_/a_215_297# 3.56e-19
C6010 _107_ _089_ 0.00335f
C6011 _325_/a_27_47# _101_ 0.00168f
C6012 net9 net16 0.00341f
C6013 _324_/a_1283_21# _152_/a_68_297# 0.00189f
C6014 net44 _017_ -2.21e-19
C6015 net13 mask\[3\] 0.109f
C6016 _325_/a_1462_47# net13 4.27e-19
C6017 output16/a_27_47# net16 0.0158f
C6018 clkbuf_2_0__f_clk/a_110_47# _319_/a_193_47# 5.02e-20
C6019 _326_/a_543_47# _253_/a_81_21# 0.00344f
C6020 _275_/a_299_297# trim_mask\[3\] 5.11e-19
C6021 _275_/a_81_21# net50 0.00416f
C6022 _275_/a_384_47# trim_val\[3\] 3.91e-19
C6023 _341_/a_193_47# _053_ 0.0171f
C6024 net34 _057_ 0.00266f
C6025 _048_ _260_/a_93_21# 4.7e-21
C6026 trim_mask\[0\] _062_ 0.245f
C6027 trim[2] trim_val\[2\] 0.00257f
C6028 output17/a_27_47# net17 0.0165f
C6029 clk net15 0.0472f
C6030 _328_/a_193_47# _328_/a_761_289# -0.0157f
C6031 _328_/a_27_47# _328_/a_543_47# -0.00454f
C6032 _153_/a_27_47# _044_ 0.0132f
C6033 _237_/a_439_47# _099_ 0.00174f
C6034 _237_/a_218_47# _092_ 9.49e-19
C6035 _119_ _279_/a_396_47# 0.00329f
C6036 _328_/a_761_289# net9 0.00368f
C6037 _192_/a_639_47# _049_ 2.36e-20
C6038 _304_/a_193_47# net2 1.14e-20
C6039 _270_/a_59_75# _112_ 0.0275f
C6040 _270_/a_145_75# net49 2.9e-19
C6041 _322_/a_1108_47# _205_/a_27_47# 0.00157f
C6042 _041_ _076_ 0.0928f
C6043 net3 _090_ 0.0948f
C6044 VPWR _279_/a_206_47# 4.21e-19
C6045 _331_/a_1462_47# trim_mask\[4\] 0.00102f
C6046 _228_/a_79_21# clone7/a_27_47# 2.84e-20
C6047 clknet_2_2__leaf_clk _028_ 0.00261f
C6048 _025_ trim_mask\[4\] 0.016f
C6049 _051_ _075_ 0.141f
C6050 trim[2] net16 4.03e-19
C6051 trim_mask\[4\] _260_/a_93_21# 0.0707f
C6052 _306_/a_543_47# _204_/a_75_212# 3.36e-19
C6053 calibrate _096_ 0.00876f
C6054 VPWR _325_/a_639_47# 5.51e-19
C6055 _317_/a_761_289# _014_ 6.4e-19
C6056 _317_/a_543_47# clknet_2_0__leaf_clk 0.0306f
C6057 _317_/a_193_47# net45 -3.96e-19
C6058 _103_ _227_/a_109_93# 0.0392f
C6059 _237_/a_76_199# _281_/a_103_199# 4.52e-20
C6060 _067_ _108_ 2.97e-19
C6061 _232_/a_32_297# _243_/a_27_297# 0.0115f
C6062 VPWR trim[3] 0.234f
C6063 net4 net15 0.384f
C6064 _327_/a_193_47# _257_/a_27_297# 2.21e-20
C6065 _135_ clkc 2.25e-19
C6066 _047_ net46 6.63e-19
C6067 _322_/a_193_47# mask\[3\] 0.625f
C6068 _248_/a_373_47# net53 0.00338f
C6069 VPWR _158_/a_68_297# 0.028f
C6070 mask\[1\] _245_/a_373_47# -2.91e-19
C6071 net43 _283_/a_75_212# 0.0336f
C6072 net16 _132_ 4.18e-20
C6073 _189_/a_408_47# clone1/a_27_47# 1.76e-20
C6074 _290_/a_207_413# output36/a_27_47# 2.71e-21
C6075 _058_ cal_count\[3\] 0.00167f
C6076 VPWR _182_/a_27_47# 0.0474f
C6077 _324_/a_193_47# mask\[4\] 1.34e-20
C6078 _094_ _337_/a_805_47# 0.00271f
C6079 net13 _169_/a_373_53# 6.93e-19
C6080 mask\[7\] _314_/a_761_289# 2.25e-19
C6081 net13 net54 0.0449f
C6082 net43 _007_ 2.63e-19
C6083 _312_/a_193_47# _155_/a_68_297# 1.03e-20
C6084 VPWR _099_ 0.0698f
C6085 _169_/a_215_311# net41 3.77e-20
C6086 output25/a_27_47# _082_ 3.65e-19
C6087 _257_/a_27_297# _058_ 3.18e-19
C6088 net12 _306_/a_639_47# 0.00108f
C6089 output32/a_27_47# trim_mask\[0\] 7.18e-21
C6090 _321_/a_193_47# _247_/a_27_297# 1.24e-19
C6091 _321_/a_27_47# _247_/a_109_297# 3.77e-20
C6092 _322_/a_27_47# mask\[4\] 5.48e-19
C6093 _325_/a_1462_47# net43 -9.14e-19
C6094 net43 mask\[3\] 0.0301f
C6095 _312_/a_1462_47# net19 9.63e-20
C6096 _226_/a_27_47# _098_ 1.11e-20
C6097 _103_ net42 0.039f
C6098 _320_/a_543_47# _017_ 4.29e-19
C6099 _320_/a_448_47# mask\[2\] 1.38e-19
C6100 trim_mask\[1\] net33 2.41e-19
C6101 _272_/a_299_297# _056_ 9.9e-20
C6102 _071_ cal_itt\[3\] 1.65e-19
C6103 _078_ _315_/a_27_47# 6.64e-20
C6104 net22 _315_/a_761_289# 9.38e-20
C6105 _253_/a_299_297# _310_/a_1283_21# 2.28e-19
C6106 _253_/a_81_21# _310_/a_1108_47# 4.33e-19
C6107 en_co_clk clkbuf_2_3__f_clk/a_110_47# 6.9e-19
C6108 VPWR _169_/a_215_311# 0.00771f
C6109 trim_mask\[1\] _336_/a_761_289# 4.87e-20
C6110 _090_ _241_/a_388_297# 3.97e-19
C6111 _321_/a_27_47# _146_/a_68_297# 8.23e-19
C6112 _040_ _246_/a_27_297# 0.0849f
C6113 _050_ _260_/a_250_297# 0.00209f
C6114 clknet_0_clk _226_/a_27_47# 5.47e-20
C6115 output8/a_27_47# trim_val\[2\] 1.29e-20
C6116 _318_/a_193_47# state\[1\] 2.44e-21
C6117 _318_/a_1283_21# net45 0.0523f
C6118 net8 _272_/a_384_47# 3.26e-19
C6119 _048_ net3 0.869f
C6120 _305_/a_1108_47# _069_ 3.66e-20
C6121 _134_ en_co_clk 0.0584f
C6122 net25 _101_ 1.56e-20
C6123 net45 net30 0.0259f
C6124 net42 _105_ 7.62e-19
C6125 _304_/a_193_47# _123_ 0.00196f
C6126 trim_mask\[0\] _332_/a_193_47# 0.00645f
C6127 net30 rebuffer3/a_75_212# 2.94e-19
C6128 _273_/a_59_75# _334_/a_27_47# 0.00722f
C6129 _326_/a_1108_47# _023_ 1.26e-19
C6130 _326_/a_448_47# _102_ 3.52e-20
C6131 _294_/a_68_297# _130_ 0.0697f
C6132 net31 trim_mask\[0\] 3.14e-19
C6133 clone1/a_27_47# _170_/a_81_21# 8.07e-20
C6134 net52 _158_/a_68_297# 8.6e-20
C6135 _041_ _286_/a_505_21# 0.0215f
C6136 _286_/a_505_21# _338_/a_1182_261# 6.11e-20
C6137 output8/a_27_47# net16 2.4e-20
C6138 _103_ _054_ 5.3e-21
C6139 _219_/a_109_297# mask\[4\] 4.12e-19
C6140 _324_/a_193_47# _020_ 3.29e-20
C6141 _324_/a_1283_21# mask\[5\] 0.00542f
C6142 VPWR _246_/a_27_297# 0.028f
C6143 en_co_clk _130_ 3.39e-20
C6144 _103_ net30 0.0276f
C6145 _337_/a_1108_47# net51 5.9e-20
C6146 _161_/a_68_297# net34 0.0078f
C6147 net24 mask\[0\] 3.77e-20
C6148 _065_ net30 0.634f
C6149 _078_ clknet_2_0__leaf_clk 0.006f
C6150 net22 net45 0.155f
C6151 _340_/a_1182_261# net2 3.27e-20
C6152 net37 _055_ 0.0027f
C6153 output24/a_27_47# net24 0.0264f
C6154 VPWR _327_/a_1270_413# 8e-20
C6155 _172_/a_150_297# _108_ 5.76e-19
C6156 _079_ _210_/a_113_297# 1.68e-20
C6157 net13 net27 0.074f
C6158 _317_/a_1462_47# net45 5.4e-19
C6159 _317_/a_639_47# state\[1\] 1.48e-19
C6160 _103_ _168_/a_27_413# 3.34e-21
C6161 _237_/a_505_21# en_co_clk 5.93e-19
C6162 cal_itt\[0\] fanout47/a_27_47# 0.00255f
C6163 _136_ _111_ 0.0028f
C6164 _122_ net37 7.04e-21
C6165 _232_/a_220_297# net55 7.38e-19
C6166 _232_/a_304_297# _096_ 3.87e-19
C6167 net21 _045_ 0.00973f
C6168 _105_ net30 0.0135f
C6169 _315_/a_1283_21# _315_/a_1108_47# 5.68e-32
C6170 clknet_2_2__leaf_clk _279_/a_314_297# 6e-20
C6171 net27 output28/a_27_47# 1.41e-19
C6172 _327_/a_27_47# _025_ 5.29e-19
C6173 net19 _152_/a_68_297# 0.00139f
C6174 trim_mask\[2\] _334_/a_543_47# 2.23e-19
C6175 _232_/a_32_297# _337_/a_193_47# 3.63e-22
C6176 trim_mask\[0\] _113_ 3.43e-19
C6177 _319_/a_761_289# _049_ 9.8e-19
C6178 _094_ _121_ 0.0342f
C6179 _064_ _026_ 9.4e-21
C6180 _064_ VPWR 0.483f
C6181 _319_/a_27_47# net30 1.48e-19
C6182 net22 _065_ 8.97e-21
C6183 trim[2] _176_/a_27_47# 8.02e-19
C6184 output33/a_27_47# net33 0.0557f
C6185 _164_/a_161_47# _099_ 6.81e-20
C6186 net23 _246_/a_27_297# 5.34e-20
C6187 _243_/a_373_47# _049_ 1.84e-19
C6188 net43 result[4] 7.88e-19
C6189 _053_ net41 8.1e-20
C6190 _104_ _257_/a_109_47# 5.15e-20
C6191 _147_/a_27_47# cal_count\[0\] 2.04e-19
C6192 _239_/a_694_21# net55 1.38e-19
C6193 net4 _124_ 0.00181f
C6194 _321_/a_27_47# _018_ 0.152f
C6195 _301_/a_47_47# net46 3.11e-20
C6196 _309_/a_1283_21# mask\[2\] 1.21e-20
C6197 ctlp[7] clknet_2_1__leaf_clk 1.53e-19
C6198 trim_mask\[0\] net2 1.07e-20
C6199 _209_/a_27_47# _205_/a_27_47# 0.0152f
C6200 _042_ _035_ 2.32e-20
C6201 _334_/a_1270_413# net34 5.17e-20
C6202 trim_mask\[2\] _335_/a_193_47# 1.44e-20
C6203 _065_ _072_ 0.128f
C6204 _341_/a_27_47# net46 -8.16e-19
C6205 mask\[4\] net21 2.5e-19
C6206 VPWR _084_ 0.235f
C6207 _246_/a_109_47# _101_ 3.78e-19
C6208 _246_/a_27_297# net52 0.0303f
C6209 en_co_clk cal_count\[3\] 0.00244f
C6210 _078_ _315_/a_1217_47# 6.12e-20
C6211 _102_ _074_ 0.415f
C6212 VPWR _053_ 1.91f
C6213 _274_/a_75_212# net46 0.0272f
C6214 _041_ _068_ 0.0507f
C6215 clknet_2_0__leaf_clk _315_/a_639_47# 1.44e-19
C6216 _321_/a_543_47# _042_ 0.0026f
C6217 _000_ mask\[4\] 3.63e-20
C6218 _004_ _315_/a_27_47# 1.61e-20
C6219 _189_/a_218_47# trim_mask\[0\] 8.43e-21
C6220 net43 fanout43/a_27_47# 0.0227f
C6221 net44 _311_/a_761_289# -0.00137f
C6222 _306_/a_193_47# rebuffer6/a_27_47# 3.16e-21
C6223 _194_/a_113_297# net30 7.16e-19
C6224 ctln[4] net18 0.00336f
C6225 mask\[2\] net53 0.0021f
C6226 _107_ _279_/a_490_47# 5.99e-19
C6227 _092_ net19 0.00741f
C6228 _321_/a_651_413# clknet_2_1__leaf_clk 0.0045f
C6229 _093_ _316_/a_193_47# 6.32e-20
C6230 calibrate _316_/a_761_289# 6.54e-20
C6231 trim_mask\[0\] _332_/a_1462_47# 0.00222f
C6232 trim[1] _055_ 0.00585f
C6233 net43 net27 0.021f
C6234 _124_ _122_ 0.00765f
C6235 _231_/a_161_47# _092_ 0.0664f
C6236 VPWR _057_ 1.64f
C6237 fanout46/a_27_47# net4 0.0135f
C6238 _026_ _057_ 0.00227f
C6239 VPWR _208_/a_535_374# -1.35e-19
C6240 _340_/a_1182_261# _123_ 0.0391f
C6241 clkbuf_2_1__f_clk/a_110_47# _282_/a_68_297# 1.45e-21
C6242 _136_ _135_ 0.185f
C6243 _281_/a_103_199# _090_ 0.0158f
C6244 net43 _222_/a_113_297# 1.63e-19
C6245 clknet_2_1__leaf_clk _313_/a_543_47# 0.0347f
C6246 cal_itt\[0\] _287_/a_75_212# 0.00199f
C6247 _189_/a_408_47# _051_ -6.94e-36
C6248 _236_/a_109_297# _095_ 5.38e-19
C6249 cal_count\[0\] _338_/a_1032_413# 0.00601f
C6250 _052_ _098_ 0.141f
C6251 _286_/a_505_21# net18 4.43e-19
C6252 _262_/a_465_47# _105_ 0.00164f
C6253 _002_ _067_ 1.66e-21
C6254 _110_ _047_ 2.45e-20
C6255 _074_ _006_ 0.227f
C6256 _064_ _063_ 0.0396f
C6257 _002_ _070_ 9.91e-19
C6258 _106_ _227_/a_209_311# 5.89e-20
C6259 _341_/a_193_47# _300_/a_47_47# 2.39e-19
C6260 _192_/a_27_47# _096_ 4.47e-19
C6261 cal_itt\[2\] net55 1.23e-20
C6262 _335_/a_27_47# net18 2.82e-20
C6263 net43 rebuffer5/a_161_47# 0.0504f
C6264 _322_/a_448_47# mask\[2\] 0.00264f
C6265 _206_/a_206_47# _049_ 2.08e-19
C6266 _058_ _333_/a_761_289# 6.41e-19
C6267 net34 _332_/a_1108_47# 4.6e-20
C6268 _107_ _092_ 0.0107f
C6269 clknet_0_clk _052_ 1.9e-20
C6270 _058_ _265_/a_299_297# 0.00973f
C6271 fanout45/a_27_47# _317_/a_27_47# 9.76e-20
C6272 VPWR _226_/a_109_47# -3.26e-19
C6273 _074_ _010_ 0.033f
C6274 _079_ net45 0.004f
C6275 _004_ clknet_2_0__leaf_clk 0.107f
C6276 trim_mask\[0\] trim_val\[1\] 8.27e-22
C6277 net47 clknet_2_1__leaf_clk -4.67e-20
C6278 _327_/a_651_413# clknet_2_2__leaf_clk 9.04e-19
C6279 cal_itt\[3\] _202_/a_79_21# 4.21e-22
C6280 _053_ _063_ 0.478f
C6281 cal_count\[2\] _131_ 0.595f
C6282 _212_/a_113_297# mask\[1\] 0.00523f
C6283 _329_/a_448_47# _027_ 2e-20
C6284 _329_/a_1108_47# net46 0.0296f
C6285 net43 _306_/a_27_47# 1.21e-19
C6286 VPWR _330_/a_448_47# 0.00283f
C6287 cal_itt\[2\] _067_ 3.46e-19
C6288 cal_itt\[2\] _070_ 0.0638f
C6289 mask\[5\] net19 0.033f
C6290 _337_/a_1283_21# _049_ 0.0176f
C6291 _259_/a_109_47# trim_mask\[4\] 7.59e-20
C6292 _104_ _260_/a_250_297# 6.25e-20
C6293 VPWR _085_ 0.167f
C6294 net49 _172_/a_150_297# 3.05e-19
C6295 _314_/a_543_47# net14 0.00272f
C6296 trim_mask\[0\] _227_/a_209_311# 0.0374f
C6297 net12 clknet_2_1__leaf_clk 1.46f
C6298 _048_ _281_/a_103_199# 0.017f
C6299 _341_/a_1217_47# net46 -1.9e-19
C6300 net16 net32 1.21e-20
C6301 mask\[2\] _016_ 2.53e-20
C6302 mask\[0\] _319_/a_805_47# 0.00218f
C6303 _321_/a_543_47# _022_ 8.25e-19
C6304 net54 net3 0.195f
C6305 _321_/a_27_47# _078_ 6.69e-19
C6306 _319_/a_1108_47# net45 0.00151f
C6307 _319_/a_651_413# clknet_2_0__leaf_clk 0.00604f
C6308 calibrate _098_ 0.247f
C6309 _307_/a_193_47# _039_ 0.00143f
C6310 _286_/a_439_47# clknet_2_3__leaf_clk 3.34e-19
C6311 _051_ _227_/a_296_53# 1.93e-20
C6312 _305_/a_639_47# net44 7.55e-19
C6313 mask\[6\] _313_/a_1283_21# 1.6e-20
C6314 _308_/a_193_47# _074_ 0.028f
C6315 ctln[5] net19 0.00146f
C6316 mask\[0\] _337_/a_193_47# 5.23e-20
C6317 clknet_2_0__leaf_clk _096_ 0.00191f
C6318 net27 _312_/a_1108_47# 0.00178f
C6319 _300_/a_47_47# _133_ 4.7e-21
C6320 state\[2\] _107_ 0.0225f
C6321 _053_ _260_/a_346_47# 8.87e-19
C6322 _188_/a_27_47# clkc 7.28e-19
C6323 result[6] _314_/a_27_47# 0.00742f
C6324 net28 _314_/a_761_289# 0.00719f
C6325 _104_ trim_val\[3\] 5.05e-20
C6326 _059_ _087_ 6.38e-19
C6327 _064_ net50 0.465f
C6328 state\[2\] _166_/a_161_47# 0.0585f
C6329 _263_/a_79_21# _226_/a_27_47# 2.58e-19
C6330 _309_/a_27_47# _310_/a_193_47# 0.00127f
C6331 _309_/a_193_47# _310_/a_27_47# 6.43e-21
C6332 calibrate clknet_0_clk 1.42e-19
C6333 _120_ _090_ 0.0263f
C6334 clknet_2_1__leaf_clk net44 0.0461f
C6335 _326_/a_27_47# net43 0.0079f
C6336 VPWR _306_/a_1270_413# 4.74e-20
C6337 _319_/a_1108_47# _065_ 8.33e-19
C6338 _327_/a_1283_21# _109_ 1.29e-19
C6339 VPWR _161_/a_68_297# 0.0165f
C6340 _297_/a_129_47# net40 0.00189f
C6341 _056_ net33 0.0724f
C6342 _200_/a_80_21# net4 0.00116f
C6343 VPWR _314_/a_543_47# 0.0125f
C6344 _341_/a_761_289# _135_ 1.11e-20
C6345 _341_/a_1108_47# net2 2.97e-19
C6346 cal_count\[0\] _130_ 7.12e-22
C6347 _019_ mask\[2\] 0.3f
C6348 clknet_2_3__leaf_clk _108_ 1.78e-19
C6349 clk _318_/a_27_47# 0.0539f
C6350 clkbuf_0_clk/a_110_47# net30 0.00164f
C6351 net15 _101_ 0.749f
C6352 _066_ rebuffer3/a_75_212# 1.04e-19
C6353 _042_ _041_ 4.99e-19
C6354 _061_ _134_ 0.0033f
C6355 VPWR rebuffer4/a_27_47# 0.0671f
C6356 net31 trimb[2] 3.03e-20
C6357 _336_/a_27_47# _336_/a_761_289# -0.0169f
C6358 clknet_2_1__leaf_clk _003_ 3.91e-19
C6359 _102_ net26 0.408f
C6360 net9 _340_/a_562_413# 6.51e-19
C6361 output23/a_27_47# _308_/a_193_47# 2.18e-19
C6362 net12 _239_/a_474_297# 0.0104f
C6363 _185_/a_68_297# _092_ 5.9e-22
C6364 _007_ _082_ 0.025f
C6365 _307_/a_651_413# _074_ 0.00467f
C6366 _280_/a_75_212# net46 0.00431f
C6367 _059_ _263_/a_297_47# 0.00551f
C6368 _326_/a_651_413# net28 7.39e-20
C6369 net33 clkc 2.25e-19
C6370 _325_/a_1108_47# mask\[5\] 1.74e-20
C6371 _026_ _027_ 1.14e-19
C6372 VPWR _027_ 0.385f
C6373 _339_/a_1602_47# cal_count\[0\] 0.0475f
C6374 fanout43/a_27_47# _080_ 8.51e-19
C6375 _066_ _065_ 0.0196f
C6376 net4 _318_/a_27_47# 5.02e-19
C6377 net50 _057_ 8.88e-20
C6378 _050_ _281_/a_253_297# 3.07e-19
C6379 _243_/a_27_297# _100_ 0.0176f
C6380 cal_itt\[0\] _284_/a_68_297# 1.11e-19
C6381 _110_ _274_/a_75_212# 0.0044f
C6382 mask\[3\] _082_ 0.00334f
C6383 _089_ _062_ 5.29e-21
C6384 _087_ _075_ 0.00266f
C6385 _304_/a_651_413# _065_ 9.08e-20
C6386 _034_ _099_ 1.39e-21
C6387 _290_/a_27_413# output40/a_27_47# 0.0126f
C6388 net43 _314_/a_448_47# 1.1e-20
C6389 _317_/a_27_47# _316_/a_651_413# 2.78e-20
C6390 clk _317_/a_1270_413# 8.78e-20
C6391 net2 _339_/a_476_47# 1.28e-19
C6392 VPWR _195_/a_218_47# -4.07e-19
C6393 _282_/a_68_297# net30 1.63e-19
C6394 _169_/a_109_53# _185_/a_68_297# 0.00167f
C6395 trim_mask\[4\] _330_/a_27_47# 1.35e-21
C6396 clknet_2_2__leaf_clk _330_/a_1108_47# 0.0234f
C6397 VPWR _326_/a_1270_413# 1.23e-19
C6398 _329_/a_1270_413# _031_ 3.59e-20
C6399 VPWR _334_/a_1270_413# 5.03e-20
C6400 _048_ _120_ 0.0423f
C6401 _123_ _298_/a_78_199# 0.0124f
C6402 _327_/a_193_47# _058_ 0.042f
C6403 _328_/a_1108_47# trim_mask\[0\] 5.76e-19
C6404 clkbuf_0_clk/a_110_47# _072_ 0.0135f
C6405 fanout47/a_27_47# _069_ 0.0024f
C6406 _237_/a_76_199# clkbuf_2_0__f_clk/a_110_47# 8.03e-19
C6407 _258_/a_109_297# net9 7.53e-20
C6408 _092_ _118_ 9.2e-20
C6409 _015_ _099_ 3.09e-20
C6410 _331_/a_1108_47# _052_ 2.8e-19
C6411 net43 _310_/a_761_289# 0.00801f
C6412 mask\[1\] _246_/a_109_297# 1.35e-19
C6413 _325_/a_543_47# net27 1.05e-19
C6414 _071_ clk 6.42e-20
C6415 _330_/a_651_413# net19 0.00323f
C6416 net4 _317_/a_1270_413# 1.46e-19
C6417 net22 _282_/a_68_297# 1.48e-20
C6418 _335_/a_543_47# _119_ 1.05e-20
C6419 net14 _310_/a_805_47# 5.85e-19
C6420 _078_ _313_/a_651_413# 4.99e-19
C6421 _324_/a_761_289# _311_/a_1283_21# 5.29e-20
C6422 _324_/a_193_47# _311_/a_1108_47# 7.02e-21
C6423 _093_ net14 0.0132f
C6424 net30 _204_/a_75_212# 0.0371f
C6425 _048_ _076_ 1.71e-19
C6426 VPWR _300_/a_47_47# 0.0721f
C6427 net13 net51 4.16e-20
C6428 _064_ _181_/a_150_297# 4.36e-20
C6429 _337_/a_651_413# net45 6.88e-20
C6430 VPWR _335_/a_448_47# 0.0181f
C6431 _323_/a_761_289# net26 3.76e-20
C6432 _239_/a_474_297# _003_ 7.81e-21
C6433 _323_/a_448_47# _042_ 0.0161f
C6434 VPWR _311_/a_193_47# -0.28f
C6435 _053_ _279_/a_396_47# 0.00233f
C6436 _015_ _169_/a_215_311# 5.91e-19
C6437 _061_ cal_count\[3\] 5.28e-20
C6438 _097_ net4 0.00243f
C6439 _071_ net4 1.18e-21
C6440 mask\[2\] _205_/a_27_47# 3.88e-19
C6441 _239_/a_27_297# _098_ 0.00146f
C6442 VPWR _332_/a_1108_47# 0.00506f
C6443 _194_/a_113_297# _066_ 0.00178f
C6444 _121_ _192_/a_174_21# 7.67e-21
C6445 _255_/a_27_47# _051_ 6.49e-19
C6446 _093_ net41 1.4e-19
C6447 _074_ valid 0.0171f
C6448 _074_ net20 0.00949f
C6449 VPWR _029_ 0.0903f
C6450 _110_ _329_/a_1108_47# 2.85e-19
C6451 net12 _318_/a_805_47# 1.31e-19
C6452 _042_ net18 0.169f
C6453 _074_ net53 0.0143f
C6454 _290_/a_207_413# trimb[1] 7.14e-19
C6455 _326_/a_1270_413# net52 5.26e-21
C6456 net9 _338_/a_1602_47# 0.00333f
C6457 trim_mask\[2\] net48 0.0468f
C6458 _336_/a_543_47# _264_/a_27_297# 8.17e-20
C6459 output21/a_27_47# output20/a_27_47# 4.46e-21
C6460 result[1] _308_/a_448_47# 6.45e-20
C6461 _023_ _078_ 3.55e-19
C6462 _281_/a_337_297# _092_ 0.0013f
C6463 _339_/a_476_47# _123_ 0.0325f
C6464 net43 _305_/a_27_47# 0.625f
C6465 VPWR _310_/a_805_47# 4.15e-19
C6466 VPWR _093_ 0.653f
C6467 _204_/a_75_212# _072_ 2.13e-20
C6468 _340_/a_956_413# cal_count\[2\] 1.2e-20
C6469 _275_/a_81_21# _335_/a_543_47# 0.0059f
C6470 net47 _065_ 0.453f
C6471 _143_/a_150_297# _065_ 8.49e-22
C6472 calibrate _331_/a_1108_47# 7.33e-19
C6473 _188_/a_27_47# _136_ 3.66e-21
C6474 clknet_2_0__leaf_clk _316_/a_761_289# 6.07e-21
C6475 net45 _316_/a_27_47# 0.00846f
C6476 _337_/a_27_47# _096_ 0.00163f
C6477 _235_/a_382_297# net3 2.21e-19
C6478 _014_ _316_/a_193_47# 0.0222f
C6479 cal_itt\[0\] _341_/a_761_289# 1.25e-20
C6480 net12 net45 0.0673f
C6481 _266_/a_68_297# _108_ 0.00179f
C6482 clk wire42/a_75_212# 0.00295f
C6483 net43 net51 0.382f
C6484 _101_ _311_/a_543_47# 3.18e-21
C6485 _128_ cal_count\[0\] 0.0168f
C6486 _104_ trim_val\[4\] 0.0488f
C6487 _309_/a_193_47# clknet_2_1__leaf_clk 0.0019f
C6488 VPWR _285_/a_113_47# -1.08e-19
C6489 _327_/a_1462_47# _058_ 2.66e-19
C6490 _328_/a_1283_21# trim_mask\[2\] 6.44e-20
C6491 net24 _081_ 0.164f
C6492 _020_ mask\[4\] 8.9e-20
C6493 net12 _103_ 8.81e-21
C6494 clknet_2_2__leaf_clk _052_ 2.54e-20
C6495 _052_ _260_/a_584_47# 0.00318f
C6496 _311_/a_805_47# net53 2.96e-19
C6497 mask\[1\] _017_ 0.00367f
C6498 clknet_0_clk _203_/a_59_75# 0.00228f
C6499 net46 net19 0.00497f
C6500 _115_ net48 0.0183f
C6501 net12 _065_ 0.0165f
C6502 _134_ net16 0.335f
C6503 clknet_0_clk _192_/a_27_47# 0.0127f
C6504 _175_/a_68_297# rebuffer1/a_75_212# 0.0215f
C6505 _333_/a_1283_21# net37 9e-19
C6506 cal_itt\[0\] clknet_0_clk 0.00304f
C6507 _333_/a_193_47# rebuffer1/a_75_212# 1.72e-20
C6508 _333_/a_27_47# _332_/a_27_47# 5.12e-19
C6509 _259_/a_373_47# _104_ 0.00109f
C6510 _324_/a_27_47# _042_ 7.87e-20
C6511 net44 net45 0.00208f
C6512 VPWR _032_ 0.0765f
C6513 _008_ _074_ 0.00334f
C6514 _306_/a_27_47# fanout44/a_27_47# 3.47e-21
C6515 _307_/a_1283_21# _210_/a_113_297# 3.48e-20
C6516 _259_/a_27_297# _330_/a_27_47# 1.16e-20
C6517 VPWR _305_/a_1270_413# -2.07e-19
C6518 net50 _027_ 0.002f
C6519 trim_mask\[3\] net46 0.0625f
C6520 net26 clknet_2_3__leaf_clk 8.28e-19
C6521 VPWR _311_/a_1462_47# 7.21e-20
C6522 output22/a_27_47# net22 0.0133f
C6523 _051_ _336_/a_27_47# 5.67e-19
C6524 _324_/a_1283_21# clknet_2_1__leaf_clk 9.42e-19
C6525 _289_/a_68_297# trimb[4] 1.71e-19
C6526 _329_/a_543_47# net9 0.00535f
C6527 output34/a_27_47# _334_/a_27_47# 4.36e-20
C6528 net33 _172_/a_68_297# 0.00219f
C6529 _136_ net33 3.56e-20
C6530 _335_/a_1108_47# clknet_2_2__leaf_clk 8.02e-20
C6531 _335_/a_27_47# trim_mask\[4\] 1.83e-22
C6532 net16 _130_ 0.0061f
C6533 net43 _224_/a_199_47# 1.59e-19
C6534 _302_/a_109_297# _066_ 0.0635f
C6535 calibrate _263_/a_79_21# 3.97e-19
C6536 clkbuf_0_clk/a_110_47# _230_/a_59_75# 8.11e-20
C6537 _107_ net46 0.00233f
C6538 _110_ _280_/a_75_212# 7.08e-22
C6539 net15 _241_/a_297_47# 0.00587f
C6540 output29/a_27_47# net14 0.0211f
C6541 _304_/a_27_47# _136_ 0.00313f
C6542 net44 _065_ 0.752f
C6543 _067_ _070_ 0.0659f
C6544 output39/a_27_47# net34 4.68e-19
C6545 _058_ en_co_clk 9.63e-19
C6546 _333_/a_1108_47# net46 -1.41e-19
C6547 _243_/a_109_47# clone7/a_27_47# 1.5e-19
C6548 _237_/a_505_21# _049_ 8.24e-19
C6549 _323_/a_1283_21# _150_/a_27_47# 2.18e-19
C6550 net45 _003_ 1.36e-21
C6551 ctln[3] net18 2.83e-20
C6552 mask\[3\] _076_ 7.04e-19
C6553 _304_/a_27_47# _284_/a_68_297# 1.21e-20
C6554 _083_ _311_/a_193_47# 5.05e-19
C6555 _303_/a_193_47# net26 4.16e-20
C6556 _332_/a_1283_21# clknet_2_2__leaf_clk 2.36e-21
C6557 _059_ _099_ 0.0305f
C6558 result[1] _005_ 0.077f
C6559 _341_/a_27_47# rebuffer3/a_75_212# 2.11e-19
C6560 _122_ cal_count\[2\] 0.136f
C6561 _264_/a_27_297# _106_ 0.00629f
C6562 _304_/a_761_289# net47 2.67e-19
C6563 cal_itt\[2\] clknet_2_3__leaf_clk 2.4e-19
C6564 _111_ clknet_2_2__leaf_clk 0.0731f
C6565 _164_/a_161_47# _093_ 0.0694f
C6566 net43 _305_/a_1217_47# -5.37e-19
C6567 net13 _318_/a_193_47# 0.0212f
C6568 net16 _339_/a_1602_47# 0.00389f
C6569 _308_/a_1283_21# net22 8.92e-21
C6570 _308_/a_761_289# _078_ 3.77e-19
C6571 trim_mask\[0\] _100_ 1.03e-20
C6572 _321_/a_27_47# _321_/a_639_47# -0.0015f
C6573 mask\[6\] net14 4.06e-22
C6574 _037_ cal_count\[2\] 2.99e-19
C6575 _319_/a_1108_47# _282_/a_68_297# 4.85e-20
C6576 net50 _335_/a_448_47# 7.97e-20
C6577 clkbuf_2_0__f_clk/a_110_47# _090_ 0.00855f
C6578 net44 _319_/a_27_47# 3.16e-20
C6579 _308_/a_27_47# clknet_2_0__leaf_clk 0.0323f
C6580 _262_/a_193_297# clkbuf_2_3__f_clk/a_110_47# 0.00178f
C6581 _065_ _003_ 0.0016f
C6582 _299_/a_27_413# cal_count\[2\] 0.0242f
C6583 _019_ _074_ 7.53e-20
C6584 clk _202_/a_79_21# 1.37e-19
C6585 _060_ en_co_clk 0.00965f
C6586 _317_/a_448_47# net14 1.74e-19
C6587 _314_/a_27_47# _158_/a_68_297# 2.64e-21
C6588 _307_/a_193_47# _315_/a_1108_47# 5.53e-21
C6589 _307_/a_1108_47# _315_/a_193_47# 5.53e-21
C6590 net45 _316_/a_1217_47# -1.47e-19
C6591 _341_/a_27_47# _065_ 0.0135f
C6592 VPWR _272_/a_384_47# -1.05e-19
C6593 _119_ _170_/a_81_21# 5.69e-21
C6594 _051_ _096_ 4.33e-21
C6595 trim[1] _333_/a_1283_21# 3.74e-20
C6596 _250_/a_27_297# _101_ 0.00747f
C6597 clknet_2_0__leaf_clk clknet_0_clk 0.822f
C6598 _306_/a_1283_21# _092_ 1.19e-19
C6599 _337_/a_27_47# _337_/a_639_47# -0.0015f
C6600 _313_/a_27_47# _313_/a_193_47# -0.324f
C6601 cal_itt\[0\] _303_/a_27_47# 1.17e-19
C6602 cal_count\[3\] _049_ 5.13e-20
C6603 result[4] result[5] 0.049f
C6604 _320_/a_543_47# net45 4.02e-20
C6605 _320_/a_1108_47# clknet_2_0__leaf_clk 1.96e-19
C6606 VPWR output29/a_27_47# 0.0655f
C6607 net9 _339_/a_381_47# 0.00292f
C6608 output32/a_27_47# _109_ 4.83e-20
C6609 net46 _279_/a_27_47# 0.00143f
C6610 VPWR _171_/a_27_47# 0.108f
C6611 net16 cal_count\[3\] 2.33e-19
C6612 _053_ _193_/a_109_297# 1.93e-19
C6613 _074_ _312_/a_805_47# 2.48e-21
C6614 VPWR _239_/a_277_297# -0.0103f
C6615 _287_/a_75_212# _338_/a_193_47# 0.00801f
C6616 _078_ _140_/a_68_297# 0.00199f
C6617 _064_ _278_/a_109_297# 5.72e-19
C6618 net26 net53 0.132f
C6619 net4 _194_/a_199_47# 2.28e-19
C6620 _331_/a_27_47# _049_ 2.8e-20
C6621 net47 _043_ 0.0686f
C6622 trim_mask\[0\] _264_/a_27_297# 5.26e-21
C6623 _097_ _237_/a_535_374# 1.33e-19
C6624 net4 _336_/a_1108_47# 0.00131f
C6625 _062_ _092_ 0.0592f
C6626 _075_ _099_ 3.69e-19
C6627 _324_/a_761_289# _021_ 1.27e-19
C6628 _312_/a_193_47# _221_/a_109_297# 8.06e-20
C6629 _333_/a_651_413# rebuffer2/a_75_212# 1.13e-19
C6630 _333_/a_1270_413# _108_ 2.09e-19
C6631 _181_/a_68_297# net46 2.99e-19
C6632 _320_/a_543_47# _065_ 8.11e-20
C6633 _307_/a_805_47# net22 7.15e-19
C6634 _307_/a_1270_413# _078_ 1.06e-19
C6635 _064_ _330_/a_543_47# 1.16e-21
C6636 _104_ _330_/a_193_47# 1.8e-20
C6637 VPWR mask\[6\] 0.427f
C6638 trim_val\[0\] _332_/a_1283_21# 0.0101f
C6639 _109_ _332_/a_193_47# 0.00209f
C6640 output16/a_27_47# net39 0.01f
C6641 _307_/a_1283_21# net45 0.0133f
C6642 _307_/a_448_47# clknet_2_0__leaf_clk 0.00107f
C6643 trim[3] _334_/a_1108_47# 4.32e-19
C6644 _111_ trim_val\[0\] 4.54e-20
C6645 VPWR _317_/a_448_47# -0.00293f
C6646 _315_/a_193_47# net14 0.0145f
C6647 _038_ _066_ 0.256f
C6648 net27 result[5] 0.00273f
C6649 clkbuf_2_0__f_clk/a_110_47# _048_ 0.012f
C6650 _094_ _095_ 0.0016f
C6651 _304_/a_651_413# _038_ 2.17e-20
C6652 _304_/a_1217_47# _136_ 1.02e-19
C6653 _101_ _009_ 5.33e-21
C6654 _316_/a_1283_21# _096_ 6.93e-20
C6655 _338_/a_27_47# _067_ 1.25e-19
C6656 VPWR _203_/a_145_75# -4.82e-19
C6657 output36/a_27_47# trimb[1] 6.66e-20
C6658 trimb[0] output37/a_27_47# 0.00178f
C6659 _304_/a_543_47# _122_ 0.0129f
C6660 net4 _035_ 3.57e-20
C6661 VPWR _192_/a_505_280# -1.72e-19
C6662 _341_/a_193_47# _304_/a_193_47# 1.89e-21
C6663 _341_/a_27_47# _304_/a_761_289# 9.3e-20
C6664 cal_itt\[1\] VPWR 0.579f
C6665 _315_/a_193_47# net41 2.66e-21
C6666 _340_/a_1032_413# net47 0.00241f
C6667 _037_ _304_/a_543_47# 2.7e-19
C6668 _060_ _235_/a_297_47# 1.12e-19
C6669 ctln[7] _318_/a_805_47# 2.48e-20
C6670 net13 _318_/a_1462_47# 1.57e-19
C6671 _108_ _279_/a_314_297# 0.00313f
C6672 _259_/a_27_297# _335_/a_27_47# 2.31e-19
C6673 net50 _032_ 0.0063f
C6674 _113_ _109_ 3.58e-19
C6675 _262_/a_193_297# cal_count\[3\] 5.67e-19
C6676 clknet_2_1__leaf_clk net19 5.46e-19
C6677 _043_ net44 1.13e-20
C6678 _074_ _205_/a_27_47# 0.00604f
C6679 _008_ net26 0.317f
C6680 _129_ _131_ 0.00885f
C6681 _059_ _053_ 4.32e-20
C6682 net24 net14 0.00633f
C6683 state\[2\] _062_ 2.69e-21
C6684 _014_ net14 3.31e-19
C6685 _309_/a_1108_47# _078_ 0.0499f
C6686 _010_ _223_/a_109_297# 0.0011f
C6687 clone1/a_27_47# _098_ 0.0229f
C6688 clk fanout45/a_27_47# 0.00263f
C6689 _128_ net16 0.0758f
C6690 _110_ net19 0.0477f
C6691 VPWR _315_/a_193_47# -0.115f
C6692 clkbuf_0_clk/a_110_47# net47 3.95e-19
C6693 _237_/a_505_21# state\[1\] 3.95e-20
C6694 mask\[6\] net52 0.201f
C6695 _309_/a_761_289# net24 0.0191f
C6696 _337_/a_761_289# net44 6.81e-19
C6697 net35 net37 0.0143f
C6698 _068_ _190_/a_27_47# 0.00106f
C6699 net28 _225_/a_109_297# 3.5e-19
C6700 cal_itt\[0\] _303_/a_1217_47# 1.13e-19
C6701 _309_/a_193_47# net45 2.05e-19
C6702 _336_/a_448_47# clkbuf_2_2__f_clk/a_110_47# 9.38e-19
C6703 _291_/a_35_297# _290_/a_207_413# 0.0019f
C6704 _304_/a_27_47# clknet_0_clk 1.69e-20
C6705 VPWR _318_/a_639_47# 0.001f
C6706 _112_ clknet_2_2__leaf_clk 0.00632f
C6707 _082_ _310_/a_761_289# 0.00213f
C6708 net25 _310_/a_1108_47# 0.0513f
C6709 mask\[3\] _310_/a_1283_21# 0.00292f
C6710 _035_ _122_ 3.09e-20
C6711 net46 _118_ 6.17e-20
C6712 _116_ trim_val\[3\] 0.00302f
C6713 _110_ trim_mask\[3\] 0.121f
C6714 _327_/a_1283_21# net46 0.0151f
C6715 _294_/a_150_297# _129_ 1.39e-19
C6716 ctln[7] net45 3.98e-19
C6717 _304_/a_27_47# _339_/a_27_47# 2.67e-20
C6718 clknet_0_clk clone1/a_27_47# 1.68e-20
C6719 _035_ _338_/a_381_47# 0.00385f
C6720 _076_ rebuffer5/a_161_47# 0.0222f
C6721 _258_/a_109_297# _033_ 6.44e-20
C6722 _162_/a_27_47# _055_ 1.54e-20
C6723 net24 _040_ 1.22e-19
C6724 _189_/a_27_47# _050_ 0.0399f
C6725 _014_ net41 0.00917f
C6726 fanout45/a_27_47# net4 0.0551f
C6727 _312_/a_448_47# _009_ 0.00196f
C6728 _110_ _107_ 0.0146f
C6729 _328_/a_639_47# VPWR 3.07e-19
C6730 _330_/a_27_47# _330_/a_639_47# -0.0015f
C6731 cal_itt\[1\] _063_ 0.257f
C6732 _288_/a_59_75# net37 0.00414f
C6733 _291_/a_35_297# _289_/a_68_297# 3.32e-19
C6734 VPWR net24 1.33f
C6735 _059_ _226_/a_109_47# 8.6e-21
C6736 _064_ _195_/a_505_21# 1.39e-19
C6737 _306_/a_27_47# _076_ 0.0196f
C6738 VPWR _014_ 0.624f
C6739 _304_/a_193_47# _133_ 0.0012f
C6740 _019_ net26 6.44e-20
C6741 net10 output9/a_27_47# 3.69e-20
C6742 _328_/a_193_47# _025_ 9.1e-19
C6743 VPWR output39/a_27_47# 0.0495f
C6744 net9 _025_ 9.33e-19
C6745 net47 _038_ 4.05e-20
C6746 _322_/a_543_47# net45 4.28e-20
C6747 _341_/a_193_47# _302_/a_27_297# 4.26e-20
C6748 _341_/a_27_47# _302_/a_109_297# 5.29e-20
C6749 net45 _331_/a_543_47# 0.00173f
C6750 _242_/a_297_47# _049_ 0.00675f
C6751 _326_/a_761_289# net27 4.37e-19
C6752 _326_/a_27_47# result[5] 0.00691f
C6753 clkbuf_2_0__f_clk/a_110_47# _283_/a_75_212# 3.13e-21
C6754 net43 _086_ 0.011f
C6755 clkbuf_0_clk/a_110_47# net44 0.00349f
C6756 _083_ mask\[6\] 6.36e-20
C6757 _164_/a_161_47# _192_/a_505_280# 1.86e-20
C6758 _321_/a_1283_21# _320_/a_193_47# 1.97e-19
C6759 _218_/a_113_297# _078_ 0.0315f
C6760 _208_/a_76_199# rebuffer4/a_27_47# 5.21e-19
C6761 _321_/a_1108_47# _320_/a_27_47# 3.64e-21
C6762 _297_/a_129_47# _132_ -5.62e-19
C6763 trim_val\[2\] _175_/a_150_297# 7.85e-19
C6764 _325_/a_193_47# _042_ 2.83e-19
C6765 clknet_2_1__leaf_clk _155_/a_68_297# 0.0393f
C6766 _143_/a_68_297# _041_ 0.00382f
C6767 _340_/a_1602_47# _122_ 0.00134f
C6768 _112_ _333_/a_651_413# 8.3e-19
C6769 net49 _333_/a_1270_413# 1.1e-19
C6770 net47 _338_/a_476_47# 0.051f
C6771 _337_/a_27_47# clknet_0_clk 0.0239f
C6772 trim[1] net35 0.0359f
C6773 _235_/a_297_47# en_co_clk 0.00145f
C6774 _258_/a_109_297# _024_ 6.81e-20
C6775 net13 _243_/a_373_47# 1.99e-19
C6776 _325_/a_1108_47# clknet_2_1__leaf_clk 5.88e-20
C6777 _093_ _034_ 1.2e-21
C6778 _104_ _335_/a_193_47# 0.0025f
C6779 _340_/a_1602_47# _037_ 5.93e-20
C6780 fanout46/a_27_47# trim_val\[4\] 0.00159f
C6781 _239_/a_474_297# _107_ 0.00144f
C6782 net23 net24 3.22e-19
C6783 _110_ _279_/a_27_47# 0.00639f
C6784 net16 _175_/a_150_297# 3.12e-19
C6785 _243_/a_27_297# net41 2.57e-19
C6786 _327_/a_448_47# _111_ 9.03e-20
C6787 _328_/a_27_47# trim_val\[3\] 8.55e-21
C6788 net16 _333_/a_761_289# 0.00842f
C6789 result[4] _310_/a_1283_21# 3.24e-19
C6790 mask\[7\] _023_ 4.85e-19
C6791 mask\[4\] _311_/a_1108_47# 0.0402f
C6792 net16 _265_/a_299_297# 0.00719f
C6793 VPWR _315_/a_1462_47# 4.59e-19
C6794 net12 _204_/a_75_212# 0.00856f
C6795 _313_/a_448_47# _010_ 0.00355f
C6796 _033_ clkbuf_2_2__f_clk/a_110_47# 0.065f
C6797 _058_ _332_/a_639_47# 8.33e-19
C6798 _050_ _227_/a_109_93# 1.83e-20
C6799 _334_/a_1108_47# _057_ 2.11e-20
C6800 _189_/a_218_47# _092_ 0.00259f
C6801 _015_ _093_ 0.0433f
C6802 VPWR _243_/a_27_297# -0.0126f
C6803 clknet_2_1__leaf_clk _248_/a_109_297# 6.27e-22
C6804 net24 net52 0.0116f
C6805 _110_ _181_/a_68_297# 3.09e-19
C6806 _328_/a_1283_21# _333_/a_27_47# 8.44e-21
C6807 _314_/a_27_47# _085_ 1.58e-21
C6808 _340_/a_27_47# _339_/a_476_47# 1.06e-20
C6809 net31 comp 0.149f
C6810 _340_/a_476_47# _339_/a_27_47# 8.3e-21
C6811 clk _316_/a_651_413# 1.11e-19
C6812 _316_/a_27_47# _316_/a_448_47# -0.00719f
C6813 mask\[1\] clknet_2_1__leaf_clk 0.00928f
C6814 _041_ net4 0.0577f
C6815 _297_/a_47_47# _131_ 3.37e-19
C6816 net44 _204_/a_75_212# 1.06e-20
C6817 _171_/a_27_47# _279_/a_396_47# 2.25e-20
C6818 _330_/a_543_47# _027_ 0.0336f
C6819 _330_/a_761_289# net46 -0.0067f
C6820 _336_/a_27_47# _119_ 0.0126f
C6821 output27/a_27_47# _074_ 2.17e-20
C6822 net43 _319_/a_761_289# -0.00611f
C6823 _067_ clknet_2_3__leaf_clk 0.0407f
C6824 clknet_2_3__leaf_clk _070_ 2.49e-20
C6825 _323_/a_1108_47# net47 0.00305f
C6826 net42 _050_ 0.00488f
C6827 _158_/a_150_297# net29 2.03e-19
C6828 _232_/a_32_297# _092_ 0.00648f
C6829 VPWR _336_/a_543_47# 0.0132f
C6830 _328_/a_1270_413# clknet_2_2__leaf_clk 2.74e-19
C6831 VPWR _304_/a_193_47# 0.0302f
C6832 _007_ _042_ 0.00131f
C6833 _340_/a_1182_261# _133_ 9.84e-20
C6834 mask\[6\] _155_/a_150_297# 2.29e-19
C6835 _340_/a_652_21# clknet_2_3__leaf_clk 9.5e-21
C6836 _341_/a_1283_21# _136_ 0.00872f
C6837 _341_/a_27_47# _038_ 0.0854f
C6838 _048_ cal_itt\[3\] 2.38e-19
C6839 _051_ _098_ 0.00265f
C6840 _020_ _311_/a_1108_47# 1.4e-20
C6841 _042_ _249_/a_27_297# 0.0295f
C6842 _041_ _122_ 0.0417f
C6843 _325_/a_193_47# _022_ 0.111f
C6844 _325_/a_448_47# mask\[6\] 0.0248f
C6845 _204_/a_75_212# _003_ 0.00223f
C6846 _338_/a_1182_261# _122_ 0.00536f
C6847 _319_/a_193_47# _101_ 0.00234f
C6848 mask\[3\] _042_ 0.754f
C6849 _169_/a_109_53# _232_/a_32_297# 1.51e-20
C6850 net47 _338_/a_1224_47# 8.53e-19
C6851 _303_/a_193_47# _067_ 9.32e-21
C6852 net3 _192_/a_639_47# 0.00129f
C6853 _314_/a_27_47# _314_/a_543_47# -1.48e-19
C6854 _303_/a_193_47# _070_ 1.44e-19
C6855 _258_/a_373_47# trim_mask\[2\] 5.31e-19
C6856 _239_/a_694_21# _095_ 1.94e-20
C6857 net13 _321_/a_1283_21# 0.0043f
C6858 _037_ _041_ 1.72e-20
C6859 _051_ clknet_0_clk 1.46f
C6860 output21/a_27_47# VPWR 0.0969f
C6861 _048_ _262_/a_205_47# 3.16e-19
C6862 _050_ _054_ 0.0156f
C6863 net13 _337_/a_1283_21# 2.47e-19
C6864 _110_ _118_ 0.0398f
C6865 _050_ net30 4.74e-19
C6866 net2 comp 0.00749f
C6867 _110_ _327_/a_1283_21# 4.67e-19
C6868 _040_ _337_/a_193_47# 4.4e-20
C6869 _236_/a_109_297# clknet_2_0__leaf_clk 1.15e-20
C6870 _336_/a_193_47# _266_/a_68_297# 2.02e-21
C6871 _104_ _189_/a_27_47# 6.3e-22
C6872 VPWR _319_/a_805_47# 1.2e-19
C6873 _168_/a_27_413# _050_ 0.0376f
C6874 VPWR _321_/a_193_47# 0.0182f
C6875 _065_ net19 0.00893f
C6876 _330_/a_1108_47# _108_ 5.54e-22
C6877 clknet_2_0__leaf_clk _209_/a_27_47# 3.24e-21
C6878 _323_/a_1108_47# net44 5.49e-20
C6879 trim[4] _332_/a_1283_21# 4.74e-19
C6880 _305_/a_193_47# en_co_clk 3.91e-21
C6881 _336_/a_543_47# _063_ 2.94e-21
C6882 output33/a_27_47# trim[3] 6.66e-20
C6883 trim[2] output34/a_27_47# 0.00212f
C6884 state\[2\] _232_/a_32_297# 1.3e-19
C6885 net47 _339_/a_1182_261# -0.00352f
C6886 VPWR _337_/a_193_47# -0.0383f
C6887 _267_/a_59_75# _332_/a_27_47# 0.00126f
C6888 _304_/a_193_47# _063_ 0.00209f
C6889 _323_/a_193_47# _323_/a_543_47# -0.0129f
C6890 _258_/a_109_47# net18 2.46e-19
C6891 _105_ net19 0.0167f
C6892 _316_/a_27_47# _013_ 0.0849f
C6893 _061_ en_co_clk 0.00756f
C6894 net4 net18 4.59e-22
C6895 _195_/a_439_47# _062_ 5.31e-19
C6896 _189_/a_408_47# _053_ 1.94e-19
C6897 _097_ _241_/a_297_47# 0.0499f
C6898 trim_mask\[2\] _274_/a_75_212# 0.036f
C6899 _192_/a_174_21# _095_ 0.0458f
C6900 _103_ _107_ 0.0467f
C6901 _089_ _100_ 0.243f
C6902 _087_ _096_ 3.13e-20
C6903 VPWR _302_/a_27_297# 0.0275f
C6904 ctlp[0] _314_/a_639_47# 3.92e-20
C6905 _305_/a_27_47# _076_ 0.0104f
C6906 _308_/a_193_47# _006_ 4.59e-21
C6907 _308_/a_543_47# _081_ 7.83e-20
C6908 _292_/a_78_199# _340_/a_1182_261# 0.00813f
C6909 _122_ _298_/a_493_297# 3.43e-19
C6910 _306_/a_193_47# _305_/a_193_47# 3.79e-20
C6911 _306_/a_761_289# _305_/a_27_47# 1.38e-19
C6912 _064_ trim_mask\[1\] 0.133f
C6913 _001_ _065_ 0.326f
C6914 _326_/a_543_47# _310_/a_193_47# 5.84e-21
C6915 _326_/a_193_47# _310_/a_543_47# 1.44e-20
C6916 _326_/a_27_47# _310_/a_1283_21# 3.63e-19
C6917 net43 _321_/a_1283_21# 0.0124f
C6918 VPWR _106_ 0.16f
C6919 _338_/a_27_47# clknet_2_3__leaf_clk 0.568f
C6920 output20/a_27_47# _312_/a_193_47# 0.00122f
C6921 _320_/a_27_47# _320_/a_193_47# -0.0563f
C6922 _334_/a_1283_21# net46 1.53e-20
C6923 _107_ _105_ 0.00862f
C6924 state\[2\] _227_/a_209_311# 4.33e-19
C6925 _266_/a_68_297# net55 5.3e-21
C6926 VPWR _340_/a_1182_261# -0.00119f
C6927 _329_/a_27_47# _274_/a_75_212# 8.25e-21
C6928 net43 _313_/a_27_47# 0.00973f
C6929 _341_/a_1217_47# _038_ 1.94e-20
C6930 _059_ _093_ 9.99e-21
C6931 _315_/a_1108_47# _241_/a_105_352# 5.06e-20
C6932 _336_/a_193_47# _028_ 6.93e-20
C6933 _336_/a_761_289# clknet_2_2__leaf_clk 0.00214f
C6934 _237_/a_76_199# net4 5.62e-20
C6935 _328_/a_27_47# trim_val\[4\] 3.04e-21
C6936 _058_ net16 0.0446f
C6937 net51 _076_ 0.0912f
C6938 _122_ net18 0.155f
C6939 _319_/a_1270_413# _016_ 1.55e-20
C6940 result[5] _224_/a_199_47# 5.81e-21
C6941 net17 _339_/a_193_47# 1.07e-20
C6942 _325_/a_639_47# _078_ 1.55e-19
C6943 _188_/a_27_47# trim_val\[0\] 1.76e-19
C6944 _321_/a_193_47# net52 0.0131f
C6945 _321_/a_543_47# _101_ 0.0338f
C6946 _190_/a_27_47# cal_itt\[3\] 0.0147f
C6947 _306_/a_761_289# net51 2.89e-19
C6948 _338_/a_381_47# net18 0.00126f
C6949 _081_ _140_/a_150_297# 0.00117f
C6950 _341_/a_193_47# _341_/a_1108_47# -0.00656f
C6951 _341_/a_27_47# _341_/a_448_47# -0.00656f
C6952 net31 _161_/a_150_297# 2.19e-20
C6953 _122_ _129_ 0.00432f
C6954 _320_/a_639_47# net44 -7.75e-19
C6955 _088_ _052_ 0.0304f
C6956 _263_/a_382_297# net55 0.00139f
C6957 _263_/a_297_47# _096_ 1.97e-20
C6958 _037_ net18 1.21e-20
C6959 _104_ _227_/a_109_93# 0.00139f
C6960 net47 _303_/a_1283_21# 0.0655f
C6961 _303_/a_193_47# _338_/a_27_47# 0.00228f
C6962 _303_/a_27_47# _338_/a_193_47# 7.98e-21
C6963 _071_ _190_/a_655_47# 6.61e-21
C6964 _231_/a_161_47# _194_/a_113_297# 3.63e-19
C6965 _335_/a_761_289# net46 0.0226f
C6966 _335_/a_543_47# _027_ 5.87e-19
C6967 _328_/a_761_289# _058_ 0.0021f
C6968 _274_/a_75_212# _115_ 0.00885f
C6969 _053_ _170_/a_81_21# 0.0382f
C6970 _060_ _049_ 0.00176f
C6971 _299_/a_27_413# _129_ 0.00788f
C6972 output27/a_27_47# net26 5.05e-21
C6973 mask\[0\] _092_ 2e-19
C6974 net27 _042_ 9.12e-20
C6975 _329_/a_1108_47# trim_mask\[2\] 0.00166f
C6976 _026_ trim_mask\[0\] 1.75e-20
C6977 VPWR trim_mask\[0\] 2.81f
C6978 VPWR _321_/a_1462_47# 2.24e-19
C6979 _286_/a_76_199# cal_count\[0\] 9.76e-19
C6980 _286_/a_218_374# _124_ 2.88e-19
C6981 net3 _243_/a_373_47# 1.2e-19
C6982 _339_/a_1032_413# _122_ 0.00357f
C6983 _332_/a_193_47# net46 0.568f
C6984 _194_/a_113_297# _107_ 5.69e-20
C6985 _110_ _330_/a_761_289# 2.26e-19
C6986 _258_/a_109_297# _257_/a_27_297# 1.18e-19
C6987 clkbuf_2_1__f_clk/a_110_47# net15 0.11f
C6988 VPWR _313_/a_1270_413# 3.73e-20
C6989 net47 _339_/a_1296_47# -7.83e-19
C6990 VPWR _337_/a_1462_47# 2.55e-19
C6991 net31 net46 9.91e-19
C6992 _106_ _063_ 0.0362f
C6993 _336_/a_1283_21# _107_ 3.14e-19
C6994 _199_/a_109_297# _070_ 1.38e-19
C6995 _307_/a_27_47# _307_/a_543_47# -0.00172f
C6996 _307_/a_193_47# _307_/a_761_289# -0.00659f
C6997 _104_ net42 1.36e-20
C6998 mask\[1\] net45 0.124f
C6999 trim_val\[0\] net33 0.0273f
C7000 _304_/a_761_289# _001_ 6.85e-20
C7001 _298_/a_78_199# _133_ 0.0954f
C7002 _310_/a_193_47# _310_/a_1108_47# -0.00817f
C7003 _156_/a_27_47# _009_ 1.44e-19
C7004 _329_/a_27_47# _329_/a_1108_47# -3.92e-19
C7005 _185_/a_68_297# net45 3.5e-20
C7006 net21 _313_/a_193_47# 8.73e-19
C7007 _046_ _313_/a_543_47# 2.94e-19
C7008 _159_/a_27_47# _313_/a_651_413# 8.84e-19
C7009 _335_/a_27_47# _335_/a_639_47# -0.0014f
C7010 state\[2\] _318_/a_1108_47# 0.00213f
C7011 _303_/a_1108_47# net4 1.61e-19
C7012 trimb[2] net34 0.0773f
C7013 _043_ net19 0.0119f
C7014 net26 _208_/a_218_374# 6.87e-20
C7015 _036_ _340_/a_1182_261# 7.23e-19
C7016 _023_ net28 2.04e-20
C7017 _301_/a_285_47# clknet_2_3__leaf_clk 0.0449f
C7018 _320_/a_651_413# clknet_0_clk 4.43e-19
C7019 mask\[1\] _065_ 0.00925f
C7020 _326_/a_651_413# _074_ 0.0022f
C7021 _313_/a_1108_47# _312_/a_27_47# 1.26e-20
C7022 _313_/a_1283_21# _312_/a_193_47# 9.64e-21
C7023 VPWR _338_/a_652_21# -0.00108f
C7024 _239_/a_694_21# _226_/a_27_47# 0.00111f
C7025 _341_/a_543_47# clknet_2_3__leaf_clk 0.0431f
C7026 _309_/a_448_47# _081_ 2.48e-21
C7027 _309_/a_1283_21# _006_ 4.1e-20
C7028 calibrate _088_ 0.218f
C7029 state\[0\] _192_/a_174_21# 1.68e-21
C7030 _113_ net46 0.14f
C7031 _323_/a_193_47# _303_/a_761_289# 4e-21
C7032 _323_/a_27_47# _303_/a_543_47# 1.23e-20
C7033 _323_/a_543_47# _303_/a_27_47# 1.92e-20
C7034 _323_/a_761_289# _303_/a_193_47# 1.8e-21
C7035 _316_/a_1108_47# net41 0.0403f
C7036 VPWR _340_/a_1296_47# 5.16e-19
C7037 _104_ _054_ 0.0343f
C7038 net43 _313_/a_1217_47# -3.08e-19
C7039 _329_/a_1108_47# _115_ 5.13e-21
C7040 _339_/a_27_47# _339_/a_652_21# -0.00883f
C7041 fanout46/a_27_47# _335_/a_193_47# 1.22e-19
C7042 net13 _320_/a_27_47# 0.00721f
C7043 _104_ net30 0.499f
C7044 _322_/a_761_289# _041_ 5.07e-21
C7045 _308_/a_1283_21# _307_/a_1283_21# 5.14e-19
C7046 trim_mask\[0\] _063_ 0.271f
C7047 net4 _191_/a_27_297# 8.17e-19
C7048 _307_/a_27_47# _138_/a_27_47# 0.0025f
C7049 rebuffer3/a_75_212# _118_ 1.4e-20
C7050 _336_/a_543_47# _279_/a_396_47# 0.00228f
C7051 _336_/a_1283_21# _279_/a_27_47# 0.00531f
C7052 _326_/a_543_47# _224_/a_113_297# 2.12e-19
C7053 _108_ rebuffer2/a_75_212# 0.0178f
C7054 _050_ _319_/a_1108_47# 3.91e-20
C7055 VPWR _316_/a_1108_47# 0.0275f
C7056 _104_ _168_/a_27_413# 7.15e-20
C7057 _332_/a_193_47# _332_/a_448_47# -0.00779f
C7058 _303_/a_1108_47# _338_/a_381_47# 5.79e-20
C7059 net2 net46 1.9e-19
C7060 _029_ _332_/a_761_289# 9.46e-20
C7061 _111_ _108_ 0.0474f
C7062 _294_/a_68_297# net16 2.83e-19
C7063 en_co_clk _049_ 0.459f
C7064 trimb[1] trimb[4] 0.0486f
C7065 _051_ _263_/a_79_21# 0.0135f
C7066 clk _331_/a_805_47# 5.18e-19
C7067 _185_/a_68_297# _243_/a_109_297# 7.35e-20
C7068 _162_/a_27_47# _333_/a_1283_21# 0.00139f
C7069 net16 en_co_clk 0.045f
C7070 trim_mask\[2\] _280_/a_75_212# 0.0345f
C7071 _339_/a_193_47# clknet_2_3__leaf_clk 4.7e-19
C7072 _110_ _062_ 3.13e-19
C7073 _181_/a_68_297# _336_/a_1283_21# 0.00107f
C7074 clkbuf_2_2__f_clk/a_110_47# _331_/a_27_47# 3.93e-19
C7075 net50 _106_ 2.39e-21
C7076 _333_/a_543_47# net32 1.22e-19
C7077 _319_/a_1283_21# _283_/a_75_212# 8.51e-19
C7078 _326_/a_193_47# _251_/a_27_297# 5.49e-20
C7079 _324_/a_805_47# net44 5.85e-19
C7080 _090_ clone7/a_27_47# 6.18e-19
C7081 _332_/a_1462_47# net46 -9.14e-19
C7082 net15 _317_/a_193_47# 0.0174f
C7083 _292_/a_78_199# _298_/a_78_199# 8.87e-19
C7084 cal_itt\[0\] _278_/a_27_47# 6.48e-20
C7085 _105_ _118_ 0.00226f
C7086 _258_/a_27_297# _025_ 0.00121f
C7087 clkbuf_0_clk/a_110_47# net19 0.0206f
C7088 _041_ _101_ 0.0098f
C7089 net3 _337_/a_1283_21# 6.01e-19
C7090 _256_/a_373_47# trim_mask\[4\] 2.84e-19
C7091 _078_ _084_ 0.00517f
C7092 _025_ _024_ 6.82e-20
C7093 _306_/a_193_47# _049_ 4.22e-19
C7094 _308_/a_543_47# net14 0.00542f
C7095 _326_/a_1283_21# clknet_2_1__leaf_clk 4.23e-20
C7096 _308_/a_1108_47# _138_/a_27_47# 1.9e-19
C7097 VPWR _323_/a_1283_21# 0.0185f
C7098 _322_/a_639_47# net44 0.00179f
C7099 VPWR _298_/a_78_199# 0.0353f
C7100 _074_ _310_/a_639_47# 0.00204f
C7101 _314_/a_1283_21# net29 0.0368f
C7102 _300_/a_377_297# net2 0.00429f
C7103 _060_ state\[1\] 0.0926f
C7104 output29/a_27_47# _314_/a_27_47# 0.0106f
C7105 _309_/a_193_47# _308_/a_1283_21# 5.28e-20
C7106 _309_/a_27_47# _308_/a_1108_47# 4.8e-19
C7107 _074_ calibrate 0.233f
C7108 _030_ _029_ 3.04e-21
C7109 net4 _090_ 3.3e-20
C7110 net43 _320_/a_27_47# 2.28e-20
C7111 net21 _313_/a_1462_47# 1.36e-19
C7112 _335_/a_543_47# _032_ 0.00157f
C7113 _051_ clknet_2_2__leaf_clk 5.36e-19
C7114 _128_ _338_/a_1602_47# 3.23e-20
C7115 net12 _242_/a_79_21# 0.00775f
C7116 _015_ _243_/a_27_297# 0.00484f
C7117 _325_/a_448_47# _321_/a_193_47# 6.78e-20
C7118 _305_/a_27_47# _305_/a_761_289# -0.0166f
C7119 _299_/a_27_413# _297_/a_47_47# 3.62e-19
C7120 net36 net33 0.157f
C7121 _288_/a_59_75# cal_count\[2\] 8.42e-19
C7122 _325_/a_543_47# _313_/a_27_47# 8.17e-21
C7123 _325_/a_27_47# _313_/a_543_47# 3.71e-21
C7124 _255_/a_27_47# _053_ 0.00554f
C7125 trim_val\[1\] net46 0.031f
C7126 ctlp[3] net16 2.35e-19
C7127 net44 _312_/a_761_289# 0.00347f
C7128 _291_/a_285_47# net47 1.21e-20
C7129 VPWR _341_/a_1108_47# 0.0101f
C7130 clkbuf_0_clk/a_110_47# _001_ 6.44e-21
C7131 net2 _332_/a_448_47# 1.91e-19
C7132 net50 trim_mask\[0\] 0.00851f
C7133 _303_/a_193_47# clknet_2_3__leaf_clk 0.587f
C7134 clknet_2_0__leaf_clk mask\[2\] 8.35e-19
C7135 net13 _320_/a_1217_47# 1.84e-20
C7136 _149_/a_68_297# mask\[4\] 0.0371f
C7137 _230_/a_145_75# _092_ 0.00232f
C7138 _117_ _335_/a_27_47# 0.00205f
C7139 _116_ _335_/a_193_47# 3.56e-20
C7140 _110_ _335_/a_761_289# 1.39e-20
C7141 _305_/a_761_289# net51 4.95e-19
C7142 net43 _307_/a_193_47# 2.76e-19
C7143 _272_/a_81_21# _334_/a_651_413# 5.04e-20
C7144 trim_val\[2\] _334_/a_193_47# 2.37e-19
C7145 net55 _095_ 0.0478f
C7146 _194_/a_113_297# _118_ 3.83e-19
C7147 _100_ _092_ 9.61e-20
C7148 _096_ _099_ 0.28f
C7149 result[7] net15 1.8e-20
C7150 VPWR _308_/a_543_47# 0.0341f
C7151 clk _048_ 0.137f
C7152 _140_/a_68_297# _245_/a_27_297# 7.94e-19
C7153 net15 net30 0.429f
C7154 _336_/a_1283_21# _118_ 1.64e-20
C7155 _336_/a_1108_47# trim_val\[4\] 3.75e-19
C7156 _306_/a_27_47# cal_itt\[3\] 1.58e-19
C7157 _106_ _279_/a_396_47# 0.00425f
C7158 _048_ clone7/a_27_47# 2.01e-20
C7159 clknet_0_clk _119_ 0.0394f
C7160 _038_ _231_/a_161_47# 1.62e-19
C7161 _228_/a_79_21# _054_ 1.26e-20
C7162 _052_ _170_/a_299_297# 0.025f
C7163 _228_/a_297_47# _049_ 0.0486f
C7164 result[5] _086_ 3.98e-19
C7165 net27 _011_ 0.0592f
C7166 net16 _334_/a_193_47# 3.08e-20
C7167 _110_ _332_/a_193_47# 0.00146f
C7168 _042_ _310_/a_761_289# 2.1e-20
C7169 _303_/a_27_47# _303_/a_761_289# -0.0166f
C7170 _169_/a_215_311# _096_ 6.38e-21
C7171 VPWR _320_/a_1270_413# -1.61e-19
C7172 clk trim_mask\[4\] 0.00945f
C7173 _110_ net31 6.29e-20
C7174 _087_ _098_ 0.0462f
C7175 ctlp[0] result[7] 0.144f
C7176 VPWR _339_/a_476_47# 0.0193f
C7177 clknet_2_1__leaf_clk _310_/a_448_47# 0.0289f
C7178 _064_ _336_/a_27_47# 8.59e-21
C7179 _328_/a_1283_21# _267_/a_59_75# 3.41e-19
C7180 VPWR output13/a_27_47# 0.114f
C7181 _048_ net4 0.00405f
C7182 net15 net22 4.98e-20
C7183 _326_/a_27_47# _022_ 6.41e-22
C7184 _078_ _085_ 0.00369f
C7185 _326_/a_1108_47# mask\[6\] 6.58e-20
C7186 VPWR _140_/a_150_297# 0.00142f
C7187 _175_/a_68_297# _055_ 3.39e-19
C7188 _333_/a_193_47# _055_ 1.23e-19
C7189 clknet_2_3__leaf_clk net53 1.23e-20
C7190 net13 _322_/a_27_47# 0.0193f
C7191 _308_/a_543_47# net23 6.34e-19
C7192 _308_/a_448_47# net43 3e-19
C7193 _308_/a_651_413# _005_ 1.23e-20
C7194 net9 _334_/a_761_289# 3.21e-19
C7195 output35/a_27_47# _131_ 4.38e-22
C7196 _258_/a_109_47# trim_mask\[4\] 1.17e-19
C7197 net49 rebuffer2/a_75_212# 0.00489f
C7198 _337_/a_193_47# _034_ 0.0752f
C7199 net4 trim_mask\[4\] 0.0156f
C7200 _112_ _108_ 0.00294f
C7201 net49 _332_/a_1283_21# 1.28e-21
C7202 _112_ _332_/a_543_47# 1.87e-20
C7203 VPWR _307_/a_639_47# 4.04e-19
C7204 trim_mask\[1\] _029_ 5.78e-21
C7205 _338_/a_476_47# _001_ 2.17e-20
C7206 state\[1\] en_co_clk 6.36e-19
C7207 _127_ net37 0.00111f
C7208 trim[0] _112_ 1.79e-20
C7209 _329_/a_805_47# _026_ 3.24e-19
C7210 _329_/a_805_47# VPWR 1.87e-19
C7211 _053_ _336_/a_27_47# 0.00136f
C7212 _256_/a_27_297# trim_val\[4\] 5.6e-20
C7213 trim_mask\[0\] _279_/a_396_47# 0.0296f
C7214 _110_ _113_ 0.255f
C7215 net9 _286_/a_505_21# 2.47e-19
C7216 VPWR trimb[2] 0.252f
C7217 _309_/a_448_47# net14 0.00314f
C7218 _263_/a_297_47# _098_ 1.51e-19
C7219 _313_/a_193_47# _045_ 1.48e-20
C7220 state\[2\] _100_ 0.00152f
C7221 _321_/a_448_47# mask\[3\] 1.66e-20
C7222 cal_itt\[1\] _195_/a_505_21# 0.0052f
C7223 cal_itt\[0\] _195_/a_218_374# 8.73e-20
C7224 _094_ _192_/a_27_47# 3.55e-19
C7225 _129_ _297_/a_285_47# 0.0265f
C7226 _048_ _073_ 7.12e-19
C7227 clknet_2_1__leaf_clk _247_/a_27_297# 0.0724f
C7228 _057_ _056_ 8.97e-20
C7229 _309_/a_193_47# _309_/a_651_413# -0.00701f
C7230 _125_ _131_ 3e-21
C7231 _311_/a_27_47# net26 0.0437f
C7232 net5 output35/a_27_47# 0.00159f
C7233 _042_ _311_/a_1283_21# 7.31e-20
C7234 net2 clknet_2_1__leaf_clk 0.0109f
C7235 _114_ net46 0.0171f
C7236 _322_/a_27_47# _322_/a_193_47# -0.17f
C7237 _309_/a_1283_21# _245_/a_109_297# 7.64e-22
C7238 _309_/a_1108_47# _245_/a_27_297# 3.74e-22
C7239 trim_mask\[0\] _181_/a_150_297# 9.24e-19
C7240 net43 rebuffer6/a_27_47# 9.98e-21
C7241 trim_mask\[3\] trim_mask\[2\] 0.0993f
C7242 _331_/a_27_47# _331_/a_193_47# -0.182f
C7243 _306_/a_448_47# clknet_2_0__leaf_clk 1.99e-19
C7244 calibrate _170_/a_299_297# 0.0408f
C7245 VPWR _303_/a_543_47# 0.0258f
C7246 _110_ net2 1.31e-20
C7247 _269_/a_81_21# trim_val\[1\] 0.0368f
C7248 _078_ _314_/a_543_47# 6.41e-19
C7249 net12 _050_ 0.0242f
C7250 _323_/a_1108_47# net19 0.0132f
C7251 _126_ net37 0.458f
C7252 _239_/a_694_21# calibrate 9.72e-20
C7253 _321_/a_1108_47# mask\[4\] 1.5e-19
C7254 net35 _162_/a_27_47# 6.06e-22
C7255 trim_val\[2\] _334_/a_1462_47# 6.42e-19
C7256 _294_/a_150_297# _125_ 2.38e-20
C7257 _081_ _212_/a_113_297# 1.76e-20
C7258 _306_/a_1217_47# cal_itt\[3\] 1.52e-19
C7259 _266_/a_68_297# clknet_2_3__leaf_clk 3.57e-20
C7260 _036_ _339_/a_476_47# 7.8e-19
C7261 cal_count\[1\] _339_/a_1182_261# 0.00358f
C7262 mask\[3\] _143_/a_68_297# 3.51e-21
C7263 _319_/a_761_289# _120_ 2.43e-20
C7264 _329_/a_27_47# trim_mask\[3\] 0.00556f
C7265 _062_ rebuffer3/a_75_212# 9.39e-20
C7266 _324_/a_27_47# _101_ 2.95e-20
C7267 clk _190_/a_27_47# 1.17e-19
C7268 VPWR _309_/a_448_47# -0.00316f
C7269 _291_/a_35_297# trimb[1] 6.6e-19
C7270 _276_/a_145_75# _110_ 0.00165f
C7271 _276_/a_59_75# _116_ 0.042f
C7272 _326_/a_27_47# _011_ 1.73e-19
C7273 _326_/a_761_289# _086_ 6.54e-20
C7274 net20 net53 3.24e-20
C7275 _328_/a_1108_47# net46 0.0251f
C7276 state\[0\] net55 0.00109f
C7277 net28 result[6] 0.0317f
C7278 _050_ net44 4.63e-19
C7279 _131_ net40 0.0122f
C7280 VPWR _339_/a_1224_47# 8.97e-20
C7281 VPWR _245_/a_373_47# -1.06e-19
C7282 trim[4] net33 3.24e-19
C7283 _104_ _336_/a_639_47# 0.00118f
C7284 _060_ _337_/a_1108_47# 3.21e-21
C7285 _103_ _062_ 2.33e-19
C7286 net54 _337_/a_448_47# 5.27e-21
C7287 _039_ _049_ 1.46e-19
C7288 _324_/a_651_413# net53 6.01e-19
C7289 net16 cal_count\[0\] 0.081f
C7290 trim_val\[3\] net18 0.00706f
C7291 mask\[7\] _158_/a_68_297# 0.0301f
C7292 _065_ _062_ 1.86e-19
C7293 _235_/a_297_47# state\[1\] 4.89e-22
C7294 _094_ clknet_2_0__leaf_clk 0.0325f
C7295 _237_/a_535_374# _090_ 0.00106f
C7296 clknet_2_1__leaf_clk _221_/a_109_297# 0.00422f
C7297 _005_ net43 4.29e-19
C7298 net13 net21 0.0411f
C7299 _238_/a_75_212# calibrate 0.0273f
C7300 _321_/a_27_47# mask\[2\] 8.74e-19
C7301 VPWR _324_/a_639_47# 8.07e-19
C7302 _294_/a_150_297# net40 4.26e-19
C7303 _105_ _062_ 2.74e-19
C7304 calibrate _192_/a_174_21# 4.35e-21
C7305 _050_ _003_ 3.51e-20
C7306 _322_/a_448_47# net53 5.51e-21
C7307 net5 net40 1.96e-19
C7308 _110_ trim_val\[1\] 8.48e-19
C7309 clknet_2_1__leaf_clk net29 0.00238f
C7310 mask\[6\] _247_/a_109_297# 5.16e-21
C7311 _309_/a_639_47# net43 6.04e-19
C7312 _061_ net16 2.82e-19
C7313 _327_/a_1108_47# trim_mask\[0\] 0.00486f
C7314 _327_/a_761_289# _024_ 0.00253f
C7315 _053_ _304_/a_639_47# 8.12e-19
C7316 _089_ net41 4.47e-19
C7317 _195_/a_76_199# _065_ 8.83e-20
C7318 net23 _245_/a_373_47# 0.00101f
C7319 net45 _137_/a_68_297# 0.00161f
C7320 _316_/a_543_47# _095_ 4.5e-19
C7321 _053_ _340_/a_193_47# 1.6e-19
C7322 output11/a_27_47# output12/a_27_47# 4.72e-21
C7323 VPWR _322_/a_1270_413# 7.33e-20
C7324 VPWR _331_/a_1270_413# 6.95e-20
C7325 _314_/a_448_47# _011_ 0.00445f
C7326 net55 _226_/a_27_47# 5.75e-19
C7327 _078_ _311_/a_193_47# 5.67e-20
C7328 _074_ _315_/a_27_47# 0.0275f
C7329 _258_/a_109_297# _058_ 2.93e-19
C7330 _324_/a_193_47# _312_/a_1108_47# 1.89e-19
C7331 _324_/a_761_289# _312_/a_1283_21# 9.96e-21
C7332 VPWR _089_ 0.0737f
C7333 _257_/a_27_297# _025_ 0.0083f
C7334 _331_/a_27_47# _260_/a_93_21# 4.97e-21
C7335 VPWR _218_/a_199_47# 9.64e-20
C7336 net49 _112_ 5.7e-19
C7337 net48 _269_/a_299_297# 1.06e-19
C7338 _272_/a_299_297# net49 9.52e-20
C7339 _008_ net20 7.12e-22
C7340 _245_/a_373_47# net52 0.00168f
C7341 _245_/a_109_297# _016_ 0.00284f
C7342 _008_ net53 0.028f
C7343 VPWR _312_/a_193_47# 0.00679f
C7344 net15 _319_/a_1108_47# 9.63e-19
C7345 net54 clone7/a_27_47# 0.0136f
C7346 _074_ _225_/a_109_297# 0.00107f
C7347 _121_ _095_ 7.97e-19
C7348 output7/a_27_47# net6 3.17e-21
C7349 _308_/a_448_47# _080_ 7.37e-19
C7350 net27 _313_/a_761_289# 2.51e-21
C7351 clknet_2_0__leaf_clk _244_/a_27_297# 0.0417f
C7352 cal_itt\[1\] _305_/a_1108_47# 3.79e-21
C7353 _194_/a_113_297# _062_ 4.43e-19
C7354 output15/a_27_47# net29 8.41e-19
C7355 _237_/a_535_374# _048_ 3.1e-19
C7356 VPWR _275_/a_299_297# 0.0235f
C7357 _336_/a_1283_21# _062_ 3.55e-19
C7358 _237_/a_505_21# net3 0.0158f
C7359 _064_ _136_ 2.37e-19
C7360 _093_ _078_ 4.53e-21
C7361 net43 net21 0.0413f
C7362 _012_ net22 9.79e-21
C7363 net54 net4 1.14e-19
C7364 _313_/a_1108_47# _084_ 1.37e-20
C7365 _059_ _337_/a_193_47# 3.64e-19
C7366 _074_ clknet_2_0__leaf_clk 0.167f
C7367 _337_/a_1108_47# en_co_clk 0.049f
C7368 _303_/a_1283_21# net19 1.08e-19
C7369 ctln[1] clknet_2_0__leaf_clk 4.53e-21
C7370 _033_ _330_/a_27_47# 6.44e-20
C7371 cal _316_/a_193_47# 2.27e-19
C7372 net1 _316_/a_27_47# 3.65e-20
C7373 _015_ _316_/a_1108_47# 3.41e-20
C7374 net3 output41/a_27_47# 9.02e-19
C7375 _254_/a_109_297# net42 5.63e-19
C7376 net8 net46 0.041f
C7377 _341_/a_193_47# _092_ 7.25e-19
C7378 _270_/a_59_75# _029_ 7.15e-20
C7379 _053_ _136_ 0.0545f
C7380 _337_/a_1283_21# _076_ 0.00101f
C7381 _336_/a_193_47# _052_ 1.27e-20
C7382 _263_/a_79_21# _087_ 0.00945f
C7383 _019_ net53 0.00779f
C7384 _110_ _114_ 0.00628f
C7385 _053_ _284_/a_68_297# 0.0136f
C7386 _099_ _098_ 0.0122f
C7387 mask\[6\] _018_ 3.93e-20
C7388 net8 _334_/a_639_47# 7.53e-19
C7389 _325_/a_761_289# net13 0.00324f
C7390 VPWR _291_/a_285_297# 5.5e-20
C7391 VPWR _213_/a_109_297# 8.7e-19
C7392 _088_ clone1/a_27_47# 0.00314f
C7393 _104_ net12 0.034f
C7394 _119_ clknet_2_2__leaf_clk 0.358f
C7395 _190_/a_465_47# clkbuf_2_3__f_clk/a_110_47# 1.07e-20
C7396 _250_/a_373_47# _021_ 0.00113f
C7397 output23/a_27_47# clknet_2_0__leaf_clk 0.00967f
C7398 _312_/a_805_47# net20 4.97e-19
C7399 _237_/a_76_199# _241_/a_297_47# 7.48e-20
C7400 clknet_0_clk _099_ 2.05e-20
C7401 _323_/a_27_47# mask\[5\] 9.28e-19
C7402 _308_/a_1283_21# mask\[1\] 0.00118f
C7403 calibrate _315_/a_805_47# 3.62e-20
C7404 _012_ _315_/a_651_413# 1.08e-20
C7405 _336_/a_1108_47# _335_/a_193_47# 3.03e-19
C7406 net9 _042_ 3.59e-19
C7407 _322_/a_448_47# _019_ 0.00364f
C7408 net24 _146_/a_68_297# 0.00108f
C7409 _212_/a_113_297# net14 0.0087f
C7410 _331_/a_761_289# trim_mask\[4\] 5.6e-19
C7411 _331_/a_448_47# _028_ 0.0145f
C7412 clknet_2_1__leaf_clk mask\[0\] 1.88e-19
C7413 state\[0\] _316_/a_543_47# 1.56e-19
C7414 net33 _108_ 0.34f
C7415 output24/a_27_47# clknet_2_1__leaf_clk 2.58e-19
C7416 _110_ _328_/a_1108_47# 3.3e-20
C7417 _320_/a_639_47# mask\[1\] 7.19e-21
C7418 _002_ _203_/a_59_75# 5.1e-20
C7419 _189_/a_27_47# wire42/a_75_212# 4.96e-20
C7420 trim[0] net33 0.00267f
C7421 _321_/a_651_413# net15 1.36e-20
C7422 net2 _065_ 0.887f
C7423 _336_/a_761_289# _108_ 0.00893f
C7424 output15/a_27_47# ctlp[1] 0.0174f
C7425 _005_ _080_ 0.0683f
C7426 _305_/a_1283_21# _065_ 6.43e-20
C7427 net18 trim_val\[4\] 1.73e-21
C7428 trim_val\[2\] net16 0.111f
C7429 _094_ _337_/a_27_47# 0.222f
C7430 _327_/a_543_47# net18 0.00215f
C7431 _052_ net55 0.0806f
C7432 _097_ _317_/a_193_47# 4.42e-21
C7433 _323_/a_1270_413# mask\[4\] 2.86e-20
C7434 _318_/a_193_47# _318_/a_543_47# -0.0129f
C7435 _218_/a_199_47# _083_ 0.0015f
C7436 _306_/a_27_47# clk 1.37e-20
C7437 comp net34 0.108f
C7438 _019_ _008_ -1.01e-24
C7439 _309_/a_27_47# _007_ 1.26e-19
C7440 _325_/a_761_289# net43 -0.00231f
C7441 _336_/a_805_47# net46 -0.00125f
C7442 _328_/a_639_47# trim_mask\[1\] 6.86e-21
C7443 _264_/a_27_297# net46 4.18e-20
C7444 VPWR _212_/a_113_297# 0.0526f
C7445 VPWR _333_/a_805_47# 4.56e-19
C7446 _068_ _202_/a_382_297# 4e-19
C7447 _081_ _017_ 8.78e-21
C7448 _149_/a_68_297# _311_/a_1108_47# 4.14e-20
C7449 _031_ net33 2.32e-21
C7450 clkbuf_0_clk/a_110_47# _062_ 0.00163f
C7451 VPWR _109_ 0.143f
C7452 _192_/a_174_21# _192_/a_27_47# -5.68e-32
C7453 output29/a_27_47# _078_ 1.41e-19
C7454 cal_itt\[2\] cal_itt\[0\] 0.0273f
C7455 _309_/a_27_47# mask\[3\] 1.75e-19
C7456 _309_/a_193_47# net25 3.78e-20
C7457 _050_ _331_/a_543_47# 0.00129f
C7458 clkbuf_2_1__f_clk/a_110_47# _319_/a_193_47# 0.0204f
C7459 _205_/a_27_47# net53 3.34e-19
C7460 comp _299_/a_298_297# 2.03e-19
C7461 _325_/a_193_47# _101_ 5.62e-19
C7462 _324_/a_1108_47# _152_/a_68_297# 4.78e-20
C7463 net42 _262_/a_27_47# 0.0135f
C7464 mask\[7\] _085_ 2e-19
C7465 _232_/a_32_297# _065_ 0.00109f
C7466 _125_ _122_ 8.39e-20
C7467 _275_/a_299_297# net50 0.00252f
C7468 _275_/a_384_47# trim_mask\[3\] 0.00122f
C7469 VPWR _152_/a_68_297# 0.0251f
C7470 _064_ clknet_0_clk 1.04e-19
C7471 _047_ net37 0.454f
C7472 net15 _316_/a_27_47# 2.99e-20
C7473 clkbuf_0_clk/a_110_47# _195_/a_76_199# 0.011f
C7474 _328_/a_193_47# _328_/a_543_47# -0.0231f
C7475 _328_/a_27_47# _328_/a_1283_21# -9.15e-20
C7476 mask\[6\] _078_ 0.216f
C7477 _337_/a_27_47# _244_/a_27_297# 4.58e-20
C7478 _210_/a_113_297# mask\[0\] 2.22e-19
C7479 _210_/a_199_47# net22 1.55e-19
C7480 net23 _212_/a_113_297# 0.00131f
C7481 _097_ net30 4.53e-21
C7482 _053_ _098_ 4.65e-21
C7483 _328_/a_543_47# net9 0.00272f
C7484 _123_ _065_ 0.0142f
C7485 _033_ _335_/a_27_47# 5.24e-22
C7486 _337_/a_1462_47# _075_ 6.2e-19
C7487 _107_ _242_/a_79_21# 0.0112f
C7488 _270_/a_145_75# _112_ 6.69e-19
C7489 _125_ _299_/a_27_413# 1.04e-19
C7490 net28 _158_/a_68_297# 0.0184f
C7491 _041_ _077_ 5.12e-20
C7492 _071_ net30 1.26e-19
C7493 net9 ctln[3] 0.00737f
C7494 _321_/a_27_47# _074_ 2.72e-20
C7495 VPWR _279_/a_490_47# -8.24e-19
C7496 net12 _228_/a_79_21# 0.00707f
C7497 trim_mask\[4\] _260_/a_250_297# 0.0758f
C7498 _306_/a_27_47# _073_ 2.64e-20
C7499 calibrate net55 0.404f
C7500 _093_ _096_ 0.119f
C7501 net13 mask\[4\] 0.0131f
C7502 VPWR _325_/a_805_47# 3.44e-19
C7503 _317_/a_543_47# _014_ 0.00226f
C7504 _317_/a_1283_21# clknet_2_0__leaf_clk 0.0495f
C7505 _317_/a_761_289# net45 2.73e-19
C7506 _306_/a_543_47# _041_ 1.18e-21
C7507 _103_ _227_/a_209_311# 0.046f
C7508 _232_/a_32_297# _243_/a_109_297# 8.58e-19
C7509 _053_ clknet_0_clk 0.0952f
C7510 _262_/a_27_47# net30 0.00193f
C7511 _092_ net41 5.14e-20
C7512 _322_/a_761_289# mask\[3\] 0.0505f
C7513 VPWR _158_/a_150_297# 2.05e-19
C7514 _325_/a_543_47# net21 0.00162f
C7515 net13 _220_/a_199_47# 2.21e-20
C7516 _315_/a_543_47# net30 4.91e-21
C7517 _333_/a_1283_21# _175_/a_68_297# 1.68e-20
C7518 net15 net44 2.1e-21
C7519 _094_ _337_/a_1217_47# 3.29e-19
C7520 _122_ net40 5.85e-20
C7521 net13 _060_ 0.202f
C7522 mask\[7\] _314_/a_543_47# 0.00299f
C7523 _238_/a_75_212# clknet_2_0__leaf_clk 0.00103f
C7524 _051_ _094_ 9.78e-22
C7525 comp _133_ 5.22e-20
C7526 clknet_2_0__leaf_clk _192_/a_174_21# 8.64e-21
C7527 _110_ net8 5.18e-21
C7528 VPWR _092_ 2.68f
C7529 _257_/a_109_297# _058_ 2.86e-19
C7530 net42 wire42/a_75_212# 0.041f
C7531 net12 _306_/a_805_47# 4.47e-19
C7532 trim_val\[3\] trim_mask\[4\] 3.15e-20
C7533 _320_/a_27_47# _076_ 2.2e-21
C7534 _037_ net40 3.14e-19
C7535 _051_ _088_ 1.53e-19
C7536 _321_/a_193_47# _247_/a_109_297# 1.21e-19
C7537 _322_/a_193_47# mask\[4\] 0.0011f
C7538 _299_/a_27_413# net40 0.00526f
C7539 cal net14 0.0197f
C7540 net49 net33 1.57e-20
C7541 _320_/a_651_413# mask\[2\] 4.21e-20
C7542 _320_/a_1283_21# _017_ 3.61e-20
C7543 trim_val\[2\] _176_/a_27_47# 0.0044f
C7544 _071_ _072_ 0.0341f
C7545 _078_ _315_/a_193_47# 1.25e-19
C7546 net22 _315_/a_543_47# 8.02e-19
C7547 _253_/a_299_297# _310_/a_1108_47# 6.39e-20
C7548 trim[1] _047_ 0.122f
C7549 VPWR _169_/a_109_53# 0.0151f
C7550 _290_/a_207_413# net33 0.00314f
C7551 trim_mask\[1\] _336_/a_543_47# 5.37e-21
C7552 _321_/a_193_47# _146_/a_68_297# 4.27e-20
C7553 _249_/a_27_297# _101_ 0.019f
C7554 _303_/a_651_413# mask\[4\] 4.61e-20
C7555 _040_ _246_/a_109_297# 7.16e-19
C7556 _050_ _260_/a_256_47# 0.00128f
C7557 state\[1\] _049_ 6.95e-20
C7558 _318_/a_1108_47# net45 0.00586f
C7559 mask\[3\] _101_ 0.201f
C7560 trim_mask\[0\] _332_/a_761_289# 0.0255f
C7561 en net3 0.00365f
C7562 _326_/a_448_47# _023_ 0.00445f
C7563 _326_/a_651_413# _102_ 1.19e-19
C7564 _326_/a_1270_413# mask\[7\] 1.46e-19
C7565 net43 mask\[4\] 9.74e-20
C7566 _211_/a_109_297# net30 5.38e-19
C7567 output7/a_27_47# clk 0.00341f
C7568 wire42/a_75_212# net30 1.1e-19
C7569 _340_/a_193_47# _285_/a_113_47# 5.7e-21
C7570 cal net41 0.0709f
C7571 state\[2\] net41 2.15e-19
C7572 _136_ _300_/a_47_47# 0.0118f
C7573 clone1/a_27_47# _170_/a_299_297# 4.68e-19
C7574 _309_/a_27_47# fanout43/a_27_47# 1.41e-19
C7575 _041_ _286_/a_218_374# 9.13e-19
C7576 net47 _124_ 0.0145f
C7577 _286_/a_505_21# _338_/a_1032_413# 0.00227f
C7578 _324_/a_1108_47# mask\[5\] 0.00329f
C7579 VPWR _246_/a_109_297# -2.98e-19
C7580 _200_/a_80_21# _230_/a_59_75# 0.0212f
C7581 _262_/a_27_47# _262_/a_465_47# -1.78e-33
C7582 _051_ _108_ 1.4e-20
C7583 VPWR mask\[5\] 1.39f
C7584 net24 _078_ 0.506f
C7585 mask\[0\] net45 0.203f
C7586 _320_/a_543_47# net15 6.38e-19
C7587 _340_/a_1032_413# net2 1.06e-19
C7588 _063_ _092_ 0.367f
C7589 state\[2\] VPWR 0.575f
C7590 VPWR cal 0.152f
C7591 VPWR _327_/a_639_47# 5.1e-19
C7592 _263_/a_79_21# _099_ 0.0441f
C7593 _079_ _210_/a_199_47# 9.05e-20
C7594 output7/a_27_47# net4 0.0341f
C7595 _317_/a_805_47# state\[1\] 9.25e-20
C7596 _322_/a_1283_21# mask\[5\] 5.3e-21
C7597 output31/a_27_47# _055_ 0.224f
C7598 net13 _222_/a_199_47# 3.31e-21
C7599 _136_ _029_ 0.0046f
C7600 _237_/a_505_21# _120_ 0.00182f
C7601 _232_/a_304_297# net55 4.17e-20
C7602 net9 _131_ 7.01e-21
C7603 state\[2\] _331_/a_1283_21# 6.97e-19
C7604 _325_/a_1270_413# _019_ 8.1e-21
C7605 _327_/a_193_47# _025_ 8.86e-20
C7606 net19 _152_/a_150_297# 1.13e-19
C7607 trim_mask\[2\] _334_/a_1283_21# 4.78e-20
C7608 _104_ _280_/a_75_212# 0.0245f
C7609 _101_ _220_/a_113_297# 1.76e-20
C7610 _050_ _107_ 0.0466f
C7611 clkbuf_0_clk/a_110_47# net2 3.61e-20
C7612 _319_/a_543_47# _049_ 8.73e-19
C7613 net13 en_co_clk 0.0537f
C7614 _324_/a_543_47# net27 2e-19
C7615 mask\[0\] _065_ 6.95e-19
C7616 _319_/a_193_47# net30 9.05e-20
C7617 _110_ _264_/a_27_297# 0.109f
C7618 _305_/a_1283_21# clkbuf_0_clk/a_110_47# 0.00428f
C7619 _305_/a_27_47# clk 0.00415f
C7620 _166_/a_161_47# _050_ 0.0255f
C7621 net23 _246_/a_109_297# 7.55e-20
C7622 _312_/a_1108_47# _045_ 9.55e-21
C7623 VPWR ctln[5] 0.0216f
C7624 trimb[0] net16 1.1e-19
C7625 net34 net46 0.00589f
C7626 VPWR comp 0.189f
C7627 _025_ _058_ 0.00193f
C7628 _104_ _331_/a_543_47# 1.29e-21
C7629 _288_/a_59_75# _297_/a_47_47# 0.00179f
C7630 _331_/a_27_47# _330_/a_27_47# 0.0967f
C7631 _321_/a_193_47# _018_ 0.00522f
C7632 _329_/a_1283_21# _334_/a_27_47# 1.95e-20
C7633 _309_/a_1108_47# mask\[2\] 6.47e-20
C7634 _302_/a_27_297# trim_mask\[1\] 1.57e-21
C7635 _341_/a_193_47# net46 -0.00277f
C7636 _246_/a_109_297# net52 0.00809f
C7637 mask\[0\] _319_/a_27_47# 0.23f
C7638 _305_/a_27_47# net4 3.13e-22
C7639 _040_ _208_/a_218_47# 3.98e-20
C7640 output6/a_27_47# ctln[0] 0.00766f
C7641 _023_ _074_ 0.175f
C7642 _086_ _011_ 0.0968f
C7643 _321_/a_27_47# net26 4.33e-20
C7644 net45 _315_/a_1270_413# -3.58e-20
C7645 _198_/a_27_47# en_co_clk 1.18e-19
C7646 _076_ rebuffer6/a_27_47# 0.0305f
C7647 _321_/a_1283_21# _042_ 0.0066f
C7648 _132_ _131_ 0.0709f
C7649 _079_ _315_/a_543_47# 8.18e-20
C7650 _040_ _017_ 0.0831f
C7651 net44 _311_/a_543_47# 0.00253f
C7652 _306_/a_761_289# rebuffer6/a_27_47# 3.83e-20
C7653 _321_/a_1270_413# clknet_2_1__leaf_clk 6.85e-20
C7654 _093_ _316_/a_761_289# 8.41e-20
C7655 _259_/a_27_297# trim_val\[3\] 7.23e-21
C7656 VPWR _208_/a_218_47# -2.69e-19
C7657 _340_/a_1032_413# _123_ 0.0867f
C7658 net43 _222_/a_199_47# 2.03e-19
C7659 clknet_2_1__leaf_clk _313_/a_1283_21# 0.0609f
C7660 _253_/a_81_21# net29 8.48e-19
C7661 cal_count\[0\] _338_/a_1602_47# 0.0142f
C7662 _286_/a_218_374# net18 7.07e-19
C7663 VPWR _017_ 0.0991f
C7664 _300_/a_285_47# _122_ 9.84e-21
C7665 _294_/a_150_297# _132_ 8.78e-19
C7666 fanout43/a_27_47# _101_ 0.00344f
C7667 net5 _132_ 0.00278f
C7668 net2 _338_/a_476_47# 2.54e-20
C7669 _341_/a_193_47# _300_/a_377_297# 1.22e-20
C7670 _192_/a_505_280# _096_ 3.38e-20
C7671 net43 en_co_clk 1.22e-20
C7672 _335_/a_193_47# net18 1.54e-19
C7673 net27 _101_ 1.61e-19
C7674 _058_ _333_/a_543_47# 0.00144f
C7675 _337_/a_27_47# _192_/a_174_21# 1.43e-21
C7676 _182_/a_27_47# trim_val\[0\] 0.0344f
C7677 cal_itt\[2\] _069_ 1.61e-19
C7678 _058_ _265_/a_384_47# 1.18e-19
C7679 fanout45/a_27_47# _317_/a_193_47# 1.34e-19
C7680 net13 _235_/a_297_47# 0.00116f
C7681 VPWR _226_/a_197_47# -2.82e-19
C7682 trim_mask\[0\] trim_mask\[1\] 0.0496f
C7683 trim_mask\[4\] trim_val\[4\] 0.261f
C7684 _301_/a_47_47# _332_/a_651_413# 5.55e-20
C7685 _211_/a_109_297# _079_ 1.66e-20
C7686 _327_/a_1270_413# clknet_2_2__leaf_clk 2.27e-20
C7687 trim_mask\[2\] _113_ 2.11e-19
C7688 net28 _085_ 0.0147f
C7689 _119_ _330_/a_1283_21# 4.21e-20
C7690 _341_/a_1283_21# _108_ 1.43e-20
C7691 net51 _073_ 2.67e-20
C7692 _101_ rebuffer5/a_161_47# 0.0034f
C7693 _072_ _202_/a_79_21# 0.0362f
C7694 _083_ mask\[5\] 0.00101f
C7695 net43 _306_/a_193_47# 5.95e-20
C7696 _212_/a_199_47# mask\[1\] 4.64e-19
C7697 _329_/a_448_47# net46 2.63e-21
C7698 VPWR _330_/a_651_413# 0.00328f
C7699 net23 _017_ 1.83e-20
C7700 cal_itt\[0\] _067_ 0.689f
C7701 trim_val\[3\] _178_/a_68_297# 0.0333f
C7702 _020_ _312_/a_1108_47# 6.99e-22
C7703 cal_itt\[0\] _070_ 0.00884f
C7704 _323_/a_651_413# _068_ 1.1e-21
C7705 output21/a_27_47# _078_ 1.82e-19
C7706 net12 _250_/a_27_297# 0.0117f
C7707 _337_/a_1108_47# _049_ 0.0107f
C7708 cal_itt\[1\] _304_/a_639_47# 1.4e-19
C7709 _068_ clkbuf_2_3__f_clk/a_110_47# 2.29e-19
C7710 _064_ clknet_2_2__leaf_clk 0.246f
C7711 _104_ _260_/a_256_47# 4.64e-19
C7712 _125_ _297_/a_285_47# 1.08e-20
C7713 _337_/a_543_47# net30 1.27e-19
C7714 _314_/a_1283_21# net14 0.00117f
C7715 trim_mask\[0\] _227_/a_296_53# 4.03e-19
C7716 _306_/a_27_47# _101_ 0.01f
C7717 _341_/a_1462_47# net46 -6.3e-19
C7718 _239_/a_694_21# _051_ 0.018f
C7719 _017_ net52 0.0157f
C7720 mask\[0\] _319_/a_1217_47# 8.79e-19
C7721 _060_ net3 0.0282f
C7722 _147_/a_27_47# _042_ 0.0402f
C7723 output36/a_27_47# net33 0.0323f
C7724 _321_/a_193_47# _078_ 3.45e-20
C7725 _319_/a_1270_413# clknet_2_0__leaf_clk 4.01e-19
C7726 _104_ net19 0.122f
C7727 _081_ clknet_2_1__leaf_clk 1e-19
C7728 _307_/a_761_289# _039_ 0.00152f
C7729 net31 net38 2.61e-20
C7730 mask\[3\] _248_/a_27_297# 0.0102f
C7731 _305_/a_805_47# net44 4.25e-19
C7732 mask\[6\] _313_/a_1108_47# 2.19e-20
C7733 _250_/a_27_297# net44 9.27e-20
C7734 _308_/a_761_289# _074_ 0.00835f
C7735 clknet_2_0__leaf_clk net55 3.53e-19
C7736 _014_ _096_ 7.19e-19
C7737 _053_ clknet_2_2__leaf_clk 0.00227f
C7738 net14 _310_/a_27_47# 0.00725f
C7739 net27 _312_/a_448_47# 5.98e-20
C7740 _233_/a_27_297# net14 0.00997f
C7741 _229_/a_27_297# _228_/a_79_21# 5.4e-20
C7742 _338_/a_476_47# _123_ 9.46e-22
C7743 _104_ trim_mask\[3\] 0.183f
C7744 result[6] _314_/a_193_47# 0.00342f
C7745 net28 _314_/a_543_47# 0.0102f
C7746 _059_ _089_ 0.0142f
C7747 _309_/a_193_47# _310_/a_193_47# 8.2e-21
C7748 _309_/a_761_289# _310_/a_27_47# 1.76e-19
C7749 _093_ clknet_0_clk 3.8e-20
C7750 mask\[7\] output29/a_27_47# 1.67e-19
C7751 _043_ _150_/a_27_47# 0.013f
C7752 _326_/a_193_47# net43 0.00792f
C7753 net10 _057_ 8.16e-19
C7754 _327_/a_1108_47# _109_ 2.67e-20
C7755 _103_ _100_ 3.7e-20
C7756 _301_/a_285_47# _135_ 5.24e-19
C7757 net12 _009_ 8.32e-19
C7758 _257_/a_27_297# _335_/a_27_47# 2.3e-20
C7759 _323_/a_27_47# clknet_2_1__leaf_clk 0.00941f
C7760 _297_/a_285_47# net40 0.00447f
C7761 VPWR _161_/a_150_297# 3.2e-19
C7762 _326_/a_639_47# net14 0.00129f
C7763 _057_ clknet_2_2__leaf_clk 2.3e-19
C7764 _104_ _107_ 0.0234f
C7765 VPWR _314_/a_1283_21# 0.0622f
C7766 _335_/a_1462_47# net18 3.94e-19
C7767 _332_/a_1283_21# clknet_2_3__leaf_clk 1.26e-21
C7768 clk _318_/a_193_47# 0.546f
C7769 _074_ _140_/a_68_297# 1.04e-20
C7770 _233_/a_27_297# net41 2.45e-20
C7771 _111_ clknet_2_3__leaf_clk 2.64e-20
C7772 net12 _318_/a_27_47# 8.01e-19
C7773 _000_ _076_ 1.78e-20
C7774 _336_/a_27_47# _336_/a_543_47# -0.00639f
C7775 _336_/a_193_47# _336_/a_761_289# -0.0118f
C7776 mask\[7\] mask\[6\] 0.224f
C7777 trim_mask\[2\] trim_val\[1\] 1.73e-20
C7778 _023_ net26 0.0652f
C7779 net9 _340_/a_956_413# 3.42e-19
C7780 _319_/a_27_47# _319_/a_448_47# -0.00642f
C7781 VPWR _310_/a_27_47# 0.0742f
C7782 net44 _009_ 0.00443f
C7783 VPWR _233_/a_27_297# 0.0532f
C7784 ctlp[5] net19 0.0054f
C7785 _276_/a_59_75# net18 4.1e-19
C7786 _026_ net46 0.00493f
C7787 _339_/a_381_47# cal_count\[0\] 0.0167f
C7788 VPWR net46 2.36f
C7789 _255_/a_27_47# _106_ 5.59e-19
C7790 net4 _318_/a_193_47# 1.57e-19
C7791 _243_/a_109_297# _100_ 1.05e-19
C7792 _243_/a_27_297# _096_ 0.00863f
C7793 _089_ _075_ 5.41e-22
C7794 _034_ _092_ 0.00377f
C7795 _317_/a_193_47# _316_/a_651_413# 5.3e-20
C7796 clk _317_/a_639_47# 5.58e-19
C7797 _317_/a_448_47# _316_/a_761_289# 1.99e-20
C7798 _317_/a_1283_21# _316_/a_1283_21# 1.13e-19
C7799 net43 _314_/a_651_413# 0.00166f
C7800 _290_/a_207_413# output40/a_27_47# 9.59e-19
C7801 net2 _339_/a_1182_261# 3.73e-21
C7802 VPWR _195_/a_439_47# 8.01e-19
C7803 cal_itt\[0\] _338_/a_27_47# 0.00494f
C7804 clknet_2_2__leaf_clk _330_/a_448_47# 0.0254f
C7805 VPWR _326_/a_639_47# 0.00132f
C7806 VPWR _334_/a_639_47# 0.00447f
C7807 _123_ _298_/a_292_297# 0.0028f
C7808 _104_ _279_/a_27_47# 1.94e-19
C7809 _327_/a_761_289# _058_ 0.0126f
C7810 net3 en_co_clk 0.0269f
C7811 _249_/a_109_47# mask\[4\] 8.82e-19
C7812 _237_/a_505_21# clkbuf_2_0__f_clk/a_110_47# 0.00244f
C7813 _097_ _316_/a_27_47# 0.00526f
C7814 _015_ _092_ 4.53e-21
C7815 mask\[1\] _246_/a_109_47# 2.54e-19
C7816 _311_/a_27_47# net53 0.0225f
C7817 net43 _310_/a_543_47# 0.00254f
C7818 _325_/a_1283_21# net27 6.09e-20
C7819 mask\[0\] _282_/a_68_297# 3.54e-19
C7820 _273_/a_59_75# trim_val\[2\] 6.49e-19
C7821 _324_/a_543_47# _311_/a_1283_21# 0.00122f
C7822 _135_ clknet_2_3__leaf_clk 0.194f
C7823 VPWR _300_/a_377_297# 3.22e-19
C7824 _087_ _088_ 4.44e-20
C7825 _104_ _181_/a_68_297# 2.89e-19
C7826 VPWR _335_/a_651_413# 0.00243f
C7827 _323_/a_543_47# net26 8.13e-19
C7828 _323_/a_651_413# _042_ 0.0262f
C7829 cal_count\[1\] net37 6.29e-19
C7830 _167_/a_161_47# state\[1\] 0.0826f
C7831 VPWR _311_/a_761_289# 0.0102f
C7832 trim_mask\[0\] _255_/a_27_47# 0.0762f
C7833 clone1/a_27_47# net55 0.0321f
C7834 _015_ _169_/a_109_53# 0.00193f
C7835 _305_/a_193_47# _198_/a_27_47# 6.08e-20
C7836 _273_/a_59_75# net16 3.67e-19
C7837 net52 _310_/a_27_47# 5.43e-22
C7838 _240_/a_109_297# _049_ 5.97e-22
C7839 _119_ _108_ 0.00681f
C7840 fanout46/a_27_47# _280_/a_75_212# 0.0197f
C7841 net46 _063_ 1.01e-21
C7842 trim_val\[3\] _334_/a_27_47# 9.05e-23
C7843 VPWR _332_/a_448_47# 6.39e-19
C7844 net9 _122_ 0.0809f
C7845 _071_ net44 2.38e-20
C7846 trim_mask\[0\] _270_/a_59_75# 2.23e-19
C7847 calibrate valid 0.00353f
C7848 net12 _318_/a_1217_47# 9.9e-20
C7849 _304_/a_27_47# _067_ 1.01e-19
C7850 net43 _039_ 0.0278f
C7851 clknet_0_clk _171_/a_27_47# 0.00186f
C7852 _336_/a_1283_21# _264_/a_27_297# 1.04e-19
C7853 _336_/a_27_47# _106_ 0.0015f
C7854 trim_mask\[2\] _114_ 0.154f
C7855 net9 _037_ 0.11f
C7856 _281_/a_253_47# _092_ 0.00833f
C7857 _339_/a_1182_261# _123_ 0.0138f
C7858 _107_ _228_/a_79_21# 0.00492f
C7859 _249_/a_109_47# _020_ 6.05e-20
C7860 net43 _305_/a_193_47# 0.612f
C7861 net47 cal_count\[2\] 8.34e-19
C7862 VPWR _310_/a_1217_47# 5.52e-20
C7863 trim[2] _055_ 1.84e-20
C7864 _041_ _072_ 5.23e-20
C7865 input1/a_75_212# cal 0.0181f
C7866 _015_ state\[2\] 8.91e-20
C7867 _008_ _311_/a_27_47# 0.147f
C7868 _322_/a_651_413# _074_ 0.00182f
C7869 _014_ _316_/a_761_289# 0.00576f
C7870 net45 _316_/a_193_47# 0.00726f
C7871 clknet_2_0__leaf_clk _316_/a_543_47# 2.38e-19
C7872 _337_/a_193_47# _096_ 6.48e-19
C7873 _337_/a_27_47# net55 2.11e-19
C7874 _235_/a_297_47# net3 0.0409f
C7875 VPWR _269_/a_81_21# 0.0649f
C7876 cal_itt\[0\] _341_/a_543_47# 5.19e-21
C7877 rstn net6 0.00668f
C7878 clknet_2_2__leaf_clk _027_ 0.0294f
C7879 clknet_2_1__leaf_clk net14 0.0168f
C7880 fanout44/a_27_47# en_co_clk 1.91e-21
C7881 _307_/a_27_47# net30 1.97e-19
C7882 _122_ _132_ 7.95e-21
C7883 _104_ _118_ 0.00748f
C7884 _309_/a_761_289# clknet_2_1__leaf_clk 9.01e-21
C7885 _328_/a_1108_47# trim_mask\[2\] 7.08e-20
C7886 _218_/a_113_297# _074_ 1.16e-20
C7887 _081_ net45 6.44e-20
C7888 _074_ _312_/a_27_47# 7.4e-19
C7889 _028_ _052_ 0.207f
C7890 _306_/a_1283_21# _050_ 5.67e-21
C7891 _311_/a_1217_47# net53 5.17e-20
C7892 trim_mask\[0\] _336_/a_27_47# 8.59e-20
C7893 _000_ _068_ 0.0121f
C7894 _299_/a_27_413# _132_ 0.0119f
C7895 _226_/a_27_47# _095_ 3.66e-19
C7896 _115_ _114_ 0.139f
C7897 _101_ net51 0.247f
C7898 clknet_2_1__leaf_clk _040_ 0.00956f
C7899 clknet_0_clk _192_/a_505_280# 0.0117f
C7900 _175_/a_150_297# rebuffer1/a_75_212# 1e-19
C7901 cal_itt\[1\] clknet_0_clk 0.0151f
C7902 _121_ clknet_2_0__leaf_clk 0.0275f
C7903 _161_/a_68_297# trim_val\[0\] 0.0576f
C7904 _333_/a_761_289# rebuffer1/a_75_212# 2.09e-20
C7905 _324_/a_193_47# _042_ 8.79e-20
C7906 _333_/a_27_47# _332_/a_193_47# 7.12e-22
C7907 _069_ _067_ 0.0456f
C7908 _307_/a_27_47# net22 0.175f
C7909 net30 net18 5.08e-20
C7910 VPWR _305_/a_639_47# 3.35e-19
C7911 _069_ _070_ 0.0359f
C7912 _127_ _129_ 1.48e-19
C7913 output35/a_27_47# net35 0.0704f
C7914 net50 net46 0.0769f
C7915 output31/a_27_47# _333_/a_1283_21# 0.00807f
C7916 net31 _333_/a_27_47# 1.1e-20
C7917 _265_/a_81_21# _332_/a_27_47# 3.01e-20
C7918 _051_ _336_/a_193_47# 0.00327f
C7919 _324_/a_1108_47# clknet_2_1__leaf_clk 0.00114f
C7920 _329_/a_1283_21# net9 3.47e-19
C7921 _050_ _062_ 0.473f
C7922 output34/a_27_47# _334_/a_193_47# 2.12e-19
C7923 net52 _310_/a_1217_47# 9.61e-21
C7924 output22/a_27_47# output24/a_27_47# 9.71e-21
C7925 _335_/a_448_47# clknet_2_2__leaf_clk 2.28e-19
C7926 input2/a_27_47# comp 0.0246f
C7927 _302_/a_109_47# _066_ 3.82e-20
C7928 calibrate _263_/a_382_297# 8.7e-21
C7929 VPWR clknet_2_1__leaf_clk 3.86f
C7930 _322_/a_27_47# _042_ 4.43e-19
C7931 _246_/a_27_297# mask\[2\] 0.0277f
C7932 _304_/a_193_47# _136_ 0.00208f
C7933 _110_ _026_ 4.25e-20
C7934 _333_/a_448_47# net46 0.0178f
C7935 _110_ VPWR 2.61f
C7936 net8 _179_/a_27_47# 0.00169f
C7937 _322_/a_1283_21# clknet_2_1__leaf_clk 5.83e-20
C7938 _323_/a_1108_47# _150_/a_27_47# 2.94e-19
C7939 _304_/a_1217_47# _067_ 1.37e-19
C7940 mask\[3\] _077_ 6.46e-21
C7941 _304_/a_193_47# _284_/a_68_297# 7.13e-21
C7942 _083_ _311_/a_761_289# 1.99e-20
C7943 _303_/a_761_289# net26 0.00133f
C7944 _059_ _092_ 0.289f
C7945 _332_/a_1108_47# clknet_2_2__leaf_clk 2.43e-21
C7946 result[1] net43 1.33e-19
C7947 mask\[1\] net15 0.00484f
C7948 _304_/a_543_47# net47 7.42e-20
C7949 cal_itt\[0\] clknet_2_3__leaf_clk 0.042f
C7950 _029_ clknet_2_2__leaf_clk 0.0802f
C7951 _126_ _129_ 0.0109f
C7952 _113_ _333_/a_27_47# 0.0141f
C7953 net43 _251_/a_27_297# 1.31e-19
C7954 net13 _049_ 0.127f
C7955 net43 _250_/a_109_47# 1.33e-20
C7956 ctln[7] _318_/a_27_47# 2.13e-19
C7957 net13 _318_/a_761_289# 0.00583f
C7958 _308_/a_1283_21# mask\[0\] 0.0103f
C7959 _308_/a_543_47# _078_ 0.00147f
C7960 _340_/a_27_47# _340_/a_1032_413# -0.00561f
C7961 _340_/a_193_47# _340_/a_1182_261# -2.22e-21
C7962 net50 _335_/a_651_413# 0.0012f
C7963 trim_val\[3\] _335_/a_639_47# 2.33e-20
C7964 net44 _319_/a_193_47# 4.35e-20
C7965 _308_/a_27_47# net24 8.97e-21
C7966 _308_/a_193_47# clknet_2_0__leaf_clk 0.00256f
C7967 _210_/a_113_297# net14 0.00505f
C7968 _299_/a_215_297# cal_count\[2\] 0.0799f
C7969 _281_/a_103_199# en_co_clk 0.0689f
C7970 net23 clknet_2_1__leaf_clk 0.00695f
C7971 _317_/a_651_413# net14 2.17e-19
C7972 calibrate _028_ 6.33e-20
C7973 net45 _316_/a_1462_47# -9.14e-19
C7974 _341_/a_193_47# _065_ 0.0116f
C7975 trim_val\[4\] net40 1.61e-20
C7976 _250_/a_109_297# _101_ 0.00127f
C7977 _306_/a_1108_47# _092_ 1.92e-19
C7978 _051_ net55 0.121f
C7979 VPWR output15/a_27_47# 0.0138f
C7980 _313_/a_27_47# _313_/a_761_289# -0.0166f
C7981 cal_itt\[0\] _303_/a_193_47# 1.47e-19
C7982 _162_/a_27_47# _047_ 0.00941f
C7983 _288_/a_59_75# _125_ 0.013f
C7984 _126_ _339_/a_1032_413# 1.28e-21
C7985 _320_/a_448_47# clknet_2_0__leaf_clk 0.00139f
C7986 _320_/a_1283_21# net45 4.09e-19
C7987 net39 net16 0.0166f
C7988 net9 _339_/a_562_413# 4.34e-19
C7989 trim_mask\[3\] fanout46/a_27_47# 0.0016f
C7990 net46 _279_/a_396_47# 7.7e-19
C7991 clknet_2_1__leaf_clk net52 0.743f
C7992 net28 mask\[6\] 0.238f
C7993 net47 _035_ 0.144f
C7994 _287_/a_75_212# _338_/a_652_21# 7.07e-19
C7995 _078_ _140_/a_150_297# 1.95e-19
C7996 VPWR _239_/a_474_297# -0.0187f
C7997 net35 net40 0.0858f
C7998 _064_ _278_/a_27_47# 0.00201f
C7999 _331_/a_193_47# _049_ 1.54e-19
C8000 _327_/a_1283_21# _267_/a_59_75# 0.0141f
C8001 _046_ net29 0.00403f
C8002 net4 _336_/a_448_47# 2.01e-20
C8003 _075_ _092_ 0.0268f
C8004 _324_/a_448_47# mask\[6\] 2.48e-21
C8005 net27 _156_/a_27_47# 3.71e-20
C8006 _324_/a_543_47# _021_ 4.34e-19
C8007 _110_ _063_ 6.44e-20
C8008 _321_/a_1283_21# _143_/a_68_297# 0.00127f
C8009 fanout46/a_27_47# _107_ 1.45e-20
C8010 _326_/a_1283_21# net25 2.65e-21
C8011 net8 trim_mask\[2\] 0.0279f
C8012 net44 _202_/a_79_21# 0.00333f
C8013 net12 _206_/a_27_93# 1.95e-19
C8014 _320_/a_1283_21# _065_ 0.00212f
C8015 _307_/a_1217_47# net22 1.27e-19
C8016 _064_ _330_/a_1283_21# 1.96e-19
C8017 _104_ _330_/a_761_289# 3.01e-20
C8018 state\[2\] _059_ 3.46e-20
C8019 trim_val\[0\] _332_/a_1108_47# 9.18e-19
C8020 VPWR _210_/a_113_297# 0.0641f
C8021 _307_/a_1108_47# net45 4.94e-19
C8022 _189_/a_27_47# _048_ 0.0101f
C8023 _239_/a_694_21# _087_ 0.0132f
C8024 _302_/a_27_297# _136_ 0.0148f
C8025 _307_/a_27_47# _079_ 2.27e-19
C8026 VPWR _317_/a_651_413# -0.00864f
C8027 _032_ clknet_2_2__leaf_clk 0.0022f
C8028 result[0] net45 3.23e-19
C8029 _315_/a_761_289# net14 0.0127f
C8030 net43 _049_ 0.006f
C8031 _302_/a_27_297# _284_/a_68_297# 5.22e-19
C8032 _251_/a_373_47# _046_ 2.01e-19
C8033 mask\[6\] _159_/a_27_47# 2.6e-19
C8034 _298_/a_215_47# _131_ 0.00144f
C8035 _094_ _099_ 5.11e-20
C8036 _288_/a_59_75# net40 0.00443f
C8037 _042_ net21 4.64e-20
C8038 output19/a_27_47# ctlp[5] 0.0188f
C8039 _088_ _099_ -1.01e-24
C8040 net44 _206_/a_27_93# 2.28e-19
C8041 _218_/a_113_297# net26 0.041f
C8042 output15/a_27_47# net52 1.33e-21
C8043 net14 output6/a_27_47# 0.0251f
C8044 _032_ net11 1.11e-19
C8045 _000_ _042_ 1.3e-20
C8046 _269_/a_81_21# _333_/a_448_47# 8.84e-19
C8047 trim_val\[1\] _333_/a_27_47# 0.00797f
C8048 _134_ _131_ 0.098f
C8049 VPWR _192_/a_476_47# -4.49e-19
C8050 _341_/a_193_47# _304_/a_761_289# 1.36e-20
C8051 _341_/a_27_47# _304_/a_543_47# 8.14e-19
C8052 net15 _281_/a_337_297# 9.27e-19
C8053 _191_/a_27_297# net30 0.00331f
C8054 _340_/a_1602_47# net47 5.68e-20
C8055 _037_ _304_/a_1283_21# 1.58e-20
C8056 _091_ net4 0.0128f
C8057 _315_/a_27_47# valid 0.0101f
C8058 _083_ clknet_2_1__leaf_clk 0.0112f
C8059 _108_ _279_/a_206_47# 0.0109f
C8060 _259_/a_109_297# _335_/a_27_47# 8.28e-19
C8061 _259_/a_27_297# _335_/a_193_47# 3.27e-19
C8062 _030_ _109_ -1.01e-24
C8063 net8 _115_ 2.98e-19
C8064 _130_ _131_ 0.152f
C8065 en_co_clk _120_ 0.129f
C8066 _007_ _310_/a_1108_47# 9.3e-21
C8067 output26/a_27_47# _310_/a_27_47# 0.0131f
C8068 net45 net14 0.0278f
C8069 _309_/a_448_47# _078_ 3.69e-19
C8070 clk _033_ 2.05e-20
C8071 _116_ net19 0.00268f
C8072 _323_/a_27_47# _043_ 3.7e-19
C8073 trimb[1] net33 6.99e-19
C8074 _337_/a_27_47# _121_ 0.0509f
C8075 VPWR _315_/a_761_289# 0.0181f
C8076 _021_ _101_ 4.46e-20
C8077 _309_/a_543_47# net24 0.0302f
C8078 _068_ _190_/a_215_47# 0.00289f
C8079 _337_/a_543_47# net44 1.27e-19
C8080 net5 _134_ 0.00203f
C8081 cal_itt\[0\] _303_/a_1462_47# 5.1e-19
C8082 _309_/a_761_289# net45 1.46e-19
C8083 _336_/a_651_413# clkbuf_2_2__f_clk/a_110_47# 0.00129f
C8084 _182_/a_27_47# _108_ 0.00233f
C8085 _304_/a_193_47# clknet_0_clk 5.02e-20
C8086 _233_/a_27_297# input1/a_75_212# 3.78e-19
C8087 _181_/a_68_297# fanout46/a_27_47# 0.00121f
C8088 net25 _310_/a_448_47# 4.37e-20
C8089 mask\[3\] _310_/a_1108_47# 0.00101f
C8090 _082_ _310_/a_543_47# 9.92e-20
C8091 VPWR _318_/a_805_47# 5.1e-19
C8092 net24 _245_/a_27_297# 0.00126f
C8093 trim_mask\[0\] _136_ 0.00162f
C8094 _200_/a_80_21# net19 0.00424f
C8095 _116_ trim_mask\[3\] 6.05e-19
C8096 _110_ net50 0.0487f
C8097 _117_ trim_val\[3\] 0.00648f
C8098 _327_/a_1108_47# net46 0.0155f
C8099 en_co_clk _076_ 0.129f
C8100 _294_/a_150_297# _130_ 9.54e-19
C8101 _104_ _062_ 4.39e-20
C8102 _035_ _338_/a_562_413# 3.7e-19
C8103 _077_ rebuffer5/a_161_47# 0.0119f
C8104 net13 state\[1\] 0.144f
C8105 ctlp[1] _046_ 0.00205f
C8106 net5 _130_ 2.21e-19
C8107 VPWR output6/a_27_47# 0.0383f
C8108 _260_/a_93_21# _049_ 0.0353f
C8109 _048_ _227_/a_109_93# 0.0208f
C8110 _040_ net45 0.0264f
C8111 net45 net41 0.413f
C8112 clknet_2_0__leaf_clk valid 0.00553f
C8113 net4 _033_ 0.0333f
C8114 net32 _055_ 0.0149f
C8115 result[1] _080_ 8.38e-19
C8116 _090_ net30 9.79e-21
C8117 output12/a_27_47# net12 0.0445f
C8118 _328_/a_805_47# VPWR 2.71e-19
C8119 net33 trimb[4] 3.24e-19
C8120 _254_/a_109_297# _107_ 6.64e-19
C8121 calibrate _095_ 0.00101f
C8122 _200_/a_80_21# _107_ 9.99e-19
C8123 trim_mask\[4\] _227_/a_109_93# 3.9e-21
C8124 _307_/a_639_47# _004_ 2.31e-19
C8125 _306_/a_193_47# _076_ 0.0151f
C8126 VPWR net45 2.99f
C8127 cal_itt\[0\] _199_/a_109_297# 4.74e-19
C8128 VPWR rebuffer3/a_75_212# 0.0512f
C8129 _328_/a_761_289# _025_ 1.82e-19
C8130 _040_ _065_ 8.69e-19
C8131 _304_/a_27_47# clknet_2_3__leaf_clk 0.236f
C8132 _322_/a_1270_413# _078_ 1.91e-19
C8133 mask\[4\] _068_ 3.07e-20
C8134 clkbuf_2_1__f_clk/a_110_47# _283_/a_75_212# 2.04e-21
C8135 clk rstn 0.0354f
C8136 net45 _331_/a_1283_21# 0.0601f
C8137 _326_/a_193_47# result[5] 7.03e-19
C8138 _326_/a_543_47# net27 5.3e-20
C8139 net42 _048_ 0.454f
C8140 _217_/a_109_297# clknet_2_1__leaf_clk 8.92e-19
C8141 _066_ net18 0.0344f
C8142 VPWR _103_ 0.0244f
C8143 _325_/a_1108_47# _250_/a_27_297# 8.86e-20
C8144 _050_ _232_/a_32_297# 6.01e-21
C8145 net43 _201_/a_113_47# 3.14e-20
C8146 _208_/a_505_21# rebuffer4/a_27_47# 0.00391f
C8147 _321_/a_1108_47# _320_/a_193_47# 4.8e-21
C8148 net47 _041_ 0.611f
C8149 clknet_2_1__leaf_clk _155_/a_150_297# 0.00148f
C8150 _337_/a_193_47# clknet_0_clk 0.0128f
C8151 net48 _333_/a_193_47# 4.16e-21
C8152 net47 _338_/a_1182_261# 0.0231f
C8153 VPWR _065_ 2.78f
C8154 _338_/a_27_47# _338_/a_193_47# -0.247f
C8155 _304_/a_651_413# net18 9.07e-20
C8156 trim_mask\[1\] _109_ 1.61e-20
C8157 _325_/a_448_47# clknet_2_1__leaf_clk 0.00239f
C8158 mask\[3\] clkbuf_2_1__f_clk/a_110_47# 8.09e-21
C8159 rstn net4 0.00228f
C8160 _104_ _335_/a_761_289# 0.00234f
C8161 _064_ _335_/a_1283_21# 0.00209f
C8162 _322_/a_1283_21# _065_ 0.00339f
C8163 _340_/a_381_47# _037_ 0.00852f
C8164 _193_/a_109_297# net46 1.51e-19
C8165 _053_ _088_ 0.00465f
C8166 net23 net45 0.0169f
C8167 VPWR _105_ 0.0103f
C8168 _110_ _279_/a_396_47# 0.00346f
C8169 net16 _333_/a_543_47# 0.0106f
C8170 result[4] _310_/a_1108_47# 2.85e-19
C8171 _102_ _023_ 2.21e-19
C8172 trim_val\[3\] net9 4.6e-19
C8173 net16 _265_/a_384_47# 8.6e-20
C8174 mask\[4\] _311_/a_448_47# 0.0249f
C8175 VPWR _319_/a_27_47# 0.065f
C8176 _048_ _054_ 1.46e-19
C8177 net12 _041_ 0.00956f
C8178 output14/a_27_47# ctlp[0] 0.0106f
C8179 trim[4] _161_/a_68_297# 0.00111f
C8180 _048_ net30 0.468f
C8181 net35 _332_/a_1270_413# 8.41e-20
C8182 _058_ _332_/a_805_47# 4.09e-19
C8183 _050_ _227_/a_209_311# 0.00104f
C8184 _064_ _108_ 0.06f
C8185 _189_/a_408_47# _092_ 0.00778f
C8186 clknet_0_clk _106_ 5.55e-20
C8187 net3 _049_ 0.0661f
C8188 VPWR _243_/a_109_297# -0.0174f
C8189 _071_ net19 4.17e-19
C8190 _320_/a_27_47# _143_/a_68_297# 8.61e-19
C8191 net45 net52 0.356f
C8192 clknet_2_0__leaf_clk _016_ 0.0814f
C8193 _328_/a_1108_47# _333_/a_27_47# 1.39e-19
C8194 _155_/a_68_297# _009_ 2.08e-21
C8195 _063_ rebuffer3/a_75_212# 6.07e-20
C8196 trim_mask\[4\] _054_ 1.48e-20
C8197 _069_ clknet_2_3__leaf_clk 4.01e-20
C8198 _340_/a_193_47# _339_/a_476_47# 5.41e-19
C8199 _340_/a_1182_261# _339_/a_27_47# 2.07e-19
C8200 _340_/a_476_47# _339_/a_193_47# 3.29e-21
C8201 _168_/a_27_413# _048_ 3.58e-20
C8202 trim_mask\[4\] net30 1.57e-19
C8203 _262_/a_27_47# net19 0.00233f
C8204 clk _316_/a_1270_413# 2.55e-20
C8205 _136_ _298_/a_78_199# 0.00209f
C8206 net25 net29 7.99e-20
C8207 _041_ net44 0.0236f
C8208 _179_/a_27_47# net34 0.013f
C8209 output34/a_27_47# trim_val\[2\] 0.0717f
C8210 net52 _065_ 0.00701f
C8211 _053_ _108_ 0.00353f
C8212 _330_/a_543_47# net46 -9.76e-19
C8213 _330_/a_1283_21# _027_ 0.0413f
C8214 _164_/a_161_47# net45 6.11e-19
C8215 _065_ _063_ 4.66e-19
C8216 cal_count\[1\] cal_count\[2\] 4.34e-19
C8217 trim_mask\[0\] _098_ 0.00401f
C8218 _336_/a_193_47# _119_ 0.00802f
C8219 _168_/a_27_413# trim_mask\[4\] 0.0309f
C8220 net43 _319_/a_543_47# -5.34e-19
C8221 net23 _319_/a_27_47# 6.85e-20
C8222 _071_ _107_ 2.52e-19
C8223 VPWR _194_/a_113_297# 0.0466f
C8224 _323_/a_448_47# net47 1.27e-21
C8225 VPWR _336_/a_1283_21# 0.0254f
C8226 _328_/a_639_47# clknet_2_2__leaf_clk 5.75e-19
C8227 VPWR _304_/a_761_289# 0.00256f
C8228 _340_/a_1032_413# _133_ 0.0121f
C8229 _105_ _063_ 0.127f
C8230 _107_ _262_/a_27_47# 0.00775f
C8231 _340_/a_476_47# clknet_2_3__leaf_clk 6.56e-19
C8232 _074_ _084_ 0.0193f
C8233 _341_/a_1108_47# _136_ 0.00705f
C8234 _341_/a_193_47# _038_ -0.0105f
C8235 _057_ _108_ 2.53e-21
C8236 trim_mask\[0\] clknet_0_clk 0.00637f
C8237 _042_ _045_ 1.83e-21
C8238 output21/a_27_47# net28 0.00665f
C8239 state\[0\] calibrate 0.00673f
C8240 _326_/a_1283_21# net15 9.71e-21
C8241 _042_ _249_/a_109_297# 0.0425f
C8242 _325_/a_761_289# _022_ 7.67e-19
C8243 _338_/a_1032_413# _122_ 0.0012f
C8244 output26/a_27_47# clknet_2_1__leaf_clk 0.0227f
C8245 _319_/a_27_47# net52 5.23e-20
C8246 _092_ _170_/a_81_21# 6.21e-19
C8247 _326_/a_193_47# _326_/a_761_289# 7.11e-33
C8248 _334_/a_27_47# _334_/a_543_47# -0.00787f
C8249 net47 net18 0.283f
C8250 net47 _338_/a_1296_47# 0.00113f
C8251 _338_/a_193_47# _338_/a_586_47# -7.91e-19
C8252 _314_/a_193_47# _314_/a_543_47# 3.55e-33
C8253 en_co_clk _068_ 0.0292f
C8254 net13 _321_/a_1108_47# 0.00106f
C8255 net42 _190_/a_27_47# 1.25e-19
C8256 _239_/a_694_21# _099_ 1.37e-20
C8257 net47 _129_ 1.66e-19
C8258 net13 _337_/a_1108_47# 0.00163f
C8259 _187_/a_27_413# net40 0.00448f
C8260 _321_/a_27_47# net53 2.51e-22
C8261 _110_ _327_/a_1108_47# 0.00254f
C8262 wire42/a_75_212# net19 4.1e-22
C8263 net13 _167_/a_161_47# 1.79e-19
C8264 _332_/a_27_47# net40 0.0196f
C8265 _336_/a_761_289# _266_/a_68_297# 4.53e-19
C8266 fanout44/a_27_47# _049_ 0.0028f
C8267 _268_/a_75_212# net40 0.0221f
C8268 net50 rebuffer3/a_75_212# 0.00292f
C8269 _042_ mask\[4\] 0.0476f
C8270 VPWR _319_/a_1217_47# 4.45e-20
C8271 fanout43/a_27_47# clkbuf_2_1__f_clk/a_110_47# 1.43e-20
C8272 VPWR _043_ 0.26f
C8273 clknet_2_1__leaf_clk _141_/a_27_47# 4.73e-19
C8274 _031_ _057_ 6.44e-20
C8275 trim_mask\[2\] net34 2.69e-19
C8276 _168_/a_207_413# _050_ 0.0609f
C8277 VPWR _321_/a_761_289# 0.0139f
C8278 net4 clkbuf_2_3__f_clk/a_110_47# 0.0209f
C8279 _253_/a_81_21# net14 0.00317f
C8280 _323_/a_448_47# net44 0.00175f
C8281 trim[4] _332_/a_1108_47# 5.6e-19
C8282 _283_/a_75_212# net30 0.0273f
C8283 _050_ mask\[0\] 9.79e-21
C8284 net47 _339_/a_1032_413# 7.04e-19
C8285 _212_/a_113_297# _078_ 0.0185f
C8286 _336_/a_1283_21# _063_ 4.46e-19
C8287 calibrate _226_/a_27_47# 8.89e-21
C8288 state\[2\] _232_/a_114_297# 2.02e-19
C8289 VPWR _337_/a_761_289# 0.00191f
C8290 _190_/a_27_47# net30 0.00291f
C8291 _326_/a_761_289# _314_/a_651_413# 1.09e-20
C8292 _107_ wire42/a_75_212# 0.00449f
C8293 _051_ clknet_2_3__leaf_clk 4.57e-19
C8294 _334_/a_193_47# rebuffer1/a_75_212# 1.5e-19
C8295 _316_/a_193_47# _013_ 0.00485f
C8296 _192_/a_174_21# _099_ 4.16e-20
C8297 _192_/a_27_47# _095_ 0.149f
C8298 net2 _208_/a_439_47# 3.89e-19
C8299 _087_ net55 0.0879f
C8300 VPWR _302_/a_109_297# -0.00347f
C8301 _305_/a_193_47# _076_ 6.5e-19
C8302 clkbuf_2_0__f_clk/a_110_47# en_co_clk 0.0217f
C8303 _327_/a_27_47# net30 9.27e-21
C8304 _291_/a_35_297# net33 0.00618f
C8305 _122_ _298_/a_215_47# 0.0162f
C8306 _292_/a_78_199# _340_/a_1032_413# 6.61e-19
C8307 net3 state\[1\] 0.00998f
C8308 _074_ _085_ 0.033f
C8309 _306_/a_543_47# _305_/a_27_47# 0.00347f
C8310 _326_/a_27_47# _310_/a_1108_47# 4.22e-22
C8311 _326_/a_761_289# _310_/a_543_47# 0.00116f
C8312 _326_/a_193_47# _310_/a_1283_21# 3.39e-19
C8313 output32/a_27_47# net37 0.00802f
C8314 net43 _321_/a_1108_47# 0.0154f
C8315 _303_/a_1462_47# _069_ 7.35e-20
C8316 _338_/a_193_47# clknet_2_3__leaf_clk 0.35f
C8317 output20/a_27_47# _312_/a_761_289# 0.0034f
C8318 output12/a_27_47# ctln[7] 4.45e-20
C8319 ctln[6] output13/a_27_47# 1.71e-19
C8320 clknet_2_1__leaf_clk _208_/a_76_199# 0.00533f
C8321 _334_/a_1108_47# net46 4.95e-19
C8322 clk output41/a_27_47# 1.65e-19
C8323 VPWR _340_/a_1032_413# -0.00678f
C8324 _329_/a_193_47# _274_/a_75_212# 1.35e-19
C8325 net43 _313_/a_193_47# 0.00757f
C8326 _134_ _122_ 0.084f
C8327 _341_/a_1462_47# _038_ 3.39e-20
C8328 _315_/a_27_47# _095_ 5.58e-22
C8329 _100_ _242_/a_79_21# 0.00506f
C8330 _336_/a_543_47# clknet_2_2__leaf_clk 0.00149f
C8331 VPWR _253_/a_81_21# 0.0212f
C8332 _113_ _267_/a_59_75# 6.11e-20
C8333 _042_ _020_ 0.0462f
C8334 net51 _077_ 1.67e-19
C8335 _270_/a_59_75# _109_ 1.23e-19
C8336 _190_/a_27_47# _072_ 3.88e-19
C8337 _190_/a_215_47# cal_itt\[3\] 1.18e-19
C8338 _306_/a_543_47# net51 1.5e-19
C8339 _321_/a_1283_21# _101_ 0.0616f
C8340 net12 _324_/a_27_47# 5.32e-19
C8341 _338_/a_562_413# net18 5.82e-19
C8342 output24/a_27_47# net25 2.02e-20
C8343 _006_ _140_/a_68_297# 4.01e-20
C8344 _341_/a_27_47# net18 0.017f
C8345 _341_/a_193_47# _341_/a_448_47# -0.00779f
C8346 clk cal_count\[3\] 1.09e-20
C8347 _301_/a_47_47# _129_ 6.02e-20
C8348 _134_ _299_/a_27_413# 1.33e-21
C8349 _122_ _130_ -4.05e-24
C8350 _320_/a_805_47# net44 -0.00125f
C8351 _263_/a_297_47# net55 0.00256f
C8352 VPWR clkbuf_0_clk/a_110_47# 0.128f
C8353 trimb[1] output40/a_27_47# 0.00214f
C8354 _341_/a_1270_413# _037_ 8.1e-21
C8355 _104_ _227_/a_209_311# 1.02e-19
C8356 output34/a_27_47# _176_/a_27_47# 0.00787f
C8357 net47 _303_/a_1108_47# 0.014f
C8358 _337_/a_1283_21# _101_ 4.33e-21
C8359 net31 net37 0.249f
C8360 _335_/a_543_47# net46 0.0341f
C8361 _032_ _330_/a_1283_21# 4.72e-19
C8362 net13 _313_/a_1462_47# 3.89e-20
C8363 _281_/a_103_199# _049_ 0.00104f
C8364 _328_/a_543_47# _058_ 0.0026f
C8365 net15 _247_/a_27_297# 0.00809f
C8366 net34 net38 0.481f
C8367 clk _331_/a_27_47# 0.0236f
C8368 _169_/a_215_311# _318_/a_651_413# 8.32e-20
C8369 _199_/a_109_297# _069_ 7.36e-19
C8370 _299_/a_27_413# _130_ 0.043f
C8371 _299_/a_215_297# _129_ 0.0274f
C8372 _329_/a_448_47# trim_mask\[2\] 8.76e-20
C8373 _074_ _314_/a_543_47# 0.00163f
C8374 net4 cal_count\[3\] 0.0122f
C8375 clknet_2_0__leaf_clk _095_ 0.0837f
C8376 _324_/a_27_47# net44 0.0194f
C8377 _027_ _108_ 8.23e-22
C8378 _286_/a_505_21# cal_count\[0\] 0.0603f
C8379 _339_/a_1602_47# _122_ 9.53e-20
C8380 _332_/a_761_289# net46 0.0153f
C8381 VPWR _282_/a_68_297# 0.00657f
C8382 _105_ _279_/a_396_47# 9.38e-20
C8383 _336_/a_1108_47# _107_ 0.00111f
C8384 output40/a_27_47# trimb[4] 0.00959f
C8385 _019_ _321_/a_27_47# 7.83e-21
C8386 _199_/a_193_297# _070_ 1.01e-19
C8387 _001_ _202_/a_79_21# 3.4e-20
C8388 _307_/a_193_47# _307_/a_543_47# -0.00264f
C8389 _307_/a_27_47# _307_/a_1283_21# -9.15e-20
C8390 output32/a_27_47# trim[1] 0.0148f
C8391 net4 _331_/a_27_47# 1.01e-19
C8392 result[2] mask\[1\] 0.00154f
C8393 _304_/a_543_47# _001_ 0.0118f
C8394 _298_/a_292_297# _133_ 0.00556f
C8395 _323_/a_543_47# clknet_2_3__leaf_clk 2.78e-20
C8396 _310_/a_193_47# _310_/a_448_47# -0.00482f
C8397 _253_/a_81_21# net52 1.82e-19
C8398 state\[0\] _317_/a_1108_47# 1.75e-19
C8399 net47 _297_/a_47_47# 1.21e-19
C8400 output22/a_27_47# result[0] 0.00895f
C8401 VPWR _179_/a_27_47# 0.0501f
C8402 net21 _313_/a_761_289# 9.46e-19
C8403 state\[2\] _318_/a_448_47# 3.21e-21
C8404 VPWR _038_ 0.0558f
C8405 cal_count\[1\] _340_/a_1602_47# 0.00724f
C8406 _122_ cal_count\[3\] 4.88e-19
C8407 _303_/a_1108_47# net44 1.56e-20
C8408 clkbuf_0_clk/a_110_47# _063_ 0.013f
C8409 VPWR _204_/a_75_212# 0.072f
C8410 _107_ _206_/a_27_93# 1.04e-19
C8411 mask\[6\] mask\[2\] 1.18e-20
C8412 _302_/a_27_297# clknet_2_2__leaf_clk 2.3e-20
C8413 net2 net37 0.61f
C8414 _313_/a_1108_47# _312_/a_193_47# 9.89e-22
C8415 VPWR _338_/a_476_47# 0.00116f
C8416 _341_/a_1283_21# clknet_2_3__leaf_clk 0.0722f
C8417 _309_/a_651_413# _081_ 8.91e-20
C8418 _309_/a_1108_47# _006_ 1.26e-19
C8419 calibrate _052_ 0.233f
C8420 _235_/a_79_21# _232_/a_32_297# 3.62e-19
C8421 _323_/a_1283_21# _303_/a_27_47# 2.93e-20
C8422 _323_/a_543_47# _303_/a_193_47# 2.56e-20
C8423 _323_/a_193_47# _303_/a_543_47# 3.24e-19
C8424 _323_/a_761_289# _303_/a_761_289# 7e-20
C8425 state\[0\] _192_/a_27_47# 1.55e-21
C8426 _037_ cal_count\[3\] 4.07e-20
C8427 trim_mask\[3\] _256_/a_27_297# 3.89e-20
C8428 _030_ net46 0.0534f
C8429 cal_itt\[2\] _053_ 3.35e-19
C8430 _066_ trim_mask\[4\] 2.16e-20
C8431 trim[1] net31 0.0412f
C8432 _316_/a_448_47# net41 0.0212f
C8433 net43 _313_/a_1462_47# -9.14e-19
C8434 fanout46/a_27_47# _335_/a_761_289# 0.00111f
C8435 _339_/a_27_47# _339_/a_476_47# -0.0251f
C8436 _339_/a_193_47# _339_/a_652_21# -0.00688f
C8437 _336_/a_639_47# trim_mask\[4\] 0.00435f
C8438 _078_ mask\[5\] 0.19f
C8439 net13 _320_/a_193_47# 0.00871f
C8440 _106_ clknet_2_2__leaf_clk 1.18e-19
C8441 _308_/a_1283_21# _307_/a_1108_47# 1.05e-20
C8442 _035_ _001_ 1.09e-19
C8443 net27 result[7] 8.81e-19
C8444 _051_ _266_/a_68_297# 4.76e-20
C8445 net15 net29 0.0176f
C8446 _015_ net45 0.0232f
C8447 clknet_2_1__leaf_clk _314_/a_27_47# 0.162f
C8448 _307_/a_193_47# _138_/a_27_47# 0.00105f
C8449 _336_/a_543_47# _279_/a_204_297# 4.32e-20
C8450 _336_/a_1108_47# _279_/a_27_47# 7.96e-19
C8451 _034_ _065_ 0.148f
C8452 output22/a_27_47# net14 1.67e-19
C8453 VPWR _316_/a_448_47# 0.00228f
C8454 _332_/a_193_47# _332_/a_651_413# -0.00701f
C8455 _332_/a_1108_47# _108_ 8.3e-20
C8456 _288_/a_59_75# _132_ 9.11e-19
C8457 _029_ _108_ 0.104f
C8458 _029_ _332_/a_543_47# 4.58e-19
C8459 _050_ _100_ 8.69e-21
C8460 _120_ _049_ 0.0916f
C8461 _146_/a_68_297# _310_/a_27_47# 4.56e-21
C8462 fanout43/a_27_47# net22 4.37e-22
C8463 _127_ _125_ 0.0731f
C8464 state\[2\] _255_/a_27_47# 3.59e-21
C8465 _162_/a_27_47# _333_/a_1108_47# 0.00116f
C8466 ctlp[0] net29 4.27e-19
C8467 ctln[6] _331_/a_1270_413# 1.07e-21
C8468 _305_/a_193_47# _068_ 2.12e-20
C8469 _141_/a_27_47# net45 0.0379f
C8470 ctln[2] trim[3] 2.75e-19
C8471 _251_/a_373_47# net15 5.93e-19
C8472 _015_ _065_ 2.22e-19
C8473 _026_ trim_mask\[2\] 0.0592f
C8474 _333_/a_1283_21# net32 0.00146f
C8475 net26 _085_ 1.3e-20
C8476 _319_/a_1108_47# _283_/a_75_212# 0.00442f
C8477 VPWR trim_mask\[2\] 0.826f
C8478 _326_/a_193_47# _251_/a_109_297# 1.92e-20
C8479 _324_/a_1217_47# net44 2.37e-19
C8480 net12 _090_ 0.0052f
C8481 _200_/a_80_21# _062_ 0.0146f
C8482 net7 _317_/a_27_47# 1.44e-20
C8483 net15 _317_/a_761_289# 0.0136f
C8484 _076_ _049_ 0.0557f
C8485 net3 _337_/a_1108_47# 6.9e-20
C8486 trim_mask\[0\] clknet_2_2__leaf_clk 0.0931f
C8487 trim_val\[1\] net37 8.1e-20
C8488 _306_/a_761_289# _049_ 4.88e-20
C8489 _326_/a_1108_47# clknet_2_1__leaf_clk 0.00135f
C8490 _306_/a_27_47# net30 6.46e-21
C8491 _167_/a_161_47# net3 0.0394f
C8492 VPWR _323_/a_1108_47# -0.00718f
C8493 _013_ net14 3.23e-20
C8494 cal _315_/a_639_47# 3.17e-19
C8495 _314_/a_1108_47# net29 0.0114f
C8496 _322_/a_805_47# net44 0.00114f
C8497 VPWR _298_/a_292_297# -5.21e-19
C8498 state\[0\] clknet_2_0__leaf_clk 2.17e-20
C8499 _329_/a_27_47# _026_ 0.0414f
C8500 _074_ _310_/a_805_47# 7.09e-19
C8501 _128_ _122_ 0.0321f
C8502 _309_/a_27_47# _308_/a_448_47# 5.28e-21
C8503 _309_/a_193_47# _308_/a_1108_47# 7.29e-21
C8504 _309_/a_543_47# _308_/a_543_47# 5.29e-20
C8505 _329_/a_27_47# VPWR 0.104f
C8506 _074_ _093_ 1.57e-19
C8507 output29/a_27_47# _314_/a_193_47# 0.00864f
C8508 _126_ _125_ 0.272f
C8509 VPWR output22/a_27_47# 0.0828f
C8510 net43 _320_/a_193_47# 0.00113f
C8511 cal_count\[1\] _041_ 0.0426f
C8512 _335_/a_1283_21# _032_ 1.97e-20
C8513 _051_ _028_ 0.156f
C8514 _015_ _243_/a_109_297# 2.1e-19
C8515 _305_/a_27_47# _305_/a_543_47# -0.00936f
C8516 _305_/a_193_47# _305_/a_761_289# -0.0145f
C8517 _299_/a_215_297# _297_/a_47_47# 4.73e-20
C8518 _127_ net40 1.19e-19
C8519 _277_/a_75_212# _057_ 6.35e-20
C8520 en_co_clk cal_itt\[3\] 1.08e-19
C8521 _280_/a_75_212# net18 6.73e-20
C8522 _325_/a_193_47# _313_/a_543_47# 2.85e-21
C8523 _325_/a_761_289# _313_/a_761_289# 3.75e-20
C8524 _325_/a_543_47# _313_/a_193_47# 3.45e-20
C8525 net30 sample 0.00301f
C8526 _072_ rebuffer5/a_161_47# 4.08e-21
C8527 net30 net40 0.00175f
C8528 trim_mask\[1\] net46 0.045f
C8529 net44 _312_/a_543_47# 0.002f
C8530 _078_ _017_ 1.16e-19
C8531 VPWR _341_/a_448_47# -0.00467f
C8532 trim_val\[3\] _258_/a_27_297# 1.39e-19
C8533 _310_/a_193_47# net29 9.97e-20
C8534 _013_ net41 0.107f
C8535 net24 mask\[2\] 0.598f
C8536 _320_/a_27_47# _101_ 7.48e-21
C8537 VPWR _115_ 0.254f
C8538 _303_/a_761_289# clknet_2_3__leaf_clk 0.0429f
C8539 net13 _320_/a_1462_47# 5.11e-19
C8540 _149_/a_150_297# mask\[4\] 5.78e-19
C8541 _117_ _335_/a_193_47# 8.94e-20
C8542 _116_ _335_/a_761_289# 1.75e-20
C8543 _110_ _335_/a_543_47# 0.00158f
C8544 _257_/a_373_47# net18 1.51e-19
C8545 _309_/a_1283_21# _140_/a_68_297# 0.00109f
C8546 _305_/a_543_47# net51 0.00137f
C8547 _030_ _269_/a_81_21# 0.00419f
C8548 _321_/a_1283_21# _248_/a_27_297# 0.0186f
C8549 ctlp[1] net15 0.0339f
C8550 net43 _307_/a_761_289# 3.38e-19
C8551 trim_val\[2\] _334_/a_761_289# 0.00131f
C8552 net48 _334_/a_27_47# 0.00996f
C8553 _002_ rebuffer4/a_27_47# 1.05e-19
C8554 _320_/a_639_47# _040_ 0.00474f
C8555 _096_ _092_ 0.229f
C8556 net55 _099_ 0.103f
C8557 _194_/a_199_47# _118_ 9.57e-20
C8558 _018_ _310_/a_27_47# 2.75e-21
C8559 VPWR _308_/a_1283_21# 0.0747f
C8560 _327_/a_27_47# _066_ 1.59e-20
C8561 _140_/a_68_297# _245_/a_109_297# 5.91e-20
C8562 output22/a_27_47# net23 3.74e-20
C8563 net22 sample 2.63e-19
C8564 _336_/a_1108_47# _118_ 8.28e-20
C8565 _328_/a_1283_21# net40 1.77e-21
C8566 _065_ _208_/a_76_199# 0.103f
C8567 _306_/a_27_47# _072_ 2.88e-19
C8568 _306_/a_193_47# cal_itt\[3\] 2.53e-19
C8569 _337_/a_27_47# _095_ 0.00525f
C8570 _106_ _279_/a_204_297# 0.00183f
C8571 net12 _048_ 0.489f
C8572 clk en 0.0348f
C8573 VPWR _013_ 0.17f
C8574 _292_/a_78_199# _339_/a_1182_261# 0.0121f
C8575 _126_ net40 0.234f
C8576 _088_ _171_/a_27_47# 5.46e-19
C8577 _110_ _332_/a_761_289# 7.59e-20
C8578 _041_ net19 0.013f
C8579 VPWR net38 0.142f
C8580 trim_mask\[0\] trim_val\[0\] 0.394f
C8581 _042_ _310_/a_543_47# 5.03e-21
C8582 _303_/a_27_47# _303_/a_543_47# -0.00454f
C8583 _303_/a_193_47# _303_/a_761_289# -0.0105f
C8584 _239_/a_27_297# _052_ 2.78e-19
C8585 _169_/a_215_311# net55 1.35e-20
C8586 _169_/a_109_53# _096_ 8.02e-19
C8587 VPWR _320_/a_639_47# 8.7e-19
C8588 VPWR _339_/a_1182_261# 0.0122f
C8589 net12 trim_mask\[4\] 0.0958f
C8590 _124_ _123_ 0.0129f
C8591 _064_ _336_/a_193_47# 3.71e-20
C8592 clknet_2_1__leaf_clk _310_/a_651_413# 0.0278f
C8593 net15 mask\[0\] 0.124f
C8594 _071_ _062_ 2.92e-19
C8595 _048_ net44 2e-20
C8596 _333_/a_761_289# _055_ 2.51e-21
C8597 clknet_0_clk _089_ 2.95e-21
C8598 net13 _322_/a_193_47# 0.0153f
C8599 net9 _334_/a_543_47# 4.91e-19
C8600 _308_/a_1283_21# net23 0.00142f
C8601 _258_/a_373_47# trim_mask\[4\] 1.19e-19
C8602 ctlp[6] _312_/a_448_47# 7.83e-20
C8603 _112_ rebuffer2/a_75_212# 1.37e-19
C8604 _337_/a_761_289# _034_ 3.46e-19
C8605 trim_mask\[1\] _332_/a_448_47# 1.91e-20
C8606 net49 _332_/a_1108_47# 2.02e-19
C8607 _136_ _109_ 0.00114f
C8608 trim_val\[2\] rebuffer1/a_75_212# 0.00255f
C8609 _262_/a_27_47# _062_ 3.41e-21
C8610 _041_ _001_ 8.1e-20
C8611 _059_ net45 1.18e-20
C8612 _338_/a_1182_261# _001_ 5.8e-20
C8613 VPWR _307_/a_805_47# 2.38e-19
C8614 _329_/a_1217_47# _026_ 7.86e-21
C8615 _309_/a_27_47# _005_ 9.51e-20
C8616 _294_/a_68_297# _131_ 0.0477f
C8617 _301_/a_47_47# _265_/a_81_21# 1.43e-20
C8618 _329_/a_1217_47# VPWR 6.3e-20
C8619 _256_/a_27_297# _118_ 2.6e-19
C8620 trim_mask\[0\] _279_/a_204_297# 0.0551f
C8621 _256_/a_109_297# trim_val\[4\] 9.23e-20
C8622 _110_ _030_ 0.00981f
C8623 comp clkc 0.0375f
C8624 net43 _320_/a_1462_47# 1.48e-19
C8625 _309_/a_651_413# net14 0.00184f
C8626 _171_/a_27_47# _108_ 1.1e-19
C8627 en_co_clk _131_ 0.00178f
C8628 _094_ _192_/a_505_280# 5.63e-20
C8629 net16 rebuffer1/a_75_212# 0.0176f
C8630 cal_itt\[0\] _195_/a_535_374# 6.42e-19
C8631 cal_itt\[1\] _195_/a_218_374# 9.79e-19
C8632 net43 net13 0.126f
C8633 clknet_2_1__leaf_clk _247_/a_109_297# 0.00436f
C8634 _311_/a_193_47# net26 0.554f
C8635 cal_count\[1\] _129_ 0.0153f
C8636 _059_ _065_ 0.00213f
C8637 _309_/a_1108_47# _245_/a_109_297# 6.06e-22
C8638 _322_/a_27_47# _322_/a_761_289# -0.0169f
C8639 _256_/a_373_47# _058_ 2.63e-19
C8640 net50 trim_mask\[2\] 0.00675f
C8641 _305_/a_1108_47# clknet_2_1__leaf_clk 9.63e-21
C8642 _331_/a_27_47# _331_/a_761_289# -0.00784f
C8643 calibrate _170_/a_384_47# 7.93e-19
C8644 VPWR _303_/a_1283_21# 0.0551f
C8645 _269_/a_299_297# trim_val\[1\] 0.0498f
C8646 _269_/a_81_21# trim_mask\[1\] 0.0607f
C8647 _146_/a_68_297# clknet_2_1__leaf_clk 0.0653f
C8648 _323_/a_448_47# net19 0.00137f
C8649 ctln[2] _057_ 0.0674f
C8650 _239_/a_27_297# calibrate 0.0201f
C8651 net5 en_co_clk 6.94e-19
C8652 net9 _332_/a_27_47# 4.94e-19
C8653 net9 _268_/a_75_212# 0.00327f
C8654 _033_ trim_val\[4\] 5.22e-21
C8655 net35 net32 2.58e-19
C8656 _306_/a_1462_47# cal_itt\[3\] 6.42e-19
C8657 _101_ rebuffer6/a_27_47# 3.72e-21
C8658 net43 _198_/a_27_47# 7.84e-20
C8659 cal_count\[1\] _339_/a_1032_413# 0.0124f
C8660 _036_ _339_/a_1182_261# 9.37e-20
C8661 _319_/a_543_47# _120_ 1.27e-19
C8662 _319_/a_1283_21# en_co_clk 2.97e-21
C8663 _329_/a_193_47# trim_mask\[3\] 0.003f
C8664 _051_ _095_ 6.97e-20
C8665 _224_/a_113_297# net29 0.002f
C8666 net7 net6 0.00138f
C8667 _324_/a_193_47# _101_ 5.02e-20
C8668 mask\[6\] _074_ 0.491f
C8669 _079_ sample 0.00111f
C8670 _078_ _310_/a_27_47# 0.00749f
C8671 VPWR _309_/a_651_413# -0.00793f
C8672 wire42/a_75_212# _062_ 4.31e-19
C8673 net19 net18 3.97e-19
C8674 _276_/a_59_75# _117_ 0.00538f
C8675 _328_/a_448_47# net46 4.11e-19
C8676 _326_/a_193_47# _011_ 0.00135f
C8677 _326_/a_543_47# _086_ 0.00197f
C8678 _291_/a_117_297# trimb[1] 2.67e-19
C8679 _277_/a_75_212# _027_ 3.83e-21
C8680 output24/a_27_47# _310_/a_193_47# 5.71e-21
C8681 _053_ net55 0.0461f
C8682 _064_ _067_ 0.0242f
C8683 VPWR _339_/a_1296_47# 1.86e-19
C8684 _231_/a_161_47# net18 1.49e-19
C8685 _136_ _092_ 0.148f
C8686 _104_ _336_/a_805_47# 4.96e-19
C8687 _104_ _264_/a_27_297# 6.77e-21
C8688 trim_mask\[3\] net18 0.692f
C8689 mask\[7\] _158_/a_150_297# 9.44e-19
C8690 net12 _249_/a_27_297# 0.00691f
C8691 _328_/a_1283_21# _271_/a_75_212# 2.79e-19
C8692 _322_/a_27_47# _101_ 0.0181f
C8693 net12 mask\[3\] 0.011f
C8694 _305_/a_27_47# net30 4.23e-20
C8695 _034_ _282_/a_68_297# 1.49e-19
C8696 _238_/a_75_212# _093_ 0.0377f
C8697 net44 _283_/a_75_212# 3.92e-21
C8698 _321_/a_193_47# mask\[2\] 0.00815f
C8699 VPWR _324_/a_805_47# 4.08e-19
C8700 _107_ net18 2.1e-20
C8701 calibrate _192_/a_27_47# 2.36e-20
C8702 _093_ _192_/a_174_21# 8.93e-19
C8703 _338_/a_1296_47# _001_ 1.29e-19
C8704 _053_ _067_ 0.0272f
C8705 _110_ trim_mask\[1\] 0.0802f
C8706 _001_ net18 0.00937f
C8707 _041_ mask\[1\] 0.0171f
C8708 _053_ _070_ 1.58e-19
C8709 _309_/a_805_47# net43 6.2e-19
C8710 _024_ trim_val\[4\] 1.29e-20
C8711 _258_/a_27_297# _327_/a_543_47# 1.14e-20
C8712 _323_/a_193_47# _152_/a_68_297# 1.58e-20
C8713 output20/a_27_47# ctlp[5] 5.22e-20
C8714 _327_/a_448_47# trim_mask\[0\] 7.47e-20
C8715 _327_/a_543_47# _024_ 0.00402f
C8716 _053_ _304_/a_805_47# 6.41e-19
C8717 _195_/a_505_21# _065_ 2.68e-19
C8718 clkbuf_2_0__f_clk/a_110_47# _049_ 0.0271f
C8719 _005_ _101_ 2.24e-20
C8720 net44 _249_/a_27_297# 2.04e-19
C8721 net45 _137_/a_150_297# 1.59e-19
C8722 _316_/a_1283_21# _095_ 4.44e-20
C8723 _270_/a_59_75# net46 1.89e-20
C8724 _053_ _340_/a_652_21# 2.67e-20
C8725 ctlp[7] net27 1.3e-20
C8726 net51 net30 8.47e-20
C8727 VPWR _322_/a_639_47# 4.88e-19
C8728 clknet_2_1__leaf_clk _018_ 0.0945f
C8729 VPWR _331_/a_639_47# 1.22e-19
C8730 _314_/a_651_413# _011_ 0.00105f
C8731 _312_/a_27_47# net20 0.0263f
C8732 mask\[3\] net44 0.294f
C8733 net28 _312_/a_193_47# 1.5e-20
C8734 _078_ _311_/a_761_289# 1.33e-20
C8735 _219_/a_109_297# _101_ 9.22e-19
C8736 _312_/a_27_47# net53 1.2e-19
C8737 VPWR _046_ 0.555f
C8738 _076_ _202_/a_297_47# 6.01e-21
C8739 _074_ _315_/a_193_47# 0.0166f
C8740 calibrate _315_/a_27_47# 0.00331f
C8741 _324_/a_543_47# _312_/a_1283_21# 0.00141f
C8742 _257_/a_109_297# _025_ 1.7e-19
C8743 _058_ net4 4.91e-20
C8744 _324_/a_27_47# net19 3.72e-19
C8745 _331_/a_193_47# _260_/a_93_21# 5.77e-21
C8746 _010_ _158_/a_68_297# 2.42e-19
C8747 _060_ clk 1.07e-20
C8748 _272_/a_81_21# _272_/a_384_47# 2.22e-34
C8749 VPWR _312_/a_761_289# -0.00107f
C8750 net15 _319_/a_448_47# 0.00961f
C8751 _327_/a_639_47# _136_ 3.85e-19
C8752 net4 mask\[4\] 1.18e-20
C8753 _060_ clone7/a_27_47# 0.078f
C8754 net12 net54 3.08e-20
C8755 _305_/a_27_47# _072_ 0.0117f
C8756 _305_/a_193_47# cal_itt\[3\] 6.76e-21
C8757 _071_ net2 1.4e-19
C8758 _235_/a_79_21# _100_ 3.23e-20
C8759 _187_/a_212_413# cal_count\[2\] 3.89e-19
C8760 output35/a_27_47# _047_ 0.00251f
C8761 net27 _313_/a_543_47# 2.25e-20
C8762 cal_itt\[2\] _305_/a_1270_413# 9.87e-20
C8763 _071_ _305_/a_1283_21# 0.0266f
C8764 _237_/a_218_47# _048_ 1.16e-19
C8765 _229_/a_27_297# _090_ 0.00623f
C8766 _327_/a_27_47# _341_/a_27_47# 4.43e-21
C8767 _066_ net40 4.32e-20
C8768 VPWR _242_/a_79_21# -0.0142f
C8769 VPWR _275_/a_384_47# -2.75e-19
C8770 _228_/a_79_21# _100_ 0.0112f
C8771 _078_ _310_/a_1217_47# 3.02e-19
C8772 _068_ _201_/a_113_47# 1.96e-19
C8773 _060_ net4 1.05e-19
C8774 cal_count\[1\] _297_/a_47_47# 5.21e-20
C8775 _056_ net46 4.84e-20
C8776 net24 _074_ 0.05f
C8777 net51 _072_ 2.5e-20
C8778 _303_/a_1108_47# net19 0.00455f
C8779 _337_/a_448_47# en_co_clk 5.36e-19
C8780 calibrate clknet_2_0__leaf_clk 0.0216f
C8781 _074_ _014_ 1.05e-21
C8782 net54 net44 1.35e-20
C8783 net13 net3 0.0105f
C8784 _033_ _330_/a_193_47# 4.32e-20
C8785 _336_/a_27_47# net46 4.72e-20
C8786 state\[0\] _051_ 0.205f
C8787 cal _316_/a_761_289# 2.1e-20
C8788 net1 _316_/a_193_47# 6.22e-20
C8789 VPWR _333_/a_27_47# 0.022f
C8790 _322_/a_1217_47# _101_ 2.21e-19
C8791 input3/a_75_212# valid 9.25e-19
C8792 _008_ _218_/a_113_297# 0.15f
C8793 _270_/a_59_75# _332_/a_448_47# 4.39e-20
C8794 _341_/a_761_289# _092_ 1.29e-21
C8795 net52 _046_ 1.65e-19
C8796 _101_ net21 3.33e-21
C8797 _062_ _206_/a_27_93# 0.00558f
C8798 _337_/a_1108_47# _076_ 0.00105f
C8799 _053_ _284_/a_150_297# 3.68e-19
C8800 _092_ _098_ 0.0892f
C8801 _097_ _232_/a_32_297# 3.18e-20
C8802 net8 _334_/a_805_47# 4.44e-19
C8803 _325_/a_543_47# net13 0.00146f
C8804 _303_/a_1108_47# _001_ 2.64e-20
C8805 _053_ _338_/a_27_47# 1.98e-21
C8806 _052_ clone1/a_27_47# 4.47e-19
C8807 _119_ _028_ 2.08e-20
C8808 _280_/a_75_212# trim_mask\[4\] 2.45e-20
C8809 _190_/a_655_47# clkbuf_2_3__f_clk/a_110_47# 2.98e-21
C8810 _038_ _193_/a_109_297# 0.00313f
C8811 ctln[5] ctln[6] 0.00305f
C8812 _277_/a_75_212# _032_ 0.00264f
C8813 _251_/a_27_297# _022_ 0.00181f
C8814 trim_mask\[0\] _278_/a_27_47# 6.4e-21
C8815 mask\[6\] net26 1.39e-19
C8816 _312_/a_1217_47# net20 8.49e-20
C8817 net12 net27 0.331f
C8818 clknet_0_clk _092_ 0.206f
C8819 _323_/a_193_47# mask\[5\] 6.07e-19
C8820 _308_/a_1108_47# mask\[1\] 1.87e-20
C8821 _048_ _229_/a_27_297# 0.00561f
C8822 _212_/a_199_47# net14 3.92e-19
C8823 net2 cal_count\[2\] 0.118f
C8824 _331_/a_543_47# trim_mask\[4\] 3.65e-19
C8825 _331_/a_651_413# _028_ 0.00136f
C8826 _257_/a_373_47# trim_mask\[4\] 1.57e-19
C8827 _051_ _226_/a_27_47# 0.0397f
C8828 clk en_co_clk 0.00988f
C8829 clknet_2_1__leaf_clk _078_ 0.0378f
C8830 VPWR _325_/a_27_47# 0.016f
C8831 state\[0\] _316_/a_1283_21# 0.00225f
C8832 net33 rebuffer2/a_75_212# 1.19e-19
C8833 en_co_clk clone7/a_27_47# 0.00156f
C8834 _332_/a_1283_21# net33 5.11e-20
C8835 net12 rebuffer5/a_161_47# 0.00721f
C8836 _107_ _191_/a_27_297# 9.44e-19
C8837 _305_/a_1217_47# _072_ 5.94e-21
C8838 _189_/a_218_47# wire42/a_75_212# 8.25e-21
C8839 _325_/a_1283_21# _322_/a_27_47# 1.42e-20
C8840 _336_/a_543_47# _108_ 4.04e-19
C8841 net27 net44 0.104f
C8842 net43 _080_ 0.00271f
C8843 rebuffer4/a_27_47# _070_ 5.08e-20
C8844 net18 _118_ 1.71e-19
C8845 net46 _173_/a_27_47# 5.03e-19
C8846 _094_ _337_/a_193_47# 0.0221f
C8847 _327_/a_1283_21# net18 2.81e-19
C8848 _189_/a_408_47# _103_ 2.68e-19
C8849 _313_/a_448_47# _085_ 1.78e-19
C8850 _323_/a_639_47# mask\[4\] 4.1e-19
C8851 _188_/a_27_47# _135_ 1.17e-19
C8852 _050_ net41 1.45e-20
C8853 net4 en_co_clk 0.125f
C8854 net10 _275_/a_299_297# 4.27e-19
C8855 net47 net40 1.13e-20
C8856 _306_/a_1108_47# clkbuf_0_clk/a_110_47# 2.75e-19
C8857 _306_/a_193_47# clk 2.25e-19
C8858 net13 fanout44/a_27_47# 0.00419f
C8859 state\[2\] _098_ 0.0595f
C8860 net12 _306_/a_27_47# 0.0176f
C8861 net44 rebuffer5/a_161_47# 6.17e-19
C8862 _322_/a_27_47# _248_/a_27_297# 2.75e-19
C8863 _144_/a_27_47# net37 1.83e-21
C8864 _328_/a_805_47# trim_mask\[1\] 4.53e-21
C8865 _325_/a_543_47# net43 0.00795f
C8866 _336_/a_1217_47# net46 -3.08e-19
C8867 net5 _061_ 0.00282f
C8868 input1/a_75_212# _013_ 2.53e-20
C8869 VPWR _212_/a_199_47# -1.32e-19
C8870 VPWR _333_/a_1217_47# 3.36e-20
C8871 _195_/a_218_47# _067_ 1.53e-20
C8872 VPWR _050_ 0.853f
C8873 net25 net14 0.00744f
C8874 _068_ _202_/a_297_47# 2.69e-19
C8875 calibrate clone1/a_27_47# 0.0484f
C8876 output32/a_27_47# _162_/a_27_47# 4.49e-19
C8877 trim_mask\[1\] rebuffer3/a_75_212# 8.85e-19
C8878 state\[2\] clknet_0_clk 5.82e-21
C8879 _192_/a_174_21# _192_/a_505_280# -1.42e-32
C8880 ctlp[6] _156_/a_27_47# 0.001f
C8881 _110_ _270_/a_59_75# 0.0511f
C8882 _309_/a_761_289# net25 1.47e-19
C8883 _309_/a_193_47# mask\[3\] 1.96e-19
C8884 cal_itt\[2\] cal_itt\[1\] 0.011f
C8885 clkbuf_2_1__f_clk/a_110_47# _319_/a_761_289# 0.00668f
C8886 _122_ en_co_clk 0.465f
C8887 _106_ _088_ 3.91e-20
C8888 _107_ _090_ 0.00633f
C8889 _325_/a_761_289# _101_ 1.37e-19
C8890 _325_/a_27_47# net52 0.00612f
C8891 _306_/a_27_47# net44 0.0081f
C8892 net42 _262_/a_109_297# 0.00567f
C8893 _003_ rebuffer5/a_161_47# 2.29e-19
C8894 _326_/a_1283_21# _253_/a_299_297# 0.00155f
C8895 output21/a_27_47# _074_ 0.0289f
C8896 _166_/a_161_47# _090_ 1.39e-20
C8897 _123_ cal_count\[2\] 0.277f
C8898 _275_/a_384_47# net50 3.6e-19
C8899 _294_/a_68_297# _299_/a_27_413# 0.00519f
C8900 _341_/a_543_47# _053_ 3.23e-19
C8901 VPWR _152_/a_150_297# 3.1e-19
C8902 _037_ en_co_clk 3.09e-20
C8903 _135_ net33 2.17e-20
C8904 clkbuf_2_2__f_clk/a_110_47# _330_/a_27_47# 0.0293f
C8905 trim[2] net48 2.08e-19
C8906 _049_ cal_itt\[3\] 2.9e-21
C8907 _103_ _170_/a_81_21# 3.65e-19
C8908 clk net7 0.0053f
C8909 net15 _316_/a_193_47# 2.68e-19
C8910 _328_/a_27_47# _328_/a_1108_47# -2.98e-20
C8911 en_co_clk _299_/a_27_413# 1.69e-19
C8912 net2 _202_/a_79_21# 0.0392f
C8913 _337_/a_193_47# _244_/a_27_297# 2.43e-20
C8914 net23 _212_/a_199_47# 0.0015f
C8915 _210_/a_113_297# _078_ 0.00196f
C8916 _210_/a_199_47# mask\[0\] 0.00146f
C8917 _235_/a_297_47# clone7/a_27_47# 8.79e-20
C8918 _328_/a_1283_21# net9 0.0067f
C8919 output31/a_27_47# _047_ 2.51e-19
C8920 net31 _162_/a_27_47# 0.042f
C8921 _305_/a_1283_21# _202_/a_79_21# 0.0114f
C8922 _304_/a_543_47# net2 3.56e-20
C8923 _107_ _242_/a_382_297# 3.55e-19
C8924 _033_ _335_/a_193_47# 6.71e-22
C8925 net24 net26 6.35e-21
C8926 _288_/a_59_75# _130_ 8.84e-22
C8927 _227_/a_209_311# wire42/a_75_212# 7.99e-20
C8928 net28 _158_/a_150_297# 3.76e-19
C8929 cal_count\[3\] trim_val\[4\] 1.44e-20
C8930 _228_/a_297_47# clone7/a_27_47# 3.22e-20
C8931 _321_/a_193_47# _074_ 1.2e-19
C8932 trim_mask\[4\] _260_/a_256_47# 4.14e-20
C8933 _306_/a_193_47# _073_ 0.00579f
C8934 _306_/a_27_47# _003_ 0.0362f
C8935 _093_ net55 0.0155f
C8936 VPWR net25 0.328f
C8937 VPWR _325_/a_1217_47# 1.19e-19
C8938 _317_/a_1283_21# _014_ 1.29e-20
C8939 _317_/a_27_47# state\[1\] 1.02e-19
C8940 _317_/a_1108_47# clknet_2_0__leaf_clk 0.0701f
C8941 _317_/a_543_47# net45 8.79e-20
C8942 _081_ net15 4.63e-20
C8943 _302_/a_27_297# _108_ 6.25e-19
C8944 _048_ net19 0.0218f
C8945 net43 fanout44/a_27_47# 0.0499f
C8946 _103_ _227_/a_296_53# 1.66e-19
C8947 output22/a_27_47# output30/a_27_47# 7.06e-19
C8948 _262_/a_109_297# net30 1.47e-19
C8949 _257_/a_27_297# trim_val\[4\] 0.00148f
C8950 net4 net7 0.0774f
C8951 _322_/a_543_47# mask\[3\] 0.0512f
C8952 _259_/a_27_297# _280_/a_75_212# 6.15e-20
C8953 _307_/a_1283_21# fanout43/a_27_47# 3.85e-22
C8954 _106_ _108_ 0.00823f
C8955 _325_/a_1283_21# net21 0.0015f
C8956 trim_mask\[0\] _088_ 0.0141f
C8957 _110_ _336_/a_27_47# 0.0106f
C8958 trim_mask\[4\] net19 0.00699f
C8959 _324_/a_543_47# mask\[4\] 1.92e-20
C8960 _064_ clknet_2_3__leaf_clk 0.211f
C8961 _094_ _337_/a_1462_47# 2.57e-19
C8962 _333_/a_27_47# _333_/a_448_47# -0.00676f
C8963 _010_ _085_ 0.102f
C8964 _301_/a_47_47# net40 0.00154f
C8965 mask\[7\] _314_/a_1283_21# 0.00165f
C8966 _238_/a_75_212# _014_ 0.00786f
C8967 net46 _172_/a_68_297# 0.00178f
C8968 clknet_2_0__leaf_clk _192_/a_27_47# 3.69e-20
C8969 _136_ net46 0.0557f
C8970 _341_/a_27_47# net40 4.38e-21
C8971 _048_ _107_ 0.175f
C8972 _257_/a_109_47# _058_ 1.22e-19
C8973 net2 _035_ 4.55e-20
C8974 _320_/a_27_47# _077_ 3.13e-20
C8975 net12 _306_/a_1217_47# 8.28e-20
C8976 trim_mask\[3\] trim_mask\[4\] 0.352f
C8977 net4 _286_/a_76_199# 7.84e-21
C8978 _051_ _052_ 0.00898f
C8979 _166_/a_161_47# _048_ 7.08e-20
C8980 _322_/a_761_289# mask\[4\] 2.91e-20
C8981 _299_/a_215_297# net40 0.00375f
C8982 _050_ _164_/a_161_47# 5.94e-19
C8983 net43 _082_ 0.00876f
C8984 net23 net25 2.16e-22
C8985 _126_ _132_ 9.98e-21
C8986 _320_/a_1270_413# mask\[2\] 1.03e-21
C8987 _320_/a_1108_47# _017_ 1.49e-19
C8988 net1 net14 0.0299f
C8989 _248_/a_27_297# net21 8.05e-21
C8990 _053_ clknet_2_3__leaf_clk 1.13f
C8991 _107_ trim_mask\[4\] 0.0049f
C8992 VPWR _169_/a_301_53# -1.01e-19
C8993 trim_mask\[1\] _336_/a_1283_21# 3.51e-19
C8994 clknet_2_0__leaf_clk _315_/a_27_47# 0.0373f
C8995 _087_ _095_ 3.83e-20
C8996 _101_ _045_ 7.28e-21
C8997 _296_/a_113_47# cal_count\[2\] 2.23e-20
C8998 _285_/a_113_47# _067_ 1.96e-20
C8999 _040_ _246_/a_109_47# 0.00443f
C9000 _050_ _260_/a_346_47# 8.98e-19
C9001 _191_/a_27_297# _118_ 7.13e-19
C9002 net25 net52 3.65e-19
C9003 _109_ clknet_2_2__leaf_clk 0.00148f
C9004 trim_mask\[0\] _108_ 0.203f
C9005 trim_mask\[0\] _332_/a_543_47# 0.00719f
C9006 _274_/a_75_212# _334_/a_27_47# 6.05e-21
C9007 _326_/a_1270_413# _102_ 5.01e-20
C9008 _326_/a_639_47# mask\[7\] 1.47e-19
C9009 _286_/a_76_199# _122_ 0.0108f
C9010 _136_ _300_/a_377_297# 6.58e-19
C9011 net1 net41 0.0625f
C9012 _185_/a_68_297# _090_ 1.5e-21
C9013 _309_/a_193_47# fanout43/a_27_47# 3.37e-20
C9014 _041_ _286_/a_535_374# 3.12e-19
C9015 net16 _131_ 0.0107f
C9016 net15 _316_/a_1462_47# 2.71e-19
C9017 _324_/a_543_47# _020_ 7.24e-20
C9018 _324_/a_448_47# mask\[5\] 7.84e-20
C9019 VPWR _246_/a_109_47# -7.39e-19
C9020 _239_/a_27_297# clone1/a_27_47# 7.83e-20
C9021 _192_/a_174_21# _243_/a_27_297# 4.67e-19
C9022 mask\[4\] _101_ 0.227f
C9023 _078_ net45 0.412f
C9024 net34 net37 2.05f
C9025 _340_/a_1602_47# net2 4.96e-19
C9026 VPWR net1 0.0318f
C9027 output24/a_27_47# result[2] 0.00476f
C9028 _104_ net41 1.28e-20
C9029 VPWR _327_/a_805_47# 2.51e-19
C9030 _263_/a_79_21# _092_ 0.00326f
C9031 _317_/a_1217_47# state\[1\] 1.2e-19
C9032 _136_ _332_/a_448_47# 0.00156f
C9033 net5 net16 3.66e-20
C9034 trim_mask\[4\] _279_/a_27_47# 0.0227f
C9035 state\[2\] _331_/a_1108_47# 6.44e-20
C9036 output27/a_27_47# result[6] 7.93e-20
C9037 result[5] output28/a_27_47# 6.68e-19
C9038 ctlp[2] output39/a_27_47# 0.0101f
C9039 output16/a_27_47# trimb[3] 6.54e-19
C9040 _035_ _123_ 1.21e-19
C9041 _051_ calibrate 0.00542f
C9042 trim_mask\[2\] _334_/a_1108_47# 8.01e-19
C9043 _232_/a_32_297# _337_/a_543_47# 5.02e-21
C9044 _319_/a_1283_21# _049_ 0.00262f
C9045 _110_ _336_/a_1217_47# 1.59e-19
C9046 _104_ _026_ 0.00511f
C9047 _078_ _065_ 0.274f
C9048 _324_/a_1283_21# net27 0.00397f
C9049 _104_ VPWR 1.31f
C9050 _162_/a_27_47# trim_val\[1\] 3.66e-20
C9051 _305_/a_193_47# clk 0.00448f
C9052 _305_/a_1108_47# clkbuf_0_clk/a_110_47# 0.00789f
C9053 _312_/a_448_47# _045_ 2.21e-19
C9054 net23 _246_/a_109_47# 3.31e-21
C9055 net20 _084_ 0.00131f
C9056 net12 _305_/a_27_47# 5.89e-19
C9057 _062_ net18 2.2e-19
C9058 _335_/a_27_47# clkbuf_2_2__f_clk/a_110_47# 9.57e-20
C9059 _325_/a_27_47# _325_/a_448_47# -0.0012f
C9060 net55 _171_/a_27_47# 4.04e-19
C9061 _084_ net53 6.92e-21
C9062 _181_/a_68_297# trim_mask\[4\] 0.0366f
C9063 cal_itt\[0\] _304_/a_27_47# 2.9e-21
C9064 net4 cal_count\[0\] 2.07e-19
C9065 _331_/a_193_47# _330_/a_27_47# 0.00133f
C9066 _331_/a_27_47# _330_/a_193_47# 0.00133f
C9067 trim_val\[0\] _109_ 0.00385f
C9068 _255_/a_27_47# _103_ 0.00498f
C9069 _269_/a_81_21# _172_/a_68_297# 0.00128f
C9070 _321_/a_761_289# _018_ 1.1e-20
C9071 _302_/a_109_297# trim_mask\[1\] 2.79e-21
C9072 net13 _076_ 1.04e-20
C9073 _341_/a_761_289# net46 -0.00406f
C9074 _185_/a_68_297# _048_ 8.76e-22
C9075 _078_ _319_/a_27_47# 1.06e-21
C9076 mask\[0\] _319_/a_193_47# 0.0251f
C9077 trim_mask\[3\] _327_/a_27_47# 1.68e-20
C9078 _305_/a_193_47# net4 6.04e-21
C9079 _040_ _208_/a_439_47# 2.37e-20
C9080 _321_/a_193_47# net26 1.99e-19
C9081 net12 net51 0.0437f
C9082 clknet_2_0__leaf_clk _315_/a_1217_47# 2.56e-19
C9083 _321_/a_1108_47# _042_ 0.016f
C9084 _307_/a_27_47# _137_/a_68_297# 3.94e-21
C9085 _020_ _101_ 0.00736f
C9086 _305_/a_27_47# net44 0.0191f
C9087 _255_/a_27_47# _105_ 1.18e-19
C9088 net44 _311_/a_1283_21# 0.00579f
C9089 _306_/a_543_47# rebuffer6/a_27_47# 4.26e-21
C9090 state\[2\] _263_/a_79_21# 7.14e-20
C9091 _321_/a_639_47# clknet_2_1__leaf_clk 0.00108f
C9092 _327_/a_27_47# _107_ 0.00192f
C9093 calibrate _316_/a_1283_21# 5.86e-20
C9094 _093_ _316_/a_543_47# 5.04e-20
C9095 trim[1] net34 0.0403f
C9096 net43 result[5] 7.57e-19
C9097 _259_/a_109_297# trim_val\[3\] 1.23e-20
C9098 _259_/a_27_297# trim_mask\[3\] 0.0886f
C9099 cal_count\[0\] _122_ 0.0263f
C9100 VPWR _208_/a_439_47# 2.35e-19
C9101 _340_/a_1602_47# _123_ 0.00883f
C9102 clknet_2_1__leaf_clk _313_/a_1108_47# 0.0614f
C9103 _236_/a_109_297# _092_ 0.00351f
C9104 net15 net14 6.76e-20
C9105 VPWR ctlp[5] 0.179f
C9106 _301_/a_285_47# _300_/a_47_47# 1.53e-19
C9107 _301_/a_47_47# _300_/a_285_47# 1.53e-19
C9108 net44 net51 0.158f
C9109 _037_ cal_count\[0\] 2.17e-20
C9110 _104_ _063_ 4.99e-20
C9111 net37 _133_ 2.9e-20
C9112 _048_ _118_ 3.3e-20
C9113 _341_/a_27_47# _300_/a_285_47# 6.92e-21
C9114 cal_count\[0\] _299_/a_27_413# 4.7e-20
C9115 net43 _120_ 5.67e-20
C9116 net9 _066_ 2.45e-20
C9117 _337_/a_27_47# _192_/a_27_47# 3.85e-20
C9118 _187_/a_27_413# _134_ 6.26e-19
C9119 ctlp[0] net14 0.00192f
C9120 cal_itt\[0\] _069_ 0.176f
C9121 fanout47/a_27_47# _065_ 1e-19
C9122 VPWR _226_/a_303_47# -9.65e-20
C9123 _110_ _136_ 5.58e-19
C9124 _004_ net45 0.00446f
C9125 _134_ _332_/a_27_47# 2.04e-20
C9126 trim_mask\[0\] net49 5.76e-20
C9127 trim_mask\[4\] _118_ 0.0192f
C9128 state\[2\] clknet_2_2__leaf_clk 2.67e-22
C9129 net15 _040_ 0.0123f
C9130 state\[2\] _260_/a_584_47# 0.00134f
C9131 net15 net41 0.00739f
C9132 en_co_clk _101_ 0.00249f
C9133 net43 _076_ 0.00837f
C9134 _119_ _330_/a_1108_47# 7.31e-20
C9135 net51 _003_ 0.00476f
C9136 cal_itt\[3\] _202_/a_297_47# 1.98e-21
C9137 _187_/a_212_413# _129_ 7.67e-22
C9138 _228_/a_79_21# net41 9.74e-20
C9139 mask\[7\] clknet_2_1__leaf_clk 0.00293f
C9140 _091_ net30 1.3e-19
C9141 net54 _107_ 9.96e-19
C9142 net21 _156_/a_27_47# 1.65e-19
C9143 net43 _306_/a_761_289# 1.24e-20
C9144 VPWR _330_/a_1270_413# 2.57e-19
C9145 cal_itt\[1\] _067_ 0.258f
C9146 trim_mask\[3\] _178_/a_68_297# 0.00411f
C9147 trim_val\[3\] _178_/a_150_297# 1.12e-19
C9148 cal_itt\[1\] _070_ 1.5e-19
C9149 net12 _250_/a_109_297# 0.00775f
C9150 _216_/a_113_297# net25 0.0134f
C9151 _087_ _226_/a_27_47# 0.00102f
C9152 VPWR _267_/a_59_75# 0.0138f
C9153 cal_itt\[2\] _106_ 1.12e-20
C9154 _337_/a_448_47# _049_ 0.009f
C9155 net31 _129_ 1.41e-20
C9156 cal_itt\[1\] _304_/a_805_47# 8.64e-20
C9157 _104_ _260_/a_346_47# 4.68e-19
C9158 VPWR net15 1.74f
C9159 VPWR _235_/a_79_21# 0.0039f
C9160 _188_/a_27_47# net33 0.00552f
C9161 _314_/a_1108_47# net14 0.00242f
C9162 trim_mask\[0\] _227_/a_368_53# 9.85e-19
C9163 cal_count\[1\] _125_ 0.072f
C9164 VPWR _228_/a_79_21# 0.00568f
C9165 _306_/a_193_47# _101_ 0.00382f
C9166 _239_/a_27_297# _051_ -5.55e-35
C9167 mask\[0\] _319_/a_1462_47# 0.00198f
C9168 _050_ _034_ 2.82e-20
C9169 net3 _281_/a_103_199# 1.3e-20
C9170 _320_/a_27_47# clkbuf_2_1__f_clk/a_110_47# 0.013f
C9171 VPWR ctlp[0] 0.0908f
C9172 _307_/a_543_47# _039_ 6.6e-19
C9173 _325_/a_1283_21# mask\[4\] 3.75e-20
C9174 mask\[3\] _248_/a_109_297# 0.0036f
C9175 _308_/a_543_47# _074_ 0.0157f
C9176 ctln[5] net11 0.00713f
C9177 net45 _096_ 1.24e-19
C9178 net27 _312_/a_651_413# 2.35e-19
C9179 _053_ _028_ 2.45e-19
C9180 net14 _310_/a_193_47# 0.0102f
C9181 net2 _298_/a_493_297# 2.43e-20
C9182 net27 net19 0.0249f
C9183 _041_ _123_ 0.0407f
C9184 _233_/a_109_297# net14 0.00183f
C9185 _033_ net30 2.25e-21
C9186 _338_/a_1182_261# _123_ 3.03e-20
C9187 _300_/a_47_47# clknet_2_3__leaf_clk 0.0435f
C9188 _337_/a_27_47# clknet_2_0__leaf_clk 0.171f
C9189 result[6] _314_/a_761_289# 4.99e-19
C9190 net28 _314_/a_1283_21# 2.21e-19
C9191 _191_/a_27_297# _062_ 0.0366f
C9192 _104_ net50 0.363f
C9193 _015_ _050_ 6.2e-21
C9194 _309_/a_543_47# _310_/a_27_47# 1.16e-20
C9195 _309_/a_27_47# _310_/a_543_47# 1.17e-20
C9196 mask\[3\] mask\[1\] 9.14e-20
C9197 net23 net15 0.00814f
C9198 _326_/a_761_289# net43 0.00904f
C9199 _152_/a_68_297# _044_ 0.00346f
C9200 VPWR _306_/a_805_47# 6.92e-20
C9201 _257_/a_27_297# _335_/a_193_47# 3.18e-22
C9202 _323_/a_193_47# clknet_2_1__leaf_clk 0.00116f
C9203 _189_/a_27_47# clkbuf_2_3__f_clk/a_110_47# 0.01f
C9204 cal_itt\[2\] trim_mask\[0\] 1.07e-20
C9205 _168_/a_27_413# _033_ 2.41e-20
C9206 _326_/a_805_47# net14 6.71e-19
C9207 _248_/a_27_297# mask\[4\] 0.00535f
C9208 _095_ _099_ 0.0338f
C9209 net2 net18 0.0112f
C9210 _065_ _096_ 2.11e-19
C9211 _341_/a_1283_21# _135_ 1.09e-19
C9212 VPWR _314_/a_1108_47# 0.0383f
C9213 cal_count\[1\] net40 0.0105f
C9214 VPWR net37 0.288f
C9215 _332_/a_1108_47# clknet_2_3__leaf_clk 1.88e-21
C9216 clk _049_ 0.483f
C9217 _051_ _203_/a_59_75# 7.77e-20
C9218 clk _318_/a_761_289# 0.0185f
C9219 _268_/a_75_212# cal_count\[3\] 2.44e-19
C9220 net15 net52 0.228f
C9221 net12 _318_/a_193_47# 8.6e-19
C9222 net2 _129_ 0.0365f
C9223 net9 net47 0.131f
C9224 _308_/a_1270_413# _039_ 1.6e-20
C9225 _051_ _192_/a_27_47# 3.56e-21
C9226 _336_/a_193_47# _336_/a_543_47# -0.00598f
C9227 _102_ mask\[6\] 0.00305f
C9228 trim_mask\[2\] trim_mask\[1\] 0.0266f
C9229 _314_/a_27_47# _046_ 6.7e-21
C9230 net9 _340_/a_1140_413# 1.65e-19
C9231 _319_/a_193_47# _319_/a_448_47# -0.00297f
C9232 _253_/a_81_21# _078_ 0.011f
C9233 _138_/a_27_47# _039_ 0.0126f
C9234 _307_/a_639_47# _074_ 0.00166f
C9235 output26/a_27_47# net25 3.74e-20
C9236 VPWR _310_/a_193_47# -0.289f
C9237 _326_/a_639_47# net28 1.7e-19
C9238 VPWR _233_/a_109_297# -0.0166f
C9239 net4 _049_ 2.26e-19
C9240 _340_/a_27_47# cal_count\[2\] 0.00347f
C9241 _024_ net30 1.38e-20
C9242 _327_/a_27_47# _118_ 1.7e-20
C9243 _050_ _281_/a_253_47# 8.07e-19
C9244 _327_/a_27_47# _327_/a_1283_21# -1.12e-19
C9245 _164_/a_161_47# net15 0.00151f
C9246 _243_/a_27_297# net55 0.0652f
C9247 _243_/a_109_297# _096_ 0.00538f
C9248 net12 _021_ 7.98e-19
C9249 net43 _314_/a_1270_413# 1.12e-19
C9250 _304_/a_639_47# _065_ 1.91e-19
C9251 clk _317_/a_805_47# 2.74e-19
C9252 _329_/a_27_47# trim_mask\[1\] 8.3e-22
C9253 _317_/a_1108_47# _316_/a_1283_21# 3.54e-22
C9254 net2 _339_/a_1032_413# 2.56e-20
C9255 cal_itt\[0\] _338_/a_193_47# 6.21e-19
C9256 _119_ _052_ 2.32e-21
C9257 _185_/a_68_297# net54 0.00954f
C9258 _028_ _330_/a_448_47# 1.13e-20
C9259 clknet_2_2__leaf_clk _330_/a_651_413# 0.00252f
C9260 _331_/a_448_47# _027_ 9.25e-21
C9261 VPWR _326_/a_805_47# 6.77e-19
C9262 _340_/a_193_47# _065_ 1.53e-20
C9263 trim_val\[2\] _055_ 5.25e-19
C9264 VPWR _334_/a_805_47# 0.0022f
C9265 _017_ _209_/a_27_47# 7.14e-22
C9266 clknet_2_1__leaf_clk clknet_0_clk 0.00445f
C9267 _058_ trim_val\[4\] 0.00626f
C9268 _104_ _279_/a_396_47# 0.0821f
C9269 result[3] _310_/a_27_47# 0.00348f
C9270 _327_/a_543_47# _058_ 0.0112f
C9271 output10/a_27_47# ctln[4] 0.00976f
C9272 net27 _155_/a_68_297# 3.65e-20
C9273 net3 _120_ 2.04e-19
C9274 _231_/a_161_47# net40 4.22e-19
C9275 _320_/a_1108_47# clknet_2_1__leaf_clk 6.67e-22
C9276 net47 _132_ 4.97e-20
C9277 _110_ clknet_0_clk 1.84e-21
C9278 _097_ _316_/a_193_47# 0.00178f
C9279 net16 _055_ 8.2e-22
C9280 VPWR _124_ 0.0937f
C9281 mask\[1\] _246_/a_373_47# 1.91e-20
C9282 net43 _310_/a_1283_21# 0.0593f
C9283 _311_/a_193_47# net53 0.0181f
C9284 _330_/a_639_47# net19 8.45e-19
C9285 mask\[6\] _010_ 3.7e-19
C9286 _021_ net44 0.00643f
C9287 mask\[0\] _282_/a_150_297# 6.75e-20
C9288 _303_/a_651_413# _068_ 2.26e-19
C9289 _049_ _073_ 6.44e-20
C9290 _115_ trim_mask\[1\] 1.95e-19
C9291 _335_/a_1108_47# _119_ 1.34e-21
C9292 _078_ _313_/a_639_47# 1.01e-19
C9293 trim[1] VPWR 0.159f
C9294 net16 _122_ 0.0236f
C9295 _012_ net14 0.0159f
C9296 _324_/a_1283_21# _311_/a_1283_21# 3.86e-20
C9297 _123_ net18 0.00946f
C9298 VPWR _300_/a_129_47# -5.9e-19
C9299 net35 _058_ 0.00316f
C9300 _089_ _088_ 5.01e-19
C9301 _087_ _052_ 3.07e-19
C9302 _337_/a_639_47# net45 3.56e-20
C9303 VPWR _335_/a_1270_413# 1.18e-19
C9304 _306_/a_1283_21# _048_ 3.18e-20
C9305 _323_/a_1270_413# _042_ 3.5e-19
C9306 net43 _068_ 1.05e-19
C9307 _309_/a_448_47# _074_ 0.0102f
C9308 VPWR _311_/a_543_47# 0.015f
C9309 _051_ clknet_2_0__leaf_clk 3.44e-19
C9310 output10/a_27_47# _335_/a_27_47# 3.61e-19
C9311 _015_ _169_/a_301_53# 2.51e-20
C9312 _053_ _279_/a_314_297# 1.27e-20
C9313 _123_ _129_ 8.37e-20
C9314 net16 _299_/a_27_413# 0.00306f
C9315 _239_/a_474_297# _098_ 6.99e-20
C9316 _136_ rebuffer3/a_75_212# 0.0027f
C9317 net14 _224_/a_113_297# 5.51e-19
C9318 _121_ _192_/a_505_280# 9.37e-20
C9319 VPWR _332_/a_651_413# -5.12e-19
C9320 fanout43/a_27_47# mask\[1\] 0.0536f
C9321 _026_ fanout46/a_27_47# 4.89e-21
C9322 net9 _301_/a_47_47# 4.82e-20
C9323 VPWR fanout46/a_27_47# 0.0596f
C9324 mask\[5\] _044_ 0.149f
C9325 _303_/a_1108_47# net2 4.77e-21
C9326 _093_ valid 9.09e-19
C9327 _012_ net41 9.64e-19
C9328 _048_ _062_ 0.0949f
C9329 _284_/a_68_297# rebuffer3/a_75_212# 2.15e-21
C9330 net12 _318_/a_1462_47# 3.18e-19
C9331 _304_/a_193_47# _067_ 2.16e-19
C9332 net9 _341_/a_27_47# 0.00101f
C9333 _218_/a_113_297# _311_/a_27_47# 3e-20
C9334 _336_/a_1108_47# _264_/a_27_297# 1.59e-20
C9335 _336_/a_193_47# _106_ 7.03e-20
C9336 net42 clkbuf_2_3__f_clk/a_110_47# 0.00341f
C9337 clkbuf_0_clk/a_110_47# fanout47/a_27_47# 2.1e-19
C9338 state\[0\] _099_ 3.09e-20
C9339 _339_/a_1032_413# _123_ 0.0695f
C9340 _107_ _228_/a_382_297# 2.25e-19
C9341 _230_/a_59_75# _091_ 0.0189f
C9342 _249_/a_373_47# _020_ 0.00113f
C9343 net43 _305_/a_761_289# 0.0367f
C9344 VPWR _310_/a_1462_47# 2.01e-19
C9345 _136_ _065_ 0.0334f
C9346 trim_mask\[4\] _062_ 1.19e-20
C9347 VPWR _012_ 0.66f
C9348 input1/a_75_212# net1 0.00337f
C9349 _275_/a_299_297# _335_/a_1283_21# 7.21e-20
C9350 _059_ _050_ 0.239f
C9351 _156_/a_27_47# _045_ 0.0153f
C9352 _284_/a_68_297# _065_ 0.0654f
C9353 _008_ _311_/a_193_47# 0.0835f
C9354 net10 net46 3.81e-20
C9355 net45 _316_/a_761_289# -6.9e-19
C9356 clknet_2_0__leaf_clk _316_/a_1283_21# 3.04e-21
C9357 clk state\[1\] 0.00418f
C9358 _169_/a_215_311# state\[0\] 0.0259f
C9359 _337_/a_193_47# net55 1.84e-19
C9360 _014_ _316_/a_543_47# 0.0124f
C9361 VPWR _269_/a_299_297# 0.0241f
C9362 _028_ _027_ 0.00438f
C9363 cal_count\[0\] _297_/a_285_47# 2.37e-20
C9364 clknet_2_2__leaf_clk net46 0.837f
C9365 state\[1\] clone7/a_27_47# 0.00516f
C9366 output37/a_27_47# _126_ 0.0104f
C9367 net43 clkbuf_2_0__f_clk/a_110_47# 4.53e-20
C9368 _307_/a_193_47# net30 1.28e-19
C9369 calibrate _087_ 0.0116f
C9370 VPWR _224_/a_113_297# 0.0524f
C9371 _309_/a_543_47# clknet_2_1__leaf_clk 5.3e-20
C9372 net2 _297_/a_47_47# 0.00997f
C9373 output32/a_27_47# _265_/a_81_21# 2.75e-20
C9374 net13 _042_ 0.0188f
C9375 net24 _006_ 0.0752f
C9376 result[2] _081_ 5.8e-19
C9377 clkbuf_2_3__f_clk/a_110_47# net30 0.00182f
C9378 _074_ _312_/a_193_47# 2.25e-19
C9379 _304_/a_1270_413# _035_ 1.07e-21
C9380 _097_ _316_/a_1462_47# 1.03e-19
C9381 clknet_2_1__leaf_clk _245_/a_27_297# 0.00291f
C9382 output38/a_27_47# net16 0.00105f
C9383 _306_/a_1108_47# _050_ 5.7e-20
C9384 _181_/a_68_297# net40 4.36e-20
C9385 net4 state\[1\] 0.483f
C9386 _299_/a_215_297# _132_ 0.00272f
C9387 _226_/a_27_47# _099_ 2.83e-19
C9388 _326_/a_1108_47# _325_/a_27_47# 3.16e-20
C9389 _161_/a_150_297# trim_val\[0\] 7.82e-19
C9390 _106_ net55 0.00401f
C9391 _333_/a_543_47# rebuffer1/a_75_212# 3.33e-19
C9392 _333_/a_193_47# _332_/a_193_47# 5.9e-22
C9393 net28 clknet_2_1__leaf_clk 0.242f
C9394 _307_/a_27_47# mask\[0\] 0.0111f
C9395 _307_/a_193_47# net22 0.21f
C9396 VPWR _305_/a_805_47# 1.7e-19
C9397 VPWR _250_/a_27_297# 0.124f
C9398 net31 _333_/a_193_47# 9.64e-20
C9399 _265_/a_81_21# _332_/a_193_47# 0.00351f
C9400 _051_ _336_/a_761_289# 1.05e-20
C9401 _324_/a_448_47# clknet_2_1__leaf_clk 8.22e-19
C9402 _329_/a_1108_47# net9 0.0115f
C9403 _050_ _075_ 0.0571f
C9404 _179_/a_27_47# _056_ 6.48e-19
C9405 _176_/a_27_47# _055_ 3.12e-22
C9406 net52 _310_/a_1462_47# 5.5e-20
C9407 _322_/a_1283_21# _250_/a_27_297# 9.71e-22
C9408 _302_/a_27_297# _067_ 0.00366f
C9409 _051_ clone1/a_27_47# 5.88e-20
C9410 _322_/a_193_47# _042_ 7.52e-20
C9411 _246_/a_109_297# mask\[2\] 0.0351f
C9412 _304_/a_761_289# _136_ 0.00121f
C9413 net34 cal_count\[2\] 7.97e-20
C9414 _116_ VPWR 0.129f
C9415 _322_/a_1108_47# clknet_2_1__leaf_clk 1.12e-19
C9416 _304_/a_1462_47# _067_ 4.31e-19
C9417 _304_/a_761_289# _284_/a_68_297# 1.96e-20
C9418 _083_ _311_/a_543_47# 5.28e-20
C9419 _303_/a_543_47# net26 3.75e-20
C9420 trim_val\[0\] net46 0.00323f
C9421 net42 cal_count\[3\] 9.22e-20
C9422 clknet_2_1__leaf_clk _159_/a_27_47# 8.29e-20
C9423 _332_/a_448_47# clknet_2_2__leaf_clk 0.00155f
C9424 VPWR _254_/a_109_297# 0.00112f
C9425 _304_/a_1283_21# net47 0.00784f
C9426 _062_ _190_/a_27_47# 2.48e-19
C9427 cal_itt\[1\] clknet_2_3__leaf_clk 0.00118f
C9428 _200_/a_80_21# VPWR 0.0202f
C9429 _311_/a_1283_21# net19 0.00189f
C9430 _113_ _333_/a_193_47# 6.65e-20
C9431 _030_ _333_/a_27_47# 0.248f
C9432 ctln[7] _318_/a_193_47# 3.63e-20
C9433 net13 _318_/a_543_47# 0.0122f
C9434 _308_/a_1108_47# mask\[0\] 0.00229f
C9435 _308_/a_1283_21# _078_ 0.00166f
C9436 result[3] clknet_2_1__leaf_clk 0.0234f
C9437 net43 _042_ 0.377f
C9438 output15/a_27_47# net28 2.54e-19
C9439 trim_mask\[0\] net55 0.0104f
C9440 _340_/a_27_47# _340_/a_1602_47# -1.94e-19
C9441 _340_/a_193_47# _340_/a_1032_413# -9.67e-21
C9442 _074_ _213_/a_109_297# 0.0012f
C9443 net50 _335_/a_1270_413# 1.41e-19
C9444 trim_val\[3\] _335_/a_805_47# 2.13e-20
C9445 _308_/a_193_47# net24 5.52e-22
C9446 net44 _319_/a_761_289# 5.86e-20
C9447 _210_/a_199_47# net14 1.81e-19
C9448 _318_/a_27_47# net41 1.75e-20
C9449 _308_/a_761_289# clknet_2_0__leaf_clk 6.24e-20
C9450 _308_/a_27_47# net45 2.93e-20
C9451 _299_/a_298_297# cal_count\[2\] 3.59e-19
C9452 _281_/a_103_199# _120_ 0.00823f
C9453 _281_/a_253_297# en_co_clk 0.00324f
C9454 net18 _150_/a_27_47# 0.00337f
C9455 _294_/a_68_297# _288_/a_59_75# 1.56e-20
C9456 VPWR _009_ 0.0178f
C9457 state\[0\] _053_ 0.00132f
C9458 _341_/a_761_289# _065_ 4.41e-19
C9459 _118_ net40 0.00482f
C9460 _327_/a_1283_21# net40 5.37e-20
C9461 net15 _034_ 1.23e-19
C9462 _251_/a_27_297# _101_ 0.034f
C9463 _103_ _098_ 0.0872f
C9464 _250_/a_109_47# _101_ 0.00184f
C9465 net45 clknet_0_clk 0.0745f
C9466 _313_/a_193_47# _313_/a_761_289# -0.0105f
C9467 _313_/a_27_47# _313_/a_543_47# -0.00936f
C9468 cal_itt\[0\] _303_/a_761_289# 1.93e-19
C9469 net13 _022_ 1.44e-20
C9470 net9 _339_/a_956_413# 2.92e-19
C9471 _320_/a_1108_47# net45 1.03e-19
C9472 VPWR _318_/a_27_47# 0.104f
C9473 cal_count\[3\] net30 0.00416f
C9474 net50 fanout46/a_27_47# 1.66e-20
C9475 trim_mask\[2\] _056_ 4.58e-19
C9476 _047_ net32 0.147f
C9477 _232_/a_32_297# _090_ 0.0413f
C9478 mask\[6\] net20 1.84e-19
C9479 _097_ net14 1.49e-20
C9480 _287_/a_75_212# _338_/a_476_47# 3.15e-19
C9481 trim_mask\[0\] _067_ 0.0124f
C9482 mask\[6\] net53 0.00571f
C9483 _103_ clknet_0_clk 0.00673f
C9484 trim_mask\[2\] _336_/a_27_47# 2.46e-19
C9485 _327_/a_1108_47# _267_/a_59_75# 3.19e-19
C9486 _140_/a_68_297# clknet_2_0__leaf_clk 5.04e-20
C9487 net4 _336_/a_651_413# 0.00382f
C9488 _324_/a_1283_21# _021_ 6.94e-21
C9489 _321_/a_1108_47# _143_/a_68_297# 5.65e-20
C9490 clknet_0_clk _065_ 0.288f
C9491 _326_/a_1108_47# net25 8.95e-20
C9492 net33 output40/a_27_47# 0.00169f
C9493 net44 _202_/a_382_297# 2.86e-19
C9494 output23/a_27_47# _213_/a_109_297# 5.98e-20
C9495 net12 _206_/a_206_47# 1.84e-20
C9496 _320_/a_1108_47# _065_ 6.09e-19
C9497 _307_/a_1462_47# net22 5.12e-19
C9498 _064_ _330_/a_1108_47# 8.48e-20
C9499 _104_ _330_/a_543_47# 3.39e-20
C9500 _328_/a_27_47# _026_ 8.37e-20
C9501 _328_/a_27_47# VPWR -0.00349f
C9502 _109_ _108_ 0.00222f
C9503 VPWR _210_/a_199_47# -3.33e-19
C9504 _200_/a_80_21# _063_ 0.0782f
C9505 _189_/a_218_47# _048_ 8.38e-19
C9506 _307_/a_448_47# net45 1.84e-21
C9507 _239_/a_694_21# _089_ 1.88e-19
C9508 trim[3] _334_/a_651_413# 5.61e-20
C9509 _168_/a_27_413# _331_/a_27_47# 6.84e-19
C9510 _308_/a_27_47# _319_/a_27_47# 1.75e-19
C9511 _302_/a_109_297# _136_ 0.00245f
C9512 clknet_0_clk _105_ 0.0125f
C9513 VPWR _317_/a_1270_413# -1.9e-19
C9514 _307_/a_193_47# _079_ 4.88e-19
C9515 _315_/a_543_47# net14 0.00521f
C9516 _097_ net41 3.65e-19
C9517 trim[4] comp 6.05e-20
C9518 net15 _141_/a_27_47# 0.00199f
C9519 output22/a_27_47# _004_ 0.00117f
C9520 _005_ net30 5.05e-20
C9521 _133_ cal_count\[2\] 0.308f
C9522 _094_ _092_ 0.105f
C9523 mask\[2\] _017_ 0.0214f
C9524 _319_/a_27_47# clknet_0_clk 0.00149f
C9525 _074_ _212_/a_113_297# 0.0208f
C9526 clkbuf_2_0__f_clk/a_110_47# net3 0.0132f
C9527 _293_/a_81_21# _041_ 0.00233f
C9528 _320_/a_193_47# _319_/a_1283_21# 8.37e-21
C9529 _088_ _092_ 6.57e-20
C9530 _052_ _099_ 1.41e-19
C9531 net44 _206_/a_206_47# 1.57e-19
C9532 _218_/a_199_47# net26 1.86e-19
C9533 _110_ net10 1.95e-20
C9534 VPWR _097_ 0.247f
C9535 _115_ _056_ 4.69e-21
C9536 trim_val\[1\] _175_/a_68_297# 5.65e-19
C9537 net12 _337_/a_1283_21# 8.78e-19
C9538 _167_/a_161_47# clk 0.00238f
C9539 trim_val\[1\] _333_/a_193_47# 4.9e-19
C9540 trim_mask\[1\] _333_/a_27_47# 0.0168f
C9541 _341_/a_193_47# _304_/a_543_47# 9.04e-20
C9542 _101_ _049_ 0.00159f
C9543 VPWR _192_/a_548_47# -5.31e-19
C9544 _071_ VPWR 0.258f
C9545 _110_ clknet_2_2__leaf_clk 1.01f
C9546 net15 _281_/a_253_47# 0.00261f
C9547 net43 _022_ 0.00404f
C9548 output14/a_27_47# net27 2.42e-20
C9549 _340_/a_381_47# net47 1.05e-20
C9550 _037_ _304_/a_1108_47# 7.95e-20
C9551 _315_/a_193_47# valid 0.00582f
C9552 _269_/a_81_21# trim_val\[0\] 2.93e-19
C9553 _005_ net22 0.00141f
C9554 _108_ _279_/a_490_47# 0.00671f
C9555 _048_ _232_/a_32_297# 4.6e-19
C9556 _259_/a_27_297# _335_/a_761_289# 2.67e-19
C9557 _259_/a_109_297# _335_/a_193_47# 4.56e-19
C9558 _008_ mask\[6\] 6.33e-21
C9559 _128_ _127_ 0.0062f
C9560 _308_/a_1217_47# net45 6.07e-20
C9561 VPWR _262_/a_27_47# 0.0714f
C9562 result[2] net14 6.6e-20
C9563 _007_ _310_/a_448_47# 0.0023f
C9564 output26/a_27_47# _310_/a_193_47# 2.68e-19
C9565 _253_/a_81_21# mask\[7\] 0.00126f
C9566 _309_/a_651_413# _078_ 0.00281f
C9567 _110_ net11 2.59e-19
C9568 _117_ net19 5.71e-21
C9569 _144_/a_27_47# _041_ 0.0257f
C9570 _323_/a_193_47# _043_ 7e-20
C9571 _187_/a_27_413# _058_ 1.98e-20
C9572 _167_/a_161_47# net4 0.0473f
C9573 _337_/a_193_47# _121_ 7.28e-19
C9574 _211_/a_109_297# net14 9.08e-19
C9575 VPWR _315_/a_543_47# 0.0319f
C9576 _309_/a_1283_21# net24 0.0733f
C9577 _068_ _190_/a_465_47# 0.00437f
C9578 _337_/a_1283_21# net44 0.0107f
C9579 _230_/a_59_75# clkbuf_2_3__f_clk/a_110_47# 0.0067f
C9580 output28/a_27_47# _011_ 0.00175f
C9581 _309_/a_543_47# net45 1.49e-19
C9582 _182_/a_27_47# _332_/a_1283_21# 0.0125f
C9583 _058_ _332_/a_27_47# 0.00986f
C9584 net43 cal_itt\[3\] 1.33e-20
C9585 _233_/a_109_297# input1/a_75_212# 7.12e-21
C9586 VPWR _318_/a_1217_47# 2.19e-19
C9587 _082_ _310_/a_1283_21# 3.18e-19
C9588 trimb[0] output38/a_27_47# 6.66e-20
C9589 output36/a_27_47# trimb[2] 0.00188f
C9590 _058_ _268_/a_75_212# 0.00368f
C9591 _200_/a_209_297# net19 0.00228f
C9592 net45 _245_/a_27_297# 0.0631f
C9593 _116_ net50 0.00151f
C9594 _117_ trim_mask\[3\] 6.22e-19
C9595 input2/a_27_47# net37 4.62e-20
C9596 _327_/a_448_47# net46 6.52e-19
C9597 _092_ _108_ 7.49e-20
C9598 cal_itt\[1\] _266_/a_68_297# 8.13e-20
C9599 _162_/a_27_47# net34 2.42e-20
C9600 _260_/a_250_297# _049_ 0.0201f
C9601 _048_ _227_/a_209_311# 0.0748f
C9602 _341_/a_27_47# _091_ 0.00191f
C9603 _189_/a_408_47# _050_ 0.00111f
C9604 _028_ _171_/a_27_47# 4.32e-20
C9605 _128_ _126_ 3.32e-19
C9606 state\[2\] _088_ 0.00635f
C9607 ctlp[6] ctlp[7] 0.0358f
C9608 mask\[1\] net51 5.71e-20
C9609 _328_/a_1217_47# VPWR 1.2e-20
C9610 _292_/a_78_199# cal_count\[2\] 1.5e-19
C9611 _071_ _063_ 0.0685f
C9612 calibrate _099_ 4.75e-19
C9613 _093_ _095_ 1.33e-19
C9614 trim_mask\[4\] _227_/a_209_311# 8.9e-21
C9615 _291_/a_285_297# _289_/a_68_297# 6.54e-21
C9616 _308_/a_1108_47# _319_/a_448_47# 4.21e-21
C9617 _136_ _038_ 0.0457f
C9618 _066_ clkbuf_2_3__f_clk/a_110_47# 5.74e-19
C9619 _200_/a_209_297# _107_ 4.95e-20
C9620 VPWR result[2] 0.185f
C9621 _110_ trim_val\[0\] 0.00507f
C9622 net3 _317_/a_27_47# 1.33e-19
C9623 _306_/a_761_289# _076_ 3.26e-20
C9624 _019_ mask\[6\] 1.18e-20
C9625 cal_itt\[0\] _199_/a_193_297# 3.23e-19
C9626 _328_/a_543_47# _025_ 5.66e-19
C9627 _038_ _284_/a_68_297# 0.00282f
C9628 _304_/a_193_47# clknet_2_3__leaf_clk 0.16f
C9629 VPWR _211_/a_109_297# -6.77e-20
C9630 _303_/a_1283_21# fanout47/a_27_47# 0.0139f
C9631 mask\[3\] _247_/a_27_297# 0.113f
C9632 VPWR wire42/a_75_212# 0.0137f
C9633 _262_/a_27_47# _063_ 0.018f
C9634 _078_ _046_ 0.357f
C9635 VPWR cal_count\[2\] 0.297f
C9636 net45 _331_/a_1108_47# 0.0184f
C9637 _326_/a_761_289# result[5] 9.44e-20
C9638 _169_/a_215_311# calibrate 1.25e-21
C9639 _097_ _164_/a_161_47# 0.00108f
C9640 net43 _011_ 1.73e-19
C9641 _325_/a_1108_47# _250_/a_109_297# 7.36e-20
C9642 _321_/a_1283_21# _320_/a_543_47# 1.26e-21
C9643 net25 _146_/a_68_297# 0.0219f
C9644 _325_/a_543_47# _042_ 0.00153f
C9645 _021_ _312_/a_651_413# 6.03e-21
C9646 _340_/a_562_413# _122_ 7.19e-20
C9647 net13 _319_/a_1283_21# 5.1e-19
C9648 _112_ _333_/a_639_47# 6.26e-19
C9649 net49 _333_/a_805_47# 6.71e-19
C9650 _337_/a_761_289# clknet_0_clk 2.53e-20
C9651 net48 _333_/a_761_289# 6.02e-21
C9652 trim_val\[2\] _333_/a_1283_21# 1.8e-20
C9653 net47 _338_/a_1032_413# 0.0296f
C9654 _338_/a_27_47# _338_/a_652_21# -0.00445f
C9655 _293_/a_81_21# _129_ 0.00305f
C9656 cal_count\[1\] _132_ 1.61e-19
C9657 _325_/a_651_413# clknet_2_1__leaf_clk 5.87e-19
C9658 _059_ _228_/a_79_21# 2.24e-19
C9659 output32/a_27_47# output35/a_27_47# 0.003f
C9660 _104_ _335_/a_543_47# 1.71e-19
C9661 _064_ _335_/a_1108_47# 0.00192f
C9662 _322_/a_1108_47# _065_ 3.11e-20
C9663 _340_/a_562_413# _037_ 1.08e-19
C9664 _050_ _170_/a_81_21# 0.0186f
C9665 _327_/a_639_47# _108_ 3.69e-19
C9666 _326_/a_27_47# output14/a_27_47# 4.86e-21
C9667 net23 result[2] 4.23e-19
C9668 _335_/a_27_47# _330_/a_27_47# 9.7e-19
C9669 _053_ _052_ 0.0087f
C9670 _110_ _279_/a_204_297# 0.00536f
C9671 _328_/a_27_47# net50 5.21e-21
C9672 _340_/a_27_47# _129_ 1.16e-20
C9673 result[4] _310_/a_448_47# 6.75e-19
C9674 _000_ _072_ 6.77e-22
C9675 trim_mask\[3\] net9 0.0183f
C9676 _305_/a_448_47# _092_ 4.12e-20
C9677 _061_ net35 0.0122f
C9678 _230_/a_59_75# cal_count\[3\] 3.92e-20
C9679 VPWR _319_/a_193_47# -0.00541f
C9680 _226_/a_303_47# _075_ 2.17e-19
C9681 _074_ mask\[5\] 5.12e-19
C9682 _062_ net40 0.0233f
C9683 _058_ _332_/a_1217_47# 9.77e-20
C9684 _293_/a_81_21# _339_/a_1032_413# 1.08e-19
C9685 trim_mask\[2\] _172_/a_68_297# 1.33e-19
C9686 _012_ input1/a_75_212# 5.56e-21
C9687 _074_ cal 0.00431f
C9688 VPWR _243_/a_109_47# -8.41e-19
C9689 _144_/a_27_47# _129_ 0.00317f
C9690 _320_/a_193_47# _143_/a_68_297# 0.00162f
C9691 _328_/a_27_47# _333_/a_448_47# 1.96e-21
C9692 _328_/a_1108_47# _333_/a_193_47# 6.92e-20
C9693 net15 _314_/a_27_47# 1.97e-21
C9694 net9 _001_ 0.00129f
C9695 trim_mask\[0\] _301_/a_285_47# 1.56e-19
C9696 net31 output35/a_27_47# 0.00667f
C9697 _063_ wire42/a_75_212# 1.25e-20
C9698 VPWR _197_/a_113_297# 0.0204f
C9699 _340_/a_1032_413# _339_/a_27_47# 4.51e-20
C9700 _340_/a_652_21# _339_/a_476_47# 4.14e-22
C9701 _340_/a_1182_261# _339_/a_193_47# 1.55e-19
C9702 _340_/a_476_47# _339_/a_652_21# 4.26e-20
C9703 _340_/a_27_47# _339_/a_1032_413# 2.42e-20
C9704 _168_/a_207_413# _048_ 2.41e-23
C9705 _187_/a_27_413# en_co_clk 0.00525f
C9706 _043_ _303_/a_27_47# 0.00115f
C9707 clk clkbuf_2_2__f_clk/a_110_47# 0.00318f
C9708 clkbuf_0_clk/a_110_47# clknet_0_clk 0.122f
C9709 _136_ _298_/a_292_297# 6.7e-20
C9710 _302_/a_27_297# clknet_2_3__leaf_clk 0.0472f
C9711 _330_/a_1108_47# _027_ 0.0566f
C9712 _330_/a_1283_21# net46 0.058f
C9713 ctlp[0] _314_/a_27_47# 0.00196f
C9714 clkbuf_2_0__f_clk/a_110_47# _281_/a_103_199# 0.0142f
C9715 _066_ cal_count\[3\] 0.0657f
C9716 net43 _319_/a_1283_21# 0.0347f
C9717 net23 _319_/a_193_47# 8.7e-20
C9718 trim[4] net46 5.7e-19
C9719 _168_/a_207_413# trim_mask\[4\] 0.0619f
C9720 _144_/a_27_47# _339_/a_1032_413# 4.27e-19
C9721 VPWR _194_/a_199_47# -2.69e-19
C9722 VPWR _202_/a_79_21# 0.0164f
C9723 net12 _320_/a_27_47# 1.15e-21
C9724 input3/a_75_212# clknet_2_0__leaf_clk 1.56e-19
C9725 VPWR _336_/a_1108_47# 0.0367f
C9726 _328_/a_805_47# clknet_2_2__leaf_clk 2.34e-19
C9727 net31 _125_ 0.00536f
C9728 _106_ clknet_2_3__leaf_clk 4.29e-19
C9729 VPWR _304_/a_543_47# 0.0109f
C9730 net25 _018_ 0.00104f
C9731 _340_/a_1602_47# _133_ 0.00808f
C9732 _107_ _262_/a_109_297# 0.00217f
C9733 _341_/a_761_289# _038_ 0.00104f
C9734 _341_/a_448_47# _136_ 0.00158f
C9735 net45 clknet_2_2__leaf_clk 0.00324f
C9736 output21/a_27_47# net20 6.94e-19
C9737 clknet_2_2__leaf_clk rebuffer3/a_75_212# 9.57e-19
C9738 _270_/a_59_75# _333_/a_27_47# 0.00308f
C9739 net4 clkbuf_2_2__f_clk/a_110_47# 0.214f
C9740 _053_ calibrate 0.145f
C9741 state\[0\] _093_ 0.0554f
C9742 _326_/a_1108_47# net15 2.21e-20
C9743 _325_/a_543_47# _022_ 4.57e-19
C9744 _325_/a_1108_47# _021_ 1.91e-20
C9745 ctlp[6] net44 2.53e-19
C9746 _319_/a_193_47# net52 8.1e-20
C9747 _325_/a_27_47# _078_ 0.0104f
C9748 _082_ _042_ 0.00156f
C9749 net54 _232_/a_32_297# 0.0606f
C9750 _239_/a_694_21# _092_ 0.0334f
C9751 _320_/a_27_47# net44 -7.05e-19
C9752 VPWR _206_/a_27_93# 0.0144f
C9753 clknet_2_2__leaf_clk _065_ 0.00202f
C9754 _187_/a_212_413# net40 0.0142f
C9755 net13 _337_/a_448_47# 0.00342f
C9756 _335_/a_448_47# _330_/a_1108_47# 2.39e-19
C9757 output35/a_27_47# net2 4.69e-19
C9758 _197_/a_113_297# _063_ 0.0474f
C9759 _321_/a_193_47# net53 7.04e-20
C9760 _040_ _337_/a_543_47# 8.12e-20
C9761 _332_/a_193_47# net40 0.0137f
C9762 VPWR _035_ 0.0551f
C9763 _336_/a_543_47# _266_/a_68_297# 1.1e-20
C9764 net31 net40 2.27e-19
C9765 VPWR _319_/a_1462_47# 1.14e-19
C9766 _105_ clknet_2_2__leaf_clk 4.87e-20
C9767 trim_mask\[0\] clknet_2_3__leaf_clk 0.324f
C9768 VPWR _256_/a_27_297# 0.0701f
C9769 ctln[4] _335_/a_27_47# 3.44e-19
C9770 _168_/a_297_47# _050_ 0.00186f
C9771 VPWR _321_/a_543_47# 0.02f
C9772 _323_/a_651_413# net44 5.32e-19
C9773 _320_/a_1283_21# _041_ 1.05e-19
C9774 net2 rebuffer5/a_161_47# 5.89e-19
C9775 _305_/a_543_47# en_co_clk 4.11e-21
C9776 _012_ output30/a_27_47# 1.46e-19
C9777 _333_/a_1283_21# _176_/a_27_47# 1.3e-19
C9778 net47 _339_/a_1602_47# 3.88e-20
C9779 VPWR _337_/a_543_47# 0.0149f
C9780 VPWR _162_/a_27_47# 0.0851f
C9781 net2 _125_ 0.0331f
C9782 _293_/a_81_21# _297_/a_47_47# 2.03e-20
C9783 _323_/a_193_47# _323_/a_1108_47# -0.00656f
C9784 net13 _143_/a_68_297# 9.7e-19
C9785 _189_/a_27_47# en_co_clk 4.84e-21
C9786 _316_/a_761_289# _013_ 3.21e-20
C9787 fanout45/a_27_47# net41 5.27e-20
C9788 _192_/a_505_280# _095_ 0.0569f
C9789 _192_/a_174_21# _092_ 0.00143f
C9790 _192_/a_27_47# _099_ 3.79e-20
C9791 cal_itt\[2\] _092_ 0.0943f
C9792 state\[2\] _170_/a_299_297# 0.00523f
C9793 _090_ _100_ 0.179f
C9794 _089_ net55 3.16e-19
C9795 _065_ _209_/a_27_47# 0.0703f
C9796 _015_ _318_/a_27_47# 0.037f
C9797 VPWR _302_/a_109_47# -0.00104f
C9798 _308_/a_543_47# _006_ 8.48e-20
C9799 _308_/a_1108_47# _081_ 3.75e-21
C9800 clkbuf_2_0__f_clk/a_110_47# _120_ 0.0439f
C9801 _033_ _280_/a_75_212# 0.00207f
C9802 _291_/a_117_297# net33 0.00159f
C9803 mask\[0\] _283_/a_75_212# 4.16e-20
C9804 _104_ trim_mask\[1\] 0.138f
C9805 _306_/a_543_47# _305_/a_193_47# 0.00115f
C9806 _306_/a_1283_21# _305_/a_27_47# 9.58e-19
C9807 _326_/a_543_47# _310_/a_543_47# 1.3e-20
C9808 _326_/a_193_47# _310_/a_1108_47# 4.77e-21
C9809 _326_/a_761_289# _310_/a_1283_21# 1.09e-20
C9810 _323_/a_27_47# net18 6.31e-21
C9811 net13 clk 0.015f
C9812 net43 _321_/a_448_47# 0.0248f
C9813 net47 cal_count\[3\] 9.79e-21
C9814 VPWR fanout45/a_27_47# 0.0604f
C9815 _338_/a_652_21# clknet_2_3__leaf_clk 0.0268f
C9816 output20/a_27_47# _312_/a_543_47# 0.0111f
C9817 _320_/a_193_47# _320_/a_761_289# -0.00517f
C9818 _320_/a_27_47# _320_/a_543_47# -0.0049f
C9819 net13 clone7/a_27_47# 0.00466f
C9820 clknet_2_1__leaf_clk _208_/a_505_21# 0.00601f
C9821 _334_/a_448_47# net46 0.0179f
C9822 _316_/a_27_47# output41/a_27_47# 1.6e-21
C9823 VPWR _340_/a_1602_47# 5.7e-19
C9824 output32/a_27_47# output31/a_27_47# 1.88e-19
C9825 _104_ _170_/a_81_21# 0.0544f
C9826 output24/a_27_47# _007_ 4.85e-19
C9827 net43 _313_/a_761_289# -0.00363f
C9828 _315_/a_27_47# _099_ 1.82e-20
C9829 _315_/a_1108_47# _241_/a_297_47# 2e-20
C9830 _301_/a_47_47# _134_ 0.00864f
C9831 _058_ net30 0.00133f
C9832 mask\[5\] net26 0.00797f
C9833 _336_/a_543_47# _028_ 4.82e-20
C9834 _336_/a_1283_21# clknet_2_2__leaf_clk 0.00137f
C9835 VPWR _253_/a_299_297# 0.0732f
C9836 _035_ _063_ 8.42e-20
C9837 net35 net16 0.0519f
C9838 clknet_2_1__leaf_clk mask\[2\] 0.387f
C9839 net34 _129_ 9.43e-20
C9840 net27 net29 0.284f
C9841 _341_/a_1108_47# _301_/a_285_47# 3.78e-20
C9842 net2 net40 0.0254f
C9843 mask\[3\] mask\[0\] 1.07e-20
C9844 net25 _078_ 0.407f
C9845 _161_/a_68_297# _332_/a_1283_21# 0.00113f
C9846 _327_/a_1283_21# net9 0.0171f
C9847 _321_/a_1108_47# _101_ 0.0581f
C9848 _190_/a_465_47# cal_itt\[3\] 8.18e-20
C9849 _338_/a_956_413# net18 7.18e-19
C9850 output22/a_27_47# _308_/a_27_47# 0.0131f
C9851 net12 _324_/a_193_47# 3.78e-20
C9852 _341_/a_193_47# _341_/a_651_413# -0.00701f
C9853 _341_/a_193_47# net18 0.00307f
C9854 net13 net4 0.00859f
C9855 _320_/a_1217_47# net44 -5.37e-19
C9856 _134_ _299_/a_215_297# 0.00177f
C9857 _036_ _035_ 4.23e-21
C9858 net47 _303_/a_448_47# 3.26e-21
C9859 _337_/a_1108_47# _101_ 1.38e-19
C9860 _337_/a_543_47# net52 3.49e-21
C9861 VPWR output12/a_27_47# 0.129f
C9862 _336_/a_448_47# net19 0.00617f
C9863 _337_/a_27_47# _263_/a_297_47# 1.6e-20
C9864 _032_ _330_/a_1108_47# 0.00731f
C9865 _335_/a_1283_21# net46 0.0892f
C9866 net15 _247_/a_109_297# 0.00362f
C9867 _281_/a_253_297# _049_ 3.38e-21
C9868 _328_/a_1283_21# _058_ 0.0034f
C9869 _321_/a_1462_47# net53 2.16e-19
C9870 _053_ _170_/a_384_47# 1.26e-19
C9871 clk _331_/a_193_47# 0.0195f
C9872 output31/a_27_47# net31 0.0404f
C9873 _199_/a_193_297# _069_ 4.24e-19
C9874 _304_/a_1283_21# _231_/a_161_47# 0.00128f
C9875 _258_/a_27_297# _280_/a_75_212# 0.02f
C9876 net12 _322_/a_27_47# 6.71e-21
C9877 _299_/a_298_297# _129_ 0.0269f
C9878 _299_/a_215_297# _130_ 0.0398f
C9879 _125_ _123_ 1.37e-21
C9880 net51 _062_ 7.83e-21
C9881 net12 _331_/a_27_47# 1.36e-19
C9882 net28 _313_/a_639_47# 0.00432f
C9883 _266_/a_68_297# _106_ 0.0507f
C9884 net44 rebuffer6/a_27_47# 0.00106f
C9885 ctlp[7] net21 0.0261f
C9886 _339_/a_1032_413# net34 4.15e-21
C9887 net50 _336_/a_1108_47# 1.67e-20
C9888 _333_/a_27_47# _173_/a_27_47# 1.35e-20
C9889 _048_ _100_ 0.21f
C9890 ctln[4] _335_/a_1217_47# 6.4e-20
C9891 _324_/a_193_47# net44 0.0216f
C9892 _014_ _095_ 0.118f
C9893 clknet_2_0__leaf_clk _099_ 3.7e-20
C9894 en_co_clk _227_/a_109_93# 2.05e-21
C9895 _332_/a_543_47# net46 0.03f
C9896 net46 _108_ 0.0945f
C9897 net4 _198_/a_27_47# 0.0121f
C9898 _110_ _330_/a_1283_21# 0.0103f
C9899 _051_ _119_ 4.4e-20
C9900 _324_/a_27_47# _323_/a_27_47# 8.63e-20
C9901 VPWR _313_/a_805_47# 3.71e-20
C9902 _336_/a_448_47# _107_ 5.02e-19
C9903 _019_ _321_/a_193_47# 1.38e-19
C9904 _001_ _202_/a_382_297# 1.78e-20
C9905 _307_/a_27_47# _307_/a_1108_47# -2.98e-20
C9906 net4 _331_/a_193_47# 1.66e-19
C9907 net43 clk 0.00926f
C9908 _037_ _339_/a_381_47# 1.56e-19
C9909 _064_ cal_itt\[0\] 2.64e-19
C9910 _050_ _336_/a_27_47# 2.14e-19
C9911 _323_/a_1283_21# clknet_2_3__leaf_clk 7.04e-22
C9912 _298_/a_493_297# _133_ 9.81e-19
C9913 result[0] _307_/a_27_47# 0.0108f
C9914 input1/a_75_212# _315_/a_543_47# 2.16e-20
C9915 _310_/a_193_47# _310_/a_651_413# -0.00701f
C9916 clknet_2_3__leaf_clk _298_/a_78_199# 1.63e-19
C9917 _041_ _040_ 4.32e-20
C9918 _074_ _310_/a_27_47# 0.0175f
C9919 _314_/a_27_47# _224_/a_113_297# 0.00106f
C9920 _322_/a_27_47# net44 0.00469f
C9921 _233_/a_27_297# _074_ 0.0123f
C9922 _046_ _313_/a_1108_47# 6.99e-20
C9923 net21 _313_/a_543_47# 0.00136f
C9924 _128_ net47 0.0987f
C9925 _051_ _331_/a_651_413# 2.87e-19
C9926 state\[2\] _318_/a_651_413# 9.5e-19
C9927 net12 _219_/a_109_297# 4.53e-19
C9928 _301_/a_47_47# cal_count\[3\] 3.02e-19
C9929 _048_ _264_/a_27_297# 0.00146f
C9930 _311_/a_27_47# _311_/a_193_47# -0.0518f
C9931 _303_/a_448_47# net44 4.4e-19
C9932 _231_/a_161_47# _091_ 0.0199f
C9933 _123_ net40 1.12e-20
C9934 output9/a_27_47# _057_ 0.0557f
C9935 _051_ _087_ 0.316f
C9936 net43 net4 2.72e-21
C9937 _097_ _281_/a_253_47# 2.12e-19
C9938 net42 en_co_clk 2.04e-20
C9939 _326_/a_639_47# _074_ 0.00132f
C9940 VPWR _041_ 1.46f
C9941 _341_/a_27_47# cal_count\[3\] 0.0348f
C9942 _302_/a_109_297# clknet_2_2__leaf_clk 5.41e-20
C9943 trim_mask\[0\] _266_/a_68_297# 9.75e-19
C9944 _338_/a_1056_47# clknet_2_3__leaf_clk 2.82e-19
C9945 VPWR _338_/a_1182_261# -0.00497f
C9946 _341_/a_1108_47# clknet_2_3__leaf_clk 0.0465f
C9947 _309_/a_1270_413# _081_ 2.96e-20
C9948 _309_/a_448_47# _006_ 0.0023f
C9949 state\[0\] _192_/a_505_280# 3.6e-21
C9950 _323_/a_1283_21# _303_/a_193_47# 3.34e-19
C9951 _323_/a_543_47# _303_/a_761_289# 4.73e-19
C9952 _323_/a_1108_47# _303_/a_27_47# 4.49e-21
C9953 _031_ net46 0.437f
C9954 trim_mask\[3\] _256_/a_109_297# 1.18e-20
C9955 cal_itt\[0\] _053_ 0.037f
C9956 net50 _256_/a_27_297# 0.00768f
C9957 trim_mask\[1\] _267_/a_59_75# 2.13e-21
C9958 clknet_2_0__leaf_clk _246_/a_27_297# 0.0312f
C9959 _315_/a_1462_47# _095_ 1.1e-19
C9960 _315_/a_1217_47# _099_ 2.14e-20
C9961 _339_/a_193_47# _339_/a_476_47# -0.0164f
C9962 _129_ _133_ 0.106f
C9963 fanout46/a_27_47# _335_/a_543_47# 1.78e-19
C9964 net13 _320_/a_761_289# 0.00446f
C9965 _336_/a_805_47# trim_mask\[4\] 0.00213f
C9966 _322_/a_1283_21# _041_ 7.76e-20
C9967 _306_/a_448_47# clknet_2_1__leaf_clk 2.39e-19
C9968 _264_/a_27_297# trim_mask\[4\] 5.68e-19
C9969 _187_/a_27_413# _061_ 0.00275f
C9970 _243_/a_27_297# _095_ 8.62e-21
C9971 _091_ _107_ 0.00135f
C9972 _271_/a_75_212# _113_ 0.0232f
C9973 clknet_2_1__leaf_clk _314_/a_193_47# 0.0234f
C9974 _307_/a_27_47# net14 0.0096f
C9975 _336_/a_543_47# _279_/a_314_297# 5.26e-20
C9976 _326_/a_27_47# net29 1.88e-19
C9977 VPWR _316_/a_651_413# 2.6e-19
C9978 mask\[7\] _046_ 0.00373f
C9979 net47 _000_ 0.00782f
C9980 _332_/a_448_47# _108_ 0.0154f
C9981 trim[3] net33 0.00119f
C9982 _033_ net19 0.00928f
C9983 _029_ _332_/a_1283_21# 1.04e-20
C9984 _337_/a_1283_21# _107_ 2.03e-19
C9985 _050_ _096_ 0.0653f
C9986 net15 _018_ 0.00157f
C9987 _146_/a_68_297# _310_/a_193_47# 2.8e-20
C9988 net43 _073_ 1.23e-19
C9989 _182_/a_27_47# net33 0.00559f
C9990 _111_ _029_ 0.0058f
C9991 fanout43/a_27_47# mask\[0\] 0.00867f
C9992 en_co_clk net30 0.00826f
C9993 _339_/a_1032_413# _133_ 7.58e-21
C9994 clk _260_/a_93_21# 2.46e-19
C9995 trim_mask\[3\] _033_ 4.38e-20
C9996 net12 net21 2.37e-20
C9997 _333_/a_1108_47# net32 5.89e-19
C9998 _324_/a_1462_47# net44 3.49e-19
C9999 _200_/a_209_297# _062_ 0.00129f
C10000 net7 _317_/a_193_47# 1.8e-20
C10001 net15 _317_/a_543_47# 0.00815f
C10002 _333_/a_27_47# _172_/a_68_297# 3.35e-19
C10003 net43 _214_/a_199_47# 1.37e-20
C10004 _104_ _255_/a_27_47# 3.79e-19
C10005 _041_ net52 0.00218f
C10006 input2/a_27_47# cal_count\[2\] 9.26e-21
C10007 _041_ _063_ 1.61e-20
C10008 _033_ _107_ 0.00183f
C10009 _306_/a_543_47# _049_ 3.01e-20
C10010 _326_/a_448_47# clknet_2_1__leaf_clk 0.00313f
C10011 _308_/a_1108_47# net14 4.01e-19
C10012 net4 _260_/a_93_21# 7.28e-20
C10013 _306_/a_193_47# net30 2.7e-20
C10014 comp output5/a_27_47# 0.00409f
C10015 VPWR _323_/a_448_47# -0.00161f
C10016 VPWR _307_/a_27_47# 0.0688f
C10017 cal _315_/a_805_47# 4.66e-20
C10018 _290_/a_27_413# net37 3.35e-19
C10019 output31/a_27_47# trim_val\[1\] 0.00829f
C10020 trim[0] _269_/a_81_21# 1.8e-19
C10021 VPWR _298_/a_493_297# -2.93e-19
C10022 state\[0\] _014_ 1.06e-20
C10023 _314_/a_448_47# net29 8.96e-20
C10024 _322_/a_1217_47# net44 8.76e-19
C10025 _300_/a_47_47# _135_ 0.00613f
C10026 _300_/a_285_47# net2 0.00153f
C10027 _329_/a_193_47# _026_ 0.0104f
C10028 output38/a_27_47# net39 0.0374f
C10029 _329_/a_193_47# VPWR 0.045f
C10030 calibrate _093_ 1.33f
C10031 _110_ _334_/a_448_47# 1.14e-20
C10032 _305_/a_27_47# net2 1.9e-19
C10033 net43 _320_/a_761_289# 2.8e-19
C10034 _036_ _041_ 0.00246f
C10035 _335_/a_1108_47# _032_ 1.92e-19
C10036 _214_/a_113_297# _101_ 0.00483f
C10037 net12 _242_/a_297_47# 4.52e-19
C10038 _325_/a_448_47# _321_/a_543_47# 1.3e-20
C10039 _313_/a_27_47# _155_/a_68_297# 3.73e-21
C10040 _305_/a_27_47# _305_/a_1283_21# -9.15e-20
C10041 _305_/a_193_47# _305_/a_543_47# -0.0113f
C10042 _299_/a_298_297# _297_/a_47_47# 5.42e-19
C10043 en_co_clk _072_ 1.19e-19
C10044 _000_ net44 0.024f
C10045 _325_/a_761_289# _313_/a_543_47# 4.07e-20
C10046 _325_/a_543_47# _313_/a_761_289# 3.29e-20
C10047 _038_ clknet_2_2__leaf_clk 1.8e-20
C10048 _272_/a_81_21# net46 0.00853f
C10049 net49 net46 0.0204f
C10050 _306_/a_27_47# mask\[0\] 4.4e-20
C10051 net44 _312_/a_1283_21# 0.00854f
C10052 VPWR net18 1.12f
C10053 VPWR _341_/a_651_413# -0.00947f
C10054 trim_val\[3\] _258_/a_109_297# 3.19e-20
C10055 trim_mask\[3\] _258_/a_27_297# 0.00419f
C10056 _320_/a_193_47# _101_ 3.1e-20
C10057 _303_/a_543_47# clknet_2_3__leaf_clk 0.0335f
C10058 net2 net51 0.0602f
C10059 net45 mask\[2\] 6.57e-20
C10060 _116_ _335_/a_543_47# 0.00144f
C10061 _117_ _335_/a_761_289# 0.00241f
C10062 _110_ _335_/a_1283_21# 3.09e-19
C10063 VPWR _129_ 0.366f
C10064 _309_/a_1108_47# _140_/a_68_297# 1.48e-19
C10065 _321_/a_1108_47# _248_/a_27_297# 7.15e-19
C10066 net43 _307_/a_543_47# 1.29e-20
C10067 _114_ _334_/a_27_47# 8.99e-20
C10068 trim_val\[2\] _334_/a_543_47# 0.00627f
C10069 net48 _334_/a_193_47# 6.36e-19
C10070 _076_ cal_itt\[3\] 1.53e-20
C10071 _320_/a_805_47# _040_ 0.00239f
C10072 net55 _092_ 0.222f
C10073 VPWR _308_/a_1108_47# 0.0361f
C10074 _307_/a_1217_47# net14 2.97e-20
C10075 _024_ _107_ 6.14e-21
C10076 mask\[0\] sample 1.96e-19
C10077 _306_/a_761_289# cal_itt\[3\] 3.97e-19
C10078 _306_/a_193_47# _072_ 3.02e-19
C10079 _065_ _208_/a_505_21# 0.0389f
C10080 _337_/a_27_47# _099_ 8.76e-22
C10081 _337_/a_193_47# _095_ 0.00207f
C10082 _106_ _279_/a_314_297# 3.92e-19
C10083 clk net3 0.00563f
C10084 _083_ _041_ 3.53e-21
C10085 _292_/a_78_199# _339_/a_1032_413# 0.00155f
C10086 _228_/a_297_47# _054_ 7.75e-20
C10087 result[5] _011_ 5.91e-19
C10088 net3 clone7/a_27_47# 1.92e-20
C10089 _052_ _171_/a_27_47# 4.28e-20
C10090 _110_ _332_/a_543_47# 1.5e-20
C10091 mask\[2\] _065_ 1.79e-20
C10092 _071_ _306_/a_1108_47# 1.73e-20
C10093 _110_ _108_ 0.0421f
C10094 VPWR _237_/a_76_199# 0.00494f
C10095 net26 _310_/a_27_47# 1.7e-19
C10096 rebuffer3/a_75_212# _278_/a_27_47# 2.1e-20
C10097 _042_ _310_/a_1283_21# 2.13e-19
C10098 _303_/a_193_47# _303_/a_543_47# -0.0102f
C10099 _239_/a_277_297# _052_ 2.72e-19
C10100 _169_/a_109_53# net55 1.7e-20
C10101 _325_/a_27_47# mask\[7\] 6.45e-19
C10102 VPWR _320_/a_805_47# 4.48e-19
C10103 state\[0\] _243_/a_27_297# 0.0209f
C10104 _058_ _066_ 0.00225f
C10105 net54 _100_ 0.0442f
C10106 VPWR _339_/a_1032_413# 0.0246f
C10107 output33/a_27_47# net37 6.98e-21
C10108 _181_/a_68_297# _033_ 3.76e-22
C10109 _104_ _336_/a_27_47# 0.267f
C10110 clknet_2_1__leaf_clk _310_/a_1270_413# 6.5e-19
C10111 _074_ clknet_2_1__leaf_clk 0.473f
C10112 ctlp[7] _045_ 0.0227f
C10113 _067_ _092_ 0.0862f
C10114 net15 _078_ 0.00631f
C10115 _133_ _297_/a_47_47# 0.00514f
C10116 net3 net4 0.416f
C10117 _300_/a_285_47# _123_ 1.36e-19
C10118 net34 _175_/a_68_297# 0.00256f
C10119 output14/a_27_47# _086_ 0.00109f
C10120 _333_/a_543_47# _055_ 1.88e-20
C10121 net34 _333_/a_193_47# 2.12e-20
C10122 net13 _322_/a_761_289# 9.37e-19
C10123 _319_/a_27_47# mask\[2\] 7.21e-21
C10124 _308_/a_1108_47# net23 1e-18
C10125 trim_mask\[2\] clknet_2_2__leaf_clk 0.59f
C10126 ctlp[6] net19 1.79e-21
C10127 _238_/a_75_212# _233_/a_27_297# 5.09e-20
C10128 _337_/a_543_47# _034_ 0.00135f
C10129 _242_/a_79_21# _098_ 0.0614f
C10130 _063_ net18 2.7e-19
C10131 VPWR _324_/a_27_47# 0.0402f
C10132 net43 _138_/a_27_47# 0.0341f
C10133 _338_/a_1032_413# _001_ 2.61e-19
C10134 VPWR _307_/a_1217_47# 5.67e-20
C10135 _105_ _278_/a_27_47# 8.14e-20
C10136 _091_ _118_ 1.49e-21
C10137 cal_count\[1\] _134_ 2.26e-21
C10138 _329_/a_1462_47# VPWR 2.5e-19
C10139 _309_/a_27_47# net43 0.00681f
C10140 _256_/a_109_297# _118_ 5.6e-20
C10141 _024_ _279_/a_27_47# 1.08e-20
C10142 trim_mask\[0\] _279_/a_314_297# 0.0472f
C10143 _187_/a_27_413# net16 0.0078f
C10144 _110_ _031_ 0.188f
C10145 _053_ _304_/a_27_47# 0.0108f
C10146 _257_/a_27_297# _280_/a_75_212# 1.85e-19
C10147 state\[2\] net55 0.0104f
C10148 cal_itt\[1\] _195_/a_535_374# 1.1e-19
C10149 cal_itt\[0\] _195_/a_218_47# 2.23e-19
C10150 net16 _332_/a_27_47# 0.0122f
C10151 _053_ clone1/a_27_47# 0.0101f
C10152 _329_/a_27_47# clknet_2_2__leaf_clk 0.032f
C10153 clknet_2_1__leaf_clk _247_/a_109_47# 3.7e-19
C10154 net16 _268_/a_75_212# 1.21e-20
C10155 _057_ net33 4.43e-21
C10156 _311_/a_761_289# net26 0.0191f
C10157 cal_count\[1\] _130_ 0.00126f
C10158 output15/a_27_47# _074_ 3.47e-20
C10159 _322_/a_193_47# _322_/a_761_289# -0.0133f
C10160 _322_/a_27_47# _322_/a_543_47# -0.00157f
C10161 _024_ _181_/a_68_297# 9.19e-21
C10162 _305_/a_448_47# clknet_2_1__leaf_clk 4.84e-20
C10163 _331_/a_193_47# _331_/a_761_289# -0.00609f
C10164 _331_/a_27_47# _331_/a_543_47# -0.00297f
C10165 _306_/a_448_47# net45 4.42e-22
C10166 VPWR _303_/a_1108_47# 0.0034f
C10167 _078_ _314_/a_1108_47# 7.59e-21
C10168 calibrate _171_/a_27_47# 1.26e-19
C10169 _269_/a_299_297# trim_mask\[1\] 0.00102f
C10170 _269_/a_81_21# net49 7.82e-20
C10171 _269_/a_384_47# trim_val\[1\] 1.99e-19
C10172 _146_/a_150_297# clknet_2_1__leaf_clk 0.00154f
C10173 VPWR output25/a_27_47# 0.0718f
C10174 _323_/a_651_413# net19 0.00193f
C10175 net13 _101_ 0.0171f
C10176 _239_/a_277_297# calibrate 0.003f
C10177 _058_ _047_ 2.25e-19
C10178 clkbuf_2_3__f_clk/a_110_47# net19 0.018f
C10179 net9 _332_/a_193_47# 2.35e-19
C10180 trim[1] output33/a_27_47# 7.46e-20
C10181 _115_ clknet_2_2__leaf_clk 8.04e-20
C10182 _015_ fanout45/a_27_47# 6.02e-20
C10183 cal_count\[1\] _339_/a_1602_47# 0.026f
C10184 _036_ _339_/a_1032_413# 2.02e-20
C10185 _237_/a_76_199# _164_/a_161_47# 5.85e-19
C10186 _319_/a_1108_47# en_co_clk 3.26e-22
C10187 _230_/a_59_75# en_co_clk 0.0101f
C10188 _329_/a_761_289# trim_mask\[3\] 8.85e-19
C10189 _329_/a_193_47# net50 3.78e-20
C10190 _224_/a_199_47# net29 5.38e-19
C10191 _051_ _099_ 0.012f
C10192 _306_/a_448_47# _065_ 2.9e-20
C10193 _336_/a_1283_21# _278_/a_27_47# 2.4e-21
C10194 _078_ _310_/a_193_47# 0.00812f
C10195 VPWR _309_/a_1270_413# 2.37e-19
C10196 _186_/a_109_297# _100_ 0.00279f
C10197 _291_/a_285_297# trimb[1] 5.07e-19
C10198 _277_/a_75_212# net46 0.00127f
C10199 mask\[7\] net25 4.43e-19
C10200 _127_ cal_count\[0\] 0.0648f
C10201 _093_ _317_/a_1108_47# 8.22e-22
C10202 VPWR _191_/a_27_297# 0.118f
C10203 _107_ clkbuf_2_3__f_clk/a_110_47# 0.0141f
C10204 _001_ _298_/a_215_47# 2.78e-21
C10205 _336_/a_1283_21# _330_/a_1283_21# 7.1e-20
C10206 _188_/a_27_47# _161_/a_68_297# 1.06e-20
C10207 _053_ _069_ 0.00188f
C10208 net30 _039_ 9.56e-19
C10209 _169_/a_215_311# _051_ 0.0381f
C10210 net50 net18 1.09f
C10211 net12 _249_/a_109_297# 0.00238f
C10212 _328_/a_193_47# _113_ 8.33e-20
C10213 _328_/a_1108_47# _271_/a_75_212# 4.38e-19
C10214 _328_/a_27_47# _030_ 2.88e-20
C10215 _322_/a_193_47# _101_ 0.0138f
C10216 VPWR _297_/a_47_47# 0.0587f
C10217 net47 mask\[4\] 0.242f
C10218 _187_/a_212_413# _132_ 8.94e-20
C10219 _094_ net45 1.73e-20
C10220 _237_/a_439_47# _090_ 5.52e-19
C10221 net9 _113_ 3.21e-20
C10222 net4 _190_/a_465_47# 1.89e-21
C10223 _305_/a_193_47# net30 1.22e-19
C10224 _321_/a_761_289# mask\[2\] 2.7e-19
C10225 VPWR _324_/a_1217_47# 1.16e-19
C10226 en_co_clk _066_ 2.69e-21
C10227 _093_ _192_/a_27_47# 1.76e-20
C10228 _189_/a_27_47# _049_ 4.05e-19
C10229 net31 _132_ 0.00487f
C10230 _110_ _272_/a_81_21# 4.04e-19
C10231 _303_/a_1108_47# _063_ 1.29e-21
C10232 _110_ net49 8.81e-19
C10233 mask\[3\] _081_ 2.32e-20
C10234 clkbuf_2_1__f_clk/a_110_47# _049_ 0.00147f
C10235 _068_ cal_itt\[3\] 3.49e-19
C10236 output8/a_27_47# _334_/a_1283_21# 9.9e-19
C10237 net8 _334_/a_27_47# 0.013f
C10238 _293_/a_81_21# _125_ 0.0586f
C10239 net28 _046_ 0.389f
C10240 _309_/a_1217_47# net43 -3.08e-19
C10241 _024_ _118_ 1.14e-20
C10242 _126_ cal_count\[0\] 0.147f
C10243 net22 _039_ 0.399f
C10244 _327_/a_651_413# trim_mask\[0\] 2.51e-19
C10245 _327_/a_1283_21# _024_ 2.09e-19
C10246 _295_/a_113_47# cal_count\[2\] 5.18e-19
C10247 _090_ net41 0.00615f
C10248 net44 _045_ 2.82e-20
C10249 net43 _101_ 0.139f
C10250 _094_ _065_ 0.191f
C10251 _316_/a_1283_21# _099_ 5.48e-21
C10252 net44 _249_/a_109_297# 2.66e-20
C10253 _305_/a_639_47# _002_ 0.00467f
C10254 net16 _332_/a_1217_47# 1.59e-19
C10255 _103_ _088_ 0.121f
C10256 _316_/a_1108_47# _095_ 9.99e-20
C10257 _053_ _340_/a_476_47# 5.85e-20
C10258 _218_/a_199_47# net53 4.92e-21
C10259 VPWR _322_/a_805_47# 2.57e-19
C10260 net9 net2 0.0285f
C10261 VPWR _331_/a_805_47# 5.66e-20
C10262 net12 mask\[4\] 0.105f
C10263 _050_ _098_ 0.115f
C10264 _312_/a_193_47# net20 0.0347f
C10265 _078_ _311_/a_543_47# 4.13e-20
C10266 _312_/a_193_47# net53 5.31e-20
C10267 calibrate _315_/a_193_47# 0.259f
C10268 _093_ _315_/a_27_47# 8.32e-20
C10269 _074_ _315_/a_761_289# 0.00545f
C10270 cal_itt\[0\] _285_/a_113_47# 6.84e-20
C10271 _002_ clknet_2_1__leaf_clk 0.00753f
C10272 _324_/a_1283_21# _312_/a_1283_21# 9.77e-20
C10273 _324_/a_543_47# _312_/a_1108_47# 4.48e-20
C10274 _161_/a_68_297# net33 0.00612f
C10275 VPWR _090_ 1.02f
C10276 _324_/a_193_47# net19 5.02e-19
C10277 _059_ _206_/a_27_93# 0.00252f
C10278 _331_/a_761_289# _260_/a_93_21# 7.97e-21
C10279 clknet_2_1__leaf_clk net26 0.105f
C10280 net12 _220_/a_199_47# 2.76e-19
C10281 _050_ clknet_0_clk 0.783f
C10282 _191_/a_27_297# _063_ -2.53e-20
C10283 _327_/a_805_47# _136_ 1.89e-19
C10284 _327_/a_448_47# _038_ 2.76e-19
C10285 _159_/a_27_47# _046_ 0.0167f
C10286 VPWR _312_/a_543_47# -6.39e-19
C10287 net15 _319_/a_651_413# 0.00187f
C10288 _094_ _319_/a_27_47# 3.12e-21
C10289 cal_count\[3\] net19 0.00666f
C10290 _144_/a_27_47# _125_ 0.00216f
C10291 net12 _060_ 2.45e-20
C10292 _320_/a_27_47# mask\[1\] 0.00683f
C10293 _305_/a_193_47# _072_ 0.134f
C10294 mask\[0\] net51 6.26e-20
C10295 _311_/a_1108_47# _072_ 2.67e-20
C10296 _231_/a_161_47# cal_count\[3\] 0.0022f
C10297 _064_ _051_ 0.00148f
C10298 _108_ rebuffer3/a_75_212# 0.0427f
C10299 net47 _020_ 0.00425f
C10300 _121_ _092_ 1.03e-21
C10301 _235_/a_79_21# _096_ 0.00268f
C10302 net15 _096_ 0.00182f
C10303 net44 mask\[4\] 0.42f
C10304 net27 _313_/a_1283_21# 1.17e-20
C10305 net45 _244_/a_27_297# 6.53e-19
C10306 _071_ _305_/a_1108_47# 2.83e-19
C10307 _293_/a_81_21# net40 0.00278f
C10308 _237_/a_439_47# _048_ 3.71e-19
C10309 _331_/a_27_47# net19 0.00294f
C10310 trim[1] _270_/a_59_75# 2.55e-20
C10311 VPWR _242_/a_382_297# -0.00102f
C10312 _228_/a_382_297# _100_ 6.54e-20
C10313 _237_/a_535_374# net3 2.81e-19
C10314 _078_ _310_/a_1462_47# 2.33e-19
C10315 _264_/a_27_297# net40 1.87e-19
C10316 _303_/a_639_47# _000_ 9.32e-19
C10317 _309_/a_27_47# _080_ 5.04e-20
C10318 net2 _132_ 0.00922f
C10319 _058_ _301_/a_47_47# 2.94e-19
C10320 _059_ _337_/a_543_47# 4.42e-20
C10321 _093_ clknet_2_0__leaf_clk 0.0107f
C10322 net37 clkc 5.01e-19
C10323 trim_mask\[3\] _257_/a_27_297# 3.91e-19
C10324 _074_ net45 0.0117f
C10325 _337_/a_651_413# en_co_clk 1.93e-19
C10326 calibrate _014_ 0.00963f
C10327 _303_/a_448_47# net19 0.0028f
C10328 _107_ cal_count\[3\] 0.00455f
C10329 _065_ _108_ 8.54e-20
C10330 _128_ cal_count\[1\] 0.18f
C10331 _001_ cal_count\[3\] 3.63e-20
C10332 _336_/a_193_47# net46 -0.00219f
C10333 _328_/a_27_47# trim_mask\[1\] 0.0505f
C10334 _065_ _244_/a_27_297# 0.00484f
C10335 _048_ net41 2.36e-19
C10336 VPWR _175_/a_68_297# -0.00333f
C10337 _053_ _051_ 0.0391f
C10338 cal _316_/a_543_47# 5.95e-20
C10339 _227_/a_109_93# _049_ 0.00546f
C10340 net12 _020_ 5.58e-20
C10341 VPWR _333_/a_193_47# 0.0558f
C10342 fanout47/a_27_47# _124_ 2.13e-19
C10343 clkbuf_2_2__f_clk/a_110_47# trim_val\[4\] 1.41e-19
C10344 _341_/a_543_47# _092_ 4.93e-21
C10345 VPWR _265_/a_81_21# 0.0399f
C10346 _075_ _206_/a_27_93# 0.0152f
C10347 _078_ _224_/a_113_297# 0.0024f
C10348 _144_/a_27_47# net40 2.09e-19
C10349 net9 _123_ 0.0156f
C10350 _337_/a_448_47# _076_ 3.97e-20
C10351 _320_/a_1283_21# mask\[3\] 4.04e-19
C10352 _336_/a_543_47# _052_ 1.55e-20
C10353 _074_ _065_ 0.0445f
C10354 VPWR _048_ 1.2f
C10355 net8 _334_/a_1217_47# 5.59e-19
C10356 _325_/a_1283_21# net13 0.0175f
C10357 net47 en_co_clk 1.35e-19
C10358 clk _330_/a_27_47# 0.00365f
C10359 _053_ _338_/a_193_47# 1.27e-21
C10360 _091_ _062_ 0.00153f
C10361 net44 _020_ 0.0153f
C10362 _251_/a_109_297# _022_ 8.39e-19
C10363 _325_/a_27_47# net28 9.8e-20
C10364 _026_ trim_mask\[4\] 1.16e-19
C10365 output23/a_27_47# net45 6.32e-21
C10366 VPWR trim_mask\[4\] 0.879f
C10367 _312_/a_1462_47# net20 1.27e-19
C10368 _250_/a_27_297# _078_ 0.00401f
C10369 net42 _049_ 0.0459f
C10370 _164_/a_161_47# _090_ 0.00462f
C10371 _337_/a_1283_21# _062_ 4.43e-19
C10372 clkbuf_2_3__f_clk/a_110_47# _118_ 2.47e-19
C10373 _331_/a_639_47# clknet_2_2__leaf_clk 2.44e-19
C10374 _331_/a_1283_21# trim_mask\[4\] 0.0295f
C10375 _260_/a_93_21# _260_/a_250_297# -6.97e-22
C10376 net13 _248_/a_27_297# 0.0128f
C10377 VPWR _325_/a_193_47# 0.0247f
C10378 calibrate _243_/a_27_297# 0.0313f
C10379 state\[0\] _316_/a_1108_47# 0.00218f
C10380 net4 _330_/a_27_47# 2.28e-19
C10381 trim_val\[2\] net48 0.0604f
C10382 net12 en_co_clk 0.013f
C10383 _332_/a_1108_47# net33 1.36e-19
C10384 _194_/a_113_297# _108_ 5.02e-19
C10385 _110_ _277_/a_75_212# 0.0273f
C10386 _123_ _132_ 9.06e-21
C10387 _321_/a_639_47# net15 1.49e-19
C10388 _325_/a_1283_21# _322_/a_193_47# 1.15e-20
C10389 _336_/a_1283_21# _108_ 0.00369f
C10390 _325_/a_27_47# _159_/a_27_47# 4.34e-20
C10391 _181_/a_68_297# cal_count\[3\] 1.25e-21
C10392 net48 net16 0.22f
C10393 _094_ _337_/a_761_289# 0.0133f
C10394 _327_/a_1108_47# net18 5.62e-19
C10395 _253_/a_81_21# _314_/a_193_47# 2.75e-22
C10396 _323_/a_805_47# mask\[4\] 2.83e-19
C10397 _287_/a_75_212# _124_ 0.0642f
C10398 _035_ _286_/a_218_47# 6.37e-20
C10399 _049_ _054_ 0.243f
C10400 _323_/a_27_47# net27 4.72e-19
C10401 _127_ net16 0.00342f
C10402 _318_/a_193_47# _318_/a_1108_47# -0.00656f
C10403 net30 _049_ 0.0182f
C10404 output10/a_27_47# trim_val\[3\] 0.0101f
C10405 net36 net38 0.0522f
C10406 _306_/a_761_289# clk 6.33e-21
C10407 clknet_2_3__leaf_clk _092_ 0.0956f
C10408 _048_ _063_ 0.268f
C10409 _007_ net14 7.62e-19
C10410 output35/a_27_47# net34 0.018f
C10411 net12 _306_/a_193_47# 0.0173f
C10412 net44 en_co_clk 0.164f
C10413 _000_ net19 0.0338f
C10414 _086_ net29 0.0497f
C10415 _136_ _267_/a_59_75# 7.02e-19
C10416 _012_ _004_ 0.00219f
C10417 _322_/a_193_47# _248_/a_27_297# 3.05e-19
C10418 _325_/a_1283_21# net43 -0.00626f
C10419 _312_/a_1283_21# net19 0.00166f
C10420 _322_/a_27_47# _248_/a_109_297# 2.38e-19
C10421 _336_/a_1462_47# net46 -9.14e-19
C10422 _168_/a_27_413# _049_ 1.45e-19
C10423 _195_/a_439_47# _067_ 0.00112f
C10424 VPWR _333_/a_1462_47# 8.45e-20
C10425 cal_itt\[1\] _203_/a_59_75# 5.31e-20
C10426 mask\[3\] net14 2.84e-21
C10427 trim_mask\[4\] _063_ 1.61e-20
C10428 net20 _152_/a_68_297# 1.58e-20
C10429 _110_ _270_/a_145_75# 0.00123f
C10430 cal_itt\[0\] cal_itt\[1\] 0.632f
C10431 net22 _049_ 2.83e-19
C10432 _309_/a_761_289# mask\[3\] 9.58e-19
C10433 _309_/a_543_47# net25 3.39e-19
C10434 _309_/a_27_47# _082_ 5.57e-20
C10435 _104_ _098_ 8.66e-21
C10436 _322_/a_27_47# mask\[1\] 2.06e-20
C10437 _164_/a_161_47# _048_ 0.014f
C10438 _333_/a_27_47# clknet_2_2__leaf_clk 0.00154f
C10439 _050_ _331_/a_1108_47# 7.7e-19
C10440 _140_/a_68_297# _246_/a_27_297# 7.2e-21
C10441 output32/a_27_47# net32 0.0423f
C10442 trim[1] _173_/a_27_47# 0.00392f
C10443 clkbuf_2_1__f_clk/a_110_47# _319_/a_543_47# 0.0132f
C10444 _125_ net34 0.0132f
C10445 input2/a_27_47# _129_ 3.05e-19
C10446 _305_/a_1108_47# _197_/a_113_297# 8.6e-23
C10447 _301_/a_47_47# en_co_clk 0.00143f
C10448 _325_/a_193_47# net52 5.69e-20
C10449 _325_/a_543_47# _101_ 2.6e-19
C10450 net16 _126_ 0.00142f
C10451 mask\[7\] net15 0.0158f
C10452 net42 _262_/a_193_297# 0.0041f
C10453 _306_/a_193_47# net44 0.00297f
C10454 en_co_clk _003_ 9.3e-20
C10455 clkbuf_2_0__f_clk/a_110_47# _319_/a_1283_21# 0.00124f
C10456 net43 _248_/a_27_297# 8.88e-19
C10457 VPWR _283_/a_75_212# 0.0332f
C10458 _341_/a_27_47# en_co_clk 2.39e-19
C10459 _104_ clknet_0_clk 0.0857f
C10460 mask\[3\] _040_ 3.21e-20
C10461 VPWR _190_/a_27_47# 0.0272f
C10462 clkbuf_2_2__f_clk/a_110_47# _330_/a_193_47# 0.0169f
C10463 trim[2] _114_ 9.22e-20
C10464 net47 _286_/a_76_199# 2.22e-19
C10465 _049_ _072_ 1.81e-20
C10466 _328_/a_27_47# _328_/a_448_47# -0.00297f
C10467 _328_/a_193_47# _328_/a_1108_47# -0.00656f
C10468 VPWR _007_ 0.458f
C10469 net2 _202_/a_382_297# 7.04e-20
C10470 _305_/a_1108_47# _202_/a_79_21# 6.84e-19
C10471 _005_ mask\[1\] 2.2e-19
C10472 _210_/a_199_47# _078_ 0.00106f
C10473 _328_/a_1108_47# net9 0.0101f
C10474 _239_/a_694_21# _103_ 4.25e-20
C10475 _107_ _242_/a_297_47# 0.00311f
C10476 _076_ _073_ 7.03e-20
C10477 VPWR _249_/a_27_297# 0.0375f
C10478 _193_/a_109_297# net18 6.37e-19
C10479 _296_/a_113_47# _132_ 1.07e-19
C10480 cal_count\[3\] _118_ 0.0221f
C10481 net12 _228_/a_297_47# 8.49e-19
C10482 net31 net32 0.0992f
C10483 trim_mask\[4\] _260_/a_346_47# 3.96e-19
C10484 _327_/a_639_47# clknet_2_3__leaf_clk 3.69e-20
C10485 VPWR _327_/a_27_47# 0.0789f
C10486 _026_ _327_/a_27_47# 2.01e-20
C10487 _136_ net37 2.66e-20
C10488 VPWR _325_/a_1462_47# 1.68e-19
C10489 _306_/a_193_47# _003_ 0.00324f
C10490 _307_/a_27_47# output30/a_27_47# 0.0123f
C10491 VPWR mask\[3\] 1.56f
C10492 _302_/a_109_297# _108_ 9.02e-19
C10493 _317_/a_1108_47# _014_ 5.47e-21
C10494 _317_/a_193_47# state\[1\] 1.09e-20
C10495 _317_/a_448_47# clknet_2_0__leaf_clk 0.017f
C10496 _317_/a_1283_21# net45 0.0584f
C10497 mask\[5\] _153_/a_27_47# 0.00284f
C10498 _103_ _227_/a_368_53# 2.7e-19
C10499 _322_/a_1283_21# _249_/a_27_297# 1.05e-20
C10500 _237_/a_76_199# _281_/a_253_47# 9.7e-19
C10501 net21 _155_/a_68_297# 0.00231f
C10502 _262_/a_193_297# net30 6.47e-19
C10503 _315_/a_27_47# _315_/a_193_47# -0.0189f
C10504 _212_/a_113_297# _016_ 5.52e-20
C10505 net34 net40 0.002f
C10506 _322_/a_1283_21# mask\[3\] 0.041f
C10507 _058_ _280_/a_75_212# 1.64e-19
C10508 _307_/a_1108_47# fanout43/a_27_47# 4.94e-22
C10509 _050_ _263_/a_79_21# 5.24e-20
C10510 output25/a_27_47# output26/a_27_47# 5.69e-19
C10511 _002_ _065_ 0.0293f
C10512 _325_/a_651_413# _046_ 4.66e-20
C10513 _325_/a_1108_47# net21 0.00558f
C10514 trim_mask\[0\] _052_ 1.94e-25
C10515 _094_ _282_/a_68_297# 0.0449f
C10516 _110_ _336_/a_193_47# 0.0134f
C10517 _065_ net26 2.68e-20
C10518 _259_/a_27_297# _026_ 3.79e-20
C10519 _259_/a_27_297# VPWR 0.0883f
C10520 clk _335_/a_27_47# 1.35e-21
C10521 mask\[7\] _314_/a_1108_47# 8.56e-19
C10522 _238_/a_75_212# net45 0.0324f
C10523 net23 _007_ 3.02e-20
C10524 fanout44/a_27_47# _101_ 8.89e-19
C10525 clknet_2_0__leaf_clk _192_/a_505_280# 1.98e-21
C10526 comp trimb[4] 0.0482f
C10527 trim_val\[0\] _333_/a_27_47# 2.17e-20
C10528 net18 _278_/a_109_297# 1.3e-20
C10529 result[3] net25 0.00318f
C10530 net54 net41 0.407f
C10531 result[4] net14 8.01e-20
C10532 net12 _306_/a_1462_47# 1.18e-19
C10533 net50 trim_mask\[4\] 0.0786f
C10534 _320_/a_761_289# _076_ 3.49e-21
C10535 _320_/a_193_47# _077_ 0.00176f
C10536 _299_/a_298_297# net40 0.00128f
C10537 net23 mask\[3\] 2.04e-20
C10538 _334_/a_27_47# net34 2.68e-20
C10539 _320_/a_448_47# _017_ 0.00202f
C10540 _063_ _190_/a_27_47# 0.00437f
C10541 _248_/a_109_297# net21 2.6e-21
C10542 VPWR _220_/a_113_297# 0.0655f
C10543 net22 _315_/a_1108_47# 8.95e-21
C10544 net4 _335_/a_27_47# 2.87e-19
C10545 _253_/a_81_21# _074_ 0.0581f
C10546 VPWR _169_/a_373_53# -3.18e-19
C10547 _234_/a_109_297# mask\[0\] 4.5e-19
C10548 trim_mask\[1\] _336_/a_1108_47# 2.78e-19
C10549 VPWR net54 0.227f
C10550 _192_/a_174_21# _065_ 0.0156f
C10551 _014_ _315_/a_27_47# 1.2e-20
C10552 clknet_2_0__leaf_clk _315_/a_193_47# 0.00951f
C10553 _125_ _133_ 4.17e-21
C10554 cal_itt\[2\] _065_ 0.00575f
C10555 _087_ _099_ 0.106f
C10556 _249_/a_109_47# _101_ 0.00454f
C10557 _050_ clknet_2_2__leaf_clk 0.00221f
C10558 _040_ _246_/a_373_47# 0.00356f
C10559 _050_ _260_/a_584_47# 1.85e-20
C10560 trim_mask\[0\] rebuffer2/a_75_212# 2.87e-20
C10561 mask\[3\] net52 0.188f
C10562 _082_ _101_ 8.79e-21
C10563 fanout43/a_27_47# net14 0.00189f
C10564 trim_mask\[0\] _332_/a_1283_21# 0.107f
C10565 _273_/a_59_75# _334_/a_543_47# 2.63e-20
C10566 _326_/a_805_47# mask\[7\] 9e-20
C10567 cal_itt\[2\] _105_ 9.08e-20
C10568 mask\[5\] net20 0.0649f
C10569 _286_/a_505_21# _122_ 7.4e-19
C10570 trim_mask\[0\] _111_ 0.226f
C10571 VPWR _178_/a_68_297# 0.0208f
C10572 cal valid 0.0947f
C10573 mask\[5\] net53 0.114f
C10574 _136_ _300_/a_129_47# 0.00104f
C10575 net27 net14 0.00986f
C10576 trimb[3] net16 3.69e-19
C10577 _041_ _286_/a_218_47# 0.0019f
C10578 _110_ net55 8.54e-21
C10579 net47 cal_count\[0\] 0.268f
C10580 clk _068_ 2.05e-20
C10581 _324_/a_1283_21# _020_ 8.91e-19
C10582 VPWR _246_/a_373_47# -1.79e-19
C10583 _006_ _310_/a_27_47# 1.34e-21
C10584 VPWR result[4] 0.0909f
C10585 net15 clknet_0_clk 0.0846f
C10586 _048_ _279_/a_396_47# 0.00276f
C10587 _235_/a_79_21# clknet_0_clk 8.61e-20
C10588 result[2] _078_ 4.7e-20
C10589 trim_mask\[0\] calibrate 4.16e-20
C10590 _328_/a_27_47# _336_/a_27_47# 1.59e-21
C10591 _236_/a_109_297# _050_ 0.00217f
C10592 _072_ _201_/a_113_47# 2.29e-19
C10593 VPWR _327_/a_1217_47# 1.49e-19
C10594 _263_/a_297_47# _099_ 0.0373f
C10595 net24 clknet_2_0__leaf_clk 1.23e-19
C10596 _004_ _210_/a_199_47# 1.84e-21
C10597 _038_ _108_ 1.47e-19
C10598 _317_/a_1462_47# state\[1\] 6.42e-19
C10599 clknet_2_0__leaf_clk _014_ 0.0967f
C10600 _062_ clkbuf_2_3__f_clk/a_110_47# 0.159f
C10601 output31/a_27_47# net34 0.0251f
C10602 _133_ net40 0.00147f
C10603 result[0] sample 0.0473f
C10604 _074_ _313_/a_639_47# 1.35e-20
C10605 input2/a_27_47# _297_/a_47_47# 1.11e-19
C10606 _256_/a_27_297# trim_mask\[1\] 0.015f
C10607 trim_mask\[4\] _279_/a_396_47# 6.28e-19
C10608 _025_ trim_val\[4\] 1.11e-20
C10609 net8 net9 0.00149f
C10610 net4 _068_ 0.00707f
C10611 _051_ _093_ 1.44e-20
C10612 _327_/a_543_47# _025_ 9.83e-21
C10613 _064_ _119_ 0.0152f
C10614 _319_/a_1108_47# _049_ 0.00215f
C10615 _110_ _336_/a_1462_47# 2.04e-19
C10616 _324_/a_1108_47# net27 0.00103f
C10617 VPWR fanout43/a_27_47# 0.0977f
C10618 _015_ _090_ 6.44e-20
C10619 output15/a_27_47# _223_/a_109_297# 5.98e-20
C10620 _305_/a_761_289# clk 3.45e-19
C10621 net12 _305_/a_193_47# 3.97e-19
C10622 VPWR output35/a_27_47# 0.136f
C10623 _083_ mask\[3\] 6.93e-20
C10624 _040_ rebuffer5/a_161_47# 1.1e-20
C10625 trim_val\[1\] net32 0.00288f
C10626 VPWR net27 0.906f
C10627 _313_/a_27_47# net29 0.00312f
C10628 _195_/a_76_199# clkbuf_2_3__f_clk/a_110_47# 1.49e-19
C10629 cal_itt\[1\] _304_/a_27_47# 1.02e-19
C10630 cal_itt\[0\] _304_/a_193_47# 2.67e-20
C10631 VPWR _222_/a_113_297# 0.0728f
C10632 _331_/a_193_47# _330_/a_193_47# 0.00469f
C10633 _321_/a_543_47# _018_ 2.12e-19
C10634 _269_/a_299_297# _172_/a_68_297# 0.00615f
C10635 net8 trim[2] 2.25e-19
C10636 trim_mask\[0\] _135_ 2.05e-20
C10637 net13 _077_ 2.18e-20
C10638 trim_mask\[2\] _335_/a_1283_21# 2.02e-20
C10639 _008_ mask\[5\] 1.37e-19
C10640 _053_ _119_ 0.00168f
C10641 _341_/a_543_47# net46 1.58e-19
C10642 _246_/a_373_47# net52 7.28e-19
C10643 VPWR _186_/a_109_297# -0.0017f
C10644 mask\[0\] _319_/a_761_289# 0.0221f
C10645 _078_ _319_/a_193_47# 1.47e-21
C10646 _043_ net26 8.16e-19
C10647 net50 _327_/a_27_47# 0.00315f
C10648 _321_/a_27_47# mask\[6\] 6.01e-19
C10649 net14 sample 8.01e-20
C10650 VPWR rebuffer5/a_161_47# 0.0694f
C10651 _058_ net19 2.29e-20
C10652 _321_/a_448_47# _042_ 2.86e-19
C10653 _307_/a_193_47# _137_/a_68_297# 1.18e-19
C10654 VPWR _125_ 0.161f
C10655 _305_/a_193_47# net44 0.0117f
C10656 net31 output37/a_27_47# 0.0146f
C10657 net23 fanout43/a_27_47# 0.0294f
C10658 net44 _311_/a_1108_47# -0.00124f
C10659 _322_/a_1283_21# rebuffer5/a_161_47# 1.06e-20
C10660 mask\[4\] net19 0.0812f
C10661 _048_ _034_ 2.06e-21
C10662 trim_mask\[2\] _108_ 0.167f
C10663 _321_/a_805_47# clknet_2_1__leaf_clk 4.26e-19
C10664 _327_/a_193_47# _107_ 5.4e-21
C10665 _093_ _316_/a_1283_21# 9.52e-20
C10666 _115_ _334_/a_448_47# 5.13e-19
C10667 trim_mask\[3\] _058_ 4.79e-21
C10668 _259_/a_109_297# trim_mask\[3\] 0.00883f
C10669 _064_ _275_/a_81_21# 1.27e-19
C10670 _259_/a_27_297# net50 0.0102f
C10671 _323_/a_27_47# _311_/a_1283_21# 9.27e-19
C10672 _340_/a_381_47# _123_ 0.0144f
C10673 _281_/a_253_47# _090_ 9.8e-19
C10674 clknet_2_1__leaf_clk _313_/a_448_47# 0.0149f
C10675 _053_ _087_ 3.09e-20
C10676 mask\[7\] _224_/a_113_297# 2.22e-19
C10677 _286_/a_218_47# net18 3.63e-19
C10678 VPWR _306_/a_27_47# 0.0881f
C10679 _327_/a_1108_47# _265_/a_81_21# 4.92e-20
C10680 _312_/a_27_47# _084_ 0.0128f
C10681 _326_/a_27_47# net14 0.00737f
C10682 fanout43/a_27_47# net52 6.06e-19
C10683 _097_ _096_ 0.00344f
C10684 _058_ _107_ 4.44e-19
C10685 _015_ _048_ 2.39e-20
C10686 _305_/a_761_289# _073_ 2.27e-20
C10687 _341_/a_1283_21# _300_/a_47_47# 2.14e-19
C10688 _322_/a_639_47# mask\[2\] 4.73e-19
C10689 net27 net52 3.96e-19
C10690 _058_ _333_/a_1108_47# 3.95e-19
C10691 _217_/a_109_297# _007_ 0.00408f
C10692 _042_ _143_/a_68_297# 7.6e-19
C10693 net15 _245_/a_27_297# 6.52e-19
C10694 output33/a_27_47# _162_/a_27_47# 2.14e-20
C10695 _187_/a_212_413# _134_ 6.6e-19
C10696 _061_ _301_/a_47_47# 5.51e-19
C10697 cal_itt\[1\] _069_ 0.0957f
C10698 cal_count\[3\] _062_ 0.0484f
C10699 VPWR sample 0.201f
C10700 VPWR net40 1.82f
C10701 trim_mask\[0\] _112_ 1.56e-19
C10702 _253_/a_81_21# net26 0.0495f
C10703 net9 _340_/a_27_47# 0.019f
C10704 _134_ _332_/a_193_47# 4.73e-20
C10705 state\[2\] _028_ 0.00598f
C10706 _155_/a_68_297# _045_ 6.76e-19
C10707 trim_mask\[2\] _031_ 0.12f
C10708 _007_ _216_/a_113_297# 2.9e-19
C10709 net28 net15 0.0994f
C10710 net31 _134_ 4.59e-22
C10711 _119_ _330_/a_448_47# 4.88e-19
C10712 _313_/a_1108_47# _009_ 4.04e-20
C10713 net52 rebuffer5/a_161_47# 0.00512f
C10714 _072_ _202_/a_297_47# 3.5e-19
C10715 output22/a_27_47# _074_ 0.00596f
C10716 _060_ _107_ 0.00674f
C10717 _102_ clknet_2_1__leaf_clk 1.34e-19
C10718 net43 _306_/a_543_47# 1.25e-19
C10719 _002_ clkbuf_0_clk/a_110_47# 0.00165f
C10720 _329_/a_1270_413# net46 1.61e-19
C10721 net46 clknet_2_3__leaf_clk 0.374f
C10722 VPWR _330_/a_639_47# 4.33e-19
C10723 _115_ _108_ 0.00253f
C10724 _339_/a_27_47# _124_ 2.96e-21
C10725 net50 _178_/a_68_297# 8.75e-19
C10726 _275_/a_81_21# _057_ 1.13e-19
C10727 output8/a_27_47# net8 0.0121f
C10728 _294_/a_68_297# cal_count\[1\] 4.41e-21
C10729 output37/a_27_47# net2 3.29e-20
C10730 _020_ net19 0.0017f
C10731 net12 _250_/a_109_47# 3.88e-20
C10732 _214_/a_113_297# clkbuf_2_1__f_clk/a_110_47# 1.49e-19
C10733 _216_/a_113_297# mask\[3\] 0.00226f
C10734 _216_/a_199_47# net25 5.39e-20
C10735 _089_ _226_/a_27_47# 2.73e-19
C10736 _337_/a_651_413# _049_ 0.00244f
C10737 VPWR _267_/a_145_75# -3.02e-19
C10738 clk _317_/a_27_47# 0.00834f
C10739 _104_ clknet_2_2__leaf_clk 0.0678f
C10740 net31 _130_ 0.00142f
C10741 cal_itt\[1\] _304_/a_1217_47# 1.09e-19
C10742 VPWR _235_/a_382_297# -7e-19
C10743 _104_ _260_/a_584_47# 0.00189f
C10744 ctlp[0] net28 0.0759f
C10745 VPWR _326_/a_27_47# 0.0514f
C10746 _101_ _076_ 0.036f
C10747 _329_/a_27_47# _031_ 8.51e-20
C10748 VPWR _334_/a_27_47# 0.0955f
C10749 _051_ _171_/a_27_47# 0.0094f
C10750 VPWR _228_/a_382_297# -9.84e-19
C10751 _048_ _281_/a_253_47# 0.00302f
C10752 _306_/a_27_47# net52 2.88e-20
C10753 _306_/a_761_289# _101_ 1.05e-20
C10754 _320_/a_193_47# clkbuf_2_1__f_clk/a_110_47# 0.00198f
C10755 net5 _131_ 0.00988f
C10756 _276_/a_59_75# clkbuf_2_2__f_clk/a_110_47# 2.09e-21
C10757 _006_ clknet_2_1__leaf_clk 0.00374f
C10758 _307_/a_1283_21# _039_ 0.0346f
C10759 _325_/a_1108_47# mask\[4\] 7.84e-19
C10760 net27 _083_ 2.92e-21
C10761 net24 _321_/a_27_47# 1.24e-20
C10762 cal_itt\[2\] clkbuf_0_clk/a_110_47# 0.0416f
C10763 _320_/a_1283_21# net51 2e-20
C10764 net4 _317_/a_27_47# 0.0101f
C10765 _321_/a_193_47# clknet_2_0__leaf_clk 9.79e-21
C10766 net45 net55 1.01e-19
C10767 net14 _310_/a_761_289# 0.0115f
C10768 net27 _312_/a_1270_413# 8.03e-20
C10769 net2 _298_/a_215_47# 0.00118f
C10770 _233_/a_109_47# net14 9.7e-20
C10771 output22/a_27_47# output23/a_27_47# 5.69e-19
C10772 _074_ _013_ 1.14e-20
C10773 _338_/a_1032_413# _123_ 6.77e-19
C10774 _300_/a_377_297# clknet_2_3__leaf_clk 2.43e-21
C10775 _181_/a_68_297# _058_ 0.00155f
C10776 _115_ _031_ 0.00172f
C10777 _337_/a_193_47# clknet_2_0__leaf_clk 0.109f
C10778 result[6] _314_/a_543_47# 8.65e-19
C10779 net28 _314_/a_1108_47# 1.46e-19
C10780 net47 net16 7.59e-20
C10781 _059_ _090_ 0.0303f
C10782 _309_/a_27_47# _310_/a_1283_21# 1.17e-19
C10783 _283_/a_75_212# _034_ 0.00249f
C10784 _063_ net40 4.59e-19
C10785 clknet_2_1__leaf_clk _010_ 0.0338f
C10786 _326_/a_543_47# net43 0.00396f
C10787 VPWR _306_/a_1217_47# 7.1e-20
C10788 _103_ net55 0.0766f
C10789 _134_ net2 0.501f
C10790 _257_/a_109_297# _335_/a_193_47# 5.17e-22
C10791 _323_/a_761_289# clknet_2_1__leaf_clk 2.53e-19
C10792 en_co_clk net19 0.00479f
C10793 cal_itt\[0\] trim_mask\[0\] 7.46e-19
C10794 _341_/a_1108_47# _135_ 2.01e-19
C10795 _065_ net55 7.5e-20
C10796 _095_ _092_ 0.337f
C10797 VPWR _314_/a_448_47# 0.00137f
C10798 _231_/a_161_47# en_co_clk 0.00148f
C10799 clk _318_/a_543_47# 0.0298f
C10800 output26/a_27_47# _007_ 0.00126f
C10801 _233_/a_27_297# valid 0.00378f
C10802 net12 _049_ 0.214f
C10803 net12 _318_/a_761_289# 9.81e-19
C10804 output31/a_27_47# VPWR 4.12e-19
C10805 net2 _130_ 0.124f
C10806 _326_/a_27_47# net52 3.61e-19
C10807 _105_ net55 0.0334f
C10808 trim_mask\[2\] net49 1.51e-19
C10809 trim_mask\[2\] _272_/a_81_21# 0.054f
C10810 net9 _340_/a_586_47# 7.81e-19
C10811 _253_/a_299_297# _078_ 0.00324f
C10812 _304_/a_27_47# _304_/a_193_47# -0.079f
C10813 _169_/a_215_311# _099_ 1.08e-21
C10814 _325_/a_27_47# mask\[2\] 1.68e-19
C10815 _307_/a_805_47# _074_ 6.43e-19
C10816 _307_/a_639_47# calibrate 2.23e-20
C10817 _119_ _027_ 6.44e-20
C10818 VPWR _310_/a_761_289# 0.0152f
C10819 _326_/a_805_47# net28 2.68e-20
C10820 VPWR _233_/a_109_47# -9.1e-19
C10821 _340_/a_193_47# cal_count\[2\] 8.14e-20
C10822 _001_ en_co_clk 6.44e-20
C10823 output7/a_27_47# VPWR 0.0642f
C10824 _067_ _065_ 0.0259f
C10825 net4 _318_/a_543_47# 1.8e-20
C10826 _065_ _070_ 0.657f
C10827 _327_/a_27_47# _327_/a_1108_47# -2.98e-20
C10828 _327_/a_193_47# _327_/a_1283_21# -9.43e-20
C10829 output15/a_27_47# _010_ 0.0629f
C10830 _243_/a_109_297# net55 0.0372f
C10831 _090_ _075_ 6.42e-21
C10832 _304_/a_805_47# _065_ 3.02e-20
C10833 net44 _049_ 0.0558f
C10834 clk _317_/a_1217_47# 5.25e-20
C10835 _317_/a_651_413# _316_/a_543_47# 3.6e-21
C10836 net2 _339_/a_1602_47# 3.98e-20
C10837 _185_/a_68_297# _060_ 0.0267f
C10838 VPWR _326_/a_1217_47# 1.17e-19
C10839 VPWR _271_/a_75_212# 0.00951f
C10840 VPWR _334_/a_1217_47# 1.01e-19
C10841 _059_ _048_ 0.0254f
C10842 _123_ _298_/a_215_47# 8.14e-19
C10843 _267_/a_59_75# clknet_2_2__leaf_clk 0.0181f
C10844 _254_/a_109_297# _098_ 0.002f
C10845 _104_ _279_/a_204_297# 5.82e-19
C10846 _058_ _118_ 0.00858f
C10847 _327_/a_1283_21# _058_ 0.0143f
C10848 net2 rebuffer6/a_27_47# 4.99e-20
C10849 clk cal_itt\[3\] 0.0472f
C10850 _238_/a_75_212# _316_/a_448_47# 5.77e-19
C10851 _097_ _316_/a_761_289# 1.11e-19
C10852 trim_mask\[1\] net18 0.204f
C10853 _311_/a_761_289# net53 0.00351f
C10854 net43 _310_/a_1108_47# 0.0202f
C10855 _330_/a_805_47# net19 3.89e-19
C10856 net13 clkbuf_2_1__f_clk/a_110_47# 2.91e-19
C10857 net50 net40 0.0315f
C10858 net4 _317_/a_1217_47# 5.18e-19
C10859 _134_ _123_ 2.37e-20
C10860 _274_/a_75_212# trim_val\[2\] 1.82e-19
C10861 _049_ _003_ 1.6e-19
C10862 _115_ _272_/a_81_21# 0.00215f
C10863 _273_/a_59_75# net48 4.38e-19
C10864 net2 cal_count\[3\] 0.0537f
C10865 _324_/a_1108_47# _311_/a_1283_21# 1.27e-20
C10866 _301_/a_47_47# net16 0.0132f
C10867 _089_ _052_ 0.00686f
C10868 VPWR _300_/a_285_47# 0.00391f
C10869 _200_/a_80_21# clknet_0_clk 4.96e-19
C10870 _266_/a_68_297# net46 2.34e-20
C10871 _337_/a_805_47# net45 5.61e-21
C10872 VPWR _335_/a_639_47# 7.26e-19
C10873 _323_/a_1108_47# net26 7.59e-19
C10874 VPWR _305_/a_27_47# 0.066f
C10875 _309_/a_651_413# _074_ 1.23e-20
C10876 VPWR _311_/a_1283_21# 0.0168f
C10877 _040_ net51 0.00283f
C10878 output10/a_27_47# _335_/a_193_47# 2.95e-19
C10879 _015_ net54 0.00246f
C10880 net4 cal_itt\[3\] 7.46e-21
C10881 _274_/a_75_212# net16 6.84e-19
C10882 net16 _299_/a_215_297# 0.0116f
C10883 ctln[4] trim_val\[3\] 0.00181f
C10884 VPWR _332_/a_1270_413# -1.76e-19
C10885 _088_ _242_/a_79_21# 1.81e-20
C10886 _194_/a_113_297# _067_ 0.0118f
C10887 _304_/a_27_47# _302_/a_27_297# 2.43e-20
C10888 _041_ _078_ 0.409f
C10889 _048_ _075_ 0.0203f
C10890 _287_/a_75_212# _035_ 0.0138f
C10891 _110_ clknet_2_3__leaf_clk 1.07e-20
C10892 output26/a_27_47# result[4] 0.00962f
C10893 _290_/a_207_413# net38 4.06e-21
C10894 VPWR net51 0.338f
C10895 _188_/a_27_47# trim_mask\[0\] 3.43e-20
C10896 _136_ cal_count\[2\] 9.64e-19
C10897 net9 _338_/a_956_413# 1.21e-19
C10898 net9 _341_/a_193_47# 0.00198f
C10899 clkbuf_2_2__f_clk/a_110_47# net30 5.18e-19
C10900 _336_/a_761_289# _106_ 6.44e-20
C10901 clk net6 0.00704f
C10902 _107_ _228_/a_297_47# 7.76e-19
C10903 trim[3] _057_ 3.31e-19
C10904 _334_/a_1108_47# _175_/a_68_297# 2.85e-20
C10905 net43 _305_/a_543_47# 0.0334f
C10906 _267_/a_59_75# trim_val\[0\] 3.87e-19
C10907 trim[2] net34 0.0157f
C10908 _073_ cal_itt\[3\] 0.0364f
C10909 _321_/a_27_47# _321_/a_193_47# -0.32f
C10910 trim_val\[3\] _335_/a_27_47# 0.0124f
C10911 _284_/a_150_297# _065_ 0.00156f
C10912 net28 _224_/a_113_297# 0.0628f
C10913 _008_ _311_/a_761_289# 6.55e-19
C10914 _286_/a_76_199# _001_ 1.8e-19
C10915 net43 clkbuf_2_1__f_clk/a_110_47# 0.00886f
C10916 clknet_2_0__leaf_clk _316_/a_1108_47# 2.11e-21
C10917 _014_ _316_/a_1283_21# 3.34e-20
C10918 net45 _316_/a_543_47# 0.00238f
C10919 calibrate _331_/a_1270_413# 2.39e-20
C10920 _338_/a_27_47# _065_ 1.44e-20
C10921 _169_/a_215_311# _053_ 0.00359f
C10922 _169_/a_109_53# state\[0\] 0.034f
C10923 _337_/a_761_289# net55 0.00343f
C10924 _337_/a_543_47# _096_ 4.24e-19
C10925 VPWR _269_/a_384_47# -2.23e-19
C10926 net34 _132_ 0.0169f
C10927 rstn ctln[0] 2.27e-19
C10928 net4 net6 0.0663f
C10929 _074_ _046_ 5.07e-20
C10930 _305_/a_27_47# net52 5.39e-21
C10931 _051_ _243_/a_27_297# 2.4e-20
C10932 _305_/a_27_47# _063_ 4.88e-21
C10933 _337_/a_27_47# _337_/a_193_47# -0.0515f
C10934 _307_/a_1283_21# _049_ 1.66e-19
C10935 _101_ _311_/a_448_47# 2.57e-21
C10936 cal_count\[1\] cal_count\[0\] 0.112f
C10937 _307_/a_761_289# net30 4.59e-21
C10938 calibrate _089_ 0.0219f
C10939 output26/a_27_47# net27 7.85e-21
C10940 _123_ cal_count\[3\] 1.48e-19
C10941 VPWR _224_/a_199_47# -1.42e-19
C10942 _309_/a_1283_21# clknet_2_1__leaf_clk 5.21e-21
C10943 _329_/a_1108_47# net16 6.01e-21
C10944 _128_ net2 0.0683f
C10945 trim_mask\[0\] net33 0.0121f
C10946 _074_ _312_/a_761_289# 1.75e-20
C10947 _238_/a_75_212# _013_ 0.0027f
C10948 trim_mask\[0\] _336_/a_761_289# 1.49e-20
C10949 net47 _149_/a_68_297# 0.00372f
C10950 _262_/a_27_47# _098_ 1.07e-20
C10951 _032_ _119_ 2.87e-21
C10952 _299_/a_298_297# _132_ 8.29e-19
C10953 _226_/a_27_47# _092_ 0.0669f
C10954 net52 net51 0.228f
C10955 _326_/a_27_47# _216_/a_113_297# 5.86e-22
C10956 _326_/a_1108_47# _325_/a_193_47# 1.29e-20
C10957 _071_ clknet_0_clk 0.0306f
C10958 _121_ net45 2.82e-20
C10959 fanout45/a_27_47# _096_ 5.43e-19
C10960 clknet_2_1__leaf_clk net20 0.0971f
C10961 _333_/a_27_47# _332_/a_543_47# 2.44e-21
C10962 _333_/a_27_47# _108_ 0.00562f
C10963 _324_/a_543_47# _042_ 8.95e-20
C10964 clknet_2_1__leaf_clk net53 0.87f
C10965 VPWR _305_/a_1217_47# 9.49e-21
C10966 _307_/a_27_47# _078_ 0.00861f
C10967 _307_/a_193_47# mask\[0\] 0.00201f
C10968 _307_/a_761_289# net22 0.0371f
C10969 trim_mask\[0\] clone1/a_27_47# 9.29e-20
C10970 VPWR _250_/a_109_297# 0.00823f
C10971 trim_val\[0\] net37 0.0153f
C10972 _158_/a_68_297# _085_ 1.59e-19
C10973 _265_/a_299_297# _332_/a_193_47# 4.56e-20
C10974 _265_/a_81_21# _332_/a_761_289# 3.19e-19
C10975 state\[2\] state\[0\] 0.00797f
C10976 _051_ _336_/a_543_47# 4.44e-21
C10977 net9 _133_ 1.33e-19
C10978 _329_/a_448_47# net9 0.00125f
C10979 _041_ fanout47/a_27_47# 0.0425f
C10980 clknet_0_clk _262_/a_27_47# 0.00311f
C10981 _335_/a_543_47# trim_mask\[4\] 4.33e-20
C10982 _322_/a_1283_21# _250_/a_109_297# 1.33e-21
C10983 _136_ _194_/a_199_47# 1.49e-19
C10984 _302_/a_109_297# _067_ 0.00139f
C10985 _121_ _065_ 0.26f
C10986 _304_/a_543_47# _136_ 0.00126f
C10987 _000_ net2 9.24e-22
C10988 _117_ VPWR 0.0327f
C10989 ctln[2] _179_/a_27_47# 0.00504f
C10990 output8/a_27_47# net34 8.93e-19
C10991 _064_ _053_ 0.0826f
C10992 _304_/a_543_47# _284_/a_68_297# 4.89e-19
C10993 net9 _341_/a_1462_47# 4.41e-20
C10994 _083_ _311_/a_1283_21# 7.61e-22
C10995 _122_ _131_ 0.0065f
C10996 fanout46/a_27_47# clknet_2_2__leaf_clk 0.105f
C10997 _305_/a_193_47# net19 1.43e-20
C10998 _304_/a_1108_47# net47 0.0177f
C10999 cal_itt\[1\] _261_/a_113_47# 2.8e-20
C11000 _094_ _050_ 0.00885f
C11001 net28 _009_ 8.18e-21
C11002 _062_ _190_/a_215_47# 7.64e-19
C11003 _311_/a_1108_47# net19 5.66e-19
C11004 _200_/a_209_297# VPWR -0.0168f
C11005 _030_ _333_/a_193_47# 0.111f
C11006 _113_ _333_/a_761_289# 7.33e-21
C11007 net43 _251_/a_109_47# 3.35e-21
C11008 net13 _318_/a_1283_21# 0.00214f
C11009 ctln[7] _318_/a_761_289# 8.2e-20
C11010 net13 net30 0.0102f
C11011 _308_/a_1108_47# _078_ 0.0125f
C11012 _050_ _088_ 0.121f
C11013 _037_ _131_ 1.12e-19
C11014 _340_/a_193_47# _340_/a_1602_47# -4.7e-21
C11015 _340_/a_27_47# _340_/a_381_47# -0.00396f
C11016 _030_ _265_/a_81_21# 2.45e-19
C11017 net50 _335_/a_639_47# 3.14e-19
C11018 _275_/a_81_21# _032_ 6.04e-19
C11019 net44 _319_/a_543_47# 2.16e-20
C11020 _308_/a_27_47# result[2] 9.42e-19
C11021 _308_/a_193_47# net45 9.57e-19
C11022 _308_/a_543_47# clknet_2_0__leaf_clk 7.75e-19
C11023 _149_/a_68_297# net44 1.91e-19
C11024 output28/a_27_47# result[7] 0.0564f
C11025 _299_/a_27_413# _131_ 0.0156f
C11026 _299_/a_382_47# cal_count\[2\] 8.88e-19
C11027 _133_ _132_ 0.00409f
C11028 wire42/a_75_212# _098_ 0.0126f
C11029 _281_/a_253_297# _120_ 6.75e-19
C11030 _281_/a_337_297# en_co_clk 0.00424f
C11031 clkbuf_0_clk/a_110_47# _067_ 0.00733f
C11032 _059_ net54 0.216f
C11033 _128_ _123_ 0.2f
C11034 cal_count\[0\] _001_ 4.97e-19
C11035 clkbuf_0_clk/a_110_47# _070_ 0.00201f
C11036 _341_/a_543_47# _065_ 0.00413f
C11037 _251_/a_109_297# _101_ 0.0497f
C11038 _119_ _171_/a_27_47# 2.72e-19
C11039 _008_ clknet_2_1__leaf_clk 0.116f
C11040 _313_/a_193_47# _313_/a_543_47# -0.0102f
C11041 cal_itt\[0\] _303_/a_543_47# 1.64e-19
C11042 _071_ _303_/a_27_47# 1.33e-19
C11043 _042_ _101_ 0.0277f
C11044 _110_ _266_/a_68_297# 6.83e-19
C11045 trim[1] trim_val\[0\] 0.00234f
C11046 VPWR _318_/a_193_47# -0.276f
C11047 clknet_0_clk wire42/a_75_212# 8.82e-22
C11048 _325_/a_27_47# _074_ 1.71e-20
C11049 _232_/a_114_297# _090_ 0.00662f
C11050 _326_/a_27_47# output26/a_27_47# 3.9e-19
C11051 _041_ _287_/a_75_212# 0.0515f
C11052 _294_/a_150_297# _299_/a_27_413# 1.95e-19
C11053 _208_/a_76_199# rebuffer5/a_161_47# 0.00349f
C11054 clknet_2_1__leaf_clk _016_ 0.0775f
C11055 _331_/a_193_47# _054_ 1.63e-22
C11056 _331_/a_543_47# _049_ 1.15e-19
C11057 trim_mask\[2\] _336_/a_193_47# 6.73e-20
C11058 net24 _140_/a_68_297# 1.86e-19
C11059 _024_ _264_/a_27_297# 2.56e-20
C11060 _324_/a_1108_47# _021_ 7.95e-20
C11061 input2/a_27_47# net40 2.19e-20
C11062 _326_/a_1108_47# mask\[3\] 1.09e-21
C11063 _333_/a_1217_47# _108_ 2.9e-19
C11064 _307_/a_1217_47# _078_ 5.09e-19
C11065 _307_/a_1462_47# mask\[0\] 3.18e-19
C11066 _104_ _330_/a_1283_21# 0.00112f
C11067 _328_/a_193_47# _026_ 1.18e-19
C11068 VPWR _021_ 0.0456f
C11069 _328_/a_193_47# VPWR -0.298f
C11070 _330_/a_27_47# _330_/a_193_47# -0.292f
C11071 trim_val\[0\] _332_/a_651_413# 4.58e-20
C11072 _200_/a_209_297# _063_ 0.0069f
C11073 _189_/a_408_47# _048_ 1.44e-19
C11074 _026_ net9 0.0184f
C11075 _308_/a_27_47# _319_/a_193_47# 1.77e-21
C11076 _308_/a_193_47# _319_/a_27_47# 8.25e-20
C11077 _302_/a_109_47# _136_ 1.26e-19
C11078 _051_ _106_ 5.03e-19
C11079 trim[3] _334_/a_1270_413# 1.63e-20
C11080 _168_/a_207_413# _331_/a_27_47# 1.17e-19
C11081 VPWR net9 0.941f
C11082 _111_ _109_ 8.27e-19
C11083 _306_/a_27_47# _208_/a_76_199# 1.43e-20
C11084 _307_/a_761_289# _079_ 3.2e-19
C11085 _307_/a_27_47# _004_ 0.037f
C11086 VPWR _317_/a_639_47# 1.75e-20
C11087 VPWR output16/a_27_47# 0.0706f
C11088 clknet_2_3__leaf_clk rebuffer3/a_75_212# 1.9e-19
C11089 _315_/a_1283_21# net14 1.52e-19
C11090 _304_/a_27_47# _298_/a_78_199# 6.77e-20
C11091 _060_ _062_ 0.0644f
C11092 _038_ _067_ 3.04e-20
C11093 net43 result[7] 9.52e-20
C11094 net43 net30 0.156f
C11095 net36 net37 0.00645f
C11096 _319_/a_193_47# clknet_0_clk 0.00163f
C11097 _074_ _212_/a_199_47# 4.22e-19
C11098 output36/a_27_47# net38 0.0398f
C11099 _019_ clknet_2_1__leaf_clk 0.00835f
C11100 _320_/a_193_47# _319_/a_1108_47# 9.6e-21
C11101 _218_/a_113_297# mask\[6\] 2.62e-20
C11102 _052_ _092_ 3.03e-19
C11103 _304_/a_448_47# _122_ 0.0014f
C11104 ctlp[7] _313_/a_1462_47# 1.98e-20
C11105 ctlp[6] output20/a_27_47# 0.0443f
C11106 _086_ net14 0.0147f
C11107 net12 _337_/a_1108_47# 2.05e-19
C11108 _336_/a_27_47# net18 7.34e-22
C11109 trim_mask\[1\] _175_/a_68_297# 1.33e-19
C11110 mask\[6\] _312_/a_27_47# 5.53e-20
C11111 _198_/a_27_47# _072_ 8.68e-20
C11112 trim_mask\[1\] _333_/a_193_47# 0.00414f
C11113 net49 _333_/a_27_47# 0.0136f
C11114 trim_val\[1\] _333_/a_761_289# 9.6e-19
C11115 _065_ clknet_2_3__leaf_clk 0.305f
C11116 VPWR _192_/a_639_47# -4.73e-19
C11117 _116_ clknet_2_2__leaf_clk 2.26e-20
C11118 VPWR trim[2] 0.277f
C11119 output32/a_27_47# _058_ 0.0029f
C11120 _037_ _304_/a_448_47# 2.13e-19
C11121 _315_/a_761_289# valid 9.39e-19
C11122 net43 net22 2.63e-19
C11123 _005_ mask\[0\] 3.99e-20
C11124 _259_/a_27_297# _335_/a_543_47# 0.00351f
C11125 net42 _260_/a_93_21# 5.04e-19
C11126 _005_ output24/a_27_47# 7.02e-19
C11127 _186_/a_109_297# _059_ 3.87e-19
C11128 _308_/a_1462_47# net45 5.4e-19
C11129 VPWR _262_/a_109_297# 0.00534f
C11130 VPWR _132_ 0.455f
C11131 _253_/a_299_297# mask\[7\] 0.00859f
C11132 _309_/a_1270_413# _078_ 9.62e-20
C11133 trim_mask\[0\] _051_ 0.0104f
C11134 _116_ net11 5.63e-20
C11135 cal_count\[1\] net16 0.0384f
C11136 _187_/a_212_413# _058_ 7.15e-20
C11137 _323_/a_761_289# _043_ 2.03e-21
C11138 mask\[1\] _039_ 1.8e-20
C11139 output30/a_27_47# sample 0.0106f
C11140 VPWR _315_/a_1283_21# 0.059f
C11141 clknet_0_clk _202_/a_79_21# 2.29e-19
C11142 _022_ _101_ 0.0143f
C11143 _303_/a_193_47# _065_ 1.73e-20
C11144 _309_/a_1108_47# net24 0.0577f
C11145 _068_ _190_/a_655_47# 0.0412f
C11146 _337_/a_1108_47# net44 0.0261f
C11147 _048_ _170_/a_81_21# 2.47e-19
C11148 _309_/a_1283_21# net45 1.36e-20
C11149 VPWR _234_/a_109_297# 4.65e-20
C11150 _058_ _332_/a_193_47# 0.00777f
C11151 net43 _072_ 0.0964f
C11152 _278_/a_109_297# net40 6.04e-19
C11153 net25 _310_/a_1270_413# 2.35e-19
C11154 net15 mask\[2\] 0.291f
C11155 _051_ _337_/a_1462_47# 3.32e-20
C11156 VPWR _318_/a_1462_47# 0.00178f
C11157 trim_mask\[1\] trim_mask\[4\] 0.0742f
C11158 _074_ net25 0.123f
C11159 _200_/a_209_47# net19 6.7e-19
C11160 net31 _058_ 5.96e-20
C11161 net45 _245_/a_109_297# 0.0535f
C11162 net27 _314_/a_27_47# 0.00152f
C11163 _117_ net50 9.65e-19
C11164 _327_/a_651_413# net46 0.00109f
C11165 _287_/a_75_212# net18 2.08e-19
C11166 clkbuf_2_0__f_clk/a_110_47# _241_/a_297_47# 1.08e-19
C11167 trim_mask\[4\] _170_/a_81_21# 1.48e-20
C11168 _260_/a_256_47# _049_ 0.00179f
C11169 _260_/a_93_21# _054_ 0.00149f
C11170 VPWR _086_ 0.0472f
C11171 _048_ _227_/a_296_53# 1.17e-19
C11172 _341_/a_193_47# _091_ 2.12e-20
C11173 net45 valid 3.94e-19
C11174 _036_ net9 0.18f
C11175 net34 net32 0.459f
C11176 state\[2\] _052_ 0.346f
C11177 _064_ _027_ 0.00133f
C11178 clknet_0_clk _206_/a_27_93# 0.0422f
C11179 output12/a_27_47# ctln[6] 0.0141f
C11180 _328_/a_1462_47# VPWR 1.46e-19
C11181 _077_ _076_ 0.00498f
C11182 calibrate _092_ 0.0617f
C11183 _093_ _099_ 0.0555f
C11184 _305_/a_1108_47# _190_/a_27_47# 4.06e-20
C11185 _194_/a_113_297# clknet_2_3__leaf_clk 0.0227f
C11186 _200_/a_209_47# _107_ 1.42e-19
C11187 net19 _049_ 1.21e-20
C11188 en_co_clk _062_ 0.114f
C11189 net3 _317_/a_193_47# 8.87e-20
C11190 _306_/a_543_47# _076_ 0.00105f
C11191 output33/a_27_47# _175_/a_68_297# 0.001f
C11192 trimb[3] net39 0.0114f
C11193 _328_/a_1283_21# _025_ 6.78e-21
C11194 _264_/a_27_297# clkbuf_2_3__f_clk/a_110_47# 4.03e-20
C11195 _328_/a_27_47# clknet_2_2__leaf_clk 0.629f
C11196 _304_/a_761_289# clknet_2_3__leaf_clk 0.00101f
C11197 _113_ _058_ 0.00723f
C11198 _303_/a_1108_47# fanout47/a_27_47# 0.0021f
C11199 mask\[3\] _247_/a_109_297# 0.0478f
C11200 _065_ net53 1.47e-19
C11201 _262_/a_109_297# _063_ 8.95e-19
C11202 _104_ _088_ 0.102f
C11203 clk net4 0.0808f
C11204 VPWR output8/a_27_47# 0.0726f
C11205 net45 _331_/a_448_47# 1.09e-20
C11206 _326_/a_543_47# result[5] 2.17e-19
C11207 net4 clone7/a_27_47# 2.18e-20
C11208 _035_ _339_/a_27_47# 2.25e-20
C11209 _215_/a_109_297# _081_ 7.96e-20
C11210 _237_/a_76_199# _096_ 1.91e-19
C11211 _325_/a_27_47# net26 9.87e-21
C11212 net13 _319_/a_1108_47# 3.56e-36
C11213 net49 _333_/a_1217_47# 1.84e-19
C11214 net25 _146_/a_150_297# 2.14e-19
C11215 mask\[3\] _146_/a_68_297# 0.0153f
C11216 _340_/a_956_413# _122_ 3.06e-19
C11217 _337_/a_543_47# clknet_0_clk 1.84e-19
C11218 net47 _338_/a_1602_47# 0.0528f
C11219 _293_/a_299_297# _129_ 0.00178f
C11220 _338_/a_27_47# _338_/a_476_47# -0.014f
C11221 _338_/a_193_47# _338_/a_652_21# -0.00688f
C11222 _059_ _235_/a_382_297# 5.19e-20
C11223 en_co_clk _195_/a_76_199# 0.0344f
C11224 result[2] result[3] 0.037f
C11225 _107_ _049_ 0.0962f
C11226 _340_/a_193_47# net18 1.81e-20
C11227 _112_ _109_ 0.00155f
C11228 _104_ _335_/a_1283_21# 8.76e-20
C11229 _327_/a_805_47# _108_ 1.45e-19
C11230 _050_ _170_/a_299_297# 0.00539f
C11231 _326_/a_193_47# output14/a_27_47# 3.39e-21
C11232 _335_/a_27_47# _330_/a_193_47# 0.00461f
C11233 _110_ _279_/a_314_297# 0.004f
C11234 _327_/a_639_47# _111_ 1.76e-19
C11235 _340_/a_193_47# _129_ 0.00163f
C11236 net43 _079_ 2.56e-19
C11237 clk _073_ 0.00414f
C11238 _282_/a_68_297# _121_ 8.78e-19
C11239 _042_ _248_/a_27_297# 5.2e-19
C11240 VPWR _319_/a_761_289# 0.0207f
C11241 _262_/a_27_47# clknet_2_2__leaf_clk 7.63e-20
C11242 _313_/a_639_47# _010_ 5e-19
C11243 _104_ _108_ 0.0175f
C11244 _293_/a_299_297# _339_/a_1032_413# 4.14e-20
C11245 calibrate cal 0.0111f
C11246 state\[2\] calibrate 0.62f
C11247 _074_ net1 0.0392f
C11248 VPWR _243_/a_373_47# -4.51e-19
C11249 net45 _016_ 0.0528f
C11250 trim[4] net37 0.00207f
C11251 _141_/a_27_47# net51 3.52e-20
C11252 _326_/a_27_47# _314_/a_27_47# 0.002f
C11253 VPWR _197_/a_199_47# 5.18e-19
C11254 _340_/a_1032_413# _339_/a_193_47# 2.36e-20
C11255 _340_/a_476_47# _339_/a_476_47# 0.00255f
C11256 _340_/a_193_47# _339_/a_1032_413# 1.02e-20
C11257 _303_/a_27_47# _035_ 1.88e-19
C11258 _327_/a_27_47# trim_mask\[1\] 6.42e-19
C11259 _316_/a_27_47# _316_/a_639_47# -0.0015f
C11260 _187_/a_212_413# en_co_clk 0.0132f
C11261 _043_ _303_/a_193_47# 5.52e-19
C11262 _136_ _298_/a_493_297# 1.66e-20
C11263 _302_/a_109_297# clknet_2_3__leaf_clk 7.57e-20
C11264 _330_/a_448_47# _027_ 0.0145f
C11265 _330_/a_1108_47# net46 -0.00525f
C11266 output14/a_27_47# _314_/a_651_413# 1.74e-19
C11267 ctlp[0] _314_/a_193_47# 0.00268f
C11268 net31 en_co_clk 2.05e-20
C11269 net43 _319_/a_1108_47# -0.0178f
C11270 _168_/a_297_47# trim_mask\[4\] 3.87e-19
C11271 _144_/a_27_47# _339_/a_1602_47# 2.69e-19
C11272 VPWR _202_/a_382_297# 2.11e-19
C11273 _058_ trim_val\[1\] 7.73e-19
C11274 _259_/a_27_297# trim_mask\[1\] 6.42e-20
C11275 _323_/a_1270_413# net47 -3.58e-20
C11276 _199_/a_109_297# _065_ 0.00221f
C11277 VPWR _336_/a_448_47# 0.00103f
C11278 _106_ _261_/a_113_47# 7.22e-21
C11279 _050_ _192_/a_174_21# 0.00136f
C11280 _328_/a_1217_47# clknet_2_2__leaf_clk 1.2e-21
C11281 VPWR _304_/a_1283_21# 0.0435f
C11282 mask\[3\] _018_ 0.163f
C11283 _340_/a_27_47# cal_count\[3\] 1.3e-20
C11284 _107_ _262_/a_193_297# 0.00229f
C11285 _340_/a_1032_413# clknet_2_3__leaf_clk 9.51e-21
C11286 _136_ net18 0.0321f
C11287 _341_/a_543_47# _038_ 0.0078f
C11288 _341_/a_651_413# _136_ 0.00138f
C11289 _255_/a_27_47# _048_ 0.00344f
C11290 net45 _028_ 0.0283f
C11291 _094_ net15 0.00573f
C11292 _235_/a_79_21# _094_ 0.00594f
C11293 net51 _208_/a_76_199# 0.00203f
C11294 _325_/a_1283_21# _022_ 4.61e-20
C11295 _325_/a_639_47# mask\[6\] 0.00432f
C11296 _284_/a_68_297# net18 0.00837f
C11297 _319_/a_1283_21# _101_ 8.24e-20
C11298 _319_/a_27_47# _016_ 0.0228f
C11299 net25 net26 0.00158f
C11300 _325_/a_193_47# _078_ 7.8e-19
C11301 _270_/a_59_75# _265_/a_81_21# 0.00111f
C11302 _037_ _122_ 0.00898f
C11303 _241_/a_388_297# net30 3.79e-19
C11304 net54 _232_/a_114_297# 0.003f
C11305 _060_ _232_/a_32_297# 0.0107f
C11306 _303_/a_1283_21# _067_ 2.4e-21
C11307 _303_/a_1283_21# _070_ 2.2e-20
C11308 _239_/a_27_297# _092_ 0.0722f
C11309 _239_/a_474_297# _095_ 2.97e-20
C11310 mask\[6\] _158_/a_68_297# 6.03e-19
C11311 _320_/a_193_47# net44 -0.0028f
C11312 _122_ _299_/a_27_413# 1.63e-20
C11313 _228_/a_79_21# _088_ 0.00196f
C11314 clkbuf_0_clk/a_110_47# clknet_2_3__leaf_clk 5.7e-20
C11315 VPWR _206_/a_206_47# -7.44e-19
C11316 trim[1] trim[4] 0.0419f
C11317 _187_/a_297_47# net40 7.44e-19
C11318 net13 _337_/a_651_413# 0.00431f
C11319 _274_/a_75_212# _273_/a_59_75# 0.00216f
C11320 _110_ _327_/a_651_413# 6.5e-21
C11321 _037_ _299_/a_27_413# 5.48e-21
C11322 _185_/a_68_297# _049_ 3.65e-19
C11323 output37/a_27_47# net34 0.0167f
C11324 _332_/a_761_289# net40 3.26e-19
C11325 _294_/a_68_297# net2 0.0191f
C11326 fanout44/a_27_47# net30 1.5e-19
C11327 VPWR _091_ 0.0978f
C11328 VPWR _256_/a_109_297# -0.0119f
C11329 ctln[4] _335_/a_193_47# 3.05e-19
C11330 VPWR _321_/a_1283_21# 0.0444f
C11331 _041_ clknet_0_clk 2.41e-20
C11332 net2 en_co_clk 0.09f
C11333 output27/a_27_47# clknet_2_1__leaf_clk 0.0124f
C11334 fanout46/a_27_47# _330_/a_1283_21# 0.00774f
C11335 trim[4] _332_/a_651_413# 1.32e-19
C11336 _041_ _339_/a_27_47# 0.0381f
C11337 VPWR _313_/a_27_47# 0.0266f
C11338 net47 _339_/a_381_47# 1.31e-20
C11339 VPWR _337_/a_1283_21# 0.0143f
C11340 _304_/a_1283_21# _063_ 0.00322f
C11341 _267_/a_59_75# _108_ 9.5e-19
C11342 _323_/a_193_47# _323_/a_448_47# -0.00482f
C11343 net13 _143_/a_150_297# 5.75e-20
C11344 ctlp[7] net43 1.17e-19
C11345 _293_/a_81_21# _128_ 3.86e-19
C11346 VPWR net32 0.258f
C11347 _316_/a_543_47# _013_ 8.33e-19
C11348 clkbuf_2_1__f_clk/a_110_47# _120_ 4.98e-20
C11349 _192_/a_27_47# _092_ 0.0198f
C11350 _192_/a_476_47# _095_ 2.62e-21
C11351 cal_itt\[0\] _092_ 0.0807f
C11352 state\[2\] _170_/a_384_47# 8.2e-20
C11353 _090_ _096_ 0.285f
C11354 _335_/a_27_47# _335_/a_193_47# -2.27e-31
C11355 output20/a_27_47# net21 4.43e-21
C11356 _015_ _318_/a_193_47# 0.0373f
C11357 _038_ clknet_2_3__leaf_clk 0.0816f
C11358 VPWR _302_/a_373_47# -7.36e-19
C11359 _032_ _057_ 3.05e-20
C11360 _149_/a_68_297# net19 0.013f
C11361 _291_/a_285_297# net33 0.00361f
C11362 _306_/a_193_47# net2 1.04e-20
C11363 _106_ _119_ 0.00412f
C11364 state\[2\] _239_/a_27_297# 3.98e-20
C11365 _074_ net15 0.00832f
C11366 _215_/a_109_297# net14 0.00101f
C11367 _306_/a_1108_47# _305_/a_27_47# 1.65e-19
C11368 _306_/a_1283_21# _305_/a_193_47# 0.00444f
C11369 _323_/a_193_47# net18 6.64e-20
C11370 _263_/a_79_21# _206_/a_27_93# 4.86e-19
C11371 _134_ net34 1.5e-20
C11372 VPWR _033_ 0.523f
C11373 ctln[1] net15 0.00218f
C11374 _338_/a_476_47# clknet_2_3__leaf_clk 0.0467f
C11375 _320_/a_27_47# _320_/a_1283_21# 1.78e-33
C11376 _320_/a_193_47# _320_/a_543_47# -0.0129f
C11377 _007_ _078_ 1.77e-19
C11378 net12 net13 0.0452f
C11379 _316_/a_193_47# output41/a_27_47# 9.62e-20
C11380 _104_ _170_/a_299_297# 0.021f
C11381 net47 _198_/a_27_47# 1.02e-19
C11382 VPWR _340_/a_381_47# -5.12e-19
C11383 net43 _337_/a_651_413# 1e-19
C11384 net43 _313_/a_543_47# 0.00564f
C11385 _301_/a_377_297# _134_ 0.00106f
C11386 _315_/a_761_289# _095_ 1.86e-20
C11387 _315_/a_193_47# _099_ 7.61e-21
C11388 net55 _242_/a_79_21# 0.048f
C11389 _336_/a_27_47# trim_mask\[4\] 0.229f
C11390 _336_/a_1108_47# clknet_2_2__leaf_clk 0.00144f
C11391 _078_ _249_/a_27_297# 9.33e-19
C11392 VPWR _253_/a_384_47# -6.88e-20
C11393 _128_ _144_/a_27_47# 0.00276f
C11394 _328_/a_27_47# _327_/a_448_47# 9.89e-21
C11395 ctlp[0] _074_ 0.00279f
C11396 net34 _130_ 0.0128f
C11397 _308_/a_27_47# _307_/a_27_47# 5.57e-19
C11398 _091_ _063_ 0.0143f
C11399 _232_/a_32_297# en_co_clk 0.00613f
C11400 mask\[3\] _078_ 0.157f
C11401 _161_/a_68_297# _332_/a_1108_47# 5.3e-19
C11402 _190_/a_655_47# cal_itt\[3\] 1.55e-20
C11403 _306_/a_1108_47# net51 1.37e-21
C11404 _327_/a_1108_47# net9 0.00184f
C11405 _321_/a_448_47# _101_ 0.0198f
C11406 output22/a_27_47# _308_/a_193_47# 2.68e-19
C11407 _338_/a_1140_413# net18 3.91e-19
C11408 net37 _108_ 1.02e-19
C11409 _134_ _299_/a_298_297# 4.26e-21
C11410 _320_/a_1462_47# net44 4.31e-19
C11411 _303_/a_27_47# _041_ 2.19e-19
C11412 net47 _303_/a_651_413# 7.12e-19
C11413 _303_/a_1283_21# _338_/a_27_47# 7.36e-19
C11414 _065_ _205_/a_27_47# 0.0507f
C11415 _337_/a_193_47# _263_/a_297_47# 1.46e-20
C11416 _336_/a_651_413# net19 0.00269f
C11417 net13 net44 0.217f
C11418 _328_/a_1108_47# _058_ 0.00215f
C11419 _123_ en_co_clk 5.23e-20
C11420 _335_/a_1108_47# net46 0.0319f
C11421 net15 _247_/a_109_47# 9.36e-19
C11422 _304_/a_1108_47# net19 1.83e-21
C11423 clk _331_/a_761_289# 0.00262f
C11424 _290_/a_27_413# _125_ 0.0449f
C11425 _053_ _171_/a_27_47# 0.0358f
C11426 _238_/a_75_212# net1 1.02e-19
C11427 net12 _322_/a_193_47# 3.45e-20
C11428 net12 _331_/a_193_47# 1.35e-19
C11429 _299_/a_298_297# _130_ 0.0196f
C11430 trim_mask\[0\] _119_ 0.0387f
C11431 net28 _313_/a_805_47# 0.0021f
C11432 VPWR _215_/a_109_297# -0.00105f
C11433 _333_/a_193_47# _173_/a_27_47# 1.92e-19
C11434 VPWR _258_/a_27_297# 0.0163f
C11435 _026_ _258_/a_27_297# 0.00217f
C11436 VPWR _024_ 0.201f
C11437 _048_ _096_ 0.021f
C11438 VPWR _147_/a_27_47# 0.0915f
C11439 net46 rebuffer2/a_75_212# 2.15e-19
C11440 VPWR rstn 0.124f
C11441 _324_/a_761_289# net44 0.011f
C11442 clknet_2_0__leaf_clk _092_ 0.144f
C11443 _014_ _099_ 0.0359f
C11444 net45 _095_ 0.0222f
C11445 _332_/a_1283_21# net46 0.00368f
C11446 net4 _198_/a_109_47# 1.92e-19
C11447 mask\[6\] _084_ 0.0364f
C11448 _110_ _330_/a_1108_47# 0.0152f
C11449 _116_ _330_/a_1283_21# 1.78e-20
C11450 _111_ net46 0.00637f
C11451 _033_ _063_ 1.18e-21
C11452 _324_/a_193_47# _323_/a_27_47# 0.00123f
C11453 _041_ _339_/a_586_47# 0.0018f
C11454 _143_/a_68_297# _101_ 1.1e-20
C11455 _137_/a_68_297# _039_ 6.66e-19
C11456 VPWR _313_/a_1217_47# 3.99e-20
C11457 _078_ _220_/a_113_297# 0.0161f
C11458 net13 _003_ 1.12e-20
C11459 _256_/a_27_297# clknet_2_2__leaf_clk 0.0116f
C11460 _336_/a_651_413# _107_ 5.99e-19
C11461 net2 _286_/a_76_199# 2.09e-21
C11462 _109_ net33 9.17e-21
C11463 _064_ cal_itt\[1\] 0.00142f
C11464 _298_/a_215_47# _133_ 0.00284f
C11465 _304_/a_1108_47# _001_ 6.56e-21
C11466 _050_ _336_/a_193_47# 9.32e-20
C11467 net12 net43 0.00841f
C11468 result[0] _307_/a_193_47# 0.001f
C11469 cal _315_/a_27_47# 0.00255f
C11470 _253_/a_384_47# net52 8.16e-20
C11471 _322_/a_193_47# net44 0.00495f
C11472 _185_/a_68_297# state\[1\] 2.14e-19
C11473 _074_ _310_/a_193_47# 0.015f
C11474 mask\[4\] _150_/a_27_47# 0.049f
C11475 _314_/a_193_47# _224_/a_113_297# 1.97e-19
C11476 _339_/a_27_47# _129_ 4.2e-20
C11477 net47 _297_/a_129_47# 2.49e-20
C11478 trim_mask\[0\] _087_ 3.44e-21
C11479 _233_/a_109_297# _074_ 0.00526f
C11480 _233_/a_27_297# calibrate 0.0455f
C11481 _065_ _095_ 0.178f
C11482 trim_mask\[1\] net40 8.96e-22
C11483 _046_ _313_/a_448_47# 1.64e-19
C11484 net21 _313_/a_1283_21# 0.00744f
C11485 state\[2\] _318_/a_1270_413# 8.41e-20
C11486 _290_/a_27_413# net40 1.87e-20
C11487 _134_ _133_ 0.00631f
C11488 _301_/a_377_297# cal_count\[3\] 6.02e-20
C11489 _303_/a_651_413# net44 3.05e-19
C11490 _051_ _089_ 0.00231f
C11491 _326_/a_805_47# _074_ 5.87e-19
C11492 trim[1] _108_ 3.27e-19
C11493 net31 cal_count\[0\] 6.25e-20
C11494 _341_/a_193_47# cal_count\[3\] 0.547f
C11495 VPWR _338_/a_1032_413# -0.00127f
C11496 _338_/a_1224_47# clknet_2_3__leaf_clk 1.82e-19
C11497 input2/a_27_47# _132_ 0.00127f
C11498 _341_/a_448_47# clknet_2_3__leaf_clk 0.016f
C11499 result[4] _078_ 5.53e-20
C11500 state\[0\] _192_/a_476_47# 3.57e-20
C11501 _323_/a_1108_47# _303_/a_193_47# 0.00107f
C11502 _323_/a_543_47# _303_/a_543_47# 1.15e-19
C11503 _323_/a_1283_21# _303_/a_761_289# 2.87e-20
C11504 _323_/a_448_47# _303_/a_27_47# 1.6e-20
C11505 cal_itt\[1\] _053_ 0.00161f
C11506 net50 _256_/a_109_297# 0.0024f
C11507 trim[1] trim[0] 0.0363f
C11508 net43 net44 0.0814f
C11509 clknet_2_0__leaf_clk _246_/a_109_297# 1.16e-20
C11510 _315_/a_1462_47# _099_ 5.67e-20
C11511 _339_/a_27_47# _339_/a_1032_413# -0.00554f
C11512 _339_/a_193_47# _339_/a_1182_261# -2.22e-21
C11513 _130_ _133_ 3.75e-19
C11514 _336_/a_1217_47# trim_mask\[4\] 9.77e-19
C11515 net13 _320_/a_543_47# 0.00303f
C11516 _306_/a_651_413# clknet_2_1__leaf_clk 7.92e-19
C11517 _276_/a_59_75# _335_/a_27_47# 0.00105f
C11518 _330_/a_27_47# net30 6.12e-20
C11519 _187_/a_212_413# _061_ 0.0509f
C11520 trim_mask\[1\] _334_/a_27_47# 1.41e-20
C11521 trim_val\[1\] _334_/a_193_47# 5.84e-22
C11522 result[5] result[7] 7.15e-19
C11523 _320_/a_27_47# _040_ 0.359f
C11524 _243_/a_109_297# _095_ 8.87e-21
C11525 _243_/a_27_297# _099_ 9.67e-21
C11526 _271_/a_75_212# _030_ 0.00288f
C11527 cal clknet_2_0__leaf_clk 0.00552f
C11528 clknet_2_1__leaf_clk _314_/a_761_289# 4.07e-20
C11529 output29/a_27_47# _085_ 9.81e-20
C11530 _307_/a_193_47# net14 0.0105f
C11531 _336_/a_448_47# _279_/a_396_47# 6.19e-19
C11532 _326_/a_193_47# net29 1.03e-19
C11533 VPWR _316_/a_1270_413# -1.11e-34
C11534 net31 _061_ 1.31e-19
C11535 _332_/a_651_413# _108_ 0.00129f
C11536 ctlp[6] VPWR 0.445f
C11537 fanout46/a_27_47# _108_ 1.48e-20
C11538 _135_ net46 6e-20
C11539 _029_ _332_/a_1108_47# 5.34e-21
C11540 _050_ net55 0.128f
C11541 _032_ _027_ 5.79e-20
C11542 _104_ _277_/a_75_212# 3.86e-19
C11543 _146_/a_150_297# _310_/a_193_47# 1.9e-20
C11544 VPWR output37/a_27_47# 0.0992f
C11545 fanout43/a_27_47# _078_ 0.053f
C11546 net43 _003_ 0.00181f
C11547 _120_ net30 1.38e-19
C11548 VPWR _320_/a_27_47# 0.0148f
C11549 fanout44/a_27_47# _319_/a_1108_47# 7.24e-20
C11550 _339_/a_1602_47# _133_ 6.44e-21
C11551 net12 _322_/a_1462_47# 3.73e-19
C11552 _286_/a_76_199# _123_ 0.0152f
C11553 net27 _078_ 0.445f
C11554 net50 _033_ 2.07e-20
C11555 mask\[6\] _085_ 0.023f
C11556 _162_/a_27_47# trim_val\[0\] 6.71e-21
C11557 _333_/a_448_47# net32 6.05e-20
C11558 net15 net26 0.0071f
C11559 _322_/a_27_47# _320_/a_1283_21# 0.00137f
C11560 _078_ _222_/a_113_297# 0.00237f
C11561 _175_/a_68_297# _172_/a_68_297# 0.0129f
C11562 net7 _317_/a_761_289# 4.61e-20
C11563 _333_/a_193_47# _172_/a_68_297# 3.32e-19
C11564 _076_ net30 0.0106f
C11565 net49 net37 1.62e-19
C11566 net2 cal_count\[0\] 1.05e-19
C11567 net22 _120_ 0.00171f
C11568 _136_ _265_/a_81_21# 8.24e-20
C11569 output12/a_27_47# net11 0.00102f
C11570 _269_/a_299_297# _108_ 9.71e-20
C11571 clone1/a_27_47# _092_ 1.19e-19
C11572 _078_ rebuffer5/a_161_47# 5.39e-19
C11573 VPWR _307_/a_193_47# 0.0143f
C11574 VPWR _323_/a_651_413# -0.00809f
C11575 _290_/a_207_413# net37 0.0104f
C11576 output31/a_27_47# trim_mask\[1\] 0.00105f
C11577 trim[0] _269_/a_299_297# 1.79e-19
C11578 _322_/a_1462_47# net44 9.59e-19
C11579 VPWR _298_/a_215_47# 0.005f
C11580 _329_/a_761_289# _026_ 7.06e-19
C11581 state\[0\] net45 0.00434f
C11582 _314_/a_651_413# net29 9.55e-19
C11583 _309_/a_1283_21# _308_/a_1283_21# 4.89e-20
C11584 _309_/a_193_47# _308_/a_651_413# 4.01e-21
C11585 _309_/a_651_413# _308_/a_193_47# 2.17e-21
C11586 _300_/a_377_297# _135_ 4.39e-19
C11587 _329_/a_761_289# VPWR 0.0193f
C11588 VPWR clkbuf_2_3__f_clk/a_110_47# 0.0504f
C11589 _074_ _012_ 0.0813f
C11590 net43 _320_/a_543_47# 1.01e-19
C11591 net23 _320_/a_27_47# 1.89e-20
C11592 _305_/a_193_47# net2 1.92e-19
C11593 _238_/a_75_212# net15 4.65e-20
C11594 _046_ _010_ 9.53e-19
C11595 _214_/a_199_47# _101_ 3.77e-19
C11596 _335_/a_448_47# _032_ 0.00455f
C11597 _015_ _243_/a_373_47# 5.24e-19
C11598 _313_/a_193_47# _155_/a_68_297# 5.89e-21
C11599 output20/a_27_47# _045_ 6.23e-19
C11600 _305_/a_27_47# _305_/a_1108_47# -2.98e-20
C11601 _299_/a_27_413# _297_/a_285_47# 4.23e-20
C11602 _062_ _049_ 0.0151f
C11603 VPWR _134_ 0.374f
C11604 _325_/a_543_47# _313_/a_543_47# 0.00153f
C11605 _061_ net2 1.78e-19
C11606 _112_ net46 0.00936f
C11607 _272_/a_299_297# net46 0.00102f
C11608 net44 _312_/a_1108_47# 0.0107f
C11609 _306_/a_193_47# mask\[0\] 7.13e-21
C11610 VPWR _341_/a_1270_413# -2.31e-19
C11611 trim_mask\[3\] _258_/a_109_297# 0.00149f
C11612 net50 _258_/a_27_297# 0.00128f
C11613 _310_/a_543_47# net29 4.49e-22
C11614 _323_/a_27_47# _000_ 4.43e-20
C11615 state\[0\] _065_ 2.46e-21
C11616 net50 _024_ 2.32e-20
C11617 net14 output41/a_27_47# 0.00326f
C11618 _320_/a_27_47# net52 0.00489f
C11619 _013_ valid 6.4e-21
C11620 clknet_2_1__leaf_clk _311_/a_27_47# 0.0322f
C11621 clknet_2_0__leaf_clk _017_ 0.123f
C11622 _303_/a_1283_21# clknet_2_3__leaf_clk 0.0739f
C11623 _319_/a_639_47# _092_ 1.66e-20
C11624 _117_ _335_/a_543_47# 1.78e-19
C11625 _110_ _335_/a_1108_47# 1.75e-19
C11626 VPWR _130_ 0.239f
C11627 _271_/a_75_212# trim_mask\[1\] 0.118f
C11628 _321_/a_1108_47# _248_/a_109_297# 2.52e-19
C11629 net43 _307_/a_1283_21# 2.34e-20
C11630 _114_ _334_/a_193_47# 5.54e-20
C11631 trim_val\[2\] _334_/a_1283_21# 0.00479f
C11632 _076_ _072_ 0.00276f
C11633 _320_/a_1217_47# _040_ 0.00102f
C11634 net13 ctln[7] 0.0872f
C11635 VPWR _308_/a_448_47# 0.00314f
C11636 _078_ sample 1.76e-19
C11637 _033_ _279_/a_396_47# 0.00101f
C11638 _065_ _208_/a_218_374# 0.00203f
C11639 _306_/a_543_47# cal_itt\[3\] 3.33e-19
C11640 _306_/a_761_289# _072_ 1.19e-19
C11641 _337_/a_27_47# _092_ 0.00189f
C11642 _337_/a_193_47# _099_ 7.41e-21
C11643 net3 _316_/a_27_47# 1.24e-19
C11644 _110_ rebuffer2/a_75_212# 9.17e-19
C11645 net16 _334_/a_1283_21# 0.00492f
C11646 net26 _310_/a_193_47# 8.49e-20
C11647 _250_/a_27_297# _074_ 3.55e-20
C11648 VPWR _237_/a_505_21# 0.0644f
C11649 output41/a_27_47# net41 0.028f
C11650 state\[2\] clone1/a_27_47# 0.0082f
C11651 _042_ _310_/a_1108_47# 1.99e-19
C11652 _239_/a_474_297# _052_ 1.88e-19
C11653 trim[1] net49 1.86e-19
C11654 _110_ _111_ 0.00137f
C11655 state\[0\] _243_/a_109_297# 1.27e-19
C11656 _325_/a_193_47# mask\[7\] 1.79e-19
C11657 _325_/a_27_47# _102_ 3.99e-21
C11658 VPWR _320_/a_1217_47# 2.71e-20
C11659 _090_ _098_ 1.75e-19
C11660 _060_ _100_ 0.312f
C11661 net54 _096_ 0.376f
C11662 VPWR _339_/a_1602_47# 0.0182f
C11663 output9/a_27_47# net46 1.71e-19
C11664 cal_count\[0\] _123_ 0.206f
C11665 _063_ clkbuf_2_3__f_clk/a_110_47# 0.0504f
C11666 _104_ _336_/a_193_47# 0.287f
C11667 clknet_2_1__leaf_clk _310_/a_639_47# 9.94e-19
C11668 comp net33 3.24e-19
C11669 _137_/a_68_297# _049_ 1.37e-19
C11670 _058_ _264_/a_27_297# 0.0014f
C11671 _133_ _297_/a_377_297# 8.42e-19
C11672 output31/a_27_47# output33/a_27_47# 0.0523f
C11673 fanout44/a_27_47# _337_/a_651_413# 5.72e-20
C11674 net34 _175_/a_150_297# 2.58e-19
C11675 _326_/a_27_47# _078_ 0.00936f
C11676 VPWR output41/a_27_47# 0.0793f
C11677 _333_/a_1283_21# _055_ 0.0274f
C11678 clknet_0_clk _090_ 9.53e-21
C11679 net13 _322_/a_543_47# 0.00836f
C11680 _128_ _133_ 5.69e-19
C11681 VPWR rebuffer6/a_27_47# 0.067f
C11682 _041_ _209_/a_27_47# 3.39e-20
C11683 _308_/a_448_47# net23 5e-20
C11684 _308_/a_639_47# net43 7.29e-19
C11685 net9 _334_/a_1108_47# 2.52e-20
C11686 net3 net44 1.09e-20
C11687 _322_/a_27_47# _040_ 1.61e-20
C11688 _337_/a_1283_21# _034_ 7.08e-20
C11689 _005_ net14 8.37e-20
C11690 net48 rebuffer1/a_75_212# 0.00258f
C11691 _112_ _332_/a_448_47# 1.93e-19
C11692 VPWR _324_/a_193_47# 0.0328f
C11693 clkbuf_2_2__f_clk/a_110_47# net19 0.0269f
C11694 VPWR _307_/a_1462_47# 2.57e-19
C11695 _309_/a_193_47# net43 0.00412f
C11696 VPWR cal_count\[3\] 2.62f
C11697 _187_/a_212_413# net16 0.00604f
C11698 _327_/a_448_47# _256_/a_27_297# 6.81e-19
C11699 _053_ _304_/a_193_47# 0.00902f
C11700 _309_/a_639_47# net14 0.00144f
C11701 _107_ _240_/a_109_297# 2.8e-19
C11702 trim_mask\[3\] clkbuf_2_2__f_clk/a_110_47# 1.5e-20
C11703 cal_itt\[1\] _195_/a_218_47# 1.04e-19
C11704 _308_/a_1283_21# _016_ 1.83e-20
C11705 cal_itt\[0\] _195_/a_439_47# 7.96e-19
C11706 net16 _332_/a_193_47# 0.0169f
C11707 VPWR _322_/a_27_47# 0.0662f
C11708 _074_ _009_ 0.00872f
C11709 _329_/a_193_47# clknet_2_2__leaf_clk 0.00122f
C11710 clknet_2_1__leaf_clk _247_/a_373_47# 1.25e-19
C11711 VPWR _257_/a_27_297# 0.0314f
C11712 VPWR _331_/a_27_47# 0.0349f
C11713 _314_/a_27_47# _086_ 0.00916f
C11714 net31 net16 4.4e-20
C11715 _311_/a_543_47# net26 0.0301f
C11716 _325_/a_27_47# _010_ 5.33e-19
C11717 _233_/a_27_297# _315_/a_27_47# 1.81e-19
C11718 _309_/a_27_47# _101_ 5.47e-20
C11719 trim_mask\[0\] _182_/a_27_47# 2.95e-19
C11720 _322_/a_193_47# _322_/a_543_47# -0.0181f
C11721 clkbuf_2_2__f_clk/a_110_47# _107_ 0.00242f
C11722 _331_/a_27_47# _331_/a_1283_21# -9.15e-20
C11723 _331_/a_193_47# _331_/a_543_47# -0.00702f
C11724 net10 net18 0.139f
C11725 VPWR _303_/a_448_47# 0.00107f
C11726 _104_ net55 0.0665f
C11727 _269_/a_81_21# _112_ 0.00251f
C11728 _269_/a_299_297# net49 0.00153f
C11729 _269_/a_384_47# trim_mask\[1\] 0.00147f
C11730 _048_ _098_ 0.127f
C11731 _323_/a_1270_413# net19 1.39e-19
C11732 trim_mask\[0\] _099_ 8.74e-21
C11733 _327_/a_27_47# _136_ 0.00263f
C11734 clknet_2_2__leaf_clk net18 0.123f
C11735 net9 _332_/a_761_289# 8.16e-20
C11736 VPWR _005_ 0.096f
C11737 _282_/a_68_297# _095_ 4.78e-19
C11738 _068_ net30 0.00285f
C11739 _036_ _339_/a_1602_47# 1.37e-20
C11740 _048_ clknet_0_clk 0.0719f
C11741 _237_/a_505_21# _164_/a_161_47# 0.00601f
C11742 trim_mask\[4\] _098_ 1.66e-20
C11743 _329_/a_543_47# trim_mask\[3\] 0.00103f
C11744 _230_/a_145_75# en_co_clk 1.15e-19
C11745 VPWR _219_/a_109_297# 0.00228f
C11746 _051_ _092_ 0.0918f
C11747 net43 _322_/a_543_47# 2.97e-20
C11748 _113_ net16 0.00136f
C11749 _004_ sample 0.0175f
C11750 _078_ _310_/a_761_289# 1.96e-19
C11751 _064_ _302_/a_27_297# 3.11e-19
C11752 VPWR _309_/a_639_47# 4.66e-19
C11753 net37 output5/a_27_47# 6.9e-20
C11754 en_co_clk _100_ 8.95e-19
C11755 _328_/a_1270_413# net46 -2.06e-19
C11756 _050_ _121_ 4.53e-21
C11757 mask\[7\] mask\[3\] 5.1e-19
C11758 _102_ net25 2.7e-20
C11759 output25/a_27_47# result[3] 0.0103f
C11760 cal_count\[3\] _063_ 0.168f
C11761 _292_/a_78_199# _128_ 0.0854f
C11762 clknet_0_clk trim_mask\[4\] 0.0177f
C11763 _064_ _106_ 0.00126f
C11764 _336_/a_1283_21# _330_/a_1108_47# 8.54e-21
C11765 _336_/a_1108_47# _330_/a_1283_21# 1.45e-19
C11766 _169_/a_109_53# _051_ 0.0198f
C11767 net12 _249_/a_109_47# 8.77e-19
C11768 fanout44/a_27_47# net44 0.00684f
C11769 _328_/a_193_47# _030_ 0.0025f
C11770 _322_/a_761_289# _101_ 0.00355f
C11771 _326_/a_1217_47# _078_ 2.97e-20
C11772 _322_/a_27_47# net52 1.87e-19
C11773 clkc net40 1.65e-19
C11774 clkbuf_2_2__f_clk/a_110_47# _279_/a_27_47# 8.19e-20
C11775 _251_/a_27_297# net29 5.81e-21
C11776 net2 net16 0.203f
C11777 net9 _030_ 3.65e-20
C11778 net4 _190_/a_655_47# 0.00167f
C11779 _005_ net23 0.0439f
C11780 VPWR _128_ 0.554f
C11781 _305_/a_761_289# net30 1.72e-20
C11782 _053_ _302_/a_27_297# 0.0625f
C11783 _238_/a_75_212# _012_ 1.22e-19
C11784 net45 _052_ 1.21e-19
C11785 _321_/a_543_47# mask\[2\] 6.01e-19
C11786 VPWR _324_/a_1462_47# 3.61e-19
C11787 _110_ _112_ 0.154f
C11788 _110_ _272_/a_299_297# 1.47e-19
C11789 net25 _006_ 1.92e-19
C11790 _068_ _072_ 0.015f
C11791 _293_/a_299_297# _125_ 2.07e-19
C11792 _309_/a_1462_47# net43 -9.14e-19
C11793 output8/a_27_47# _334_/a_1108_47# 0.00177f
C11794 net8 _334_/a_193_47# 0.0163f
C11795 mask\[0\] _039_ 0.0317f
C11796 _327_/a_1270_413# trim_mask\[0\] 7.89e-20
C11797 _327_/a_1108_47# _024_ 0.00102f
C11798 net4 trim_val\[4\] 0.0023f
C11799 _053_ _106_ 8.4e-19
C11800 _195_/a_535_374# _065_ 1.25e-20
C11801 _305_/a_805_47# _002_ 0.0023f
C11802 net16 _332_/a_1462_47# 2.04e-19
C11803 _103_ _052_ 9.12e-20
C11804 fanout44/a_27_47# _003_ 1.15e-19
C11805 _316_/a_1283_21# _092_ 4.55e-19
C11806 clkbuf_2_0__f_clk/a_110_47# net30 0.0321f
C11807 VPWR _322_/a_1217_47# 7.57e-20
C11808 _329_/a_1462_47# clknet_2_2__leaf_clk 4.85e-19
C11809 VPWR _331_/a_1217_47# 6.18e-20
C11810 _250_/a_27_297# net26 2.73e-20
C11811 _312_/a_761_289# net20 0.0042f
C11812 _214_/a_113_297# mask\[1\] 0.0423f
C11813 _323_/a_193_47# _249_/a_27_297# 1.81e-20
C11814 VPWR net21 0.509f
C11815 _308_/a_761_289# _212_/a_113_297# 0.00133f
C11816 _074_ _315_/a_543_47# 0.016f
C11817 calibrate _315_/a_761_289# 0.0238f
C11818 _093_ _315_/a_193_47# 1.05e-19
C11819 state\[2\] _051_ 0.601f
C11820 _309_/a_1217_47# _101_ 9.27e-21
C11821 _064_ trim_mask\[0\] 0.303f
C11822 _161_/a_150_297# net33 3.83e-19
C11823 _257_/a_373_47# _025_ -1.67e-20
C11824 _324_/a_761_289# net19 2.59e-19
C11825 clkbuf_2_3__f_clk/a_110_47# _279_/a_396_47# 6.1e-19
C11826 _331_/a_543_47# _260_/a_93_21# 7.88e-19
C11827 VPWR _000_ 0.0391f
C11828 _317_/a_27_47# _317_/a_193_47# -0.0061f
C11829 trim_val\[2\] trim_val\[1\] 0.0161f
C11830 VPWR _312_/a_1283_21# 0.0467f
C11831 _327_/a_1217_47# _136_ 7.17e-20
C11832 _277_/a_75_212# fanout46/a_27_47# 3e-19
C11833 _232_/a_32_297# _049_ 0.0148f
C11834 _320_/a_193_47# mask\[1\] 0.402f
C11835 _305_/a_761_289# _072_ 0.0264f
C11836 _305_/a_543_47# cal_itt\[3\] 6.56e-19
C11837 clkbuf_2_0__f_clk/a_110_47# net22 1.84e-20
C11838 net13 _107_ 5.96e-20
C11839 _078_ net51 0.00111f
C11840 output31/a_27_47# _056_ 1.1e-19
C11841 net31 _176_/a_27_47# 5.31e-19
C11842 _321_/a_193_47# _085_ 3.94e-21
C11843 _198_/a_27_47# net19 0.00225f
C11844 net15 net55 1.07e-20
C11845 _235_/a_79_21# net55 0.013f
C11846 net13 _166_/a_161_47# 1.58e-19
C11847 _111_ rebuffer3/a_75_212# 1.05e-21
C11848 en net14 0.0186f
C11849 result[4] mask\[7\] 5.8e-20
C11850 net16 trim_val\[1\] 0.0116f
C11851 _293_/a_299_297# net40 0.0103f
C11852 _331_/a_193_47# net19 0.00104f
C11853 net50 cal_count\[3\] 0.0229f
C11854 _189_/a_27_47# cal_itt\[3\] 2.17e-19
C11855 _087_ _089_ 0.0912f
C11856 VPWR _242_/a_297_47# -0.00207f
C11857 _228_/a_79_21# net55 3.8e-20
C11858 _058_ net34 7.39e-20
C11859 _323_/a_27_47# mask\[4\] 0.00764f
C11860 trim_mask\[0\] _053_ 0.396f
C11861 _303_/a_805_47# _000_ 3.81e-19
C11862 _283_/a_75_212# clknet_0_clk 0.00409f
C11863 net16 _123_ 0.036f
C11864 clknet_0_clk _190_/a_27_47# 0.0106f
C11865 result[2] _074_ 0.00705f
C11866 output35/a_27_47# _136_ 4.5e-19
C11867 _059_ _337_/a_1283_21# 4.91e-20
C11868 net33 net46 0.0155f
C11869 trim_mask\[3\] _257_/a_109_297# 1.15e-19
C11870 _337_/a_1270_413# en_co_clk 7.91e-20
C11871 net50 _257_/a_27_297# 0.00549f
C11872 _093_ _014_ 0.0073f
C11873 calibrate net45 0.157f
C11874 _303_/a_651_413# net19 0.00477f
C11875 _128_ _036_ 0.0103f
C11876 _312_/a_27_47# _312_/a_193_47# -0.009f
C11877 _074_ _211_/a_109_297# 0.00107f
C11878 _328_/a_193_47# trim_mask\[1\] 0.554f
C11879 _336_/a_761_289# net46 -0.00669f
C11880 VPWR _175_/a_150_297# 1.52e-19
C11881 net5 _187_/a_27_413# 1.94e-19
C11882 _024_ _193_/a_109_297# 1.86e-19
C11883 net1 _316_/a_543_47# 1.71e-20
C11884 VPWR _333_/a_761_289# 0.0104f
C11885 _227_/a_209_311# _049_ 0.0102f
C11886 net9 trim_mask\[1\] 0.00869f
C11887 net43 net19 4.36e-20
C11888 _219_/a_109_297# _083_ 3.99e-21
C11889 _341_/a_1283_21# _092_ 1.81e-21
C11890 _075_ _206_/a_206_47# 0.00341f
C11891 VPWR _265_/a_299_297# 0.0793f
C11892 _103_ calibrate 0.00146f
C11893 _078_ _224_/a_199_47# 7.62e-19
C11894 _200_/a_80_21# cal_itt\[2\] 0.02f
C11895 _337_/a_651_413# _076_ 1.38e-19
C11896 calibrate _065_ 3.98e-20
C11897 mask\[7\] net27 0.0419f
C11898 _263_/a_79_21# _090_ 0.022f
C11899 net8 _334_/a_1462_47# 4.63e-19
C11900 VPWR en 0.168f
C11901 _325_/a_1108_47# net13 0.0152f
C11902 _319_/a_193_47# _244_/a_27_297# 3.22e-20
C11903 clk _330_/a_193_47# 0.00144f
C11904 _288_/a_59_75# _122_ 5.33e-20
C11905 _053_ _338_/a_652_21# 9.89e-22
C11906 net31 trimb[0] 0.00722f
C11907 output23/a_27_47# result[2] 7.83e-19
C11908 result[1] output24/a_27_47# 0.00235f
C11909 clknet_2_1__leaf_clk _225_/a_109_297# 4.44e-19
C11910 _320_/a_27_47# _141_/a_27_47# 3.45e-19
C11911 _094_ _206_/a_27_93# 3.47e-19
C11912 _250_/a_109_297# _078_ 7.17e-19
C11913 _323_/a_27_47# _020_ 0.155f
C11914 _323_/a_543_47# mask\[5\] 4.63e-19
C11915 _308_/a_651_413# mask\[1\] 2.4e-19
C11916 net54 _098_ 1.04e-19
C11917 _320_/a_1283_21# mask\[4\] 7.02e-20
C11918 _337_/a_1283_21# _075_ 0.0308f
C11919 _337_/a_1108_47# _062_ 9.67e-20
C11920 _041_ _208_/a_505_21# 3.19e-20
C11921 _321_/a_27_47# _310_/a_27_47# 5.48e-21
C11922 cal_count\[3\] _279_/a_396_47# 9.29e-19
C11923 _331_/a_1108_47# trim_mask\[4\] 0.00262f
C11924 _331_/a_639_47# _028_ 0.00129f
C11925 _331_/a_805_47# clknet_2_2__leaf_clk 8.94e-20
C11926 output31/a_27_47# _173_/a_27_47# 0.00944f
C11927 _051_ _226_/a_197_47# 2.74e-19
C11928 _093_ _243_/a_27_297# 0.0328f
C11929 calibrate _243_/a_109_297# 0.0473f
C11930 _260_/a_93_21# _260_/a_256_47# -3.48e-20
C11931 net13 _248_/a_109_297# 0.00833f
C11932 VPWR _325_/a_761_289# 0.00298f
C11933 state\[0\] _316_/a_448_47# 1.44e-20
C11934 net4 _330_/a_193_47# 2.27e-19
C11935 trim_val\[2\] _114_ 0.0134f
C11936 _041_ mask\[2\] 0.271f
C11937 clknet_2_1__leaf_clk clknet_2_0__leaf_clk 0.028f
C11938 _091_ _195_/a_505_21# 0.00583f
C11939 _116_ _277_/a_75_212# 0.0372f
C11940 net54 clknet_0_clk 4.49e-20
C11941 _325_/a_1108_47# _322_/a_193_47# 2.21e-19
C11942 _336_/a_1108_47# _108_ 2.38e-19
C11943 _136_ net40 0.0317f
C11944 net13 mask\[1\] 0.0277f
C11945 _325_/a_193_47# _159_/a_27_47# 2.65e-20
C11946 _071_ _002_ 3.17e-21
C11947 _114_ net16 8.85e-19
C11948 clkbuf_2_0__f_clk/a_110_47# _079_ 8.04e-21
C11949 _094_ _337_/a_543_47# 0.038f
C11950 _327_/a_448_47# net18 0.0021f
C11951 net13 _185_/a_68_297# 0.00304f
C11952 _284_/a_68_297# net40 2.83e-21
C11953 _253_/a_81_21# _314_/a_761_289# 1.88e-22
C11954 _035_ _286_/a_439_47# 3.12e-20
C11955 _323_/a_1217_47# mask\[4\] 5.2e-19
C11956 _323_/a_193_47# net27 1.6e-19
C11957 _318_/a_193_47# _318_/a_448_47# -0.00482f
C11958 net12 _076_ 0.619f
C11959 output10/a_27_47# trim_mask\[3\] 0.0104f
C11960 _306_/a_543_47# clk 3.57e-21
C11961 VPWR _241_/a_105_352# 0.0112f
C11962 _048_ _263_/a_79_21# 0.0191f
C11963 net12 _306_/a_761_289# 0.00389f
C11964 _320_/a_27_47# _208_/a_76_199# 3.03e-21
C11965 _136_ _267_/a_145_75# 1.14e-19
C11966 _322_/a_761_289# _248_/a_27_297# 0.00173f
C11967 _322_/a_193_47# _248_/a_109_297# 3.84e-19
C11968 _325_/a_1108_47# net43 -0.0143f
C11969 _312_/a_1108_47# net19 6.62e-19
C11970 net42 cal_itt\[3\] 2.24e-19
C11971 _232_/a_32_297# state\[1\] 8.56e-19
C11972 _168_/a_207_413# _049_ 0.00139f
C11973 _294_/a_68_297# net34 3.27e-20
C11974 _238_/a_75_212# _097_ 0.00544f
C11975 _210_/a_113_297# _315_/a_27_47# 3.34e-20
C11976 _043_ _311_/a_27_47# 8.03e-22
C11977 net34 en_co_clk 1.13e-19
C11978 _107_ _260_/a_93_21# 0.00214f
C11979 _192_/a_174_21# _192_/a_548_47# -8.51e-21
C11980 mask\[0\] _049_ 0.0198f
C11981 cal_itt\[2\] _071_ 0.441f
C11982 _322_/a_193_47# mask\[1\] 2e-21
C11983 _309_/a_543_47# mask\[3\] 0.00691f
C11984 output33/a_27_47# trim[2] 0.00959f
C11985 trim_mask\[0\] _161_/a_68_297# 0.00319f
C11986 _333_/a_193_47# clknet_2_2__leaf_clk 1e-19
C11987 net44 _076_ 0.148f
C11988 clkbuf_2_1__f_clk/a_110_47# _319_/a_1283_21# 0.00615f
C11989 _308_/a_27_47# fanout43/a_27_47# 0.00358f
C11990 input2/a_27_47# _130_ 0.0114f
C11991 _325_/a_761_289# net52 1.3e-20
C11992 _325_/a_1283_21# _101_ 0.00102f
C11993 _301_/a_377_297# en_co_clk 5.5e-20
C11994 mask\[3\] _245_/a_27_297# 1.03e-19
C11995 _102_ net15 7.88e-20
C11996 _306_/a_761_289# net44 0.00164f
C11997 _265_/a_81_21# clknet_2_2__leaf_clk 0.00101f
C11998 _256_/a_27_297# _108_ 1.48e-19
C11999 _293_/a_81_21# cal_count\[0\] 0.0585f
C12000 clkbuf_2_0__f_clk/a_110_47# _319_/a_1108_47# 1.63e-20
C12001 _326_/a_651_413# _253_/a_81_21# 6.67e-19
C12002 _326_/a_27_47# mask\[7\] 0.0131f
C12003 cal_itt\[2\] _262_/a_27_47# 1.31e-19
C12004 _341_/a_193_47# en_co_clk 5.4e-20
C12005 input1/a_75_212# output41/a_27_47# 0.00329f
C12006 _048_ clknet_2_2__leaf_clk 2.04e-20
C12007 VPWR _190_/a_215_47# -0.00217f
C12008 clkbuf_2_2__f_clk/a_110_47# _330_/a_761_289# 0.00656f
C12009 net47 _286_/a_505_21# 0.0104f
C12010 _162_/a_27_47# _108_ 0.00185f
C12011 _328_/a_193_47# _328_/a_448_47# -0.00779f
C12012 net2 _202_/a_297_47# 0.0404f
C12013 _021_ _078_ 5.51e-21
C12014 net30 cal_itt\[3\] 0.176f
C12015 _340_/a_27_47# cal_count\[0\] 3.14e-19
C12016 net43 mask\[1\] 0.144f
C12017 _119_ _279_/a_490_47# 1.7e-19
C12018 _328_/a_448_47# net9 5.07e-19
C12019 _305_/a_1283_21# _202_/a_297_47# 3e-19
C12020 _239_/a_27_297# _103_ 7.91e-19
C12021 net10 trim_mask\[4\] 5.9e-22
C12022 _033_ _335_/a_543_47# 1.35e-19
C12023 VPWR _045_ 0.29f
C12024 _076_ _003_ 0.149f
C12025 VPWR _249_/a_109_297# -0.0176f
C12026 _321_/a_448_47# _310_/a_1108_47# 2e-21
C12027 _248_/a_27_297# _101_ 0.0925f
C12028 _210_/a_113_297# clknet_2_0__leaf_clk 0.0654f
C12029 _321_/a_543_47# _074_ 4.42e-20
C12030 clknet_2_2__leaf_clk trim_mask\[4\] 0.559f
C12031 trim_mask\[4\] _260_/a_584_47# 1.83e-20
C12032 _306_/a_761_289# _003_ 2.33e-20
C12033 _306_/a_543_47# _073_ 9.17e-19
C12034 _307_/a_193_47# output30/a_27_47# 6.7e-19
C12035 VPWR _327_/a_193_47# -0.0118f
C12036 _317_/a_448_47# _014_ 0.00455f
C12037 _317_/a_761_289# state\[1\] 2.01e-19
C12038 _317_/a_651_413# clknet_2_0__leaf_clk 0.0267f
C12039 _317_/a_1108_47# net45 0.00804f
C12040 state\[0\] _013_ 7.07e-20
C12041 output31/a_27_47# _172_/a_68_297# 0.001f
C12042 _144_/a_27_47# cal_count\[0\] 0.0451f
C12043 _262_/a_205_47# net30 1.49e-19
C12044 _257_/a_109_47# trim_val\[4\] 4.68e-19
C12045 _110_ net33 1.3e-20
C12046 _322_/a_1108_47# mask\[3\] 0.057f
C12047 result[3] _007_ 0.00262f
C12048 _051_ net46 1.84e-21
C12049 net15 _121_ 0.0264f
C12050 _094_ _282_/a_150_297# 7.8e-19
C12051 _026_ _058_ 4.85e-19
C12052 _110_ _336_/a_761_289# 0.00634f
C12053 _259_/a_109_297# _026_ 1.11e-19
C12054 VPWR _058_ 1.05f
C12055 _104_ clknet_2_3__leaf_clk 1.02e-19
C12056 _259_/a_109_297# VPWR 0.00164f
C12057 net15 _010_ 0.00749f
C12058 _329_/a_27_47# _330_/a_1108_47# 2.73e-20
C12059 _125_ _339_/a_27_47# 2.29e-20
C12060 VPWR mask\[4\] 0.198f
C12061 trim_val\[0\] _333_/a_193_47# 1.49e-20
C12062 result[3] mask\[3\] 1.45e-19
C12063 _060_ net41 0.0735f
C12064 _320_/a_761_289# _077_ 4.25e-20
C12065 _030_ net32 3.33e-21
C12066 _306_/a_27_47# clknet_0_clk 1.07e-20
C12067 _265_/a_81_21# trim_val\[0\] 0.0409f
C12068 cal_itt\[3\] _072_ 0.255f
C12069 result[7] _011_ 0.00565f
C12070 _322_/a_1283_21# mask\[4\] 0.0114f
C12071 _299_/a_382_47# net40 2.78e-19
C12072 _063_ _190_/a_215_47# 0.0481f
C12073 _334_/a_193_47# net34 2.5e-19
C12074 _114_ _176_/a_27_47# 1.25e-20
C12075 _166_/a_161_47# net3 3.74e-21
C12076 VPWR _220_/a_199_47# 4.24e-19
C12077 mask\[0\] _315_/a_1108_47# 6.28e-21
C12078 net4 _335_/a_193_47# 0.00102f
C12079 _023_ _310_/a_27_47# 6.27e-19
C12080 _253_/a_299_297# _074_ 0.0478f
C12081 VPWR _060_ 0.189f
C12082 _192_/a_27_47# _065_ 0.0136f
C12083 net47 _068_ 3.15e-19
C12084 _087_ _092_ 0.0261f
C12085 _089_ _099_ 9.94e-20
C12086 clknet_2_0__leaf_clk _315_/a_761_289# 0.00145f
C12087 _014_ _315_/a_193_47# 0.00248f
C12088 net45 _315_/a_27_47# 0.00178f
C12089 cal_itt\[0\] _065_ 0.0235f
C12090 _249_/a_373_47# _101_ 5.79e-19
C12091 _050_ _028_ 0.182f
C12092 net8 trim_val\[2\] 0.179f
C12093 _318_/a_1270_413# net45 -3.58e-20
C12094 _159_/a_27_47# _220_/a_113_297# 1.62e-21
C12095 _321_/a_27_47# clknet_2_1__leaf_clk 0.19f
C12096 trim_mask\[0\] _332_/a_1108_47# 0.0462f
C12097 _326_/a_1217_47# mask\[7\] 7.28e-19
C12098 _078_ _086_ 0.00284f
C12099 _286_/a_218_374# _122_ 7.33e-19
C12100 trim_mask\[0\] _029_ 0.00237f
C12101 VPWR _178_/a_150_297# 1.12e-19
C12102 _136_ _300_/a_285_47# 0.00637f
C12103 net1 valid 0.0364f
C12104 _314_/a_1108_47# _010_ 1.93e-21
C12105 _041_ _286_/a_439_47# 0.00175f
C12106 net8 net16 0.0137f
C12107 _124_ _338_/a_27_47# 2.26e-20
C12108 _324_/a_1108_47# _020_ 0.00287f
C12109 _006_ _310_/a_193_47# 1.06e-20
C12110 fanout43/a_27_47# _245_/a_27_297# 0.0216f
C12111 _002_ _202_/a_79_21# 0.00349f
C12112 VPWR _020_ 0.13f
C12113 VPWR _327_/a_1462_47# 2.34e-19
C12114 _263_/a_297_47# _092_ 0.0243f
C12115 clknet_2_0__leaf_clk net45 0.853f
C12116 _059_ _237_/a_505_21# 7.37e-21
C12117 _074_ _313_/a_805_47# 1.15e-20
C12118 cal_count\[3\] _278_/a_109_297# 9.2e-19
C12119 _256_/a_109_297# trim_mask\[1\] 0.00191f
C12120 trim_mask\[4\] _279_/a_204_297# 5.72e-20
C12121 net27 net28 0.41f
C12122 _143_/a_68_297# clkbuf_2_1__f_clk/a_110_47# 5.14e-19
C12123 _327_/a_27_47# clknet_2_2__leaf_clk 0.0668f
C12124 _190_/a_465_47# net19 0.00242f
C12125 result[3] result[4] 0.0472f
C12126 _313_/a_193_47# _221_/a_109_297# 6.1e-21
C12127 net44 _068_ 0.0278f
C12128 _319_/a_1283_21# net30 1.19e-19
C12129 _162_/a_27_47# net49 5.55e-21
C12130 _218_/a_113_297# mask\[5\] 9e-21
C12131 state\[2\] _087_ 0.00261f
C12132 net54 _263_/a_79_21# 0.00284f
C12133 trim[2] _056_ 0.00662f
C12134 _274_/a_75_212# rebuffer1/a_75_212# 1.32e-20
C12135 output21/a_27_47# mask\[6\] 0.00634f
C12136 cal_itt\[0\] _194_/a_113_297# 3.46e-19
C12137 _100_ _049_ 0.0119f
C12138 net12 _305_/a_761_289# 7.74e-20
C12139 mask\[5\] _312_/a_27_47# 1.04e-19
C12140 cal_itt\[2\] _202_/a_79_21# 0.00272f
C12141 clknet_2_0__leaf_clk _065_ 0.113f
C12142 en_co_clk net41 3.57e-19
C12143 _081_ _039_ 9.79e-21
C12144 _313_/a_193_47# net29 0.0017f
C12145 _259_/a_27_297# clknet_2_2__leaf_clk 5.1e-19
C12146 cal_itt\[1\] _304_/a_193_47# 1.53e-19
C12147 VPWR _222_/a_199_47# -1.05e-19
C12148 _189_/a_27_47# clk 0.0122f
C12149 output14/a_27_47# output28/a_27_47# 0.00151f
C12150 _269_/a_299_297# _172_/a_150_297# 8.01e-20
C12151 _321_/a_1283_21# _018_ 4.83e-21
C12152 _074_ _041_ 0.0864f
C12153 _294_/a_68_297# VPWR 0.00585f
C12154 trim_mask\[2\] _335_/a_1108_47# 5.98e-21
C12155 _341_/a_1283_21# net46 0.0148f
C12156 net27 _159_/a_27_47# 0.0334f
C12157 mask\[0\] _319_/a_543_47# 0.036f
C12158 VPWR en_co_clk 6.29f
C12159 _080_ mask\[1\] 0.00324f
C12160 trimb[1] net37 0.00242f
C12161 _321_/a_193_47# mask\[6\] 7.54e-20
C12162 _185_/a_68_297# net3 7.88e-22
C12163 _321_/a_543_47# net26 6.88e-20
C12164 _319_/a_27_47# clknet_2_0__leaf_clk 0.62f
C12165 _321_/a_651_413# _042_ 0.00176f
C12166 _307_/a_193_47# _137_/a_150_297# 5.99e-20
C12167 _083_ mask\[4\] 0.284f
C12168 _305_/a_761_289# net44 0.0065f
C12169 cal_count\[0\] net34 1.94e-19
C12170 trim_mask\[2\] rebuffer2/a_75_212# 6.01e-22
C12171 net44 _311_/a_448_47# 5.66e-19
C12172 _134_ _295_/a_113_47# 1.68e-19
C12173 _293_/a_81_21# net16 0.00959f
C12174 _322_/a_1108_47# rebuffer5/a_161_47# 2.12e-19
C12175 state\[2\] _263_/a_297_47# 1.72e-20
C12176 _321_/a_1217_47# clknet_2_1__leaf_clk 8.36e-20
C12177 _104_ _266_/a_68_297# 0.00161f
C12178 net50 _058_ 0.0378f
C12179 _259_/a_109_297# net50 0.00887f
C12180 _259_/a_109_47# trim_mask\[3\] 0.00453f
C12181 _064_ _275_/a_299_297# 1.87e-19
C12182 _323_/a_193_47# _311_/a_1283_21# 1.72e-19
C12183 _323_/a_27_47# _311_/a_1108_47# 5.58e-19
C12184 _340_/a_562_413# _123_ 0.00221f
C12185 _276_/a_59_75# net4 7.64e-22
C12186 clknet_2_1__leaf_clk _313_/a_651_413# 0.00144f
C12187 mask\[7\] _224_/a_199_47# 0.00145f
C12188 _286_/a_439_47# net18 2.47e-19
C12189 VPWR _306_/a_193_47# 0.0353f
C12190 net7 net14 3.57e-21
C12191 _327_/a_1108_47# _265_/a_299_297# 1.68e-20
C12192 _312_/a_193_47# _084_ 2.63e-19
C12193 _097_ net55 1.31e-20
C12194 _326_/a_193_47# net14 0.00884f
C12195 _178_/a_68_297# clknet_2_2__leaf_clk 3.17e-20
C12196 _061_ net34 6.04e-19
C12197 net37 trimb[4] 0.00207f
C12198 _341_/a_1108_47# _300_/a_47_47# 3.89e-19
C12199 _305_/a_543_47# _073_ 4.8e-21
C12200 _110_ _051_ 3.65e-20
C12201 _329_/a_1108_47# rebuffer1/a_75_212# 2.03e-20
C12202 _335_/a_1283_21# net18 0.00776f
C12203 _322_/a_805_47# mask\[2\] 1.81e-19
C12204 net35 _333_/a_1283_21# 1.16e-19
C12205 cal input3/a_75_212# 0.00459f
C12206 net43 output14/a_27_47# 0.0031f
C12207 net15 _245_/a_109_297# 4.09e-19
C12208 net47 _042_ 0.0705f
C12209 net16 _144_/a_27_47# 0.0102f
C12210 _214_/a_113_297# _247_/a_27_297# 5.11e-20
C12211 _182_/a_27_47# _109_ 1.08e-19
C12212 fanout45/a_27_47# _317_/a_1283_21# 0.00344f
C12213 _262_/a_27_47# net55 0.0368f
C12214 VPWR ctlp[3] 0.11f
C12215 _050_ _095_ 0.501f
C12216 net8 _176_/a_27_47# 2.96e-19
C12217 _258_/a_27_297# trim_mask\[1\] 2.65e-19
C12218 _253_/a_299_297# net26 6.75e-19
C12219 _134_ _332_/a_761_289# 2.32e-19
C12220 _024_ trim_mask\[1\] 8.08e-20
C12221 trim[2] _173_/a_27_47# 8.78e-19
C12222 net9 _340_/a_193_47# 0.0212f
C12223 _198_/a_27_47# _062_ 6.55e-20
C12224 _307_/a_27_47# _074_ 0.0166f
C12225 en_co_clk _063_ 0.0175f
C12226 _108_ net18 0.192f
C12227 clk _227_/a_109_93# 0.00819f
C12228 _315_/a_1283_21# _096_ 8.71e-21
C12229 _326_/a_27_47# net28 9.15e-20
C12230 _228_/a_297_47# net41 4.1e-20
C12231 _023_ clknet_2_1__leaf_clk 0.184f
C12232 net43 _306_/a_1283_21# 0.00135f
C12233 VPWR _330_/a_805_47# 2.28e-19
C12234 _339_/a_193_47# _124_ 1.29e-20
C12235 trim_mask\[0\] _171_/a_27_47# 3.71e-19
C12236 _071_ _067_ 0.0156f
C12237 _275_/a_299_297# _057_ 2.45e-19
C12238 _071_ _070_ 1.97e-19
C12239 net12 _250_/a_373_47# 0.00129f
C12240 _216_/a_199_47# mask\[3\] 0.00132f
C12241 _087_ _226_/a_197_47# 3.03e-20
C12242 _304_/a_27_47# _065_ 0.0109f
C12243 cal_itt\[1\] _106_ 8.72e-20
C12244 _337_/a_1270_413# _049_ 1.04e-19
C12245 net12 _042_ 0.00452f
C12246 _317_/a_27_47# _316_/a_27_47# 5.3e-21
C12247 clk _317_/a_193_47# 0.00965f
C12248 _104_ _028_ 1.08e-20
C12249 cal_itt\[1\] _304_/a_1462_47# 4.99e-19
C12250 _103_ clone1/a_27_47# 0.00696f
C12251 VPWR net7 0.214f
C12252 VPWR _235_/a_297_47# -6.55e-19
C12253 fanout44/a_27_47# mask\[1\] 9.97e-21
C12254 VPWR _326_/a_193_47# 0.0221f
C12255 _314_/a_651_413# net14 0.00311f
C12256 _101_ _077_ 0.00277f
C12257 _329_/a_193_47# _031_ 1.39e-19
C12258 VPWR _334_/a_193_47# 0.0342f
C12259 VPWR _228_/a_297_47# -0.00239f
C12260 _164_/a_161_47# en_co_clk 9.44e-19
C12261 net4 _227_/a_109_93# 1.04e-21
C12262 _306_/a_543_47# _101_ 4.44e-21
C12263 _239_/a_474_297# _051_ 0.00233f
C12264 _321_/a_1283_21# _078_ 1.24e-21
C12265 clknet_0_clk net51 1.07e-20
C12266 _307_/a_1108_47# _039_ 0.0336f
C12267 net42 clk 0.0128f
C12268 VPWR _286_/a_76_199# 0.00297f
C12269 _124_ clknet_2_3__leaf_clk 2.19e-19
C12270 _330_/a_27_47# net19 0.0187f
C12271 net4 _317_/a_193_47# 0.0134f
C12272 _321_/a_761_289# clknet_2_0__leaf_clk 1.49e-20
C12273 cal_itt\[0\] clkbuf_0_clk/a_110_47# 0.0265f
C12274 result[0] _039_ 2.93e-19
C12275 state\[1\] _100_ 0.0265f
C12276 _335_/a_27_47# _280_/a_75_212# 2.42e-20
C12277 _078_ _313_/a_27_47# 0.00921f
C12278 net14 _310_/a_543_47# 0.00416f
C12279 _042_ net44 0.0115f
C12280 _233_/a_373_47# net14 7.15e-19
C12281 calibrate _013_ 0.0224f
C12282 _338_/a_1602_47# _123_ 4.3e-20
C12283 _300_/a_129_47# clknet_2_3__leaf_clk 0.00307f
C12284 _181_/a_150_297# _058_ 4.66e-19
C12285 _337_/a_27_47# net45 2.29e-20
C12286 _337_/a_761_289# clknet_2_0__leaf_clk 6.55e-19
C12287 net55 wire42/a_75_212# 0.00638f
C12288 net28 _314_/a_448_47# 0.0037f
C12289 _309_/a_27_47# _310_/a_1108_47# 3.96e-19
C12290 _309_/a_193_47# _310_/a_1283_21# 5.38e-20
C12291 trim_mask\[3\] _330_/a_27_47# 5.23e-20
C12292 _326_/a_1283_21# net43 1.67e-19
C12293 VPWR _306_/a_1462_47# 1.48e-19
C12294 _323_/a_543_47# clknet_2_1__leaf_clk 1.49e-19
C12295 cal_itt\[1\] trim_mask\[0\] 7.2e-20
C12296 _248_/a_109_47# mask\[4\] 0.00184f
C12297 net9 _136_ 0.0501f
C12298 _099_ _092_ 0.266f
C12299 VPWR _314_/a_651_413# 0.00121f
C12300 _002_ _041_ 3.63e-20
C12301 clk _054_ 0.00996f
C12302 clk _318_/a_1283_21# 0.031f
C12303 _041_ net26 5.16e-20
C12304 _337_/a_27_47# _065_ 0.0302f
C12305 _233_/a_109_297# valid 0.00145f
C12306 clk net30 1.03f
C12307 net15 _016_ 0.0382f
C12308 net12 _318_/a_543_47# 7.82e-19
C12309 _290_/a_27_413# output37/a_27_47# 0.011f
C12310 _069_ _065_ 0.0747f
C12311 _326_/a_193_47# net52 0.00214f
C12312 _336_/a_27_47# _336_/a_448_47# -0.00346f
C12313 trim_mask\[2\] _112_ 6.44e-20
C12314 trim_mask\[2\] _272_/a_299_297# 5.7e-20
C12315 net9 _340_/a_796_47# 5.14e-19
C12316 net14 _039_ 0.00234f
C12317 _253_/a_384_47# _078_ 5.45e-19
C12318 _319_/a_1283_21# _319_/a_1108_47# -2.84e-32
C12319 _319_/a_27_47# _319_/a_639_47# -0.0015f
C12320 output35/a_27_47# trim_val\[0\] 6.59e-20
C12321 _169_/a_215_311# _092_ 1.18e-21
C12322 _325_/a_193_47# mask\[2\] 9.95e-20
C12323 _307_/a_805_47# calibrate 3.52e-21
C12324 _209_/a_27_47# rebuffer5/a_161_47# 0.0197f
C12325 _168_/a_27_413# clk 0.00939f
C12326 _119_ net46 0.0655f
C12327 VPWR _310_/a_543_47# 7.17e-19
C12328 cal_itt\[0\] _038_ 6.38e-20
C12329 VPWR _233_/a_373_47# -2.5e-19
C12330 clknet_2_2__leaf_clk net40 0.0226f
C12331 trim_mask\[4\] _278_/a_27_47# 2.53e-20
C12332 _340_/a_652_21# cal_count\[2\] 1.56e-19
C12333 _339_/a_1140_413# cal_count\[0\] 1.36e-19
C12334 net4 net30 0.0619f
C12335 _327_/a_27_47# _327_/a_448_47# -0.00373f
C12336 _243_/a_109_47# net55 8.55e-19
C12337 state\[0\] _050_ 5.44e-19
C12338 cal_itt\[2\] _041_ 5.23e-20
C12339 _304_/a_1217_47# _065_ 2.55e-19
C12340 clk _317_/a_1462_47# 2.24e-19
C12341 cal_itt\[0\] _338_/a_476_47# 3.8e-19
C12342 input4/a_27_47# output6/a_27_47# 1.74e-20
C12343 clknet_2_2__leaf_clk _330_/a_639_47# 0.00497f
C12344 trim_mask\[4\] _330_/a_1283_21# 4.53e-19
C12345 trim_val\[2\] net34 0.0981f
C12346 VPWR _326_/a_1462_47# 0.00178f
C12347 _292_/a_78_199# cal_count\[0\] 1.96e-20
C12348 _036_ _286_/a_76_199# 8.26e-20
C12349 _107_ _076_ 2.89e-19
C12350 _267_/a_145_75# clknet_2_2__leaf_clk 3.94e-19
C12351 _168_/a_27_413# net4 3.44e-21
C12352 _019_ net15 -1.01e-36
C12353 _104_ _279_/a_314_297# 6.76e-19
C12354 _327_/a_1108_47# _058_ 0.0142f
C12355 output25/a_27_47# _074_ 4.25e-19
C12356 clk _072_ 0.207f
C12357 _334_/a_27_47# clknet_2_2__leaf_clk 0.0207f
C12358 _097_ _316_/a_543_47# 3.7e-19
C12359 net16 net34 0.0142f
C12360 net12 cal_itt\[3\] 0.012f
C12361 state\[2\] _099_ 1.26e-19
C12362 VPWR cal_count\[0\] 0.336f
C12363 _094_ _090_ 2.67e-20
C12364 net43 _310_/a_448_47# 3e-19
C12365 _311_/a_543_47# net53 0.00637f
C12366 _303_/a_639_47# _068_ 2.23e-19
C12367 VPWR _039_ 0.456f
C12368 _273_/a_59_75# _114_ 0.0371f
C12369 _115_ _272_/a_299_297# 5.06e-19
C12370 _115_ _112_ 0.00388f
C12371 result[0] result[1] 0.0489f
C12372 net30 _073_ 0.348f
C12373 _282_/a_68_297# clknet_2_0__leaf_clk 0.0127f
C12374 _090_ _088_ 1.46e-20
C12375 VPWR _335_/a_805_47# 3.65e-19
C12376 _197_/a_113_297# _067_ 0.00155f
C12377 VPWR _305_/a_193_47# -0.0425f
C12378 _322_/a_193_47# _247_/a_27_297# 1.58e-20
C12379 net2 _198_/a_27_47# 3.03e-20
C12380 _275_/a_81_21# net46 1.21e-19
C12381 trim_mask\[3\] _330_/a_1217_47# 1.1e-19
C12382 _051_ net45 0.00193f
C12383 VPWR _311_/a_1108_47# -0.00144f
C12384 state\[2\] _169_/a_215_311# 0.0157f
C12385 _015_ _060_ 0.0675f
C12386 _064_ _092_ 0.00523f
C12387 _050_ _226_/a_27_47# 6.6e-19
C12388 _101_ _310_/a_1108_47# 1.33e-21
C12389 net16 _299_/a_298_297# 0.00289f
C12390 VPWR _061_ 0.0542f
C12391 net44 cal_itt\[3\] 0.0603f
C12392 trim_val\[0\] net40 3.63e-20
C12393 mask\[7\] _086_ 0.00401f
C12394 ctln[4] trim_mask\[3\] 1.69e-19
C12395 _194_/a_199_47# _067_ 4.04e-19
C12396 VPWR _332_/a_639_47# 0.00379f
C12397 _052_ _242_/a_79_21# 0.0196f
C12398 _126_ _122_ 1.19e-19
C12399 _304_/a_193_47# _302_/a_27_297# 3.45e-21
C12400 _304_/a_27_47# _302_/a_109_297# 4.56e-21
C12401 _103_ _051_ 0.0432f
C12402 net9 _301_/a_129_47# 9.57e-21
C12403 net55 _206_/a_27_93# 1.27e-19
C12404 _012_ valid 0.0086f
C12405 _337_/a_1217_47# _065_ 9.91e-20
C12406 net13 _232_/a_32_297# 0.00856f
C12407 _202_/a_79_21# _070_ 0.00627f
C12408 net9 _338_/a_1140_413# 1.04e-19
C12409 net43 _247_/a_27_297# 4.34e-21
C12410 net23 _039_ 1.96e-19
C12411 _051_ _065_ 8.6e-23
C12412 net9 _341_/a_761_289# 7.52e-19
C12413 net3 _062_ 0.00358f
C12414 _336_/a_27_47# _033_ 0.0355f
C12415 _336_/a_543_47# _106_ 7.17e-19
C12416 _335_/a_27_47# net19 0.00104f
C12417 net43 net2 3.18e-20
C12418 _339_/a_381_47# _123_ 0.0146f
C12419 _322_/a_1108_47# net51 3.81e-20
C12420 _053_ _092_ 0.0183f
C12421 mask\[3\] mask\[2\] 0.0187f
C12422 _200_/a_80_21# clknet_2_3__leaf_clk 0.00128f
C12423 net5 _047_ 4.5e-19
C12424 result[1] net14 5.96e-20
C12425 _289_/a_68_297# _129_ 0.00941f
C12426 _126_ _299_/a_27_413# 4.82e-20
C12427 net43 _305_/a_1283_21# 0.00716f
C12428 _003_ cal_itt\[3\] 2.56e-19
C12429 _073_ _072_ 3.27e-19
C12430 _058_ _193_/a_109_297# 2.5e-19
C12431 _321_/a_27_47# _321_/a_761_289# -0.0166f
C12432 trim_mask\[3\] _335_/a_27_47# 0.002f
C12433 trim_val\[3\] _335_/a_193_47# 6.48e-19
C12434 output28/a_27_47# net29 2.96e-19
C12435 _094_ _048_ 0.00253f
C12436 _008_ _311_/a_543_47# 4.27e-19
C12437 _286_/a_505_21# _001_ 1.03e-19
C12438 _338_/a_193_47# _065_ 1.8e-20
C12439 trim_mask\[1\] cal_count\[3\] 2.64e-20
C12440 _014_ _316_/a_1108_47# 0.00182f
C12441 clknet_2_0__leaf_clk _316_/a_448_47# 9.35e-19
C12442 net45 _316_/a_1283_21# -0.00315f
C12443 _337_/a_543_47# net55 0.00186f
C12444 _169_/a_301_53# state\[0\] 1.53e-19
C12445 cal_itt\[0\] _341_/a_448_47# 7.48e-21
C12446 net27 _044_ 0.00603f
C12447 _048_ _088_ 0.217f
C12448 clkbuf_0_clk/a_110_47# _304_/a_27_47# 8.33e-21
C12449 _320_/a_27_47# _078_ 3.44e-19
C12450 _305_/a_193_47# _063_ 7.72e-20
C12451 _101_ _311_/a_651_413# 2.69e-21
C12452 _036_ cal_count\[0\] 0.083f
C12453 _307_/a_543_47# net30 1.21e-19
C12454 net9 _339_/a_27_47# 0.0159f
C12455 _309_/a_1108_47# clknet_2_1__leaf_clk 3.88e-21
C12456 net2 _297_/a_129_47# 5.79e-19
C12457 _257_/a_27_297# trim_mask\[1\] 0.0961f
C12458 mask\[1\] _076_ 2.4e-19
C12459 result[2] _006_ 8.61e-19
C12460 net16 _133_ 0.0261f
C12461 _034_ en_co_clk 5.03e-19
C12462 _271_/a_75_212# clknet_2_2__leaf_clk 0.0696f
C12463 _074_ _312_/a_543_47# 3.22e-20
C12464 clkbuf_2_1__f_clk/a_110_47# _101_ 0.0272f
C12465 trim_mask\[4\] _088_ 1.03e-19
C12466 _250_/a_27_297# net53 0.0241f
C12467 trim_mask\[0\] _336_/a_543_47# 4.83e-20
C12468 _173_/a_27_47# net32 0.0217f
C12469 net47 _149_/a_150_297# 2.47e-19
C12470 _333_/a_27_47# rebuffer2/a_75_212# 4.72e-20
C12471 VPWR result[1] 0.188f
C12472 _175_/a_68_297# _108_ 0.0279f
C12473 _326_/a_193_47# _216_/a_113_297# 7.22e-21
C12474 _333_/a_193_47# _108_ 0.00776f
C12475 mask\[5\] _084_ 0.0617f
C12476 _068_ net19 0.276f
C12477 _324_/a_1283_21# _042_ 2.73e-20
C12478 result[6] clknet_2_1__leaf_clk 0.0373f
C12479 calibrate _242_/a_79_21# 0.00237f
C12480 _307_/a_193_47# _078_ 0.0115f
C12481 _307_/a_761_289# mask\[0\] 7.07e-20
C12482 _307_/a_543_47# net22 0.015f
C12483 _259_/a_27_297# _330_/a_1283_21# 0.00828f
C12484 VPWR _305_/a_1462_47# 3.12e-19
C12485 VPWR _251_/a_27_297# 0.0704f
C12486 _328_/a_1283_21# _329_/a_1283_21# 1.06e-19
C12487 VPWR _250_/a_109_47# -3.87e-19
C12488 _015_ en_co_clk 6.27e-19
C12489 _265_/a_81_21# _108_ 0.00859f
C12490 _265_/a_81_21# _332_/a_543_47# 0.00114f
C12491 state\[2\] _053_ 0.129f
C12492 _329_/a_651_413# net9 0.00203f
C12493 output34/a_27_47# _334_/a_1283_21# 9e-19
C12494 net34 _176_/a_27_47# 0.0156f
C12495 clknet_0_clk _262_/a_109_297# 0.00374f
C12496 _335_/a_1283_21# trim_mask\[4\] 7.62e-19
C12497 output22/a_27_47# clknet_2_0__leaf_clk 0.0311f
C12498 net43 net29 0.0608f
C12499 _302_/a_109_47# _067_ 1.47e-19
C12500 _048_ _108_ 0.00102f
C12501 _322_/a_543_47# _042_ 3.29e-20
C12502 _110_ _119_ 0.00786f
C12503 _235_/a_79_21# _095_ 0.00715f
C12504 net15 _095_ 0.0835f
C12505 _246_/a_27_297# _017_ 0.00919f
C12506 _304_/a_27_47# _038_ 1.35e-20
C12507 _277_/a_75_212# net18 8.68e-19
C12508 _138_/a_27_47# net30 9.28e-20
C12509 _333_/a_639_47# net46 0.00232f
C12510 _237_/a_439_47# _049_ 7.78e-20
C12511 _255_/a_27_47# clkbuf_2_3__f_clk/a_110_47# 1.92e-20
C12512 _083_ _311_/a_1108_47# 1.65e-20
C12513 _001_ _068_ 1.8e-20
C12514 output25/a_27_47# net26 6.71e-20
C12515 trim_mask\[4\] _108_ 0.183f
C12516 result[1] net23 0.00306f
C12517 net20 _009_ 0.0217f
C12518 _304_/a_448_47# net47 -2.34e-19
C12519 _062_ _190_/a_465_47# 0.00215f
C12520 _200_/a_209_47# VPWR -7.92e-19
C12521 _071_ clknet_2_3__leaf_clk 7.99e-20
C12522 _009_ net53 1.32e-20
C12523 _030_ _333_/a_761_289# 7.67e-19
C12524 _113_ _333_/a_543_47# 3.51e-20
C12525 net43 _251_/a_373_47# 6.22e-20
C12526 ctln[7] _318_/a_543_47# 1.28e-19
C12527 net13 _318_/a_1108_47# 0.00312f
C12528 _230_/a_59_75# net4 0.012f
C12529 _218_/a_113_297# clknet_2_1__leaf_clk 5.24e-19
C12530 _050_ _052_ 0.349f
C12531 _340_/a_27_47# _340_/a_562_413# -0.0012f
C12532 _340_/a_193_47# _340_/a_381_47# -5.68e-19
C12533 _319_/a_193_47# _121_ 3.72e-20
C12534 _040_ _049_ 2.28e-19
C12535 net50 _335_/a_805_47# 2.13e-19
C12536 clknet_2_1__leaf_clk _312_/a_27_47# 0.0695f
C12537 _308_/a_543_47# net24 7.21e-21
C12538 _049_ net41 0.0018f
C12539 net44 _319_/a_1283_21# 1.61e-19
C12540 net8 _273_/a_59_75# 7.89e-20
C12541 _318_/a_761_289# net41 2.4e-20
C12542 _308_/a_1283_21# clknet_2_0__leaf_clk 1.65e-19
C12543 net22 _138_/a_27_47# 0.0015f
C12544 _262_/a_27_47# clknet_2_3__leaf_clk 1.87e-19
C12545 _008_ _250_/a_27_297# 2.07e-21
C12546 _299_/a_215_297# _131_ 0.0538f
C12547 _281_/a_253_47# en_co_clk 5.79e-19
C12548 _281_/a_337_297# _120_ 8.29e-19
C12549 _059_ _060_ 0.596f
C12550 _338_/a_796_47# _065_ 1.61e-20
C12551 clknet_2_0__leaf_clk _013_ 0.0347f
C12552 VPWR trim_val\[2\] 0.349f
C12553 _292_/a_78_199# net16 5.04e-19
C12554 _323_/a_27_47# _149_/a_68_297# 7.54e-19
C12555 _337_/a_27_47# _282_/a_68_297# 6.09e-19
C12556 _251_/a_27_297# net52 0.0839f
C12557 net5 _301_/a_47_47# 7.27e-20
C12558 _306_/a_1270_413# _092_ 5.17e-21
C12559 _313_/a_193_47# _313_/a_1283_21# -9.9e-20
C12560 cal_itt\[0\] _303_/a_1283_21# 0.00609f
C12561 net27 mask\[2\] 4.53e-21
C12562 net31 output34/a_27_47# 1.78e-19
C12563 net9 _339_/a_586_47# 2.06e-19
C12564 _320_/a_639_47# clknet_2_0__leaf_clk 3.68e-19
C12565 VPWR _049_ 0.988f
C12566 trimb[0] net34 0.0659f
C12567 VPWR _318_/a_761_289# 0.0123f
C12568 _325_/a_193_47# _074_ 9.03e-20
C12569 net13 mask\[0\] 0.00197f
C12570 trim_mask\[0\] _302_/a_27_297# 4.91e-21
C12571 _110_ _275_/a_81_21# 0.0625f
C12572 _276_/a_59_75# trim_val\[3\] 2.68e-19
C12573 trim_mask\[2\] net33 0.00626f
C12574 VPWR net16 1.84f
C12575 _232_/a_220_297# _090_ 0.00378f
C12576 _035_ _338_/a_27_47# 0.0112f
C12577 _289_/a_68_297# _297_/a_47_47# 4.35e-19
C12578 net4 _066_ 2.22e-19
C12579 trim_mask\[2\] _336_/a_761_289# 1.41e-21
C12580 _078_ rebuffer6/a_27_47# 9.27e-20
C12581 net51 _209_/a_27_47# 0.00296f
C12582 _140_/a_68_297# net45 3.35e-20
C12583 trim_mask\[0\] _106_ 0.152f
C12584 trim[3] net46 1.66e-19
C12585 _324_/a_448_47# _021_ 0.00226f
C12586 _324_/a_193_47# _078_ 1.08e-20
C12587 _333_/a_1462_47# _108_ 3.59e-19
C12588 _104_ _330_/a_1108_47# 5.9e-20
C12589 _328_/a_761_289# VPWR 0.0104f
C12590 _330_/a_27_47# _330_/a_761_289# -0.0166f
C12591 ctln[5] _330_/a_448_47# 4.12e-20
C12592 _200_/a_209_47# _063_ 0.00187f
C12593 _307_/a_1270_413# net45 -2.06e-19
C12594 _168_/a_207_413# _331_/a_193_47# 2.79e-21
C12595 _308_/a_193_47# _319_/a_193_47# 0.00148f
C12596 _302_/a_373_47# _136_ 3.16e-19
C12597 _029_ _109_ 7.06e-19
C12598 _227_/a_209_311# _260_/a_93_21# 4.03e-19
C12599 VPWR _317_/a_805_47# 5.66e-20
C12600 output35/a_27_47# trim[4] 0.00977f
C12601 _307_/a_543_47# _079_ 4.49e-19
C12602 _307_/a_193_47# _004_ 0.00546f
C12603 _100_ _240_/a_109_297# 6.37e-19
C12604 _315_/a_1108_47# net14 0.00637f
C12605 mask\[7\] _313_/a_27_47# 6.7e-19
C12606 _304_/a_193_47# _298_/a_78_199# 4.02e-20
C12607 _060_ _075_ 0.0648f
C12608 _322_/a_27_47# _078_ 0.0041f
C12609 clknet_2_3__leaf_clk cal_count\[2\] 3.1e-20
C12610 _319_/a_761_289# clknet_0_clk 0.00127f
C12611 _050_ calibrate 0.501f
C12612 output38/a_27_47# trimb[3] 9.86e-19
C12613 trimb[2] output39/a_27_47# 0.00275f
C12614 _041_ _067_ 2.26e-20
C12615 _304_/a_651_413# _122_ 0.00442f
C12616 _041_ _070_ 6.58e-20
C12617 _115_ net33 1.51e-21
C12618 _336_/a_193_47# net18 8.89e-21
C12619 mask\[6\] _312_/a_193_47# 3.48e-20
C12620 _051_ clkbuf_0_clk/a_110_47# 4.12e-20
C12621 _112_ _333_/a_27_47# 0.0184f
C12622 trim_mask\[1\] _333_/a_761_289# 7.01e-19
C12623 net49 _333_/a_193_47# 0.0129f
C12624 trim_val\[1\] _333_/a_543_47# 0.00171f
C12625 net52 _049_ 2.01e-19
C12626 _063_ _049_ 9.1e-20
C12627 _117_ clknet_2_2__leaf_clk 8.95e-22
C12628 _101_ net30 4.32e-20
C12629 state\[0\] net15 0.0042f
C12630 _042_ net19 0.0106f
C12631 _037_ _304_/a_651_413# 2.26e-19
C12632 net54 _094_ 0.00268f
C12633 _315_/a_543_47# valid 0.00124f
C12634 net43 mask\[0\] 0.6f
C12635 _005_ _078_ 2.11e-19
C12636 _127_ _297_/a_285_47# 7.44e-21
C12637 _259_/a_27_297# _335_/a_1283_21# 3.08e-19
C12638 _327_/a_27_47# _108_ 0.03f
C12639 _105_ _261_/a_113_47# 2.27e-19
C12640 _134_ clkc 2.48e-19
C12641 net54 _088_ 6.12e-21
C12642 VPWR _262_/a_193_297# 0.00304f
C12643 _059_ en_co_clk 0.091f
C12644 _232_/a_32_297# net3 0.00234f
C12645 _219_/a_109_297# _078_ 0.00526f
C12646 _308_/a_448_47# _004_ 1.79e-20
C12647 _007_ _074_ 0.0698f
C12648 _253_/a_299_297# _102_ 7.3e-19
C12649 _253_/a_384_47# mask\[7\] 3.46e-19
C12650 _253_/a_81_21# _023_ 0.00209f
C12651 net38 net33 0.0369f
C12652 _309_/a_639_47# _078_ 9.62e-19
C12653 _117_ net11 1.72e-19
C12654 _323_/a_543_47# _043_ 1.57e-20
C12655 _187_/a_297_47# _058_ 1.5e-19
C12656 _090_ _192_/a_174_21# 4.94e-20
C12657 VPWR _315_/a_1108_47# 0.0124f
C12658 _309_/a_448_47# net24 0.0164f
C12659 _337_/a_448_47# net44 3.99e-20
C12660 net28 _086_ 0.106f
C12661 _074_ _249_/a_27_297# 4.66e-19
C12662 net35 _332_/a_27_47# 7.94e-19
C12663 _058_ _332_/a_761_289# 0.00357f
C12664 clkbuf_2_2__f_clk/a_110_47# _264_/a_27_297# 5.39e-21
C12665 _278_/a_27_47# net40 2.08e-19
C12666 _024_ _136_ 7.49e-19
C12667 _239_/a_694_21# _048_ 0.052f
C12668 _074_ mask\[3\] 0.116f
C12669 _200_/a_303_47# net19 0.00109f
C12670 net27 _314_/a_193_47# 8.02e-20
C12671 _327_/a_1270_413# net46 1.29e-19
C12672 _035_ _338_/a_586_47# 3.33e-19
C12673 _126_ _297_/a_285_47# 2.58e-20
C12674 _260_/a_346_47# _049_ 3.59e-20
C12675 _047_ _055_ 3.3e-20
C12676 _048_ _227_/a_368_53# 3.75e-19
C12677 state\[1\] net41 0.00658f
C12678 VPWR _201_/a_113_47# -4.43e-20
C12679 clk _316_/a_27_47# 2.74e-19
C12680 trim[4] net40 0.00188f
C12681 net47 net4 0.0212f
C12682 net12 clk 0.0267f
C12683 clknet_0_clk _206_/a_206_47# 4.75e-19
C12684 _064_ net46 0.0173f
C12685 net12 clone7/a_27_47# 1.4e-20
C12686 VPWR _176_/a_27_47# 0.086f
C12687 _048_ _317_/a_1283_21# 1.69e-19
C12688 output23/a_27_47# _007_ 4.13e-20
C12689 _093_ _092_ 1.08e-19
C12690 _194_/a_199_47# clknet_2_3__leaf_clk 5.14e-19
C12691 _200_/a_303_47# _107_ 8.43e-20
C12692 _168_/a_207_413# _260_/a_93_21# 0.016f
C12693 en_co_clk _075_ 0.17f
C12694 VPWR state\[1\] 0.17f
C12695 net10 net9 2.17e-19
C12696 _328_/a_1108_47# _025_ 7.13e-20
C12697 _328_/a_193_47# clknet_2_2__leaf_clk 0.595f
C12698 _322_/a_1217_47# _078_ 1.61e-19
C12699 _304_/a_543_47# clknet_2_3__leaf_clk 0.00312f
C12700 _030_ _058_ 0.00101f
C12701 _082_ _247_/a_27_297# 1.82e-20
C12702 _104_ _052_ 0.434f
C12703 _340_/a_1182_261# _298_/a_78_199# 0.00134f
C12704 _262_/a_193_297# _063_ 0.0256f
C12705 _078_ net21 0.427f
C12706 net9 clknet_2_2__leaf_clk 0.185f
C12707 _074_ _220_/a_113_297# 3.15e-19
C12708 net12 net4 0.00967f
C12709 net45 _331_/a_651_413# 0.00133f
C12710 _326_/a_1283_21# result[5] 1.47e-19
C12711 _035_ _339_/a_193_47# 7.63e-21
C12712 _257_/a_27_297# _336_/a_27_47# 6.17e-21
C12713 net47 _122_ 0.1f
C12714 clk net44 0.00764f
C12715 _067_ net18 0.0225f
C12716 _237_/a_505_21# _096_ 0.0498f
C12717 _048_ _192_/a_174_21# 0.0324f
C12718 _053_ net46 6.57e-19
C12719 cal_itt\[2\] _048_ 2.04e-20
C12720 _325_/a_193_47# net26 4.29e-20
C12721 mask\[3\] _146_/a_150_297# 2.27e-19
C12722 _325_/a_1108_47# _042_ 1.08e-19
C12723 _340_/a_1140_413# _122_ 2.73e-19
C12724 _041_ _338_/a_27_47# 4.85e-19
C12725 _337_/a_1283_21# clknet_0_clk 2.34e-19
C12726 net47 _338_/a_381_47# 0.0215f
C12727 _338_/a_193_47# _338_/a_476_47# -0.0183f
C12728 _059_ _235_/a_297_47# 1.17e-19
C12729 en_co_clk _195_/a_505_21# 0.0307f
C12730 _037_ net47 0.00229f
C12731 net13 _100_ 0.00763f
C12732 _325_/a_639_47# clknet_2_1__leaf_clk 3.39e-19
C12733 _059_ _228_/a_297_47# 8.65e-21
C12734 _186_/a_109_297# _088_ 9.11e-21
C12735 _104_ _335_/a_1108_47# 7.7e-20
C12736 _327_/a_1217_47# _108_ 3.22e-20
C12737 _326_/a_761_289# output14/a_27_47# 2.73e-21
C12738 _110_ _279_/a_206_47# 0.00264f
C12739 _057_ net46 1.95e-19
C12740 _327_/a_805_47# _111_ 1.11e-19
C12741 net16 _333_/a_448_47# 0.00323f
C12742 _340_/a_652_21# _129_ 2.33e-21
C12743 clknet_2_1__leaf_clk _158_/a_68_297# 0.00905f
C12744 _005_ _004_ 0.00243f
C12745 _239_/a_27_297# _050_ 0.0164f
C12746 _035_ clknet_2_3__leaf_clk 0.107f
C12747 result[4] _074_ 2.42e-19
C12748 clk _003_ 2.86e-19
C12749 mask\[4\] _311_/a_639_47# 0.00428f
C12750 _042_ _248_/a_109_297# 3.94e-19
C12751 net19 cal_itt\[3\] 4.96e-20
C12752 net12 _073_ 0.00478f
C12753 VPWR _319_/a_543_47# 0.0273f
C12754 _313_/a_805_47# _010_ 2.14e-19
C12755 VPWR _149_/a_68_297# 0.0289f
C12756 _120_ _137_/a_68_297# 2.11e-20
C12757 _033_ clknet_0_clk 0.00723f
C12758 VPWR trimb[0] 0.252f
C12759 calibrate net1 0.00394f
C12760 _042_ mask\[1\] 0.00296f
C12761 _326_/a_27_47# _314_/a_193_47# 3.41e-19
C12762 _326_/a_193_47# _314_/a_27_47# 7.79e-19
C12763 _327_/a_193_47# trim_mask\[1\] 9.96e-21
C12764 net17 _041_ 1.18e-20
C12765 _303_/a_193_47# _035_ 1.09e-21
C12766 _187_/a_297_47# en_co_clk 6.97e-19
C12767 _074_ fanout43/a_27_47# 1.42e-19
C12768 _104_ calibrate 0.0487f
C12769 _049_ _279_/a_396_47# 1.43e-19
C12770 net44 _073_ 6.49e-20
C12771 _136_ _298_/a_215_47# 0.00109f
C12772 _081_ _214_/a_113_297# 3.44e-19
C12773 _302_/a_109_47# clknet_2_3__leaf_clk 0.00176f
C12774 _136_ clkbuf_2_3__f_clk/a_110_47# 8.86e-19
C12775 _330_/a_651_413# _027_ 8.49e-19
C12776 _330_/a_448_47# net46 9.44e-22
C12777 ctlp[0] _314_/a_761_289# 9.95e-19
C12778 _164_/a_161_47# state\[1\] 2.13e-19
C12779 net27 _074_ 0.119f
C12780 cal_count\[1\] _131_ 1.02e-20
C12781 _244_/a_27_297# rebuffer5/a_161_47# 8.58e-19
C12782 net43 _319_/a_448_47# 3.2e-20
C12783 _074_ _222_/a_113_297# 1.18e-19
C12784 VPWR _202_/a_297_47# 0.00149f
C12785 _259_/a_109_297# trim_mask\[1\] 1.38e-20
C12786 _199_/a_193_297# _065_ 0.00156f
C12787 _058_ trim_mask\[1\] 0.00544f
C12788 output24/a_27_47# _080_ 8.56e-20
C12789 VPWR _336_/a_651_413# 0.00146f
C12790 _050_ _192_/a_27_47# 8.37e-19
C12791 _328_/a_1462_47# clknet_2_2__leaf_clk 2.16e-19
C12792 _303_/a_1283_21# _069_ 4.45e-19
C12793 VPWR _304_/a_1108_47# 0.02f
C12794 _136_ _134_ 0.00441f
C12795 _007_ net26 0.00175f
C12796 _000_ fanout47/a_27_47# 1.13e-19
C12797 _340_/a_193_47# cal_count\[3\] 1.07e-20
C12798 _107_ _262_/a_205_47# 1.29e-19
C12799 _341_/a_1283_21# _038_ 1.39e-19
C12800 _341_/a_1270_413# _136_ 8.32e-20
C12801 _235_/a_382_297# _094_ 0.0014f
C12802 _249_/a_27_297# net26 8.35e-19
C12803 net51 _208_/a_505_21# 0.144f
C12804 clknet_2_1__leaf_clk _246_/a_27_297# 0.00409f
C12805 _325_/a_1108_47# _022_ 1.61e-19
C12806 _325_/a_805_47# mask\[6\] 0.00211f
C12807 _319_/a_1108_47# _101_ 7.56e-20
C12808 _319_/a_543_47# net52 6.98e-19
C12809 _319_/a_193_47# _016_ 0.0715f
C12810 _341_/a_27_47# _122_ 5.3e-19
C12811 _284_/a_150_297# net18 4.94e-19
C12812 _073_ _003_ 0.00156f
C12813 mask\[3\] net26 0.00358f
C12814 _325_/a_761_289# _078_ 1.14e-21
C12815 _241_/a_297_47# net30 7.26e-20
C12816 _306_/a_27_47# _244_/a_27_297# 0.0129f
C12817 net54 _232_/a_220_297# 0.00188f
C12818 _334_/a_27_47# _334_/a_448_47# -0.00752f
C12819 _303_/a_1108_47# _067_ 5.17e-21
C12820 _338_/a_27_47# net18 0.016f
C12821 _303_/a_1108_47# _070_ 2.47e-19
C12822 _239_/a_277_297# _092_ 0.0588f
C12823 _320_/a_761_289# net44 -0.0067f
C12824 _122_ _299_/a_215_297# 1.87e-19
C12825 mask\[6\] _158_/a_150_297# 1.07e-19
C12826 output23/a_27_47# fanout43/a_27_47# 1.78e-20
C12827 _228_/a_382_297# _088_ 0.00112f
C12828 _228_/a_79_21# _052_ 0.00929f
C12829 cal_itt\[2\] _190_/a_27_47# 0.0397f
C12830 net13 _337_/a_1270_413# 6.96e-20
C12831 net13 _313_/a_1283_21# 4.31e-19
C12832 _185_/a_150_297# _049_ 3.24e-20
C12833 _332_/a_543_47# net40 7.76e-19
C12834 _108_ net40 1.01f
C12835 net28 _313_/a_27_47# 0.209f
C12836 _161_/a_68_297# net46 0.00116f
C12837 _167_/a_161_47# net41 1.11e-19
C12838 VPWR _256_/a_109_47# -9.67e-19
C12839 VPWR _321_/a_1108_47# 0.0172f
C12840 _034_ _049_ 0.0137f
C12841 _323_/a_639_47# net44 4.2e-19
C12842 _110_ _064_ 0.00401f
C12843 clone1/a_27_47# _242_/a_79_21# 7.45e-19
C12844 trim[4] _332_/a_1270_413# 9.46e-21
C12845 _041_ _339_/a_193_47# 0.275f
C12846 _074_ sample 0.0136f
C12847 _333_/a_27_47# net33 2.82e-20
C12848 net47 _339_/a_562_413# 2.38e-19
C12849 VPWR _337_/a_1108_47# 0.00156f
C12850 VPWR _313_/a_193_47# 0.0267f
C12851 _267_/a_145_75# _108_ 1.73e-19
C12852 _304_/a_1108_47# _063_ 0.00103f
C12853 _323_/a_193_47# _323_/a_651_413# -0.00701f
C12854 _111_ _267_/a_59_75# 2.9e-19
C12855 VPWR _167_/a_161_47# 0.0862f
C12856 _050_ clknet_2_0__leaf_clk 0.115f
C12857 _334_/a_1283_21# rebuffer1/a_75_212# 6.81e-19
C12858 net17 net18 0.0821f
C12859 clknet_2_1__leaf_clk _084_ 0.277f
C12860 _068_ _062_ 0.0311f
C12861 _097_ _095_ 9.72e-19
C12862 fanout44/a_27_47# mask\[0\] 4.45e-19
C12863 _192_/a_505_280# _092_ 5.22e-19
C12864 _192_/a_548_47# _095_ 1.35e-20
C12865 net8 _333_/a_543_47# 9.56e-21
C12866 _159_/a_27_47# _313_/a_27_47# 3.54e-20
C12867 net2 _076_ 0.353f
C12868 _136_ cal_count\[3\] 0.193f
C12869 cal_itt\[1\] _092_ 0.00235f
C12870 _090_ net55 0.339f
C12871 _015_ _318_/a_761_289# 6.55e-19
C12872 net30 trim_val\[4\] 6.05e-20
C12873 _027_ net46 0.282f
C12874 _149_/a_150_297# net19 4.36e-19
C12875 _292_/a_215_47# _340_/a_1032_413# 8.4e-19
C12876 _306_/a_761_289# net2 3.19e-21
C12877 _284_/a_68_297# cal_count\[3\] 2.16e-19
C12878 _110_ _053_ 4.68e-19
C12879 calibrate net15 0.00828f
C12880 _235_/a_79_21# calibrate 1.35e-20
C12881 _306_/a_1283_21# _305_/a_761_289# 0.00118f
C12882 _306_/a_1108_47# _305_/a_193_47# 2.86e-19
C12883 _326_/a_543_47# _310_/a_1108_47# 1.16e-20
C12884 _326_/a_1283_21# _310_/a_1283_21# 1.51e-20
C12885 _326_/a_651_413# _310_/a_193_47# 2.21e-20
C12886 _320_/a_27_47# clknet_0_clk 3.01e-19
C12887 ctln[7] clk 1.18e-20
C12888 net43 _321_/a_1270_413# -2.06e-19
C12889 _326_/a_27_47# _074_ 0.019f
C12890 _041_ clknet_2_3__leaf_clk 0.011f
C12891 _338_/a_1182_261# clknet_2_3__leaf_clk 0.0623f
C12892 result[4] net26 0.00273f
C12893 calibrate _228_/a_79_21# 0.0432f
C12894 clknet_2_1__leaf_clk _208_/a_535_374# 3.1e-19
C12895 net54 _192_/a_174_21# 6.74e-19
C12896 VPWR _340_/a_562_413# -7.6e-19
C12897 _104_ _170_/a_384_47# 3.55e-19
C12898 net43 _313_/a_1283_21# -0.0079f
C12899 mask\[6\] mask\[5\] 0.017f
C12900 _195_/a_76_199# _068_ 6.49e-19
C12901 _329_/a_1283_21# _274_/a_75_212# 0.0112f
C12902 _078_ _045_ 7.44e-19
C12903 _141_/a_27_47# _049_ 4.22e-19
C12904 net55 _242_/a_382_297# 0.00129f
C12905 _336_/a_193_47# trim_mask\[4\] 0.0256f
C12906 _078_ _249_/a_109_297# 1.15e-19
C12907 _110_ _057_ 0.0685f
C12908 _308_/a_193_47# _307_/a_27_47# 6.5e-21
C12909 _308_/a_27_47# _307_/a_193_47# 1.21e-19
C12910 _104_ _239_/a_27_297# 1.47e-22
C12911 result[5] net29 6.48e-20
C12912 _232_/a_114_297# en_co_clk 4.78e-19
C12913 _321_/a_651_413# _101_ 8.49e-19
C12914 _306_/a_448_47# net51 6.51e-21
C12915 _334_/a_27_47# _031_ 0.0341f
C12916 net37 rebuffer2/a_75_212# 1.32e-20
C12917 _303_/a_193_47# _041_ 1.89e-19
C12918 net47 _303_/a_1270_413# -2.55e-20
C12919 _303_/a_1108_47# _338_/a_27_47# 3.5e-19
C12920 _303_/a_1283_21# _338_/a_193_47# 1.98e-19
C12921 _300_/a_47_47# net46 6.86e-20
C12922 _337_/a_1283_21# _263_/a_79_21# 7.38e-22
C12923 _268_/a_75_212# _332_/a_27_47# 5.61e-20
C12924 clknet_0_clk clkbuf_2_3__f_clk/a_110_47# 0.0209f
C12925 _335_/a_448_47# net46 0.00515f
C12926 _281_/a_253_47# _049_ 8.9e-20
C12927 _328_/a_448_47# _058_ 0.00115f
C12928 clk _331_/a_543_47# 0.00889f
C12929 state\[0\] _318_/a_27_47# 0.00104f
C12930 _060_ _318_/a_448_47# 3.19e-20
C12931 _290_/a_207_413# _125_ 0.0669f
C12932 output31/a_27_47# trim[0] 0.00927f
C12933 _258_/a_109_47# _280_/a_75_212# 3.49e-20
C12934 net12 _331_/a_761_289# 7.17e-20
C12935 net28 _313_/a_1217_47# 8.92e-19
C12936 net27 net26 1.42e-19
C12937 net4 _280_/a_75_212# 3.38e-19
C12938 _078_ mask\[4\] 0.083f
C12939 net8 output34/a_27_47# 0.00119f
C12940 _329_/a_639_47# trim_mask\[2\] 1.57e-19
C12941 _074_ _314_/a_448_47# 1.14e-19
C12942 VPWR _258_/a_109_297# -0.00489f
C12943 _048_ net55 0.907f
C12944 _324_/a_543_47# net44 0.0102f
C12945 _014_ _092_ 5.33e-19
C12946 net45 _099_ 0.0026f
C12947 _332_/a_1108_47# net46 0.0494f
C12948 net3 _100_ 3.82e-21
C12949 net4 _198_/a_181_47# 4.12e-19
C12950 _308_/a_27_47# _308_/a_448_47# -0.00373f
C12951 _029_ net46 0.041f
C12952 _116_ _330_/a_1108_47# 1.53e-20
C12953 _041_ _339_/a_796_47# 0.00181f
C12954 clknet_2_1__leaf_clk _085_ 0.196f
C12955 _078_ _220_/a_199_47# 1.28e-19
C12956 VPWR _313_/a_1462_47# 8.13e-20
C12957 _002_ rebuffer5/a_161_47# 2.85e-20
C12958 _256_/a_109_297# clknet_2_2__leaf_clk 0.00629f
C12959 net4 _331_/a_543_47# 1.41e-19
C12960 trim_mask\[4\] net55 6.4e-20
C12961 _304_/a_448_47# _001_ 0.0214f
C12962 result[0] _307_/a_761_289# 5.27e-19
C12963 cal _315_/a_193_47# 0.00305f
C12964 net1 _315_/a_27_47# 4.25e-19
C12965 _169_/a_215_311# net45 2.97e-19
C12966 _074_ _310_/a_761_289# 0.0091f
C12967 net39 net34 0.0575f
C12968 _322_/a_761_289# net44 0.0197f
C12969 net47 _297_/a_285_47# 1.15e-19
C12970 _233_/a_27_297# _093_ 0.0437f
C12971 _233_/a_109_297# calibrate 0.0282f
C12972 _289_/a_68_297# _125_ 0.00518f
C12973 _126_ _288_/a_59_75# 0.0258f
C12974 _065_ _099_ 3.14e-19
C12975 _041_ net53 0.106f
C12976 net21 _313_/a_1108_47# 0.00661f
C12977 _046_ _313_/a_651_413# 4.33e-19
C12978 _051_ _331_/a_639_47# 2.63e-19
C12979 state\[2\] _318_/a_639_47# 2.38e-19
C12980 _321_/a_1108_47# _083_ 4.68e-23
C12981 _325_/a_27_47# _321_/a_27_47# 1.3e-21
C12982 _270_/a_59_75# _058_ 0.00281f
C12983 _050_ clone1/a_27_47# 0.00933f
C12984 output7/a_27_47# ctln[1] 0.0105f
C12985 net43 _081_ 0.00795f
C12986 _290_/a_207_413# net40 1.78e-19
C12987 _311_/a_193_47# _311_/a_761_289# -0.00517f
C12988 _311_/a_27_47# _311_/a_543_47# -0.00482f
C12989 _306_/a_27_47# _002_ 0.00358f
C12990 trim[1] rebuffer2/a_75_212# 2.73e-19
C12991 net12 _101_ 0.0151f
C12992 _341_/a_761_289# cal_count\[3\] 0.0186f
C12993 state\[0\] _097_ 4.23e-21
C12994 _338_/a_1296_47# clknet_2_3__leaf_clk 3.98e-19
C12995 _135_ net37 1.53e-20
C12996 VPWR _338_/a_1602_47# 0.00364f
C12997 clknet_2_3__leaf_clk net18 0.0822f
C12998 _341_/a_651_413# clknet_2_3__leaf_clk 0.00499f
C12999 _323_/a_1283_21# _303_/a_543_47# 3.62e-19
C13000 _323_/a_27_47# _303_/a_651_413# 4.77e-20
C13001 _323_/a_651_413# _303_/a_27_47# 2.28e-20
C13002 net50 _256_/a_109_47# 2.29e-19
C13003 _067_ trim_mask\[4\] 6.2e-21
C13004 _316_/a_639_47# net41 0.0043f
C13005 VPWR _273_/a_59_75# 0.0192f
C13006 _339_/a_193_47# _339_/a_1032_413# -9.67e-21
C13007 _129_ trimb[4] 0.00203f
C13008 net13 _320_/a_1283_21# 0.0124f
C13009 _078_ _020_ 3.53e-21
C13010 _336_/a_1462_47# trim_mask\[4\] 0.00226f
C13011 _033_ clknet_2_2__leaf_clk 0.759f
C13012 clknet_2_3__leaf_clk _129_ 3e-21
C13013 _276_/a_59_75# _335_/a_193_47# 1.13e-21
C13014 VPWR output18/a_27_47# 0.0623f
C13015 _187_/a_297_47# _061_ 9.21e-19
C13016 cal_count\[3\] _098_ 1.22e-20
C13017 trim_mask\[1\] _334_/a_193_47# 1.13e-20
C13018 output15/a_27_47# _085_ 0.0257f
C13019 VPWR _240_/a_109_297# -5.4e-19
C13020 _272_/a_81_21# _334_/a_27_47# 4.16e-20
C13021 _320_/a_193_47# _040_ 0.0371f
C13022 VPWR _214_/a_113_297# 0.0464f
C13023 _096_ _241_/a_105_352# 1.46e-19
C13024 clknet_2_1__leaf_clk _314_/a_543_47# 6.19e-19
C13025 _307_/a_761_289# net14 0.00982f
C13026 cal _014_ 3e-20
C13027 net1 clknet_2_0__leaf_clk 1.47e-19
C13028 _015_ state\[1\] 0.0493f
C13029 _307_/a_1283_21# _138_/a_27_47# 0.00116f
C13030 _051_ _242_/a_79_21# 2.03e-20
C13031 _336_/a_651_413# _279_/a_396_47# 6.53e-20
C13032 _326_/a_761_289# net29 7.76e-20
C13033 mask\[1\] _319_/a_1283_21# 9.46e-20
C13034 VPWR _316_/a_639_47# 1.96e-19
C13035 _228_/a_382_297# _170_/a_299_297# 3.58e-19
C13036 _289_/a_68_297# net40 0.00492f
C13037 net44 _101_ 0.158f
C13038 clknet_0_clk cal_count\[3\] 1.76e-20
C13039 cal_itt\[2\] _306_/a_27_47# 2.48e-21
C13040 clknet_2_1__leaf_clk rebuffer4/a_27_47# 0.012f
C13041 _059_ _049_ 0.00658f
C13042 _029_ _332_/a_448_47# 0.00235f
C13043 VPWR clkbuf_2_2__f_clk/a_110_47# 0.0544f
C13044 _032_ net46 0.0294f
C13045 _169_/a_109_53# _243_/a_27_297# 6.94e-21
C13046 _244_/a_27_297# net51 0.00395f
C13047 VPWR _320_/a_193_47# -0.209f
C13048 net2 _068_ 0.00928f
C13049 _047_ _333_/a_1283_21# 0.0012f
C13050 _339_/a_1032_413# trimb[4] 2.64e-22
C13051 _050_ _337_/a_27_47# 1.51e-19
C13052 trim_mask\[2\] _119_ 0.104f
C13053 _286_/a_505_21# _123_ 0.0371f
C13054 _305_/a_1283_21# _068_ 6.01e-19
C13055 _322_/a_27_47# clknet_0_clk 1.13e-19
C13056 _064_ rebuffer3/a_75_212# 0.00294f
C13057 clknet_0_clk _331_/a_27_47# 0.0133f
C13058 _322_/a_193_47# _320_/a_1283_21# 1.65e-20
C13059 _322_/a_27_47# _320_/a_1108_47# 3.32e-20
C13060 _326_/a_1108_47# _251_/a_27_297# 2.95e-19
C13061 _326_/a_27_47# net26 0.00144f
C13062 _323_/a_448_47# net53 1.6e-21
C13063 _200_/a_303_47# _062_ 3.3e-19
C13064 trim_val\[0\] net32 1.68e-19
C13065 net7 _317_/a_543_47# 1.06e-19
C13066 net15 _317_/a_1108_47# 0.0035f
C13067 _074_ net51 5.04e-19
C13068 _101_ _003_ 5.74e-19
C13069 _308_/a_27_47# _005_ 0.0798f
C13070 clk net19 0.039f
C13071 _110_ _027_ 0.00725f
C13072 _258_/a_27_297# clknet_2_2__leaf_clk 0.0569f
C13073 _024_ clknet_2_2__leaf_clk 0.153f
C13074 mask\[0\] _120_ 0.00193f
C13075 trim_val\[1\] rebuffer1/a_75_212# 8.86e-20
C13076 _308_/a_651_413# net14 0.00291f
C13077 output35/a_27_47# output5/a_27_47# 3.56e-20
C13078 VPWR _323_/a_1270_413# -1.52e-19
C13079 VPWR _307_/a_761_289# 0.00267f
C13080 _290_/a_297_47# net37 0.00147f
C13081 _053_ net45 5.85e-20
C13082 _314_/a_1270_413# net29 1.14e-19
C13083 cal_count\[1\] _122_ 0.113f
C13084 _329_/a_543_47# _026_ 0.00188f
C13085 output29/a_27_47# _314_/a_1283_21# 5.15e-19
C13086 _329_/a_543_47# VPWR 0.033f
C13087 _053_ rebuffer3/a_75_212# 1.3e-19
C13088 calibrate _012_ 0.189f
C13089 net23 _320_/a_193_47# 6.01e-21
C13090 net43 _320_/a_1283_21# 3.85e-19
C13091 state\[2\] _243_/a_27_297# 5.29e-21
C13092 _321_/a_27_47# net25 9.67e-20
C13093 _305_/a_27_47# _305_/a_448_47# -0.00642f
C13094 _305_/a_193_47# _305_/a_1108_47# -0.00656f
C13095 _064_ _105_ 3.99e-19
C13096 _075_ _049_ 0.119f
C13097 _250_/a_27_297# _311_/a_27_47# 1.96e-20
C13098 net4 net19 0.346f
C13099 _309_/a_27_47# _309_/a_193_47# -0.019f
C13100 clk _107_ 0.0308f
C13101 cal_count\[1\] _299_/a_27_413# 4.98e-21
C13102 _103_ _053_ 9.49e-19
C13103 _272_/a_384_47# net46 1.37e-19
C13104 _231_/a_161_47# net4 0.005f
C13105 net44 _312_/a_448_47# 3.52e-19
C13106 _310_/a_1283_21# net29 1.08e-21
C13107 trim_mask\[3\] _258_/a_109_47# 0.0017f
C13108 _275_/a_81_21# trim_mask\[2\] 2.87e-21
C13109 _323_/a_193_47# _000_ 2.54e-19
C13110 _053_ _065_ 0.218f
C13111 _320_/a_193_47# net52 0.00316f
C13112 net24 _017_ 0.00128f
C13113 clknet_2_1__leaf_clk _311_/a_193_47# 0.00342f
C13114 trim_mask\[3\] net4 9.76e-21
C13115 _303_/a_1108_47# clknet_2_3__leaf_clk 0.0604f
C13116 _319_/a_805_47# _092_ 2.63e-21
C13117 _019_ _041_ 8.1e-20
C13118 _110_ _335_/a_448_47# 0.00206f
C13119 _305_/a_448_47# net51 0.00158f
C13120 net43 _307_/a_1108_47# 1.76e-19
C13121 _005_ _307_/a_448_47# 2.65e-19
C13122 _114_ _334_/a_761_289# 0.00204f
C13123 trim_val\[2\] _334_/a_1108_47# 0.00116f
C13124 _320_/a_1462_47# _040_ 6.28e-19
C13125 _053_ _105_ 0.0933f
C13126 VPWR _308_/a_651_413# 0.00229f
C13127 result[0] net43 6.17e-20
C13128 _306_/a_1283_21# cal_itt\[3\] 0.00464f
C13129 _306_/a_543_47# _072_ 1.35e-19
C13130 net4 _107_ 0.0857f
C13131 _065_ _208_/a_535_374# 0.00104f
C13132 _337_/a_193_47# _092_ 5.56e-19
C13133 _337_/a_543_47# _095_ 3.65e-19
C13134 net13 _040_ 0.171f
C13135 net3 _316_/a_193_47# 1.57e-20
C13136 net13 net41 0.00634f
C13137 _128_ _339_/a_27_47# 6.99e-19
C13138 net4 _001_ 0.0163f
C13139 _166_/a_161_47# net4 0.0367f
C13140 net16 _334_/a_1108_47# 2.65e-19
C13141 VPWR _237_/a_218_374# 2.64e-19
C13142 _250_/a_109_297# _074_ 9.52e-21
C13143 trim_mask\[0\] _109_ 0.103f
C13144 _303_/a_27_47# _303_/a_448_47# -0.00297f
C13145 trim[1] _112_ 4.99e-21
C13146 _110_ _029_ 1.78e-19
C13147 VPWR _320_/a_1462_47# 6.24e-19
C13148 net54 net55 0.395f
C13149 _060_ _096_ 0.0587f
C13150 _290_/a_27_413# cal_count\[0\] 7.71e-19
C13151 _064_ _194_/a_113_297# 0.0042f
C13152 VPWR _339_/a_381_47# -7.23e-19
C13153 _302_/a_27_297# _092_ 0.0121f
C13154 _064_ _336_/a_1283_21# 2.96e-19
C13155 _104_ _336_/a_761_289# 0.0473f
C13156 _324_/a_27_47# net20 0.0134f
C13157 _062_ cal_itt\[3\] 2.91e-19
C13158 _051_ _050_ 0.507f
C13159 VPWR net13 1.11f
C13160 _324_/a_27_47# net53 0.0107f
C13161 _048_ _121_ 1.12e-20
C13162 _326_/a_193_47# _078_ 0.0225f
C13163 output14/a_27_47# _011_ 1.29e-19
C13164 ctlp[0] _225_/a_109_297# 4.39e-19
C13165 _333_/a_1108_47# _055_ 0.00518f
C13166 net15 clknet_2_0__leaf_clk 0.153f
C13167 _106_ _092_ 2.91e-20
C13168 _104_ clone1/a_27_47# 1.3e-19
C13169 VPWR output28/a_27_47# 0.044f
C13170 net9 _334_/a_448_47# 3.67e-19
C13171 _308_/a_651_413# net23 9.76e-19
C13172 _308_/a_805_47# net43 5.25e-19
C13173 _001_ _122_ 0.589f
C13174 _337_/a_1108_47# _034_ 1.97e-19
C13175 _242_/a_297_47# _098_ 0.0523f
C13176 _322_/a_193_47# _040_ 1.3e-20
C13177 net43 net14 2.29f
C13178 VPWR _324_/a_761_289# 0.0151f
C13179 _059_ state\[1\] 0.00785f
C13180 VPWR net39 0.0374f
C13181 _053_ _194_/a_113_297# 2.1e-19
C13182 _143_/a_68_297# mask\[1\] 0.00832f
C13183 _195_/a_76_199# cal_itt\[3\] 4.72e-20
C13184 _309_/a_761_289# net43 -2.12e-19
C13185 _024_ _279_/a_204_297# 6.23e-22
C13186 trim_mask\[0\] _279_/a_490_47# 3.36e-19
C13187 _037_ _001_ 7.89e-19
C13188 _187_/a_297_47# net16 4.92e-19
C13189 net4 _279_/a_27_47# 5.29e-20
C13190 _042_ _247_/a_27_297# 0.0322f
C13191 _053_ _304_/a_761_289# 0.00917f
C13192 VPWR _198_/a_27_47# 0.0264f
C13193 _313_/a_1108_47# _045_ 7.2e-20
C13194 cal_itt\[1\] _195_/a_439_47# 9.57e-19
C13195 _308_/a_1108_47# _016_ 6.48e-19
C13196 _005_ _245_/a_27_297# 7.7e-20
C13197 _305_/a_27_47# _002_ 0.152f
C13198 net16 _332_/a_761_289# 0.00716f
C13199 VPWR _322_/a_193_47# -0.16f
C13200 _329_/a_761_289# clknet_2_2__leaf_clk 4.82e-20
C13201 _314_/a_193_47# _086_ 8.56e-20
C13202 VPWR _257_/a_109_297# 1.05e-19
C13203 VPWR _331_/a_193_47# 0.035f
C13204 net9 _335_/a_1283_21# 1.72e-19
C13205 _311_/a_1283_21# net26 0.0499f
C13206 _189_/a_27_47# _227_/a_109_93# 2.21e-20
C13207 _325_/a_193_47# _010_ 3.98e-19
C13208 _015_ _167_/a_161_47# 0.0131f
C13209 net43 _040_ 8.69e-20
C13210 _233_/a_109_297# _315_/a_27_47# 1.46e-19
C13211 _233_/a_27_297# _315_/a_193_47# 9.55e-19
C13212 en_co_clk clkc 0.00312f
C13213 _309_/a_193_47# _101_ 2.73e-19
C13214 _320_/a_27_47# _209_/a_27_47# 2.73e-21
C13215 _331_/a_27_47# _331_/a_1108_47# -2.98e-20
C13216 _041_ _205_/a_27_47# 0.0753f
C13217 VPWR _303_/a_651_413# 0.00128f
C13218 _269_/a_299_297# _112_ 0.00116f
C13219 _323_/a_639_47# net19 8.84e-19
C13220 _110_ _032_ 0.111f
C13221 cal_itt\[0\] _124_ 7.19e-19
C13222 _291_/a_35_297# _129_ 7.54e-21
C13223 _002_ net51 0.0071f
C13224 _327_/a_193_47# _136_ 0.0014f
C13225 trim_mask\[0\] _092_ 0.00122f
C13226 net13 net52 0.0204f
C13227 net35 _047_ 2.85e-19
C13228 net9 _332_/a_543_47# 5.4e-20
C13229 net9 _108_ 0.0117f
C13230 _094_ _234_/a_109_297# 0.00165f
C13231 _324_/a_27_47# _008_ 2.16e-20
C13232 VPWR net43 2.29f
C13233 trim[3] _179_/a_27_47# 7.28e-19
C13234 output34/a_27_47# net34 0.0248f
C13235 _337_/a_1462_47# _092_ 3.4e-20
C13236 cal_itt\[2\] _305_/a_27_47# 0.00128f
C13237 net3 _316_/a_1462_47# 9.82e-20
C13238 _036_ _339_/a_381_47# 0.00819f
C13239 _030_ net16 0.00367f
C13240 _058_ _172_/a_68_297# 1.31e-19
C13241 _189_/a_27_47# net42 1.7e-19
C13242 _058_ _136_ 0.153f
C13243 VPWR _309_/a_805_47# 2.95e-19
C13244 _064_ _302_/a_109_297# 0.00114f
C13245 _186_/a_109_297# net55 2.48e-19
C13246 _303_/a_27_47# _000_ 0.0291f
C13247 en_co_clk _096_ 0.0308f
C13248 _185_/a_68_297# net4 5.8e-20
C13249 _328_/a_639_47# net46 8.55e-19
C13250 _102_ mask\[3\] 1.05e-19
C13251 _023_ net25 1.3e-20
C13252 net24 _310_/a_27_47# 2.97e-21
C13253 net13 _164_/a_161_47# 4.35e-19
C13254 _292_/a_292_297# _128_ 0.00566f
C13255 trim[2] _108_ 4.34e-20
C13256 _336_/a_1108_47# _330_/a_1108_47# 6.38e-21
C13257 _198_/a_27_47# _063_ 0.0778f
C13258 _169_/a_301_53# _051_ 3.97e-19
C13259 trim[0] trim[2] 0.0391f
C13260 _065_ rebuffer4/a_27_47# 0.0332f
C13261 _328_/a_761_289# _030_ 7.31e-20
C13262 _322_/a_543_47# _101_ 0.00139f
C13263 _322_/a_193_47# net52 5.82e-23
C13264 VPWR _297_/a_129_47# -7.45e-19
C13265 _007_ _006_ 0.00117f
C13266 _188_/a_27_47# net37 0.0139f
C13267 clkbuf_2_2__f_clk/a_110_47# _279_/a_396_47# 0.00226f
C13268 _265_/a_81_21# clknet_2_3__leaf_clk 3.16e-21
C13269 net9 _031_ 7.5e-19
C13270 net43 net23 0.043f
C13271 _226_/a_27_47# _206_/a_27_93# 6.99e-19
C13272 _305_/a_543_47# net30 8.41e-21
C13273 ctlp[7] _156_/a_27_47# 3.27e-19
C13274 _283_/a_75_212# _121_ 0.0102f
C13275 _097_ calibrate 0.0132f
C13276 _321_/a_1283_21# mask\[2\] 0.00221f
C13277 _189_/a_27_47# _054_ 3.69e-21
C13278 _189_/a_408_47# _049_ 9.24e-19
C13279 _048_ clknet_2_3__leaf_clk 2.42e-19
C13280 _189_/a_27_47# net30 0.00307f
C13281 _134_ trim_val\[0\] 1.07e-20
C13282 net8 _334_/a_761_289# 0.00805f
C13283 net28 net21 0.0199f
C13284 _293_/a_384_47# _125_ 0.0015f
C13285 clkbuf_2_1__f_clk/a_110_47# net30 3.38e-20
C13286 state\[2\] trim_mask\[0\] 0.00126f
C13287 state\[0\] fanout45/a_27_47# 4.75e-21
C13288 _078_ _039_ 0.2f
C13289 _327_/a_639_47# trim_mask\[0\] 5.51e-21
C13290 _327_/a_448_47# _024_ 0.0128f
C13291 net4 _118_ 0.00759f
C13292 output10/a_27_47# VPWR 0.0691f
C13293 net43 net52 0.151f
C13294 _305_/a_1217_47# _002_ 0.00102f
C13295 net43 _063_ 0.00244f
C13296 _026_ _025_ 0.00206f
C13297 VPWR _322_/a_1462_47# 0.00178f
C13298 VPWR _331_/a_1462_47# 7.03e-20
C13299 _250_/a_109_297# net26 5.73e-20
C13300 VPWR _025_ 0.0114f
C13301 trim_mask\[4\] clknet_2_3__leaf_clk 1.03e-21
C13302 _312_/a_543_47# net20 0.00959f
C13303 VPWR _260_/a_93_21# 0.00317f
C13304 _308_/a_543_47# _212_/a_113_297# 4.65e-19
C13305 _093_ _315_/a_761_289# 1.4e-19
C13306 _012_ _315_/a_27_47# 0.0374f
C13307 calibrate _315_/a_543_47# 0.00737f
C13308 _309_/a_1462_47# _101_ 4.66e-20
C13309 _324_/a_1108_47# _312_/a_1108_47# 4.89e-20
C13310 mask\[6\] clknet_2_1__leaf_clk 0.125f
C13311 clkbuf_2_3__f_clk/a_110_47# _279_/a_204_297# 2.91e-21
C13312 _257_/a_27_297# clknet_2_2__leaf_clk 0.0282f
C13313 _331_/a_27_47# clknet_2_2__leaf_clk 0.0409f
C13314 _324_/a_543_47# net19 6.58e-20
C13315 _053_ clkbuf_0_clk/a_110_47# 8.73e-19
C13316 net33 net37 0.841f
C13317 net2 cal_itt\[3\] 2.98e-22
C13318 _327_/a_1462_47# _136_ 1.06e-19
C13319 _159_/a_27_47# net21 0.00333f
C13320 VPWR _312_/a_1108_47# 0.0149f
C13321 net15 _319_/a_639_47# 7.77e-19
C13322 _232_/a_114_297# _049_ 2.35e-19
C13323 _320_/a_761_289# mask\[1\] 0.0192f
C13324 net42 _227_/a_109_93# 2.25e-19
C13325 _305_/a_543_47# _072_ 0.00622f
C13326 _305_/a_1283_21# cal_itt\[3\] 1.82e-20
C13327 clkbuf_2_0__f_clk/a_110_47# mask\[0\] 0.00815f
C13328 _321_/a_27_47# net15 0.0128f
C13329 _074_ _086_ 0.0331f
C13330 _104_ _051_ 0.00947f
C13331 _235_/a_382_297# net55 8.92e-19
C13332 trim_val\[3\] _280_/a_75_212# 4.87e-21
C13333 result[4] _102_ 2.99e-20
C13334 cal_itt\[2\] _305_/a_1217_47# 1.19e-20
C13335 net3 net14 0.0121f
C13336 net16 trim_mask\[1\] 0.0189f
C13337 _189_/a_27_47# _072_ 5.62e-20
C13338 _189_/a_218_47# cal_itt\[3\] 1.94e-19
C13339 net15 _337_/a_27_47# 2.65e-20
C13340 _235_/a_79_21# _337_/a_27_47# 5.73e-21
C13341 _080_ net14 0.00104f
C13342 _067_ net40 3.32e-19
C13343 _320_/a_1283_21# fanout44/a_27_47# 2.76e-20
C13344 trim[1] _188_/a_27_47# 8.91e-21
C13345 output8/a_27_47# _108_ 9.16e-20
C13346 net8 rebuffer1/a_75_212# 4.41e-20
C13347 trim[4] net32 0.00269f
C13348 _170_/a_81_21# _049_ 0.0483f
C13349 _323_/a_193_47# mask\[4\] 0.00134f
C13350 net31 _131_ 0.0059f
C13351 clknet_0_clk _190_/a_215_47# 2.56e-19
C13352 _058_ _301_/a_129_47# 7.04e-20
C13353 _059_ _337_/a_1108_47# 4.98e-19
C13354 net50 _257_/a_109_297# 0.00363f
C13355 _337_/a_639_47# en_co_clk 4.18e-19
C13356 _303_/a_1270_413# net19 9.48e-20
C13357 _012_ clknet_2_0__leaf_clk 0.00553f
C13358 _093_ net45 0.0295f
C13359 calibrate _211_/a_109_297# 2.18e-19
C13360 _033_ _330_/a_1283_21# 1.15e-20
C13361 _336_/a_543_47# net46 -9.92e-19
C13362 _328_/a_27_47# _112_ 2.47e-21
C13363 _328_/a_761_289# trim_mask\[1\] 0.0188f
C13364 net5 _187_/a_212_413# 6.96e-19
C13365 _227_/a_296_53# _049_ 1.28e-19
C13366 _227_/a_109_93# _054_ 7.34e-20
C13367 VPWR _333_/a_543_47# 0.0201f
C13368 _087_ _242_/a_79_21# 5.14e-20
C13369 output15/a_27_47# mask\[6\] 5.65e-21
C13370 _291_/a_35_297# _297_/a_47_47# 1.75e-19
C13371 _227_/a_109_93# net30 0.00138f
C13372 net3 net41 0.00983f
C13373 fanout47/a_27_47# cal_count\[0\] 1.46e-20
C13374 _341_/a_1108_47# _092_ 8.65e-22
C13375 VPWR _265_/a_384_47# -1.33e-19
C13376 _136_ en_co_clk 0.00657f
C13377 _200_/a_80_21# cal_itt\[0\] 0.0302f
C13378 _200_/a_209_297# cal_itt\[2\] 0.00592f
C13379 net31 net5 0.0416f
C13380 _053_ _038_ 0.0563f
C13381 net12 _156_/a_27_47# 2.04e-19
C13382 _337_/a_1270_413# _076_ 3.59e-20
C13383 _093_ _065_ 0.0062f
C13384 _284_/a_68_297# en_co_clk 0.0135f
C13385 _263_/a_382_297# _090_ 0.00164f
C13386 _168_/a_27_413# _227_/a_109_93# 1.68e-19
C13387 mask\[7\] _222_/a_199_47# 5.21e-21
C13388 VPWR net3 2.49f
C13389 _288_/a_145_75# _122_ 5.55e-20
C13390 _053_ _338_/a_476_47# 9.6e-21
C13391 VPWR _080_ 0.181f
C13392 trim[1] net33 0.00648f
C13393 result[1] _078_ 4.11e-20
C13394 _190_/a_27_47# clknet_2_3__leaf_clk 3.8e-20
C13395 _179_/a_27_47# _057_ 0.0249f
C13396 trim[2] _272_/a_81_21# 2e-19
C13397 output33/a_27_47# trim_val\[2\] 0.00947f
C13398 _004_ _039_ 1.08e-19
C13399 _320_/a_193_47# _141_/a_27_47# 0.00913f
C13400 _250_/a_109_47# _078_ 1.96e-19
C13401 _237_/a_76_199# _095_ 0.00196f
C13402 net42 _054_ 1.86e-19
C13403 _323_/a_193_47# _020_ 0.00933f
C13404 _285_/a_113_47# _065_ 8.6e-21
C13405 net42 net30 0.00662f
C13406 _060_ _098_ 3.68e-19
C13407 _320_/a_1108_47# mask\[4\] 8.26e-21
C13408 _337_/a_1108_47# _075_ 0.00231f
C13409 _064_ trim_mask\[2\] 0.385f
C13410 _321_/a_27_47# _310_/a_193_47# 1.7e-22
C13411 _321_/a_193_47# _310_/a_27_47# 1.77e-21
C13412 net2 _131_ 0.072f
C13413 _135_ cal_count\[2\] 7.17e-20
C13414 _331_/a_448_47# trim_mask\[4\] 1.05e-19
C13415 _331_/a_805_47# _028_ 6.71e-19
C13416 _331_/a_1217_47# clknet_2_2__leaf_clk 2.72e-20
C13417 _051_ _226_/a_303_47# 7.24e-19
C13418 output33/a_27_47# net16 7.09e-19
C13419 _327_/a_27_47# clknet_2_3__leaf_clk 3.43e-20
C13420 _260_/a_93_21# _260_/a_346_47# -3.48e-20
C13421 net13 _248_/a_109_47# 6.47e-19
C13422 VPWR _325_/a_543_47# 0.0061f
C13423 _093_ _243_/a_109_297# 0.00354f
C13424 net4 _330_/a_761_289# 0.00111f
C13425 _309_/a_27_47# mask\[1\] 5.17e-20
C13426 net24 clknet_2_1__leaf_clk 0.0488f
C13427 _117_ _277_/a_75_212# 0.0342f
C13428 net42 _168_/a_27_413# 3.84e-21
C13429 _060_ clknet_0_clk 1.05e-20
C13430 _048_ _266_/a_68_297# 0.0478f
C13431 VPWR output34/a_27_47# 0.0626f
C13432 net23 _080_ 0.186f
C13433 net27 _010_ 1.37e-19
C13434 _325_/a_761_289# _159_/a_27_47# 0.00118f
C13435 _042_ _150_/a_27_47# 0.0295f
C13436 _064_ _329_/a_27_47# 3.82e-21
C13437 _094_ _337_/a_1283_21# 6.51e-19
C13438 _010_ _222_/a_113_297# 0.00151f
C13439 net13 _185_/a_150_297# 3.34e-19
C13440 _323_/a_1462_47# mask\[4\] 0.00237f
C13441 _287_/a_75_212# cal_count\[0\] 4.82e-19
C13442 _051_ net15 2.07e-20
C13443 net5 net2 9.9e-19
C13444 _051_ _235_/a_79_21# 1.18e-20
C13445 _318_/a_193_47# _318_/a_651_413# -0.00701f
C13446 net12 _077_ 0.00266f
C13447 net30 _054_ 0.00711f
C13448 output10/a_27_47# net50 0.00167f
C13449 _306_/a_1283_21# clk 0.0142f
C13450 _061_ clkc 4.9e-19
C13451 _302_/a_27_297# net46 4.03e-20
C13452 _266_/a_68_297# trim_mask\[4\] 1.75e-20
C13453 VPWR _241_/a_388_297# 6.64e-19
C13454 net12 _306_/a_543_47# 0.00752f
C13455 net50 _025_ 9.84e-20
C13456 _011_ net29 0.00552f
C13457 _050_ _119_ 2.53e-20
C13458 _080_ net52 2.07e-22
C13459 _325_/a_448_47# net43 0.00299f
C13460 net43 _216_/a_113_297# 3.67e-19
C13461 net13 _034_ 0.00173f
C13462 net42 _072_ 1.06e-20
C13463 _320_/a_27_47# mask\[2\] 0.00131f
C13464 _289_/a_68_297# _132_ 0.00342f
C13465 _106_ net46 9.94e-21
C13466 _168_/a_297_47# _049_ 7.02e-19
C13467 _168_/a_27_413# _054_ 0.00299f
C13468 trim_mask\[2\] _057_ 2.32e-20
C13469 _082_ net14 0.00888f
C13470 _210_/a_113_297# _315_/a_193_47# 3.16e-20
C13471 _168_/a_27_413# net30 0.00119f
C13472 clk _062_ 0.0102f
C13473 _107_ _260_/a_250_297# 0.0013f
C13474 _127_ _126_ 0.00987f
C13475 _309_/a_761_289# _082_ 5.07e-21
C13476 cal_itt\[0\] _071_ 6.03e-19
C13477 _322_/a_761_289# mask\[1\] 2.24e-20
C13478 trim_val\[3\] net19 5.82e-23
C13479 _333_/a_761_289# clknet_2_2__leaf_clk 1.54e-20
C13480 _303_/a_27_47# mask\[4\] 9.47e-20
C13481 net44 _077_ 0.00501f
C13482 net22 net30 0.0562f
C13483 VPWR fanout44/a_27_47# 0.0766f
C13484 clkbuf_2_1__f_clk/a_110_47# _319_/a_1108_47# 0.00376f
C13485 _308_/a_193_47# fanout43/a_27_47# 0.00553f
C13486 _318_/a_27_47# clknet_2_0__leaf_clk 0.0142f
C13487 _164_/a_161_47# net3 0.0238f
C13488 _325_/a_543_47# net52 5.95e-20
C13489 _325_/a_1108_47# _101_ 2.63e-19
C13490 mask\[3\] _245_/a_109_297# 2.59e-20
C13491 _091_ _108_ 3.2e-20
C13492 _015_ net13 0.171f
C13493 _306_/a_543_47# net44 0.00118f
C13494 _256_/a_109_297# _108_ 7.11e-19
C13495 net26 _086_ 6.86e-21
C13496 _293_/a_299_297# cal_count\[0\] 0.0317f
C13497 cal_itt\[2\] _262_/a_109_297# 7.66e-20
C13498 _326_/a_27_47# _102_ 7.75e-20
C13499 _326_/a_193_47# mask\[7\] 0.0141f
C13500 _050_ _087_ 6.6e-20
C13501 _329_/a_27_47# _057_ 1.44e-20
C13502 trim_val\[3\] trim_mask\[3\] 0.413f
C13503 _123_ _131_ 2.67e-19
C13504 _341_/a_448_47# _053_ 2.94e-20
C13505 _249_/a_27_297# net53 0.0809f
C13506 VPWR _190_/a_465_47# -3.62e-19
C13507 _048_ _028_ 8.13e-20
C13508 _162_/a_27_47# rebuffer2/a_75_212# 3.09e-20
C13509 clkbuf_2_2__f_clk/a_110_47# _330_/a_543_47# 0.00978f
C13510 net4 _062_ 0.34f
C13511 _047_ _332_/a_27_47# 1.63e-20
C13512 mask\[3\] net53 0.00172f
C13513 net15 _316_/a_1283_21# 0.0144f
C13514 _328_/a_193_47# _328_/a_651_413# -0.00701f
C13515 net30 _072_ 0.00455f
C13516 _103_ _171_/a_27_47# 1.75e-19
C13517 _340_/a_193_47# cal_count\[0\] 4.99e-21
C13518 _305_/a_27_47# _067_ 1.18e-20
C13519 _305_/a_27_47# _070_ 3.36e-21
C13520 _305_/a_1108_47# _202_/a_297_47# 3.77e-19
C13521 _328_/a_651_413# net9 0.00125f
C13522 net32 _108_ 2.14e-19
C13523 VPWR _249_/a_109_47# -3.5e-19
C13524 net13 _141_/a_27_47# 0.00464f
C13525 _248_/a_109_297# _101_ 0.0266f
C13526 _028_ trim_mask\[4\] 0.0918f
C13527 trim[0] net32 0.00352f
C13528 trim_mask\[0\] net46 0.351f
C13529 VPWR _327_/a_761_289# 0.0166f
C13530 _306_/a_1283_21# _073_ 0.00125f
C13531 _306_/a_543_47# _003_ 2.39e-19
C13532 VPWR _082_ 0.292f
C13533 _302_/a_373_47# _108_ 8.63e-21
C13534 _317_/a_448_47# net45 1.84e-21
C13535 _317_/a_543_47# state\[1\] 1.69e-19
C13536 _317_/a_1270_413# clknet_2_0__leaf_clk 6.2e-19
C13537 output16/a_27_47# ctlp[2] 0.00883f
C13538 _115_ _057_ 1.61e-20
C13539 clknet_0_clk en_co_clk 0.0377f
C13540 _074_ _313_/a_27_47# 0.0119f
C13541 _315_/a_193_47# _315_/a_761_289# -0.00541f
C13542 _257_/a_373_47# trim_val\[4\] 2.41e-20
C13543 _270_/a_59_75# net16 0.00339f
C13544 net4 _195_/a_76_199# 0.0136f
C13545 mask\[1\] _101_ 0.267f
C13546 _322_/a_448_47# mask\[3\] 0.0168f
C13547 _033_ _108_ 6.2e-21
C13548 net51 _070_ 1.36e-20
C13549 net43 _034_ 0.021f
C13550 _050_ _263_/a_297_47# 2.23e-20
C13551 _110_ _336_/a_543_47# 0.00179f
C13552 trimb[1] _125_ 0.00521f
C13553 _259_/a_109_47# VPWR -9.77e-19
C13554 _333_/a_1283_21# _333_/a_1108_47# 5.68e-32
C13555 _333_/a_27_47# _333_/a_639_47# -0.00188f
C13556 _303_/a_27_47# _020_ 0.00106f
C13557 _062_ _073_ 5.27e-20
C13558 _329_/a_193_47# _330_/a_1108_47# 1.79e-21
C13559 output33/a_27_47# _176_/a_27_47# 0.00817f
C13560 _097_ clknet_2_0__leaf_clk 1.42e-19
C13561 fanout44/a_27_47# net52 4.86e-20
C13562 _046_ _158_/a_68_297# 7.47e-19
C13563 _320_/a_1283_21# _076_ 5.33e-20
C13564 _320_/a_543_47# _077_ 2.5e-20
C13565 _306_/a_193_47# clknet_0_clk 8.12e-20
C13566 _265_/a_299_297# trim_val\[0\] 6.27e-19
C13567 calibrate fanout45/a_27_47# 1.6e-20
C13568 net27 _153_/a_27_47# 0.00138f
C13569 output21/a_27_47# clknet_2_1__leaf_clk 7.72e-20
C13570 _322_/a_1108_47# mask\[4\] 1.63e-20
C13571 _063_ _190_/a_465_47# 0.0154f
C13572 trim_val\[2\] _056_ 0.215f
C13573 _334_/a_761_289# net34 5.32e-21
C13574 _008_ _249_/a_27_297# 1.5e-20
C13575 _330_/a_1108_47# net18 1.78e-36
C13576 _078_ _315_/a_1108_47# 1.81e-19
C13577 _023_ _310_/a_193_47# 4.6e-19
C13578 VPWR _281_/a_103_199# 0.0284f
C13579 _192_/a_505_280# _065_ 0.00195f
C13580 _014_ _315_/a_761_289# 1.89e-20
C13581 net45 _315_/a_193_47# -9.81e-19
C13582 clknet_2_0__leaf_clk _315_/a_543_47# 0.00107f
C13583 cal_itt\[1\] _065_ 0.00318f
C13584 _089_ _092_ 1.2e-20
C13585 _090_ _095_ 0.132f
C13586 _125_ trimb[4] 0.00214f
C13587 _296_/a_113_47# _131_ 7.51e-19
C13588 trim[4] _130_ 2.59e-20
C13589 net16 _056_ 0.00292f
C13590 _321_/a_193_47# clknet_2_1__leaf_clk 0.131f
C13591 trim_mask\[0\] _332_/a_448_47# 5.1e-19
C13592 _024_ _108_ 0.0014f
C13593 output32/a_27_47# _055_ 6.66e-22
C13594 cal_itt\[1\] _105_ 4.25e-19
C13595 _326_/a_1462_47# mask\[7\] 0.00136f
C13596 _079_ net30 0.0937f
C13597 _286_/a_535_374# _122_ 2.48e-19
C13598 result[5] net14 8.01e-20
C13599 _124_ _338_/a_193_47# 1.13e-19
C13600 _242_/a_79_21# _099_ 5.38e-19
C13601 net37 output40/a_27_47# 0.00597f
C13602 _324_/a_639_47# mask\[5\] 1.48e-19
C13603 _006_ _310_/a_761_289# 2.15e-19
C13604 _074_ _215_/a_109_297# 0.00107f
C13605 _305_/a_1217_47# _067_ 2.25e-21
C13606 net5 _296_/a_113_47# 1.24e-19
C13607 _061_ _136_ 0.00202f
C13608 _322_/a_27_47# mask\[2\] 0.0965f
C13609 net16 clkc 3e-20
C13610 net34 rebuffer1/a_75_212# 4.93e-19
C13611 net24 net45 2.76e-20
C13612 result[2] clknet_2_0__leaf_clk 0.00281f
C13613 _079_ net22 0.152f
C13614 _014_ net45 0.345f
C13615 _187_/a_27_413# _301_/a_47_47# 0.0264f
C13616 cal_itt\[0\] _197_/a_113_297# 0.0641f
C13617 net31 _055_ 0.131f
C13618 trimb[4] net40 0.00278f
C13619 _211_/a_109_297# clknet_2_0__leaf_clk 0.00371f
C13620 cal_count\[3\] _278_/a_27_47# 1.1e-19
C13621 _256_/a_109_47# trim_mask\[1\] 0.00171f
C13622 clknet_2_3__leaf_clk net40 0.00271f
C13623 _122_ _332_/a_193_47# 8.3e-20
C13624 trim_mask\[0\] _269_/a_81_21# 3.76e-20
C13625 net27 net20 0.0479f
C13626 _301_/a_47_47# _332_/a_27_47# 7.08e-21
C13627 trim_mask\[4\] _279_/a_314_297# 1.27e-19
C13628 net8 ctln[3] 2.28e-19
C13629 _327_/a_193_47# clknet_2_2__leaf_clk 0.114f
C13630 _019_ mask\[3\] 0.0341f
C13631 net27 net53 1.42e-19
C13632 _104_ _119_ 0.103f
C13633 _190_/a_655_47# net19 0.00661f
C13634 clk net2 2.48e-20
C13635 _319_/a_651_413# _049_ 2.26e-19
C13636 net13 _059_ 0.00434f
C13637 _110_ _106_ 0.0826f
C13638 _218_/a_199_47# mask\[5\] 1.96e-20
C13639 _319_/a_1108_47# net30 1.04e-20
C13640 _060_ _263_/a_79_21# 0.0144f
C13641 net54 _263_/a_382_297# 2.94e-19
C13642 state\[2\] _089_ 3.47e-21
C13643 _305_/a_1283_21# clk 0.00454f
C13644 _329_/a_27_47# _027_ 2.54e-19
C13645 VPWR _330_/a_27_47# 0.0149f
C13646 _339_/a_27_47# _286_/a_76_199# 5.71e-21
C13647 _048_ _095_ 0.0407f
C13648 _312_/a_639_47# _045_ 1.15e-19
C13649 _096_ _049_ 0.0741f
C13650 net24 _065_ 3.63e-21
C13651 cal_itt\[0\] _194_/a_199_47# 2.4e-19
C13652 mask\[5\] _312_/a_193_47# 1.47e-20
C13653 net12 _305_/a_543_47# 3.3e-19
C13654 _323_/a_27_47# _068_ 1.08e-20
C13655 net49 net32 1.42e-20
C13656 VPWR result[5] 0.144f
C13657 _058_ clknet_2_2__leaf_clk 0.0751f
C13658 _259_/a_109_297# clknet_2_2__leaf_clk 6.37e-21
C13659 cal_itt\[1\] _304_/a_761_289# 1.88e-19
C13660 _189_/a_218_47# clk 0.00292f
C13661 _321_/a_1108_47# _018_ 2.29e-21
C13662 cal_count\[1\] _288_/a_59_75# 0.0268f
C13663 _292_/a_493_297# _125_ 2.04e-21
C13664 net2 net4 0.00902f
C13665 _341_/a_1108_47# net46 -0.00937f
C13666 mask\[0\] _319_/a_1283_21# 0.0494f
C13667 VPWR _120_ 0.137f
C13668 net6 ctln[0] 0.0627f
C13669 _040_ _076_ 3.91e-20
C13670 net45 _315_/a_1462_47# 5.4e-19
C13671 _319_/a_193_47# clknet_2_0__leaf_clk 0.605f
C13672 _321_/a_1270_413# _042_ 2.02e-19
C13673 _325_/a_1108_47# _248_/a_27_297# 4.4e-20
C13674 _305_/a_543_47# net44 0.00943f
C13675 output11/a_27_47# net19 2.97e-19
C13676 net44 _311_/a_651_413# 0.00125f
C13677 _293_/a_299_297# net16 0.00195f
C13678 _107_ trim_val\[4\] 9.3e-19
C13679 _259_/a_109_47# net50 9.28e-19
C13680 _104_ _275_/a_81_21# 6.99e-22
C13681 _064_ _275_/a_384_47# 8.95e-20
C13682 _259_/a_373_47# trim_mask\[3\] 0.00244f
C13683 output28/a_27_47# _314_/a_27_47# 0.0132f
C13684 _189_/a_27_47# net44 3.35e-21
C13685 net3 _034_ 2.54e-21
C13686 VPWR _076_ 0.621f
C13687 _340_/a_956_413# _123_ 0.00237f
C13688 _110_ trim_mask\[0\] 0.0683f
C13689 net13 _075_ 2.54e-20
C13690 clknet_2_1__leaf_clk _313_/a_1270_413# 3.05e-19
C13691 clkbuf_2_1__f_clk/a_110_47# net44 0.00139f
C13692 state\[0\] _090_ 1.04e-19
C13693 cal_itt\[0\] _035_ 0.0171f
C13694 _340_/a_193_47# net16 1.08e-20
C13695 VPWR _306_/a_761_289# 0.015f
C13696 _008_ net27 9.66e-23
C13697 _312_/a_761_289# _084_ 2.17e-20
C13698 valid sample 0.0379f
C13699 net2 _122_ 0.244f
C13700 _301_/a_285_47# _300_/a_285_47# 0.00178f
C13701 _326_/a_761_289# net14 0.00502f
C13702 fanout43/a_27_47# _016_ 2.63e-19
C13703 _176_/a_27_47# _056_ 0.0264f
C13704 net43 _059_ 1.7e-19
C13705 _065_ _243_/a_27_297# 1.46e-19
C13706 _335_/a_1108_47# net18 0.00662f
C13707 _322_/a_1217_47# mask\[2\] 3.77e-21
C13708 clkbuf_2_3__f_clk/a_110_47# _108_ 1.24e-19
C13709 _058_ _333_/a_651_413# 6.29e-19
C13710 net35 _333_/a_1108_47# 3.91e-20
C13711 _037_ net2 1.05e-19
C13712 _015_ net3 0.0538f
C13713 net2 _299_/a_27_413# 9.13e-19
C13714 _061_ _301_/a_129_47# 2.39e-19
C13715 _071_ _069_ 4.41e-20
C13716 _058_ trim_val\[0\] 0.0634f
C13717 net33 cal_count\[2\] 3.22e-19
C13718 fanout45/a_27_47# _317_/a_1108_47# 6.5e-20
C13719 _232_/a_32_297# net4 2.27e-21
C13720 _050_ _099_ 2.42e-19
C13721 mask\[7\] _251_/a_27_297# 0.0115f
C13722 _253_/a_384_47# net26 0.00117f
C13723 mask\[3\] _205_/a_27_47# 5.26e-20
C13724 net9 _340_/a_652_21# 0.00712f
C13725 _134_ _332_/a_543_47# 1.86e-19
C13726 _134_ _108_ 3.3e-20
C13727 _217_/a_109_297# _082_ 3.1e-19
C13728 _307_/a_193_47# _074_ 0.0168f
C13729 clk _227_/a_209_311# 5.87e-19
C13730 _315_/a_1108_47# _096_ 4.88e-19
C13731 en_co_clk _263_/a_79_21# 3.16e-19
C13732 _326_/a_193_47# net28 4.64e-20
C13733 _111_ net18 7.79e-21
C13734 _279_/a_27_47# trim_val\[4\] 0.0299f
C13735 net43 _306_/a_1108_47# 1.11e-19
C13736 VPWR _330_/a_1217_47# 8.79e-20
C13737 _339_/a_27_47# cal_count\[0\] 0.491f
C13738 output8/a_27_47# ctln[2] 0.0108f
C13739 _169_/a_215_311# _050_ 3.11e-19
C13740 _216_/a_113_297# _082_ 0.00941f
C13741 _090_ _226_/a_27_47# 8.61e-20
C13742 _087_ _226_/a_303_47# 9.6e-20
C13743 _304_/a_193_47# _065_ 0.0205f
C13744 _337_/a_639_47# _049_ 7.11e-19
C13745 _317_/a_193_47# _316_/a_27_47# 6.94e-21
C13746 clk _317_/a_761_289# 0.00393f
C13747 _317_/a_27_47# _316_/a_193_47# 1.35e-20
C13748 net43 _314_/a_27_47# 0.0144f
C13749 clknet_2_0__leaf_clk _206_/a_27_93# 5.13e-20
C13750 ctlp[0] result[6] 4.71e-19
C13751 trim_val\[1\] _055_ 0.112f
C13752 VPWR _326_/a_761_289# 0.0124f
C13753 net52 _076_ 0.0165f
C13754 _051_ _318_/a_27_47# 9.02e-20
C13755 _329_/a_761_289# _031_ 1.76e-19
C13756 trim_val\[2\] _172_/a_68_297# 5.43e-19
C13757 VPWR _334_/a_761_289# 0.019f
C13758 _019_ net27 4.53e-21
C13759 VPWR ctln[4] 0.0197f
C13760 _164_/a_161_47# _120_ 5.12e-20
C13761 net4 _227_/a_209_311# 2.66e-21
C13762 _181_/a_68_297# trim_val\[4\] 0.029f
C13763 state\[0\] _048_ 0.0114f
C13764 net3 _281_/a_253_47# 2.32e-20
C13765 _320_/a_543_47# clkbuf_2_1__f_clk/a_110_47# 4.44e-19
C13766 _046_ _085_ 0.0687f
C13767 _321_/a_1108_47# _078_ 1.62e-20
C13768 net16 _172_/a_68_297# 0.00115f
C13769 _307_/a_448_47# _039_ 1.22e-19
C13770 VPWR _286_/a_505_21# -0.0105f
C13771 _291_/a_35_297# _125_ 0.023f
C13772 _136_ net16 0.0255f
C13773 _330_/a_193_47# net19 0.0203f
C13774 _123_ _122_ 0.539f
C13775 cal_itt\[1\] clkbuf_0_clk/a_110_47# 0.0143f
C13776 _308_/a_448_47# _074_ 0.00411f
C13777 net12 net42 2.81e-20
C13778 net4 _317_/a_761_289# 0.00189f
C13779 state\[1\] _096_ 2.16e-19
C13780 _127_ net47 1.52e-20
C13781 _335_/a_193_47# _280_/a_75_212# 5.89e-20
C13782 _078_ _313_/a_193_47# 8.12e-19
C13783 _093_ _013_ 0.0321f
C13784 _300_/a_285_47# clknet_2_3__leaf_clk 0.0447f
C13785 _087_ _228_/a_79_21# 0.0111f
C13786 _101_ _062_ 3.72e-20
C13787 _337_/a_193_47# net45 2.77e-20
C13788 _337_/a_543_47# clknet_2_0__leaf_clk 0.00278f
C13789 VPWR _335_/a_27_47# 0.105f
C13790 result[6] _314_/a_1108_47# 1.96e-19
C13791 net28 _314_/a_651_413# 0.00362f
C13792 _037_ _123_ 0.0114f
C13793 _309_/a_761_289# _310_/a_1283_21# 3.87e-22
C13794 _323_/a_27_47# _042_ 0.05f
C13795 _309_/a_27_47# _310_/a_448_47# 1.58e-20
C13796 trim_mask\[3\] _330_/a_193_47# 8.52e-21
C13797 _326_/a_1108_47# net43 1.05e-19
C13798 _123_ _299_/a_27_413# 5.11e-22
C13799 _257_/a_27_297# _335_/a_1283_21# 1.03e-20
C13800 _323_/a_1283_21# clknet_2_1__leaf_clk 1.09e-20
C13801 _248_/a_373_47# mask\[4\] -6.68e-19
C13802 VPWR _314_/a_1270_413# 6.93e-20
C13803 cal_count\[3\] _108_ 0.00102f
C13804 _302_/a_27_297# rebuffer3/a_75_212# 1.03e-19
C13805 VPWR rebuffer1/a_75_212# 0.04f
C13806 clk _318_/a_1108_47# 0.0526f
C13807 _337_/a_193_47# _065_ 0.00349f
C13808 _236_/a_109_297# en_co_clk 2.11e-19
C13809 _233_/a_109_47# valid 1.39e-19
C13810 net28 _310_/a_543_47# 1.51e-20
C13811 mask\[5\] _152_/a_68_297# 0.0729f
C13812 _048_ _226_/a_27_47# 0.0335f
C13813 net12 _054_ 2.18e-21
C13814 _135_ _129_ 7.86e-20
C13815 net12 _318_/a_1283_21# 0.00577f
C13816 _290_/a_207_413# output37/a_27_47# 0.00114f
C13817 _074_ rebuffer6/a_27_47# 7.09e-21
C13818 net12 net30 0.011f
C13819 net9 _338_/a_27_47# 2.21e-19
C13820 _326_/a_761_289# net52 2.03e-19
C13821 fanout45/a_27_47# clknet_2_0__leaf_clk 4.69e-20
C13822 _257_/a_27_297# _108_ 1.61e-21
C13823 trim_mask\[2\] _272_/a_384_47# 0.00125f
C13824 _291_/a_35_297# net40 2.3e-20
C13825 result[1] _308_/a_27_47# 0.0203f
C13826 net9 _340_/a_1056_47# 3.98e-19
C13827 _324_/a_193_47# _074_ 8.1e-21
C13828 _304_/a_27_47# _304_/a_543_47# -0.00259f
C13829 _325_/a_761_289# mask\[2\] 1.27e-19
C13830 net54 _095_ 0.172f
C13831 _168_/a_207_413# clk 0.0154f
C13832 VPWR _310_/a_1283_21# 0.0466f
C13833 _302_/a_27_297# _065_ 0.0274f
C13834 trim_val\[4\] _118_ 0.304f
C13835 _340_/a_476_47# cal_count\[2\] 2.99e-20
C13836 _103_ _106_ 0.00163f
C13837 _327_/a_193_47# _327_/a_448_47# -0.00373f
C13838 _053_ _050_ 0.183f
C13839 _322_/a_27_47# _074_ 0.00841f
C13840 _304_/a_1462_47# _065_ 4.06e-19
C13841 VPWR _068_ 0.68f
C13842 cal_itt\[0\] _041_ 0.0129f
C13843 trim_val\[0\] en_co_clk 7.78e-20
C13844 net44 net30 0.0123f
C13845 clknet_2_2__leaf_clk _330_/a_805_47# 0.00252f
C13846 trim_mask\[4\] _330_/a_1108_47# 1.95e-22
C13847 _051_ _318_/a_1217_47# 5.08e-20
C13848 output27/a_27_47# _007_ 8.94e-20
C13849 _036_ _286_/a_505_21# 0.00106f
C13850 _168_/a_207_413# net4 8.59e-22
C13851 clkbuf_2_0__f_clk/a_110_47# net14 7.11e-22
C13852 _106_ _105_ 0.14f
C13853 _327_/a_448_47# _058_ 0.00438f
C13854 _059_ net3 0.0264f
C13855 _197_/a_113_297# _069_ 0.00932f
C13856 _334_/a_193_47# clknet_2_2__leaf_clk 0.00381f
C13857 _097_ _316_/a_1283_21# 5.84e-19
C13858 net9 net17 0.0215f
C13859 state\[2\] _092_ 2.44e-20
C13860 net12 _072_ 0.00247f
C13861 _311_/a_1283_21# net53 2.38e-20
C13862 trim_mask\[0\] rebuffer3/a_75_212# 3.37e-21
C13863 _205_/a_27_47# rebuffer5/a_161_47# 1.96e-19
C13864 _005_ _074_ 0.0772f
C13865 _274_/a_75_212# net48 1.93e-19
C13866 _162_/a_27_47# net33 0.00588f
C13867 _301_/a_129_47# net16 0.00162f
C13868 _090_ _052_ 1.32e-19
C13869 net30 _003_ 0.0681f
C13870 _282_/a_150_297# clknet_2_0__leaf_clk 8.17e-21
C13871 VPWR _335_/a_1217_47# 6.15e-20
C13872 _322_/a_193_47# _247_/a_109_297# 1.26e-20
C13873 _197_/a_199_47# _067_ 6.92e-19
C13874 VPWR _305_/a_761_289# 0.0157f
C13875 _197_/a_199_47# _070_ 3.51e-21
C13876 _275_/a_299_297# net46 6.39e-20
C13877 trim_mask\[3\] _330_/a_1462_47# 4.97e-19
C13878 _309_/a_639_47# _074_ 2.64e-19
C13879 VPWR _311_/a_448_47# -0.00272f
C13880 trim_mask\[0\] _103_ 0.232f
C13881 state\[2\] _169_/a_109_53# 1.05e-19
C13882 _305_/a_1108_47# _198_/a_27_47# 5.62e-20
C13883 net52 _310_/a_1283_21# 3.73e-19
C13884 _098_ _049_ 0.0909f
C13885 _051_ wire42/a_75_212# 2.15e-20
C13886 net16 _299_/a_382_47# 4.83e-19
C13887 net44 _072_ 0.477f
C13888 fanout46/a_27_47# _119_ 0.0686f
C13889 VPWR _332_/a_805_47# 0.00186f
C13890 _052_ _242_/a_382_297# 0.00147f
C13891 _304_/a_761_289# _302_/a_27_297# 4.37e-21
C13892 net9 _301_/a_285_47# 9.99e-20
C13893 _020_ _044_ 1.01e-19
C13894 _202_/a_382_297# _070_ 4.2e-19
C13895 net13 _232_/a_114_297# 0.00141f
C13896 VPWR clkbuf_2_0__f_clk/a_110_47# 0.106f
C13897 _068_ _063_ 0.647f
C13898 trim_mask\[0\] _105_ 0.00879f
C13899 clknet_0_clk _049_ 0.0925f
C13900 _304_/a_1283_21# _067_ 0.013f
C13901 output9/a_27_47# net18 5.56e-21
C13902 net9 _341_/a_543_47# 1.97e-19
C13903 _041_ clknet_2_0__leaf_clk 4.53e-21
C13904 _336_/a_193_47# _033_ 0.0412f
C13905 clk ctln[0] 0.0136f
C13906 output23/a_27_47# _005_ 0.0668f
C13907 _335_/a_193_47# net19 2.89e-20
C13908 _339_/a_562_413# _123_ 0.00224f
C13909 cal_itt\[2\] clkbuf_2_3__f_clk/a_110_47# 0.00843f
C13910 _289_/a_150_297# _129_ 3.83e-19
C13911 _289_/a_68_297# _130_ 3.28e-21
C13912 net43 _305_/a_1108_47# 0.0211f
C13913 net16 _339_/a_27_47# 6.15e-20
C13914 _214_/a_113_297# _078_ 0.0816f
C13915 _003_ _072_ 6.33e-20
C13916 _321_/a_27_47# _321_/a_543_47# -0.00936f
C13917 _321_/a_193_47# _321_/a_761_289# -0.0105f
C13918 net43 _146_/a_68_297# 0.0294f
C13919 net50 _335_/a_27_47# 0.00398f
C13920 trim_mask\[3\] _335_/a_193_47# 0.00315f
C13921 trim_val\[3\] _335_/a_761_289# 4.26e-20
C13922 _234_/a_109_297# _121_ 3.7e-19
C13923 _247_/a_27_297# _101_ 0.0482f
C13924 _042_ net14 1.65e-20
C13925 _008_ _311_/a_1283_21# 3.61e-20
C13926 _317_/a_27_47# net14 8.86e-19
C13927 _014_ _316_/a_448_47# 0.00439f
C13928 net45 _316_/a_1108_47# -0.00104f
C13929 _338_/a_652_21# _065_ 7.36e-20
C13930 _307_/a_27_47# _315_/a_27_47# 2.09e-19
C13931 net2 _101_ 3.53e-21
C13932 _169_/a_373_53# state\[0\] 2.78e-19
C13933 _329_/a_1108_47# net48 2.35e-20
C13934 state\[0\] net54 0.051f
C13935 cal_itt\[0\] net18 4.6e-19
C13936 net4 ctln[0] 0.0219f
C13937 _074_ net21 0.473f
C13938 _048_ _052_ 0.0522f
C13939 clkbuf_0_clk/a_110_47# _304_/a_193_47# 1.02e-19
C13940 _059_ fanout44/a_27_47# 1.22e-21
C13941 _167_/a_161_47# _096_ 4.21e-21
C13942 _320_/a_193_47# _078_ 3.94e-19
C13943 _305_/a_761_289# _063_ 4.1e-20
C13944 output32/a_27_47# _333_/a_1283_21# 9.15e-19
C13945 _337_/a_27_47# _337_/a_543_47# -0.00482f
C13946 _307_/a_1283_21# net30 6.9e-19
C13947 calibrate _090_ 0.0169f
C13948 output26/a_27_47# result[5] 0.00311f
C13949 result[4] output27/a_27_47# 1.02e-19
C13950 net2 _297_/a_285_47# 0.00117f
C13951 net9 _339_/a_193_47# 0.0164f
C13952 _309_/a_448_47# clknet_2_1__leaf_clk 2.63e-20
C13953 _257_/a_109_297# trim_mask\[1\] 0.00583f
C13954 mask\[1\] _077_ 4.87e-19
C13955 _091_ _067_ 0.00473f
C13956 clknet_2_1__leaf_clk _245_/a_373_47# 1.69e-19
C13957 trim_mask\[0\] _194_/a_113_297# 0.0371f
C13958 net28 _251_/a_27_297# 0.00115f
C13959 trim_mask\[4\] _052_ 0.144f
C13960 _250_/a_109_297# net53 0.00431f
C13961 trim_mask\[0\] _336_/a_1283_21# 5.37e-20
C13962 _317_/a_27_47# net41 1.11e-20
C13963 _333_/a_193_47# rebuffer2/a_75_212# 3.4e-20
C13964 _324_/a_193_47# net26 2.1e-21
C13965 _175_/a_150_297# _108_ 5.09e-19
C13966 _064_ _104_ 0.67f
C13967 _333_/a_193_47# _332_/a_1283_21# 5.72e-21
C13968 _333_/a_761_289# _108_ 0.00569f
C13969 _324_/a_1108_47# _042_ 1.03e-19
C13970 calibrate _242_/a_382_297# 2.4e-19
C13971 _307_/a_543_47# mask\[0\] 2.09e-20
C13972 _307_/a_1283_21# net22 0.0765f
C13973 _307_/a_761_289# _078_ 0.00235f
C13974 _259_/a_27_297# _330_/a_1108_47# 3.98e-19
C13975 _328_/a_1283_21# _329_/a_1108_47# 1.18e-19
C13976 _328_/a_1108_47# _329_/a_1283_21# 5.34e-20
C13977 VPWR _251_/a_109_297# -0.0145f
C13978 VPWR _250_/a_373_47# 3.11e-20
C13979 _029_ _333_/a_27_47# 2.08e-20
C13980 net15 _158_/a_68_297# 8.23e-19
C13981 _034_ _076_ 1.79e-20
C13982 net31 _333_/a_1283_21# 0.0177f
C13983 _265_/a_299_297# _332_/a_543_47# 9.16e-20
C13984 _265_/a_299_297# _108_ 0.0219f
C13985 _307_/a_27_47# clknet_2_0__leaf_clk 0.0258f
C13986 _324_/a_639_47# clknet_2_1__leaf_clk 3.14e-19
C13987 VPWR _042_ 6.28f
C13988 _329_/a_1270_413# net9 1.44e-19
C13989 output34/a_27_47# _334_/a_1108_47# 5.37e-19
C13990 net9 clknet_2_3__leaf_clk 0.162f
C13991 clknet_0_clk _262_/a_193_297# 7.06e-19
C13992 _111_ _265_/a_81_21# 3.52e-20
C13993 _335_/a_1108_47# trim_mask\[4\] 4.24e-19
C13994 VPWR _317_/a_27_47# 0.0621f
C13995 _322_/a_27_47# net26 1.42e-20
C13996 output27/a_27_47# net27 0.0218f
C13997 clkbuf_2_0__f_clk/a_110_47# _164_/a_161_47# 5.09e-19
C13998 _235_/a_382_297# _095_ 1.16e-19
C13999 _235_/a_79_21# _099_ 6.65e-20
C14000 net15 _099_ 0.0134f
C14001 _246_/a_109_297# _017_ 0.00219f
C14002 _304_/a_193_47# _038_ 7.11e-21
C14003 _304_/a_1108_47# _136_ 5.64e-19
C14004 result[1] result[3] 0.00269f
C14005 _333_/a_805_47# net46 6.28e-20
C14006 net34 _131_ 0.0115f
C14007 _100_ clone7/a_27_47# 0.0701f
C14008 _104_ _053_ 0.802f
C14009 net43 _018_ 0.192f
C14010 output36/a_27_47# output37/a_27_47# 0.00254f
C14011 _083_ _311_/a_448_47# 4.21e-20
C14012 _109_ net46 3.12e-20
C14013 _332_/a_639_47# clknet_2_2__leaf_clk 5.75e-19
C14014 _273_/a_59_75# _056_ 8.32e-21
C14015 _051_ _206_/a_27_93# 0.0228f
C14016 _062_ _190_/a_655_47# 0.0401f
C14017 _200_/a_303_47# VPWR -9.05e-19
C14018 _048_ calibrate 0.12f
C14019 _113_ _333_/a_1283_21# 3.12e-21
C14020 _030_ _333_/a_543_47# 4.57e-19
C14021 _230_/a_145_75# net4 7.2e-19
C14022 net13 _318_/a_448_47# 0.00562f
C14023 _308_/a_651_413# _078_ 8.7e-19
C14024 _340_/a_27_47# _340_/a_956_413# -0.00135f
C14025 _275_/a_384_47# _032_ 7.95e-20
C14026 net50 _335_/a_1217_47# 1.51e-19
C14027 clknet_2_1__leaf_clk _312_/a_193_47# 0.0248f
C14028 net44 _319_/a_1108_47# 1.96e-19
C14029 net8 _273_/a_145_75# 1.62e-20
C14030 _128_ _290_/a_207_413# 3.1e-21
C14031 _308_/a_1108_47# clknet_2_0__leaf_clk 0.00133f
C14032 _219_/a_109_297# net26 1.97e-19
C14033 net5 net34 0.217f
C14034 _062_ trim_val\[4\] 8.95e-19
C14035 _014_ _013_ 0.0694f
C14036 _314_/a_1108_47# _158_/a_68_297# 7.54e-20
C14037 calibrate trim_mask\[4\] 0.0443f
C14038 _276_/a_59_75# net19 5.08e-21
C14039 _292_/a_292_297# net16 1.54e-20
C14040 _323_/a_193_47# _149_/a_68_297# 1.55e-20
C14041 _337_/a_193_47# _282_/a_68_297# 2.71e-19
C14042 _251_/a_373_47# _101_ 3.04e-19
C14043 _251_/a_109_297# net52 0.0411f
C14044 _309_/a_27_47# output24/a_27_47# 8.25e-19
C14045 _237_/a_76_199# clknet_2_0__leaf_clk 4.11e-20
C14046 net5 _301_/a_377_297# 5.38e-20
C14047 _195_/a_76_199# _190_/a_655_47# 6.49e-20
C14048 _313_/a_27_47# _313_/a_448_47# -0.00642f
C14049 _313_/a_193_47# _313_/a_1108_47# 1.42e-32
C14050 cal_itt\[0\] _303_/a_1108_47# 8.04e-19
C14051 cal_itt\[1\] _303_/a_1283_21# 4.77e-20
C14052 _336_/a_27_47# clkbuf_2_2__f_clk/a_110_47# 0.0189f
C14053 _042_ net52 0.0113f
C14054 _320_/a_805_47# clknet_2_0__leaf_clk 1.55e-19
C14055 _025_ trim_mask\[1\] 0.12f
C14056 _216_/a_113_297# _310_/a_1283_21# 0.00123f
C14057 net9 _339_/a_796_47# 2.99e-19
C14058 net15 _246_/a_27_297# 0.0109f
C14059 VPWR _318_/a_543_47# 0.0087f
C14060 net13 _078_ 0.0381f
C14061 output39/a_27_47# net38 4.96e-20
C14062 _110_ _275_/a_299_297# 0.0517f
C14063 _116_ _275_/a_81_21# 0.00305f
C14064 _276_/a_59_75# trim_mask\[3\] 2e-20
C14065 _276_/a_145_75# trim_val\[3\] 1.39e-20
C14066 _135_ _265_/a_81_21# 2.87e-21
C14067 _232_/a_304_297# _090_ 0.00148f
C14068 _021_ net20 1.25e-19
C14069 _189_/a_27_47# _107_ 0.00319f
C14070 _035_ _338_/a_193_47# 0.112f
C14071 _021_ net53 0.054f
C14072 _331_/a_543_47# _054_ 1.12e-20
C14073 trim_mask\[2\] _336_/a_543_47# 1.15e-20
C14074 _260_/a_93_21# _170_/a_81_21# 4.36e-19
C14075 net4 _336_/a_805_47# 4.25e-19
C14076 _128_ _289_/a_68_297# 2.16e-20
C14077 _312_/a_27_47# _009_ 0.212f
C14078 net4 _264_/a_27_297# 0.00976f
C14079 VPWR _022_ 0.118f
C14080 _328_/a_543_47# VPWR 0.0128f
C14081 _330_/a_27_47# _330_/a_543_47# -0.00936f
C14082 _330_/a_193_47# _330_/a_761_289# -0.0105f
C14083 _208_/a_76_199# _076_ 0.0236f
C14084 _200_/a_303_47# _063_ 0.00116f
C14085 _041_ _069_ 1.36e-19
C14086 _051_ fanout45/a_27_47# 3.53e-19
C14087 _302_/a_27_297# _038_ 0.0029f
C14088 VPWR ctln[3] 0.0154f
C14089 net46 _092_ 9.46e-20
C14090 _307_/a_761_289# _004_ 0.00175f
C14091 VPWR _317_/a_1217_47# 2.84e-20
C14092 mask\[7\] _313_/a_193_47# 2.26e-19
C14093 _304_/a_193_47# _298_/a_292_297# 8.14e-21
C14094 _322_/a_193_47# _078_ 0.0036f
C14095 mask\[6\] _046_ 0.075f
C14096 _133_ _131_ 0.00247f
C14097 net21 net26 2.96e-20
C14098 _319_/a_543_47# clknet_0_clk 8.27e-19
C14099 _050_ _093_ 2.32e-20
C14100 _326_/a_27_47# output27/a_27_47# 3.72e-19
C14101 _249_/a_27_297# _311_/a_27_47# 0.0111f
C14102 VPWR cal_itt\[3\] 0.204f
C14103 _341_/a_27_47# _066_ 0.0126f
C14104 _227_/a_109_93# net19 5.86e-21
C14105 _000_ net26 5.23e-20
C14106 net14 net6 0.00948f
C14107 _083_ _042_ 8.1e-20
C14108 _011_ net14 0.00251f
C14109 net51 _205_/a_27_47# 9.02e-20
C14110 _340_/a_27_47# _122_ 0.00249f
C14111 _112_ _333_/a_193_47# 0.0105f
C14112 trim_mask\[1\] _333_/a_543_47# 7.04e-19
C14113 net49 _333_/a_761_289# 0.0106f
C14114 trim_val\[1\] _333_/a_1283_21# 0.043f
C14115 net33 _129_ 2.66e-19
C14116 _293_/a_81_21# _299_/a_27_413# 9.18e-21
C14117 _304_/a_27_47# net18 0.00548f
C14118 trim[1] _182_/a_27_47# 0.00212f
C14119 output32/a_27_47# net35 0.00348f
C14120 _263_/a_79_21# _049_ 9.78e-19
C14121 _315_/a_448_47# net41 5.39e-20
C14122 _340_/a_1140_413# net47 -5.38e-19
C14123 _037_ _304_/a_1270_413# 8.96e-21
C14124 _060_ _094_ 1.56e-20
C14125 _315_/a_1283_21# valid 1.44e-19
C14126 net43 _078_ 2.58f
C14127 _259_/a_27_297# _335_/a_1108_47# 0.00164f
C14128 _259_/a_109_297# _335_/a_1283_21# 3.4e-19
C14129 _327_/a_193_47# _108_ 0.00281f
C14130 _340_/a_27_47# _037_ 0.0477f
C14131 _060_ _088_ 5.91e-21
C14132 net54 _052_ 1.63e-20
C14133 cal_count\[1\] _127_ 1.22e-19
C14134 _327_/a_27_47# _111_ 1.77e-19
C14135 _327_/a_1283_21# _268_/a_75_212# 0.01f
C14136 VPWR _262_/a_205_47# -4.58e-20
C14137 _253_/a_299_297# _023_ 9.1e-19
C14138 _309_/a_805_47# _078_ 0.00136f
C14139 _187_/a_212_413# net35 0.025f
C14140 _107_ _227_/a_109_93# 0.00575f
C14141 _090_ _192_/a_27_47# 5.02e-20
C14142 fanout45/a_27_47# _316_/a_1283_21# 0.0122f
C14143 _323_/a_1283_21# _043_ 0.0167f
C14144 VPWR _315_/a_448_47# 0.00423f
C14145 _074_ _045_ 0.158f
C14146 _022_ net52 0.00265f
C14147 _309_/a_651_413# net24 0.0265f
C14148 _337_/a_651_413# net44 7.12e-19
C14149 _074_ _249_/a_109_297# 3.35e-20
C14150 _313_/a_27_47# _010_ 0.0352f
C14151 cal_itt\[2\] _000_ 0.00363f
C14152 output17/a_27_47# ctlp[3] 0.00841f
C14153 net35 _332_/a_193_47# 8.54e-19
C14154 mask\[0\] _101_ 0.0411f
C14155 _058_ _332_/a_543_47# 0.00456f
C14156 _058_ _108_ 0.228f
C14157 net42 net19 5.45e-21
C14158 _233_/a_27_297# cal 0.00651f
C14159 _304_/a_1108_47# clknet_0_clk 1.9e-19
C14160 _082_ _310_/a_651_413# 9.17e-19
C14161 net55 clkbuf_2_3__f_clk/a_110_47# 1.03e-19
C14162 trim_mask\[0\] _038_ 3.83e-20
C14163 _239_/a_27_297# _048_ 1.64e-19
C14164 net31 net35 1.68e-19
C14165 net27 _314_/a_761_289# 3.66e-19
C14166 _327_/a_639_47# net46 4.64e-19
C14167 VPWR net6 0.188f
C14168 VPWR _011_ 0.382f
C14169 cal_count\[1\] _126_ 0.0948f
C14170 clk _316_/a_193_47# 6.05e-19
C14171 mask\[1\] clkbuf_2_1__f_clk/a_110_47# 0.0121f
C14172 net16 clknet_2_2__leaf_clk 1.2e-19
C14173 _239_/a_27_297# trim_mask\[4\] 1.85e-21
C14174 fanout47/a_27_47# _198_/a_27_47# 2.81e-20
C14175 _063_ cal_itt\[3\] 0.00277f
C14176 _149_/a_68_297# _303_/a_27_47# 5.08e-21
C14177 _104_ _027_ 0.145f
C14178 net47 net44 6.3e-19
C14179 net42 _107_ 0.0111f
C14180 _074_ mask\[4\] 0.189f
C14181 _292_/a_215_47# cal_count\[2\] 4.49e-19
C14182 _069_ net18 1.21e-20
C14183 _067_ clkbuf_2_3__f_clk/a_110_47# 0.00377f
C14184 _110_ _109_ 0.0292f
C14185 net30 net19 0.00891f
C14186 _304_/a_448_47# _133_ 8.76e-21
C14187 _328_/a_448_47# _025_ 0.00249f
C14188 _328_/a_761_289# clknet_2_2__leaf_clk 0.0443f
C14189 _322_/a_1462_47# _078_ 5.11e-19
C14190 _304_/a_1283_21# clknet_2_3__leaf_clk 4.73e-20
C14191 mask\[3\] _247_/a_373_47# 5.58e-19
C14192 _217_/a_109_297# _042_ 4.64e-22
C14193 _340_/a_1032_413# _298_/a_78_199# 0.00129f
C14194 _231_/a_161_47# net30 7.08e-21
C14195 _236_/a_109_297# _049_ 7.62e-20
C14196 VPWR _131_ 0.137f
C14197 _048_ _203_/a_59_75# 1.4e-20
C14198 net45 _331_/a_1270_413# 1.41e-19
C14199 _326_/a_1108_47# result[5] 1.11e-19
C14200 net15 _085_ 0.46f
C14201 _257_/a_27_297# _336_/a_193_47# 1.28e-19
C14202 clkbuf_2_0__f_clk/a_110_47# _034_ 4.34e-20
C14203 net54 calibrate 0.0341f
C14204 _215_/a_109_297# _006_ 0.00424f
C14205 _237_/a_505_21# net55 3.76e-21
C14206 _325_/a_27_47# mask\[6\] 0.151f
C14207 _048_ _192_/a_27_47# 0.0194f
C14208 cal_itt\[0\] _048_ -1.01e-24
C14209 net12 net44 0.0433f
C14210 _075_ _076_ 0.00538f
C14211 _041_ _338_/a_193_47# 1.06e-19
C14212 _216_/a_113_297# _042_ 4.09e-19
C14213 _337_/a_1108_47# clknet_0_clk 8.64e-21
C14214 clknet_2_0__leaf_clk _090_ 0.00154f
C14215 net47 _338_/a_562_413# 1.12e-19
C14216 _341_/a_27_47# net47 3.98e-21
C14217 en_co_clk _195_/a_218_374# 0.0029f
C14218 _094_ en_co_clk 0.112f
C14219 trim_mask\[2\] trim_mask\[0\] 2.63e-20
C14220 _107_ _054_ 0.00434f
C14221 _147_/a_27_47# net17 0.0045f
C14222 net35 net2 1.98e-20
C14223 net13 _096_ 0.649f
C14224 _107_ net30 0.239f
C14225 _294_/a_150_297# VPWR -6.63e-19
C14226 _064_ _335_/a_1270_413# 6.72e-20
C14227 _327_/a_1462_47# _108_ 4.2e-20
C14228 en_co_clk _088_ 9.79e-21
C14229 _015_ clkbuf_2_0__f_clk/a_110_47# 3.35e-20
C14230 _326_/a_543_47# output14/a_27_47# 1.43e-20
C14231 _050_ _171_/a_27_47# 0.0108f
C14232 _110_ _279_/a_490_47# 1.61e-20
C14233 VPWR net5 0.304f
C14234 _327_/a_1217_47# _111_ 1.58e-19
C14235 net16 _333_/a_651_413# 0.0056f
C14236 _340_/a_476_47# _129_ 6.87e-21
C14237 _239_/a_277_297# _050_ 7.3e-19
C14238 clknet_2_1__leaf_clk _158_/a_150_297# 6.18e-21
C14239 result[4] _310_/a_639_47# 3.91e-19
C14240 mask\[4\] _311_/a_805_47# 0.00207f
C14241 net16 trim_val\[0\] 0.0338f
C14242 net27 _311_/a_27_47# 1.98e-21
C14243 _168_/a_27_413# _107_ 0.00152f
C14244 VPWR _319_/a_1283_21# 0.0221f
C14245 net19 _072_ 7.43e-19
C14246 net12 _003_ 0.181f
C14247 _091_ clknet_2_3__leaf_clk 0.0011f
C14248 _053_ _124_ 1.67e-20
C14249 _313_/a_1217_47# _010_ 4.2e-20
C14250 VPWR _149_/a_150_297# 3.49e-19
C14251 _256_/a_109_297# clknet_2_3__leaf_clk 1.28e-20
C14252 _093_ net1 0.00103f
C14253 cal_count\[3\] net55 6.92e-20
C14254 _064_ fanout46/a_27_47# 0.00164f
C14255 output33/a_27_47# output34/a_27_47# 0.00243f
C14256 _314_/a_1108_47# _085_ 1.44e-20
C14257 net33 _297_/a_47_47# 0.0046f
C14258 net2 _288_/a_59_75# 0.057f
C14259 _326_/a_27_47# _314_/a_761_289# 4.89e-21
C14260 _326_/a_193_47# _314_/a_193_47# 6.68e-19
C14261 _303_/a_761_289# _035_ 7.91e-22
C14262 _341_/a_193_47# net4 1.23e-21
C14263 _043_ _303_/a_543_47# 7.66e-19
C14264 net44 _003_ 0.00506f
C14265 en_co_clk _108_ 7.36e-21
C14266 _302_/a_373_47# clknet_2_3__leaf_clk 0.00164f
C14267 net30 _279_/a_27_47# 7.15e-20
C14268 _330_/a_1270_413# _027_ 3.05e-19
C14269 ctlp[0] _314_/a_543_47# 0.00126f
C14270 _001_ _072_ 1.65e-20
C14271 net34 _055_ 0.161f
C14272 clkbuf_2_0__f_clk/a_110_47# _281_/a_253_47# 2.55e-19
C14273 en_co_clk _244_/a_27_297# 3.94e-20
C14274 _048_ clknet_2_0__leaf_clk 7.83e-20
C14275 _336_/a_1108_47# _119_ 3.82e-20
C14276 _067_ cal_count\[3\] 0.0363f
C14277 _080_ _078_ 5.82e-19
C14278 net35 trim_val\[1\] 0.00225f
C14279 _323_/a_543_47# _041_ 7.81e-21
C14280 _058_ net49 0.00402f
C14281 VPWR _336_/a_1270_413# 4.96e-19
C14282 _213_/a_109_297# net45 5.77e-21
C14283 _050_ _192_/a_505_280# 0.0264f
C14284 _303_/a_1108_47# _069_ 0.00103f
C14285 VPWR _304_/a_448_47# 0.00233f
C14286 _082_ _018_ 9.07e-20
C14287 net4 _316_/a_1462_47# 4.88e-20
C14288 _340_/a_652_21# cal_count\[3\] 8.19e-20
C14289 _107_ _262_/a_465_47# 3.06e-19
C14290 _340_/a_381_47# clknet_2_3__leaf_clk 0.00224f
C14291 _341_/a_1108_47# _038_ 3.1e-19
C14292 _341_/a_639_47# _136_ 9.98e-19
C14293 _186_/a_109_297# calibrate 0.00292f
C14294 _235_/a_297_47# _094_ 1.11e-19
C14295 _249_/a_109_297# net26 6.35e-20
C14296 _025_ _336_/a_27_47# 2.56e-21
C14297 clknet_2_1__leaf_clk _246_/a_109_297# 0.00544f
C14298 _325_/a_448_47# _022_ 0.00211f
C14299 _325_/a_1217_47# mask\[6\] 8.65e-19
C14300 _319_/a_761_289# _016_ 3.37e-19
C14301 _341_/a_193_47# _122_ 5.13e-19
C14302 _325_/a_543_47# _078_ 0.00122f
C14303 _161_/a_68_297# net37 0.00916f
C14304 _190_/a_27_47# _203_/a_59_75# 0.0134f
C14305 _306_/a_193_47# _244_/a_27_297# 3.15e-19
C14306 net54 _232_/a_304_297# 0.0016f
C14307 _015_ _317_/a_27_47# 9.18e-22
C14308 _338_/a_193_47# net18 0.0121f
C14309 clknet_2_1__leaf_clk mask\[5\] 0.0811f
C14310 _320_/a_27_47# _121_ 2.11e-20
C14311 _239_/a_474_297# _092_ 0.0755f
C14312 _228_/a_297_47# _088_ 1.57e-19
C14313 _320_/a_543_47# net44 -9.76e-19
C14314 _228_/a_382_297# _052_ 0.00143f
C14315 cal_itt\[2\] _190_/a_215_47# 0.0111f
C14316 cal_itt\[0\] _190_/a_27_47# 2.61e-20
C14317 _104_ _032_ 3.44e-21
C14318 net13 _313_/a_1108_47# 0.00232f
C14319 net13 _337_/a_639_47# 0.00101f
C14320 _321_/a_1283_21# net53 0.00285f
C14321 _169_/a_215_311# _318_/a_27_47# 2.83e-20
C14322 _332_/a_1283_21# net40 1.44e-20
C14323 _288_/a_59_75# _123_ 2.1e-21
C14324 mask\[4\] net26 0.591f
C14325 net28 _313_/a_193_47# 0.0253f
C14326 _111_ net40 0.0034f
C14327 _239_/a_694_21# _060_ 1.71e-19
C14328 _161_/a_150_297# net46 1.6e-19
C14329 VPWR _256_/a_373_47# -6.01e-19
C14330 _306_/a_1108_47# _068_ 9.75e-21
C14331 VPWR _321_/a_448_47# 0.00188f
C14332 _323_/a_805_47# net44 1.74e-19
C14333 clone1/a_27_47# _242_/a_382_297# 2.88e-19
C14334 net33 _175_/a_68_297# 0.0158f
C14335 _250_/a_27_297# _084_ 4.16e-19
C14336 mask\[1\] net22 1.8e-20
C14337 _333_/a_193_47# net33 1.54e-19
C14338 _041_ _339_/a_652_21# 0.0173f
C14339 VPWR _313_/a_761_289# 0.0207f
C14340 net36 net16 2.74e-19
C14341 net47 _339_/a_956_413# 4.53e-19
C14342 VPWR _337_/a_448_47# 7.64e-19
C14343 _212_/a_113_297# net45 0.00109f
C14344 _029_ _267_/a_59_75# 1.07e-19
C14345 _111_ _267_/a_145_75# 1.69e-19
C14346 _298_/a_78_199# _298_/a_292_297# -1.09e-21
C14347 clk net14 0.0521f
C14348 _334_/a_1108_47# rebuffer1/a_75_212# 3.8e-20
C14349 _316_/a_1108_47# _013_ 4.03e-21
C14350 _143_/a_68_297# _040_ 6.46e-21
C14351 _097_ _099_ 0.0211f
C14352 fanout44/a_27_47# _078_ 5.71e-21
C14353 _192_/a_639_47# _095_ 1.24e-19
C14354 _054_ _118_ 8.99e-21
C14355 net2 _077_ 8.99e-20
C14356 _237_/a_76_199# _316_/a_1283_21# 1.98e-19
C14357 _159_/a_27_47# _313_/a_193_47# 6.61e-20
C14358 _335_/a_27_47# _335_/a_543_47# -0.00214f
C14359 _015_ _318_/a_543_47# 8.44e-19
C14360 net30 _118_ 0.141f
C14361 output38/a_27_47# net34 0.0944f
C14362 _306_/a_543_47# net2 2.27e-20
C14363 trim[1] _161_/a_68_297# 2.18e-19
C14364 clkbuf_2_2__f_clk/a_110_47# clknet_0_clk 0.019f
C14365 _292_/a_215_47# _340_/a_1602_47# 6.57e-19
C14366 _122_ _133_ 0.109f
C14367 _337_/a_27_47# _090_ 5.41e-22
C14368 _093_ net15 0.00808f
C14369 _306_/a_193_47# _305_/a_448_47# 2.4e-19
C14370 _306_/a_1283_21# _305_/a_543_47# 1.1e-19
C14371 _326_/a_1283_21# _310_/a_1108_47# 3.98e-19
C14372 _326_/a_1108_47# _310_/a_1283_21# 3.09e-21
C14373 _320_/a_193_47# clknet_0_clk 9.18e-19
C14374 net43 _321_/a_639_47# 0.00354f
C14375 _283_/a_75_212# clknet_2_0__leaf_clk 0.0101f
C14376 ctln[1] net7 0.0086f
C14377 output37/a_27_47# trimb[1] 0.00971f
C14378 _326_/a_193_47# _074_ 0.0206f
C14379 VPWR _143_/a_68_297# 0.0182f
C14380 _338_/a_1032_413# clknet_2_3__leaf_clk 0.0853f
C14381 _320_/a_193_47# _320_/a_1108_47# -0.00656f
C14382 _320_/a_27_47# _320_/a_448_47# -0.00676f
C14383 net12 ctln[7] 0.00247f
C14384 _129_ output40/a_27_47# 2.28e-19
C14385 net4 net14 1.54e-19
C14386 _309_/a_27_47# _081_ 0.00169f
C14387 _037_ _133_ 0.0109f
C14388 _048_ clone1/a_27_47# 0.0259f
C14389 calibrate _228_/a_382_297# 0.00142f
C14390 _334_/a_639_47# net46 0.00323f
C14391 _060_ _192_/a_174_21# 2.07e-20
C14392 net54 _192_/a_27_47# 0.0079f
C14393 _200_/a_80_21# _053_ 0.0384f
C14394 clk net41 3.86e-20
C14395 VPWR _340_/a_956_413# -5.48e-19
C14396 _189_/a_27_47# _306_/a_1283_21# 5.38e-22
C14397 _329_/a_1108_47# _274_/a_75_212# 0.00253f
C14398 net43 _313_/a_1108_47# -0.0235f
C14399 _301_/a_285_47# _134_ 7.11e-33
C14400 _315_/a_1283_21# _095_ 8.55e-19
C14401 _020_ net26 3.23e-19
C14402 _299_/a_27_413# _133_ 3.3e-19
C14403 net55 _242_/a_297_47# 2.28e-19
C14404 _104_ _171_/a_27_47# 0.0483f
C14405 _336_/a_448_47# _028_ 4.1e-20
C14406 _336_/a_761_289# trim_mask\[4\] 0.0221f
C14407 clone7/a_27_47# net41 0.00163f
C14408 clknet_2_1__leaf_clk _017_ 6.06e-19
C14409 _116_ _057_ 6.5e-20
C14410 _328_/a_1283_21# _327_/a_1283_21# 1.65e-19
C14411 _308_/a_193_47# _307_/a_193_47# 0.0016f
C14412 _135_ net40 7.13e-19
C14413 _232_/a_220_297# en_co_clk 2.85e-19
C14414 _009_ _084_ 0.102f
C14415 _082_ _078_ 0.0538f
C14416 _230_/a_59_75# _107_ 2.31e-19
C14417 _306_/a_651_413# net51 3.67e-19
C14418 _321_/a_448_47# net52 6.06e-21
C14419 _321_/a_1270_413# _101_ 3.07e-19
C14420 _334_/a_193_47# _031_ 0.00405f
C14421 _338_/a_796_47# net18 4.63e-19
C14422 trim_mask\[4\] clone1/a_27_47# 9.23e-21
C14423 _000_ _070_ 6.75e-20
C14424 net24 net25 1.32e-20
C14425 mask\[3\] clknet_2_0__leaf_clk 1.61e-20
C14426 _332_/a_1108_47# net37 4.63e-20
C14427 VPWR clk 4.07f
C14428 _066_ net19 8.99e-21
C14429 _332_/a_27_47# _332_/a_193_47# -0.221f
C14430 net47 _303_/a_639_47# 5.51e-21
C14431 output34/a_27_47# _056_ 7.29e-19
C14432 _303_/a_1108_47# _338_/a_193_47# 9.13e-19
C14433 _337_/a_1270_413# _101_ 8.97e-21
C14434 _189_/a_27_47# _062_ 0.0498f
C14435 VPWR clone7/a_27_47# 0.00398f
C14436 _337_/a_1108_47# _263_/a_79_21# 3.12e-19
C14437 net4 net41 1.15e-19
C14438 _336_/a_639_47# net19 7.16e-19
C14439 ctlp[4] net18 0.00492f
C14440 _339_/a_1032_413# output40/a_27_47# 1.1e-20
C14441 _231_/a_161_47# _066_ 0.00683f
C14442 _328_/a_651_413# _058_ 5.41e-19
C14443 _335_/a_651_413# net46 0.0046f
C14444 _064_ _328_/a_27_47# 3.82e-21
C14445 _094_ _039_ 1.23e-20
C14446 output37/a_27_47# trimb[4] 2.97e-20
C14447 state\[0\] _318_/a_193_47# 4.22e-20
C14448 clk _331_/a_1283_21# 5.3e-21
C14449 _290_/a_297_47# _125_ 0.00172f
C14450 net12 _331_/a_543_47# 5.19e-20
C14451 net28 _313_/a_1462_47# 0.002f
C14452 _329_/a_805_47# trim_mask\[2\] 9.76e-20
C14453 VPWR _258_/a_109_47# -0.00104f
C14454 net43 mask\[7\] 0.0334f
C14455 _324_/a_1283_21# net44 0.00602f
C14456 VPWR net4 3.93f
C14457 net45 _092_ 0.00188f
C14458 net12 _229_/a_27_297# 0.00101f
C14459 _048_ _337_/a_27_47# 1.76e-20
C14460 _332_/a_448_47# net46 0.0162f
C14461 net3 _096_ 0.027f
C14462 fanout46/a_27_47# _027_ 2.72e-19
C14463 _308_/a_193_47# _308_/a_448_47# -0.00373f
C14464 _333_/a_1462_47# net33 7.82e-19
C14465 _041_ _339_/a_1056_47# 0.00208f
C14466 _143_/a_68_297# net52 0.00329f
C14467 _336_/a_639_47# _107_ 2.69e-19
C14468 _019_ _321_/a_1283_21# 0.002f
C14469 _304_/a_651_413# _001_ 1.44e-20
C14470 _103_ _092_ 0.0113f
C14471 _113_ _332_/a_27_47# 1.61e-20
C14472 result[0] _307_/a_543_47# 0.00117f
C14473 cal _315_/a_761_289# 6.15e-19
C14474 net1 _315_/a_193_47# 0.00824f
C14475 _322_/a_543_47# net44 0.00563f
C14476 clknet_2_3__leaf_clk _298_/a_215_47# 1.91e-20
C14477 _169_/a_109_53# net45 4.09e-21
C14478 _074_ _310_/a_543_47# 0.0136f
C14479 _314_/a_543_47# _224_/a_113_297# 9.8e-19
C14480 _292_/a_78_199# _122_ 0.0137f
C14481 clkbuf_2_3__f_clk/a_110_47# clknet_2_3__leaf_clk 0.0019f
C14482 _233_/a_109_297# _093_ 9.13e-19
C14483 _289_/a_150_297# _125_ 2.24e-19
C14484 _065_ _092_ 0.0108f
C14485 _046_ _313_/a_1270_413# 7.93e-21
C14486 net21 _313_/a_448_47# 5.49e-20
C14487 _214_/a_113_297# _245_/a_27_297# 2.2e-20
C14488 VPWR _055_ 0.294f
C14489 cal_count\[1\] net47 1.48e-20
C14490 _270_/a_145_75# _058_ 3.85e-20
C14491 net13 _098_ 2.72e-21
C14492 state\[2\] _318_/a_805_47# 1.41e-19
C14493 _325_/a_193_47# _321_/a_27_47# 5.65e-19
C14494 _325_/a_27_47# _321_/a_193_47# 2.01e-19
C14495 VPWR _122_ 0.532f
C14496 _134_ clknet_2_3__leaf_clk 0.0566f
C14497 clk _063_ 7.88e-20
C14498 _311_/a_193_47# _311_/a_543_47# -0.0129f
C14499 _306_/a_193_47# _002_ 0.00792f
C14500 _187_/a_27_413# net2 5.73e-21
C14501 _051_ _090_ 0.202f
C14502 VPWR _073_ 0.198f
C14503 _105_ _092_ 2.75e-20
C14504 _269_/a_81_21# net46 2.74e-20
C14505 output17/a_27_47# net16 5.69e-19
C14506 _341_/a_543_47# cal_count\[3\] 0.0299f
C14507 VPWR _338_/a_381_47# 1.32e-19
C14508 _341_/a_1270_413# clknet_2_3__leaf_clk 8.2e-20
C14509 en_co_clk _192_/a_174_21# 0.0229f
C14510 cal_itt\[2\] en_co_clk 0.253f
C14511 _323_/a_651_413# _303_/a_193_47# 1.92e-21
C14512 _323_/a_1108_47# _303_/a_543_47# 3.42e-20
C14513 net2 _332_/a_27_47# 2.97e-19
C14514 net13 clknet_0_clk 0.0596f
C14515 trim_mask\[0\] _242_/a_79_21# 2.03e-20
C14516 _071_ _053_ 0.00497f
C14517 _316_/a_805_47# net41 0.00208f
C14518 VPWR _037_ 0.889f
C14519 VPWR _273_/a_145_75# -6.36e-20
C14520 ctlp[6] net20 0.0765f
C14521 _339_/a_193_47# _339_/a_1602_47# -4.7e-21
C14522 _339_/a_27_47# _339_/a_381_47# -0.00538f
C14523 _033_ _028_ 7.86e-20
C14524 net13 _320_/a_1108_47# 0.014f
C14525 _081_ _101_ 0.024f
C14526 VPWR _299_/a_27_413# 0.0394f
C14527 _227_/a_109_93# _062_ 6.61e-21
C14528 _272_/a_299_297# _334_/a_27_47# 2.64e-20
C14529 _272_/a_81_21# _334_/a_193_47# 4.54e-19
C14530 _320_/a_761_289# _040_ 0.0236f
C14531 VPWR _214_/a_199_47# -4.76e-19
C14532 _053_ _262_/a_27_47# 0.0129f
C14533 trim[4] net16 4.7e-20
C14534 _074_ _039_ 4.18e-20
C14535 clknet_2_1__leaf_clk _314_/a_1283_21# 2.14e-20
C14536 output29/a_27_47# net15 1.16e-20
C14537 _307_/a_543_47# net14 0.00307f
C14538 net1 _014_ 1.44e-20
C14539 cal net45 3.14e-19
C14540 state\[2\] net45 0.0706f
C14541 net4 _063_ 0.0356f
C14542 _307_/a_1108_47# _138_/a_27_47# 8.52e-19
C14543 _051_ _242_/a_382_297# 1.34e-21
C14544 _326_/a_543_47# net29 1.9e-19
C14545 mask\[1\] _319_/a_1108_47# 2.41e-19
C14546 trim_mask\[0\] _333_/a_27_47# 4.34e-20
C14547 _332_/a_639_47# _108_ 0.00129f
C14548 _289_/a_150_297# net40 2.58e-19
C14549 output27/a_27_47# _086_ 8.35e-19
C14550 cal_itt\[2\] _306_/a_193_47# 8.89e-21
C14551 net47 net19 0.152f
C14552 _146_/a_68_297# _310_/a_1283_21# 9.04e-19
C14553 trimb[2] net38 0.00263f
C14554 VPWR _320_/a_761_289# 0.00188f
C14555 state\[2\] _103_ 0.00629f
C14556 _198_/a_27_47# clknet_0_clk 1.31e-19
C14557 _181_/a_68_297# _066_ 1.06e-20
C14558 _050_ _337_/a_193_47# 1.33e-19
C14559 ctlp[0] output29/a_27_47# 6.9e-19
C14560 output14/a_27_47# result[7] 0.0905f
C14561 _286_/a_218_374# _123_ 0.00109f
C14562 clknet_2_1__leaf_clk _310_/a_27_47# 0.0902f
C14563 _305_/a_1108_47# _068_ 1.61e-21
C14564 clknet_0_clk _331_/a_193_47# 0.00248f
C14565 result[5] _078_ 4.73e-20
C14566 _164_/a_161_47# net4 3.57e-20
C14567 mask\[6\] net15 0.0927f
C14568 ctlp[7] _155_/a_68_297# 0.00111f
C14569 _322_/a_193_47# _320_/a_1108_47# 5.87e-21
C14570 _322_/a_761_289# _320_/a_1283_21# 1.22e-19
C14571 _319_/a_1283_21# _034_ 1.22e-20
C14572 _316_/a_1283_21# _090_ 9.09e-20
C14573 _326_/a_1108_47# _251_/a_109_297# 1.24e-19
C14574 net42 _062_ 7.43e-19
C14575 _326_/a_193_47# net26 1.15e-20
C14576 trimb[0] net36 0.0043f
C14577 net15 _317_/a_448_47# 0.00169f
C14578 cal_itt\[0\] net40 5.38e-21
C14579 _308_/a_27_47# net43 0.0167f
C14580 _308_/a_193_47# _005_ 0.0903f
C14581 _116_ _027_ 1.29e-20
C14582 _063_ _073_ 1.41e-19
C14583 _110_ net46 0.393f
C14584 _258_/a_109_297# clknet_2_2__leaf_clk 0.00682f
C14585 input2/a_27_47# _131_ 0.0115f
C14586 _051_ _048_ 0.425f
C14587 _337_/a_27_47# _283_/a_75_212# 1.36e-19
C14588 trim_mask\[1\] rebuffer1/a_75_212# 2.07e-19
C14589 _306_/a_1283_21# net30 2.19e-20
C14590 net47 _001_ 0.0223f
C14591 VPWR _307_/a_543_47# 0.0108f
C14592 VPWR _323_/a_639_47# 7.45e-19
C14593 net14 _138_/a_27_47# 0.00511f
C14594 net43 clknet_0_clk 0.152f
C14595 _036_ _122_ 0.00237f
C14596 clknet_2_0__leaf_clk rebuffer5/a_161_47# 0.005f
C14597 cal_count\[3\] clknet_2_3__leaf_clk 0.519f
C14598 _329_/a_1283_21# _026_ 1.29e-20
C14599 _329_/a_1283_21# VPWR 0.03f
C14600 output29/a_27_47# _314_/a_1108_47# 7.19e-19
C14601 _309_/a_1108_47# _308_/a_1108_47# 2.99e-21
C14602 _093_ _012_ 0.0245f
C14603 _305_/a_543_47# net2 1.86e-19
C14604 net43 _320_/a_1108_47# 5.92e-19
C14605 _315_/a_27_47# sample 0.00261f
C14606 VPWR output38/a_27_47# 0.0873f
C14607 _309_/a_27_47# net14 0.0121f
C14608 _051_ trim_mask\[4\] 0.266f
C14609 _053_ wire42/a_75_212# 1.84e-20
C14610 _321_/a_27_47# mask\[3\] 0.00649f
C14611 _321_/a_193_47# net25 6.82e-20
C14612 _305_/a_193_47# _305_/a_448_47# -0.00297f
C14613 _036_ _037_ 2.57e-20
C14614 _062_ _054_ 1.53e-22
C14615 clkbuf_2_1__f_clk/a_110_47# _247_/a_27_297# 1.56e-20
C14616 _078_ _076_ 0.0104f
C14617 _119_ net18 1.51e-19
C14618 _188_/a_27_47# output35/a_27_47# 0.00787f
C14619 en_co_clk output5/a_27_47# 2.25e-19
C14620 _062_ net30 0.148f
C14621 _325_/a_1283_21# _313_/a_1283_21# 9.75e-19
C14622 net5 input2/a_27_47# 0.00102f
C14623 cal_count\[1\] _299_/a_215_297# 1.12e-20
C14624 net44 _312_/a_651_413# 0.00133f
C14625 net12 _107_ 0.0371f
C14626 net44 net19 0.0822f
C14627 _320_/a_1283_21# _101_ 5.34e-21
C14628 _320_/a_761_289# net52 7.52e-19
C14629 _306_/a_27_47# clknet_2_0__leaf_clk 0.0146f
C14630 clknet_2_1__leaf_clk _311_/a_761_289# 7.33e-21
C14631 _303_/a_448_47# clknet_2_3__leaf_clk 0.0138f
C14632 net12 _166_/a_161_47# 0.00737f
C14633 _110_ _335_/a_651_413# 7.89e-21
C14634 _305_/a_651_413# net51 7.46e-20
C14635 _271_/a_75_212# _112_ 7.61e-19
C14636 trim_val\[2\] _334_/a_448_47# 7.84e-20
C14637 _018_ _310_/a_1283_21# 3.75e-19
C14638 VPWR _308_/a_1270_413# 1.14e-19
C14639 _094_ _049_ 0.0783f
C14640 _273_/a_59_75# clknet_2_2__leaf_clk 0.00184f
C14641 _128_ trimb[1] 1.84e-19
C14642 _195_/a_76_199# net30 8.82e-21
C14643 _306_/a_1283_21# _072_ 0.00214f
C14644 _306_/a_1108_47# cal_itt\[3\] 0.0014f
C14645 _065_ _208_/a_218_47# 0.00117f
C14646 _337_/a_543_47# _099_ 1.53e-21
C14647 _337_/a_761_289# _092_ 1.3e-19
C14648 _266_/a_68_297# clkbuf_2_3__f_clk/a_110_47# 9.54e-19
C14649 _264_/a_27_297# trim_val\[4\] 3.83e-19
C14650 result[1] _074_ 0.00166f
C14651 net3 _316_/a_761_289# 2.15e-19
C14652 VPWR _138_/a_27_47# 0.0626f
C14653 _292_/a_215_47# _339_/a_1032_413# 1.16e-19
C14654 _128_ _339_/a_193_47# 8.08e-20
C14655 trim_mask\[0\] _050_ 3.24e-20
C14656 clknet_2_0__leaf_clk sample 0.236f
C14657 _088_ _049_ 0.0514f
C14658 _260_/a_93_21# _098_ 2.07e-21
C14659 net13 net28 3.54e-20
C14660 ctlp[2] ctlp[3] 0.00303f
C14661 _017_ _065_ 6.2e-21
C14662 net26 _310_/a_543_47# 2.08e-19
C14663 VPWR _237_/a_535_374# -2.59e-20
C14664 output41/a_27_47# valid 0.00805f
C14665 VPWR _309_/a_27_47# 0.0718f
C14666 _042_ _310_/a_651_413# 1.29e-20
C14667 _281_/a_103_199# _096_ 2.67e-20
C14668 _303_/a_193_47# _303_/a_448_47# -0.00297f
C14669 state\[0\] _243_/a_373_47# 6.15e-20
C14670 _325_/a_543_47# mask\[7\] 2.6e-20
C14671 _060_ net55 0.0944f
C14672 output28/a_27_47# net28 0.0296f
C14673 _290_/a_207_413# cal_count\[0\] 0.00352f
C14674 rebuffer6/a_27_47# net53 0.0129f
C14675 VPWR _339_/a_562_413# -6.69e-19
C14676 _341_/a_27_47# _231_/a_161_47# 4.77e-19
C14677 _302_/a_109_297# _092_ 0.00153f
C14678 output35/a_27_47# net33 0.0075f
C14679 _064_ _336_/a_1108_47# 1.31e-19
C14680 _104_ _336_/a_543_47# 0.0247f
C14681 net54 _337_/a_27_47# 0.00143f
C14682 clkbuf_2_2__f_clk/a_110_47# clknet_2_2__leaf_clk 0.0844f
C14683 _324_/a_193_47# net20 5.31e-21
C14684 _062_ _072_ 5.18e-20
C14685 _336_/a_27_47# _330_/a_27_47# 4.35e-20
C14686 _324_/a_193_47# net53 0.00258f
C14687 _019_ _320_/a_27_47# 1.79e-19
C14688 _053_ _197_/a_113_297# 3.07e-19
C14689 net30 _137_/a_68_297# 0.00208f
C14690 _275_/a_81_21# net18 0.00275f
C14691 _326_/a_1108_47# _022_ 4.8e-20
C14692 _326_/a_805_47# mask\[6\] 1.94e-21
C14693 net24 net15 0.00618f
C14694 _326_/a_761_289# _078_ 0.0108f
C14695 net34 _333_/a_1283_21# 0.00138f
C14696 _333_/a_448_47# _055_ 8.27e-22
C14697 net15 _014_ 0.0791f
C14698 net12 _325_/a_1108_47# 7.56e-21
C14699 _308_/a_1270_413# net23 5.16e-20
C14700 _308_/a_1217_47# net43 9.72e-19
C14701 _128_ clknet_2_3__leaf_clk 1.4e-20
C14702 net9 _334_/a_651_413# 4.52e-19
C14703 net13 _159_/a_27_47# 2.62e-19
C14704 _337_/a_448_47# _034_ 0.00166f
C14705 trim_val\[2\] _108_ 0.0396f
C14706 VPWR _324_/a_543_47# 0.0178f
C14707 clkbuf_2_2__f_clk/a_110_47# net11 2.35e-20
C14708 _322_/a_27_47# net53 2.38e-20
C14709 output23/a_27_47# result[1] 0.00859f
C14710 _110_ _269_/a_81_21# 0.00291f
C14711 _341_/a_27_47# _001_ 5.83e-20
C14712 _053_ _194_/a_199_47# 0.00139f
C14713 _309_/a_543_47# net43 0.00393f
C14714 _125_ net33 0.401f
C14715 _309_/a_27_47# net23 3.7e-20
C14716 _108_ _049_ 2.47e-20
C14717 _289_/a_68_297# cal_count\[0\] 4.41e-19
C14718 net22 _137_/a_68_297# 0.0166f
C14719 net4 _279_/a_396_47# 0.0117f
C14720 _042_ _247_/a_109_297# 0.0466f
C14721 _053_ _304_/a_543_47# 0.0172f
C14722 net31 _127_ 3.67e-20
C14723 VPWR _198_/a_109_47# -1.62e-19
C14724 _005_ _245_/a_109_297# 5e-20
C14725 net16 _332_/a_543_47# 0.00336f
C14726 _244_/a_27_297# _049_ 7.59e-19
C14727 net16 _108_ 0.253f
C14728 clkbuf_0_clk/a_110_47# _092_ 5e-20
C14729 _305_/a_193_47# _002_ 0.012f
C14730 VPWR _322_/a_761_289# 0.00958f
C14731 _329_/a_543_47# clknet_2_2__leaf_clk 2.28e-19
C14732 VPWR _331_/a_761_289# 0.0275f
C14733 _021_ _311_/a_27_47# 7.16e-21
C14734 _314_/a_27_47# _011_ 0.0339f
C14735 _314_/a_761_289# _086_ 1.62e-19
C14736 VPWR _257_/a_109_47# -9.67e-19
C14737 trim[0] net16 3.49e-20
C14738 _189_/a_27_47# _227_/a_209_311# 4.59e-21
C14739 _311_/a_1108_47# net26 0.0577f
C14740 _233_/a_27_297# _315_/a_761_289# 3.84e-19
C14741 _146_/a_68_297# _042_ 9.24e-19
C14742 net43 net28 0.434f
C14743 _309_/a_761_289# _101_ 1.29e-19
C14744 output20/a_27_47# _156_/a_27_47# 5.42e-20
C14745 _320_/a_193_47# _209_/a_27_47# 2.58e-19
C14746 _305_/a_639_47# clknet_2_1__leaf_clk 1.98e-20
C14747 _064_ _256_/a_27_297# 0.00741f
C14748 _324_/a_27_47# _312_/a_27_47# 1.9e-20
C14749 _331_/a_27_47# _331_/a_448_47# -0.00297f
C14750 net12 mask\[1\] 1.8e-20
C14751 VPWR _303_/a_1270_413# 7.05e-20
C14752 _000_ clknet_2_3__leaf_clk 0.0294f
C14753 _185_/a_68_297# _316_/a_27_47# 6.01e-22
C14754 _323_/a_805_47# net19 5.15e-19
C14755 _116_ _032_ 0.0668f
C14756 _219_/a_109_297# net53 8.05e-19
C14757 _327_/a_761_289# _136_ 9.25e-19
C14758 trim_val\[2\] _031_ 1.29e-19
C14759 _305_/a_27_47# _203_/a_59_75# 1.32e-21
C14760 _040_ _101_ 0.0781f
C14761 net9 _111_ 0.174f
C14762 net31 _126_ 0.00137f
C14763 _235_/a_79_21# _243_/a_27_297# 9.24e-21
C14764 _266_/a_68_297# cal_count\[3\] 8.9e-19
C14765 _023_ _007_ 2.04e-20
C14766 _308_/a_27_47# _080_ 1.26e-19
C14767 net33 net40 0.994f
C14768 cal_itt\[2\] _305_/a_193_47# 0.00164f
C14769 _329_/a_1108_47# trim_mask\[3\] 1.06e-19
C14770 output29/a_27_47# _224_/a_113_297# 1.79e-20
C14771 _058_ _172_/a_150_297# 5.6e-20
C14772 net16 _031_ 2.98e-19
C14773 net3 clknet_0_clk 8.51e-19
C14774 _078_ _310_/a_1283_21# 0.00703f
C14775 _104_ _302_/a_27_297# 4.46e-22
C14776 VPWR _309_/a_1217_47# 5.34e-19
C14777 _303_/a_193_47# _000_ -0.00347f
C14778 en_co_clk net55 0.0459f
C14779 net43 _159_/a_27_47# 0.00878f
C14780 _328_/a_805_47# net46 5.57e-19
C14781 net24 _310_/a_193_47# 2.6e-21
C14782 mask\[1\] net44 0.144f
C14783 VPWR _101_ 1.34f
C14784 _233_/a_27_297# net45 2.35e-19
C14785 _038_ _092_ 0.00838f
C14786 _292_/a_493_297# _128_ 6.9e-20
C14787 _104_ _106_ 0.00183f
C14788 net46 rebuffer3/a_75_212# 8.12e-20
C14789 net43 result[3] 6.6e-20
C14790 _169_/a_373_53# _051_ 0.00165f
C14791 net54 _051_ 0.00909f
C14792 clk input1/a_75_212# 5.57e-20
C14793 _015_ clk 0.0298f
C14794 _328_/a_1283_21# _113_ 0.0215f
C14795 _328_/a_543_47# _030_ 2.04e-20
C14796 _322_/a_1283_21# _101_ 1.38e-19
C14797 _322_/a_761_289# net52 3.59e-21
C14798 VPWR _297_/a_285_47# -0.00216f
C14799 _094_ state\[1\] 3.09e-22
C14800 clkbuf_2_2__f_clk/a_110_47# _279_/a_204_297# 6.65e-21
C14801 _053_ _302_/a_109_47# 0.00306f
C14802 _097_ _093_ 0.507f
C14803 _321_/a_1108_47# mask\[2\] 0.00121f
C14804 en_co_clk _067_ 0.0436f
C14805 en_co_clk _070_ 4.53e-21
C14806 net21 net20 0.00154f
C14807 _065_ net46 0.00145f
C14808 net8 _334_/a_543_47# 0.00525f
C14809 net21 net53 1.58e-20
C14810 _327_/a_805_47# trim_mask\[0\] 3.21e-21
C14811 _327_/a_651_413# _024_ 0.00219f
C14812 _015_ net4 0.0171f
C14813 _042_ _018_ 0.172f
C14814 _219_/a_109_297# _008_ 0.00121f
C14815 _295_/a_113_47# _131_ 1.4e-19
C14816 _230_/a_59_75# _062_ 0.00845f
C14817 net23 _101_ 0.0393f
C14818 _305_/a_1462_47# _002_ 7.49e-19
C14819 _000_ net53 0.00139f
C14820 mask\[6\] _250_/a_27_297# 0.0375f
C14821 net2 _126_ 0.0711f
C14822 net9 _135_ 4.07e-19
C14823 _312_/a_1283_21# net20 9.79e-19
C14824 VPWR _260_/a_250_297# 0.0125f
C14825 _078_ _311_/a_448_47# 1.55e-20
C14826 net13 _236_/a_109_297# 1.33e-19
C14827 _093_ _315_/a_543_47# 1.44e-19
C14828 _012_ _315_/a_193_47# 0.0449f
C14829 calibrate _315_/a_1283_21# 0.0316f
C14830 _337_/a_1283_21# _226_/a_27_47# 0.00132f
C14831 _322_/a_27_47# _019_ 0.0341f
C14832 _104_ trim_mask\[0\] 0.274f
C14833 _300_/a_47_47# cal_count\[2\] 8.29e-19
C14834 _331_/a_193_47# clknet_2_2__leaf_clk 0.00168f
C14835 _331_/a_27_47# _028_ 0.326f
C14836 _324_/a_1283_21# net19 0.00291f
C14837 clkbuf_2_3__f_clk/a_110_47# _279_/a_314_297# 2.66e-21
C14838 _257_/a_109_297# clknet_2_2__leaf_clk 2.86e-20
C14839 _280_/a_75_212# net19 1.78e-22
C14840 clkbuf_2_1__f_clk/a_110_47# mask\[0\] 3.73e-19
C14841 net48 trim_val\[1\] 9.98e-21
C14842 _317_/a_193_47# _317_/a_761_289# -0.00517f
C14843 _272_/a_81_21# trim_val\[2\] 0.0413f
C14844 net54 _316_/a_1283_21# 6.52e-20
C14845 _101_ net52 0.873f
C14846 net2 _072_ 0.234f
C14847 VPWR _312_/a_448_47# 1.22e-19
C14848 net15 _319_/a_805_47# 3.43e-19
C14849 _230_/a_59_75# _195_/a_76_199# 1.86e-19
C14850 _232_/a_220_297# _049_ 6.24e-19
C14851 _320_/a_543_47# mask\[1\] 0.0346f
C14852 _305_/a_1283_21# _072_ 0.0404f
C14853 _305_/a_1108_47# cal_itt\[3\] 4.63e-19
C14854 net42 _227_/a_209_311# 7.88e-20
C14855 clkbuf_2_0__f_clk/a_110_47# _078_ 1.16e-19
C14856 output31/a_27_47# net33 0.0052f
C14857 _321_/a_193_47# net15 0.0117f
C14858 _321_/a_543_47# _085_ 3.19e-20
C14859 _235_/a_297_47# net55 0.00705f
C14860 trim_mask\[3\] _280_/a_75_212# 6.83e-19
C14861 clknet_2_0__leaf_clk net51 0.0639f
C14862 fanout44/a_27_47# clknet_0_clk 1.96e-21
C14863 result[4] _023_ 5.22e-19
C14864 cal_itt\[2\] _305_/a_1462_47# 8.36e-19
C14865 _066_ _062_ 0.0114f
C14866 net16 net49 0.433f
C14867 _272_/a_81_21# net16 0.00258f
C14868 net15 _337_/a_193_47# 1.08e-20
C14869 _235_/a_79_21# _337_/a_193_47# 4.82e-19
C14870 _087_ _090_ 0.0429f
C14871 VPWR trim_val\[3\] 0.0499f
C14872 net35 net34 0.00132f
C14873 result[7] net29 0.00222f
C14874 _170_/a_299_297# _049_ 2.69e-19
C14875 _323_/a_761_289# mask\[4\] 0.00101f
C14876 fanout47/a_27_47# _068_ 3.24e-19
C14877 _239_/a_694_21# _049_ 0.00157f
C14878 _058_ _301_/a_285_47# 1.75e-19
C14879 _337_/a_805_47# en_co_clk 2.38e-19
C14880 _012_ _014_ 1.56e-20
C14881 mask\[6\] _009_ 4.05e-19
C14882 _303_/a_639_47# net19 0.00129f
C14883 _328_/a_543_47# trim_mask\[1\] 0.03f
C14884 _033_ _330_/a_1108_47# 5.66e-20
C14885 _336_/a_1283_21# net46 0.0406f
C14886 _336_/a_1108_47# _027_ 1.01e-21
C14887 cal _316_/a_448_47# 3.68e-20
C14888 _227_/a_209_311# _054_ 5.12e-20
C14889 _227_/a_368_53# _049_ 2.88e-19
C14890 VPWR _333_/a_1283_21# 0.014f
C14891 net9 _112_ 1.19e-20
C14892 en valid 0.00147f
C14893 _227_/a_209_311# net30 1.72e-20
C14894 _341_/a_448_47# _092_ 5.82e-21
C14895 _128_ _291_/a_35_297# 6.89e-19
C14896 _200_/a_209_297# cal_itt\[0\] 0.0294f
C14897 _200_/a_80_21# cal_itt\[1\] 0.00295f
C14898 _048_ _119_ 6.77e-19
C14899 _309_/a_27_47# _216_/a_113_297# 2.65e-20
C14900 _126_ _123_ 2.34e-21
C14901 _336_/a_448_47# _052_ 1.24e-20
C14902 _205_/a_27_47# rebuffer6/a_27_47# 2.19e-20
C14903 _023_ net27 2.27e-19
C14904 mask\[7\] result[5] 0.00214f
C14905 _284_/a_150_297# en_co_clk 8.78e-19
C14906 _107_ _229_/a_27_297# 7.58e-19
C14907 _263_/a_297_47# _090_ 1.29e-19
C14908 _083_ _101_ 0.0013f
C14909 net16 _289_/a_68_297# 5.02e-19
C14910 _168_/a_27_413# _227_/a_209_311# 6.04e-21
C14911 _168_/a_207_413# _227_/a_109_93# 2.38e-20
C14912 _325_/a_651_413# net13 5.88e-19
C14913 clk _330_/a_543_47# 1.65e-19
C14914 _053_ _041_ 2.62e-20
C14915 net43 _209_/a_27_47# 3.21e-20
C14916 _119_ trim_mask\[4\] 0.00837f
C14917 _304_/a_193_47# _124_ 5.74e-22
C14918 trim[2] _272_/a_299_297# 1.59e-19
C14919 output10/a_27_47# net10 0.0263f
C14920 _237_/a_76_199# _099_ 0.0546f
C14921 _237_/a_505_21# _095_ 0.00165f
C14922 _048_ _087_ 0.463f
C14923 _192_/a_174_21# _049_ 0.00495f
C14924 _042_ _078_ 0.0121f
C14925 _336_/a_1108_47# _335_/a_448_47# 3.67e-21
C14926 _322_/a_27_47# _205_/a_27_47# 0.0117f
C14927 output9/a_27_47# net9 0.0142f
C14928 _331_/a_1217_47# _028_ 1.84e-19
C14929 _331_/a_1462_47# clknet_2_2__leaf_clk 3.64e-20
C14930 _025_ clknet_2_2__leaf_clk 0.149f
C14931 clknet_2_2__leaf_clk _260_/a_93_21# 1.05e-20
C14932 _327_/a_193_47# clknet_2_3__leaf_clk 4.14e-19
C14933 calibrate _243_/a_373_47# 1.78e-19
C14934 net13 _248_/a_373_47# 5.63e-19
C14935 VPWR _325_/a_1283_21# 0.0366f
C14936 state\[0\] _316_/a_1270_413# 8.89e-21
C14937 net4 _330_/a_543_47# 3.94e-19
C14938 net48 _114_ 0.00155f
C14939 _059_ clone7/a_27_47# 0.00398f
C14940 _309_/a_193_47# mask\[1\] 9.34e-20
C14941 trim_mask\[0\] _267_/a_59_75# 0.0743f
C14942 clknet_2_1__leaf_clk net45 0.266f
C14943 net42 _168_/a_207_413# 2.09e-21
C14944 _048_ _266_/a_150_297# 5.59e-19
C14945 _336_/a_651_413# _108_ 3.38e-20
C14946 _325_/a_543_47# _159_/a_27_47# 1.05e-19
C14947 _058_ clknet_2_3__leaf_clk 6.52e-19
C14948 _064_ _329_/a_193_47# 5.56e-20
C14949 ctlp[1] result[7] 8.79e-20
C14950 _094_ _337_/a_1108_47# 0.004f
C14951 _010_ _222_/a_199_47# 1.01e-19
C14952 _214_/a_113_297# mask\[2\] 2.31e-19
C14953 _059_ net4 3.63e-20
C14954 mask\[4\] clknet_2_3__leaf_clk 1.27e-19
C14955 VPWR _248_/a_27_297# 0.0992f
C14956 _306_/a_1108_47# clk 0.00192f
C14957 VPWR _241_/a_297_47# -2.13e-19
C14958 clknet_2_1__leaf_clk _065_ 0.0218f
C14959 _121_ en_co_clk 0.00168f
C14960 _048_ _263_/a_297_47# 2.8e-19
C14961 net12 _306_/a_1283_21# 0.00158f
C14962 _110_ _103_ 4.07e-20
C14963 _325_/a_651_413# net43 0.00319f
C14964 _064_ net18 0.0288f
C14965 _320_/a_193_47# mask\[2\] 5.9e-19
C14966 cal _013_ 4.03e-19
C14967 _168_/a_207_413# _054_ 3.69e-20
C14968 _125_ output40/a_27_47# 0.0129f
C14969 _253_/a_81_21# _310_/a_27_47# 0.0015f
C14970 output32/a_27_47# _047_ 0.0241f
C14971 _107_ _260_/a_256_47# 2.35e-19
C14972 _192_/a_505_280# _192_/a_548_47# -2.14e-20
C14973 cal_itt\[1\] _071_ 4.59e-19
C14974 _322_/a_543_47# mask\[1\] 1.91e-19
C14975 _309_/a_543_47# _082_ 9.95e-19
C14976 _303_/a_193_47# mask\[4\] 2.28e-19
C14977 net12 _062_ 0.00931f
C14978 _333_/a_543_47# clknet_2_2__leaf_clk 4.83e-20
C14979 mask\[0\] net30 0.228f
C14980 clknet_2_1__leaf_clk _319_/a_27_47# 0.00309f
C14981 clkbuf_2_1__f_clk/a_110_47# _319_/a_448_47# 6.83e-19
C14982 _308_/a_761_289# fanout43/a_27_47# 0.00118f
C14983 _318_/a_193_47# clknet_2_0__leaf_clk 0.00367f
C14984 _325_/a_448_47# _101_ 2e-19
C14985 _306_/a_1283_21# net44 0.0633f
C14986 trim_mask\[0\] net37 0.00301f
C14987 _256_/a_109_47# _108_ 1.46e-20
C14988 _293_/a_384_47# cal_count\[0\] 7.39e-19
C14989 net20 _045_ 0.0131f
C14990 ctlp[2] net16 0.00419f
C14991 _326_/a_27_47# _023_ 0.0332f
C14992 _326_/a_193_47# _102_ 0.00182f
C14993 _326_/a_761_289# mask\[7\] 0.00354f
C14994 cal_itt\[2\] _262_/a_193_297# 2.71e-19
C14995 net43 _248_/a_373_47# 3.4e-20
C14996 _050_ _089_ 5.45e-21
C14997 _045_ net53 1.02e-19
C14998 _329_/a_193_47# _057_ 3.06e-19
C14999 trim_val\[3\] net50 0.0617f
C15000 _249_/a_109_297# net53 0.051f
C15001 _053_ net18 0.829f
C15002 _107_ net19 0.0393f
C15003 VPWR _190_/a_655_47# -9.49e-19
C15004 clkbuf_2_0__f_clk/a_110_47# _096_ 0.0044f
C15005 clknet_0_clk _330_/a_27_47# 5.66e-19
C15006 clkbuf_2_2__f_clk/a_110_47# _330_/a_1283_21# 0.0109f
C15007 ctlp[3] net17 0.00417f
C15008 _286_/a_76_199# _338_/a_27_47# 1.64e-19
C15009 _001_ net19 2.07e-19
C15010 _231_/a_161_47# _107_ 4.94e-19
C15011 net15 _316_/a_1108_47# 0.00642f
C15012 _022_ _078_ 2.81e-20
C15013 _305_/a_193_47# _067_ 6.85e-20
C15014 net22 mask\[0\] 0.17f
C15015 _305_/a_193_47# _070_ 2.92e-20
C15016 net31 _047_ 0.104f
C15017 _328_/a_1270_413# net9 1.5e-19
C15018 _336_/a_1108_47# _032_ 3.86e-21
C15019 net44 _062_ 5.01e-19
C15020 _020_ clknet_2_3__leaf_clk 0.00112f
C15021 VPWR _249_/a_373_47# -4.29e-19
C15022 _210_/a_113_297# net45 0.00159f
C15023 _340_/a_1602_47# _300_/a_47_47# 6.18e-20
C15024 _057_ net18 0.026f
C15025 VPWR trim_val\[4\] 0.102f
C15026 _026_ _327_/a_543_47# 4.33e-20
C15027 output40/a_27_47# net40 0.0513f
C15028 _306_/a_1108_47# _073_ 1.09e-19
C15029 _306_/a_1283_21# _003_ 1.29e-20
C15030 VPWR _327_/a_543_47# 0.0234f
C15031 _317_/a_1283_21# state\[1\] 0.00705f
C15032 _074_ _313_/a_193_47# 6.67e-19
C15033 clknet_0_clk _120_ 8.5e-19
C15034 cal_itt\[2\] _201_/a_113_47# 2.46e-19
C15035 _315_/a_27_47# _315_/a_1283_21# -9.15e-20
C15036 _315_/a_193_47# _315_/a_543_47# -8.58e-19
C15037 _270_/a_145_75# net16 4.09e-19
C15038 mask\[4\] net20 1.68e-22
C15039 net4 _195_/a_505_21# 7.28e-19
C15040 _322_/a_651_413# mask\[3\] 0.0227f
C15041 mask\[4\] net53 0.572f
C15042 _259_/a_27_297# _119_ 4.94e-19
C15043 _166_/a_161_47# _107_ 1.77e-19
C15044 _110_ _336_/a_1283_21# 0.00565f
C15045 VPWR net35 0.226f
C15046 _259_/a_373_47# VPWR -5.29e-19
C15047 _062_ _003_ 1.18e-20
C15048 _023_ _314_/a_448_47# 1.94e-20
C15049 _097_ _014_ 0.0205f
C15050 VPWR output11/a_27_47# 0.0473f
C15051 _249_/a_27_297# _312_/a_27_47# 3.88e-21
C15052 output36/a_27_47# net16 3.37e-19
C15053 _109_ _333_/a_27_47# 1.75e-20
C15054 _038_ net46 0.026f
C15055 result[3] _082_ 5.94e-19
C15056 _341_/a_1283_21# net40 1.69e-20
C15057 _320_/a_1283_21# _077_ 2.48e-19
C15058 _320_/a_1108_47# _076_ 0.00196f
C15059 _265_/a_384_47# trim_val\[0\] 3.13e-19
C15060 trim[1] trim_mask\[0\] 6.55e-19
C15061 _093_ fanout45/a_27_47# 2.06e-20
C15062 _322_/a_448_47# mask\[4\] 8.95e-19
C15063 _063_ _190_/a_655_47# 0.0228f
C15064 _258_/a_27_297# _335_/a_1108_47# 3.02e-20
C15065 _334_/a_543_47# net34 3.03e-21
C15066 net4 _335_/a_543_47# 3.88e-20
C15067 mask\[7\] _310_/a_1283_21# 0.00273f
C15068 en_co_clk clknet_2_3__leaf_clk 0.0129f
C15069 VPWR _281_/a_253_297# -5.04e-19
C15070 _149_/a_68_297# net26 0.00522f
C15071 net13 mask\[2\] 0.0636f
C15072 trim_mask\[1\] _336_/a_1270_413# 1.19e-20
C15073 _225_/a_109_297# _086_ 0.00114f
C15074 _192_/a_476_47# _065_ 7.4e-21
C15075 _090_ _099_ 0.07f
C15076 net45 _315_/a_761_289# 1.39e-20
C15077 clknet_2_0__leaf_clk _315_/a_1283_21# 0.00635f
C15078 _014_ _315_/a_543_47# 4.82e-21
C15079 VPWR _288_/a_59_75# 0.005f
C15080 _234_/a_109_297# clknet_2_0__leaf_clk 1.76e-21
C15081 _122_ _295_/a_113_47# 1.45e-19
C15082 _063_ trim_val\[4\] 6.93e-21
C15083 ctln[2] trim_val\[2\] 1.8e-20
C15084 net8 net48 0.0209f
C15085 _107_ _279_/a_27_47# 0.0022f
C15086 _321_/a_761_289# clknet_2_1__leaf_clk 0.00609f
C15087 _058_ _266_/a_68_297# 3.24e-19
C15088 trim_mask\[0\] _332_/a_651_413# 1.2e-19
C15089 _273_/a_59_75# _334_/a_448_47# 2.34e-19
C15090 _020_ net20 2.56e-22
C15091 _024_ _111_ 7.76e-21
C15092 _020_ net53 0.155f
C15093 _169_/a_215_311# _090_ 2.65e-21
C15094 net54 _087_ 9.32e-20
C15095 ctln[2] net16 1.33e-20
C15096 cal_count\[0\] _338_/a_27_47# 6.43e-21
C15097 _124_ _338_/a_652_21# 0.00466f
C15098 _008_ mask\[4\] 0.0966f
C15099 _242_/a_79_21# _092_ 3.06e-20
C15100 _324_/a_805_47# mask\[5\] 9.25e-20
C15101 _006_ _310_/a_543_47# 2.82e-20
C15102 fanout43/a_27_47# _245_/a_109_47# 5.73e-20
C15103 _305_/a_1462_47# _067_ 1.46e-21
C15104 _064_ _191_/a_27_297# 0.0426f
C15105 _002_ _202_/a_297_47# 0.00166f
C15106 _188_/a_27_47# _132_ 4.11e-22
C15107 _181_/a_68_297# _107_ 2.75e-20
C15108 net47 net2 0.0188f
C15109 _051_ net51 3.7e-20
C15110 _322_/a_193_47# mask\[2\] 0.0128f
C15111 trim_mask\[2\] net46 0.249f
C15112 net24 result[2] 0.0148f
C15113 net34 _332_/a_27_47# 2.82e-21
C15114 _079_ mask\[0\] 0.0294f
C15115 net9 _304_/a_27_47# 0.00441f
C15116 cal_itt\[0\] _197_/a_199_47# 0.00176f
C15117 cal_itt\[1\] _197_/a_113_297# 0.00166f
C15118 VPWR _156_/a_27_47# 0.0829f
C15119 input2/a_27_47# _297_/a_285_47# 7.66e-20
C15120 trim_mask\[4\] _279_/a_206_47# 0.00114f
C15121 _301_/a_47_47# _332_/a_193_47# 9.75e-21
C15122 net27 result[6] 9.45e-21
C15123 _327_/a_761_289# clknet_2_2__leaf_clk 5.58e-19
C15124 _319_/a_1270_413# _049_ 3.27e-20
C15125 _324_/a_1270_413# net27 1.8e-20
C15126 _319_/a_448_47# net30 5.56e-19
C15127 _047_ trim_val\[1\] 0.00257f
C15128 _253_/a_81_21# clknet_2_1__leaf_clk 6.49e-21
C15129 _060_ _263_/a_382_297# 2.06e-19
C15130 net12 net2 0.00487f
C15131 _305_/a_1108_47# clk 0.00238f
C15132 VPWR _330_/a_193_47# 0.0224f
C15133 _329_/a_193_47# _027_ 0.00194f
C15134 trim[2] net33 0.0962f
C15135 _329_/a_27_47# net46 0.0117f
C15136 _339_/a_27_47# _286_/a_505_21# 0.033f
C15137 _339_/a_193_47# _286_/a_76_199# 4.61e-20
C15138 _048_ _099_ 0.0926f
C15139 net43 mask\[2\] 8.01e-19
C15140 _312_/a_805_47# _045_ 5.01e-20
C15141 net55 _049_ 0.0429f
C15142 _275_/a_81_21# _178_/a_68_297# 0.00128f
C15143 cal_itt\[2\] _202_/a_297_47# 0.00712f
C15144 net45 _065_ 6.92e-19
C15145 _323_/a_193_47# _068_ 2.08e-22
C15146 _065_ rebuffer3/a_75_212# 9.5e-22
C15147 net17 cal_count\[0\] 9.79e-21
C15148 net19 _118_ 3.87e-20
C15149 _313_/a_543_47# net29 1.85e-22
C15150 _259_/a_109_47# clknet_2_2__leaf_clk 3.13e-21
C15151 cal_itt\[1\] _304_/a_543_47# 1.58e-19
C15152 _200_/a_80_21# _106_ 1.09e-20
C15153 _189_/a_408_47# clk 0.00194f
C15154 _321_/a_448_47# _018_ 0.00199f
C15155 _101_ _208_/a_76_199# 0.00106f
C15156 _231_/a_161_47# _118_ 3.89e-19
C15157 _019_ mask\[4\] 0.00507f
C15158 net33 _132_ 0.00629f
C15159 _030_ _055_ 1.99e-20
C15160 _008_ _020_ 3.4e-20
C15161 _027_ net18 1.1e-19
C15162 _104_ _089_ 0.00112f
C15163 _181_/a_68_297# _279_/a_27_47# 0.0158f
C15164 _341_/a_448_47# net46 1.27e-21
C15165 net50 trim_val\[4\] 7.69e-20
C15166 mask\[0\] _319_/a_1108_47# 0.0378f
C15167 state\[2\] _242_/a_79_21# 0.00202f
C15168 clkbuf_2_2__f_clk/a_110_47# _108_ 7.12e-19
C15169 _305_/a_1108_47# net4 2.22e-21
C15170 _040_ _077_ 8.91e-20
C15171 _115_ net46 0.241f
C15172 net2 net44 0.00953f
C15173 _319_/a_761_289# clknet_2_0__leaf_clk 0.0526f
C15174 _319_/a_27_47# net45 3.7e-19
C15175 _321_/a_639_47# _042_ 3.04e-19
C15176 _307_/a_1283_21# _137_/a_68_297# 0.0135f
C15177 _325_/a_1108_47# _248_/a_109_297# 5.3e-21
C15178 _286_/a_76_199# clknet_2_3__leaf_clk 0.00387f
C15179 net44 _311_/a_1270_413# 1.35e-19
C15180 _293_/a_384_47# net16 2.61e-19
C15181 _306_/a_651_413# rebuffer6/a_27_47# 6.28e-21
C15182 net27 _312_/a_27_47# 2.34e-19
C15183 _107_ _118_ 0.0151f
C15184 _233_/a_27_297# _013_ 2.65e-19
C15185 net47 _123_ 0.192f
C15186 _273_/a_59_75# _031_ 0.00952f
C15187 _264_/a_27_297# net30 0.0977f
C15188 _189_/a_218_47# net44 2.22e-22
C15189 VPWR _077_ 0.0865f
C15190 _340_/a_1140_413# _123_ 0.00163f
C15191 _053_ _090_ 2.67e-20
C15192 VPWR _306_/a_543_47# 0.0247f
C15193 _319_/a_27_47# _065_ 2.03e-19
C15194 _312_/a_543_47# _084_ 1.05e-19
C15195 _301_/a_47_47# net2 0.00226f
C15196 cal_itt\[0\] _091_ 0.134f
C15197 _322_/a_1283_21# _077_ 4.15e-20
C15198 _326_/a_543_47# net14 0.00717f
C15199 net2 _003_ 4.96e-20
C15200 _200_/a_80_21# trim_mask\[0\] 1.5e-19
C15201 clknet_0_clk _068_ 0.0251f
C15202 _241_/a_105_352# _095_ 0.0394f
C15203 _341_/a_27_47# net2 1.15e-20
C15204 _293_/a_81_21# _126_ 9.24e-20
C15205 _058_ _333_/a_1270_413# 3.76e-21
C15206 net2 _299_/a_215_297# 0.0259f
C15207 _061_ _301_/a_285_47# 2.07e-19
C15208 _308_/a_193_47# _039_ 4.38e-19
C15209 net13 _094_ 0.0763f
C15210 _102_ _251_/a_27_297# 0.00446f
C15211 mask\[7\] _251_/a_109_297# 5.7e-19
C15212 _050_ _092_ 0.882f
C15213 trim_mask\[2\] _269_/a_81_21# 1.32e-20
C15214 net9 _340_/a_476_47# 0.0153f
C15215 net4 trim_mask\[1\] 2.12e-21
C15216 _307_/a_761_289# _074_ 0.00439f
C15217 _064_ _048_ 7.4e-21
C15218 _304_/a_193_47# cal_count\[2\] 1.23e-21
C15219 output36/a_27_47# trimb[0] 0.0113f
C15220 trimb[1] cal_count\[0\] 4.96e-19
C15221 en_co_clk _263_/a_382_297# 1.73e-19
C15222 _326_/a_761_289# net28 9.18e-19
C15223 output19/a_27_47# net19 0.0144f
C15224 _325_/a_27_47# mask\[5\] 2.2e-21
C15225 net43 _306_/a_448_47# 5.43e-21
C15226 _279_/a_27_47# _118_ 0.0491f
C15227 _329_/a_1217_47# net46 9.36e-20
C15228 VPWR _330_/a_1462_47# 0.00178f
C15229 _339_/a_193_47# cal_count\[0\] 0.498f
C15230 _169_/a_109_53# _050_ 3.88e-20
C15231 _144_/a_27_47# _126_ 6.56e-22
C15232 net43 _314_/a_193_47# 0.0124f
C15233 _304_/a_761_289# _065_ 0.00475f
C15234 _337_/a_805_47# _049_ 3.28e-19
C15235 _317_/a_193_47# _316_/a_193_47# 9.38e-21
C15236 clk _317_/a_543_47# 0.00437f
C15237 _317_/a_27_47# _316_/a_761_289# 0.00112f
C15238 _064_ trim_mask\[4\] 0.18f
C15239 clknet_2_2__leaf_clk _330_/a_27_47# 0.28f
C15240 trim_mask\[1\] _055_ 0.00202f
C15241 VPWR _326_/a_543_47# 0.0155f
C15242 mask\[4\] _205_/a_27_47# 1.07e-21
C15243 net52 _077_ 5.79e-19
C15244 _051_ _318_/a_193_47# 2.52e-19
C15245 _329_/a_543_47# _031_ 1.22e-19
C15246 VPWR _334_/a_543_47# 0.0295f
C15247 _181_/a_150_297# trim_val\[4\] 8.47e-19
C15248 _053_ _048_ 0.0572f
C15249 _181_/a_68_297# _118_ 0.0224f
C15250 _106_ _262_/a_27_47# 0.00426f
C15251 _328_/a_27_47# trim_mask\[0\] 1.21e-20
C15252 clkbuf_2_0__f_clk/a_110_47# clknet_0_clk 0.0393f
C15253 cal_count\[0\] trimb[4] 5.67e-20
C15254 _307_/a_651_413# _039_ 6.5e-19
C15255 VPWR _286_/a_218_374# 2.66e-19
C15256 cal_count\[0\] clknet_2_3__leaf_clk 0.36f
C15257 _330_/a_27_47# net11 1.44e-20
C15258 _330_/a_761_289# net19 0.00452f
C15259 net4 _317_/a_543_47# 3.81e-19
C15260 _308_/a_651_413# _074_ 0.00538f
C15261 _303_/a_27_47# _068_ 0.00323f
C15262 _273_/a_59_75# _272_/a_81_21# 0.00979f
C15263 _335_/a_761_289# _280_/a_75_212# 1.36e-21
C15264 _078_ _313_/a_761_289# 6.56e-20
C15265 state\[1\] net55 0.0176f
C15266 _053_ trim_mask\[4\] 0.0186f
C15267 net14 _310_/a_1108_47# 4.01e-19
C15268 _089_ _228_/a_79_21# 0.00733f
C15269 net5 clkc 0.0661f
C15270 _337_/a_761_289# net45 4.08e-19
C15271 VPWR _335_/a_193_47# 0.0602f
C15272 _110_ trim_mask\[2\] 0.515f
C15273 result[6] _314_/a_448_47# 9.22e-19
C15274 state\[2\] _050_ 0.711f
C15275 _309_/a_651_413# _310_/a_27_47# 6.14e-21
C15276 _309_/a_543_47# _310_/a_1283_21# 9.43e-19
C15277 _237_/a_76_199# _093_ 4.41e-19
C15278 _237_/a_505_21# calibrate 5.7e-20
C15279 net43 _094_ 2.06e-20
C15280 trim_mask\[3\] _330_/a_761_289# 8.58e-21
C15281 _323_/a_193_47# _042_ 0.545f
C15282 _067_ _201_/a_113_47# 2.18e-20
C15283 _070_ _201_/a_113_47# 3.03e-20
C15284 _326_/a_448_47# net43 1.1e-20
C15285 _134_ _135_ 0.0234f
C15286 _257_/a_27_297# _335_/a_1108_47# 4.52e-21
C15287 _257_/a_109_297# _335_/a_1283_21# 8.88e-21
C15288 _323_/a_1108_47# clknet_2_1__leaf_clk 6.95e-20
C15289 _061_ clknet_2_3__leaf_clk 0.00543f
C15290 VPWR _187_/a_27_413# 0.0233f
C15291 net13 _074_ 0.13f
C15292 VPWR _314_/a_639_47# 4.68e-19
C15293 _302_/a_109_297# rebuffer3/a_75_212# 1.6e-19
C15294 _032_ net18 4.23e-19
C15295 VPWR _332_/a_27_47# 0.0703f
C15296 clk _318_/a_448_47# 0.0164f
C15297 mask\[5\] _152_/a_150_297# 9.54e-19
C15298 _111_ cal_count\[3\] 0.00281f
C15299 _337_/a_761_289# _065_ 8.96e-21
C15300 _233_/a_373_47# valid 1.33e-19
C15301 _143_/a_68_297# _078_ 0.0426f
C15302 _048_ _226_/a_109_47# 0.00218f
C15303 _110_ _329_/a_27_47# 1.2e-19
C15304 VPWR _268_/a_75_212# 0.0661f
C15305 trim_mask\[0\] _262_/a_27_47# 0.00833f
C15306 net12 _318_/a_1108_47# 0.00278f
C15307 _083_ _077_ 5.66e-20
C15308 net9 _338_/a_193_47# 5.19e-20
C15309 _326_/a_543_47# net52 1.38e-19
C15310 _326_/a_1108_47# _101_ 6.61e-20
C15311 mask\[7\] _022_ 0.00102f
C15312 result[1] _308_/a_193_47# 0.00876f
C15313 net9 _340_/a_1224_47# 1.72e-20
C15314 _106_ wire42/a_75_212# 1.27e-20
C15315 net54 _099_ 0.0742f
C15316 _060_ _095_ 3.3e-20
C15317 _168_/a_297_47# clk 7.46e-19
C15318 VPWR _310_/a_1108_47# -4.61e-19
C15319 _302_/a_109_297# _065_ 3.33e-21
C15320 _340_/a_1182_261# cal_count\[2\] 0.00355f
C15321 net4 _318_/a_448_47# 1.7e-19
C15322 net17 net16 0.00167f
C15323 net47 _150_/a_27_47# 6.57e-19
C15324 _110_ _115_ 0.00236f
C15325 _121_ _049_ 0.0172f
C15326 _322_/a_193_47# _074_ 0.0117f
C15327 calibrate _331_/a_27_47# 6.64e-20
C15328 _329_/a_1283_21# trim_mask\[1\] 1.09e-19
C15329 _169_/a_215_311# net54 6.47e-20
C15330 _209_/a_27_47# _076_ 0.00552f
C15331 clknet_2_2__leaf_clk _330_/a_1217_47# 4.62e-19
C15332 net43 _244_/a_27_297# 0.00135f
C15333 _062_ net19 0.248f
C15334 _081_ net22 3.65e-20
C15335 _127_ net34 1.73e-19
C15336 _104_ _279_/a_490_47# 0.00142f
C15337 _231_/a_161_47# _062_ 7.77e-21
C15338 _327_/a_651_413# _058_ 0.00331f
C15339 net10 ctln[4] 0.00363f
C15340 _064_ _327_/a_27_47# 4.55e-19
C15341 _197_/a_199_47# _069_ 3.8e-19
C15342 _334_/a_761_289# clknet_2_2__leaf_clk 5.11e-19
C15343 _097_ _316_/a_1108_47# 9.37e-19
C15344 _088_ _260_/a_93_21# 2.44e-19
C15345 net43 _310_/a_1270_413# -9.71e-20
C15346 _311_/a_1108_47# net53 0.00102f
C15347 clkbuf_0_clk/a_110_47# _065_ 1.79e-20
C15348 net43 _074_ 0.0393f
C15349 _274_/a_75_212# _114_ 0.00163f
C15350 mask\[0\] net44 2.97e-19
C15351 trim_mask\[0\] wire42/a_75_212# 4.51e-19
C15352 _135_ cal_count\[3\] 0.00152f
C15353 clkbuf_2_1__f_clk/a_110_47# _040_ 0.00524f
C15354 _301_/a_285_47# net16 0.00322f
C15355 _259_/a_27_297# _064_ 0.0117f
C15356 _249_/a_27_297# _084_ 1.18e-20
C15357 _195_/a_76_199# net19 7.11e-20
C15358 VPWR _335_/a_1462_47# 7.25e-20
C15359 VPWR _305_/a_543_47# 0.018f
C15360 _107_ _062_ 0.0161f
C15361 net33 net32 1.61e-19
C15362 VPWR _311_/a_651_413# -0.00888f
C15363 state\[2\] _169_/a_301_53# 1.57e-21
C15364 output10/a_27_47# _335_/a_1283_21# 1.15e-19
C15365 _327_/a_27_47# _053_ 7.36e-20
C15366 _104_ _092_ 1.49e-20
C15367 net52 _310_/a_1108_47# 9.14e-20
C15368 _126_ net34 0.00327f
C15369 _335_/a_27_47# clknet_2_2__leaf_clk 0.0137f
C15370 VPWR _189_/a_27_47# 0.0542f
C15371 VPWR clkbuf_2_1__f_clk/a_110_47# 0.0195f
C15372 mask\[7\] _011_ 2.81e-19
C15373 _282_/a_68_297# _065_ 0.0229f
C15374 VPWR _332_/a_1217_47# 1.35e-19
C15375 _052_ _242_/a_297_47# 0.00254f
C15376 _304_/a_543_47# _302_/a_27_297# 8.26e-20
C15377 net13 _232_/a_220_297# 9.18e-19
C15378 _202_/a_297_47# _070_ 5.36e-19
C15379 _276_/a_59_75# VPWR 0.0304f
C15380 _333_/a_27_47# net46 0.369f
C15381 _304_/a_1108_47# _067_ 0.0051f
C15382 net24 _041_ 0.00654f
C15383 net9 _341_/a_1283_21# 0.0146f
C15384 _336_/a_1108_47# _106_ 3.75e-20
C15385 en_co_clk _095_ 0.575f
C15386 _339_/a_956_413# _123_ 0.00243f
C15387 _320_/a_1283_21# net30 4.43e-21
C15388 trimb[1] net16 4.04e-20
C15389 cal_itt\[0\] clkbuf_2_3__f_clk/a_110_47# 0.00811f
C15390 _267_/a_59_75# _109_ 0.0177f
C15391 net43 _305_/a_448_47# 0.0145f
C15392 net16 _339_/a_193_47# 1.92e-21
C15393 _214_/a_199_47# _078_ 2.65e-19
C15394 _038_ _065_ 0.243f
C15395 net43 _146_/a_150_297# 3.43e-19
C15396 _132_ output40/a_27_47# 7.25e-21
C15397 _321_/a_193_47# _321_/a_543_47# -0.0102f
C15398 _321_/a_27_47# _321_/a_1283_21# -9.15e-20
C15399 _319_/a_27_47# _282_/a_68_297# 7.58e-19
C15400 cal net1 0.0202f
C15401 net50 _335_/a_193_47# 0.00563f
C15402 trim_mask\[3\] _335_/a_761_289# 5.63e-20
C15403 trim_val\[3\] _335_/a_543_47# 1.48e-20
C15404 _220_/a_113_297# _084_ 0.00716f
C15405 _247_/a_109_297# _101_ 0.00262f
C15406 _065_ _204_/a_75_212# 1.15e-19
C15407 _008_ _311_/a_1108_47# 1.09e-19
C15408 net23 clkbuf_2_1__f_clk/a_110_47# 0.00115f
C15409 _317_/a_193_47# net14 5.64e-19
C15410 calibrate _331_/a_1217_47# 6.96e-20
C15411 _338_/a_476_47# _065_ 4.08e-20
C15412 net5 _136_ 5.3e-20
C15413 _014_ _316_/a_651_413# 0.00325f
C15414 net45 _316_/a_448_47# 5.09e-19
C15415 cal_itt\[1\] net18 2.96e-20
C15416 _053_ net54 1.84e-19
C15417 state\[0\] _060_ 0.0789f
C15418 _094_ net3 0.0127f
C15419 clk _336_/a_27_47# 2.69e-21
C15420 trim_mask\[4\] _027_ 2.73e-19
C15421 fanout47/a_27_47# net4 0.0201f
C15422 _320_/a_761_289# _078_ 1.24e-19
C15423 _320_/a_543_47# mask\[0\] 1.57e-20
C15424 _305_/a_543_47# _063_ 1.33e-20
C15425 _337_/a_27_47# _337_/a_1283_21# -9.15e-20
C15426 _307_/a_1108_47# net30 1.86e-19
C15427 _093_ _090_ 0.0849f
C15428 net13 net26 0.0114f
C15429 net9 _339_/a_652_21# 0.0048f
C15430 _320_/a_27_47# clknet_2_0__leaf_clk 0.03f
C15431 _257_/a_109_47# trim_mask\[1\] 8.34e-19
C15432 _104_ state\[2\] 0.0326f
C15433 _256_/a_27_297# _302_/a_27_297# 3.29e-21
C15434 net16 trimb[4] 3e-20
C15435 cal_count\[1\] net2 0.742f
C15436 net16 clknet_2_3__leaf_clk 0.016f
C15437 _181_/a_68_297# _062_ 3.02e-20
C15438 clkbuf_2_1__f_clk/a_110_47# net52 0.241f
C15439 _291_/a_35_297# cal_count\[0\] 0.0397f
C15440 clknet_0_clk cal_itt\[3\] 0.0237f
C15441 trim_mask\[0\] _336_/a_1108_47# 5.1e-20
C15442 _317_/a_193_47# net41 6.96e-21
C15443 net4 _336_/a_27_47# 0.00723f
C15444 _324_/a_27_47# mask\[6\] 4.25e-20
C15445 _333_/a_761_289# rebuffer2/a_75_212# 7.71e-20
C15446 VPWR _227_/a_109_93# 9.72e-19
C15447 _333_/a_651_413# rebuffer1/a_75_212# 4.98e-20
C15448 _333_/a_193_47# _332_/a_1108_47# 1.42e-21
C15449 _333_/a_543_47# _108_ 0.0112f
C15450 calibrate _242_/a_297_47# 0.00166f
C15451 _307_/a_1283_21# mask\[0\] 0.00278f
C15452 _307_/a_1108_47# net22 0.0591f
C15453 _307_/a_543_47# _078_ 3.81e-19
C15454 _259_/a_109_297# _330_/a_1108_47# 1.52e-19
C15455 VPWR _251_/a_109_47# -6.1e-19
C15456 _109_ net37 7.01e-21
C15457 _328_/a_1108_47# _329_/a_1108_47# 4.15e-21
C15458 net31 _333_/a_1108_47# 0.00298f
C15459 _265_/a_384_47# _108_ 1.18e-19
C15460 _178_/a_68_297# _057_ 9.24e-19
C15461 result[0] net22 0.0019f
C15462 _051_ _336_/a_448_47# 8.21e-21
C15463 _307_/a_193_47# clknet_2_0__leaf_clk 0.00726f
C15464 _324_/a_805_47# clknet_2_1__leaf_clk 1.32e-19
C15465 _329_/a_639_47# net9 7.53e-19
C15466 trim[3] _334_/a_27_47# 4.94e-20
C15467 clknet_0_clk _262_/a_205_47# 1.91e-20
C15468 VPWR _317_/a_193_47# -0.294f
C15469 _060_ _226_/a_27_47# 0.02f
C15470 _322_/a_193_47# net26 2.09e-20
C15471 _298_/a_78_199# cal_count\[2\] 0.0133f
C15472 result[7] net14 0.0254f
C15473 _235_/a_79_21# _092_ 0.0527f
C15474 net15 _092_ 0.167f
C15475 _304_/a_761_289# _038_ 0.00102f
C15476 _304_/a_448_47# _136_ 4.81e-19
C15477 trimb[3] net34 0.00164f
C15478 net14 net30 0.0107f
C15479 _333_/a_1217_47# net46 2.11e-20
C15480 _293_/a_81_21# net47 1.83e-20
C15481 _096_ clone7/a_27_47# 0.00608f
C15482 net12 _100_ 0.0959f
C15483 net2 net19 0.00927f
C15484 _303_/a_651_413# net26 1.01e-19
C15485 ctlp[7] _313_/a_1283_21# 0.00107f
C15486 clknet_2_1__leaf_clk _046_ 0.0278f
C15487 net27 _084_ 0.0275f
C15488 _332_/a_805_47# clknet_2_2__leaf_clk 2.34e-19
C15489 VPWR net42 0.482f
C15490 _051_ _206_/a_206_47# 5.53e-21
C15491 cal_itt\[0\] cal_count\[3\] 8.11e-20
C15492 _269_/a_81_21# _333_/a_27_47# 0.00145f
C15493 net4 _287_/a_75_212# 1.58e-19
C15494 _304_/a_1270_413# net47 2.4e-19
C15495 _048_ _093_ 0.153f
C15496 net43 _002_ 0.311f
C15497 _030_ _333_/a_1283_21# 4.61e-20
C15498 _113_ _333_/a_1108_47# 3.38e-21
C15499 _340_/a_27_47# net47 0.00376f
C15500 _256_/a_27_297# trim_mask\[0\] 0.0931f
C15501 _315_/a_27_47# output41/a_27_47# 3.29e-20
C15502 net13 _318_/a_651_413# 0.00247f
C15503 net43 net26 0.0143f
C15504 _074_ net3 3.09e-20
C15505 _308_/a_1270_413# _078_ 1.46e-19
C15506 _074_ _080_ 0.176f
C15507 net50 _335_/a_1462_47# 1.92e-19
C15508 clknet_2_1__leaf_clk _312_/a_761_289# 4.98e-19
C15509 _094_ fanout44/a_27_47# 5.81e-20
C15510 _308_/a_1108_47# net24 3.38e-21
C15511 net4 _096_ 3.61e-21
C15512 net22 net14 0.467f
C15513 _308_/a_1283_21# net45 0.0158f
C15514 _078_ _138_/a_27_47# 0.0117f
C15515 _308_/a_448_47# clknet_2_0__leaf_clk 0.00154f
C15516 _040_ net30 1.71e-20
C15517 _018_ _101_ 0.0497f
C15518 _299_/a_382_47# _131_ 0.00298f
C15519 trim_mask\[0\] _162_/a_27_47# 0.00115f
C15520 cal_count\[1\] _123_ 0.0248f
C15521 _062_ _118_ 0.0733f
C15522 state\[0\] en_co_clk 0.00123f
C15523 _341_/a_448_47# _065_ 0.00802f
C15524 net45 _013_ 0.0718f
C15525 VPWR net48 0.252f
C15526 _309_/a_27_47# _078_ 0.0158f
C15527 _292_/a_493_297# net16 6.13e-20
C15528 net47 _144_/a_27_47# 4.17e-20
C15529 output37/a_27_47# net33 0.0101f
C15530 _337_/a_193_47# _282_/a_150_297# 1.24e-19
C15531 _188_/a_27_47# _134_ 3.59e-21
C15532 _237_/a_505_21# clknet_2_0__leaf_clk 7.15e-20
C15533 _237_/a_76_199# _014_ 7.24e-19
C15534 _313_/a_193_47# _313_/a_448_47# -0.00297f
C15535 net2 _001_ 0.148f
C15536 VPWR _127_ 0.0569f
C15537 output20/a_27_47# net44 0.00394f
C15538 cal_itt\[0\] _303_/a_448_47# 7.63e-20
C15539 cal_itt\[1\] _303_/a_1108_47# 1.16e-20
C15540 _336_/a_193_47# clkbuf_2_2__f_clk/a_110_47# 0.0151f
C15541 VPWR result[7] 0.472f
C15542 net9 _339_/a_1056_47# 2.24e-19
C15543 net15 _246_/a_109_297# 0.00523f
C15544 _320_/a_1217_47# clknet_2_0__leaf_clk 1.2e-21
C15545 _051_ _337_/a_1283_21# 7.17e-19
C15546 VPWR _054_ 0.0917f
C15547 _216_/a_113_297# _310_/a_1108_47# 0.00151f
C15548 net25 _310_/a_27_47# 0.00129f
C15549 trim[1] _109_ 6.11e-20
C15550 VPWR _318_/a_1283_21# 0.0596f
C15551 _287_/a_75_212# _122_ 8.88e-21
C15552 VPWR net30 3.93f
C15553 _116_ _275_/a_299_297# 5.83e-20
C15554 _110_ _275_/a_384_47# 7.91e-21
C15555 _276_/a_59_75# net50 4.67e-19
C15556 _117_ _275_/a_81_21# 0.014f
C15557 en_co_clk _207_/a_109_297# 0.00235f
C15558 cal_itt\[2\] net43 0.00762f
C15559 _189_/a_218_47# _107_ 6.77e-19
C15560 net28 _022_ 8.53e-19
C15561 _035_ _338_/a_652_21# 1.2e-19
C15562 output15/a_27_47# _046_ 0.00266f
C15563 _064_ net40 0.347f
C15564 trim_mask\[2\] _336_/a_1283_21# 0.00755f
C15565 _188_/a_27_47# _130_ 5.13e-22
C15566 _341_/a_193_47# _230_/a_59_75# 6.55e-21
C15567 clknet_2_0__leaf_clk output41/a_27_47# 1.81e-20
C15568 _312_/a_193_47# _009_ 0.0158f
C15569 _173_/a_27_47# _055_ 0.0152f
C15570 VPWR _168_/a_27_413# 0.0431f
C15571 state\[2\] _228_/a_79_21# 2.59e-20
C15572 output23/a_27_47# _080_ 0.00498f
C15573 _320_/a_639_47# _065_ 2.56e-20
C15574 _259_/a_27_297# _027_ 0.0104f
C15575 _104_ _330_/a_651_413# 6.03e-20
C15576 _110_ _333_/a_27_47# 6.35e-19
C15577 _328_/a_1283_21# VPWR 0.00714f
C15578 net42 _063_ 0.00632f
C15579 _208_/a_76_199# _077_ 0.0271f
C15580 _330_/a_193_47# _330_/a_543_47# -0.0102f
C15581 _208_/a_505_21# _076_ 0.0564f
C15582 VPWR net22 0.457f
C15583 _051_ _033_ 4.8e-20
C15584 calibrate _241_/a_105_352# 9.55e-20
C15585 ctlp[2] net39 0.0015f
C15586 _168_/a_207_413# _331_/a_543_47# 3.65e-21
C15587 VPWR _126_ 0.447f
C15588 _308_/a_1283_21# _319_/a_27_47# 2.4e-19
C15589 _302_/a_109_297# _038_ 1.67e-20
C15590 VPWR _317_/a_1462_47# 7.03e-20
C15591 _306_/a_761_289# _208_/a_505_21# 8.62e-21
C15592 _307_/a_543_47# _004_ 0.00153f
C15593 net55 _240_/a_109_297# 0.00361f
C15594 en_co_clk _226_/a_27_47# 0.00555f
C15595 _315_/a_651_413# net14 0.00176f
C15596 trim_val\[3\] trim_mask\[1\] 1.05e-21
C15597 _322_/a_761_289# _078_ 3.39e-21
C15598 _053_ net40 0.00149f
C15599 fanout44/a_27_47# _244_/a_27_297# 2.31e-19
C15600 _134_ net33 3.12e-20
C15601 net27 _085_ 0.0174f
C15602 _319_/a_1283_21# clknet_0_clk 0.0256f
C15603 _232_/a_32_297# _107_ 6.74e-19
C15604 _249_/a_27_297# _311_/a_193_47# 3.43e-19
C15605 _222_/a_113_297# _085_ 0.00622f
C15606 trimb[0] trimb[1] 0.0464f
C15607 VPWR _072_ 0.717f
C15608 _304_/a_639_47# _122_ 0.00166f
C15609 _341_/a_193_47# _066_ 1.06e-20
C15610 clkbuf_2_2__f_clk/a_110_47# net55 3.7e-19
C15611 _239_/a_474_297# _242_/a_79_21# 1.54e-19
C15612 _021_ _312_/a_27_47# 3.92e-20
C15613 _112_ _333_/a_761_289# 4.82e-19
C15614 net49 _333_/a_543_47# 0.00704f
C15615 trim_val\[1\] _333_/a_1108_47# 0.0199f
C15616 _340_/a_193_47# _122_ 0.00197f
C15617 _272_/a_299_297# _333_/a_761_289# 9.29e-21
C15618 net33 _130_ 0.00557f
C15619 _304_/a_193_47# net18 0.0092f
C15620 _341_/a_448_47# _304_/a_761_289# 1.91e-20
C15621 _263_/a_382_297# _049_ 2.17e-20
C15622 net52 net30 1.74e-20
C15623 _315_/a_1108_47# valid 5.38e-19
C15624 _340_/a_1182_261# _041_ 4.68e-21
C15625 _340_/a_586_47# net47 1.54e-19
C15626 _063_ net30 0.0247f
C15627 _325_/a_27_47# clknet_2_1__leaf_clk 0.0192f
C15628 net23 net22 0.00148f
C15629 _123_ _001_ 0.0103f
C15630 input4/a_27_47# rstn 0.0134f
C15631 _340_/a_193_47# _037_ 0.0228f
C15632 _327_/a_761_289# _108_ 2.33e-19
C15633 _005_ clknet_2_0__leaf_clk 0.00317f
C15634 VPWR _262_/a_465_47# -2e-19
C15635 _327_/a_193_47# _111_ 1.95e-19
C15636 _309_/a_1217_47# _078_ 0.0011f
C15637 _309_/a_1462_47# mask\[0\] 2.34e-20
C15638 fanout45/a_27_47# _316_/a_1108_47# 0.00133f
C15639 mask\[4\] _311_/a_27_47# 0.228f
C15640 _107_ _227_/a_209_311# 0.00952f
C15641 _090_ _192_/a_505_280# 0.00181f
C15642 _323_/a_1108_47# _043_ 0.00275f
C15643 mask\[1\] _247_/a_27_297# 4.05e-20
C15644 _079_ net14 0.0167f
C15645 VPWR _315_/a_651_413# -0.00431f
C15646 _058_ rebuffer2/a_75_212# 0.005f
C15647 _303_/a_1283_21# _065_ 2.22e-20
C15648 _309_/a_1270_413# net24 4.39e-19
C15649 _337_/a_1270_413# net44 5.33e-20
C15650 _149_/a_68_297# clknet_2_3__leaf_clk 6.28e-21
C15651 _313_/a_193_47# _010_ -9.8e-19
C15652 net28 _011_ 0.0751f
C15653 cal_itt\[0\] _000_ 1.21e-20
C15654 output35/a_27_47# _161_/a_68_297# 0.00583f
C15655 _078_ _101_ 1.01f
C15656 _058_ _332_/a_1283_21# 0.00241f
C15657 _048_ _171_/a_27_47# 0.00273f
C15658 _334_/a_27_47# _057_ 9.67e-20
C15659 net2 mask\[1\] 3.22e-20
C15660 _233_/a_27_297# net1 0.0286f
C15661 _233_/a_109_297# cal 0.00146f
C15662 net15 _017_ 6.48e-20
C15663 _058_ _111_ 0.0177f
C15664 _239_/a_277_297# _048_ 2.53e-20
C15665 _074_ _082_ 0.0436f
C15666 _136_ net4 3e-20
C15667 comp net37 8.58e-19
C15668 net27 _314_/a_543_47# 9.2e-20
C15669 _327_/a_805_47# net46 2.73e-19
C15670 _291_/a_35_297# net16 0.00571f
C15671 _028_ _049_ 8.92e-19
C15672 _047_ net34 0.103f
C15673 trim_mask\[4\] _171_/a_27_47# 7.91e-20
C15674 _316_/a_27_47# _316_/a_193_47# -0.00228f
C15675 clk _316_/a_761_289# 2.77e-19
C15676 _036_ _126_ -1.01e-24
C15677 _235_/a_297_47# _226_/a_27_47# 0.0143f
C15678 _063_ _072_ 0.00253f
C15679 ctln[6] clk 1.18e-20
C15680 _149_/a_68_297# _303_/a_193_47# 1.58e-19
C15681 _104_ net46 0.688f
C15682 net3 _317_/a_1283_21# 4.42e-20
C15683 _323_/a_27_47# net47 1.51e-19
C15684 _306_/a_448_47# _076_ 2.94e-20
C15685 _304_/a_27_47# cal_count\[3\] 8.79e-21
C15686 net10 ctln[3] 3.57e-21
C15687 _328_/a_543_47# clknet_2_2__leaf_clk 0.0363f
C15688 output33/a_27_47# _333_/a_1283_21# 9.71e-21
C15689 _304_/a_1108_47# clknet_2_3__leaf_clk 1.68e-19
C15690 _136_ _122_ 0.00727f
C15691 VPWR _079_ 0.0112f
C15692 _262_/a_465_47# _063_ 2.79e-19
C15693 VPWR trimb[3] 0.224f
C15694 _302_/a_27_297# net18 0.0108f
C15695 _284_/a_68_297# _122_ 0.00525f
C15696 _326_/a_448_47# result[5] 2.53e-19
C15697 _035_ _339_/a_476_47# 1.11e-21
C15698 _257_/a_109_297# _336_/a_193_47# 1.7e-19
C15699 net50 net30 3.8e-20
C15700 _037_ _136_ 0.00132f
C15701 _060_ calibrate 0.0293f
C15702 net54 _093_ 0.0229f
C15703 _325_/a_193_47# mask\[6\] 0.0252f
C15704 _048_ _192_/a_505_280# 0.0187f
C15705 _325_/a_651_413# _042_ 4.99e-19
C15706 _014_ _090_ 0.00256f
C15707 _041_ _338_/a_652_21# 1.13e-19
C15708 _337_/a_448_47# clknet_0_clk 6.06e-21
C15709 _185_/a_68_297# _232_/a_32_297# 1.12e-19
C15710 net3 _192_/a_174_21# 0.0616f
C15711 en_co_clk _195_/a_535_374# 0.00124f
C15712 _094_ _120_ 0.0625f
C15713 _306_/a_27_47# rebuffer4/a_27_47# 7.75e-22
C15714 net13 net55 0.314f
C15715 _058_ _135_ 1.25e-19
C15716 net25 clknet_2_1__leaf_clk 0.367f
C15717 _104_ _335_/a_651_413# 1.87e-19
C15718 _335_/a_27_47# _330_/a_1283_21# 0.011f
C15719 _327_/a_1462_47# _111_ 7.11e-19
C15720 _340_/a_1182_261# _129_ 5.56e-20
C15721 result[4] _310_/a_805_47# 1.99e-19
C15722 mask\[4\] _311_/a_1217_47# 8.37e-19
C15723 _168_/a_207_413# _107_ 0.0022f
C15724 en _315_/a_27_47# 1.21e-19
C15725 _094_ _076_ 5.86e-20
C15726 VPWR _319_/a_1108_47# 0.00989f
C15727 VPWR _230_/a_59_75# -0.00197f
C15728 _313_/a_1462_47# _010_ 4.67e-20
C15729 clkbuf_2_1__f_clk/a_110_47# _141_/a_27_47# 4.1e-19
C15730 net19 _150_/a_27_47# 8.67e-19
C15731 _012_ cal 0.00363f
C15732 _323_/a_27_47# net44 0.00995f
C15733 clk _098_ 3.92e-19
C15734 _103_ _242_/a_79_21# 7.62e-20
C15735 net2 _288_/a_145_75# 0.00219f
C15736 _326_/a_543_47# _314_/a_27_47# 8.69e-21
C15737 _326_/a_761_289# _314_/a_193_47# 5.17e-21
C15738 _326_/a_27_47# _314_/a_543_47# 1.17e-20
C15739 _326_/a_193_47# _314_/a_761_289# 5.38e-22
C15740 trim_mask\[1\] trim_val\[4\] 0.00357f
C15741 _340_/a_1182_261# _339_/a_1032_413# 5.58e-20
C15742 _340_/a_1032_413# _339_/a_1182_261# 7.12e-20
C15743 _051_ clkbuf_2_3__f_clk/a_110_47# 0.00607f
C15744 _128_ net33 0.00162f
C15745 _303_/a_543_47# _035_ 2.78e-21
C15746 trim_mask\[0\] net18 0.0149f
C15747 _195_/a_76_199# _062_ 0.0547f
C15748 _254_/a_109_297# _092_ 0.00184f
C15749 _200_/a_80_21# _092_ 0.0621f
C15750 _229_/a_27_297# _100_ 0.0509f
C15751 _090_ _243_/a_27_297# 8.83e-19
C15752 clk clknet_0_clk 0.188f
C15753 en_co_clk _332_/a_1283_21# 3.21e-19
C15754 net30 _279_/a_396_47# 0.00106f
C15755 output18/a_27_47# net17 1.18e-20
C15756 _330_/a_1270_413# net46 -1.22e-19
C15757 clknet_0_clk clone7/a_27_47# 4.43e-21
C15758 _048_ _014_ 1.92e-19
C15759 _336_/a_448_47# _119_ 0.0083f
C15760 result[5] _074_ 2.8e-19
C15761 net43 _319_/a_1270_413# -2.06e-19
C15762 VPWR _066_ 0.409f
C15763 en clknet_2_0__leaf_clk 6.3e-20
C15764 _058_ _112_ 0.0036f
C15765 _267_/a_59_75# net46 2.04e-20
C15766 net47 _133_ 1.57e-19
C15767 _198_/a_27_47# _067_ 0.062f
C15768 VPWR _336_/a_639_47# 5.1e-19
C15769 VPWR _304_/a_651_413# 9.34e-19
C15770 _198_/a_27_47# _070_ 0.00194f
C15771 net43 net55 0.00162f
C15772 output12/a_27_47# output13/a_27_47# 5.8e-21
C15773 _340_/a_476_47# cal_count\[3\] 1.54e-19
C15774 mask\[6\] _249_/a_27_297# 6.45e-20
C15775 _250_/a_27_297# mask\[5\] 0.0446f
C15776 _341_/a_448_47# _038_ 0.0308f
C15777 _341_/a_805_47# _136_ 4.9e-19
C15778 calibrate en_co_clk 0.00117f
C15779 _315_/a_27_47# _241_/a_105_352# 2.24e-21
C15780 _249_/a_109_47# net26 0.00123f
C15781 _025_ _336_/a_193_47# 1.26e-20
C15782 net4 clknet_0_clk 0.12f
C15783 clknet_2_1__leaf_clk _246_/a_109_47# 0.0012f
C15784 _325_/a_1462_47# mask\[6\] 0.00198f
C15785 _244_/a_27_297# _076_ 2.71e-19
C15786 mask\[6\] mask\[3\] 8.02e-19
C15787 _319_/a_543_47# _016_ 0.00131f
C15788 _300_/a_47_47# net40 0.00196f
C15789 _095_ _049_ 0.0214f
C15790 _325_/a_1283_21# _078_ 1.76e-20
C15791 _230_/a_59_75# _063_ 0.042f
C15792 _161_/a_150_297# net37 3.96e-19
C15793 _015_ _317_/a_193_47# 5.56e-20
C15794 _338_/a_652_21# net18 0.0113f
C15795 _320_/a_193_47# _121_ 1.99e-19
C15796 _341_/a_27_47# _341_/a_193_47# -0.266f
C15797 _228_/a_297_47# _052_ 0.00498f
C15798 _320_/a_1283_21# net44 0.0669f
C15799 output37/a_27_47# output40/a_27_47# 0.00222f
C15800 ctlp[7] VPWR 0.31f
C15801 cal_itt\[0\] _190_/a_215_47# 1.53e-19
C15802 cal_itt\[1\] _190_/a_27_47# 7.64e-19
C15803 cal_itt\[2\] _190_/a_465_47# 5.71e-20
C15804 net43 _067_ 0.00265f
C15805 net13 _337_/a_805_47# 4.26e-19
C15806 net43 _070_ 6.25e-20
C15807 _321_/a_1108_47# net53 4.72e-19
C15808 _169_/a_215_311# _318_/a_193_47# 2.81e-20
C15809 _332_/a_1108_47# net40 7.08e-20
C15810 _336_/a_651_413# _266_/a_68_297# 4.89e-21
C15811 net28 _313_/a_761_289# 0.022f
C15812 _029_ net40 0.0203f
C15813 _078_ _248_/a_27_297# 4.2e-21
C15814 _329_/a_27_47# trim_mask\[2\] 2.05e-19
C15815 _048_ _243_/a_27_297# 1.73e-20
C15816 clknet_0_clk _073_ 5.34e-22
C15817 VPWR _321_/a_651_413# 9.24e-19
C15818 net46 net37 1.7e-19
C15819 _339_/a_27_47# _122_ 6.27e-21
C15820 _135_ en_co_clk 0.00293f
C15821 _110_ _104_ 0.0117f
C15822 clone1/a_27_47# _242_/a_297_47# 0.0382f
C15823 _250_/a_109_297# _084_ 1.14e-19
C15824 mask\[6\] _220_/a_113_297# 0.00553f
C15825 _034_ net30 0.0547f
C15826 mask\[5\] _009_ 1.37e-19
C15827 _333_/a_1283_21# _056_ 1.36e-20
C15828 trim[2] trim[3] 0.0486f
C15829 _041_ _339_/a_476_47# 0.043f
C15830 net47 _339_/a_1140_413# 2.79e-20
C15831 mask\[1\] mask\[0\] 0.0883f
C15832 VPWR _337_/a_651_413# 9.52e-19
C15833 VPWR _313_/a_543_47# 0.0308f
C15834 VPWR _047_ 0.15f
C15835 _106_ _191_/a_27_297# 5e-19
C15836 _051_ cal_count\[3\] 1.48e-20
C15837 output24/a_27_47# mask\[1\] 2.25e-19
C15838 _037_ _339_/a_27_47# 2.81e-20
C15839 _050_ net45 4.41e-19
C15840 _260_/a_93_21# net55 3.94e-21
C15841 _293_/a_81_21# cal_count\[1\] 0.00317f
C15842 _310_/a_27_47# _310_/a_193_47# -0.0199f
C15843 _316_/a_448_47# _013_ 0.0116f
C15844 _097_ _092_ 0.0631f
C15845 trim_mask\[2\] _115_ 0.0818f
C15846 _159_/a_27_47# _313_/a_761_289# 0.00138f
C15847 _071_ _092_ 0.0264f
C15848 _292_/a_78_199# net47 0.00916f
C15849 _015_ _318_/a_1283_21# 4.1e-20
C15850 state\[2\] _318_/a_27_47# 6.04e-19
C15851 _051_ _331_/a_27_47# 0.0011f
C15852 _308_/a_651_413# _006_ 1.65e-21
C15853 _033_ _119_ 0.727f
C15854 _103_ _050_ 0.0737f
C15855 _337_/a_193_47# _090_ 2.84e-21
C15856 _306_/a_1108_47# _305_/a_543_47# 5.01e-19
C15857 _326_/a_651_413# _310_/a_543_47# 3.01e-20
C15858 _326_/a_1108_47# _310_/a_1108_47# 8.34e-21
C15859 _323_/a_1283_21# net18 3.42e-19
C15860 _320_/a_761_289# clknet_0_clk 0.00358f
C15861 _262_/a_27_47# _092_ 8.22e-20
C15862 net43 _321_/a_805_47# 8.55e-19
C15863 _326_/a_761_289# _074_ 0.00387f
C15864 _050_ _065_ 0.0226f
C15865 VPWR net47 0.723f
C15866 VPWR _143_/a_150_297# -6.52e-19
C15867 _338_/a_1602_47# clknet_2_3__leaf_clk 0.0097f
C15868 output20/a_27_47# _312_/a_651_413# 2.85e-19
C15869 _320_/a_193_47# _320_/a_448_47# -0.00363f
C15870 _042_ mask\[2\] 0.0316f
C15871 _130_ output40/a_27_47# 5.69e-21
C15872 _309_/a_193_47# _081_ 0.00817f
C15873 calibrate _228_/a_297_47# 6.83e-19
C15874 clknet_2_1__leaf_clk _208_/a_439_47# 5.61e-19
C15875 _060_ _192_/a_27_47# 1.36e-20
C15876 _334_/a_805_47# net46 4.47e-19
C15877 _200_/a_209_297# _053_ 2.12e-19
C15878 _316_/a_27_47# net41 0.19f
C15879 VPWR _340_/a_1140_413# -2.86e-19
C15880 output32/a_27_47# net31 0.00233f
C15881 net24 _007_ 3.43e-21
C15882 net43 _313_/a_448_47# 0.00195f
C15883 _189_/a_27_47# _306_/a_1108_47# 4.15e-22
C15884 _008_ _321_/a_1108_47# 1.37e-20
C15885 _315_/a_1108_47# _095_ 7.61e-19
C15886 _315_/a_1283_21# _099_ 3e-19
C15887 _129_ _298_/a_78_199# 1.27e-19
C15888 _299_/a_215_297# _133_ 4.06e-19
C15889 net12 _040_ 1.15e-20
C15890 net12 net41 5.07e-20
C15891 _336_/a_543_47# trim_mask\[4\] 0.0358f
C15892 cal_count\[1\] _144_/a_27_47# 0.0563f
C15893 net2 _062_ 1.3e-20
C15894 _117_ _057_ 7.58e-20
C15895 _328_/a_1108_47# _327_/a_1283_21# 2.15e-22
C15896 _308_/a_193_47# _307_/a_761_289# 6.96e-20
C15897 _308_/a_27_47# _307_/a_543_47# 1.1e-20
C15898 net27 output29/a_27_47# 1.35e-21
C15899 _305_/a_27_47# rebuffer4/a_27_47# 8.38e-19
C15900 net17 _339_/a_381_47# 8.46e-20
C15901 _232_/a_304_297# en_co_clk 1.27e-19
C15902 _230_/a_145_75# _107_ 8.43e-20
C15903 net24 mask\[3\] 0.0026f
C15904 _338_/a_1056_47# net18 4e-19
C15905 _050_ _319_/a_27_47# 1.58e-21
C15906 _107_ _100_ 0.0129f
C15907 VPWR _316_/a_27_47# 0.108f
C15908 rebuffer1/a_75_212# _108_ 0.0104f
C15909 _303_/a_543_47# _041_ 3.11e-20
C15910 _332_/a_27_47# _332_/a_761_289# -0.00784f
C15911 net47 _303_/a_805_47# 3.21e-21
C15912 _303_/a_27_47# _338_/a_381_47# 7.45e-21
C15913 _189_/a_27_47# _075_ 4.85e-20
C15914 net13 _121_ 3.21e-20
C15915 VPWR net12 1.3f
C15916 _337_/a_1283_21# _263_/a_297_47# 1.43e-21
C15917 _335_/a_1270_413# net46 6.96e-20
C15918 _328_/a_1270_413# _058_ 3.74e-20
C15919 _264_/a_27_297# net19 2.68e-19
C15920 state\[0\] _049_ 4.22e-19
C15921 clk _331_/a_1108_47# 9.3e-19
C15922 output14/a_27_47# net29 0.00225f
C15923 _040_ net44 0.279f
C15924 _231_/a_161_47# _264_/a_27_297# 3.44e-21
C15925 net51 rebuffer4/a_27_47# 0.00335f
C15926 _258_/a_27_297# _119_ 9.01e-19
C15927 net12 _322_/a_1283_21# 0.00904f
C15928 net27 mask\[6\] 0.348f
C15929 net12 _331_/a_1283_21# 0.00486f
C15930 output8/a_27_47# trim[3] 6.33e-19
C15931 mask\[6\] _222_/a_113_297# 3.61e-19
C15932 _329_/a_1217_47# trim_mask\[2\] 1.33e-19
C15933 _026_ _258_/a_373_47# 4.62e-20
C15934 _333_/a_1283_21# _173_/a_27_47# 4.74e-19
C15935 VPWR _258_/a_373_47# -7.36e-19
C15936 net43 _102_ 0.00624f
C15937 _324_/a_1108_47# net44 0.0112f
C15938 net3 net55 0.134f
C15939 _332_/a_651_413# net46 0.0266f
C15940 _048_ _337_/a_193_47# 1.59e-20
C15941 fanout46/a_27_47# net46 0.0192f
C15942 _207_/a_109_297# _049_ 0.00121f
C15943 wire42/a_75_212# _092_ 0.00229f
C15944 _110_ _330_/a_1270_413# 1.46e-19
C15945 clknet_2_1__leaf_clk net15 1.21f
C15946 _041_ _339_/a_1224_47# 0.00127f
C15947 _324_/a_1283_21# _323_/a_27_47# 0.00384f
C15948 VPWR net44 2.28f
C15949 _143_/a_150_297# net52 1.32e-19
C15950 _256_/a_373_47# clknet_2_2__leaf_clk 0.00102f
C15951 _336_/a_805_47# _107_ 1.48e-19
C15952 net47 _063_ 0.0107f
C15953 _019_ _321_/a_1108_47# 4.75e-19
C15954 _264_/a_27_297# _107_ 0.0246f
C15955 _308_/a_27_47# _138_/a_27_47# 0.0116f
C15956 _110_ _267_/a_59_75# 0.0266f
C15957 _094_ clkbuf_2_0__f_clk/a_110_47# 0.00233f
C15958 net9 _053_ 6.64e-20
C15959 result[0] _307_/a_1283_21# 1.48e-19
C15960 cal _315_/a_543_47# 0.00152f
C15961 _113_ _332_/a_193_47# 1.3e-20
C15962 _074_ _310_/a_1283_21# 0.0107f
C15963 mask\[7\] _101_ 0.0667f
C15964 _322_/a_1283_21# net44 0.0586f
C15965 _309_/a_27_47# _308_/a_27_47# 6.48e-21
C15966 _233_/a_373_47# calibrate 3.04e-19
C15967 _233_/a_27_297# _012_ 0.0443f
C15968 _340_/a_27_47# _001_ 1.09e-19
C15969 net31 _113_ 2.53e-20
C15970 net21 _313_/a_651_413# 2.12e-19
C15971 _036_ net47 0.0224f
C15972 _325_/a_193_47# _321_/a_193_47# 1.07e-20
C15973 _002_ _076_ 1.23e-19
C15974 net43 _006_ 8.08e-19
C15975 net26 _076_ 0.00189f
C15976 _226_/a_27_47# _049_ 6.98e-19
C15977 _048_ _106_ 0.2f
C15978 VPWR _301_/a_47_47# 0.0232f
C15979 net30 output30/a_27_47# 0.0508f
C15980 net9 _057_ 0.0755f
C15981 _187_/a_212_413# net2 1.13e-20
C15982 VPWR _003_ 0.0965f
C15983 net12 net52 4.96e-20
C15984 _022_ mask\[2\] 9.54e-25
C15985 net30 _278_/a_109_297# 8.41e-21
C15986 _269_/a_299_297# net46 0.00155f
C15987 _341_/a_1283_21# cal_count\[3\] 0.0485f
C15988 _302_/a_27_297# trim_mask\[4\] 1.27e-19
C15989 VPWR _338_/a_562_413# 4.03e-20
C15990 VPWR _341_/a_27_47# 0.0423f
C15991 _341_/a_639_47# clknet_2_3__leaf_clk 0.00133f
C15992 en_co_clk _192_/a_27_47# 0.00756f
C15993 cal_itt\[0\] en_co_clk 0.426f
C15994 net2 _332_/a_193_47# 2.47e-19
C15995 net43 _121_ 0.0321f
C15996 _316_/a_1217_47# net41 8.27e-19
C15997 net43 _010_ 0.0145f
C15998 VPWR _274_/a_75_212# 0.0904f
C15999 _339_/a_27_47# _339_/a_562_413# -0.0012f
C16000 _339_/a_193_47# _339_/a_381_47# -0.00883f
C16001 fanout46/a_27_47# _335_/a_651_413# 1.44e-19
C16002 net31 net2 0.00231f
C16003 net13 _320_/a_448_47# 3.09e-19
C16004 VPWR _299_/a_215_297# 0.0224f
C16005 _106_ trim_mask\[4\] 1.48e-20
C16006 _227_/a_209_311# _062_ 1.75e-20
C16007 output15/a_27_47# net15 0.0335f
C16008 trim_mask\[1\] _334_/a_543_47# 8.39e-22
C16009 _272_/a_81_21# _334_/a_761_289# 6.84e-20
C16010 _272_/a_299_297# _334_/a_193_47# 4.55e-20
C16011 _320_/a_543_47# _040_ 0.0357f
C16012 _096_ _241_/a_297_47# 7.33e-19
C16013 _053_ _262_/a_109_297# 0.00471f
C16014 clknet_2_1__leaf_clk _314_/a_1108_47# 4.87e-19
C16015 net1 net45 1.51e-20
C16016 net22 output30/a_27_47# 0.00146f
C16017 _051_ _242_/a_297_47# 1.36e-20
C16018 _336_/a_27_47# trim_val\[4\] 6.4e-19
C16019 _264_/a_27_297# _279_/a_27_47# 6.6e-19
C16020 VPWR _316_/a_1217_47# 3.62e-20
C16021 trim_mask\[0\] _333_/a_193_47# 1.91e-19
C16022 _332_/a_805_47# _108_ 6.71e-19
C16023 _228_/a_297_47# _170_/a_384_47# 2.15e-20
C16024 net44 net52 0.0125f
C16025 net44 _063_ 1.71e-20
C16026 _110_ net37 5.19e-20
C16027 trim_mask\[0\] _265_/a_81_21# 0.0556f
C16028 _059_ net30 1.8e-20
C16029 _146_/a_68_297# _310_/a_1108_47# 3.64e-19
C16030 output14/a_27_47# ctlp[1] 5.95e-22
C16031 _058_ net33 0.0312f
C16032 output32/a_27_47# trim_val\[1\] 1.5e-19
C16033 clk clknet_2_2__leaf_clk 0.0052f
C16034 VPWR _320_/a_543_47# 0.00138f
C16035 net54 _243_/a_27_297# 0.00149f
C16036 _339_/a_381_47# clknet_2_3__leaf_clk 6.75e-19
C16037 _104_ net45 2.79e-21
C16038 _286_/a_535_374# _123_ 0.00177f
C16039 trim_mask\[0\] _048_ 0.124f
C16040 _104_ rebuffer3/a_75_212# 2.43e-21
C16041 clknet_2_1__leaf_clk _310_/a_193_47# 0.595f
C16042 fanout44/a_27_47# net55 4.46e-19
C16043 _333_/a_639_47# net32 1.09e-19
C16044 _322_/a_543_47# _320_/a_1283_21# 1.58e-20
C16045 _326_/a_27_47# mask\[6\] 5.74e-21
C16046 en input4/a_27_47# 1.99e-20
C16047 _326_/a_761_289# net26 7.11e-20
C16048 net15 _317_/a_651_413# 0.00245f
C16049 _333_/a_1283_21# _172_/a_68_297# 2.46e-19
C16050 net12 _083_ 0.00879f
C16051 _308_/a_193_47# net43 0.0162f
C16052 _308_/a_761_289# _005_ 9.52e-19
C16053 _117_ _027_ 1.84e-20
C16054 _116_ net46 3.1e-19
C16055 ctlp[6] _312_/a_27_47# 6.16e-19
C16056 _104_ _103_ 0.00313f
C16057 _258_/a_109_47# clknet_2_2__leaf_clk 0.00309f
C16058 comp cal_count\[2\] 8.28e-20
C16059 trim_mask\[0\] trim_mask\[4\] 0.115f
C16060 cal_count\[1\] net34 1.15e-20
C16061 _306_/a_651_413# _049_ 5.46e-20
C16062 _341_/a_27_47# _063_ 2.69e-20
C16063 net49 rebuffer1/a_75_212# 2.47e-19
C16064 _308_/a_639_47# net14 7.18e-19
C16065 net4 clknet_2_2__leaf_clk 0.744f
C16066 _306_/a_1108_47# net30 6.43e-20
C16067 _119_ clkbuf_2_3__f_clk/a_110_47# 2.64e-20
C16068 VPWR _323_/a_805_47# 3.81e-19
C16069 VPWR _307_/a_1283_21# 0.0439f
C16070 clknet_2_0__leaf_clk en_co_clk 0.0128f
C16071 net31 trim_val\[1\] 0.0297f
C16072 state\[0\] state\[1\] 0.215f
C16073 _329_/a_1108_47# _026_ 3.46e-19
C16074 result[7] _314_/a_27_47# 0.00352f
C16075 _329_/a_1108_47# VPWR 0.0203f
C16076 _305_/a_1283_21# net2 1.58e-19
C16077 _266_/a_68_297# clkbuf_2_2__f_clk/a_110_47# 1.71e-19
C16078 _309_/a_193_47# net14 0.0121f
C16079 _335_/a_639_47# _032_ 3.71e-19
C16080 _321_/a_761_289# net25 4.62e-21
C16081 _321_/a_193_47# mask\[3\] 2.82e-19
C16082 _313_/a_1283_21# _155_/a_68_297# 7.54e-19
C16083 _104_ _105_ 8.7e-20
C16084 _092_ _206_/a_27_93# 5.28e-20
C16085 _078_ _077_ 0.0145f
C16086 _309_/a_193_47# _309_/a_761_289# -0.00517f
C16087 _083_ net44 0.00381f
C16088 _325_/a_1283_21# _313_/a_1108_47# 8.78e-21
C16089 cal_count\[1\] _299_/a_298_297# 6.02e-20
C16090 _061_ _135_ 5.21e-19
C16091 net44 _312_/a_1270_413# 1.41e-19
C16092 clknet_0_clk _101_ 0.00175f
C16093 VPWR _341_/a_1217_47# 3.07e-20
C16094 _323_/a_543_47# _000_ 1.96e-19
C16095 _110_ trim[1] 5.23e-20
C16096 _320_/a_1108_47# _101_ 1.13e-19
C16097 _320_/a_543_47# net52 4.37e-19
C16098 _306_/a_193_47# clknet_2_0__leaf_clk 0.00116f
C16099 clknet_2_1__leaf_clk _311_/a_543_47# 3.51e-20
C16100 _313_/a_27_47# _158_/a_68_297# 4.15e-19
C16101 _303_/a_651_413# clknet_2_3__leaf_clk 8.49e-19
C16102 _323_/a_27_47# net19 0.0156f
C16103 output8/a_27_47# _057_ 0.0648f
C16104 _327_/a_27_47# _302_/a_27_297# 8.93e-19
C16105 _188_/a_27_47# en_co_clk 0.00106f
C16106 net48 _334_/a_1108_47# 4.81e-19
C16107 _018_ _310_/a_1108_47# 5.62e-19
C16108 VPWR _308_/a_639_47# 7.36e-19
C16109 _306_/a_1108_47# _072_ 4.11e-19
C16110 _306_/a_448_47# cal_itt\[3\] 1.38e-19
C16111 _182_/a_27_47# net32 1.88e-19
C16112 _065_ _208_/a_439_47# 4.22e-21
C16113 _337_/a_1283_21# _099_ 1.09e-21
C16114 _337_/a_543_47# _092_ 3.51e-19
C16115 _264_/a_27_297# _118_ 0.0112f
C16116 _292_/a_215_47# _339_/a_1602_47# 9.75e-21
C16117 _052_ _049_ 0.419f
C16118 net13 net53 0.0143f
C16119 _110_ _332_/a_651_413# 2.02e-20
C16120 _079_ output30/a_27_47# 0.00107f
C16121 VPWR _237_/a_218_47# -4.49e-19
C16122 net26 _310_/a_1283_21# 6.96e-20
C16123 VPWR _309_/a_193_47# -0.276f
C16124 _110_ fanout46/a_27_47# 0.00447f
C16125 _050_ _282_/a_68_297# 1.25e-19
C16126 _074_ _042_ 0.448f
C16127 _328_/a_27_47# net46 0.00477f
C16128 _253_/a_81_21# net25 8.35e-19
C16129 _290_/a_297_47# cal_count\[0\] 5.23e-19
C16130 VPWR _339_/a_956_413# -5.25e-19
C16131 _341_/a_193_47# _231_/a_161_47# 3.72e-19
C16132 _302_/a_109_47# _092_ 0.0017f
C16133 _002_ _068_ 6.92e-19
C16134 _104_ _336_/a_1283_21# 0.0587f
C16135 net54 _337_/a_193_47# 3.54e-19
C16136 ctln[1] _317_/a_27_47# 1.75e-20
C16137 VPWR ctln[7] 0.0616f
C16138 _006_ _080_ 9.8e-20
C16139 _068_ net26 3.89e-20
C16140 _324_/a_761_289# net53 5.65e-19
C16141 _019_ _320_/a_193_47# 1.24e-19
C16142 _275_/a_299_297# net18 0.00664f
C16143 net30 _137_/a_150_297# 1.66e-19
C16144 net2 _123_ 0.0507f
C16145 _326_/a_543_47# _078_ 0.00326f
C16146 net7 clknet_2_0__leaf_clk 2.04e-20
C16147 net15 net45 1.2f
C16148 net13 _322_/a_448_47# 0.00788f
C16149 _294_/a_68_297# net33 0.00445f
C16150 cal_count\[1\] _133_ 0.00162f
C16151 net3 _121_ 1.77e-21
C16152 trim[4] _131_ 3.48e-21
C16153 _308_/a_1462_47# net43 9.59e-19
C16154 _337_/a_651_413# _034_ 7.15e-19
C16155 _097_ _233_/a_27_297# 7.99e-20
C16156 VPWR _324_/a_1283_21# 0.0259f
C16157 en_co_clk net33 4.99e-19
C16158 _119_ cal_count\[3\] 3.29e-21
C16159 VPWR _280_/a_75_212# 0.018f
C16160 _189_/a_27_47# _170_/a_81_21# 1.01e-20
C16161 _322_/a_193_47# net53 2.02e-19
C16162 net31 _296_/a_113_47# 1.37e-19
C16163 _110_ _269_/a_299_297# 4.72e-19
C16164 _341_/a_193_47# _001_ 2.94e-19
C16165 _309_/a_1283_21# net43 -0.00725f
C16166 _309_/a_193_47# net23 6.13e-20
C16167 _304_/a_27_47# en_co_clk 7.65e-20
C16168 output20/a_27_47# output19/a_27_47# 3.07e-21
C16169 mask\[0\] _137_/a_68_297# 0.0644f
C16170 net22 _137_/a_150_297# 1.11e-20
C16171 _327_/a_27_47# trim_mask\[0\] 8.62e-19
C16172 net4 _279_/a_204_297# 0.00404f
C16173 net16 rebuffer2/a_75_212# 0.00604f
C16174 _257_/a_27_297# _119_ 1.41e-19
C16175 VPWR _198_/a_181_47# -1.83e-19
C16176 cal_itt\[2\] _068_ 0.0725f
C16177 net15 _065_ 0.00704f
C16178 _305_/a_761_289# _002_ 0.0231f
C16179 net16 _332_/a_1283_21# 0.00684f
C16180 _277_/a_75_212# _335_/a_27_47# 2.48e-20
C16181 output21/a_27_47# net27 6.42e-21
C16182 VPWR _322_/a_543_47# 6.9e-19
C16183 net9 _300_/a_47_47# 0.00155f
C16184 _329_/a_1283_21# clknet_2_2__leaf_clk 0.0163f
C16185 _314_/a_193_47# _011_ 0.0423f
C16186 _314_/a_543_47# _086_ 9.06e-19
C16187 net16 _111_ 7.22e-22
C16188 VPWR _257_/a_373_47# -6.84e-19
C16189 VPWR _331_/a_543_47# 0.0198f
C16190 _066_ _193_/a_109_297# 0.00125f
C16191 _311_/a_448_47# net26 0.0163f
C16192 net5 trim[4] 2.79e-19
C16193 _233_/a_27_297# _315_/a_543_47# 0.00338f
C16194 _233_/a_109_297# _315_/a_761_289# 3.22e-19
C16195 _064_ _091_ 0.003f
C16196 _322_/a_193_47# _322_/a_448_47# -0.00482f
C16197 _309_/a_543_47# _101_ 3.1e-20
C16198 _259_/a_27_297# trim_mask\[0\] 4.06e-21
C16199 _064_ _256_/a_109_297# 0.00118f
C16200 net43 net53 0.0152f
C16201 _324_/a_27_47# _312_/a_193_47# 2.78e-21
C16202 _324_/a_193_47# _312_/a_27_47# 1.15e-19
C16203 _305_/a_805_47# clknet_2_1__leaf_clk 1.33e-20
C16204 VPWR _229_/a_27_297# 0.0206f
C16205 _250_/a_27_297# clknet_2_1__leaf_clk 0.045f
C16206 _331_/a_193_47# _331_/a_448_47# -0.00297f
C16207 calibrate _049_ 0.139f
C16208 VPWR _303_/a_639_47# 4.33e-19
C16209 _185_/a_68_297# _316_/a_193_47# 2.13e-20
C16210 _245_/a_27_297# _101_ 0.058f
C16211 _323_/a_1217_47# net19 2.55e-19
C16212 cal_itt\[0\] cal_count\[0\] 4.18e-21
C16213 _117_ _032_ 0.277f
C16214 net15 _319_/a_27_47# 0.0217f
C16215 _327_/a_543_47# _136_ 0.00139f
C16216 _305_/a_193_47# _203_/a_59_75# 6.15e-20
C16217 net9 _029_ 0.00231f
C16218 _081_ mask\[1\] 0.274f
C16219 _235_/a_79_21# _243_/a_109_297# 2.02e-20
C16220 _308_/a_193_47# _080_ 6.57e-20
C16221 net28 _101_ 5.23e-20
C16222 state\[2\] fanout45/a_27_47# 2.77e-20
C16223 cal_itt\[2\] _305_/a_761_289# 6.11e-19
C16224 cal_itt\[0\] _305_/a_193_47# 4.7e-21
C16225 _329_/a_448_47# trim_mask\[3\] 8.81e-19
C16226 _053_ _091_ 2.3e-19
C16227 _022_ _074_ 1.49e-19
C16228 net35 _136_ 4.2e-19
C16229 _324_/a_448_47# _101_ 4.94e-21
C16230 _078_ _310_/a_1108_47# 0.0108f
C16231 VPWR _309_/a_1462_47# 3.65e-19
C16232 _120_ net55 2.09e-21
C16233 _303_/a_761_289# _000_ 3.71e-19
C16234 _110_ _116_ 0.406f
C16235 _326_/a_448_47# _011_ 2.6e-20
C16236 _328_/a_1217_47# net46 5.14e-19
C16237 result[2] _310_/a_27_47# 7.53e-20
C16238 _337_/a_27_47# en_co_clk 0.00752f
C16239 _233_/a_109_297# net45 0.00122f
C16240 _292_/a_78_199# cal_count\[1\] 0.00271f
C16241 _292_/a_215_47# _128_ 8.6e-19
C16242 _064_ _033_ 0.00276f
C16243 _001_ _133_ 5.05e-20
C16244 clkbuf_2_0__f_clk/a_110_47# _192_/a_174_21# 4.98e-19
C16245 _198_/a_181_47# _063_ 1.28e-19
C16246 state\[0\] _167_/a_161_47# 0.00282f
C16247 input1/a_75_212# _316_/a_27_47# 4.41e-21
C16248 _060_ _051_ 0.26f
C16249 _015_ _316_/a_27_47# 3.05e-21
C16250 _328_/a_1108_47# _113_ 0.00303f
C16251 _328_/a_1283_21# _030_ 6.43e-19
C16252 _322_/a_1108_47# _101_ 0.0104f
C16253 input3/a_75_212# output41/a_27_47# 0.0101f
C16254 _270_/a_59_75# _332_/a_27_47# 7.88e-19
C16255 _219_/a_109_297# _218_/a_113_297# 1.95e-20
C16256 clkbuf_2_2__f_clk/a_110_47# _279_/a_314_297# 1.04e-20
C16257 net13 _019_ 0.105f
C16258 clknet_2_1__leaf_clk _009_ 0.113f
C16259 _135_ net16 0.00779f
C16260 VPWR cal_count\[1\] 0.728f
C16261 _305_/a_1108_47# net30 8.45e-20
C16262 _053_ _302_/a_373_47# 0.00193f
C16263 net44 _034_ 3.16e-19
C16264 _321_/a_448_47# mask\[2\] 6.41e-20
C16265 _303_/a_639_47# _063_ 3.94e-20
C16266 _082_ _006_ 0.00503f
C16267 net8 _334_/a_1283_21# 0.0111f
C16268 _323_/a_448_47# _152_/a_68_297# 1.63e-20
C16269 _327_/a_1217_47# trim_mask\[0\] 6.68e-21
C16270 _327_/a_1270_413# _024_ 4.33e-20
C16271 net43 _016_ 3.64e-19
C16272 clknet_2_0__leaf_clk _039_ 0.00324f
C16273 _053_ _340_/a_381_47# 8.64e-20
C16274 ctln[5] output12/a_27_47# 2.68e-20
C16275 mask\[6\] _250_/a_109_297# 0.0011f
C16276 _312_/a_1108_47# net20 0.00215f
C16277 VPWR _260_/a_256_47# -7.83e-19
C16278 net42 _170_/a_81_21# 7.65e-19
C16279 _042_ net26 0.0409f
C16280 _074_ _315_/a_448_47# 0.00471f
C16281 _076_ _070_ 2.23e-20
C16282 calibrate _315_/a_1108_47# 0.0532f
C16283 _012_ _315_/a_761_289# 8.16e-19
C16284 _320_/a_1283_21# _248_/a_109_297# 1.26e-21
C16285 _337_/a_1108_47# _226_/a_27_47# 9.99e-20
C16286 _064_ _258_/a_27_297# 0.00296f
C16287 _322_/a_193_47# _019_ 0.0348f
C16288 _064_ _024_ 9.91e-20
C16289 _300_/a_377_297# cal_count\[2\] 2.46e-19
C16290 _331_/a_193_47# _028_ 0.33f
C16291 _331_/a_761_289# clknet_2_2__leaf_clk 1.82e-19
C16292 _324_/a_1108_47# net19 0.00166f
C16293 clkbuf_2_1__f_clk/a_110_47# _078_ 0.0012f
C16294 _124_ _065_ 5.23e-20
C16295 _317_/a_27_47# _317_/a_1283_21# -9.15e-20
C16296 _317_/a_193_47# _317_/a_543_47# -0.0129f
C16297 net48 trim_mask\[1\] 1.98e-20
C16298 net54 _316_/a_1108_47# 2.02e-20
C16299 _060_ _316_/a_1283_21# 6.36e-21
C16300 trim_mask\[0\] output35/a_27_47# 9.4e-19
C16301 _272_/a_299_297# trim_val\[2\] 0.00842f
C16302 _143_/a_68_297# mask\[2\] 0.0432f
C16303 VPWR _312_/a_651_413# 1.95e-32
C16304 _094_ _319_/a_1283_21# 1.33e-20
C16305 net15 _319_/a_1217_47# 6.04e-20
C16306 _232_/a_304_297# _049_ 0.0014f
C16307 _110_ _328_/a_27_47# 5.55e-20
C16308 VPWR net19 1.21f
C16309 _320_/a_1283_21# mask\[1\] 0.0316f
C16310 _305_/a_1108_47# _072_ 0.059f
C16311 ctln[0] VGND 0.459f
C16312 net6 VGND 0.338f
C16313 output6/a_27_47# VGND 0.326f
C16314 sample VGND 0.177f
C16315 output30/a_27_47# VGND 0.626f
C16316 valid VGND 0.474f
C16317 net41 VGND 3.13f
C16318 output41/a_27_47# VGND 0.562f
C16319 _201_/a_113_47# VGND 9.84e-20
C16320 net40 VGND 1.81f
C16321 _278_/a_27_47# VGND 0.0727f
C16322 _278_/a_109_297# VGND -3.12e-19
C16323 net53 VGND 1.73f
C16324 rebuffer6/a_27_47# VGND 0.263f
C16325 _131_ VGND 1.23f
C16326 cal_count\[2\] VGND 0.616f
C16327 _295_/a_113_47# VGND -1.03e-21
C16328 clkc VGND 0.215f
C16329 output5/a_27_47# VGND 0.274f
C16330 trimb[4] VGND 0.225f
C16331 output40/a_27_47# VGND 0.653f
C16332 _070_ VGND 0.435f
C16333 _202_/a_297_47# VGND 0.0845f
C16334 _202_/a_382_297# VGND -5.84e-19
C16335 _202_/a_79_21# VGND 0.159f
C16336 _118_ VGND 0.291f
C16337 trim_val\[4\] VGND 0.427f
C16338 _279_/a_490_47# VGND -2.41e-19
C16339 _279_/a_206_47# VGND -0.00352f
C16340 _279_/a_314_297# VGND 0.00252f
C16341 _279_/a_204_297# VGND 0.00251f
C16342 _279_/a_396_47# VGND 0.407f
C16343 _279_/a_27_47# VGND 0.186f
C16344 _150_/a_27_47# VGND 0.235f
C16345 rebuffer5/a_161_47# VGND 0.608f
C16346 _132_ VGND 0.267f
C16347 _296_/a_113_47# VGND -1.21e-19
C16348 _072_ VGND 0.439f
C16349 cal_itt\[3\] VGND 0.59f
C16350 _203_/a_145_75# VGND 3.38e-19
C16351 _203_/a_59_75# VGND 0.18f
C16352 _084_ VGND 0.152f
C16353 _220_/a_199_47# VGND -9.41e-20
C16354 _220_/a_113_297# VGND 0.0293f
C16355 net18 VGND 2.59f
C16356 rebuffer4/a_27_47# VGND 0.248f
C16357 _297_/a_285_47# VGND 0.0387f
C16358 _297_/a_129_47# VGND 3.82e-19
C16359 _297_/a_377_297# VGND 0.00288f
C16360 _297_/a_47_47# VGND 0.313f
C16361 _003_ VGND 0.476f
C16362 _073_ VGND 0.66f
C16363 _204_/a_75_212# VGND 0.306f
C16364 _009_ VGND 0.376f
C16365 _221_/a_109_297# VGND -8.02e-19
C16366 _044_ VGND 0.356f
C16367 _152_/a_150_297# VGND -2.33e-19
C16368 _152_/a_68_297# VGND 0.179f
C16369 rebuffer3/a_75_212# VGND 0.26f
C16370 _133_ VGND 0.253f
C16371 _298_/a_215_47# VGND 0.0858f
C16372 _298_/a_493_297# VGND -2.84e-19
C16373 _298_/a_292_297# VGND -0.00126f
C16374 _298_/a_78_199# VGND 0.157f
C16375 _205_/a_27_47# VGND 0.64f
C16376 clone7/a_27_47# VGND 0.359f
C16377 _085_ VGND 0.279f
C16378 _222_/a_199_47# VGND -2.87e-19
C16379 _222_/a_113_297# VGND 0.0344f
C16380 _153_/a_27_47# VGND 0.276f
C16381 rebuffer2/a_75_212# VGND 0.296f
C16382 _130_ VGND 0.233f
C16383 _129_ VGND 0.598f
C16384 _299_/a_382_47# VGND -8.4e-19
C16385 _299_/a_298_297# VGND 0.00857f
C16386 _299_/a_215_297# VGND 0.159f
C16387 _299_/a_27_413# VGND 0.187f
C16388 _054_ VGND 0.355f
C16389 _049_ VGND 3f
C16390 _170_/a_384_47# VGND -2.58e-19
C16391 _170_/a_299_297# VGND 0.0325f
C16392 _170_/a_81_21# VGND 0.145f
C16393 _206_/a_206_47# VGND -0.00138f
C16394 _206_/a_27_93# VGND 0.176f
C16395 _039_ VGND 0.193f
C16396 _137_/a_150_297# VGND -1.25e-19
C16397 _137_/a_68_297# VGND 0.178f
C16398 net11 VGND 0.318f
C16399 net19 VGND 1.9f
C16400 _223_/a_109_297# VGND -3.5e-19
C16401 _108_ VGND 3.12f
C16402 rebuffer1/a_75_212# VGND 0.246f
C16403 _098_ VGND 0.86f
C16404 _240_/a_109_297# VGND -0.00104f
C16405 net30 VGND 1.55f
C16406 _171_/a_27_47# VGND 0.382f
C16407 _076_ VGND 0.859f
C16408 _207_/a_109_297# VGND -8.91e-19
C16409 _138_/a_27_47# VGND 0.249f
C16410 net29 VGND 1.34f
C16411 _224_/a_199_47# VGND -4.41e-19
C16412 _224_/a_113_297# VGND 0.0319f
C16413 _045_ VGND 0.482f
C16414 _155_/a_150_297# VGND -2.86e-19
C16415 _155_/a_68_297# VGND 0.151f
C16416 _092_ VGND 3.53f
C16417 _099_ VGND 1.97f
C16418 _095_ VGND 0.91f
C16419 _241_/a_297_47# VGND 0.0216f
C16420 _241_/a_388_297# VGND -8.87e-19
C16421 _241_/a_105_352# VGND 0.169f
C16422 _055_ VGND 0.219f
C16423 _172_/a_150_297# VGND -1.29e-19
C16424 _172_/a_68_297# VGND 0.163f
C16425 _310_/a_1462_47# VGND -8.75e-19
C16426 _310_/a_1217_47# VGND -4.82e-19
C16427 _310_/a_805_47# VGND 1.8e-19
C16428 _310_/a_639_47# VGND 3.35e-19
C16429 _310_/a_1270_413# VGND 4.62e-20
C16430 _310_/a_651_413# VGND 0.00625f
C16431 _310_/a_448_47# VGND 0.0148f
C16432 _310_/a_1108_47# VGND 0.129f
C16433 _310_/a_1283_21# VGND 0.291f
C16434 _310_/a_543_47# VGND 0.179f
C16435 _310_/a_761_289# VGND 0.124f
C16436 _310_/a_193_47# VGND 0.28f
C16437 _310_/a_27_47# VGND 0.542f
C16438 clknet_2_3__leaf_clk VGND 2.7f
C16439 clkbuf_2_3__f_clk/a_110_47# VGND 1.73f
C16440 _077_ VGND 0.111f
C16441 _208_/a_439_47# VGND 2.66e-19
C16442 _208_/a_218_47# VGND 8.02e-20
C16443 _208_/a_535_374# VGND 6.93e-19
C16444 _208_/a_218_374# VGND -1.61e-19
C16445 _208_/a_505_21# VGND 0.269f
C16446 _208_/a_76_199# VGND 0.151f
C16447 net14 VGND 1.4f
C16448 _011_ VGND 0.204f
C16449 _086_ VGND 0.122f
C16450 _225_/a_109_297# VGND -8.62e-19
C16451 _156_/a_27_47# VGND 0.274f
C16452 net26 VGND 3.2f
C16453 _311_/a_1462_47# VGND -8.05e-19
C16454 _311_/a_1217_47# VGND -4.08e-19
C16455 _311_/a_805_47# VGND -4.94e-19
C16456 _311_/a_639_47# VGND -0.00108f
C16457 _311_/a_1270_413# VGND 8.96e-20
C16458 _311_/a_651_413# VGND 0.00796f
C16459 _311_/a_448_47# VGND 0.0118f
C16460 _311_/a_1108_47# VGND 0.136f
C16461 _311_/a_1283_21# VGND 0.299f
C16462 _311_/a_543_47# VGND 0.176f
C16463 _311_/a_761_289# VGND 0.135f
C16464 _311_/a_193_47# VGND 0.311f
C16465 _311_/a_27_47# VGND 0.438f
C16466 _242_/a_297_47# VGND 0.0343f
C16467 _242_/a_382_297# VGND -5.32e-19
C16468 _242_/a_79_21# VGND 0.173f
C16469 net32 VGND 0.579f
C16470 _173_/a_27_47# VGND 0.213f
C16471 _190_/a_655_47# VGND 0.0277f
C16472 _190_/a_465_47# VGND 0.0109f
C16473 _190_/a_215_47# VGND 0.0163f
C16474 _190_/a_27_47# VGND 0.298f
C16475 _209_/a_27_47# VGND 0.45f
C16476 _075_ VGND 0.693f
C16477 _062_ VGND 1.34f
C16478 _226_/a_303_47# VGND -4.73e-19
C16479 _226_/a_197_47# VGND -5.42e-19
C16480 _226_/a_109_47# VGND -6.07e-19
C16481 _226_/a_27_47# VGND 0.158f
C16482 net20 VGND 1.22f
C16483 wire42/a_75_212# VGND 0.246f
C16484 _312_/a_1462_47# VGND 3.58e-19
C16485 _312_/a_1217_47# VGND 1.86e-19
C16486 _312_/a_805_47# VGND 5.48e-19
C16487 _312_/a_639_47# VGND 0.00114f
C16488 _312_/a_1270_413# VGND 1.66e-19
C16489 _312_/a_651_413# VGND 0.0118f
C16490 _312_/a_448_47# VGND 0.0207f
C16491 _312_/a_1108_47# VGND 0.158f
C16492 _312_/a_1283_21# VGND 0.324f
C16493 _312_/a_543_47# VGND 0.19f
C16494 _312_/a_761_289# VGND 0.148f
C16495 _312_/a_193_47# VGND 0.34f
C16496 _312_/a_27_47# VGND 0.561f
C16497 net55 VGND 0.859f
C16498 _096_ VGND 0.443f
C16499 _100_ VGND 0.216f
C16500 _243_/a_373_47# VGND -8.09e-19
C16501 _243_/a_109_47# VGND -0.00164f
C16502 _243_/a_109_297# VGND -6.92e-19
C16503 _243_/a_27_297# VGND 0.177f
C16504 net37 VGND 0.512f
C16505 _063_ VGND 1.25f
C16506 _191_/a_27_297# VGND 0.0593f
C16507 _260_/a_584_47# VGND -0.00127f
C16508 _260_/a_346_47# VGND -0.00146f
C16509 _260_/a_256_47# VGND -0.00132f
C16510 _260_/a_250_297# VGND 0.0356f
C16511 _260_/a_93_21# VGND 0.137f
C16512 _227_/a_368_53# VGND -5.8e-19
C16513 _227_/a_296_53# VGND -1.21e-19
C16514 _227_/a_209_311# VGND 0.126f
C16515 _227_/a_109_93# VGND 0.145f
C16516 _158_/a_150_297# VGND 4.75e-20
C16517 _158_/a_68_297# VGND 0.181f
C16518 _010_ VGND 0.344f
C16519 _313_/a_1462_47# VGND -8.44e-19
C16520 _313_/a_1217_47# VGND -4.41e-19
C16521 _313_/a_805_47# VGND -5.33e-19
C16522 _313_/a_639_47# VGND -0.00116f
C16523 _313_/a_1270_413# VGND 1.18e-19
C16524 _313_/a_651_413# VGND 0.00836f
C16525 _313_/a_448_47# VGND 0.0138f
C16526 _313_/a_1108_47# VGND 0.139f
C16527 _313_/a_1283_21# VGND 0.3f
C16528 _313_/a_543_47# VGND 0.162f
C16529 _313_/a_761_289# VGND 0.122f
C16530 _313_/a_193_47# VGND 0.319f
C16531 _313_/a_27_47# VGND 0.387f
C16532 net51 VGND 0.788f
C16533 _244_/a_27_297# VGND 0.0595f
C16534 _175_/a_150_297# VGND 1.23e-19
C16535 _175_/a_68_297# VGND 0.174f
C16536 net46 VGND 4.5f
C16537 _027_ VGND 0.244f
C16538 _330_/a_1217_47# VGND 6.9e-20
C16539 _330_/a_805_47# VGND -4.9e-19
C16540 _330_/a_639_47# VGND -0.00109f
C16541 _330_/a_1270_413# VGND 2.57e-20
C16542 _330_/a_651_413# VGND 0.00807f
C16543 _330_/a_448_47# VGND 0.0102f
C16544 _330_/a_1108_47# VGND 0.136f
C16545 _330_/a_1283_21# VGND 0.3f
C16546 _330_/a_543_47# VGND 0.163f
C16547 _330_/a_761_289# VGND 0.132f
C16548 _330_/a_193_47# VGND 0.275f
C16549 _330_/a_27_47# VGND 0.383f
C16550 cal_count\[3\] VGND 0.667f
C16551 _261_/a_113_47# VGND -7.28e-22
C16552 _065_ VGND 2.46f
C16553 _192_/a_639_47# VGND -5.47e-19
C16554 _192_/a_548_47# VGND -7.23e-19
C16555 _192_/a_476_47# VGND -7.49e-19
C16556 _192_/a_505_280# VGND 0.185f
C16557 _192_/a_27_47# VGND 0.197f
C16558 _192_/a_174_21# VGND 0.197f
C16559 clone1/a_27_47# VGND 0.281f
C16560 _052_ VGND 0.947f
C16561 _088_ VGND 0.189f
C16562 _228_/a_297_47# VGND 0.0693f
C16563 _228_/a_382_297# VGND -5.55e-19
C16564 _228_/a_79_21# VGND 0.183f
C16565 net21 VGND 0.706f
C16566 _046_ VGND 0.221f
C16567 _159_/a_27_47# VGND 0.237f
C16568 _314_/a_1217_47# VGND 9.94e-20
C16569 _314_/a_805_47# VGND 2.56e-19
C16570 _314_/a_639_47# VGND 4.79e-19
C16571 _314_/a_1270_413# VGND 1.18e-19
C16572 _314_/a_651_413# VGND 0.00755f
C16573 _314_/a_448_47# VGND 0.0176f
C16574 _314_/a_1108_47# VGND 0.161f
C16575 _314_/a_1283_21# VGND 0.351f
C16576 _314_/a_543_47# VGND 0.166f
C16577 _314_/a_761_289# VGND 0.127f
C16578 _314_/a_193_47# VGND 0.295f
C16579 _314_/a_27_47# VGND 0.496f
C16580 _016_ VGND 0.243f
C16581 net52 VGND 2.4f
C16582 _101_ VGND 1.98f
C16583 _245_/a_373_47# VGND 3.81e-19
C16584 _245_/a_109_47# VGND -0.00142f
C16585 _245_/a_109_297# VGND 0.0021f
C16586 _245_/a_27_297# VGND 0.2f
C16587 net33 VGND 1.11f
C16588 _056_ VGND 0.219f
C16589 _176_/a_27_47# VGND 0.267f
C16590 trim_mask\[4\] VGND 2.57f
C16591 _028_ VGND 0.279f
C16592 clknet_2_2__leaf_clk VGND 3.81f
C16593 _331_/a_1462_47# VGND 6.1e-19
C16594 _331_/a_1217_47# VGND 2.49e-19
C16595 _331_/a_805_47# VGND 6.94e-19
C16596 _331_/a_639_47# VGND 0.00137f
C16597 _331_/a_1270_413# VGND 1.07e-19
C16598 _331_/a_651_413# VGND 0.00785f
C16599 _331_/a_448_47# VGND 0.0175f
C16600 _331_/a_1108_47# VGND 0.166f
C16601 _331_/a_1283_21# VGND 0.337f
C16602 _331_/a_543_47# VGND 0.174f
C16603 _331_/a_761_289# VGND 0.128f
C16604 _331_/a_193_47# VGND 0.306f
C16605 _331_/a_27_47# VGND 0.531f
C16606 _105_ VGND 0.267f
C16607 _262_/a_465_47# VGND -1.84e-19
C16608 _262_/a_193_297# VGND -0.00323f
C16609 _262_/a_109_297# VGND -0.00197f
C16610 _262_/a_27_47# VGND 0.237f
C16611 _193_/a_109_297# VGND -7.17e-19
C16612 _090_ VGND 0.475f
C16613 _089_ VGND 0.24f
C16614 _087_ VGND 0.444f
C16615 _229_/a_27_297# VGND 0.0588f
C16616 _315_/a_1270_413# VGND 2.91e-20
C16617 _315_/a_651_413# VGND 0.00515f
C16618 _315_/a_448_47# VGND 0.0142f
C16619 _315_/a_1108_47# VGND 0.156f
C16620 _315_/a_1283_21# VGND 0.338f
C16621 _315_/a_543_47# VGND 0.158f
C16622 _315_/a_761_289# VGND 0.121f
C16623 _315_/a_193_47# VGND 0.292f
C16624 _315_/a_27_47# VGND 0.554f
C16625 _017_ VGND 0.161f
C16626 mask\[2\] VGND 2.46f
C16627 _246_/a_373_47# VGND -8.76e-19
C16628 _246_/a_109_47# VGND -0.00113f
C16629 _246_/a_109_297# VGND 0.00601f
C16630 _246_/a_27_297# VGND 0.194f
C16631 net38 VGND 0.503f
C16632 _332_/a_1462_47# VGND -2.63e-20
C16633 _332_/a_1217_47# VGND -4.26e-19
C16634 _332_/a_1270_413# VGND 2.69e-19
C16635 _332_/a_651_413# VGND 0.00605f
C16636 _332_/a_448_47# VGND 0.0157f
C16637 _332_/a_1108_47# VGND 0.155f
C16638 _332_/a_1283_21# VGND 0.321f
C16639 _332_/a_543_47# VGND 0.18f
C16640 _332_/a_761_289# VGND 0.123f
C16641 _332_/a_193_47# VGND 0.312f
C16642 _332_/a_27_47# VGND 0.526f
C16643 _107_ VGND 1.56f
C16644 _263_/a_297_47# VGND 0.0661f
C16645 _263_/a_382_297# VGND -7.56e-19
C16646 _263_/a_79_21# VGND 0.14f
C16647 _067_ VGND 1.76f
C16648 _066_ VGND 0.276f
C16649 _194_/a_199_47# VGND 6.23e-20
C16650 _194_/a_113_297# VGND 0.0341f
C16651 _119_ VGND 0.3f
C16652 _280_/a_75_212# VGND 0.224f
C16653 _057_ VGND 1.06f
C16654 _178_/a_150_297# VGND -3.18e-19
C16655 _178_/a_68_297# VGND 0.172f
C16656 _013_ VGND 0.337f
C16657 _316_/a_1462_47# VGND -7.5e-19
C16658 _316_/a_1217_47# VGND -3.77e-19
C16659 _316_/a_805_47# VGND 7.04e-19
C16660 _316_/a_639_47# VGND 4.52e-19
C16661 _316_/a_1270_413# VGND 1.17e-19
C16662 _316_/a_651_413# VGND 0.0147f
C16663 _316_/a_448_47# VGND 0.0124f
C16664 _316_/a_1108_47# VGND 0.139f
C16665 _316_/a_1283_21# VGND 0.313f
C16666 _316_/a_543_47# VGND 0.185f
C16667 _316_/a_761_289# VGND 0.141f
C16668 _316_/a_193_47# VGND 0.319f
C16669 _316_/a_27_47# VGND 0.418f
C16670 _018_ VGND 0.395f
C16671 _247_/a_373_47# VGND -0.00126f
C16672 _247_/a_109_47# VGND -0.00117f
C16673 _247_/a_109_297# VGND 5.82e-19
C16674 _247_/a_27_297# VGND 0.197f
C16675 _333_/a_1462_47# VGND 2.9e-19
C16676 _333_/a_1217_47# VGND 4.36e-19
C16677 _333_/a_805_47# VGND 5.23e-19
C16678 _333_/a_639_47# VGND 9.64e-19
C16679 _333_/a_1270_413# VGND 1.2e-19
C16680 _333_/a_651_413# VGND 0.00798f
C16681 _333_/a_448_47# VGND 0.0126f
C16682 _333_/a_1108_47# VGND 0.156f
C16683 _333_/a_1283_21# VGND 0.307f
C16684 _333_/a_543_47# VGND 0.173f
C16685 _333_/a_761_289# VGND 0.145f
C16686 _333_/a_193_47# VGND 0.304f
C16687 _333_/a_27_47# VGND 0.406f
C16688 _106_ VGND 0.769f
C16689 _264_/a_27_297# VGND 0.0559f
C16690 _068_ VGND 0.425f
C16691 _195_/a_439_47# VGND -2.31e-19
C16692 _195_/a_218_47# VGND -6.48e-19
C16693 _195_/a_535_374# VGND -3.69e-19
C16694 _195_/a_218_374# VGND -6.75e-19
C16695 _195_/a_505_21# VGND 0.251f
C16696 _195_/a_76_199# VGND 0.12f
C16697 _120_ VGND 0.244f
C16698 en_co_clk VGND 1.51f
C16699 _281_/a_253_47# VGND 0.0115f
C16700 _281_/a_337_297# VGND -0.00113f
C16701 _281_/a_253_297# VGND -9.14e-19
C16702 _281_/a_103_199# VGND 0.211f
C16703 clknet_0_clk VGND 3.97f
C16704 clkbuf_2_2__f_clk/a_110_47# VGND 1.71f
C16705 state\[1\] VGND 0.956f
C16706 net45 VGND 4.61f
C16707 _014_ VGND 0.587f
C16708 clknet_2_0__leaf_clk VGND 4.08f
C16709 _317_/a_1462_47# VGND 5.46e-19
C16710 _317_/a_1217_47# VGND 1.2e-19
C16711 _317_/a_805_47# VGND 7.93e-19
C16712 _317_/a_639_47# VGND 0.00364f
C16713 _317_/a_1270_413# VGND 1.01e-19
C16714 _317_/a_651_413# VGND 0.0114f
C16715 _317_/a_448_47# VGND 0.0243f
C16716 _317_/a_1108_47# VGND 0.165f
C16717 _317_/a_1283_21# VGND 0.333f
C16718 _317_/a_543_47# VGND 0.2f
C16719 _317_/a_761_289# VGND 0.144f
C16720 _317_/a_193_47# VGND 0.332f
C16721 _317_/a_27_47# VGND 0.568f
C16722 mask\[4\] VGND 2.78f
C16723 _248_/a_373_47# VGND -8.12e-19
C16724 _248_/a_109_47# VGND -0.00146f
C16725 _248_/a_109_297# VGND 2.85e-19
C16726 _248_/a_27_297# VGND 0.18f
C16727 net34 VGND 1.61f
C16728 _179_/a_27_47# VGND 0.25f
C16729 _109_ VGND 0.166f
C16730 trim_val\[0\] VGND 0.946f
C16731 _265_/a_384_47# VGND -3.83e-19
C16732 _265_/a_299_297# VGND 0.0362f
C16733 _265_/a_81_21# VGND 0.127f
C16734 _031_ VGND 0.258f
C16735 _334_/a_1462_47# VGND 0.00184f
C16736 _334_/a_1217_47# VGND 5.95e-20
C16737 _334_/a_1270_413# VGND 2.69e-19
C16738 _334_/a_651_413# VGND 0.00733f
C16739 _334_/a_448_47# VGND 0.0139f
C16740 _334_/a_1108_47# VGND 0.171f
C16741 _334_/a_1283_21# VGND 0.336f
C16742 _334_/a_543_47# VGND 0.168f
C16743 _334_/a_761_289# VGND 0.139f
C16744 _334_/a_193_47# VGND 0.31f
C16745 _334_/a_27_47# VGND 0.484f
C16746 _121_ VGND 0.199f
C16747 _282_/a_150_297# VGND -1.98e-19
C16748 _282_/a_68_297# VGND 0.152f
C16749 state\[2\] VGND 0.983f
C16750 _015_ VGND 0.457f
C16751 _318_/a_651_413# VGND 0.00472f
C16752 _318_/a_448_47# VGND 0.0157f
C16753 _318_/a_1108_47# VGND 0.156f
C16754 _318_/a_1283_21# VGND 0.336f
C16755 _318_/a_543_47# VGND 0.175f
C16756 _318_/a_761_289# VGND 0.123f
C16757 _318_/a_193_47# VGND 0.311f
C16758 _318_/a_27_47# VGND 0.567f
C16759 _020_ VGND 0.975f
C16760 mask\[5\] VGND 1.02f
C16761 _249_/a_373_47# VGND 0.00141f
C16762 _249_/a_109_47# VGND -0.00111f
C16763 _249_/a_109_297# VGND 5.35e-19
C16764 _249_/a_27_297# VGND 0.229f
C16765 _032_ VGND 0.439f
C16766 _335_/a_1462_47# VGND -8.62e-19
C16767 _335_/a_1217_47# VGND -4.26e-19
C16768 _335_/a_805_47# VGND -5.87e-19
C16769 _335_/a_639_47# VGND -0.00109f
C16770 _335_/a_1270_413# VGND 6.88e-20
C16771 _335_/a_651_413# VGND 0.0101f
C16772 _335_/a_448_47# VGND 0.014f
C16773 _335_/a_1108_47# VGND 0.136f
C16774 _335_/a_1283_21# VGND 0.307f
C16775 _335_/a_543_47# VGND 0.166f
C16776 _335_/a_761_289# VGND 0.138f
C16777 _335_/a_193_47# VGND 0.301f
C16778 _335_/a_27_47# VGND 0.525f
C16779 _266_/a_150_297# VGND -4.61e-19
C16780 _266_/a_68_297# VGND 0.156f
C16781 _069_ VGND 0.139f
C16782 _197_/a_199_47# VGND -4.12e-19
C16783 _197_/a_113_297# VGND 0.0356f
C16784 _034_ VGND 0.277f
C16785 _283_/a_75_212# VGND 0.228f
C16786 _319_/a_1462_47# VGND -8.2e-19
C16787 _319_/a_1217_47# VGND -4.2e-19
C16788 _319_/a_805_47# VGND -5.23e-19
C16789 _319_/a_639_47# VGND -0.00113f
C16790 _319_/a_1270_413# VGND 6.7e-20
C16791 _319_/a_651_413# VGND 0.00642f
C16792 _319_/a_448_47# VGND 0.01f
C16793 _319_/a_1108_47# VGND 0.133f
C16794 _319_/a_1283_21# VGND 0.297f
C16795 _319_/a_543_47# VGND 0.155f
C16796 _319_/a_761_289# VGND 0.118f
C16797 _319_/a_193_47# VGND 0.273f
C16798 _319_/a_27_47# VGND 0.413f
C16799 _033_ VGND 0.221f
C16800 _336_/a_1462_47# VGND -9.48e-19
C16801 _336_/a_1217_47# VGND -5.03e-19
C16802 _336_/a_805_47# VGND -6.6e-19
C16803 _336_/a_639_47# VGND -0.00145f
C16804 _336_/a_651_413# VGND 0.00587f
C16805 _336_/a_448_47# VGND 0.00856f
C16806 _336_/a_1108_47# VGND 0.129f
C16807 _336_/a_1283_21# VGND 0.287f
C16808 _336_/a_543_47# VGND 0.153f
C16809 _336_/a_761_289# VGND 0.117f
C16810 _336_/a_193_47# VGND 0.269f
C16811 _336_/a_27_47# VGND 0.395f
C16812 _267_/a_145_75# VGND -0.0013f
C16813 _267_/a_59_75# VGND 0.163f
C16814 _198_/a_181_47# VGND -4.01e-19
C16815 _198_/a_109_47# VGND -4.03e-19
C16816 _198_/a_27_47# VGND 0.18f
C16817 _122_ VGND 1.84f
C16818 _284_/a_150_297# VGND -1.79e-19
C16819 _284_/a_68_297# VGND 0.169f
C16820 net44 VGND 2.94f
C16821 _337_/a_1462_47# VGND 2.63e-19
C16822 _337_/a_1217_47# VGND 1.16e-19
C16823 _337_/a_805_47# VGND -5.45e-19
C16824 _337_/a_639_47# VGND -0.00123f
C16825 _337_/a_1270_413# VGND 5.36e-20
C16826 _337_/a_651_413# VGND 0.00719f
C16827 _337_/a_448_47# VGND 0.011f
C16828 _337_/a_1108_47# VGND 0.16f
C16829 _337_/a_1283_21# VGND 0.332f
C16830 _337_/a_543_47# VGND 0.159f
C16831 _337_/a_761_289# VGND 0.138f
C16832 _337_/a_193_47# VGND 0.303f
C16833 _337_/a_27_47# VGND 0.375f
C16834 _029_ VGND 0.442f
C16835 _111_ VGND 0.46f
C16836 _268_/a_75_212# VGND 0.261f
C16837 _001_ VGND 0.586f
C16838 _199_/a_193_297# VGND -6.63e-19
C16839 _199_/a_109_297# VGND -5.59e-19
C16840 _123_ VGND 0.583f
C16841 _285_/a_113_47# VGND 1.85e-19
C16842 _338_/a_1296_47# VGND -4.76e-19
C16843 _338_/a_1224_47# VGND -4.71e-19
C16844 _338_/a_1056_47# VGND -4.53e-19
C16845 _338_/a_796_47# VGND -4.19e-19
C16846 _338_/a_586_47# VGND -8.82e-19
C16847 _338_/a_1140_413# VGND 3.5e-19
C16848 _338_/a_956_413# VGND 5.62e-19
C16849 _338_/a_562_413# VGND 5.72e-19
C16850 _338_/a_381_47# VGND 0.0336f
C16851 _338_/a_1602_47# VGND 0.146f
C16852 _338_/a_1032_413# VGND 0.345f
C16853 _338_/a_1182_261# VGND 0.145f
C16854 _338_/a_476_47# VGND 0.322f
C16855 _338_/a_652_21# VGND 0.136f
C16856 _338_/a_193_47# VGND 0.228f
C16857 _338_/a_27_47# VGND 0.489f
C16858 _112_ VGND 0.28f
C16859 net49 VGND 0.422f
C16860 trim_mask\[1\] VGND 1.48f
C16861 trim_val\[1\] VGND 0.362f
C16862 _269_/a_384_47# VGND 9.75e-20
C16863 _269_/a_299_297# VGND 0.0358f
C16864 _269_/a_81_21# VGND 0.135f
C16865 _040_ VGND 1.28f
C16866 _140_/a_150_297# VGND -4.61e-19
C16867 _140_/a_68_297# VGND 0.149f
C16868 cal_count\[0\] VGND 1.19f
C16869 _124_ VGND 0.177f
C16870 _286_/a_439_47# VGND -2.64e-19
C16871 _286_/a_218_47# VGND -2.58e-19
C16872 _286_/a_535_374# VGND -1.67e-19
C16873 _286_/a_218_374# VGND -8.87e-20
C16874 _286_/a_505_21# VGND 0.253f
C16875 _286_/a_76_199# VGND 0.146f
C16876 _339_/a_1296_47# VGND -4.9e-19
C16877 _339_/a_1224_47# VGND -4.99e-19
C16878 _339_/a_1056_47# VGND -4.93e-19
C16879 _339_/a_796_47# VGND -4.72e-19
C16880 _339_/a_586_47# VGND -8.66e-19
C16881 _339_/a_1140_413# VGND 6.77e-20
C16882 _339_/a_956_413# VGND 1.87e-19
C16883 _339_/a_562_413# VGND 1.7e-19
C16884 _339_/a_381_47# VGND 0.0198f
C16885 _339_/a_1602_47# VGND 0.116f
C16886 _339_/a_1032_413# VGND 0.302f
C16887 _339_/a_1182_261# VGND 0.124f
C16888 _339_/a_476_47# VGND 0.298f
C16889 _339_/a_652_21# VGND 0.135f
C16890 _339_/a_193_47# VGND 0.199f
C16891 _339_/a_27_47# VGND 0.447f
C16892 _078_ VGND 2.56f
C16893 mask\[0\] VGND 3.46f
C16894 net22 VGND 1.06f
C16895 _210_/a_199_47# VGND -1.67e-19
C16896 _210_/a_113_297# VGND 0.0354f
C16897 _141_/a_27_47# VGND 0.259f
C16898 _035_ VGND 0.427f
C16899 _287_/a_75_212# VGND 0.226f
C16900 _004_ VGND 0.585f
C16901 _079_ VGND 0.363f
C16902 _211_/a_109_297# VGND -8.64e-19
C16903 net7 VGND 0.305f
C16904 net15 VGND 1.43f
C16905 net4 VGND 2.51f
C16906 rstn VGND 0.359f
C16907 input4/a_27_47# VGND 0.276f
C16908 clknet_2_1__leaf_clk VGND 4f
C16909 clkbuf_2_1__f_clk/a_110_47# VGND 1.69f
C16910 _125_ VGND 0.937f
C16911 _288_/a_145_75# VGND 2.67e-19
C16912 _288_/a_59_75# VGND 0.214f
C16913 fanout47/a_27_47# VGND 0.425f
C16914 mask\[1\] VGND 1.27f
C16915 _212_/a_199_47# VGND -4.91e-19
C16916 _212_/a_113_297# VGND 0.0287f
C16917 _041_ VGND 4.65f
C16918 _143_/a_150_297# VGND -2.16e-19
C16919 _143_/a_68_297# VGND 0.168f
C16920 net3 VGND 1.07f
C16921 en VGND 0.446f
C16922 input3/a_75_212# VGND 0.267f
C16923 _126_ VGND 0.541f
C16924 _289_/a_150_297# VGND -1.98e-19
C16925 _289_/a_68_297# VGND 0.17f
C16926 fanout46/a_27_47# VGND 0.557f
C16927 _080_ VGND 0.0999f
C16928 _213_/a_109_297# VGND -0.00128f
C16929 _144_/a_27_47# VGND 0.211f
C16930 comp VGND 0.28f
C16931 input2/a_27_47# VGND 0.38f
C16932 _091_ VGND 0.221f
C16933 _230_/a_145_75# VGND -0.00114f
C16934 _230_/a_59_75# VGND 0.166f
C16935 _161_/a_150_297# VGND -2.91e-19
C16936 _161_/a_68_297# VGND 0.148f
C16937 fanout45/a_27_47# VGND 0.33f
C16938 _214_/a_199_47# VGND 9.48e-19
C16939 _214_/a_113_297# VGND 0.0406f
C16940 net16 VGND 2.31f
C16941 net1 VGND 0.339f
C16942 cal VGND 0.542f
C16943 input1/a_75_212# VGND 0.264f
C16944 _135_ VGND 0.205f
C16945 net2 VGND 6.36f
C16946 _300_/a_285_47# VGND 0.0151f
C16947 _300_/a_129_47# VGND 2.25e-19
C16948 _300_/a_377_297# VGND -8.33e-19
C16949 _300_/a_47_47# VGND 0.243f
C16950 _231_/a_161_47# VGND 0.622f
C16951 _047_ VGND 0.311f
C16952 _162_/a_27_47# VGND 0.242f
C16953 fanout44/a_27_47# VGND 0.333f
C16954 _006_ VGND 0.233f
C16955 _081_ VGND 0.514f
C16956 _215_/a_109_297# VGND -1.36e-19
C16957 _042_ VGND 0.834f
C16958 _146_/a_150_297# VGND -2.84e-19
C16959 _146_/a_68_297# VGND 0.161f
C16960 _134_ VGND 0.41f
C16961 _301_/a_285_47# VGND 0.0149f
C16962 _301_/a_129_47# VGND 1.79e-19
C16963 _301_/a_377_297# VGND -0.00125f
C16964 _301_/a_47_47# VGND 0.24f
C16965 _232_/a_304_297# VGND -9.51e-19
C16966 _232_/a_220_297# VGND -0.00123f
C16967 _232_/a_114_297# VGND -0.00201f
C16968 _232_/a_32_297# VGND 0.426f
C16969 net36 VGND 0.162f
C16970 fanout43/a_27_47# VGND 0.53f
C16971 net39 VGND 0.532f
C16972 ctlp[5] VGND 0.524f
C16973 output19/a_27_47# VGND 0.332f
C16974 _082_ VGND 0.208f
C16975 mask\[3\] VGND 1.25f
C16976 net25 VGND 0.959f
C16977 _216_/a_199_47# VGND 7.32e-21
C16978 _216_/a_113_297# VGND 0.0325f
C16979 net17 VGND 1.22f
C16980 _147_/a_27_47# VGND 0.281f
C16981 _038_ VGND 0.451f
C16982 _136_ VGND 1.18f
C16983 _302_/a_373_47# VGND -0.00113f
C16984 _302_/a_109_47# VGND -0.00138f
C16985 _302_/a_109_297# VGND 0.00305f
C16986 _302_/a_27_297# VGND 0.188f
C16987 _012_ VGND 0.356f
C16988 _093_ VGND 0.623f
C16989 calibrate VGND 0.855f
C16990 _074_ VGND 4.23f
C16991 _233_/a_373_47# VGND 2.17e-19
C16992 _233_/a_109_47# VGND -0.00188f
C16993 _233_/a_109_297# VGND -1.69e-19
C16994 _233_/a_27_297# VGND 0.203f
C16995 _048_ VGND 3.31f
C16996 _164_/a_161_47# VGND 0.596f
C16997 _021_ VGND 0.435f
C16998 _250_/a_373_47# VGND 2.78e-19
C16999 _250_/a_109_47# VGND -0.00168f
C17000 _250_/a_109_297# VGND 1.7e-20
C17001 _250_/a_27_297# VGND 0.186f
C17002 _058_ VGND 1.55f
C17003 _181_/a_150_297# VGND -1.92e-19
C17004 _181_/a_68_297# VGND 0.165f
C17005 ctlp[4] VGND 0.55f
C17006 output18/a_27_47# VGND 0.337f
C17007 result[7] VGND 0.395f
C17008 output29/a_27_47# VGND 0.33f
C17009 _007_ VGND 0.235f
C17010 _217_/a_109_297# VGND -8.91e-19
C17011 _000_ VGND 0.547f
C17012 _303_/a_1462_47# VGND 2.06e-19
C17013 _303_/a_1217_47# VGND 9.86e-20
C17014 _303_/a_805_47# VGND 2.55e-19
C17015 _303_/a_639_47# VGND 5.19e-19
C17016 _303_/a_1270_413# VGND 5.06e-20
C17017 _303_/a_651_413# VGND 0.00584f
C17018 _303_/a_448_47# VGND 0.0175f
C17019 _303_/a_1108_47# VGND 0.155f
C17020 _303_/a_1283_21# VGND 0.422f
C17021 _303_/a_543_47# VGND 0.162f
C17022 _303_/a_761_289# VGND 0.128f
C17023 _303_/a_193_47# VGND 0.3f
C17024 _303_/a_27_47# VGND 0.548f
C17025 _234_/a_109_297# VGND -3.13e-19
C17026 _320_/a_1217_47# VGND -5.03e-19
C17027 _320_/a_805_47# VGND -7.16e-19
C17028 _320_/a_639_47# VGND -0.00152f
C17029 _320_/a_1270_413# VGND 5.39e-20
C17030 _320_/a_651_413# VGND 0.00834f
C17031 _320_/a_448_47# VGND 0.0136f
C17032 _320_/a_1108_47# VGND 0.147f
C17033 _320_/a_1283_21# VGND 0.303f
C17034 _320_/a_543_47# VGND 0.173f
C17035 _320_/a_761_289# VGND 0.133f
C17036 _320_/a_193_47# VGND 0.293f
C17037 _320_/a_27_47# VGND 0.377f
C17038 _022_ VGND 0.156f
C17039 mask\[6\] VGND 2.71f
C17040 _251_/a_373_47# VGND -0.00105f
C17041 _251_/a_109_47# VGND 5.56e-19
C17042 _251_/a_109_297# VGND 0.0046f
C17043 _251_/a_27_297# VGND 0.196f
C17044 net35 VGND 0.545f
C17045 _182_/a_27_47# VGND 0.245f
C17046 clkbuf_2_0__f_clk/a_110_47# VGND 1.76f
C17047 ctlp[3] VGND 0.572f
C17048 output17/a_27_47# VGND 0.314f
C17049 result[6] VGND 0.381f
C17050 net28 VGND 2.19f
C17051 output28/a_27_47# VGND 0.563f
C17052 trimb[3] VGND 0.285f
C17053 output39/a_27_47# VGND 0.578f
C17054 _083_ VGND 0.314f
C17055 _218_/a_199_47# VGND -4.56e-19
C17056 _218_/a_113_297# VGND 0.0298f
C17057 _043_ VGND 0.856f
C17058 _149_/a_150_297# VGND -3.44e-19
C17059 _149_/a_68_297# VGND 0.158f
C17060 _050_ VGND 1.51f
C17061 _166_/a_161_47# VGND 0.669f
C17062 net47 VGND 3.49f
C17063 _304_/a_1462_47# VGND 0.00184f
C17064 _304_/a_1217_47# VGND 1.88e-19
C17065 _304_/a_805_47# VGND 4.35e-19
C17066 _304_/a_639_47# VGND 7.64e-19
C17067 _304_/a_1270_413# VGND 1e-19
C17068 _304_/a_651_413# VGND 0.00897f
C17069 _304_/a_448_47# VGND 0.0156f
C17070 _304_/a_1108_47# VGND 0.172f
C17071 _304_/a_1283_21# VGND 0.349f
C17072 _304_/a_543_47# VGND 0.172f
C17073 _304_/a_761_289# VGND 0.139f
C17074 _304_/a_193_47# VGND 0.297f
C17075 _304_/a_27_47# VGND 0.495f
C17076 _094_ VGND 1.14f
C17077 _235_/a_297_47# VGND 0.0202f
C17078 _235_/a_382_297# VGND -8.23e-19
C17079 _235_/a_79_21# VGND 0.14f
C17080 _321_/a_1462_47# VGND 2.59e-19
C17081 _321_/a_1217_47# VGND -4.18e-19
C17082 _321_/a_805_47# VGND -5.21e-19
C17083 _321_/a_639_47# VGND -0.00119f
C17084 _321_/a_1270_413# VGND 8.16e-20
C17085 _321_/a_651_413# VGND 0.00904f
C17086 _321_/a_448_47# VGND 0.0094f
C17087 _321_/a_1108_47# VGND 0.15f
C17088 _321_/a_1283_21# VGND 0.301f
C17089 _321_/a_543_47# VGND 0.174f
C17090 _321_/a_761_289# VGND 0.134f
C17091 _321_/a_193_47# VGND 0.292f
C17092 _321_/a_27_47# VGND 0.38f
C17093 clk VGND 4.02f
C17094 clkbuf_0_clk/a_110_47# VGND 1.75f
C17095 ctlp[2] VGND 0.52f
C17096 output16/a_27_47# VGND 0.359f
C17097 result[5] VGND 0.274f
C17098 net27 VGND 4.14f
C17099 output27/a_27_47# VGND 0.334f
C17100 trimb[2] VGND 0.28f
C17101 output38/a_27_47# VGND 0.644f
C17102 _008_ VGND 0.181f
C17103 _219_/a_109_297# VGND -0.00126f
C17104 _002_ VGND 0.808f
C17105 _305_/a_1462_47# VGND 1.03e-19
C17106 _305_/a_1217_47# VGND -4.97e-19
C17107 _305_/a_805_47# VGND -6.53e-19
C17108 _305_/a_639_47# VGND -0.00139f
C17109 _305_/a_1270_413# VGND 3.27e-20
C17110 _305_/a_651_413# VGND 0.00576f
C17111 _305_/a_448_47# VGND 0.00947f
C17112 _305_/a_1108_47# VGND 0.135f
C17113 _305_/a_1283_21# VGND 0.298f
C17114 _305_/a_543_47# VGND 0.158f
C17115 _305_/a_761_289# VGND 0.117f
C17116 _305_/a_193_47# VGND 0.276f
C17117 _305_/a_27_47# VGND 0.448f
C17118 _236_/a_109_297# VGND -0.00122f
C17119 _051_ VGND 3.28f
C17120 _167_/a_161_47# VGND 0.649f
C17121 _023_ VGND 0.242f
C17122 _102_ VGND 0.344f
C17123 mask\[7\] VGND 1.96f
C17124 _253_/a_384_47# VGND 4.62e-20
C17125 _253_/a_299_297# VGND 0.0327f
C17126 _253_/a_81_21# VGND 0.143f
C17127 _019_ VGND 0.172f
C17128 _322_/a_1217_47# VGND -4.41e-19
C17129 _322_/a_805_47# VGND 2.55e-19
C17130 _322_/a_639_47# VGND 5.19e-19
C17131 _322_/a_1270_413# VGND 5.06e-20
C17132 _322_/a_651_413# VGND 0.00562f
C17133 _322_/a_448_47# VGND 0.0153f
C17134 _322_/a_1108_47# VGND 0.135f
C17135 _322_/a_1283_21# VGND 0.304f
C17136 _322_/a_543_47# VGND 0.178f
C17137 _322_/a_761_289# VGND 0.122f
C17138 _322_/a_193_47# VGND 0.287f
C17139 _322_/a_27_47# VGND 0.539f
C17140 _270_/a_145_75# VGND 1.46e-20
C17141 _270_/a_59_75# VGND 0.212f
C17142 ctlp[1] VGND 0.516f
C17143 output15/a_27_47# VGND 0.33f
C17144 result[4] VGND 0.233f
C17145 output26/a_27_47# VGND 0.333f
C17146 trimb[1] VGND 0.202f
C17147 output37/a_27_47# VGND 0.589f
C17148 _306_/a_1462_47# VGND 3.4e-19
C17149 _306_/a_1217_47# VGND 1.77e-19
C17150 _306_/a_805_47# VGND 0.00144f
C17151 _306_/a_639_47# VGND 0.00461f
C17152 _306_/a_1270_413# VGND 9.17e-20
C17153 _306_/a_651_413# VGND 0.0132f
C17154 _306_/a_448_47# VGND 0.0177f
C17155 _306_/a_1108_47# VGND 0.146f
C17156 _306_/a_1283_21# VGND 0.303f
C17157 _306_/a_543_47# VGND 0.191f
C17158 _306_/a_761_289# VGND 0.139f
C17159 _306_/a_193_47# VGND 0.319f
C17160 _306_/a_27_47# VGND 0.533f
C17161 _237_/a_439_47# VGND -5.32e-19
C17162 _237_/a_218_47# VGND -6.39e-19
C17163 _237_/a_535_374# VGND -2.11e-19
C17164 _237_/a_218_374# VGND -2.89e-19
C17165 _237_/a_505_21# VGND 0.302f
C17166 _237_/a_76_199# VGND 0.132f
C17167 _168_/a_297_47# VGND 4.39e-19
C17168 _168_/a_207_413# VGND 0.141f
C17169 _168_/a_27_413# VGND 0.206f
C17170 _323_/a_1462_47# VGND -8.82e-19
C17171 _323_/a_1217_47# VGND 6.19e-20
C17172 _323_/a_805_47# VGND 1.62e-19
C17173 _323_/a_639_47# VGND 3.29e-19
C17174 _323_/a_1270_413# VGND 2.27e-20
C17175 _323_/a_651_413# VGND 0.00734f
C17176 _323_/a_448_47# VGND 0.0153f
C17177 _323_/a_1108_47# VGND 0.156f
C17178 _323_/a_1283_21# VGND 0.297f
C17179 _323_/a_543_47# VGND 0.178f
C17180 _323_/a_761_289# VGND 0.138f
C17181 _323_/a_193_47# VGND 0.299f
C17182 _323_/a_27_47# VGND 0.503f
C17183 net42 VGND 0.286f
C17184 _254_/a_109_297# VGND -7.75e-19
C17185 _060_ VGND 0.822f
C17186 net54 VGND 0.742f
C17187 _185_/a_150_297# VGND -3.26e-19
C17188 _185_/a_68_297# VGND 0.158f
C17189 _037_ VGND 0.325f
C17190 _340_/a_381_47# VGND 0.0225f
C17191 _340_/a_1602_47# VGND 0.135f
C17192 _340_/a_1032_413# VGND 0.306f
C17193 _340_/a_1182_261# VGND 0.128f
C17194 _340_/a_476_47# VGND 0.309f
C17195 _340_/a_652_21# VGND 0.136f
C17196 _340_/a_193_47# VGND 0.34f
C17197 _340_/a_27_47# VGND 0.47f
C17198 _030_ VGND 0.162f
C17199 _113_ VGND 0.348f
C17200 _271_/a_75_212# VGND 0.218f
C17201 ctlp[0] VGND 0.491f
C17202 output14/a_27_47# VGND 0.591f
C17203 result[3] VGND 0.243f
C17204 output25/a_27_47# VGND 0.304f
C17205 trimb[0] VGND 0.244f
C17206 output36/a_27_47# VGND 0.624f
C17207 _307_/a_1462_47# VGND 2.63e-19
C17208 _307_/a_1217_47# VGND 5.76e-20
C17209 _307_/a_805_47# VGND 3.4e-19
C17210 _307_/a_639_47# VGND 6.34e-19
C17211 _307_/a_1270_413# VGND 3.88e-20
C17212 _307_/a_651_413# VGND 0.00839f
C17213 _307_/a_448_47# VGND 0.0175f
C17214 _307_/a_1108_47# VGND 0.155f
C17215 _307_/a_1283_21# VGND 0.317f
C17216 _307_/a_543_47# VGND 0.173f
C17217 _307_/a_761_289# VGND 0.139f
C17218 _307_/a_193_47# VGND 0.3f
C17219 _307_/a_27_47# VGND 0.549f
C17220 _097_ VGND 0.399f
C17221 _238_/a_75_212# VGND 0.24f
C17222 _053_ VGND 3.28f
C17223 state\[0\] VGND 0.812f
C17224 _169_/a_373_53# VGND -3.53e-19
C17225 _169_/a_301_53# VGND -1.2e-19
C17226 _169_/a_109_53# VGND 0.146f
C17227 _169_/a_215_311# VGND 0.239f
C17228 _324_/a_1462_47# VGND 1.11e-19
C17229 _324_/a_1217_47# VGND 6.49e-20
C17230 _324_/a_805_47# VGND 2.34e-19
C17231 _324_/a_639_47# VGND 5.12e-19
C17232 _324_/a_1270_413# VGND 3.52e-20
C17233 _324_/a_651_413# VGND 0.0084f
C17234 _324_/a_448_47# VGND 0.0179f
C17235 _324_/a_1108_47# VGND 0.144f
C17236 _324_/a_1283_21# VGND 0.314f
C17237 _324_/a_543_47# VGND 0.172f
C17238 _324_/a_761_289# VGND 0.137f
C17239 _324_/a_193_47# VGND 0.3f
C17240 _324_/a_27_47# VGND 0.512f
C17241 _103_ VGND 0.413f
C17242 _255_/a_27_47# VGND 0.0624f
C17243 _059_ VGND 0.367f
C17244 _186_/a_109_297# VGND -0.00119f
C17245 _341_/a_1462_47# VGND -7.89e-19
C17246 _341_/a_1217_47# VGND -3.93e-19
C17247 _341_/a_805_47# VGND 5.25e-19
C17248 _341_/a_639_47# VGND 0.00113f
C17249 _341_/a_1270_413# VGND 8.12e-20
C17250 _341_/a_651_413# VGND 0.00878f
C17251 _341_/a_448_47# VGND 0.00882f
C17252 _341_/a_1108_47# VGND 0.136f
C17253 _341_/a_1283_21# VGND 0.312f
C17254 _341_/a_543_47# VGND 0.186f
C17255 _341_/a_761_289# VGND 0.136f
C17256 _341_/a_193_47# VGND 0.311f
C17257 _341_/a_27_47# VGND 0.523f
C17258 _114_ VGND 0.122f
C17259 net48 VGND 0.17f
C17260 trim_val\[2\] VGND 0.744f
C17261 _272_/a_384_47# VGND -2.25e-19
C17262 _272_/a_299_297# VGND 0.033f
C17263 _272_/a_81_21# VGND 0.146f
C17264 ctln[7] VGND 0.79f
C17265 net13 VGND 1.11f
C17266 output13/a_27_47# VGND 0.649f
C17267 result[2] VGND 0.226f
C17268 net24 VGND 0.767f
C17269 output24/a_27_47# VGND 0.606f
C17270 trim[4] VGND 0.213f
C17271 output35/a_27_47# VGND 0.616f
C17272 net23 VGND 1.54f
C17273 net43 VGND 5.74f
C17274 _005_ VGND 0.182f
C17275 _308_/a_1462_47# VGND 1.41e-19
C17276 _308_/a_1217_47# VGND -4.83e-19
C17277 _308_/a_805_47# VGND 1.75e-19
C17278 _308_/a_639_47# VGND 3.2e-19
C17279 _308_/a_1270_413# VGND 3.11e-20
C17280 _308_/a_651_413# VGND 0.00526f
C17281 _308_/a_448_47# VGND 0.0148f
C17282 _308_/a_1108_47# VGND 0.132f
C17283 _308_/a_1283_21# VGND 0.313f
C17284 _308_/a_543_47# VGND 0.16f
C17285 _308_/a_761_289# VGND 0.122f
C17286 _308_/a_193_47# VGND 0.277f
C17287 _308_/a_27_47# VGND 0.539f
C17288 _239_/a_474_297# VGND 0.0238f
C17289 _239_/a_277_297# VGND 0.0192f
C17290 _239_/a_27_297# VGND 0.0442f
C17291 _239_/a_694_21# VGND 0.286f
C17292 _325_/a_1462_47# VGND -9.48e-19
C17293 _325_/a_1217_47# VGND -5.03e-19
C17294 _325_/a_805_47# VGND -7.03e-19
C17295 _325_/a_639_47# VGND -0.00151f
C17296 _325_/a_651_413# VGND 0.00788f
C17297 _325_/a_448_47# VGND 0.00886f
C17298 _325_/a_1108_47# VGND 0.132f
C17299 _325_/a_1283_21# VGND 0.316f
C17300 _325_/a_543_47# VGND 0.176f
C17301 _325_/a_761_289# VGND 0.132f
C17302 _325_/a_193_47# VGND 0.297f
C17303 _325_/a_27_47# VGND 0.448f
C17304 _024_ VGND 0.256f
C17305 trim_mask\[0\] VGND 2.82f
C17306 _256_/a_373_47# VGND -6.23e-19
C17307 _256_/a_109_47# VGND -0.00147f
C17308 _256_/a_109_297# VGND 0.00105f
C17309 _256_/a_27_297# VGND 0.197f
C17310 _061_ VGND 0.254f
C17311 _187_/a_297_47# VGND 0.0015f
C17312 _187_/a_212_413# VGND 0.285f
C17313 _187_/a_27_413# VGND 0.248f
C17314 _115_ VGND 0.211f
C17315 _273_/a_145_75# VGND -0.0013f
C17316 _273_/a_59_75# VGND 0.169f
C17317 _127_ VGND 0.254f
C17318 _290_/a_297_47# VGND 2.47e-19
C17319 _290_/a_207_413# VGND 0.132f
C17320 _290_/a_27_413# VGND 0.195f
C17321 ctln[6] VGND 0.603f
C17322 net12 VGND 2.07f
C17323 output12/a_27_47# VGND 0.675f
C17324 result[1] VGND 0.169f
C17325 output23/a_27_47# VGND 0.326f
C17326 trim[3] VGND 0.292f
C17327 output34/a_27_47# VGND 0.602f
C17328 _309_/a_1462_47# VGND -7.68e-19
C17329 _309_/a_1217_47# VGND -5.03e-19
C17330 _309_/a_805_47# VGND 4.87e-19
C17331 _309_/a_639_47# VGND 7.8e-19
C17332 _309_/a_651_413# VGND 0.008f
C17333 _309_/a_448_47# VGND 0.0169f
C17334 _309_/a_1108_47# VGND 0.132f
C17335 _309_/a_1283_21# VGND 0.29f
C17336 _309_/a_543_47# VGND 0.184f
C17337 _309_/a_761_289# VGND 0.139f
C17338 _309_/a_193_47# VGND 0.292f
C17339 _309_/a_27_47# VGND 0.564f
C17340 _326_/a_651_413# VGND 0.00471f
C17341 _326_/a_448_47# VGND 0.0157f
C17342 _326_/a_1108_47# VGND 0.152f
C17343 _326_/a_1283_21# VGND 0.317f
C17344 _326_/a_543_47# VGND 0.16f
C17345 _326_/a_761_289# VGND 0.121f
C17346 _326_/a_193_47# VGND 0.288f
C17347 _326_/a_27_47# VGND 0.498f
C17348 _025_ VGND 0.314f
C17349 _257_/a_373_47# VGND -0.001f
C17350 _257_/a_109_47# VGND -3.65e-19
C17351 _257_/a_109_297# VGND 0.00155f
C17352 _257_/a_27_297# VGND 0.187f
C17353 net5 VGND 0.32f
C17354 _188_/a_27_47# VGND 0.277f
C17355 _274_/a_75_212# VGND 0.249f
C17356 _291_/a_285_47# VGND 0.00334f
C17357 _291_/a_285_297# VGND 0.0295f
C17358 _291_/a_117_297# VGND -3.33e-19
C17359 _291_/a_35_297# VGND 0.291f
C17360 ctln[3] VGND 0.512f
C17361 net9 VGND 1.18f
C17362 output9/a_27_47# VGND 0.311f
C17363 ctln[5] VGND 0.495f
C17364 output11/a_27_47# VGND 0.338f
C17365 result[0] VGND 0.136f
C17366 output22/a_27_47# VGND 0.336f
C17367 trim[2] VGND 0.236f
C17368 output33/a_27_47# VGND 0.58f
C17369 _327_/a_1217_47# VGND 4.72e-20
C17370 _327_/a_805_47# VGND 1.72e-19
C17371 _327_/a_639_47# VGND 3.81e-19
C17372 _327_/a_1270_413# VGND 4.68e-20
C17373 _327_/a_651_413# VGND 0.00866f
C17374 _327_/a_448_47# VGND 0.0155f
C17375 _327_/a_1108_47# VGND 0.156f
C17376 _327_/a_1283_21# VGND 0.428f
C17377 _327_/a_543_47# VGND 0.181f
C17378 _327_/a_761_289# VGND 0.138f
C17379 _327_/a_193_47# VGND 0.297f
C17380 _327_/a_27_47# VGND 0.559f
C17381 trim_mask\[2\] VGND 2.77f
C17382 _258_/a_373_47# VGND -0.0012f
C17383 _258_/a_109_47# VGND -0.0014f
C17384 _258_/a_109_297# VGND 0.00155f
C17385 _258_/a_27_297# VGND 0.193f
C17386 _189_/a_408_47# VGND 0.0397f
C17387 _189_/a_218_47# VGND 0.00955f
C17388 _189_/a_27_47# VGND 0.303f
C17389 net50 VGND 0.439f
C17390 trim_mask\[3\] VGND 1.4f
C17391 trim_val\[3\] VGND 0.623f
C17392 _275_/a_384_47# VGND -2.14e-19
C17393 _275_/a_299_297# VGND 0.0331f
C17394 _275_/a_81_21# VGND 0.176f
C17395 _036_ VGND 0.208f
C17396 cal_count\[1\] VGND 0.508f
C17397 _128_ VGND 0.525f
C17398 _292_/a_215_47# VGND 0.0691f
C17399 _292_/a_493_297# VGND -2.83e-19
C17400 _292_/a_292_297# VGND -0.00118f
C17401 _292_/a_78_199# VGND 0.143f
C17402 ctln[2] VGND 0.626f
C17403 net8 VGND 0.664f
C17404 output8/a_27_47# VGND 0.352f
C17405 ctln[4] VGND 0.52f
C17406 net10 VGND 0.264f
C17407 output10/a_27_47# VGND 0.325f
C17408 ctlp[7] VGND 0.58f
C17409 output21/a_27_47# VGND 0.603f
C17410 trim[1] VGND 0.187f
C17411 output32/a_27_47# VGND 0.604f
C17412 _328_/a_1462_47# VGND -8.64e-19
C17413 _328_/a_1217_47# VGND -4.95e-19
C17414 _328_/a_805_47# VGND 3.45e-19
C17415 _328_/a_639_47# VGND 7.27e-19
C17416 _328_/a_1270_413# VGND 5.15e-20
C17417 _328_/a_651_413# VGND 0.00863f
C17418 _328_/a_448_47# VGND 0.0178f
C17419 _328_/a_1108_47# VGND 0.135f
C17420 _328_/a_1283_21# VGND 0.297f
C17421 _328_/a_543_47# VGND 0.184f
C17422 _328_/a_761_289# VGND 0.139f
C17423 _328_/a_193_47# VGND 0.314f
C17424 _328_/a_27_47# VGND 0.479f
C17425 _104_ VGND 1.6f
C17426 _064_ VGND 1.27f
C17427 _259_/a_373_47# VGND 1.83e-19
C17428 _259_/a_109_47# VGND -7.5e-19
C17429 _259_/a_109_297# VGND 0.00761f
C17430 _259_/a_27_297# VGND 0.202f
C17431 _117_ VGND 0.184f
C17432 _116_ VGND 0.231f
C17433 _110_ VGND 1.69f
C17434 _276_/a_145_75# VGND -2.95e-20
C17435 _276_/a_59_75# VGND 0.198f
C17436 _293_/a_384_47# VGND 0.00107f
C17437 _293_/a_299_297# VGND 0.0499f
C17438 _293_/a_81_21# VGND 0.164f
C17439 ctln[1] VGND 0.506f
C17440 output7/a_27_47# VGND 0.346f
C17441 ctlp[6] VGND 0.587f
C17442 output20/a_27_47# VGND 0.597f
C17443 trim[0] VGND 0.228f
C17444 net31 VGND 1.96f
C17445 output31/a_27_47# VGND 0.562f
C17446 _026_ VGND 0.418f
C17447 _329_/a_1462_47# VGND 3.57e-19
C17448 _329_/a_1217_47# VGND 6.9e-20
C17449 _329_/a_805_47# VGND 6.04e-19
C17450 _329_/a_639_47# VGND 0.00124f
C17451 _329_/a_1270_413# VGND 4.28e-20
C17452 _329_/a_651_413# VGND 0.00862f
C17453 _329_/a_448_47# VGND 0.0192f
C17454 _329_/a_1108_47# VGND 0.145f
C17455 _329_/a_1283_21# VGND 0.317f
C17456 _329_/a_543_47# VGND 0.173f
C17457 _329_/a_761_289# VGND 0.139f
C17458 _329_/a_193_47# VGND 0.317f
C17459 _329_/a_27_47# VGND 0.569f
C17460 _071_ VGND 0.2f
C17461 cal_itt\[1\] VGND 1.12f
C17462 cal_itt\[0\] VGND 1.33f
C17463 cal_itt\[2\] VGND 0.765f
C17464 _200_/a_303_47# VGND -0.00134f
C17465 _200_/a_209_47# VGND -0.00113f
C17466 _200_/a_209_297# VGND 0.00288f
C17467 _200_/a_80_21# VGND 0.189f
C17468 _277_/a_75_212# VGND 0.246f
C17469 VPWR VGND 0.482p
C17470 _294_/a_150_297# VGND -2.09e-19
C17471 _294_/a_68_297# VGND 0.157f
.ends

