magic
tech sky130B
magscale 1 2
timestamp 1694553763
<< viali >>
rect 1501 15657 1535 15691
rect 2789 15657 2823 15691
rect 6561 15657 6595 15691
rect 7941 15657 7975 15691
rect 9137 15657 9171 15691
rect 11713 15657 11747 15691
rect 13185 15657 13219 15691
rect 14381 15657 14415 15691
rect 16221 15657 16255 15691
rect 15853 15589 15887 15623
rect 1961 15453 1995 15487
rect 4629 15453 4663 15487
rect 9321 15453 9355 15487
rect 16129 15453 16163 15487
rect 1777 15385 1811 15419
rect 2329 15385 2363 15419
rect 3065 15385 3099 15419
rect 6469 15385 6503 15419
rect 8217 15385 8251 15419
rect 11621 15385 11655 15419
rect 13093 15385 13127 15419
rect 14657 15385 14691 15419
rect 15577 15385 15611 15419
rect 4813 15317 4847 15351
rect 2421 15113 2455 15147
rect 6101 15113 6135 15147
rect 8125 15113 8159 15147
rect 14841 15113 14875 15147
rect 16405 15113 16439 15147
rect 1409 15045 1443 15079
rect 1777 14977 1811 15011
rect 2145 14977 2179 15011
rect 2237 14977 2271 15011
rect 2329 14977 2363 15011
rect 3157 14977 3191 15011
rect 6193 14977 6227 15011
rect 8217 14977 8251 15011
rect 14933 14977 14967 15011
rect 16129 14977 16163 15011
rect 2973 14841 3007 14875
rect 16129 14297 16163 14331
rect 16497 14297 16531 14331
rect 1593 14025 1627 14059
rect 4905 14025 4939 14059
rect 4077 13957 4111 13991
rect 5733 13957 5767 13991
rect 1409 13889 1443 13923
rect 1869 13889 1903 13923
rect 2881 13889 2915 13923
rect 3249 13889 3283 13923
rect 3801 13889 3835 13923
rect 3893 13889 3927 13923
rect 4353 13889 4387 13923
rect 4813 13889 4847 13923
rect 5089 13889 5123 13923
rect 5365 13889 5399 13923
rect 5549 13889 5583 13923
rect 7021 13889 7055 13923
rect 7205 13889 7239 13923
rect 4445 13821 4479 13855
rect 5273 13821 5307 13855
rect 1685 13685 1719 13719
rect 4721 13685 4755 13719
rect 7113 13685 7147 13719
rect 3157 13481 3191 13515
rect 4629 13481 4663 13515
rect 9597 13481 9631 13515
rect 12909 13481 12943 13515
rect 4537 13413 4571 13447
rect 7757 13413 7791 13447
rect 9229 13413 9263 13447
rect 1409 13345 1443 13379
rect 4169 13345 4203 13379
rect 5273 13345 5307 13379
rect 7665 13345 7699 13379
rect 8033 13345 8067 13379
rect 6745 13277 6779 13311
rect 6929 13277 6963 13311
rect 7205 13277 7239 13311
rect 7297 13277 7331 13311
rect 8125 13277 8159 13311
rect 9781 13277 9815 13311
rect 11161 13277 11195 13311
rect 1685 13209 1719 13243
rect 6561 13209 6595 13243
rect 8953 13209 8987 13243
rect 11437 13209 11471 13243
rect 16129 13209 16163 13243
rect 16497 13209 16531 13243
rect 4721 13141 4755 13175
rect 7021 13141 7055 13175
rect 9413 13141 9447 13175
rect 1961 12937 1995 12971
rect 4445 12937 4479 12971
rect 7297 12937 7331 12971
rect 11989 12937 12023 12971
rect 15301 12937 15335 12971
rect 15945 12937 15979 12971
rect 16129 12937 16163 12971
rect 1777 12869 1811 12903
rect 10609 12869 10643 12903
rect 2145 12801 2179 12835
rect 2513 12801 2547 12835
rect 4629 12801 4663 12835
rect 4721 12801 4755 12835
rect 4997 12801 5031 12835
rect 5365 12801 5399 12835
rect 5457 12801 5491 12835
rect 5733 12801 5767 12835
rect 6377 12801 6411 12835
rect 7205 12801 7239 12835
rect 7389 12801 7423 12835
rect 8585 12801 8619 12835
rect 10885 12801 10919 12835
rect 11713 12801 11747 12835
rect 11897 12801 11931 12835
rect 12173 12801 12207 12835
rect 15117 12801 15151 12835
rect 15761 12801 15795 12835
rect 16037 12801 16071 12835
rect 2329 12733 2363 12767
rect 2881 12733 2915 12767
rect 7021 12733 7055 12767
rect 11529 12733 11563 12767
rect 4307 12665 4341 12699
rect 4905 12665 4939 12699
rect 5641 12665 5675 12699
rect 1501 12597 1535 12631
rect 5181 12597 5215 12631
rect 8493 12597 8527 12631
rect 9137 12597 9171 12631
rect 2329 12393 2363 12427
rect 6975 12393 7009 12427
rect 8585 12393 8619 12427
rect 11897 12393 11931 12427
rect 12541 12325 12575 12359
rect 13461 12325 13495 12359
rect 2513 12257 2547 12291
rect 2605 12257 2639 12291
rect 5549 12257 5583 12291
rect 14105 12257 14139 12291
rect 14381 12257 14415 12291
rect 2053 12189 2087 12223
rect 2697 12189 2731 12223
rect 2789 12189 2823 12223
rect 3341 12189 3375 12223
rect 3985 12189 4019 12223
rect 5181 12189 5215 12223
rect 8769 12189 8803 12223
rect 9873 12189 9907 12223
rect 12081 12189 12115 12223
rect 12173 12189 12207 12223
rect 12265 12189 12299 12223
rect 12357 12189 12391 12223
rect 12909 12189 12943 12223
rect 13277 12189 13311 12223
rect 13553 12189 13587 12223
rect 13737 12189 13771 12223
rect 13829 12189 13863 12223
rect 2973 12121 3007 12155
rect 3157 12121 3191 12155
rect 12725 12121 12759 12155
rect 1869 12053 1903 12087
rect 3801 12053 3835 12087
rect 10425 12053 10459 12087
rect 15853 12053 15887 12087
rect 5043 11849 5077 11883
rect 13921 11849 13955 11883
rect 15117 11849 15151 11883
rect 9965 11781 9999 11815
rect 12909 11781 12943 11815
rect 14749 11781 14783 11815
rect 3249 11713 3283 11747
rect 5825 11713 5859 11747
rect 7205 11713 7239 11747
rect 12357 11713 12391 11747
rect 12817 11713 12851 11747
rect 13093 11713 13127 11747
rect 14197 11713 14231 11747
rect 14933 11713 14967 11747
rect 3617 11645 3651 11679
rect 5917 11645 5951 11679
rect 6193 11645 6227 11679
rect 7113 11645 7147 11679
rect 10241 11645 10275 11679
rect 12081 11645 12115 11679
rect 14105 11645 14139 11679
rect 14289 11645 14323 11679
rect 14381 11645 14415 11679
rect 6837 11577 6871 11611
rect 8493 11509 8527 11543
rect 13277 11509 13311 11543
rect 3433 11305 3467 11339
rect 3893 11305 3927 11339
rect 6561 11305 6595 11339
rect 8585 11305 8619 11339
rect 10701 11305 10735 11339
rect 12725 11305 12759 11339
rect 14105 11305 14139 11339
rect 7481 11237 7515 11271
rect 2421 11169 2455 11203
rect 2605 11169 2639 11203
rect 2697 11169 2731 11203
rect 4353 11169 4387 11203
rect 4537 11169 4571 11203
rect 4813 11169 4847 11203
rect 9321 11169 9355 11203
rect 10977 11169 11011 11203
rect 13369 11169 13403 11203
rect 16405 11169 16439 11203
rect 1869 11101 1903 11135
rect 1961 11101 1995 11135
rect 2145 11101 2179 11135
rect 2237 11101 2271 11135
rect 2789 11101 2823 11135
rect 2881 11101 2915 11135
rect 6745 11101 6779 11135
rect 7297 11101 7331 11135
rect 7389 11101 7423 11135
rect 10241 11101 10275 11135
rect 10333 11101 10367 11135
rect 10517 11101 10551 11135
rect 14749 11101 14783 11135
rect 15761 11101 15795 11135
rect 3065 11033 3099 11067
rect 3249 11033 3283 11067
rect 5089 11033 5123 11067
rect 8401 11033 8435 11067
rect 8601 11033 8635 11067
rect 11253 11033 11287 11067
rect 15853 11033 15887 11067
rect 16129 11033 16163 11067
rect 1685 10965 1719 10999
rect 4261 10965 4295 10999
rect 8769 10965 8803 10999
rect 9965 10965 9999 10999
rect 12817 10965 12851 10999
rect 4537 10761 4571 10795
rect 6929 10761 6963 10795
rect 11805 10761 11839 10795
rect 12173 10761 12207 10795
rect 15117 10761 15151 10795
rect 1685 10693 1719 10727
rect 4997 10693 5031 10727
rect 7297 10693 7331 10727
rect 10404 10693 10438 10727
rect 10609 10693 10643 10727
rect 11161 10693 11195 10727
rect 12357 10693 12391 10727
rect 13369 10693 13403 10727
rect 10931 10659 10965 10693
rect 4353 10625 4387 10659
rect 5365 10625 5399 10659
rect 6745 10625 6779 10659
rect 9873 10625 9907 10659
rect 10057 10625 10091 10659
rect 10149 10625 10183 10659
rect 11989 10625 12023 10659
rect 12262 10647 12296 10681
rect 12587 10659 12621 10693
rect 14933 10625 14967 10659
rect 1409 10557 1443 10591
rect 4721 10557 4755 10591
rect 5181 10557 5215 10591
rect 7021 10557 7055 10591
rect 8769 10557 8803 10591
rect 9413 10557 9447 10591
rect 13093 10557 13127 10591
rect 5273 10489 5307 10523
rect 9689 10489 9723 10523
rect 10241 10489 10275 10523
rect 12725 10489 12759 10523
rect 3157 10421 3191 10455
rect 4721 10421 4755 10455
rect 5181 10421 5215 10455
rect 8861 10421 8895 10455
rect 10425 10421 10459 10455
rect 10793 10421 10827 10455
rect 10977 10421 11011 10455
rect 12541 10421 12575 10455
rect 14841 10421 14875 10455
rect 1501 10217 1535 10251
rect 6745 10217 6779 10251
rect 7021 10217 7055 10251
rect 10057 10217 10091 10251
rect 14933 10217 14967 10251
rect 6929 10081 6963 10115
rect 7573 10081 7607 10115
rect 11161 10081 11195 10115
rect 11529 10081 11563 10115
rect 1777 10013 1811 10047
rect 4629 10013 4663 10047
rect 6653 10013 6687 10047
rect 7389 10013 7423 10047
rect 9505 10013 9539 10047
rect 9689 10013 9723 10047
rect 10701 10013 10735 10047
rect 10977 10013 11011 10047
rect 11253 10013 11287 10047
rect 6929 9945 6963 9979
rect 7481 9945 7515 9979
rect 9873 9945 9907 9979
rect 14565 9945 14599 9979
rect 14749 9945 14783 9979
rect 8953 9877 8987 9911
rect 10793 9877 10827 9911
rect 13001 9877 13035 9911
rect 8953 9605 8987 9639
rect 11989 9605 12023 9639
rect 1777 9537 1811 9571
rect 4169 9537 4203 9571
rect 4537 9537 4571 9571
rect 6377 9537 6411 9571
rect 6560 9537 6594 9571
rect 6745 9537 6779 9571
rect 6929 9537 6963 9571
rect 8677 9537 8711 9571
rect 12633 9537 12667 9571
rect 13185 9537 13219 9571
rect 14105 9537 14139 9571
rect 2053 9469 2087 9503
rect 5963 9469 5997 9503
rect 6653 9469 6687 9503
rect 11069 9469 11103 9503
rect 13001 9469 13035 9503
rect 13461 9469 13495 9503
rect 13645 9469 13679 9503
rect 13737 9469 13771 9503
rect 13829 9469 13863 9503
rect 13921 9469 13955 9503
rect 14381 9469 14415 9503
rect 10517 9401 10551 9435
rect 3525 9333 3559 9367
rect 7021 9333 7055 9367
rect 10425 9333 10459 9367
rect 13369 9333 13403 9367
rect 15853 9333 15887 9367
rect 2237 9129 2271 9163
rect 5273 9129 5307 9163
rect 6653 9129 6687 9163
rect 9321 9129 9355 9163
rect 12541 9129 12575 9163
rect 13001 9129 13035 9163
rect 14289 9129 14323 9163
rect 5457 9061 5491 9095
rect 6193 9061 6227 9095
rect 9229 9061 9263 9095
rect 12817 9061 12851 9095
rect 4353 8993 4387 9027
rect 5733 8993 5767 9027
rect 6561 8993 6595 9027
rect 6745 8993 6779 9027
rect 11529 8993 11563 9027
rect 12173 8993 12207 9027
rect 1777 8925 1811 8959
rect 2421 8925 2455 8959
rect 4997 8925 5031 8959
rect 5181 8925 5215 8959
rect 6009 8925 6043 8959
rect 6653 8925 6687 8959
rect 8953 8925 8987 8959
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 11069 8925 11103 8959
rect 11713 8925 11747 8959
rect 11897 8925 11931 8959
rect 14105 8925 14139 8959
rect 16129 8925 16163 8959
rect 1409 8857 1443 8891
rect 4169 8857 4203 8891
rect 5089 8857 5123 8891
rect 7021 8857 7055 8891
rect 8769 8857 8803 8891
rect 10793 8857 10827 8891
rect 11253 8857 11287 8891
rect 12725 8857 12759 8891
rect 13185 8857 13219 8891
rect 16497 8857 16531 8891
rect 3801 8789 3835 8823
rect 4261 8789 4295 8823
rect 6285 8789 6319 8823
rect 12357 8789 12391 8823
rect 12525 8789 12559 8823
rect 12975 8789 13009 8823
rect 8953 8585 8987 8619
rect 15117 8585 15151 8619
rect 15853 8585 15887 8619
rect 5089 8517 5123 8551
rect 5273 8517 5307 8551
rect 2789 8449 2823 8483
rect 4537 8449 4571 8483
rect 4905 8449 4939 8483
rect 4997 8449 5031 8483
rect 6377 8449 6411 8483
rect 7297 8449 7331 8483
rect 8493 8449 8527 8483
rect 8585 8449 8619 8483
rect 8861 8449 8895 8483
rect 9137 8449 9171 8483
rect 9229 8449 9263 8483
rect 9413 8449 9447 8483
rect 9597 8449 9631 8483
rect 11529 8449 11563 8483
rect 13185 8449 13219 8483
rect 13369 8449 13403 8483
rect 15485 8449 15519 8483
rect 16037 8449 16071 8483
rect 16221 8449 16255 8483
rect 8677 8381 8711 8415
rect 13645 8381 13679 8415
rect 15393 8381 15427 8415
rect 15577 8381 15611 8415
rect 15669 8381 15703 8415
rect 8861 8313 8895 8347
rect 9321 8313 9355 8347
rect 4721 8245 4755 8279
rect 5273 8245 5307 8279
rect 6837 8245 6871 8279
rect 15209 8245 15243 8279
rect 3157 8041 3191 8075
rect 4905 8041 4939 8075
rect 12081 8041 12115 8075
rect 13737 8041 13771 8075
rect 4721 7973 4755 8007
rect 10885 7973 10919 8007
rect 1409 7905 1443 7939
rect 1685 7905 1719 7939
rect 4353 7905 4387 7939
rect 4813 7905 4847 7939
rect 5549 7905 5583 7939
rect 5733 7905 5767 7939
rect 7849 7905 7883 7939
rect 12357 7905 12391 7939
rect 12909 7905 12943 7939
rect 13461 7905 13495 7939
rect 14105 7905 14139 7939
rect 14657 7905 14691 7939
rect 14841 7905 14875 7939
rect 3801 7837 3835 7871
rect 3893 7837 3927 7871
rect 4077 7837 4111 7871
rect 4261 7837 4295 7871
rect 4537 7837 4571 7871
rect 5917 7837 5951 7871
rect 6101 7837 6135 7871
rect 6193 7837 6227 7871
rect 7573 7837 7607 7871
rect 9873 7837 9907 7871
rect 10057 7837 10091 7871
rect 10333 7837 10367 7871
rect 10885 7837 10919 7871
rect 11253 7837 11287 7871
rect 11345 7837 11379 7871
rect 11509 7837 11543 7871
rect 13553 7837 13587 7871
rect 15025 7837 15059 7871
rect 15209 7837 15243 7871
rect 15485 7837 15519 7871
rect 16129 7837 16163 7871
rect 5365 7769 5399 7803
rect 11897 7769 11931 7803
rect 12102 7769 12136 7803
rect 5273 7701 5307 7735
rect 6377 7701 6411 7735
rect 9229 7701 9263 7735
rect 11713 7701 11747 7735
rect 12265 7701 12299 7735
rect 13093 7701 13127 7735
rect 15301 7701 15335 7735
rect 16405 7701 16439 7735
rect 2053 7497 2087 7531
rect 3985 7497 4019 7531
rect 4445 7497 4479 7531
rect 7665 7497 7699 7531
rect 13277 7497 13311 7531
rect 2145 7429 2179 7463
rect 3868 7429 3902 7463
rect 4077 7429 4111 7463
rect 7481 7429 7515 7463
rect 11805 7429 11839 7463
rect 2513 7361 2547 7395
rect 3525 7361 3559 7395
rect 4905 7361 4939 7395
rect 7297 7361 7331 7395
rect 7849 7361 7883 7395
rect 9597 7361 9631 7395
rect 9965 7361 9999 7395
rect 10149 7361 10183 7395
rect 10425 7361 10459 7395
rect 11069 7361 11103 7395
rect 14105 7361 14139 7395
rect 2605 7293 2639 7327
rect 2697 7293 2731 7327
rect 2789 7293 2823 7327
rect 4353 7293 4387 7327
rect 10977 7293 11011 7327
rect 11529 7293 11563 7327
rect 13921 7293 13955 7327
rect 14381 7293 14415 7327
rect 11253 7225 11287 7259
rect 2329 7157 2363 7191
rect 2973 7157 3007 7191
rect 3709 7157 3743 7191
rect 4813 7157 4847 7191
rect 13369 7157 13403 7191
rect 15853 7157 15887 7191
rect 3157 6953 3191 6987
rect 5733 6953 5767 6987
rect 6634 6953 6668 6987
rect 9216 6953 9250 6987
rect 10701 6953 10735 6987
rect 13663 6953 13697 6987
rect 14565 6953 14599 6987
rect 4077 6817 4111 6851
rect 4169 6817 4203 6851
rect 4286 6817 4320 6851
rect 5089 6817 5123 6851
rect 6193 6817 6227 6851
rect 8309 6817 8343 6851
rect 8493 6817 8527 6851
rect 10885 6817 10919 6851
rect 12173 6817 12207 6851
rect 1409 6749 1443 6783
rect 3433 6749 3467 6783
rect 3617 6749 3651 6783
rect 3801 6749 3835 6783
rect 5273 6749 5307 6783
rect 5549 6749 5583 6783
rect 5917 6749 5951 6783
rect 6009 6749 6043 6783
rect 6285 6749 6319 6783
rect 6377 6749 6411 6783
rect 8217 6749 8251 6783
rect 8585 6749 8619 6783
rect 8953 6749 8987 6783
rect 11069 6749 11103 6783
rect 11253 6749 11287 6783
rect 11345 6749 11379 6783
rect 13921 6749 13955 6783
rect 14105 6749 14139 6783
rect 14381 6749 14415 6783
rect 1685 6681 1719 6715
rect 8493 6681 8527 6715
rect 14197 6681 14231 6715
rect 3249 6613 3283 6647
rect 4445 6613 4479 6647
rect 5457 6613 5491 6647
rect 8125 6613 8159 6647
rect 8677 6613 8711 6647
rect 2421 6409 2455 6443
rect 5707 6409 5741 6443
rect 9873 6409 9907 6443
rect 1409 6341 1443 6375
rect 4537 6341 4571 6375
rect 5917 6341 5951 6375
rect 7205 6341 7239 6375
rect 1777 6273 1811 6307
rect 1961 6273 1995 6307
rect 2697 6273 2731 6307
rect 4629 6273 4663 6307
rect 4813 6273 4847 6307
rect 8493 6273 8527 6307
rect 10333 6273 10367 6307
rect 2605 6205 2639 6239
rect 6561 6205 6595 6239
rect 7573 6205 7607 6239
rect 7665 6205 7699 6239
rect 7941 6205 7975 6239
rect 12081 6205 12115 6239
rect 12357 6205 12391 6239
rect 5549 6137 5583 6171
rect 2237 6069 2271 6103
rect 3249 6069 3283 6103
rect 4721 6069 4755 6103
rect 5733 6069 5767 6103
rect 7113 6069 7147 6103
rect 7849 6069 7883 6103
rect 10241 6069 10275 6103
rect 3801 5865 3835 5899
rect 5549 5865 5583 5899
rect 12173 5865 12207 5899
rect 3249 5797 3283 5831
rect 1501 5729 1535 5763
rect 4353 5729 4387 5763
rect 5181 5729 5215 5763
rect 7941 5729 7975 5763
rect 9045 5729 9079 5763
rect 4721 5661 4755 5695
rect 5023 5661 5057 5695
rect 5457 5661 5491 5695
rect 6377 5661 6411 5695
rect 6469 5661 6503 5695
rect 6653 5661 6687 5695
rect 6837 5661 6871 5695
rect 7113 5661 7147 5695
rect 10885 5661 10919 5695
rect 1777 5593 1811 5627
rect 4813 5593 4847 5627
rect 4905 5593 4939 5627
rect 6745 5593 6779 5627
rect 6975 5593 7009 5627
rect 7297 5593 7331 5627
rect 9321 5593 9355 5627
rect 16129 5593 16163 5627
rect 4537 5525 4571 5559
rect 5733 5525 5767 5559
rect 10793 5525 10827 5559
rect 16405 5525 16439 5559
rect 1593 5321 1627 5355
rect 1961 5321 1995 5355
rect 2237 5321 2271 5355
rect 5365 5321 5399 5355
rect 9873 5321 9907 5355
rect 3893 5253 3927 5287
rect 7573 5253 7607 5287
rect 9321 5253 9355 5287
rect 11145 5253 11179 5287
rect 11345 5253 11379 5287
rect 1409 5185 1443 5219
rect 2145 5185 2179 5219
rect 2421 5185 2455 5219
rect 2697 5185 2731 5219
rect 2881 5185 2915 5219
rect 3617 5185 3651 5219
rect 5825 5185 5859 5219
rect 6009 5185 6043 5219
rect 7297 5185 7331 5219
rect 9413 5185 9447 5219
rect 9505 5185 9539 5219
rect 9689 5185 9723 5219
rect 10885 5117 10919 5151
rect 13001 5117 13035 5151
rect 13277 5117 13311 5151
rect 2605 5049 2639 5083
rect 10241 5049 10275 5083
rect 10977 5049 11011 5083
rect 3157 4981 3191 5015
rect 5917 4981 5951 5015
rect 11161 4981 11195 5015
rect 11529 4981 11563 5015
rect 3525 4777 3559 4811
rect 7573 4777 7607 4811
rect 12357 4777 12391 4811
rect 7665 4709 7699 4743
rect 9183 4709 9217 4743
rect 2697 4641 2731 4675
rect 2881 4641 2915 4675
rect 3065 4641 3099 4675
rect 5825 4641 5859 4675
rect 6101 4641 6135 4675
rect 8309 4641 8343 4675
rect 8401 4641 8435 4675
rect 8493 4641 8527 4675
rect 13001 4641 13035 4675
rect 13093 4641 13127 4675
rect 13277 4641 13311 4675
rect 1961 4573 1995 4607
rect 2053 4573 2087 4607
rect 2237 4573 2271 4607
rect 2329 4573 2363 4607
rect 2973 4573 3007 4607
rect 3157 4573 3191 4607
rect 3341 4573 3375 4607
rect 7849 4573 7883 4607
rect 7941 4573 7975 4607
rect 8585 4573 8619 4607
rect 8953 4573 8987 4607
rect 10793 4573 10827 4607
rect 10885 4573 10919 4607
rect 11161 4573 11195 4607
rect 11529 4573 11563 4607
rect 11713 4573 11747 4607
rect 11989 4573 12023 4607
rect 12817 4573 12851 4607
rect 12909 4573 12943 4607
rect 13369 4573 13403 4607
rect 13553 4573 13587 4607
rect 13737 4573 13771 4607
rect 14289 4573 14323 4607
rect 16129 4573 16163 4607
rect 11345 4505 11379 4539
rect 12173 4505 12207 4539
rect 1777 4437 1811 4471
rect 8769 4437 8803 4471
rect 10149 4437 10183 4471
rect 10977 4437 11011 4471
rect 11897 4437 11931 4471
rect 14105 4437 14139 4471
rect 16405 4437 16439 4471
rect 7297 4233 7331 4267
rect 1869 4165 1903 4199
rect 3617 4165 3651 4199
rect 9781 4165 9815 4199
rect 13829 4165 13863 4199
rect 3433 4097 3467 4131
rect 3893 4097 3927 4131
rect 6653 4097 6687 4131
rect 6837 4097 6871 4131
rect 7113 4097 7147 4131
rect 7297 4097 7331 4131
rect 8309 4097 8343 4131
rect 8493 4097 8527 4131
rect 9045 4097 9079 4131
rect 11529 4097 11563 4131
rect 1593 4029 1627 4063
rect 4169 4029 4203 4063
rect 6377 4029 6411 4063
rect 6561 4029 6595 4063
rect 6745 4029 6779 4063
rect 8033 4029 8067 4063
rect 8125 4029 8159 4063
rect 8769 4029 8803 4063
rect 8861 4029 8895 4063
rect 8953 4029 8987 4063
rect 9505 4029 9539 4063
rect 14105 4029 14139 4063
rect 5641 3961 5675 3995
rect 7389 3961 7423 3995
rect 11713 3961 11747 3995
rect 3341 3893 3375 3927
rect 3801 3893 3835 3927
rect 8585 3893 8619 3927
rect 11253 3893 11287 3927
rect 12357 3893 12391 3927
rect 6285 3689 6319 3723
rect 8125 3689 8159 3723
rect 9229 3689 9263 3723
rect 9597 3553 9631 3587
rect 1777 3485 1811 3519
rect 3801 3485 3835 3519
rect 4629 3485 4663 3519
rect 5457 3485 5491 3519
rect 5641 3485 5675 3519
rect 5733 3485 5767 3519
rect 6009 3485 6043 3519
rect 6193 3485 6227 3519
rect 6469 3485 6503 3519
rect 7389 3485 7423 3519
rect 7665 3485 7699 3519
rect 9413 3485 9447 3519
rect 9689 3485 9723 3519
rect 10793 3485 10827 3519
rect 11069 3485 11103 3519
rect 11345 3485 11379 3519
rect 14105 3485 14139 3519
rect 15945 3485 15979 3519
rect 1409 3417 1443 3451
rect 5825 3417 5859 3451
rect 7757 3417 7791 3451
rect 7941 3417 7975 3451
rect 14289 3417 14323 3451
rect 3985 3349 4019 3383
rect 4445 3349 4479 3383
rect 5273 3349 5307 3383
rect 7205 3349 7239 3383
rect 7573 3349 7607 3383
rect 9781 3349 9815 3383
rect 10609 3349 10643 3383
rect 10977 3349 11011 3383
rect 11437 3349 11471 3383
rect 14473 3349 14507 3383
rect 16037 3349 16071 3383
rect 2145 3145 2179 3179
rect 8125 3145 8159 3179
rect 10241 3145 10275 3179
rect 11529 3145 11563 3179
rect 15117 3145 15151 3179
rect 1777 3077 1811 3111
rect 4077 3077 4111 3111
rect 9597 3077 9631 3111
rect 10333 3077 10367 3111
rect 10977 3077 11011 3111
rect 16129 3077 16163 3111
rect 1961 3009 1995 3043
rect 5641 3009 5675 3043
rect 5825 3009 5859 3043
rect 5917 3009 5951 3043
rect 7021 3009 7055 3043
rect 7481 3009 7515 3043
rect 9873 3009 9907 3043
rect 10517 3009 10551 3043
rect 10701 3009 10735 3043
rect 11161 3009 11195 3043
rect 13277 3009 13311 3043
rect 14933 3009 14967 3043
rect 15669 3009 15703 3043
rect 3801 2941 3835 2975
rect 5549 2941 5583 2975
rect 6837 2941 6871 2975
rect 7205 2941 7239 2975
rect 13001 2941 13035 2975
rect 1501 2805 1535 2839
rect 7297 2805 7331 2839
rect 10885 2805 10919 2839
rect 11345 2805 11379 2839
rect 15761 2805 15795 2839
rect 16405 2805 16439 2839
rect 8125 2601 8159 2635
rect 11069 2601 11103 2635
rect 11161 2533 11195 2567
rect 6377 2465 6411 2499
rect 6653 2465 6687 2499
rect 2145 2397 2179 2431
rect 3525 2397 3559 2431
rect 6101 2397 6135 2431
rect 9873 2397 9907 2431
rect 10885 2397 10919 2431
rect 11345 2397 11379 2431
rect 11805 2397 11839 2431
rect 15117 2397 15151 2431
rect 15669 2397 15703 2431
rect 16129 2397 16163 2431
rect 1777 2329 1811 2363
rect 4813 2329 4847 2363
rect 8677 2329 8711 2363
rect 3249 2261 3283 2295
rect 4537 2261 4571 2295
rect 6009 2261 6043 2295
rect 8401 2261 8435 2295
rect 9965 2261 9999 2295
rect 11897 2261 11931 2295
rect 14841 2261 14875 2295
rect 15853 2261 15887 2295
rect 16405 2261 16439 2295
<< metal1 >>
rect 944 15802 16836 15824
rect 944 15750 950 15802
rect 1002 15750 1014 15802
rect 1066 15750 1078 15802
rect 1130 15750 1142 15802
rect 1194 15750 1206 15802
rect 1258 15750 4950 15802
rect 5002 15750 5014 15802
rect 5066 15750 5078 15802
rect 5130 15750 5142 15802
rect 5194 15750 5206 15802
rect 5258 15750 8950 15802
rect 9002 15750 9014 15802
rect 9066 15750 9078 15802
rect 9130 15750 9142 15802
rect 9194 15750 9206 15802
rect 9258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 16836 15802
rect 944 15728 16836 15750
rect 1486 15648 1492 15700
rect 1544 15648 1550 15700
rect 2774 15648 2780 15700
rect 2832 15648 2838 15700
rect 5810 15648 5816 15700
rect 5868 15688 5874 15700
rect 6549 15691 6607 15697
rect 6549 15688 6561 15691
rect 5868 15660 6561 15688
rect 5868 15648 5874 15660
rect 6549 15657 6561 15660
rect 6595 15657 6607 15691
rect 6549 15651 6607 15657
rect 7834 15648 7840 15700
rect 7892 15688 7898 15700
rect 7929 15691 7987 15697
rect 7929 15688 7941 15691
rect 7892 15660 7941 15688
rect 7892 15648 7898 15660
rect 7929 15657 7941 15660
rect 7975 15657 7987 15691
rect 7929 15651 7987 15657
rect 9125 15691 9183 15697
rect 9125 15657 9137 15691
rect 9171 15688 9183 15691
rect 9306 15688 9312 15700
rect 9171 15660 9312 15688
rect 9171 15657 9183 15660
rect 9125 15651 9183 15657
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 11701 15691 11759 15697
rect 11701 15688 11713 15691
rect 11112 15660 11713 15688
rect 11112 15648 11118 15660
rect 11701 15657 11713 15660
rect 11747 15657 11759 15691
rect 11701 15651 11759 15657
rect 12802 15648 12808 15700
rect 12860 15688 12866 15700
rect 13173 15691 13231 15697
rect 13173 15688 13185 15691
rect 12860 15660 13185 15688
rect 12860 15648 12866 15660
rect 13173 15657 13185 15660
rect 13219 15657 13231 15691
rect 13173 15651 13231 15657
rect 14366 15648 14372 15700
rect 14424 15648 14430 15700
rect 16206 15648 16212 15700
rect 16264 15648 16270 15700
rect 15841 15623 15899 15629
rect 15841 15589 15853 15623
rect 15887 15620 15899 15623
rect 17402 15620 17408 15632
rect 15887 15592 17408 15620
rect 15887 15589 15899 15592
rect 15841 15583 15899 15589
rect 17402 15580 17408 15592
rect 17460 15580 17466 15632
rect 658 15444 664 15496
rect 716 15484 722 15496
rect 1949 15487 2007 15493
rect 1949 15484 1961 15487
rect 716 15456 1961 15484
rect 716 15444 722 15456
rect 1949 15453 1961 15456
rect 1995 15453 2007 15487
rect 1949 15447 2007 15453
rect 4522 15444 4528 15496
rect 4580 15484 4586 15496
rect 4617 15487 4675 15493
rect 4617 15484 4629 15487
rect 4580 15456 4629 15484
rect 4580 15444 4586 15456
rect 4617 15453 4629 15456
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 9306 15444 9312 15496
rect 9364 15444 9370 15496
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 15304 15456 16129 15484
rect 15304 15428 15332 15456
rect 16117 15453 16129 15456
rect 16163 15453 16175 15487
rect 16117 15447 16175 15453
rect 1765 15419 1823 15425
rect 1765 15385 1777 15419
rect 1811 15385 1823 15419
rect 1765 15379 1823 15385
rect 1780 15348 1808 15379
rect 2314 15376 2320 15428
rect 2372 15376 2378 15428
rect 3050 15376 3056 15428
rect 3108 15376 3114 15428
rect 6270 15416 6276 15428
rect 4724 15388 6276 15416
rect 4724 15348 4752 15388
rect 6270 15376 6276 15388
rect 6328 15376 6334 15428
rect 6454 15376 6460 15428
rect 6512 15376 6518 15428
rect 8202 15376 8208 15428
rect 8260 15376 8266 15428
rect 11606 15376 11612 15428
rect 11664 15376 11670 15428
rect 12802 15376 12808 15428
rect 12860 15416 12866 15428
rect 13081 15419 13139 15425
rect 13081 15416 13093 15419
rect 12860 15388 13093 15416
rect 12860 15376 12866 15388
rect 13081 15385 13093 15388
rect 13127 15385 13139 15419
rect 13081 15379 13139 15385
rect 14642 15376 14648 15428
rect 14700 15376 14706 15428
rect 15286 15376 15292 15428
rect 15344 15376 15350 15428
rect 15562 15376 15568 15428
rect 15620 15376 15626 15428
rect 1780 15320 4752 15348
rect 4801 15351 4859 15357
rect 4801 15317 4813 15351
rect 4847 15348 4859 15351
rect 5994 15348 6000 15360
rect 4847 15320 6000 15348
rect 4847 15317 4859 15320
rect 4801 15311 4859 15317
rect 5994 15308 6000 15320
rect 6052 15308 6058 15360
rect 1104 15258 16836 15280
rect 1104 15206 1610 15258
rect 1662 15206 1674 15258
rect 1726 15206 1738 15258
rect 1790 15206 1802 15258
rect 1854 15206 1866 15258
rect 1918 15206 5610 15258
rect 5662 15206 5674 15258
rect 5726 15206 5738 15258
rect 5790 15206 5802 15258
rect 5854 15206 5866 15258
rect 5918 15206 9610 15258
rect 9662 15206 9674 15258
rect 9726 15206 9738 15258
rect 9790 15206 9802 15258
rect 9854 15206 9866 15258
rect 9918 15206 13610 15258
rect 13662 15206 13674 15258
rect 13726 15206 13738 15258
rect 13790 15206 13802 15258
rect 13854 15206 13866 15258
rect 13918 15206 16836 15258
rect 1104 15184 16836 15206
rect 2314 15104 2320 15156
rect 2372 15144 2378 15156
rect 2409 15147 2467 15153
rect 2409 15144 2421 15147
rect 2372 15116 2421 15144
rect 2372 15104 2378 15116
rect 2409 15113 2421 15116
rect 2455 15113 2467 15147
rect 2409 15107 2467 15113
rect 6089 15147 6147 15153
rect 6089 15113 6101 15147
rect 6135 15144 6147 15147
rect 6454 15144 6460 15156
rect 6135 15116 6460 15144
rect 6135 15113 6147 15116
rect 6089 15107 6147 15113
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 8113 15147 8171 15153
rect 8113 15113 8125 15147
rect 8159 15144 8171 15147
rect 8202 15144 8208 15156
rect 8159 15116 8208 15144
rect 8159 15113 8171 15116
rect 8113 15107 8171 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 14642 15104 14648 15156
rect 14700 15144 14706 15156
rect 14829 15147 14887 15153
rect 14829 15144 14841 15147
rect 14700 15116 14841 15144
rect 14700 15104 14706 15116
rect 14829 15113 14841 15116
rect 14875 15113 14887 15147
rect 14829 15107 14887 15113
rect 16393 15147 16451 15153
rect 16393 15113 16405 15147
rect 16439 15144 16451 15147
rect 16482 15144 16488 15156
rect 16439 15116 16488 15144
rect 16439 15113 16451 15116
rect 16393 15107 16451 15113
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 1394 15036 1400 15088
rect 1452 15036 1458 15088
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 2133 15011 2191 15017
rect 2133 15008 2145 15011
rect 1811 14980 2145 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 2133 14977 2145 14980
rect 2179 14977 2191 15011
rect 2133 14971 2191 14977
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2240 14940 2268 14971
rect 2314 14968 2320 15020
rect 2372 14968 2378 15020
rect 3142 14968 3148 15020
rect 3200 14968 3206 15020
rect 6178 14968 6184 15020
rect 6236 14968 6242 15020
rect 8202 14968 8208 15020
rect 8260 14968 8266 15020
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 15008 14979 15011
rect 15286 15008 15292 15020
rect 14967 14980 15292 15008
rect 14967 14977 14979 14980
rect 14921 14971 14979 14977
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 16114 14968 16120 15020
rect 16172 14968 16178 15020
rect 11606 14940 11612 14952
rect 2240 14912 11612 14940
rect 2976 14881 3004 14912
rect 11606 14900 11612 14912
rect 11664 14900 11670 14952
rect 2961 14875 3019 14881
rect 2961 14841 2973 14875
rect 3007 14872 3019 14875
rect 3007 14844 3041 14872
rect 3007 14841 3019 14844
rect 2961 14835 3019 14841
rect 944 14714 16836 14736
rect 944 14662 950 14714
rect 1002 14662 1014 14714
rect 1066 14662 1078 14714
rect 1130 14662 1142 14714
rect 1194 14662 1206 14714
rect 1258 14662 4950 14714
rect 5002 14662 5014 14714
rect 5066 14662 5078 14714
rect 5130 14662 5142 14714
rect 5194 14662 5206 14714
rect 5258 14662 8950 14714
rect 9002 14662 9014 14714
rect 9066 14662 9078 14714
rect 9130 14662 9142 14714
rect 9194 14662 9206 14714
rect 9258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 16836 14714
rect 944 14640 16836 14662
rect 5074 14328 5080 14340
rect 2884 14300 5080 14328
rect 2884 14272 2912 14300
rect 5074 14288 5080 14300
rect 5132 14288 5138 14340
rect 15930 14288 15936 14340
rect 15988 14328 15994 14340
rect 16117 14331 16175 14337
rect 16117 14328 16129 14331
rect 15988 14300 16129 14328
rect 15988 14288 15994 14300
rect 16117 14297 16129 14300
rect 16163 14297 16175 14331
rect 16117 14291 16175 14297
rect 16485 14331 16543 14337
rect 16485 14297 16497 14331
rect 16531 14328 16543 14331
rect 16942 14328 16948 14340
rect 16531 14300 16948 14328
rect 16531 14297 16543 14300
rect 16485 14291 16543 14297
rect 16942 14288 16948 14300
rect 17000 14288 17006 14340
rect 2866 14220 2872 14272
rect 2924 14220 2930 14272
rect 3786 14220 3792 14272
rect 3844 14260 3850 14272
rect 5534 14260 5540 14272
rect 3844 14232 5540 14260
rect 3844 14220 3850 14232
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 1104 14170 16836 14192
rect 1104 14118 1610 14170
rect 1662 14118 1674 14170
rect 1726 14118 1738 14170
rect 1790 14118 1802 14170
rect 1854 14118 1866 14170
rect 1918 14118 5610 14170
rect 5662 14118 5674 14170
rect 5726 14118 5738 14170
rect 5790 14118 5802 14170
rect 5854 14118 5866 14170
rect 5918 14118 9610 14170
rect 9662 14118 9674 14170
rect 9726 14118 9738 14170
rect 9790 14118 9802 14170
rect 9854 14118 9866 14170
rect 9918 14118 13610 14170
rect 13662 14118 13674 14170
rect 13726 14118 13738 14170
rect 13790 14118 13802 14170
rect 13854 14118 13866 14170
rect 13918 14118 16836 14170
rect 1104 14096 16836 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1627 14028 3280 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 1946 13920 1952 13932
rect 1903 13892 1952 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 2866 13880 2872 13932
rect 2924 13880 2930 13932
rect 3252 13929 3280 14028
rect 3786 14016 3792 14068
rect 3844 14016 3850 14068
rect 4522 14016 4528 14068
rect 4580 14056 4586 14068
rect 4893 14059 4951 14065
rect 4893 14056 4905 14059
rect 4580 14028 4905 14056
rect 4580 14016 4586 14028
rect 4893 14025 4905 14028
rect 4939 14025 4951 14059
rect 4893 14019 4951 14025
rect 5074 14016 5080 14068
rect 5132 14056 5138 14068
rect 5132 14028 7236 14056
rect 5132 14016 5138 14028
rect 3804 13929 3832 14016
rect 4065 13991 4123 13997
rect 4065 13957 4077 13991
rect 4111 13988 4123 13991
rect 4154 13988 4160 14000
rect 4111 13960 4160 13988
rect 4111 13957 4123 13960
rect 4065 13951 4123 13957
rect 4154 13948 4160 13960
rect 4212 13988 4218 14000
rect 5721 13991 5779 13997
rect 5721 13988 5733 13991
rect 4212 13960 5120 13988
rect 4212 13948 4218 13960
rect 3237 13923 3295 13929
rect 3237 13889 3249 13923
rect 3283 13920 3295 13923
rect 3789 13923 3847 13929
rect 3789 13920 3801 13923
rect 3283 13892 3801 13920
rect 3283 13889 3295 13892
rect 3237 13883 3295 13889
rect 3789 13889 3801 13892
rect 3835 13889 3847 13923
rect 3789 13883 3847 13889
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13889 3939 13923
rect 3881 13883 3939 13889
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4522 13920 4528 13932
rect 4387 13892 4528 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 3896 13852 3924 13883
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4798 13880 4804 13932
rect 4856 13920 4862 13932
rect 5092 13929 5120 13960
rect 5184 13960 5733 13988
rect 5077 13923 5135 13929
rect 4856 13892 5028 13920
rect 4856 13880 4862 13892
rect 4246 13852 4252 13864
rect 3896 13824 4252 13852
rect 4246 13812 4252 13824
rect 4304 13852 4310 13864
rect 4433 13855 4491 13861
rect 4304 13824 4384 13852
rect 4304 13812 4310 13824
rect 4356 13784 4384 13824
rect 4433 13821 4445 13855
rect 4479 13852 4491 13855
rect 4614 13852 4620 13864
rect 4479 13824 4620 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 5000 13852 5028 13892
rect 5077 13889 5089 13923
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5184 13852 5212 13960
rect 5721 13957 5733 13960
rect 5767 13957 5779 13991
rect 5721 13951 5779 13957
rect 5350 13880 5356 13932
rect 5408 13880 5414 13932
rect 5534 13880 5540 13932
rect 5592 13920 5598 13932
rect 6730 13920 6736 13932
rect 5592 13892 6736 13920
rect 5592 13880 5598 13892
rect 6730 13880 6736 13892
rect 6788 13880 6794 13932
rect 6914 13880 6920 13932
rect 6972 13920 6978 13932
rect 7208 13929 7236 14028
rect 7009 13923 7067 13929
rect 7009 13920 7021 13923
rect 6972 13892 7021 13920
rect 6972 13880 6978 13892
rect 7009 13889 7021 13892
rect 7055 13889 7067 13923
rect 7009 13883 7067 13889
rect 7193 13923 7251 13929
rect 7193 13889 7205 13923
rect 7239 13920 7251 13923
rect 7466 13920 7472 13932
rect 7239 13892 7472 13920
rect 7239 13889 7251 13892
rect 7193 13883 7251 13889
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 5000 13824 5212 13852
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 6822 13852 6828 13864
rect 5307 13824 6828 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 5350 13784 5356 13796
rect 4356 13756 5356 13784
rect 5350 13744 5356 13756
rect 5408 13744 5414 13796
rect 1670 13676 1676 13728
rect 1728 13676 1734 13728
rect 4706 13676 4712 13728
rect 4764 13676 4770 13728
rect 7098 13676 7104 13728
rect 7156 13676 7162 13728
rect 944 13626 16836 13648
rect 944 13574 950 13626
rect 1002 13574 1014 13626
rect 1066 13574 1078 13626
rect 1130 13574 1142 13626
rect 1194 13574 1206 13626
rect 1258 13574 4950 13626
rect 5002 13574 5014 13626
rect 5066 13574 5078 13626
rect 5130 13574 5142 13626
rect 5194 13574 5206 13626
rect 5258 13574 8950 13626
rect 9002 13574 9014 13626
rect 9066 13574 9078 13626
rect 9130 13574 9142 13626
rect 9194 13574 9206 13626
rect 9258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 16836 13626
rect 944 13552 16836 13574
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 3145 13515 3203 13521
rect 3145 13512 3157 13515
rect 3108 13484 3157 13512
rect 3108 13472 3114 13484
rect 3145 13481 3157 13484
rect 3191 13512 3203 13515
rect 3326 13512 3332 13524
rect 3191 13484 3332 13512
rect 3191 13481 3203 13484
rect 3145 13475 3203 13481
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 4614 13472 4620 13524
rect 4672 13472 4678 13524
rect 4908 13484 8248 13512
rect 4525 13447 4583 13453
rect 4525 13413 4537 13447
rect 4571 13444 4583 13447
rect 4798 13444 4804 13456
rect 4571 13416 4804 13444
rect 4571 13413 4583 13416
rect 4525 13407 4583 13413
rect 4798 13404 4804 13416
rect 4856 13404 4862 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2958 13376 2964 13388
rect 1443 13348 2964 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2958 13336 2964 13348
rect 3016 13336 3022 13388
rect 4154 13336 4160 13388
rect 4212 13336 4218 13388
rect 1670 13200 1676 13252
rect 1728 13200 1734 13252
rect 4062 13240 4068 13252
rect 2898 13212 4068 13240
rect 4062 13200 4068 13212
rect 4120 13200 4126 13252
rect 4908 13240 4936 13484
rect 5350 13404 5356 13456
rect 5408 13404 5414 13456
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 7745 13447 7803 13453
rect 7745 13444 7757 13447
rect 5592 13416 7757 13444
rect 5592 13404 5598 13416
rect 7745 13413 7757 13416
rect 7791 13413 7803 13447
rect 7745 13407 7803 13413
rect 7944 13416 8156 13444
rect 5261 13379 5319 13385
rect 5261 13345 5273 13379
rect 5307 13376 5319 13379
rect 5368 13376 5396 13404
rect 5307 13348 5396 13376
rect 5307 13345 5319 13348
rect 5261 13339 5319 13345
rect 6822 13336 6828 13388
rect 6880 13336 6886 13388
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7374 13376 7380 13388
rect 7156 13348 7380 13376
rect 7156 13336 7162 13348
rect 7374 13336 7380 13348
rect 7432 13376 7438 13388
rect 7653 13379 7711 13385
rect 7653 13376 7665 13379
rect 7432 13348 7665 13376
rect 7432 13336 7438 13348
rect 7653 13345 7665 13348
rect 7699 13345 7711 13379
rect 7653 13339 7711 13345
rect 6730 13268 6736 13320
rect 6788 13268 6794 13320
rect 4632 13212 4936 13240
rect 6549 13243 6607 13249
rect 2590 13132 2596 13184
rect 2648 13172 2654 13184
rect 4632 13172 4660 13212
rect 6549 13209 6561 13243
rect 6595 13209 6607 13243
rect 6840 13240 6868 13336
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13308 6975 13311
rect 7190 13308 7196 13320
rect 6963 13280 7196 13308
rect 6963 13277 6975 13280
rect 6917 13271 6975 13277
rect 7190 13268 7196 13280
rect 7248 13268 7254 13320
rect 7285 13311 7343 13317
rect 7285 13277 7297 13311
rect 7331 13308 7343 13311
rect 7944 13308 7972 13416
rect 8021 13379 8079 13385
rect 8021 13345 8033 13379
rect 8067 13345 8079 13379
rect 8021 13339 8079 13345
rect 7331 13280 7972 13308
rect 7331 13277 7343 13280
rect 7285 13271 7343 13277
rect 7300 13240 7328 13271
rect 8036 13240 8064 13339
rect 8128 13317 8156 13416
rect 8220 13376 8248 13484
rect 9306 13472 9312 13524
rect 9364 13512 9370 13524
rect 9585 13515 9643 13521
rect 9585 13512 9597 13515
rect 9364 13484 9597 13512
rect 9364 13472 9370 13484
rect 9585 13481 9597 13484
rect 9631 13481 9643 13515
rect 9585 13475 9643 13481
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 12897 13515 12955 13521
rect 12897 13512 12909 13515
rect 12860 13484 12909 13512
rect 12860 13472 12866 13484
rect 12897 13481 12909 13484
rect 12943 13481 12955 13515
rect 12897 13475 12955 13481
rect 9217 13447 9275 13453
rect 9217 13413 9229 13447
rect 9263 13444 9275 13447
rect 10226 13444 10232 13456
rect 9263 13416 10232 13444
rect 9263 13413 9275 13416
rect 9217 13407 9275 13413
rect 10226 13404 10232 13416
rect 10284 13404 10290 13456
rect 8220 13348 9904 13376
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 6840 13212 7328 13240
rect 7392 13212 8064 13240
rect 6549 13203 6607 13209
rect 2648 13144 4660 13172
rect 4709 13175 4767 13181
rect 2648 13132 2654 13144
rect 4709 13141 4721 13175
rect 4755 13172 4767 13175
rect 4890 13172 4896 13184
rect 4755 13144 4896 13172
rect 4755 13141 4767 13144
rect 4709 13135 4767 13141
rect 4890 13132 4896 13144
rect 4948 13132 4954 13184
rect 6564 13172 6592 13203
rect 6914 13172 6920 13184
rect 6564 13144 6920 13172
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 7006 13132 7012 13184
rect 7064 13132 7070 13184
rect 7282 13132 7288 13184
rect 7340 13172 7346 13184
rect 7392 13172 7420 13212
rect 8662 13200 8668 13252
rect 8720 13240 8726 13252
rect 8941 13243 8999 13249
rect 8941 13240 8953 13243
rect 8720 13212 8953 13240
rect 8720 13200 8726 13212
rect 8941 13209 8953 13212
rect 8987 13209 8999 13243
rect 8941 13203 8999 13209
rect 7340 13144 7420 13172
rect 9401 13175 9459 13181
rect 7340 13132 7346 13144
rect 9401 13141 9413 13175
rect 9447 13172 9459 13175
rect 9784 13172 9812 13271
rect 9447 13144 9812 13172
rect 9876 13172 9904 13348
rect 10870 13268 10876 13320
rect 10928 13308 10934 13320
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 10928 13280 11161 13308
rect 10928 13268 10934 13280
rect 11149 13277 11161 13280
rect 11195 13277 11207 13311
rect 11149 13271 11207 13277
rect 11422 13200 11428 13252
rect 11480 13200 11486 13252
rect 12710 13240 12716 13252
rect 12650 13212 12716 13240
rect 12710 13200 12716 13212
rect 12768 13200 12774 13252
rect 16114 13200 16120 13252
rect 16172 13200 16178 13252
rect 16485 13243 16543 13249
rect 16485 13209 16497 13243
rect 16531 13209 16543 13243
rect 16485 13203 16543 13209
rect 13998 13172 14004 13184
rect 9876 13144 14004 13172
rect 9447 13141 9459 13144
rect 9401 13135 9459 13141
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 16500 13172 16528 13203
rect 16942 13172 16948 13184
rect 16500 13144 16948 13172
rect 16942 13132 16948 13144
rect 17000 13132 17006 13184
rect 1104 13082 16836 13104
rect 1104 13030 1610 13082
rect 1662 13030 1674 13082
rect 1726 13030 1738 13082
rect 1790 13030 1802 13082
rect 1854 13030 1866 13082
rect 1918 13030 5610 13082
rect 5662 13030 5674 13082
rect 5726 13030 5738 13082
rect 5790 13030 5802 13082
rect 5854 13030 5866 13082
rect 5918 13030 9610 13082
rect 9662 13030 9674 13082
rect 9726 13030 9738 13082
rect 9790 13030 9802 13082
rect 9854 13030 9866 13082
rect 9918 13030 13610 13082
rect 13662 13030 13674 13082
rect 13726 13030 13738 13082
rect 13790 13030 13802 13082
rect 13854 13030 13866 13082
rect 13918 13030 16836 13082
rect 1104 13008 16836 13030
rect 1946 12928 1952 12980
rect 2004 12928 2010 12980
rect 2590 12928 2596 12980
rect 2648 12928 2654 12980
rect 2866 12928 2872 12980
rect 2924 12968 2930 12980
rect 4433 12971 4491 12977
rect 4433 12968 4445 12971
rect 2924 12940 4445 12968
rect 2924 12928 2930 12940
rect 4433 12937 4445 12940
rect 4479 12937 4491 12971
rect 4433 12931 4491 12937
rect 4890 12928 4896 12980
rect 4948 12968 4954 12980
rect 4948 12940 5028 12968
rect 4948 12928 4954 12940
rect 1765 12903 1823 12909
rect 1765 12869 1777 12903
rect 1811 12900 1823 12903
rect 2608 12900 2636 12928
rect 4062 12900 4068 12912
rect 1811 12872 2636 12900
rect 3910 12872 4068 12900
rect 1811 12869 1823 12872
rect 1765 12863 1823 12869
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 2130 12792 2136 12844
rect 2188 12792 2194 12844
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 2958 12832 2964 12844
rect 2547 12804 2964 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 4338 12792 4344 12844
rect 4396 12832 4402 12844
rect 4617 12835 4675 12841
rect 4617 12832 4629 12835
rect 4396 12804 4629 12832
rect 4396 12792 4402 12804
rect 4617 12801 4629 12804
rect 4663 12801 4675 12835
rect 4617 12795 4675 12801
rect 2317 12767 2375 12773
rect 2317 12733 2329 12767
rect 2363 12764 2375 12767
rect 2363 12736 2544 12764
rect 2363 12733 2375 12736
rect 2317 12727 2375 12733
rect 2516 12640 2544 12736
rect 2866 12724 2872 12776
rect 2924 12724 2930 12776
rect 2976 12764 3004 12792
rect 3234 12764 3240 12776
rect 2976 12736 3240 12764
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 4632 12764 4660 12795
rect 4706 12792 4712 12844
rect 4764 12792 4770 12844
rect 5000 12841 5028 12940
rect 7190 12928 7196 12980
rect 7248 12928 7254 12980
rect 7282 12928 7288 12980
rect 7340 12928 7346 12980
rect 7374 12928 7380 12980
rect 7432 12928 7438 12980
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 8720 12940 10916 12968
rect 8720 12928 8726 12940
rect 5092 12872 6868 12900
rect 5092 12844 5120 12872
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12801 5043 12835
rect 4985 12795 5043 12801
rect 5074 12792 5080 12844
rect 5132 12792 5138 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 5534 12832 5540 12844
rect 5491 12804 5540 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 5368 12764 5396 12795
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 5721 12835 5779 12841
rect 5721 12801 5733 12835
rect 5767 12832 5779 12835
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 5767 12804 6377 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 6365 12801 6377 12804
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 4632 12736 5396 12764
rect 4246 12656 4252 12708
rect 4304 12705 4310 12708
rect 4304 12699 4353 12705
rect 4304 12665 4307 12699
rect 4341 12665 4353 12699
rect 4304 12659 4353 12665
rect 4893 12699 4951 12705
rect 4893 12665 4905 12699
rect 4939 12696 4951 12699
rect 5350 12696 5356 12708
rect 4939 12668 5356 12696
rect 4939 12665 4951 12668
rect 4893 12659 4951 12665
rect 4304 12656 4310 12659
rect 5350 12656 5356 12668
rect 5408 12696 5414 12708
rect 5629 12699 5687 12705
rect 5629 12696 5641 12699
rect 5408 12668 5641 12696
rect 5408 12656 5414 12668
rect 5629 12665 5641 12668
rect 5675 12665 5687 12699
rect 6840 12696 6868 12872
rect 7208 12841 7236 12928
rect 7392 12841 7420 12928
rect 10594 12860 10600 12912
rect 10652 12860 10658 12912
rect 10888 12844 10916 12940
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11480 12940 11989 12968
rect 11480 12928 11486 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 11977 12931 12035 12937
rect 15286 12928 15292 12980
rect 15344 12928 15350 12980
rect 15562 12928 15568 12980
rect 15620 12928 15626 12980
rect 15930 12928 15936 12980
rect 15988 12928 15994 12980
rect 16114 12928 16120 12980
rect 16172 12928 16178 12980
rect 15580 12900 15608 12928
rect 12406 12872 15608 12900
rect 7193 12835 7251 12841
rect 7193 12801 7205 12835
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 9306 12832 9312 12844
rect 8628 12804 9312 12832
rect 8628 12792 8634 12804
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9490 12792 9496 12844
rect 9548 12792 9554 12844
rect 10870 12792 10876 12844
rect 10928 12792 10934 12844
rect 11698 12792 11704 12844
rect 11756 12792 11762 12844
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12832 11943 12835
rect 12161 12835 12219 12841
rect 12161 12832 12173 12835
rect 11931 12804 12173 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 12161 12801 12173 12804
rect 12207 12801 12219 12835
rect 12161 12795 12219 12801
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7009 12767 7067 12773
rect 7009 12764 7021 12767
rect 6972 12736 7021 12764
rect 6972 12724 6978 12736
rect 7009 12733 7021 12736
rect 7055 12764 7067 12767
rect 7282 12764 7288 12776
rect 7055 12736 7288 12764
rect 7055 12733 7067 12736
rect 7009 12727 7067 12733
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 9600 12736 11529 12764
rect 9600 12696 9628 12736
rect 11517 12733 11529 12736
rect 11563 12764 11575 12767
rect 11790 12764 11796 12776
rect 11563 12736 11796 12764
rect 11563 12733 11575 12736
rect 11517 12727 11575 12733
rect 11790 12724 11796 12736
rect 11848 12724 11854 12776
rect 12406 12696 12434 12872
rect 15102 12792 15108 12844
rect 15160 12792 15166 12844
rect 15746 12792 15752 12844
rect 15804 12792 15810 12844
rect 15948 12832 15976 12928
rect 16025 12835 16083 12841
rect 16025 12832 16037 12835
rect 15948 12804 16037 12832
rect 16025 12801 16037 12804
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 6840 12668 9628 12696
rect 10796 12668 12434 12696
rect 5629 12659 5687 12665
rect 1486 12588 1492 12640
rect 1544 12588 1550 12640
rect 2498 12588 2504 12640
rect 2556 12628 2562 12640
rect 5074 12628 5080 12640
rect 2556 12600 5080 12628
rect 2556 12588 2562 12600
rect 5074 12588 5080 12600
rect 5132 12588 5138 12640
rect 5169 12631 5227 12637
rect 5169 12597 5181 12631
rect 5215 12628 5227 12631
rect 5534 12628 5540 12640
rect 5215 12600 5540 12628
rect 5215 12597 5227 12600
rect 5169 12591 5227 12597
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 6270 12588 6276 12640
rect 6328 12628 6334 12640
rect 8481 12631 8539 12637
rect 8481 12628 8493 12631
rect 6328 12600 8493 12628
rect 6328 12588 6334 12600
rect 8481 12597 8493 12600
rect 8527 12597 8539 12631
rect 8481 12591 8539 12597
rect 9122 12588 9128 12640
rect 9180 12588 9186 12640
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 10796 12628 10824 12668
rect 9456 12600 10824 12628
rect 9456 12588 9462 12600
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 13814 12628 13820 12640
rect 11848 12600 13820 12628
rect 11848 12588 11854 12600
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 944 12538 16836 12560
rect 944 12486 950 12538
rect 1002 12486 1014 12538
rect 1066 12486 1078 12538
rect 1130 12486 1142 12538
rect 1194 12486 1206 12538
rect 1258 12486 4950 12538
rect 5002 12486 5014 12538
rect 5066 12486 5078 12538
rect 5130 12486 5142 12538
rect 5194 12486 5206 12538
rect 5258 12486 8950 12538
rect 9002 12486 9014 12538
rect 9066 12486 9078 12538
rect 9130 12486 9142 12538
rect 9194 12486 9206 12538
rect 9258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 16836 12538
rect 944 12464 16836 12486
rect 2130 12384 2136 12436
rect 2188 12424 2194 12436
rect 2317 12427 2375 12433
rect 2317 12424 2329 12427
rect 2188 12396 2329 12424
rect 2188 12384 2194 12396
rect 2317 12393 2329 12396
rect 2363 12393 2375 12427
rect 2317 12387 2375 12393
rect 6963 12427 7021 12433
rect 6963 12393 6975 12427
rect 7009 12424 7021 12427
rect 7282 12424 7288 12436
rect 7009 12396 7288 12424
rect 7009 12393 7021 12396
rect 6963 12387 7021 12393
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 8570 12384 8576 12436
rect 8628 12384 8634 12436
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 11885 12427 11943 12433
rect 11885 12424 11897 12427
rect 11756 12396 11897 12424
rect 11756 12384 11762 12396
rect 11885 12393 11897 12396
rect 11931 12393 11943 12427
rect 14182 12424 14188 12436
rect 11885 12387 11943 12393
rect 12406 12396 14188 12424
rect 2866 12356 2872 12368
rect 2516 12328 2872 12356
rect 2516 12297 2544 12328
rect 2866 12316 2872 12328
rect 2924 12316 2930 12368
rect 7466 12316 7472 12368
rect 7524 12356 7530 12368
rect 12250 12356 12256 12368
rect 7524 12328 12256 12356
rect 7524 12316 7530 12328
rect 12250 12316 12256 12328
rect 12308 12356 12314 12368
rect 12406 12356 12434 12396
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 12308 12328 12434 12356
rect 12308 12316 12314 12328
rect 12526 12316 12532 12368
rect 12584 12316 12590 12368
rect 13449 12359 13507 12365
rect 13449 12325 13461 12359
rect 13495 12356 13507 12359
rect 13495 12328 14228 12356
rect 13495 12325 13507 12328
rect 13449 12319 13507 12325
rect 2501 12291 2559 12297
rect 2501 12257 2513 12291
rect 2547 12257 2559 12291
rect 2501 12251 2559 12257
rect 2593 12291 2651 12297
rect 2593 12257 2605 12291
rect 2639 12288 2651 12291
rect 2639 12260 3464 12288
rect 2639 12257 2651 12260
rect 2593 12251 2651 12257
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 2056 12152 2084 12183
rect 2682 12180 2688 12232
rect 2740 12180 2746 12232
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12220 2835 12223
rect 3326 12220 3332 12232
rect 2823 12192 3332 12220
rect 2823 12189 2835 12192
rect 2777 12183 2835 12189
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 2961 12155 3019 12161
rect 2961 12152 2973 12155
rect 2056 12124 2973 12152
rect 2961 12121 2973 12124
rect 3007 12121 3019 12155
rect 2961 12115 3019 12121
rect 3145 12155 3203 12161
rect 3145 12121 3157 12155
rect 3191 12152 3203 12155
rect 3436 12152 3464 12260
rect 5534 12248 5540 12300
rect 5592 12248 5598 12300
rect 5644 12260 9352 12288
rect 3878 12180 3884 12232
rect 3936 12220 3942 12232
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3936 12192 3985 12220
rect 3936 12180 3942 12192
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 4120 12192 5181 12220
rect 4120 12180 4126 12192
rect 5169 12189 5181 12192
rect 5215 12189 5227 12223
rect 5644 12220 5672 12260
rect 9324 12232 9352 12260
rect 10870 12248 10876 12300
rect 10928 12288 10934 12300
rect 11330 12288 11336 12300
rect 10928 12260 11336 12288
rect 10928 12248 10934 12260
rect 11330 12248 11336 12260
rect 11388 12288 11394 12300
rect 14093 12291 14151 12297
rect 14093 12288 14105 12291
rect 11388 12260 14105 12288
rect 11388 12248 11394 12260
rect 14093 12257 14105 12260
rect 14139 12257 14151 12291
rect 14200 12288 14228 12328
rect 14369 12291 14427 12297
rect 14369 12288 14381 12291
rect 14200 12260 14381 12288
rect 14093 12251 14151 12257
rect 14369 12257 14381 12260
rect 14415 12257 14427 12291
rect 14369 12251 14427 12257
rect 5169 12183 5227 12189
rect 5276 12192 5672 12220
rect 8757 12223 8815 12229
rect 5276 12152 5304 12192
rect 8757 12189 8769 12223
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 8772 12152 8800 12183
rect 9306 12180 9312 12232
rect 9364 12220 9370 12232
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 9364 12192 9873 12220
rect 9364 12180 9370 12192
rect 9861 12189 9873 12192
rect 9907 12220 9919 12223
rect 10962 12220 10968 12232
rect 9907 12192 10968 12220
rect 9907 12189 9919 12192
rect 9861 12183 9919 12189
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 12069 12223 12127 12229
rect 12069 12189 12081 12223
rect 12115 12189 12127 12223
rect 12069 12183 12127 12189
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 10134 12152 10140 12164
rect 3191 12124 5304 12152
rect 5828 12124 5934 12152
rect 8772 12124 10140 12152
rect 3191 12121 3203 12124
rect 3145 12115 3203 12121
rect 1857 12087 1915 12093
rect 1857 12053 1869 12087
rect 1903 12084 1915 12087
rect 1946 12084 1952 12096
rect 1903 12056 1952 12084
rect 1903 12053 1915 12056
rect 1857 12047 1915 12053
rect 1946 12044 1952 12056
rect 2004 12084 2010 12096
rect 2314 12084 2320 12096
rect 2004 12056 2320 12084
rect 2004 12044 2010 12056
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 3789 12087 3847 12093
rect 3789 12084 3801 12087
rect 3660 12056 3801 12084
rect 3660 12044 3666 12056
rect 3789 12053 3801 12056
rect 3835 12053 3847 12087
rect 3789 12047 3847 12053
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 5828 12084 5856 12124
rect 10134 12112 10140 12124
rect 10192 12112 10198 12164
rect 5500 12056 5856 12084
rect 5500 12044 5506 12056
rect 10410 12044 10416 12096
rect 10468 12044 10474 12096
rect 12084 12084 12112 12183
rect 12176 12152 12204 12183
rect 12250 12180 12256 12232
rect 12308 12180 12314 12232
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12220 12403 12223
rect 12802 12220 12808 12232
rect 12391 12192 12808 12220
rect 12391 12189 12403 12192
rect 12345 12183 12403 12189
rect 12802 12180 12808 12192
rect 12860 12220 12866 12232
rect 12897 12223 12955 12229
rect 12897 12220 12909 12223
rect 12860 12192 12909 12220
rect 12860 12180 12866 12192
rect 12897 12189 12909 12192
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12220 13323 12223
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 13311 12192 13553 12220
rect 13311 12189 13323 12192
rect 13265 12183 13323 12189
rect 13541 12189 13553 12192
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 12618 12152 12624 12164
rect 12176 12124 12624 12152
rect 12618 12112 12624 12124
rect 12676 12152 12682 12164
rect 12713 12155 12771 12161
rect 12713 12152 12725 12155
rect 12676 12124 12725 12152
rect 12676 12112 12682 12124
rect 12713 12121 12725 12124
rect 12759 12121 12771 12155
rect 13740 12152 13768 12183
rect 13814 12180 13820 12232
rect 13872 12180 13878 12232
rect 14274 12152 14280 12164
rect 13740 12124 14280 12152
rect 12713 12115 12771 12121
rect 14274 12112 14280 12124
rect 14332 12112 14338 12164
rect 15378 12112 15384 12164
rect 15436 12112 15442 12164
rect 13446 12084 13452 12096
rect 12084 12056 13452 12084
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 15010 12044 15016 12096
rect 15068 12084 15074 12096
rect 15841 12087 15899 12093
rect 15841 12084 15853 12087
rect 15068 12056 15853 12084
rect 15068 12044 15074 12056
rect 15841 12053 15853 12056
rect 15887 12053 15899 12087
rect 15841 12047 15899 12053
rect 1104 11994 16836 12016
rect 1104 11942 1610 11994
rect 1662 11942 1674 11994
rect 1726 11942 1738 11994
rect 1790 11942 1802 11994
rect 1854 11942 1866 11994
rect 1918 11942 5610 11994
rect 5662 11942 5674 11994
rect 5726 11942 5738 11994
rect 5790 11942 5802 11994
rect 5854 11942 5866 11994
rect 5918 11942 9610 11994
rect 9662 11942 9674 11994
rect 9726 11942 9738 11994
rect 9790 11942 9802 11994
rect 9854 11942 9866 11994
rect 9918 11942 13610 11994
rect 13662 11942 13674 11994
rect 13726 11942 13738 11994
rect 13790 11942 13802 11994
rect 13854 11942 13866 11994
rect 13918 11942 16836 11994
rect 1104 11920 16836 11942
rect 4522 11840 4528 11892
rect 4580 11880 4586 11892
rect 5031 11883 5089 11889
rect 5031 11880 5043 11883
rect 4580 11852 5043 11880
rect 4580 11840 4586 11852
rect 5031 11849 5043 11852
rect 5077 11849 5089 11883
rect 12526 11880 12532 11892
rect 5031 11843 5089 11849
rect 12360 11852 12532 11880
rect 5442 11812 5448 11824
rect 4646 11798 5448 11812
rect 4632 11784 5448 11798
rect 3234 11704 3240 11756
rect 3292 11744 3298 11756
rect 3292 11716 3740 11744
rect 3292 11704 3298 11716
rect 3602 11636 3608 11688
rect 3660 11636 3666 11688
rect 3712 11676 3740 11716
rect 4062 11676 4068 11688
rect 3712 11648 4068 11676
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4154 11636 4160 11688
rect 4212 11676 4218 11688
rect 4632 11676 4660 11784
rect 5442 11772 5448 11784
rect 5500 11772 5506 11824
rect 7466 11812 7472 11824
rect 5828 11784 7472 11812
rect 5828 11753 5856 11784
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 9490 11772 9496 11824
rect 9548 11772 9554 11824
rect 9953 11815 10011 11821
rect 9953 11781 9965 11815
rect 9999 11812 10011 11815
rect 10042 11812 10048 11824
rect 9999 11784 10048 11812
rect 9999 11781 10011 11784
rect 9953 11775 10011 11781
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 7190 11704 7196 11756
rect 7248 11704 7254 11756
rect 12360 11753 12388 11852
rect 12526 11840 12532 11852
rect 12584 11840 12590 11892
rect 13909 11883 13967 11889
rect 13909 11849 13921 11883
rect 13955 11880 13967 11883
rect 14274 11880 14280 11892
rect 13955 11852 14280 11880
rect 13955 11849 13967 11852
rect 13909 11843 13967 11849
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 15102 11840 15108 11892
rect 15160 11840 15166 11892
rect 12897 11815 12955 11821
rect 12897 11781 12909 11815
rect 12943 11812 12955 11815
rect 14090 11812 14096 11824
rect 12943 11784 14096 11812
rect 12943 11781 12955 11784
rect 12897 11775 12955 11781
rect 14090 11772 14096 11784
rect 14148 11772 14154 11824
rect 14737 11815 14795 11821
rect 14737 11781 14749 11815
rect 14783 11812 14795 11815
rect 14783 11784 15056 11812
rect 14783 11781 14795 11784
rect 14737 11775 14795 11781
rect 15028 11756 15056 11784
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11744 14243 11747
rect 14921 11747 14979 11753
rect 14921 11744 14933 11747
rect 14231 11716 14504 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 4212 11648 4660 11676
rect 5905 11679 5963 11685
rect 4212 11636 4218 11648
rect 5905 11645 5917 11679
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 6181 11679 6239 11685
rect 6181 11645 6193 11679
rect 6227 11676 6239 11679
rect 7101 11679 7159 11685
rect 7101 11676 7113 11679
rect 6227 11648 7113 11676
rect 6227 11645 6239 11648
rect 6181 11639 6239 11645
rect 7101 11645 7113 11648
rect 7147 11645 7159 11679
rect 7101 11639 7159 11645
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 11330 11676 11336 11688
rect 10275 11648 11336 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 5920 11608 5948 11639
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11480 11648 12081 11676
rect 11480 11636 11486 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 12250 11636 12256 11688
rect 12308 11676 12314 11688
rect 12820 11676 12848 11707
rect 12308 11648 12848 11676
rect 12308 11636 12314 11648
rect 6730 11608 6736 11620
rect 5920 11580 6736 11608
rect 6730 11568 6736 11580
rect 6788 11568 6794 11620
rect 6822 11568 6828 11620
rect 6880 11568 6886 11620
rect 12710 11568 12716 11620
rect 12768 11608 12774 11620
rect 13096 11608 13124 11707
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 14093 11679 14151 11685
rect 14093 11676 14105 11679
rect 13504 11648 14105 11676
rect 13504 11636 13510 11648
rect 14093 11645 14105 11648
rect 14139 11645 14151 11679
rect 14277 11679 14335 11685
rect 14277 11676 14289 11679
rect 14093 11639 14151 11645
rect 14200 11648 14289 11676
rect 12768 11580 13124 11608
rect 12768 11568 12774 11580
rect 14200 11552 14228 11648
rect 14277 11645 14289 11648
rect 14323 11645 14335 11679
rect 14277 11639 14335 11645
rect 14369 11679 14427 11685
rect 14369 11645 14381 11679
rect 14415 11645 14427 11679
rect 14476 11676 14504 11716
rect 14844 11716 14933 11744
rect 14844 11688 14872 11716
rect 14921 11713 14933 11716
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 15010 11704 15016 11756
rect 15068 11704 15074 11756
rect 14826 11676 14832 11688
rect 14476 11648 14832 11676
rect 14369 11639 14427 11645
rect 14384 11608 14412 11639
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 15028 11608 15056 11704
rect 14384 11580 15056 11608
rect 3234 11500 3240 11552
rect 3292 11540 3298 11552
rect 8478 11540 8484 11552
rect 3292 11512 8484 11540
rect 3292 11500 3298 11512
rect 8478 11500 8484 11512
rect 8536 11500 8542 11552
rect 13265 11543 13323 11549
rect 13265 11509 13277 11543
rect 13311 11540 13323 11543
rect 13354 11540 13360 11552
rect 13311 11512 13360 11540
rect 13311 11509 13323 11512
rect 13265 11503 13323 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 14182 11500 14188 11552
rect 14240 11500 14246 11552
rect 944 11450 16836 11472
rect 944 11398 950 11450
rect 1002 11398 1014 11450
rect 1066 11398 1078 11450
rect 1130 11398 1142 11450
rect 1194 11398 1206 11450
rect 1258 11398 4950 11450
rect 5002 11398 5014 11450
rect 5066 11398 5078 11450
rect 5130 11398 5142 11450
rect 5194 11398 5206 11450
rect 5258 11398 8950 11450
rect 9002 11398 9014 11450
rect 9066 11398 9078 11450
rect 9130 11398 9142 11450
rect 9194 11398 9206 11450
rect 9258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 16836 11450
rect 944 11376 16836 11398
rect 2866 11296 2872 11348
rect 2924 11296 2930 11348
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 3200 11308 3433 11336
rect 3200 11296 3206 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 3878 11296 3884 11348
rect 3936 11296 3942 11348
rect 6549 11339 6607 11345
rect 6549 11305 6561 11339
rect 6595 11336 6607 11339
rect 6730 11336 6736 11348
rect 6595 11308 6736 11336
rect 6595 11305 6607 11308
rect 6549 11299 6607 11305
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 8573 11339 8631 11345
rect 8573 11336 8585 11339
rect 8536 11308 8585 11336
rect 8536 11296 8542 11308
rect 8573 11305 8585 11308
rect 8619 11305 8631 11339
rect 8573 11299 8631 11305
rect 2884 11268 2912 11296
rect 2608 11240 3464 11268
rect 2608 11209 2636 11240
rect 2409 11203 2467 11209
rect 2409 11200 2421 11203
rect 2148 11172 2421 11200
rect 2148 11141 2176 11172
rect 2409 11169 2421 11172
rect 2455 11169 2467 11203
rect 2409 11163 2467 11169
rect 2593 11203 2651 11209
rect 2593 11169 2605 11203
rect 2639 11169 2651 11203
rect 2593 11163 2651 11169
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 2731 11172 3188 11200
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 1949 11135 2007 11141
rect 1949 11132 1961 11135
rect 1903 11104 1961 11132
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 1949 11101 1961 11104
rect 1995 11101 2007 11135
rect 1949 11095 2007 11101
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 2222 11092 2228 11144
rect 2280 11092 2286 11144
rect 2774 11092 2780 11144
rect 2832 11092 2838 11144
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 2884 11064 2912 11095
rect 2958 11064 2964 11076
rect 2884 11036 2964 11064
rect 2958 11024 2964 11036
rect 3016 11064 3022 11076
rect 3053 11067 3111 11073
rect 3053 11064 3065 11067
rect 3016 11036 3065 11064
rect 3016 11024 3022 11036
rect 3053 11033 3065 11036
rect 3099 11033 3111 11067
rect 3160 11064 3188 11172
rect 3436 11076 3464 11240
rect 6362 11228 6368 11280
rect 6420 11268 6426 11280
rect 7469 11271 7527 11277
rect 7469 11268 7481 11271
rect 6420 11240 7481 11268
rect 6420 11228 6426 11240
rect 7469 11237 7481 11240
rect 7515 11237 7527 11271
rect 7469 11231 7527 11237
rect 4338 11160 4344 11212
rect 4396 11160 4402 11212
rect 4522 11160 4528 11212
rect 4580 11160 4586 11212
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 8588 11200 8616 11299
rect 10410 11296 10416 11348
rect 10468 11296 10474 11348
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 10689 11339 10747 11345
rect 10689 11336 10701 11339
rect 10652 11308 10701 11336
rect 10652 11296 10658 11308
rect 10689 11305 10701 11308
rect 10735 11305 10747 11339
rect 10689 11299 10747 11305
rect 12618 11296 12624 11348
rect 12676 11336 12682 11348
rect 12713 11339 12771 11345
rect 12713 11336 12725 11339
rect 12676 11308 12725 11336
rect 12676 11296 12682 11308
rect 12713 11305 12725 11308
rect 12759 11305 12771 11339
rect 12713 11299 12771 11305
rect 10318 11228 10324 11280
rect 10376 11228 10382 11280
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 4847 11172 6868 11200
rect 8588 11172 9321 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4816 11132 4844 11163
rect 4120 11104 4844 11132
rect 4120 11092 4126 11104
rect 6730 11092 6736 11144
rect 6788 11092 6794 11144
rect 3234 11064 3240 11076
rect 3160 11036 3240 11064
rect 3053 11027 3111 11033
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 3418 11024 3424 11076
rect 3476 11024 3482 11076
rect 5074 11024 5080 11076
rect 5132 11024 5138 11076
rect 6638 11064 6644 11076
rect 6302 11036 6644 11064
rect 6638 11024 6644 11036
rect 6696 11024 6702 11076
rect 1486 10956 1492 11008
rect 1544 10996 1550 11008
rect 1673 10999 1731 11005
rect 1673 10996 1685 10999
rect 1544 10968 1685 10996
rect 1544 10956 1550 10968
rect 1673 10965 1685 10968
rect 1719 10965 1731 10999
rect 1673 10959 1731 10965
rect 4246 10956 4252 11008
rect 4304 10956 4310 11008
rect 6840 10996 6868 11172
rect 9309 11169 9321 11172
rect 9355 11169 9367 11203
rect 10336 11200 10364 11228
rect 9309 11163 9367 11169
rect 10244 11172 10364 11200
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11132 7343 11135
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 7331 11104 7389 11132
rect 7331 11101 7343 11104
rect 7285 11095 7343 11101
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 9398 11132 9404 11144
rect 7377 11095 7435 11101
rect 8680 11104 9404 11132
rect 8389 11067 8447 11073
rect 8389 11033 8401 11067
rect 8435 11064 8447 11067
rect 8478 11064 8484 11076
rect 8435 11036 8484 11064
rect 8435 11033 8447 11036
rect 8389 11027 8447 11033
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 8589 11067 8647 11073
rect 8589 11033 8601 11067
rect 8635 11064 8647 11067
rect 8680 11064 8708 11104
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 10244 11141 10272 11172
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 10428 11132 10456 11296
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 11330 11200 11336 11212
rect 11011 11172 11336 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 12728 11200 12756 11299
rect 14090 11296 14096 11348
rect 14148 11296 14154 11348
rect 13357 11203 13415 11209
rect 13357 11200 13369 11203
rect 12728 11172 13369 11200
rect 13357 11169 13369 11172
rect 13403 11169 13415 11203
rect 13357 11163 13415 11169
rect 16393 11203 16451 11209
rect 16393 11169 16405 11203
rect 16439 11200 16451 11203
rect 16482 11200 16488 11212
rect 16439 11172 16488 11200
rect 16439 11169 16451 11172
rect 16393 11163 16451 11169
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 10367 11104 10456 11132
rect 10505 11135 10563 11141
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 10505 11101 10517 11135
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 14737 11135 14795 11141
rect 14737 11101 14749 11135
rect 14783 11132 14795 11135
rect 14826 11132 14832 11144
rect 14783 11104 14832 11132
rect 14783 11101 14795 11104
rect 14737 11095 14795 11101
rect 10520 11064 10548 11095
rect 14826 11092 14832 11104
rect 14884 11092 14890 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15120 11104 15761 11132
rect 15120 11076 15148 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 8635 11036 8708 11064
rect 8772 11036 10548 11064
rect 8635 11033 8647 11036
rect 8589 11027 8647 11033
rect 7006 10996 7012 11008
rect 6840 10968 7012 10996
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 8772 11005 8800 11036
rect 11238 11024 11244 11076
rect 11296 11024 11302 11076
rect 12466 11036 12940 11064
rect 12912 11008 12940 11036
rect 15102 11024 15108 11076
rect 15160 11024 15166 11076
rect 15841 11067 15899 11073
rect 15841 11033 15853 11067
rect 15887 11064 15899 11067
rect 16117 11067 16175 11073
rect 16117 11064 16129 11067
rect 15887 11036 16129 11064
rect 15887 11033 15899 11036
rect 15841 11027 15899 11033
rect 16117 11033 16129 11036
rect 16163 11033 16175 11067
rect 16117 11027 16175 11033
rect 8757 10999 8815 11005
rect 8757 10965 8769 10999
rect 8803 10965 8815 10999
rect 8757 10959 8815 10965
rect 9950 10956 9956 11008
rect 10008 10956 10014 11008
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 11422 10996 11428 11008
rect 10652 10968 11428 10996
rect 10652 10956 10658 10968
rect 11422 10956 11428 10968
rect 11480 10956 11486 11008
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 12526 10996 12532 11008
rect 12124 10968 12532 10996
rect 12124 10956 12130 10968
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 12802 10956 12808 11008
rect 12860 10956 12866 11008
rect 12894 10956 12900 11008
rect 12952 10956 12958 11008
rect 1104 10906 16836 10928
rect 1104 10854 1610 10906
rect 1662 10854 1674 10906
rect 1726 10854 1738 10906
rect 1790 10854 1802 10906
rect 1854 10854 1866 10906
rect 1918 10854 5610 10906
rect 5662 10854 5674 10906
rect 5726 10854 5738 10906
rect 5790 10854 5802 10906
rect 5854 10854 5866 10906
rect 5918 10854 9610 10906
rect 9662 10854 9674 10906
rect 9726 10854 9738 10906
rect 9790 10854 9802 10906
rect 9854 10854 9866 10906
rect 9918 10854 13610 10906
rect 13662 10854 13674 10906
rect 13726 10854 13738 10906
rect 13790 10854 13802 10906
rect 13854 10854 13866 10906
rect 13918 10854 16836 10906
rect 1104 10832 16836 10854
rect 1486 10752 1492 10804
rect 1544 10752 1550 10804
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4396 10764 4537 10792
rect 4396 10752 4402 10764
rect 4525 10761 4537 10764
rect 4571 10792 4583 10795
rect 4571 10764 5028 10792
rect 4571 10761 4583 10764
rect 4525 10755 4583 10761
rect 1504 10724 1532 10752
rect 5000 10733 5028 10764
rect 5350 10752 5356 10804
rect 5408 10752 5414 10804
rect 6917 10795 6975 10801
rect 6917 10761 6929 10795
rect 6963 10761 6975 10795
rect 9306 10792 9312 10804
rect 6917 10755 6975 10761
rect 8588 10764 9312 10792
rect 1673 10727 1731 10733
rect 1673 10724 1685 10727
rect 1504 10696 1685 10724
rect 1673 10693 1685 10696
rect 1719 10693 1731 10727
rect 1673 10687 1731 10693
rect 4985 10727 5043 10733
rect 4985 10693 4997 10727
rect 5031 10693 5043 10727
rect 5368 10724 5396 10752
rect 4985 10687 5043 10693
rect 5092 10696 5396 10724
rect 6932 10724 6960 10755
rect 8588 10736 8616 10764
rect 9306 10752 9312 10764
rect 9364 10792 9370 10804
rect 9364 10764 11192 10792
rect 9364 10752 9370 10764
rect 7285 10727 7343 10733
rect 7285 10724 7297 10727
rect 6932 10696 7297 10724
rect 3326 10656 3332 10668
rect 2806 10628 3332 10656
rect 3326 10616 3332 10628
rect 3384 10616 3390 10668
rect 4246 10616 4252 10668
rect 4304 10656 4310 10668
rect 4341 10659 4399 10665
rect 4341 10656 4353 10659
rect 4304 10628 4353 10656
rect 4304 10616 4310 10628
rect 4341 10625 4353 10628
rect 4387 10656 4399 10659
rect 5092 10656 5120 10696
rect 7285 10693 7297 10696
rect 7331 10693 7343 10727
rect 7285 10687 7343 10693
rect 8570 10684 8576 10736
rect 8628 10684 8634 10736
rect 9398 10684 9404 10736
rect 9456 10724 9462 10736
rect 10410 10733 10416 10736
rect 10392 10727 10416 10733
rect 10392 10724 10404 10727
rect 9456 10696 10404 10724
rect 9456 10684 9462 10696
rect 10392 10693 10404 10696
rect 10468 10724 10474 10736
rect 10612 10733 10640 10764
rect 11164 10733 11192 10764
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 11296 10764 11805 10792
rect 11296 10752 11302 10764
rect 11793 10761 11805 10764
rect 11839 10761 11851 10795
rect 11793 10755 11851 10761
rect 12066 10752 12072 10804
rect 12124 10752 12130 10804
rect 12161 10795 12219 10801
rect 12161 10761 12173 10795
rect 12207 10792 12219 10795
rect 12802 10792 12808 10804
rect 12207 10764 12808 10792
rect 12207 10761 12219 10764
rect 12161 10755 12219 10761
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 13998 10752 14004 10804
rect 14056 10792 14062 10804
rect 15102 10792 15108 10804
rect 14056 10764 15108 10792
rect 14056 10752 14062 10764
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 10597 10727 10655 10733
rect 10468 10696 10548 10724
rect 10392 10687 10416 10693
rect 10410 10684 10416 10687
rect 10468 10684 10474 10696
rect 4387 10628 5120 10656
rect 5353 10659 5411 10665
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 5353 10625 5365 10659
rect 5399 10656 5411 10659
rect 6362 10656 6368 10668
rect 5399 10628 6368 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 6914 10656 6920 10668
rect 6779 10628 6920 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 8294 10616 8300 10668
rect 8352 10656 8358 10668
rect 9861 10659 9919 10665
rect 8352 10628 8418 10656
rect 8352 10616 8358 10628
rect 9861 10625 9873 10659
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 1394 10548 1400 10600
rect 1452 10548 1458 10600
rect 4709 10591 4767 10597
rect 4709 10557 4721 10591
rect 4755 10588 4767 10591
rect 4798 10588 4804 10600
rect 4755 10560 4804 10588
rect 4755 10557 4767 10560
rect 4709 10551 4767 10557
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 5169 10591 5227 10597
rect 5169 10557 5181 10591
rect 5215 10588 5227 10591
rect 6822 10588 6828 10600
rect 5215 10560 6828 10588
rect 5215 10557 5227 10560
rect 5169 10551 5227 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7006 10548 7012 10600
rect 7064 10548 7070 10600
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10588 8815 10591
rect 9398 10588 9404 10600
rect 8803 10560 9404 10588
rect 8803 10557 8815 10560
rect 8757 10551 8815 10557
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 9876 10588 9904 10619
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10045 10659 10103 10665
rect 10045 10656 10057 10659
rect 10008 10628 10057 10656
rect 10008 10616 10014 10628
rect 10045 10625 10057 10628
rect 10091 10625 10103 10659
rect 10045 10619 10103 10625
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10656 10195 10659
rect 10520 10656 10548 10696
rect 10597 10693 10609 10727
rect 10643 10693 10655 10727
rect 11149 10727 11207 10733
rect 10597 10687 10655 10693
rect 10919 10693 10977 10699
rect 10919 10659 10931 10693
rect 10965 10659 10977 10693
rect 11149 10693 11161 10727
rect 11195 10724 11207 10727
rect 11606 10724 11612 10736
rect 11195 10696 11612 10724
rect 11195 10693 11207 10696
rect 11149 10687 11207 10693
rect 11606 10684 11612 10696
rect 11664 10684 11670 10736
rect 10919 10656 10977 10659
rect 10183 10628 10364 10656
rect 10520 10653 10977 10656
rect 11977 10659 12035 10665
rect 10520 10628 10976 10653
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 10336 10600 10364 10628
rect 11977 10625 11989 10659
rect 12023 10656 12035 10659
rect 12084 10656 12112 10752
rect 12023 10628 12112 10656
rect 12250 10684 12256 10736
rect 12308 10684 12314 10736
rect 12345 10727 12403 10733
rect 12345 10693 12357 10727
rect 12391 10693 12403 10727
rect 12345 10687 12403 10693
rect 12575 10693 12633 10699
rect 12575 10690 12587 10693
rect 12250 10681 12308 10684
rect 12250 10647 12262 10681
rect 12296 10647 12308 10681
rect 12250 10641 12308 10647
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 9876 10560 10272 10588
rect 5074 10480 5080 10532
rect 5132 10520 5138 10532
rect 5261 10523 5319 10529
rect 5132 10492 5212 10520
rect 5132 10480 5138 10492
rect 2958 10412 2964 10464
rect 3016 10452 3022 10464
rect 3145 10455 3203 10461
rect 3145 10452 3157 10455
rect 3016 10424 3157 10452
rect 3016 10412 3022 10424
rect 3145 10421 3157 10424
rect 3191 10421 3203 10455
rect 3145 10415 3203 10421
rect 4706 10412 4712 10464
rect 4764 10412 4770 10464
rect 5184 10461 5212 10492
rect 5261 10489 5273 10523
rect 5307 10520 5319 10523
rect 5350 10520 5356 10532
rect 5307 10492 5356 10520
rect 5307 10489 5319 10492
rect 5261 10483 5319 10489
rect 5350 10480 5356 10492
rect 5408 10480 5414 10532
rect 9677 10523 9735 10529
rect 9677 10489 9689 10523
rect 9723 10520 9735 10523
rect 10042 10520 10048 10532
rect 9723 10492 10048 10520
rect 9723 10489 9735 10492
rect 9677 10483 9735 10489
rect 10042 10480 10048 10492
rect 10100 10480 10106 10532
rect 10244 10529 10272 10560
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 11698 10588 11704 10600
rect 10376 10560 11704 10588
rect 10376 10548 10382 10560
rect 11698 10548 11704 10560
rect 11756 10588 11762 10600
rect 12268 10588 12296 10641
rect 11756 10560 12296 10588
rect 11756 10548 11762 10560
rect 10229 10523 10287 10529
rect 10229 10489 10241 10523
rect 10275 10489 10287 10523
rect 11514 10520 11520 10532
rect 10229 10483 10287 10489
rect 10428 10492 11520 10520
rect 5169 10455 5227 10461
rect 5169 10421 5181 10455
rect 5215 10421 5227 10455
rect 5169 10415 5227 10421
rect 8846 10412 8852 10464
rect 8904 10412 8910 10464
rect 10428 10461 10456 10492
rect 11514 10480 11520 10492
rect 11572 10480 11578 10532
rect 11606 10480 11612 10532
rect 11664 10520 11670 10532
rect 12360 10520 12388 10687
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 12560 10659 12587 10690
rect 12621 10659 12633 10693
rect 13354 10684 13360 10736
rect 13412 10684 13418 10736
rect 15378 10724 15384 10736
rect 14582 10696 15384 10724
rect 15378 10684 15384 10696
rect 15436 10684 15442 10736
rect 12560 10656 12633 10659
rect 12492 10653 12633 10656
rect 12492 10628 12588 10653
rect 12492 10616 12498 10628
rect 14918 10616 14924 10668
rect 14976 10616 14982 10668
rect 13081 10591 13139 10597
rect 13081 10557 13093 10591
rect 13127 10557 13139 10591
rect 13081 10551 13139 10557
rect 11664 10492 12388 10520
rect 11664 10480 11670 10492
rect 12710 10480 12716 10532
rect 12768 10480 12774 10532
rect 10413 10455 10471 10461
rect 10413 10421 10425 10455
rect 10459 10421 10471 10455
rect 10413 10415 10471 10421
rect 10778 10412 10784 10464
rect 10836 10412 10842 10464
rect 10962 10412 10968 10464
rect 11020 10412 11026 10464
rect 12529 10455 12587 10461
rect 12529 10421 12541 10455
rect 12575 10452 12587 10455
rect 12618 10452 12624 10464
rect 12575 10424 12624 10452
rect 12575 10421 12587 10424
rect 12529 10415 12587 10421
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 13096 10452 13124 10551
rect 13538 10452 13544 10464
rect 13096 10424 13544 10452
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 14826 10412 14832 10464
rect 14884 10412 14890 10464
rect 944 10362 16836 10384
rect 944 10310 950 10362
rect 1002 10310 1014 10362
rect 1066 10310 1078 10362
rect 1130 10310 1142 10362
rect 1194 10310 1206 10362
rect 1258 10310 4950 10362
rect 5002 10310 5014 10362
rect 5066 10310 5078 10362
rect 5130 10310 5142 10362
rect 5194 10310 5206 10362
rect 5258 10310 8950 10362
rect 9002 10310 9014 10362
rect 9066 10310 9078 10362
rect 9130 10310 9142 10362
rect 9194 10310 9206 10362
rect 9258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 16836 10362
rect 944 10288 16836 10310
rect 934 10208 940 10260
rect 992 10248 998 10260
rect 1489 10251 1547 10257
rect 1489 10248 1501 10251
rect 992 10220 1501 10248
rect 992 10208 998 10220
rect 1489 10217 1501 10220
rect 1535 10217 1547 10251
rect 1489 10211 1547 10217
rect 6270 10208 6276 10260
rect 6328 10248 6334 10260
rect 6733 10251 6791 10257
rect 6733 10248 6745 10251
rect 6328 10220 6745 10248
rect 6328 10208 6334 10220
rect 6733 10217 6745 10220
rect 6779 10217 6791 10251
rect 6733 10211 6791 10217
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 6972 10220 7021 10248
rect 6972 10208 6978 10220
rect 7009 10217 7021 10220
rect 7055 10217 7067 10251
rect 7009 10211 7067 10217
rect 8846 10208 8852 10260
rect 8904 10208 8910 10260
rect 9398 10208 9404 10260
rect 9456 10208 9462 10260
rect 10045 10251 10103 10257
rect 10045 10217 10057 10251
rect 10091 10248 10103 10251
rect 10134 10248 10140 10260
rect 10091 10220 10140 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 10778 10208 10784 10260
rect 10836 10208 10842 10260
rect 11514 10208 11520 10260
rect 11572 10248 11578 10260
rect 14826 10248 14832 10260
rect 11572 10220 14832 10248
rect 11572 10208 11578 10220
rect 14826 10208 14832 10220
rect 14884 10208 14890 10260
rect 14918 10208 14924 10260
rect 14976 10208 14982 10260
rect 4798 10072 4804 10124
rect 4856 10072 4862 10124
rect 6914 10072 6920 10124
rect 6972 10072 6978 10124
rect 7558 10072 7564 10124
rect 7616 10072 7622 10124
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10044 1823 10047
rect 1811 10016 2774 10044
rect 1811 10013 1823 10016
rect 1765 10007 1823 10013
rect 2746 9908 2774 10016
rect 4614 10004 4620 10056
rect 4672 10004 4678 10056
rect 4816 10044 4844 10072
rect 5350 10044 5356 10056
rect 4816 10016 5356 10044
rect 5350 10004 5356 10016
rect 5408 10044 5414 10056
rect 6641 10047 6699 10053
rect 6641 10044 6653 10047
rect 5408 10016 6653 10044
rect 5408 10004 5414 10016
rect 6641 10013 6653 10016
rect 6687 10044 6699 10047
rect 6822 10044 6828 10056
rect 6687 10016 6828 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7377 10047 7435 10053
rect 7377 10013 7389 10047
rect 7423 10044 7435 10047
rect 8864 10044 8892 10208
rect 9416 10112 9444 10208
rect 9416 10084 9720 10112
rect 7423 10016 8892 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 9490 10004 9496 10056
rect 9548 10004 9554 10056
rect 9692 10053 9720 10084
rect 10318 10072 10324 10124
rect 10376 10112 10382 10124
rect 10376 10084 10732 10112
rect 10376 10072 10382 10084
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10013 9735 10047
rect 10594 10044 10600 10056
rect 9677 10007 9735 10013
rect 9784 10016 10600 10044
rect 6917 9979 6975 9985
rect 6917 9945 6929 9979
rect 6963 9976 6975 9979
rect 7469 9979 7527 9985
rect 7469 9976 7481 9979
rect 6963 9948 7481 9976
rect 6963 9945 6975 9948
rect 6917 9939 6975 9945
rect 7469 9945 7481 9948
rect 7515 9945 7527 9979
rect 9784 9976 9812 10016
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 10704 10053 10732 10084
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10013 10747 10047
rect 10796 10044 10824 10208
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10112 11207 10115
rect 11517 10115 11575 10121
rect 11517 10112 11529 10115
rect 11195 10084 11529 10112
rect 11195 10081 11207 10084
rect 11149 10075 11207 10081
rect 11517 10081 11529 10084
rect 11563 10081 11575 10115
rect 11517 10075 11575 10081
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10796 10016 10977 10044
rect 10689 10007 10747 10013
rect 10965 10013 10977 10016
rect 11011 10013 11023 10047
rect 10965 10007 11023 10013
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10013 11299 10047
rect 12802 10044 12808 10056
rect 12650 10030 12808 10044
rect 11241 10007 11299 10013
rect 12636 10016 12808 10030
rect 7469 9939 7527 9945
rect 7576 9948 9812 9976
rect 9861 9979 9919 9985
rect 7576 9908 7604 9948
rect 9861 9945 9873 9979
rect 9907 9976 9919 9979
rect 10318 9976 10324 9988
rect 9907 9948 10324 9976
rect 9907 9945 9919 9948
rect 9861 9939 9919 9945
rect 10318 9936 10324 9948
rect 10376 9936 10382 9988
rect 11256 9976 11284 10007
rect 11256 9948 11376 9976
rect 11348 9920 11376 9948
rect 2746 9880 7604 9908
rect 7650 9868 7656 9920
rect 7708 9908 7714 9920
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 7708 9880 8953 9908
rect 7708 9868 7714 9880
rect 8941 9877 8953 9880
rect 8987 9877 8999 9911
rect 8941 9871 8999 9877
rect 10781 9911 10839 9917
rect 10781 9877 10793 9911
rect 10827 9908 10839 9911
rect 11238 9908 11244 9920
rect 10827 9880 11244 9908
rect 10827 9877 10839 9880
rect 10781 9871 10839 9877
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 11330 9868 11336 9920
rect 11388 9868 11394 9920
rect 11514 9868 11520 9920
rect 11572 9908 11578 9920
rect 12636 9908 12664 10016
rect 12802 10004 12808 10016
rect 12860 10044 12866 10056
rect 15378 10044 15384 10056
rect 12860 10016 15384 10044
rect 12860 10004 12866 10016
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 14550 9936 14556 9988
rect 14608 9936 14614 9988
rect 14737 9979 14795 9985
rect 14737 9945 14749 9979
rect 14783 9945 14795 9979
rect 14737 9939 14795 9945
rect 11572 9880 12664 9908
rect 12989 9911 13047 9917
rect 11572 9868 11578 9880
rect 12989 9877 13001 9911
rect 13035 9908 13047 9911
rect 13446 9908 13452 9920
rect 13035 9880 13452 9908
rect 13035 9877 13047 9880
rect 12989 9871 13047 9877
rect 13446 9868 13452 9880
rect 13504 9908 13510 9920
rect 14752 9908 14780 9939
rect 13504 9880 14780 9908
rect 13504 9868 13510 9880
rect 1104 9818 16836 9840
rect 1104 9766 1610 9818
rect 1662 9766 1674 9818
rect 1726 9766 1738 9818
rect 1790 9766 1802 9818
rect 1854 9766 1866 9818
rect 1918 9766 5610 9818
rect 5662 9766 5674 9818
rect 5726 9766 5738 9818
rect 5790 9766 5802 9818
rect 5854 9766 5866 9818
rect 5918 9766 9610 9818
rect 9662 9766 9674 9818
rect 9726 9766 9738 9818
rect 9790 9766 9802 9818
rect 9854 9766 9866 9818
rect 9918 9766 13610 9818
rect 13662 9766 13674 9818
rect 13726 9766 13738 9818
rect 13790 9766 13802 9818
rect 13854 9766 13866 9818
rect 13918 9766 16836 9818
rect 1104 9744 16836 9766
rect 6914 9664 6920 9716
rect 6972 9664 6978 9716
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 11296 9676 12020 9704
rect 11296 9664 11302 9676
rect 2130 9596 2136 9648
rect 2188 9636 2194 9648
rect 6932 9636 6960 9664
rect 2188 9608 2530 9636
rect 3344 9608 4292 9636
rect 2188 9596 2194 9608
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 1765 9571 1823 9577
rect 1765 9568 1777 9571
rect 1452 9540 1777 9568
rect 1452 9528 1458 9540
rect 1765 9537 1777 9540
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 1780 9364 1808 9531
rect 3344 9512 3372 9608
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4157 9571 4215 9577
rect 4157 9568 4169 9571
rect 4120 9540 4169 9568
rect 4120 9528 4126 9540
rect 4157 9537 4169 9540
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 2038 9460 2044 9512
rect 2096 9460 2102 9512
rect 2130 9460 2136 9512
rect 2188 9500 2194 9512
rect 3326 9500 3332 9512
rect 2188 9472 3332 9500
rect 2188 9460 2194 9472
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 4080 9432 4108 9528
rect 4264 9500 4292 9608
rect 4525 9571 4583 9577
rect 4525 9537 4537 9571
rect 4571 9568 4583 9571
rect 4614 9568 4620 9580
rect 4571 9540 4620 9568
rect 4571 9537 4583 9540
rect 4525 9531 4583 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 5276 9568 5304 9622
rect 6563 9608 7420 9636
rect 5442 9568 5448 9580
rect 5276 9540 5448 9568
rect 5276 9500 5304 9540
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 6563 9577 6591 9608
rect 7392 9580 7420 9608
rect 8846 9596 8852 9648
rect 8904 9636 8910 9648
rect 8941 9639 8999 9645
rect 8941 9636 8953 9639
rect 8904 9608 8953 9636
rect 8904 9596 8910 9608
rect 8941 9605 8953 9608
rect 8987 9605 8999 9639
rect 8941 9599 8999 9605
rect 9398 9596 9404 9648
rect 9456 9596 9462 9648
rect 11992 9645 12020 9676
rect 11977 9639 12035 9645
rect 11977 9605 11989 9639
rect 12023 9605 12035 9639
rect 11977 9599 12035 9605
rect 13262 9596 13268 9648
rect 13320 9636 13326 9648
rect 13630 9636 13636 9648
rect 13320 9608 13636 9636
rect 13320 9596 13326 9608
rect 13630 9596 13636 9608
rect 13688 9596 13694 9648
rect 15378 9596 15384 9648
rect 15436 9596 15442 9648
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 6328 9540 6377 9568
rect 6328 9528 6334 9540
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 6548 9571 6606 9577
rect 6548 9537 6560 9571
rect 6594 9537 6606 9571
rect 6548 9531 6606 9537
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 6822 9528 6828 9580
rect 6880 9568 6886 9580
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 6880 9540 6929 9568
rect 6880 9528 6886 9540
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 8662 9528 8668 9580
rect 8720 9528 8726 9580
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 13173 9571 13231 9577
rect 12676 9540 13124 9568
rect 12676 9528 12682 9540
rect 4264 9472 5304 9500
rect 3436 9404 4108 9432
rect 5276 9432 5304 9472
rect 5951 9503 6009 9509
rect 5951 9469 5963 9503
rect 5997 9500 6009 9503
rect 6641 9503 6699 9509
rect 6641 9500 6653 9503
rect 5997 9472 6653 9500
rect 5997 9469 6009 9472
rect 5951 9463 6009 9469
rect 6564 9444 6592 9472
rect 6641 9469 6653 9472
rect 6687 9469 6699 9503
rect 6641 9463 6699 9469
rect 11057 9503 11115 9509
rect 11057 9469 11069 9503
rect 11103 9469 11115 9503
rect 11057 9463 11115 9469
rect 6362 9432 6368 9444
rect 5276 9404 6368 9432
rect 2682 9364 2688 9376
rect 1780 9336 2688 9364
rect 2682 9324 2688 9336
rect 2740 9364 2746 9376
rect 3436 9364 3464 9404
rect 6362 9392 6368 9404
rect 6420 9392 6426 9444
rect 6546 9392 6552 9444
rect 6604 9392 6610 9444
rect 8294 9432 8300 9444
rect 6840 9404 8300 9432
rect 2740 9336 3464 9364
rect 2740 9324 2746 9336
rect 3510 9324 3516 9376
rect 3568 9324 3574 9376
rect 6380 9364 6408 9392
rect 6840 9364 6868 9404
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 10042 9392 10048 9444
rect 10100 9432 10106 9444
rect 10505 9435 10563 9441
rect 10505 9432 10517 9435
rect 10100 9404 10517 9432
rect 10100 9392 10106 9404
rect 10505 9401 10517 9404
rect 10551 9401 10563 9435
rect 10505 9395 10563 9401
rect 6380 9336 6868 9364
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7009 9367 7067 9373
rect 7009 9364 7021 9367
rect 6972 9336 7021 9364
rect 6972 9324 6978 9336
rect 7009 9333 7021 9336
rect 7055 9364 7067 9367
rect 7558 9364 7564 9376
rect 7055 9336 7564 9364
rect 7055 9333 7067 9336
rect 7009 9327 7067 9333
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 10226 9324 10232 9376
rect 10284 9364 10290 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 10284 9336 10425 9364
rect 10284 9324 10290 9336
rect 10413 9333 10425 9336
rect 10459 9364 10471 9367
rect 11072 9364 11100 9463
rect 12802 9460 12808 9512
rect 12860 9500 12866 9512
rect 12989 9503 13047 9509
rect 12989 9500 13001 9503
rect 12860 9472 13001 9500
rect 12860 9460 12866 9472
rect 12989 9469 13001 9472
rect 13035 9469 13047 9503
rect 12989 9463 13047 9469
rect 13096 9432 13124 9540
rect 13173 9537 13185 9571
rect 13219 9537 13231 9571
rect 13173 9531 13231 9537
rect 13188 9500 13216 9531
rect 13354 9528 13360 9580
rect 13412 9568 13418 9580
rect 14093 9571 14151 9577
rect 14093 9568 14105 9571
rect 13412 9540 14105 9568
rect 13412 9528 13418 9540
rect 14093 9537 14105 9540
rect 14139 9537 14151 9571
rect 14093 9531 14151 9537
rect 13449 9503 13507 9509
rect 13449 9500 13461 9503
rect 13188 9472 13461 9500
rect 13449 9469 13461 9472
rect 13495 9469 13507 9503
rect 13449 9463 13507 9469
rect 13538 9460 13544 9512
rect 13596 9460 13602 9512
rect 13630 9460 13636 9512
rect 13688 9460 13694 9512
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 13556 9432 13584 9460
rect 13740 9432 13768 9463
rect 13814 9460 13820 9512
rect 13872 9460 13878 9512
rect 13909 9503 13967 9509
rect 13909 9469 13921 9503
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 13096 9404 13768 9432
rect 10459 9336 11100 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 11790 9324 11796 9376
rect 11848 9364 11854 9376
rect 12250 9364 12256 9376
rect 11848 9336 12256 9364
rect 11848 9324 11854 9336
rect 12250 9324 12256 9336
rect 12308 9364 12314 9376
rect 12802 9364 12808 9376
rect 12308 9336 12808 9364
rect 12308 9324 12314 9336
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 13357 9367 13415 9373
rect 13357 9333 13369 9367
rect 13403 9364 13415 9367
rect 13722 9364 13728 9376
rect 13403 9336 13728 9364
rect 13403 9333 13415 9336
rect 13357 9327 13415 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 13924 9364 13952 9463
rect 14366 9460 14372 9512
rect 14424 9460 14430 9512
rect 14550 9364 14556 9376
rect 13924 9336 14556 9364
rect 14550 9324 14556 9336
rect 14608 9364 14614 9376
rect 15841 9367 15899 9373
rect 15841 9364 15853 9367
rect 14608 9336 15853 9364
rect 14608 9324 14614 9336
rect 15841 9333 15853 9336
rect 15887 9364 15899 9367
rect 16114 9364 16120 9376
rect 15887 9336 16120 9364
rect 15887 9333 15899 9336
rect 15841 9327 15899 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 944 9274 16836 9296
rect 944 9222 950 9274
rect 1002 9222 1014 9274
rect 1066 9222 1078 9274
rect 1130 9222 1142 9274
rect 1194 9222 1206 9274
rect 1258 9222 4950 9274
rect 5002 9222 5014 9274
rect 5066 9222 5078 9274
rect 5130 9222 5142 9274
rect 5194 9222 5206 9274
rect 5258 9222 8950 9274
rect 9002 9222 9014 9274
rect 9066 9222 9078 9274
rect 9130 9222 9142 9274
rect 9194 9222 9206 9274
rect 9258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 16836 9274
rect 944 9200 16836 9222
rect 2038 9120 2044 9172
rect 2096 9160 2102 9172
rect 2225 9163 2283 9169
rect 2225 9160 2237 9163
rect 2096 9132 2237 9160
rect 2096 9120 2102 9132
rect 2225 9129 2237 9132
rect 2271 9129 2283 9163
rect 2225 9123 2283 9129
rect 5261 9163 5319 9169
rect 5261 9129 5273 9163
rect 5307 9160 5319 9163
rect 6641 9163 6699 9169
rect 5307 9132 6316 9160
rect 5307 9129 5319 9132
rect 5261 9123 5319 9129
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 3878 9024 3884 9036
rect 3568 8996 3884 9024
rect 3568 8984 3574 8996
rect 3878 8984 3884 8996
rect 3936 9024 3942 9036
rect 4341 9027 4399 9033
rect 4341 9024 4353 9027
rect 3936 8996 4353 9024
rect 3936 8984 3942 8996
rect 4341 8993 4353 8996
rect 4387 8993 4399 9027
rect 4341 8987 4399 8993
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 1946 8956 1952 8968
rect 1811 8928 1952 8956
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 1946 8916 1952 8928
rect 2004 8916 2010 8968
rect 2409 8959 2467 8965
rect 2409 8925 2421 8959
rect 2455 8956 2467 8959
rect 2455 8928 2774 8956
rect 2455 8925 2467 8928
rect 2409 8919 2467 8925
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1397 8891 1455 8897
rect 1397 8888 1409 8891
rect 992 8860 1409 8888
rect 992 8848 998 8860
rect 1397 8857 1409 8860
rect 1443 8857 1455 8891
rect 1397 8851 1455 8857
rect 2746 8820 2774 8928
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4672 8928 4997 8956
rect 4672 8916 4678 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5276 8956 5304 9123
rect 5442 9052 5448 9104
rect 5500 9052 5506 9104
rect 5994 9092 6000 9104
rect 5736 9064 6000 9092
rect 5736 9033 5764 9064
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 6181 9095 6239 9101
rect 6181 9061 6193 9095
rect 6227 9061 6239 9095
rect 6288 9092 6316 9132
rect 6641 9129 6653 9163
rect 6687 9160 6699 9163
rect 7650 9160 7656 9172
rect 6687 9132 7656 9160
rect 6687 9129 6699 9132
rect 6641 9123 6699 9129
rect 7650 9120 7656 9132
rect 7708 9120 7714 9172
rect 9309 9163 9367 9169
rect 9309 9129 9321 9163
rect 9355 9160 9367 9163
rect 9490 9160 9496 9172
rect 9355 9132 9496 9160
rect 9355 9129 9367 9132
rect 9309 9123 9367 9129
rect 9490 9120 9496 9132
rect 9548 9160 9554 9172
rect 12529 9163 12587 9169
rect 9548 9132 12434 9160
rect 9548 9120 9554 9132
rect 6288 9064 6684 9092
rect 6181 9055 6239 9061
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 8993 5779 9027
rect 6196 9024 6224 9055
rect 6196 8996 6500 9024
rect 5721 8987 5779 8993
rect 5215 8928 5304 8956
rect 5997 8959 6055 8965
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5997 8925 6009 8959
rect 6043 8956 6055 8959
rect 6043 8928 6316 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 4157 8891 4215 8897
rect 4157 8857 4169 8891
rect 4203 8888 4215 8891
rect 5077 8891 5135 8897
rect 5077 8888 5089 8891
rect 4203 8860 5089 8888
rect 4203 8857 4215 8860
rect 4157 8851 4215 8857
rect 5077 8857 5089 8860
rect 5123 8857 5135 8891
rect 5077 8851 5135 8857
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 2746 8792 3801 8820
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 4249 8823 4307 8829
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 4430 8820 4436 8832
rect 4295 8792 4436 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 6288 8829 6316 8928
rect 6362 8916 6368 8968
rect 6420 8916 6426 8968
rect 6273 8823 6331 8829
rect 6273 8789 6285 8823
rect 6319 8789 6331 8823
rect 6380 8820 6408 8916
rect 6472 8888 6500 8996
rect 6546 8984 6552 9036
rect 6604 8984 6610 9036
rect 6656 8965 6684 9064
rect 9214 9052 9220 9104
rect 9272 9052 9278 9104
rect 12250 9052 12256 9104
rect 12308 9052 12314 9104
rect 6733 9027 6791 9033
rect 6733 8993 6745 9027
rect 6779 9024 6791 9027
rect 7006 9024 7012 9036
rect 6779 8996 7012 9024
rect 6779 8993 6791 8996
rect 6733 8987 6791 8993
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7466 8984 7472 9036
rect 7524 9024 7530 9036
rect 8754 9024 8760 9036
rect 7524 8996 8760 9024
rect 7524 8984 7530 8996
rect 8754 8984 8760 8996
rect 8812 9024 8818 9036
rect 10042 9024 10048 9036
rect 8812 8996 9076 9024
rect 8812 8984 8818 8996
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 9048 8965 9076 8996
rect 9232 8996 10048 9024
rect 9232 8965 9260 8996
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 10134 8984 10140 9036
rect 10192 9024 10198 9036
rect 11514 9024 11520 9036
rect 10192 8996 11520 9024
rect 10192 8984 10198 8996
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 12161 9027 12219 9033
rect 11664 8996 11928 9024
rect 11664 8984 11670 8996
rect 11900 8968 11928 8996
rect 12161 8993 12173 9027
rect 12207 9024 12219 9027
rect 12268 9024 12296 9052
rect 12207 8996 12296 9024
rect 12207 8993 12219 8996
rect 12161 8987 12219 8993
rect 9033 8959 9091 8965
rect 9033 8925 9045 8959
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 9766 8956 9772 8968
rect 9456 8928 9772 8956
rect 9456 8916 9462 8928
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8956 11115 8959
rect 11330 8956 11336 8968
rect 11103 8928 11336 8956
rect 11103 8925 11115 8928
rect 11057 8919 11115 8925
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 11698 8916 11704 8968
rect 11756 8916 11762 8968
rect 11882 8916 11888 8968
rect 11940 8916 11946 8968
rect 12406 8956 12434 9132
rect 12529 9129 12541 9163
rect 12575 9160 12587 9163
rect 12618 9160 12624 9172
rect 12575 9132 12624 9160
rect 12575 9129 12587 9132
rect 12529 9123 12587 9129
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 12989 9163 13047 9169
rect 12989 9129 13001 9163
rect 13035 9160 13047 9163
rect 13998 9160 14004 9172
rect 13035 9132 14004 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14277 9163 14335 9169
rect 14277 9129 14289 9163
rect 14323 9160 14335 9163
rect 14366 9160 14372 9172
rect 14323 9132 14372 9160
rect 14323 9129 14335 9132
rect 14277 9123 14335 9129
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 12805 9095 12863 9101
rect 12805 9092 12817 9095
rect 12544 9064 12817 9092
rect 12544 9036 12572 9064
rect 12805 9061 12817 9064
rect 12851 9061 12863 9095
rect 12805 9055 12863 9061
rect 12526 8984 12532 9036
rect 12584 8984 12590 9036
rect 15562 9024 15568 9036
rect 12912 8996 15568 9024
rect 12912 8956 12940 8996
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 12406 8928 12940 8956
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13780 8928 14105 8956
rect 13780 8916 13786 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 16114 8916 16120 8968
rect 16172 8916 16178 8968
rect 7009 8891 7067 8897
rect 7009 8888 7021 8891
rect 6472 8860 7021 8888
rect 7009 8857 7021 8860
rect 7055 8857 7067 8891
rect 8757 8891 8815 8897
rect 7009 8851 7067 8857
rect 7116 8860 7498 8888
rect 7116 8820 7144 8860
rect 8757 8857 8769 8891
rect 8803 8888 8815 8891
rect 10781 8891 10839 8897
rect 8803 8860 9168 8888
rect 8803 8857 8815 8860
rect 8757 8851 8815 8857
rect 6380 8792 7144 8820
rect 6273 8783 6331 8789
rect 7282 8780 7288 8832
rect 7340 8820 7346 8832
rect 8772 8820 8800 8851
rect 7340 8792 8800 8820
rect 9140 8820 9168 8860
rect 10781 8857 10793 8891
rect 10827 8888 10839 8891
rect 10870 8888 10876 8900
rect 10827 8860 10876 8888
rect 10827 8857 10839 8860
rect 10781 8851 10839 8857
rect 10870 8848 10876 8860
rect 10928 8848 10934 8900
rect 11241 8891 11299 8897
rect 11241 8857 11253 8891
rect 11287 8888 11299 8891
rect 11422 8888 11428 8900
rect 11287 8860 11428 8888
rect 11287 8857 11299 8860
rect 11241 8851 11299 8857
rect 11422 8848 11428 8860
rect 11480 8848 11486 8900
rect 11900 8888 11928 8916
rect 12713 8891 12771 8897
rect 12713 8888 12725 8891
rect 11900 8860 12725 8888
rect 12713 8857 12725 8860
rect 12759 8888 12771 8891
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 12759 8860 13185 8888
rect 12759 8857 12771 8860
rect 12713 8851 12771 8857
rect 13173 8857 13185 8860
rect 13219 8857 13231 8891
rect 13173 8851 13231 8857
rect 16485 8891 16543 8897
rect 16485 8857 16497 8891
rect 16531 8888 16543 8891
rect 16758 8888 16764 8900
rect 16531 8860 16764 8888
rect 16531 8857 16543 8860
rect 16485 8851 16543 8857
rect 16758 8848 16764 8860
rect 16816 8848 16822 8900
rect 10134 8820 10140 8832
rect 9140 8792 10140 8820
rect 7340 8780 7346 8792
rect 10134 8780 10140 8792
rect 10192 8780 10198 8832
rect 11514 8780 11520 8832
rect 11572 8820 11578 8832
rect 12526 8829 12532 8832
rect 12345 8823 12403 8829
rect 12345 8820 12357 8823
rect 11572 8792 12357 8820
rect 11572 8780 11578 8792
rect 12345 8789 12357 8792
rect 12391 8789 12403 8823
rect 12345 8783 12403 8789
rect 12513 8823 12532 8829
rect 12513 8789 12525 8823
rect 12584 8820 12590 8832
rect 12963 8823 13021 8829
rect 12963 8820 12975 8823
rect 12584 8792 12975 8820
rect 12513 8783 12532 8789
rect 12526 8780 12532 8783
rect 12584 8780 12590 8792
rect 12963 8789 12975 8792
rect 13009 8789 13021 8823
rect 12963 8783 13021 8789
rect 1104 8730 16836 8752
rect 1104 8678 1610 8730
rect 1662 8678 1674 8730
rect 1726 8678 1738 8730
rect 1790 8678 1802 8730
rect 1854 8678 1866 8730
rect 1918 8678 5610 8730
rect 5662 8678 5674 8730
rect 5726 8678 5738 8730
rect 5790 8678 5802 8730
rect 5854 8678 5866 8730
rect 5918 8678 9610 8730
rect 9662 8678 9674 8730
rect 9726 8678 9738 8730
rect 9790 8678 9802 8730
rect 9854 8678 9866 8730
rect 9918 8678 13610 8730
rect 13662 8678 13674 8730
rect 13726 8678 13738 8730
rect 13790 8678 13802 8730
rect 13854 8678 13866 8730
rect 13918 8678 16836 8730
rect 1104 8656 16836 8678
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 3936 8588 5212 8616
rect 3936 8576 3942 8588
rect 4154 8508 4160 8560
rect 4212 8548 4218 8560
rect 5077 8551 5135 8557
rect 5077 8548 5089 8551
rect 4212 8520 5089 8548
rect 4212 8508 4218 8520
rect 5077 8517 5089 8520
rect 5123 8517 5135 8551
rect 5077 8511 5135 8517
rect 2682 8440 2688 8492
rect 2740 8480 2746 8492
rect 2777 8483 2835 8489
rect 2777 8480 2789 8483
rect 2740 8452 2789 8480
rect 2740 8440 2746 8452
rect 2777 8449 2789 8452
rect 2823 8449 2835 8483
rect 2777 8443 2835 8449
rect 4522 8440 4528 8492
rect 4580 8440 4586 8492
rect 4798 8440 4804 8492
rect 4856 8480 4862 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4856 8452 4905 8480
rect 4856 8440 4862 8452
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8480 5043 8483
rect 5184 8480 5212 8588
rect 5994 8576 6000 8628
rect 6052 8576 6058 8628
rect 8938 8616 8944 8628
rect 8772 8588 8944 8616
rect 5261 8551 5319 8557
rect 5261 8517 5273 8551
rect 5307 8548 5319 8551
rect 5350 8548 5356 8560
rect 5307 8520 5356 8548
rect 5307 8517 5319 8520
rect 5261 8511 5319 8517
rect 5350 8508 5356 8520
rect 5408 8548 5414 8560
rect 5534 8548 5540 8560
rect 5408 8520 5540 8548
rect 5408 8508 5414 8520
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 5031 8452 5212 8480
rect 6012 8480 6040 8576
rect 8772 8548 8800 8588
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9214 8576 9220 8628
rect 9272 8576 9278 8628
rect 11330 8576 11336 8628
rect 11388 8616 11394 8628
rect 13354 8616 13360 8628
rect 11388 8588 13360 8616
rect 11388 8576 11394 8588
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14642 8616 14648 8628
rect 14056 8588 14648 8616
rect 14056 8576 14062 8588
rect 14642 8576 14648 8588
rect 14700 8616 14706 8628
rect 15105 8619 15163 8625
rect 15105 8616 15117 8619
rect 14700 8588 15117 8616
rect 14700 8576 14706 8588
rect 15105 8585 15117 8588
rect 15151 8585 15163 8619
rect 15105 8579 15163 8585
rect 9232 8548 9260 8576
rect 10134 8548 10140 8560
rect 8496 8520 8800 8548
rect 8864 8520 9260 8548
rect 9324 8520 10140 8548
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6012 8452 6377 8480
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 8496 8489 8524 8520
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8449 8631 8483
rect 8573 8443 8631 8449
rect 2314 8372 2320 8424
rect 2372 8412 2378 8424
rect 6638 8412 6644 8424
rect 2372 8384 6644 8412
rect 2372 8372 2378 8384
rect 6638 8372 6644 8384
rect 6696 8372 6702 8424
rect 8588 8344 8616 8443
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 8864 8489 8892 8520
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 8938 8440 8944 8492
rect 8996 8440 9002 8492
rect 9122 8440 9128 8492
rect 9180 8440 9186 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8480 9275 8483
rect 9324 8480 9352 8520
rect 10134 8508 10140 8520
rect 10192 8508 10198 8560
rect 11422 8508 11428 8560
rect 11480 8548 11486 8560
rect 11480 8520 14122 8548
rect 11480 8508 11486 8520
rect 9263 8452 9352 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 9398 8440 9404 8492
rect 9456 8440 9462 8492
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8480 9643 8483
rect 9631 8452 9665 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8412 8723 8415
rect 8772 8412 8800 8440
rect 8956 8412 8984 8440
rect 8711 8384 8800 8412
rect 8864 8384 8984 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 8864 8353 8892 8384
rect 9030 8372 9036 8424
rect 9088 8412 9094 8424
rect 9600 8412 9628 8443
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11020 8452 11529 8480
rect 11020 8440 11026 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13354 8480 13360 8492
rect 13219 8452 13360 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 15120 8480 15148 8579
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 15841 8619 15899 8625
rect 15841 8616 15853 8619
rect 15804 8588 15853 8616
rect 15804 8576 15810 8588
rect 15841 8585 15853 8588
rect 15887 8585 15899 8619
rect 15841 8579 15899 8585
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 15120 8452 15485 8480
rect 15473 8449 15485 8452
rect 15519 8480 15531 8483
rect 16025 8483 16083 8489
rect 16025 8480 16037 8483
rect 15519 8452 16037 8480
rect 15519 8449 15531 8452
rect 15473 8443 15531 8449
rect 16025 8449 16037 8452
rect 16071 8449 16083 8483
rect 16025 8443 16083 8449
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 16209 8483 16267 8489
rect 16209 8480 16221 8483
rect 16172 8452 16221 8480
rect 16172 8440 16178 8452
rect 16209 8449 16221 8452
rect 16255 8449 16267 8483
rect 16209 8443 16267 8449
rect 10410 8412 10416 8424
rect 9088 8384 10416 8412
rect 9088 8372 9094 8384
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 13630 8372 13636 8424
rect 13688 8372 13694 8424
rect 13722 8372 13728 8424
rect 13780 8412 13786 8424
rect 15381 8415 15439 8421
rect 15381 8412 15393 8415
rect 13780 8384 15393 8412
rect 13780 8372 13786 8384
rect 15381 8381 15393 8384
rect 15427 8381 15439 8415
rect 15381 8375 15439 8381
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8381 15623 8415
rect 15565 8375 15623 8381
rect 15657 8415 15715 8421
rect 15657 8381 15669 8415
rect 15703 8412 15715 8415
rect 16132 8412 16160 8440
rect 15703 8384 16160 8412
rect 15703 8381 15715 8384
rect 15657 8375 15715 8381
rect 8849 8347 8907 8353
rect 8588 8316 8800 8344
rect 4246 8236 4252 8288
rect 4304 8276 4310 8288
rect 4709 8279 4767 8285
rect 4709 8276 4721 8279
rect 4304 8248 4721 8276
rect 4304 8236 4310 8248
rect 4709 8245 4721 8248
rect 4755 8245 4767 8279
rect 4709 8239 4767 8245
rect 5261 8279 5319 8285
rect 5261 8245 5273 8279
rect 5307 8276 5319 8279
rect 5350 8276 5356 8288
rect 5307 8248 5356 8276
rect 5307 8245 5319 8248
rect 5261 8239 5319 8245
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 6825 8279 6883 8285
rect 6825 8245 6837 8279
rect 6871 8276 6883 8279
rect 8662 8276 8668 8288
rect 6871 8248 8668 8276
rect 6871 8245 6883 8248
rect 6825 8239 6883 8245
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 8772 8276 8800 8316
rect 8849 8313 8861 8347
rect 8895 8313 8907 8347
rect 8849 8307 8907 8313
rect 9306 8304 9312 8356
rect 9364 8304 9370 8356
rect 10870 8344 10876 8356
rect 9416 8316 10876 8344
rect 9416 8276 9444 8316
rect 10870 8304 10876 8316
rect 10928 8304 10934 8356
rect 15580 8344 15608 8375
rect 14660 8316 15608 8344
rect 8772 8248 9444 8276
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11698 8276 11704 8288
rect 11112 8248 11704 8276
rect 11112 8236 11118 8248
rect 11698 8236 11704 8248
rect 11756 8236 11762 8288
rect 14182 8236 14188 8288
rect 14240 8276 14246 8288
rect 14660 8276 14688 8316
rect 14240 8248 14688 8276
rect 14240 8236 14246 8248
rect 15194 8236 15200 8288
rect 15252 8236 15258 8288
rect 944 8186 16836 8208
rect 944 8134 950 8186
rect 1002 8134 1014 8186
rect 1066 8134 1078 8186
rect 1130 8134 1142 8186
rect 1194 8134 1206 8186
rect 1258 8134 4950 8186
rect 5002 8134 5014 8186
rect 5066 8134 5078 8186
rect 5130 8134 5142 8186
rect 5194 8134 5206 8186
rect 5258 8134 8950 8186
rect 9002 8134 9014 8186
rect 9066 8134 9078 8186
rect 9130 8134 9142 8186
rect 9194 8134 9206 8186
rect 9258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 16836 8186
rect 944 8112 16836 8134
rect 3145 8075 3203 8081
rect 3145 8041 3157 8075
rect 3191 8072 3203 8075
rect 4154 8072 4160 8084
rect 3191 8044 4160 8072
rect 3191 8041 3203 8044
rect 3145 8035 3203 8041
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 4798 8032 4804 8084
rect 4856 8072 4862 8084
rect 4893 8075 4951 8081
rect 4893 8072 4905 8075
rect 4856 8044 4905 8072
rect 4856 8032 4862 8044
rect 4893 8041 4905 8044
rect 4939 8041 4951 8075
rect 4893 8035 4951 8041
rect 5350 8032 5356 8084
rect 5408 8032 5414 8084
rect 6638 8032 6644 8084
rect 6696 8072 6702 8084
rect 11422 8072 11428 8084
rect 6696 8044 11428 8072
rect 6696 8032 6702 8044
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 12069 8075 12127 8081
rect 12069 8041 12081 8075
rect 12115 8072 12127 8075
rect 12115 8044 12149 8072
rect 12115 8041 12127 8044
rect 12069 8035 12127 8041
rect 4709 8007 4767 8013
rect 4709 7973 4721 8007
rect 4755 8004 4767 8007
rect 5368 8004 5396 8032
rect 4755 7976 5396 8004
rect 10873 8007 10931 8013
rect 4755 7973 4767 7976
rect 4709 7967 4767 7973
rect 10873 7973 10885 8007
rect 10919 8004 10931 8007
rect 11054 8004 11060 8016
rect 10919 7976 11060 8004
rect 10919 7973 10931 7976
rect 10873 7967 10931 7973
rect 11054 7964 11060 7976
rect 11112 7964 11118 8016
rect 11348 7976 11652 8004
rect 1394 7896 1400 7948
rect 1452 7896 1458 7948
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 1719 7908 4353 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 4341 7899 4399 7905
rect 4430 7896 4436 7948
rect 4488 7936 4494 7948
rect 4801 7939 4859 7945
rect 4801 7936 4813 7939
rect 4488 7908 4813 7936
rect 4488 7896 4494 7908
rect 4801 7905 4813 7908
rect 4847 7905 4859 7939
rect 4801 7899 4859 7905
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 5537 7939 5595 7945
rect 5537 7936 5549 7939
rect 5500 7908 5549 7936
rect 5500 7896 5506 7908
rect 5537 7905 5549 7908
rect 5583 7936 5595 7939
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 5583 7908 5733 7936
rect 5583 7905 5595 7908
rect 5537 7899 5595 7905
rect 5721 7905 5733 7908
rect 5767 7936 5779 7939
rect 7282 7936 7288 7948
rect 5767 7908 7288 7936
rect 5767 7905 5779 7908
rect 5721 7899 5779 7905
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 7374 7896 7380 7948
rect 7432 7936 7438 7948
rect 7837 7939 7895 7945
rect 7837 7936 7849 7939
rect 7432 7908 7849 7936
rect 7432 7896 7438 7908
rect 7837 7905 7849 7908
rect 7883 7905 7895 7939
rect 7837 7899 7895 7905
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 3804 7800 3832 7831
rect 3878 7828 3884 7880
rect 3936 7828 3942 7880
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7868 4123 7871
rect 4154 7868 4160 7880
rect 4111 7840 4160 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 4295 7840 4537 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4525 7837 4537 7840
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 5994 7868 6000 7880
rect 5951 7840 6000 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 5353 7803 5411 7809
rect 2056 7772 2162 7800
rect 3804 7772 4292 7800
rect 2056 7744 2084 7772
rect 4264 7744 4292 7772
rect 5353 7769 5365 7803
rect 5399 7800 5411 7803
rect 5920 7800 5948 7831
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 6181 7871 6239 7877
rect 6181 7868 6193 7871
rect 6135 7840 6193 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 6181 7837 6193 7840
rect 6227 7837 6239 7871
rect 6181 7831 6239 7837
rect 7558 7828 7564 7880
rect 7616 7828 7622 7880
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7868 9919 7871
rect 9950 7868 9956 7880
rect 9907 7840 9956 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 10042 7828 10048 7880
rect 10100 7828 10106 7880
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 10192 7840 10333 7868
rect 10192 7828 10198 7840
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 10410 7828 10416 7880
rect 10468 7868 10474 7880
rect 10873 7871 10931 7877
rect 10873 7868 10885 7871
rect 10468 7840 10885 7868
rect 10468 7828 10474 7840
rect 10873 7837 10885 7840
rect 10919 7868 10931 7871
rect 11072 7868 11100 7964
rect 11348 7877 11376 7976
rect 11624 7936 11652 7976
rect 11974 7964 11980 8016
rect 12032 8004 12038 8016
rect 12084 8004 12112 8035
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 13446 8072 13452 8084
rect 12584 8044 13452 8072
rect 12584 8032 12590 8044
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 13630 8032 13636 8084
rect 13688 8072 13694 8084
rect 13725 8075 13783 8081
rect 13725 8072 13737 8075
rect 13688 8044 13737 8072
rect 13688 8032 13694 8044
rect 13725 8041 13737 8044
rect 13771 8041 13783 8075
rect 13725 8035 13783 8041
rect 15194 8032 15200 8084
rect 15252 8032 15258 8084
rect 12032 7976 12940 8004
rect 12032 7964 12038 7976
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 11624 7908 12357 7936
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 12434 7896 12440 7948
rect 12492 7896 12498 7948
rect 12912 7945 12940 7976
rect 13372 7976 14872 8004
rect 12897 7939 12955 7945
rect 12897 7905 12909 7939
rect 12943 7905 12955 7939
rect 12897 7899 12955 7905
rect 11514 7877 11520 7880
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 10919 7840 11008 7868
rect 11072 7840 11253 7868
rect 10919 7837 10931 7840
rect 10873 7831 10931 7837
rect 5399 7772 5948 7800
rect 5399 7769 5411 7772
rect 5353 7763 5411 7769
rect 2038 7692 2044 7744
rect 2096 7692 2102 7744
rect 4246 7692 4252 7744
rect 4304 7732 4310 7744
rect 4890 7732 4896 7744
rect 4304 7704 4896 7732
rect 4304 7692 4310 7704
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5261 7735 5319 7741
rect 5261 7701 5273 7735
rect 5307 7732 5319 7735
rect 6086 7732 6092 7744
rect 5307 7704 6092 7732
rect 5307 7701 5319 7704
rect 5261 7695 5319 7701
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6362 7692 6368 7744
rect 6420 7692 6426 7744
rect 9217 7735 9275 7741
rect 9217 7701 9229 7735
rect 9263 7732 9275 7735
rect 9306 7732 9312 7744
rect 9263 7704 9312 7732
rect 9263 7701 9275 7704
rect 9217 7695 9275 7701
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 10980 7732 11008 7840
rect 11241 7837 11253 7840
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11497 7871 11520 7877
rect 11497 7837 11509 7871
rect 11497 7831 11520 7837
rect 11514 7828 11520 7831
rect 11572 7828 11578 7880
rect 12452 7868 12480 7896
rect 13372 7880 13400 7976
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7936 13507 7939
rect 14093 7939 14151 7945
rect 14093 7936 14105 7939
rect 13495 7908 14105 7936
rect 13495 7905 13507 7908
rect 13449 7899 13507 7905
rect 14093 7905 14105 7908
rect 14139 7905 14151 7939
rect 14093 7899 14151 7905
rect 14642 7896 14648 7948
rect 14700 7896 14706 7948
rect 14844 7945 14872 7976
rect 14829 7939 14887 7945
rect 14829 7905 14841 7939
rect 14875 7905 14887 7939
rect 15212 7936 15240 8032
rect 14829 7899 14887 7905
rect 15028 7908 15240 7936
rect 11624 7840 12480 7868
rect 11624 7732 11652 7840
rect 11882 7760 11888 7812
rect 11940 7760 11946 7812
rect 12100 7809 12128 7840
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 15028 7877 15056 7908
rect 13541 7871 13599 7877
rect 13541 7837 13553 7871
rect 13587 7868 13599 7871
rect 15013 7871 15071 7877
rect 13587 7840 14136 7868
rect 13587 7837 13599 7840
rect 13541 7831 13599 7837
rect 12090 7803 12148 7809
rect 12090 7769 12102 7803
rect 12136 7769 12148 7803
rect 13556 7800 13584 7831
rect 12090 7763 12148 7769
rect 12176 7772 13584 7800
rect 10980 7704 11652 7732
rect 11698 7692 11704 7744
rect 11756 7692 11762 7744
rect 11790 7692 11796 7744
rect 11848 7732 11854 7744
rect 12176 7732 12204 7772
rect 14108 7744 14136 7840
rect 15013 7837 15025 7871
rect 15059 7837 15071 7871
rect 15013 7831 15071 7837
rect 15197 7871 15255 7877
rect 15197 7837 15209 7871
rect 15243 7868 15255 7871
rect 15473 7871 15531 7877
rect 15473 7868 15485 7871
rect 15243 7840 15485 7868
rect 15243 7837 15255 7840
rect 15197 7831 15255 7837
rect 15473 7837 15485 7840
rect 15519 7837 15531 7871
rect 15473 7831 15531 7837
rect 15562 7828 15568 7880
rect 15620 7868 15626 7880
rect 16117 7871 16175 7877
rect 16117 7868 16129 7871
rect 15620 7840 16129 7868
rect 15620 7828 15626 7840
rect 16117 7837 16129 7840
rect 16163 7837 16175 7871
rect 16117 7831 16175 7837
rect 11848 7704 12204 7732
rect 12253 7735 12311 7741
rect 11848 7692 11854 7704
rect 12253 7701 12265 7735
rect 12299 7732 12311 7735
rect 12618 7732 12624 7744
rect 12299 7704 12624 7732
rect 12299 7701 12311 7704
rect 12253 7695 12311 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 13081 7735 13139 7741
rect 13081 7732 13093 7735
rect 12860 7704 13093 7732
rect 12860 7692 12866 7704
rect 13081 7701 13093 7704
rect 13127 7732 13139 7735
rect 13354 7732 13360 7744
rect 13127 7704 13360 7732
rect 13127 7701 13139 7704
rect 13081 7695 13139 7701
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 14090 7692 14096 7744
rect 14148 7692 14154 7744
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 15289 7735 15347 7741
rect 15289 7732 15301 7735
rect 14884 7704 15301 7732
rect 14884 7692 14890 7704
rect 15289 7701 15301 7704
rect 15335 7701 15347 7735
rect 15289 7695 15347 7701
rect 16393 7735 16451 7741
rect 16393 7701 16405 7735
rect 16439 7732 16451 7735
rect 16758 7732 16764 7744
rect 16439 7704 16764 7732
rect 16439 7701 16451 7704
rect 16393 7695 16451 7701
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 1104 7642 16836 7664
rect 1104 7590 1610 7642
rect 1662 7590 1674 7642
rect 1726 7590 1738 7642
rect 1790 7590 1802 7642
rect 1854 7590 1866 7642
rect 1918 7590 5610 7642
rect 5662 7590 5674 7642
rect 5726 7590 5738 7642
rect 5790 7590 5802 7642
rect 5854 7590 5866 7642
rect 5918 7590 9610 7642
rect 9662 7590 9674 7642
rect 9726 7590 9738 7642
rect 9790 7590 9802 7642
rect 9854 7590 9866 7642
rect 9918 7590 13610 7642
rect 13662 7590 13674 7642
rect 13726 7590 13738 7642
rect 13790 7590 13802 7642
rect 13854 7590 13866 7642
rect 13918 7590 16836 7642
rect 1104 7568 16836 7590
rect 2038 7488 2044 7540
rect 2096 7488 2102 7540
rect 3973 7531 4031 7537
rect 3973 7497 3985 7531
rect 4019 7528 4031 7531
rect 4154 7528 4160 7540
rect 4019 7500 4160 7528
rect 4019 7497 4031 7500
rect 3973 7491 4031 7497
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4246 7488 4252 7540
rect 4304 7488 4310 7540
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7497 4491 7531
rect 4433 7491 4491 7497
rect 2133 7463 2191 7469
rect 2133 7429 2145 7463
rect 2179 7460 2191 7463
rect 2314 7460 2320 7472
rect 2179 7432 2320 7460
rect 2179 7429 2191 7432
rect 2133 7423 2191 7429
rect 2314 7420 2320 7432
rect 2372 7420 2378 7472
rect 3878 7469 3884 7472
rect 3856 7463 3884 7469
rect 3856 7460 3868 7463
rect 2424 7432 3868 7460
rect 2424 7324 2452 7432
rect 3856 7429 3868 7432
rect 3856 7423 3884 7429
rect 3878 7420 3884 7423
rect 3936 7420 3942 7472
rect 4065 7463 4123 7469
rect 4065 7429 4077 7463
rect 4111 7460 4123 7463
rect 4264 7460 4292 7488
rect 4111 7432 4292 7460
rect 4111 7429 4123 7432
rect 4065 7423 4123 7429
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 3142 7392 3148 7404
rect 2547 7364 3148 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 3142 7352 3148 7364
rect 3200 7392 3206 7404
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 3200 7364 3525 7392
rect 3200 7352 3206 7364
rect 3513 7361 3525 7364
rect 3559 7361 3571 7395
rect 3513 7355 3571 7361
rect 4448 7336 4476 7491
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 7616 7500 7665 7528
rect 7616 7488 7622 7500
rect 7653 7497 7665 7500
rect 7699 7497 7711 7531
rect 7653 7491 7711 7497
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 11756 7500 11836 7528
rect 11756 7488 11762 7500
rect 7469 7463 7527 7469
rect 7469 7460 7481 7463
rect 6104 7432 7481 7460
rect 6104 7404 6132 7432
rect 7469 7429 7481 7432
rect 7515 7460 7527 7463
rect 9214 7460 9220 7472
rect 7515 7432 9220 7460
rect 7515 7429 7527 7432
rect 7469 7423 7527 7429
rect 9214 7420 9220 7432
rect 9272 7420 9278 7472
rect 10686 7460 10692 7472
rect 10060 7432 10692 7460
rect 10060 7404 10088 7432
rect 10686 7420 10692 7432
rect 10744 7460 10750 7472
rect 11808 7469 11836 7500
rect 11974 7488 11980 7540
rect 12032 7528 12038 7540
rect 13265 7531 13323 7537
rect 13265 7528 13277 7531
rect 12032 7500 13277 7528
rect 12032 7488 12038 7500
rect 13265 7497 13277 7500
rect 13311 7497 13323 7531
rect 13265 7491 13323 7497
rect 11793 7463 11851 7469
rect 10744 7432 11100 7460
rect 10744 7420 10750 7432
rect 4890 7352 4896 7404
rect 4948 7352 4954 7404
rect 5350 7352 5356 7404
rect 5408 7392 5414 7404
rect 5408 7364 5488 7392
rect 5408 7352 5414 7364
rect 2593 7327 2651 7333
rect 2593 7324 2605 7327
rect 2424 7296 2605 7324
rect 2593 7293 2605 7296
rect 2639 7293 2651 7327
rect 2593 7287 2651 7293
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7293 2743 7327
rect 2685 7287 2743 7293
rect 2777 7327 2835 7333
rect 2777 7293 2789 7327
rect 2823 7324 2835 7327
rect 3970 7324 3976 7336
rect 2823 7296 3976 7324
rect 2823 7293 2835 7296
rect 2777 7287 2835 7293
rect 2700 7256 2728 7287
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4341 7327 4399 7333
rect 4341 7293 4353 7327
rect 4387 7293 4399 7327
rect 4341 7287 4399 7293
rect 4154 7256 4160 7268
rect 2700 7228 4160 7256
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 4356 7256 4384 7287
rect 4430 7284 4436 7336
rect 4488 7284 4494 7336
rect 5460 7324 5488 7364
rect 6086 7352 6092 7404
rect 6144 7352 6150 7404
rect 7282 7352 7288 7404
rect 7340 7352 7346 7404
rect 7558 7352 7564 7404
rect 7616 7392 7622 7404
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 7616 7364 7849 7392
rect 7616 7352 7622 7364
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 9490 7352 9496 7404
rect 9548 7392 9554 7404
rect 9585 7395 9643 7401
rect 9585 7392 9597 7395
rect 9548 7364 9597 7392
rect 9548 7352 9554 7364
rect 9585 7361 9597 7364
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7392 10011 7395
rect 10042 7392 10048 7404
rect 9999 7364 10048 7392
rect 9999 7361 10011 7364
rect 9953 7355 10011 7361
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 10134 7352 10140 7404
rect 10192 7352 10198 7404
rect 10410 7352 10416 7404
rect 10468 7352 10474 7404
rect 11072 7401 11100 7432
rect 11793 7429 11805 7463
rect 11839 7429 11851 7463
rect 13446 7460 13452 7472
rect 13018 7432 13452 7460
rect 11793 7423 11851 7429
rect 13446 7420 13452 7432
rect 13504 7460 13510 7472
rect 13504 7432 14858 7460
rect 13504 7420 13510 7432
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 5460 7296 10977 7324
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 10965 7287 11023 7293
rect 10980 7256 11008 7287
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 11204 7296 11529 7324
rect 11204 7284 11210 7296
rect 11517 7293 11529 7296
rect 11563 7293 11575 7327
rect 11882 7324 11888 7336
rect 11517 7287 11575 7293
rect 11624 7296 11888 7324
rect 4356 7228 4568 7256
rect 10980 7228 11100 7256
rect 2314 7148 2320 7200
rect 2372 7148 2378 7200
rect 2866 7148 2872 7200
rect 2924 7188 2930 7200
rect 2961 7191 3019 7197
rect 2961 7188 2973 7191
rect 2924 7160 2973 7188
rect 2924 7148 2930 7160
rect 2961 7157 2973 7160
rect 3007 7157 3019 7191
rect 2961 7151 3019 7157
rect 3326 7148 3332 7200
rect 3384 7188 3390 7200
rect 3697 7191 3755 7197
rect 3697 7188 3709 7191
rect 3384 7160 3709 7188
rect 3384 7148 3390 7160
rect 3697 7157 3709 7160
rect 3743 7157 3755 7191
rect 4540 7188 4568 7228
rect 4801 7191 4859 7197
rect 4801 7188 4813 7191
rect 4540 7160 4813 7188
rect 3697 7151 3755 7157
rect 4801 7157 4813 7160
rect 4847 7188 4859 7191
rect 5534 7188 5540 7200
rect 4847 7160 5540 7188
rect 4847 7157 4859 7160
rect 4801 7151 4859 7157
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 10962 7188 10968 7200
rect 7616 7160 10968 7188
rect 7616 7148 7622 7160
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 11072 7188 11100 7228
rect 11238 7216 11244 7268
rect 11296 7256 11302 7268
rect 11624 7256 11652 7296
rect 11882 7284 11888 7296
rect 11940 7284 11946 7336
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 13909 7327 13967 7333
rect 13909 7324 13921 7327
rect 12492 7296 13921 7324
rect 12492 7284 12498 7296
rect 13909 7293 13921 7296
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 13998 7284 14004 7336
rect 14056 7324 14062 7336
rect 14108 7324 14136 7355
rect 14056 7296 14136 7324
rect 14369 7327 14427 7333
rect 14056 7284 14062 7296
rect 14369 7293 14381 7327
rect 14415 7324 14427 7327
rect 14826 7324 14832 7336
rect 14415 7296 14832 7324
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 11296 7228 11652 7256
rect 11296 7216 11302 7228
rect 12526 7188 12532 7200
rect 11072 7160 12532 7188
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12802 7148 12808 7200
rect 12860 7188 12866 7200
rect 13357 7191 13415 7197
rect 13357 7188 13369 7191
rect 12860 7160 13369 7188
rect 12860 7148 12866 7160
rect 13357 7157 13369 7160
rect 13403 7157 13415 7191
rect 13357 7151 13415 7157
rect 15841 7191 15899 7197
rect 15841 7157 15853 7191
rect 15887 7188 15899 7191
rect 16114 7188 16120 7200
rect 15887 7160 16120 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 944 7098 16836 7120
rect 944 7046 950 7098
rect 1002 7046 1014 7098
rect 1066 7046 1078 7098
rect 1130 7046 1142 7098
rect 1194 7046 1206 7098
rect 1258 7046 4950 7098
rect 5002 7046 5014 7098
rect 5066 7046 5078 7098
rect 5130 7046 5142 7098
rect 5194 7046 5206 7098
rect 5258 7046 8950 7098
rect 9002 7046 9014 7098
rect 9066 7046 9078 7098
rect 9130 7046 9142 7098
rect 9194 7046 9206 7098
rect 9258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 16836 7098
rect 944 7024 16836 7046
rect 3142 6944 3148 6996
rect 3200 6944 3206 6996
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 5721 6987 5779 6993
rect 3936 6956 4292 6984
rect 3936 6944 3942 6956
rect 3160 6916 3188 6944
rect 3160 6888 4108 6916
rect 2406 6808 2412 6860
rect 2464 6848 2470 6860
rect 4080 6857 4108 6888
rect 4065 6851 4123 6857
rect 2464 6820 3464 6848
rect 2464 6808 2470 6820
rect 3436 6789 3464 6820
rect 4065 6817 4077 6851
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 4154 6808 4160 6860
rect 4212 6808 4218 6860
rect 4264 6857 4292 6956
rect 5721 6953 5733 6987
rect 5767 6984 5779 6987
rect 6270 6984 6276 6996
rect 5767 6956 6276 6984
rect 5767 6953 5779 6956
rect 5721 6947 5779 6953
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 6622 6987 6680 6993
rect 6622 6984 6634 6987
rect 6420 6956 6634 6984
rect 6420 6944 6426 6956
rect 6622 6953 6634 6956
rect 6668 6953 6680 6987
rect 6622 6947 6680 6953
rect 9204 6987 9262 6993
rect 9204 6953 9216 6987
rect 9250 6984 9262 6987
rect 9306 6984 9312 6996
rect 9250 6956 9312 6984
rect 9250 6953 9262 6956
rect 9204 6947 9262 6953
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 10686 6944 10692 6996
rect 10744 6944 10750 6996
rect 12434 6984 12440 6996
rect 12406 6944 12440 6984
rect 12492 6944 12498 6996
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 13538 6984 13544 6996
rect 12676 6956 13544 6984
rect 12676 6944 12682 6956
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 13651 6987 13709 6993
rect 13651 6953 13663 6987
rect 13697 6984 13709 6987
rect 14553 6987 14611 6993
rect 14553 6984 14565 6987
rect 13697 6956 14565 6984
rect 13697 6953 13709 6956
rect 13651 6947 13709 6953
rect 14553 6953 14565 6956
rect 14599 6953 14611 6987
rect 14553 6947 14611 6953
rect 8110 6876 8116 6928
rect 8168 6916 8174 6928
rect 8168 6888 8432 6916
rect 8168 6876 8174 6888
rect 4264 6851 4332 6857
rect 4264 6820 4286 6851
rect 4274 6817 4286 6820
rect 4320 6817 4332 6851
rect 4274 6811 4332 6817
rect 4614 6808 4620 6860
rect 4672 6848 4678 6860
rect 4982 6848 4988 6860
rect 4672 6820 4988 6848
rect 4672 6808 4678 6820
rect 4982 6808 4988 6820
rect 5040 6848 5046 6860
rect 5077 6851 5135 6857
rect 5077 6848 5089 6851
rect 5040 6820 5089 6848
rect 5040 6808 5046 6820
rect 5077 6817 5089 6820
rect 5123 6817 5135 6851
rect 5626 6848 5632 6860
rect 5077 6811 5135 6817
rect 5460 6820 5632 6848
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 1412 6712 1440 6743
rect 3602 6740 3608 6792
rect 3660 6740 3666 6792
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6780 3847 6783
rect 3835 6752 3924 6780
rect 3835 6749 3847 6752
rect 3789 6743 3847 6749
rect 1673 6715 1731 6721
rect 1412 6684 1532 6712
rect 1504 6656 1532 6684
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 1946 6712 1952 6724
rect 1719 6684 1952 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 1946 6672 1952 6684
rect 2004 6672 2010 6724
rect 3142 6712 3148 6724
rect 2898 6684 3148 6712
rect 3142 6672 3148 6684
rect 3200 6672 3206 6724
rect 3896 6656 3924 6752
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 4028 6752 5273 6780
rect 4028 6740 4034 6752
rect 5261 6749 5273 6752
rect 5307 6780 5319 6783
rect 5460 6780 5488 6820
rect 5626 6808 5632 6820
rect 5684 6848 5690 6860
rect 6181 6851 6239 6857
rect 5684 6820 6040 6848
rect 5684 6808 5690 6820
rect 6012 6792 6040 6820
rect 6181 6817 6193 6851
rect 6227 6848 6239 6851
rect 8297 6851 8355 6857
rect 8297 6848 8309 6851
rect 6227 6820 8309 6848
rect 6227 6817 6239 6820
rect 6181 6811 6239 6817
rect 8297 6817 8309 6820
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 5307 6752 5488 6780
rect 5537 6783 5595 6789
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5537 6749 5549 6783
rect 5583 6780 5595 6783
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5583 6752 5917 6780
rect 5583 6749 5595 6752
rect 5537 6743 5595 6749
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 5350 6712 5356 6724
rect 4724 6684 5356 6712
rect 4724 6656 4752 6684
rect 5350 6672 5356 6684
rect 5408 6712 5414 6724
rect 5552 6712 5580 6743
rect 5994 6740 6000 6792
rect 6052 6740 6058 6792
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 5408 6684 5580 6712
rect 6288 6712 6316 6743
rect 6362 6740 6368 6792
rect 6420 6740 6426 6792
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8018 6712 8024 6724
rect 6288 6684 6776 6712
rect 7866 6684 8024 6712
rect 5408 6672 5414 6684
rect 6748 6656 6776 6684
rect 8018 6672 8024 6684
rect 8076 6672 8082 6724
rect 8220 6656 8248 6743
rect 1486 6604 1492 6656
rect 1544 6604 1550 6656
rect 3234 6604 3240 6656
rect 3292 6604 3298 6656
rect 3878 6604 3884 6656
rect 3936 6604 3942 6656
rect 4433 6647 4491 6653
rect 4433 6613 4445 6647
rect 4479 6644 4491 6647
rect 4706 6644 4712 6656
rect 4479 6616 4712 6644
rect 4479 6613 4491 6616
rect 4433 6607 4491 6613
rect 4706 6604 4712 6616
rect 4764 6604 4770 6656
rect 5442 6604 5448 6656
rect 5500 6604 5506 6656
rect 6730 6604 6736 6656
rect 6788 6604 6794 6656
rect 7282 6604 7288 6656
rect 7340 6644 7346 6656
rect 8110 6644 8116 6656
rect 7340 6616 8116 6644
rect 7340 6604 7346 6616
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 8202 6604 8208 6656
rect 8260 6604 8266 6656
rect 8312 6644 8340 6811
rect 8404 6780 8432 6888
rect 11054 6876 11060 6928
rect 11112 6916 11118 6928
rect 11974 6916 11980 6928
rect 11112 6888 11980 6916
rect 11112 6876 11118 6888
rect 11974 6876 11980 6888
rect 12032 6876 12038 6928
rect 12406 6916 12434 6944
rect 12268 6888 12434 6916
rect 8481 6851 8539 6857
rect 8481 6817 8493 6851
rect 8527 6848 8539 6851
rect 9950 6848 9956 6860
rect 8527 6820 8800 6848
rect 8527 6817 8539 6820
rect 8481 6811 8539 6817
rect 8772 6792 8800 6820
rect 8864 6820 9956 6848
rect 8573 6783 8631 6789
rect 8573 6780 8585 6783
rect 8404 6752 8585 6780
rect 8573 6749 8585 6752
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 8754 6740 8760 6792
rect 8812 6740 8818 6792
rect 8481 6715 8539 6721
rect 8481 6681 8493 6715
rect 8527 6712 8539 6715
rect 8864 6712 8892 6820
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 10410 6848 10416 6860
rect 10336 6820 10416 6848
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6749 8999 6783
rect 10336 6766 10364 6820
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 10870 6808 10876 6860
rect 10928 6808 10934 6860
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12268 6848 12296 6888
rect 12894 6848 12900 6860
rect 12207 6820 12296 6848
rect 12406 6820 12900 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 8941 6743 8999 6749
rect 8527 6684 8892 6712
rect 8527 6681 8539 6684
rect 8481 6675 8539 6681
rect 8665 6647 8723 6653
rect 8665 6644 8677 6647
rect 8312 6616 8677 6644
rect 8665 6613 8677 6616
rect 8711 6613 8723 6647
rect 8956 6644 8984 6743
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 11057 6783 11115 6789
rect 11057 6780 11069 6783
rect 10560 6752 11069 6780
rect 10560 6740 10566 6752
rect 11057 6749 11069 6752
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11238 6740 11244 6792
rect 11296 6740 11302 6792
rect 11333 6783 11391 6789
rect 11333 6749 11345 6783
rect 11379 6780 11391 6783
rect 12406 6780 12434 6820
rect 12894 6808 12900 6820
rect 12952 6848 12958 6860
rect 12952 6820 14228 6848
rect 12952 6808 12958 6820
rect 11379 6752 12434 6780
rect 13909 6783 13967 6789
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 13909 6749 13921 6783
rect 13955 6780 13967 6783
rect 13998 6780 14004 6792
rect 13955 6752 14004 6780
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 14090 6740 14096 6792
rect 14148 6740 14154 6792
rect 11146 6712 11152 6724
rect 10612 6684 11152 6712
rect 9398 6644 9404 6656
rect 8956 6616 9404 6644
rect 8665 6607 8723 6613
rect 9398 6604 9404 6616
rect 9456 6644 9462 6656
rect 10612 6644 10640 6684
rect 11146 6672 11152 6684
rect 11204 6672 11210 6724
rect 14200 6721 14228 6820
rect 14369 6783 14427 6789
rect 14369 6749 14381 6783
rect 14415 6749 14427 6783
rect 14369 6743 14427 6749
rect 14185 6715 14243 6721
rect 13202 6684 13492 6712
rect 13464 6656 13492 6684
rect 14185 6681 14197 6715
rect 14231 6681 14243 6715
rect 14185 6675 14243 6681
rect 9456 6616 10640 6644
rect 9456 6604 9462 6616
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 13446 6644 13452 6656
rect 12676 6616 13452 6644
rect 12676 6604 12682 6616
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 13538 6604 13544 6656
rect 13596 6644 13602 6656
rect 14384 6644 14412 6743
rect 13596 6616 14412 6644
rect 13596 6604 13602 6616
rect 1104 6554 16836 6576
rect 1104 6502 1610 6554
rect 1662 6502 1674 6554
rect 1726 6502 1738 6554
rect 1790 6502 1802 6554
rect 1854 6502 1866 6554
rect 1918 6502 5610 6554
rect 5662 6502 5674 6554
rect 5726 6502 5738 6554
rect 5790 6502 5802 6554
rect 5854 6502 5866 6554
rect 5918 6502 9610 6554
rect 9662 6502 9674 6554
rect 9726 6502 9738 6554
rect 9790 6502 9802 6554
rect 9854 6502 9866 6554
rect 9918 6502 13610 6554
rect 13662 6502 13674 6554
rect 13726 6502 13738 6554
rect 13790 6502 13802 6554
rect 13854 6502 13866 6554
rect 13918 6502 16836 6554
rect 1104 6480 16836 6502
rect 2314 6400 2320 6452
rect 2372 6400 2378 6452
rect 2406 6400 2412 6452
rect 2464 6400 2470 6452
rect 4798 6400 4804 6452
rect 4856 6400 4862 6452
rect 5350 6400 5356 6452
rect 5408 6440 5414 6452
rect 5695 6443 5753 6449
rect 5695 6440 5707 6443
rect 5408 6412 5707 6440
rect 5408 6400 5414 6412
rect 5695 6409 5707 6412
rect 5741 6409 5753 6443
rect 5695 6403 5753 6409
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 5868 6412 8340 6440
rect 5868 6400 5874 6412
rect 934 6332 940 6384
rect 992 6372 998 6384
rect 1397 6375 1455 6381
rect 1397 6372 1409 6375
rect 992 6344 1409 6372
rect 992 6332 998 6344
rect 1397 6341 1409 6344
rect 1443 6341 1455 6375
rect 1397 6335 1455 6341
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6304 2007 6307
rect 2332 6304 2360 6400
rect 4522 6332 4528 6384
rect 4580 6332 4586 6384
rect 4816 6372 4844 6400
rect 4632 6344 4844 6372
rect 5905 6375 5963 6381
rect 4632 6313 4660 6344
rect 5905 6341 5917 6375
rect 5951 6372 5963 6375
rect 6086 6372 6092 6384
rect 5951 6344 6092 6372
rect 5951 6341 5963 6344
rect 5905 6335 5963 6341
rect 6086 6332 6092 6344
rect 6144 6332 6150 6384
rect 7193 6375 7251 6381
rect 7193 6341 7205 6375
rect 7239 6372 7251 6375
rect 7466 6372 7472 6384
rect 7239 6344 7472 6372
rect 7239 6341 7251 6344
rect 7193 6335 7251 6341
rect 1995 6276 2360 6304
rect 2685 6307 2743 6313
rect 1995 6273 2007 6276
rect 1949 6267 2007 6273
rect 2685 6273 2697 6307
rect 2731 6273 2743 6307
rect 2685 6267 2743 6273
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6304 4859 6307
rect 4982 6304 4988 6316
rect 4847 6276 4988 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 1780 6236 1808 6267
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 1780 6208 2605 6236
rect 2593 6205 2605 6208
rect 2639 6205 2651 6239
rect 2700 6236 2728 6267
rect 4982 6264 4988 6276
rect 5040 6304 5046 6316
rect 7208 6304 7236 6335
rect 7466 6332 7472 6344
rect 7524 6332 7530 6384
rect 8202 6372 8208 6384
rect 7576 6344 8208 6372
rect 5040 6276 7236 6304
rect 5040 6264 5046 6276
rect 6549 6239 6607 6245
rect 2700 6208 6500 6236
rect 2593 6199 2651 6205
rect 4430 6168 4436 6180
rect 2240 6140 4436 6168
rect 2240 6109 2268 6140
rect 4430 6128 4436 6140
rect 4488 6128 4494 6180
rect 5442 6128 5448 6180
rect 5500 6128 5506 6180
rect 5534 6128 5540 6180
rect 5592 6168 5598 6180
rect 5810 6168 5816 6180
rect 5592 6140 5816 6168
rect 5592 6128 5598 6140
rect 5810 6128 5816 6140
rect 5868 6128 5874 6180
rect 6472 6168 6500 6208
rect 6549 6205 6561 6239
rect 6595 6236 6607 6239
rect 6730 6236 6736 6248
rect 6595 6208 6736 6236
rect 6595 6205 6607 6208
rect 6549 6199 6607 6205
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7576 6245 7604 6344
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 8312 6372 8340 6412
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 9306 6440 9312 6452
rect 8812 6412 9312 6440
rect 8812 6400 8818 6412
rect 9306 6400 9312 6412
rect 9364 6440 9370 6452
rect 9861 6443 9919 6449
rect 9861 6440 9873 6443
rect 9364 6412 9873 6440
rect 9364 6400 9370 6412
rect 9861 6409 9873 6412
rect 9907 6409 9919 6443
rect 9861 6403 9919 6409
rect 10502 6400 10508 6452
rect 10560 6400 10566 6452
rect 10686 6400 10692 6452
rect 10744 6400 10750 6452
rect 10520 6372 10548 6400
rect 8312 6344 10548 6372
rect 8110 6264 8116 6316
rect 8168 6304 8174 6316
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8168 6276 8493 6304
rect 8168 6264 8174 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6304 10379 6307
rect 10704 6304 10732 6400
rect 16022 6304 16028 6316
rect 10367 6276 10732 6304
rect 12084 6276 16028 6304
rect 10367 6273 10379 6276
rect 10321 6267 10379 6273
rect 12084 6245 12112 6276
rect 16022 6264 16028 6276
rect 16080 6264 16086 6316
rect 7561 6239 7619 6245
rect 7561 6236 7573 6239
rect 7156 6208 7573 6236
rect 7156 6196 7162 6208
rect 7561 6205 7573 6208
rect 7607 6205 7619 6239
rect 7561 6199 7619 6205
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6236 7711 6239
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 7699 6208 7941 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 7929 6205 7941 6208
rect 7975 6205 7987 6239
rect 7929 6199 7987 6205
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 12084 6168 12112 6199
rect 12342 6196 12348 6248
rect 12400 6196 12406 6248
rect 6472 6140 12112 6168
rect 2225 6103 2283 6109
rect 2225 6069 2237 6103
rect 2271 6069 2283 6103
rect 2225 6063 2283 6069
rect 3237 6103 3295 6109
rect 3237 6069 3249 6103
rect 3283 6100 3295 6103
rect 3786 6100 3792 6112
rect 3283 6072 3792 6100
rect 3283 6069 3295 6072
rect 3237 6063 3295 6069
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 4706 6060 4712 6112
rect 4764 6060 4770 6112
rect 5460 6100 5488 6128
rect 5721 6103 5779 6109
rect 5721 6100 5733 6103
rect 5460 6072 5733 6100
rect 5721 6069 5733 6072
rect 5767 6069 5779 6103
rect 5721 6063 5779 6069
rect 7098 6060 7104 6112
rect 7156 6060 7162 6112
rect 7834 6060 7840 6112
rect 7892 6060 7898 6112
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 9582 6100 9588 6112
rect 8352 6072 9588 6100
rect 8352 6060 8358 6072
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 10229 6103 10287 6109
rect 10229 6069 10241 6103
rect 10275 6100 10287 6103
rect 12434 6100 12440 6112
rect 10275 6072 12440 6100
rect 10275 6069 10287 6072
rect 10229 6063 10287 6069
rect 12434 6060 12440 6072
rect 12492 6100 12498 6112
rect 12710 6100 12716 6112
rect 12492 6072 12716 6100
rect 12492 6060 12498 6072
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 944 6010 16836 6032
rect 944 5958 950 6010
rect 1002 5958 1014 6010
rect 1066 5958 1078 6010
rect 1130 5958 1142 6010
rect 1194 5958 1206 6010
rect 1258 5958 4950 6010
rect 5002 5958 5014 6010
rect 5066 5958 5078 6010
rect 5130 5958 5142 6010
rect 5194 5958 5206 6010
rect 5258 5958 8950 6010
rect 9002 5958 9014 6010
rect 9066 5958 9078 6010
rect 9130 5958 9142 6010
rect 9194 5958 9206 6010
rect 9258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 16836 6010
rect 944 5936 16836 5958
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 3660 5868 3801 5896
rect 3660 5856 3666 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 3789 5859 3847 5865
rect 4706 5856 4712 5908
rect 4764 5856 4770 5908
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5537 5899 5595 5905
rect 5537 5896 5549 5899
rect 5316 5868 5549 5896
rect 5316 5856 5322 5868
rect 5537 5865 5549 5868
rect 5583 5896 5595 5899
rect 5994 5896 6000 5908
rect 5583 5868 6000 5896
rect 5583 5865 5595 5868
rect 5537 5859 5595 5865
rect 5994 5856 6000 5868
rect 6052 5896 6058 5908
rect 6822 5896 6828 5908
rect 6052 5868 6828 5896
rect 6052 5856 6058 5868
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 10318 5896 10324 5908
rect 8956 5868 10324 5896
rect 3237 5831 3295 5837
rect 3237 5797 3249 5831
rect 3283 5828 3295 5831
rect 3878 5828 3884 5840
rect 3283 5800 3884 5828
rect 3283 5797 3295 5800
rect 3237 5791 3295 5797
rect 3878 5788 3884 5800
rect 3936 5828 3942 5840
rect 3936 5800 4384 5828
rect 3936 5788 3942 5800
rect 1486 5720 1492 5772
rect 1544 5760 1550 5772
rect 3786 5760 3792 5772
rect 1544 5732 3792 5760
rect 1544 5720 1550 5732
rect 3786 5720 3792 5732
rect 3844 5720 3850 5772
rect 4356 5769 4384 5800
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5729 4399 5763
rect 4724 5760 4752 5856
rect 7098 5828 7104 5840
rect 5184 5800 7104 5828
rect 5184 5769 5212 5800
rect 7098 5788 7104 5800
rect 7156 5788 7162 5840
rect 5169 5763 5227 5769
rect 4724 5732 4936 5760
rect 4341 5723 4399 5729
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 4908 5692 4936 5732
rect 5169 5729 5181 5763
rect 5215 5729 5227 5763
rect 6086 5760 6092 5772
rect 5169 5723 5227 5729
rect 5460 5732 6092 5760
rect 5011 5695 5069 5701
rect 5011 5692 5023 5695
rect 4908 5664 5023 5692
rect 5011 5661 5023 5664
rect 5057 5661 5069 5695
rect 5011 5655 5069 5661
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 5460 5701 5488 5732
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 7282 5760 7288 5772
rect 6656 5732 7288 5760
rect 5445 5695 5503 5701
rect 5445 5661 5457 5695
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 1765 5627 1823 5633
rect 1765 5593 1777 5627
rect 1811 5593 1823 5627
rect 3142 5624 3148 5636
rect 2990 5596 3148 5624
rect 1765 5587 1823 5593
rect 1780 5556 1808 5587
rect 3142 5584 3148 5596
rect 3200 5584 3206 5636
rect 4801 5627 4859 5633
rect 4801 5624 4813 5627
rect 3252 5596 4813 5624
rect 1946 5556 1952 5568
rect 1780 5528 1952 5556
rect 1946 5516 1952 5528
rect 2004 5516 2010 5568
rect 2590 5516 2596 5568
rect 2648 5556 2654 5568
rect 3252 5556 3280 5596
rect 4801 5593 4813 5596
rect 4847 5593 4859 5627
rect 4801 5587 4859 5593
rect 4893 5627 4951 5633
rect 4893 5593 4905 5627
rect 4939 5624 4951 5627
rect 5276 5624 5304 5652
rect 4939 5596 5304 5624
rect 6104 5624 6132 5720
rect 6656 5701 6684 5732
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 7926 5720 7932 5772
rect 7984 5760 7990 5772
rect 8956 5760 8984 5868
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 11146 5856 11152 5908
rect 11204 5896 11210 5908
rect 12161 5899 12219 5905
rect 12161 5896 12173 5899
rect 11204 5868 12173 5896
rect 11204 5856 11210 5868
rect 12161 5865 12173 5868
rect 12207 5896 12219 5899
rect 13446 5896 13452 5908
rect 12207 5868 13452 5896
rect 12207 5865 12219 5868
rect 12161 5859 12219 5865
rect 13446 5856 13452 5868
rect 13504 5896 13510 5908
rect 13998 5896 14004 5908
rect 13504 5868 14004 5896
rect 13504 5856 13510 5868
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 7984 5732 8984 5760
rect 9033 5763 9091 5769
rect 7984 5720 7990 5732
rect 9033 5729 9045 5763
rect 9079 5760 9091 5763
rect 9398 5760 9404 5772
rect 9079 5732 9404 5760
rect 9079 5729 9091 5732
rect 9033 5723 9091 5729
rect 9398 5720 9404 5732
rect 9456 5720 9462 5772
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 9732 5732 12434 5760
rect 9732 5720 9738 5732
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 6457 5695 6515 5701
rect 6457 5692 6469 5695
rect 6411 5664 6469 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 6457 5661 6469 5664
rect 6503 5661 6515 5695
rect 6457 5655 6515 5661
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 6822 5652 6828 5704
rect 6880 5652 6886 5704
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5692 7159 5695
rect 7190 5692 7196 5704
rect 7147 5664 7196 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 10410 5652 10416 5704
rect 10468 5652 10474 5704
rect 10873 5695 10931 5701
rect 10873 5661 10885 5695
rect 10919 5692 10931 5695
rect 10962 5692 10968 5704
rect 10919 5664 10968 5692
rect 10919 5661 10931 5664
rect 10873 5655 10931 5661
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 6104 5596 6684 5624
rect 4939 5593 4951 5596
rect 4893 5587 4951 5593
rect 6656 5568 6684 5596
rect 6730 5584 6736 5636
rect 6788 5584 6794 5636
rect 6963 5627 7021 5633
rect 6963 5593 6975 5627
rect 7009 5624 7021 5627
rect 7285 5627 7343 5633
rect 7285 5624 7297 5627
rect 7009 5596 7297 5624
rect 7009 5593 7021 5596
rect 6963 5587 7021 5593
rect 7285 5593 7297 5596
rect 7331 5593 7343 5627
rect 7285 5587 7343 5593
rect 9309 5627 9367 5633
rect 9309 5593 9321 5627
rect 9355 5593 9367 5627
rect 12406 5624 12434 5732
rect 16117 5627 16175 5633
rect 16117 5624 16129 5627
rect 12406 5596 16129 5624
rect 9309 5587 9367 5593
rect 16117 5593 16129 5596
rect 16163 5593 16175 5627
rect 16117 5587 16175 5593
rect 2648 5528 3280 5556
rect 2648 5516 2654 5528
rect 4522 5516 4528 5568
rect 4580 5516 4586 5568
rect 5721 5559 5779 5565
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 6086 5556 6092 5568
rect 5767 5528 6092 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 6638 5516 6644 5568
rect 6696 5556 6702 5568
rect 8386 5556 8392 5568
rect 6696 5528 8392 5556
rect 6696 5516 6702 5528
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 9324 5556 9352 5587
rect 9950 5556 9956 5568
rect 9324 5528 9956 5556
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10781 5559 10839 5565
rect 10781 5525 10793 5559
rect 10827 5556 10839 5559
rect 10870 5556 10876 5568
rect 10827 5528 10876 5556
rect 10827 5525 10839 5528
rect 10781 5519 10839 5525
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 16393 5559 16451 5565
rect 16393 5525 16405 5559
rect 16439 5556 16451 5559
rect 16482 5556 16488 5568
rect 16439 5528 16488 5556
rect 16439 5525 16451 5528
rect 16393 5519 16451 5525
rect 16482 5516 16488 5528
rect 16540 5516 16546 5568
rect 1104 5466 16836 5488
rect 1104 5414 1610 5466
rect 1662 5414 1674 5466
rect 1726 5414 1738 5466
rect 1790 5414 1802 5466
rect 1854 5414 1866 5466
rect 1918 5414 5610 5466
rect 5662 5414 5674 5466
rect 5726 5414 5738 5466
rect 5790 5414 5802 5466
rect 5854 5414 5866 5466
rect 5918 5414 9610 5466
rect 9662 5414 9674 5466
rect 9726 5414 9738 5466
rect 9790 5414 9802 5466
rect 9854 5414 9866 5466
rect 9918 5414 13610 5466
rect 13662 5414 13674 5466
rect 13726 5414 13738 5466
rect 13790 5414 13802 5466
rect 13854 5414 13866 5466
rect 13918 5414 16836 5466
rect 1104 5392 16836 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 1596 5284 1624 5315
rect 1946 5312 1952 5364
rect 2004 5312 2010 5364
rect 2038 5312 2044 5364
rect 2096 5352 2102 5364
rect 2225 5355 2283 5361
rect 2225 5352 2237 5355
rect 2096 5324 2237 5352
rect 2096 5312 2102 5324
rect 2225 5321 2237 5324
rect 2271 5321 2283 5355
rect 2225 5315 2283 5321
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 3510 5352 3516 5364
rect 2556 5324 3516 5352
rect 2556 5312 2562 5324
rect 2590 5284 2596 5296
rect 1596 5256 2596 5284
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 750 5176 756 5228
rect 808 5216 814 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 808 5188 1409 5216
rect 808 5176 814 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2148 5148 2176 5179
rect 2406 5176 2412 5228
rect 2464 5176 2470 5228
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 2774 5216 2780 5228
rect 2731 5188 2780 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 2884 5225 2912 5324
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 4522 5352 4528 5364
rect 3896 5324 4528 5352
rect 3786 5284 3792 5296
rect 3620 5256 3792 5284
rect 3620 5225 3648 5256
rect 3786 5244 3792 5256
rect 3844 5244 3850 5296
rect 3896 5293 3924 5324
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 5258 5312 5264 5364
rect 5316 5312 5322 5364
rect 5353 5355 5411 5361
rect 5353 5321 5365 5355
rect 5399 5352 5411 5355
rect 6730 5352 6736 5364
rect 5399 5324 6736 5352
rect 5399 5321 5411 5324
rect 5353 5315 5411 5321
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 8386 5312 8392 5364
rect 8444 5352 8450 5364
rect 9861 5355 9919 5361
rect 8444 5324 9352 5352
rect 8444 5312 8450 5324
rect 3881 5287 3939 5293
rect 3881 5253 3893 5287
rect 3927 5253 3939 5287
rect 5276 5284 5304 5312
rect 7561 5287 7619 5293
rect 5276 5256 5856 5284
rect 3881 5247 3939 5253
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5185 2927 5219
rect 2869 5179 2927 5185
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5185 3663 5219
rect 5350 5216 5356 5228
rect 5014 5202 5356 5216
rect 3605 5179 3663 5185
rect 5000 5188 5356 5202
rect 3234 5148 3240 5160
rect 2148 5120 3240 5148
rect 3234 5108 3240 5120
rect 3292 5108 3298 5160
rect 2593 5083 2651 5089
rect 2593 5049 2605 5083
rect 2639 5080 2651 5083
rect 3326 5080 3332 5092
rect 2639 5052 3332 5080
rect 2639 5049 2651 5052
rect 2593 5043 2651 5049
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 3142 4972 3148 5024
rect 3200 5012 3206 5024
rect 5000 5012 5028 5188
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5828 5225 5856 5256
rect 7561 5253 7573 5287
rect 7607 5284 7619 5287
rect 7834 5284 7840 5296
rect 7607 5256 7840 5284
rect 7607 5253 7619 5256
rect 7561 5247 7619 5253
rect 7834 5244 7840 5256
rect 7892 5244 7898 5296
rect 8018 5244 8024 5296
rect 8076 5244 8082 5296
rect 9324 5293 9352 5324
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 9950 5352 9956 5364
rect 9907 5324 9956 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 11072 5324 11376 5352
rect 9309 5287 9367 5293
rect 9309 5253 9321 5287
rect 9355 5284 9367 5287
rect 11072 5284 11100 5324
rect 11348 5293 11376 5324
rect 12618 5312 12624 5364
rect 12676 5352 12682 5364
rect 12802 5352 12808 5364
rect 12676 5324 12808 5352
rect 12676 5312 12682 5324
rect 12802 5312 12808 5324
rect 12860 5312 12866 5364
rect 9355 5256 11100 5284
rect 11133 5287 11191 5293
rect 9355 5253 9367 5256
rect 9309 5247 9367 5253
rect 11133 5253 11145 5287
rect 11179 5284 11191 5287
rect 11333 5287 11391 5293
rect 11179 5253 11192 5284
rect 11133 5247 11192 5253
rect 11333 5253 11345 5287
rect 11379 5253 11391 5287
rect 12636 5284 12664 5312
rect 12558 5256 12664 5284
rect 11333 5247 11391 5253
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6012 5148 6040 5179
rect 6362 5176 6368 5228
rect 6420 5216 6426 5228
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 6420 5188 7297 5216
rect 6420 5176 6426 5188
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5185 9459 5219
rect 9401 5179 9459 5185
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5185 9551 5219
rect 9493 5179 9551 5185
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5216 9735 5219
rect 9723 5188 11008 5216
rect 9723 5185 9735 5188
rect 9677 5179 9735 5185
rect 6638 5148 6644 5160
rect 6012 5120 6644 5148
rect 6638 5108 6644 5120
rect 6696 5148 6702 5160
rect 6914 5148 6920 5160
rect 6696 5120 6920 5148
rect 6696 5108 6702 5120
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7190 5108 7196 5160
rect 7248 5148 7254 5160
rect 9416 5148 9444 5179
rect 7248 5120 9444 5148
rect 7248 5108 7254 5120
rect 9508 5080 9536 5179
rect 10318 5108 10324 5160
rect 10376 5108 10382 5160
rect 10870 5108 10876 5160
rect 10928 5108 10934 5160
rect 10229 5083 10287 5089
rect 10229 5080 10241 5083
rect 5736 5052 7420 5080
rect 5736 5024 5764 5052
rect 3200 4984 5028 5012
rect 3200 4972 3206 4984
rect 5718 4972 5724 5024
rect 5776 4972 5782 5024
rect 5905 5015 5963 5021
rect 5905 4981 5917 5015
rect 5951 5012 5963 5015
rect 6362 5012 6368 5024
rect 5951 4984 6368 5012
rect 5951 4981 5963 4984
rect 5905 4975 5963 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 7392 5012 7420 5052
rect 9324 5052 10241 5080
rect 9324 5024 9352 5052
rect 10229 5049 10241 5052
rect 10275 5049 10287 5083
rect 10229 5043 10287 5049
rect 8846 5012 8852 5024
rect 7392 4984 8852 5012
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 9306 4972 9312 5024
rect 9364 4972 9370 5024
rect 10336 5012 10364 5108
rect 10980 5089 11008 5188
rect 11164 5160 11192 5247
rect 11146 5108 11152 5160
rect 11204 5108 11210 5160
rect 12618 5108 12624 5160
rect 12676 5148 12682 5160
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12676 5120 13001 5148
rect 12676 5108 12682 5120
rect 12989 5117 13001 5120
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 13265 5151 13323 5157
rect 13265 5117 13277 5151
rect 13311 5148 13323 5151
rect 13446 5148 13452 5160
rect 13311 5120 13452 5148
rect 13311 5117 13323 5120
rect 13265 5111 13323 5117
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 10965 5083 11023 5089
rect 10965 5049 10977 5083
rect 11011 5049 11023 5083
rect 10965 5043 11023 5049
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 10336 4984 11161 5012
rect 11149 4981 11161 4984
rect 11195 4981 11207 5015
rect 11149 4975 11207 4981
rect 11514 4972 11520 5024
rect 11572 4972 11578 5024
rect 944 4922 16836 4944
rect 944 4870 950 4922
rect 1002 4870 1014 4922
rect 1066 4870 1078 4922
rect 1130 4870 1142 4922
rect 1194 4870 1206 4922
rect 1258 4870 4950 4922
rect 5002 4870 5014 4922
rect 5066 4870 5078 4922
rect 5130 4870 5142 4922
rect 5194 4870 5206 4922
rect 5258 4870 8950 4922
rect 9002 4870 9014 4922
rect 9066 4870 9078 4922
rect 9130 4870 9142 4922
rect 9194 4870 9206 4922
rect 9258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 16836 4922
rect 944 4848 16836 4870
rect 3418 4808 3424 4820
rect 2884 4780 3424 4808
rect 2884 4681 2912 4780
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 3510 4768 3516 4820
rect 3568 4768 3574 4820
rect 6270 4808 6276 4820
rect 5828 4780 6276 4808
rect 5718 4740 5724 4752
rect 2976 4712 5724 4740
rect 2685 4675 2743 4681
rect 2685 4672 2697 4675
rect 2240 4644 2697 4672
rect 2240 4613 2268 4644
rect 2685 4641 2697 4644
rect 2731 4641 2743 4675
rect 2685 4635 2743 4641
rect 2869 4675 2927 4681
rect 2869 4641 2881 4675
rect 2915 4641 2927 4675
rect 2869 4635 2927 4641
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4604 2007 4607
rect 2041 4607 2099 4613
rect 2041 4604 2053 4607
rect 1995 4576 2053 4604
rect 1995 4573 2007 4576
rect 1949 4567 2007 4573
rect 2041 4573 2053 4576
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2314 4564 2320 4616
rect 2372 4564 2378 4616
rect 2976 4613 3004 4712
rect 5718 4700 5724 4712
rect 5776 4700 5782 4752
rect 5828 4684 5856 4780
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 7926 4808 7932 4820
rect 7607 4780 7932 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8294 4768 8300 4820
rect 8352 4768 8358 4820
rect 8570 4768 8576 4820
rect 8628 4808 8634 4820
rect 11146 4808 11152 4820
rect 8628 4780 11152 4808
rect 8628 4768 8634 4780
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 11514 4768 11520 4820
rect 11572 4768 11578 4820
rect 12342 4768 12348 4820
rect 12400 4768 12406 4820
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 12986 4808 12992 4820
rect 12768 4780 12992 4808
rect 12768 4768 12774 4780
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 7653 4743 7711 4749
rect 7653 4740 7665 4743
rect 7116 4712 7665 4740
rect 3050 4632 3056 4684
rect 3108 4632 3114 4684
rect 5810 4632 5816 4684
rect 5868 4632 5874 4684
rect 6086 4632 6092 4684
rect 6144 4632 6150 4684
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 7116 4672 7144 4712
rect 7653 4709 7665 4712
rect 7699 4709 7711 4743
rect 8312 4740 8340 4768
rect 9171 4743 9229 4749
rect 9171 4740 9183 4743
rect 8312 4712 9183 4740
rect 7653 4703 7711 4709
rect 9171 4709 9183 4712
rect 9217 4709 9229 4743
rect 9171 4703 9229 4709
rect 10318 4700 10324 4752
rect 10376 4740 10382 4752
rect 11422 4740 11428 4752
rect 10376 4712 11428 4740
rect 10376 4700 10382 4712
rect 11422 4700 11428 4712
rect 11480 4700 11486 4752
rect 6880 4644 7144 4672
rect 6880 4632 6886 4644
rect 7282 4632 7288 4684
rect 7340 4672 7346 4684
rect 7340 4644 7880 4672
rect 7340 4632 7346 4644
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4573 3019 4607
rect 2961 4567 3019 4573
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 2976 4536 3004 4567
rect 2832 4508 3004 4536
rect 3160 4536 3188 4567
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 3329 4607 3387 4613
rect 3329 4604 3341 4607
rect 3292 4576 3341 4604
rect 3292 4564 3298 4576
rect 3329 4573 3341 4576
rect 3375 4573 3387 4607
rect 3329 4567 3387 4573
rect 7190 4564 7196 4616
rect 7248 4604 7254 4616
rect 7742 4604 7748 4616
rect 7248 4576 7748 4604
rect 7248 4564 7254 4576
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 7852 4613 7880 4644
rect 8294 4632 8300 4684
rect 8352 4632 8358 4684
rect 8386 4632 8392 4684
rect 8444 4632 8450 4684
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 9306 4672 9312 4684
rect 8527 4644 9312 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 11054 4672 11060 4684
rect 10704 4644 11060 4672
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 3160 4508 3372 4536
rect 2832 4496 2838 4508
rect 3344 4480 3372 4508
rect 5534 4496 5540 4548
rect 5592 4496 5598 4548
rect 7944 4536 7972 4567
rect 8570 4564 8576 4616
rect 8628 4564 8634 4616
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 7484 4508 7972 4536
rect 1765 4471 1823 4477
rect 1765 4437 1777 4471
rect 1811 4468 1823 4471
rect 1946 4468 1952 4480
rect 1811 4440 1952 4468
rect 1811 4437 1823 4440
rect 1765 4431 1823 4437
rect 1946 4428 1952 4440
rect 2004 4428 2010 4480
rect 3326 4428 3332 4480
rect 3384 4428 3390 4480
rect 5552 4468 5580 4496
rect 7484 4468 7512 4508
rect 8110 4496 8116 4548
rect 8168 4536 8174 4548
rect 8956 4536 8984 4567
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 10704 4604 10732 4644
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11532 4672 11560 4768
rect 12526 4700 12532 4752
rect 12584 4740 12590 4752
rect 14182 4740 14188 4752
rect 12584 4712 13124 4740
rect 12584 4700 12590 4712
rect 11164 4644 12020 4672
rect 9088 4576 10732 4604
rect 9088 4564 9094 4576
rect 10778 4564 10784 4616
rect 10836 4564 10842 4616
rect 10870 4564 10876 4616
rect 10928 4564 10934 4616
rect 11164 4613 11192 4644
rect 11992 4613 12020 4644
rect 12986 4632 12992 4684
rect 13044 4632 13050 4684
rect 13096 4681 13124 4712
rect 13188 4712 14188 4740
rect 13081 4675 13139 4681
rect 13081 4641 13093 4675
rect 13127 4641 13139 4675
rect 13081 4635 13139 4641
rect 11149 4607 11207 4613
rect 11149 4573 11161 4607
rect 11195 4573 11207 4607
rect 11517 4607 11575 4613
rect 11517 4604 11529 4607
rect 11149 4567 11207 4573
rect 11256 4576 11529 4604
rect 8168 4508 8984 4536
rect 8168 4496 8174 4508
rect 10502 4496 10508 4548
rect 10560 4536 10566 4548
rect 11256 4536 11284 4576
rect 11517 4573 11529 4576
rect 11563 4573 11575 4607
rect 11517 4567 11575 4573
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4573 12035 4607
rect 11977 4567 12035 4573
rect 10560 4508 11284 4536
rect 11333 4539 11391 4545
rect 10560 4496 10566 4508
rect 11333 4505 11345 4539
rect 11379 4536 11391 4539
rect 11716 4536 11744 4567
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12805 4607 12863 4613
rect 12805 4604 12817 4607
rect 12492 4576 12817 4604
rect 12492 4564 12498 4576
rect 12805 4573 12817 4576
rect 12851 4573 12863 4607
rect 12805 4567 12863 4573
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4604 12955 4607
rect 13188 4604 13216 4712
rect 14182 4700 14188 4712
rect 14240 4700 14246 4752
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4672 13323 4675
rect 13311 4644 13584 4672
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 12943 4576 13216 4604
rect 12943 4573 12955 4576
rect 12897 4567 12955 4573
rect 13354 4564 13360 4616
rect 13412 4564 13418 4616
rect 13556 4613 13584 4644
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4604 13783 4607
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13771 4576 14289 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 16114 4564 16120 4616
rect 16172 4564 16178 4616
rect 12161 4539 12219 4545
rect 12161 4536 12173 4539
rect 11379 4508 11744 4536
rect 11808 4508 12173 4536
rect 11379 4505 11391 4508
rect 11333 4499 11391 4505
rect 5552 4440 7512 4468
rect 8757 4471 8815 4477
rect 8757 4437 8769 4471
rect 8803 4468 8815 4471
rect 9950 4468 9956 4480
rect 8803 4440 9956 4468
rect 8803 4437 8815 4440
rect 8757 4431 8815 4437
rect 9950 4428 9956 4440
rect 10008 4428 10014 4480
rect 10134 4428 10140 4480
rect 10192 4428 10198 4480
rect 10962 4428 10968 4480
rect 11020 4468 11026 4480
rect 11808 4468 11836 4508
rect 12161 4505 12173 4508
rect 12207 4505 12219 4539
rect 12161 4499 12219 4505
rect 11020 4440 11836 4468
rect 11020 4428 11026 4440
rect 11882 4428 11888 4480
rect 11940 4428 11946 4480
rect 14090 4428 14096 4480
rect 14148 4428 14154 4480
rect 16393 4471 16451 4477
rect 16393 4437 16405 4471
rect 16439 4468 16451 4471
rect 16758 4468 16764 4480
rect 16439 4440 16764 4468
rect 16439 4437 16451 4440
rect 16393 4431 16451 4437
rect 16758 4428 16764 4440
rect 16816 4428 16822 4480
rect 1104 4378 16836 4400
rect 1104 4326 1610 4378
rect 1662 4326 1674 4378
rect 1726 4326 1738 4378
rect 1790 4326 1802 4378
rect 1854 4326 1866 4378
rect 1918 4326 5610 4378
rect 5662 4326 5674 4378
rect 5726 4326 5738 4378
rect 5790 4326 5802 4378
rect 5854 4326 5866 4378
rect 5918 4326 9610 4378
rect 9662 4326 9674 4378
rect 9726 4326 9738 4378
rect 9790 4326 9802 4378
rect 9854 4326 9866 4378
rect 9918 4326 13610 4378
rect 13662 4326 13674 4378
rect 13726 4326 13738 4378
rect 13790 4326 13802 4378
rect 13854 4326 13866 4378
rect 13918 4326 16836 4378
rect 1104 4304 16836 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 2832 4236 3648 4264
rect 2832 4224 2838 4236
rect 1857 4199 1915 4205
rect 1857 4165 1869 4199
rect 1903 4196 1915 4199
rect 1946 4196 1952 4208
rect 1903 4168 1952 4196
rect 1903 4165 1915 4168
rect 1857 4159 1915 4165
rect 1946 4156 1952 4168
rect 2004 4156 2010 4208
rect 3142 4196 3148 4208
rect 3082 4168 3148 4196
rect 3142 4156 3148 4168
rect 3200 4156 3206 4208
rect 3620 4205 3648 4236
rect 3896 4236 6040 4264
rect 3605 4199 3663 4205
rect 3605 4165 3617 4199
rect 3651 4165 3663 4199
rect 3605 4159 3663 4165
rect 3326 4088 3332 4140
rect 3384 4128 3390 4140
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 3384 4100 3433 4128
rect 3384 4088 3390 4100
rect 3421 4097 3433 4100
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 3786 4088 3792 4140
rect 3844 4128 3850 4140
rect 3896 4137 3924 4236
rect 6012 4208 6040 4236
rect 7282 4224 7288 4276
rect 7340 4224 7346 4276
rect 8386 4224 8392 4276
rect 8444 4264 8450 4276
rect 8444 4236 9168 4264
rect 8444 4224 8450 4236
rect 5442 4196 5448 4208
rect 5382 4168 5448 4196
rect 5442 4156 5448 4168
rect 5500 4196 5506 4208
rect 5500 4168 5948 4196
rect 5500 4156 5506 4168
rect 3881 4131 3939 4137
rect 3881 4128 3893 4131
rect 3844 4100 3893 4128
rect 3844 4088 3850 4100
rect 3881 4097 3893 4100
rect 3927 4097 3939 4131
rect 5920 4128 5948 4168
rect 5994 4156 6000 4208
rect 6052 4156 6058 4208
rect 7006 4196 7012 4208
rect 6104 4168 7012 4196
rect 6104 4128 6132 4168
rect 7006 4156 7012 4168
rect 7064 4156 7070 4208
rect 7300 4196 7328 4224
rect 7300 4168 8340 4196
rect 6641 4131 6699 4137
rect 6641 4128 6653 4131
rect 5920 4100 6132 4128
rect 6472 4100 6653 4128
rect 3881 4091 3939 4097
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4060 1639 4063
rect 3804 4060 3832 4088
rect 6472 4072 6500 4100
rect 6641 4097 6653 4100
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 6822 4088 6828 4140
rect 6880 4088 6886 4140
rect 7101 4131 7159 4137
rect 7101 4126 7113 4131
rect 7024 4098 7113 4126
rect 1627 4032 3832 4060
rect 4157 4063 4215 4069
rect 1627 4029 1639 4032
rect 1581 4023 1639 4029
rect 4157 4029 4169 4063
rect 4203 4060 4215 4063
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 4203 4032 6377 4060
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 6454 4020 6460 4072
rect 6512 4020 6518 4072
rect 6546 4020 6552 4072
rect 6604 4020 6610 4072
rect 6730 4020 6736 4072
rect 6788 4020 6794 4072
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 5629 3995 5687 4001
rect 5629 3992 5641 3995
rect 5592 3964 5641 3992
rect 5592 3952 5598 3964
rect 5629 3961 5641 3964
rect 5675 3961 5687 3995
rect 6564 3992 6592 4020
rect 7024 3992 7052 4098
rect 7101 4097 7113 4098
rect 7147 4126 7159 4131
rect 7285 4131 7343 4137
rect 7147 4098 7236 4126
rect 7147 4097 7159 4098
rect 7101 4091 7159 4097
rect 7208 4060 7236 4098
rect 7285 4097 7297 4131
rect 7331 4128 7343 4131
rect 7374 4128 7380 4140
rect 7331 4100 7380 4128
rect 7331 4097 7343 4100
rect 7285 4091 7343 4097
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 8312 4137 8340 4168
rect 8297 4131 8355 4137
rect 7944 4100 8248 4128
rect 7944 4060 7972 4100
rect 7208 4032 7972 4060
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 8067 4032 8125 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8113 4029 8125 4032
rect 8159 4029 8171 4063
rect 8220 4060 8248 4100
rect 8297 4097 8309 4131
rect 8343 4128 8355 4131
rect 8386 4128 8392 4140
rect 8343 4100 8392 4128
rect 8343 4097 8355 4100
rect 8297 4091 8355 4097
rect 8386 4088 8392 4100
rect 8444 4088 8450 4140
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8527 4100 9045 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 8570 4060 8576 4072
rect 8220 4032 8576 4060
rect 8113 4023 8171 4029
rect 6564 3964 7052 3992
rect 5629 3955 5687 3961
rect 7190 3952 7196 4004
rect 7248 3992 7254 4004
rect 7377 3995 7435 4001
rect 7377 3992 7389 3995
rect 7248 3964 7389 3992
rect 7248 3952 7254 3964
rect 7377 3961 7389 3964
rect 7423 3961 7435 3995
rect 7377 3955 7435 3961
rect 8036 3936 8064 4023
rect 8570 4020 8576 4032
rect 8628 4060 8634 4072
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 8628 4032 8769 4060
rect 8628 4020 8634 4032
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 8849 4063 8907 4069
rect 8849 4029 8861 4063
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 8941 4063 8999 4069
rect 8941 4029 8953 4063
rect 8987 4060 8999 4063
rect 9140 4060 9168 4236
rect 9950 4224 9956 4276
rect 10008 4224 10014 4276
rect 11882 4224 11888 4276
rect 11940 4224 11946 4276
rect 9769 4199 9827 4205
rect 9769 4165 9781 4199
rect 9815 4196 9827 4199
rect 9968 4196 9996 4224
rect 9815 4168 9996 4196
rect 9815 4165 9827 4168
rect 9769 4159 9827 4165
rect 11517 4131 11575 4137
rect 8987 4032 9168 4060
rect 8987 4029 8999 4032
rect 8941 4023 8999 4029
rect 3326 3884 3332 3936
rect 3384 3884 3390 3936
rect 3789 3927 3847 3933
rect 3789 3893 3801 3927
rect 3835 3924 3847 3927
rect 3878 3924 3884 3936
rect 3835 3896 3884 3924
rect 3835 3893 3847 3896
rect 3789 3887 3847 3893
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 8018 3884 8024 3936
rect 8076 3884 8082 3936
rect 8570 3884 8576 3936
rect 8628 3884 8634 3936
rect 8864 3924 8892 4023
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9493 4063 9551 4069
rect 9493 4060 9505 4063
rect 9456 4032 9505 4060
rect 9456 4020 9462 4032
rect 9493 4029 9505 4032
rect 9539 4029 9551 4063
rect 9493 4023 9551 4029
rect 10410 4020 10416 4072
rect 10468 4060 10474 4072
rect 10888 4060 10916 4114
rect 11517 4097 11529 4131
rect 11563 4128 11575 4131
rect 11900 4128 11928 4224
rect 13817 4199 13875 4205
rect 13817 4165 13829 4199
rect 13863 4196 13875 4199
rect 14090 4196 14096 4208
rect 13863 4168 14096 4196
rect 13863 4165 13875 4168
rect 13817 4159 13875 4165
rect 14090 4156 14096 4168
rect 14148 4156 14154 4208
rect 12710 4128 12716 4140
rect 11563 4100 11928 4128
rect 11992 4100 12716 4128
rect 11563 4097 11575 4100
rect 11517 4091 11575 4097
rect 11992 4060 12020 4100
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 12618 4060 12624 4072
rect 10468 4032 12020 4060
rect 12406 4032 12624 4060
rect 10468 4020 10474 4032
rect 11701 3995 11759 4001
rect 11701 3961 11713 3995
rect 11747 3992 11759 3995
rect 12406 3992 12434 4032
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 14093 4063 14151 4069
rect 14093 4060 14105 4063
rect 13504 4032 14105 4060
rect 13504 4020 13510 4032
rect 14093 4029 14105 4032
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 11747 3964 12434 3992
rect 11747 3961 11759 3964
rect 11701 3955 11759 3961
rect 10134 3924 10140 3936
rect 8864 3896 10140 3924
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 10836 3896 11253 3924
rect 10836 3884 10842 3896
rect 11241 3893 11253 3896
rect 11287 3893 11299 3927
rect 11241 3887 11299 3893
rect 12345 3927 12403 3933
rect 12345 3893 12357 3927
rect 12391 3924 12403 3927
rect 12434 3924 12440 3936
rect 12391 3896 12440 3924
rect 12391 3893 12403 3896
rect 12345 3887 12403 3893
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 944 3834 16836 3856
rect 944 3782 950 3834
rect 1002 3782 1014 3834
rect 1066 3782 1078 3834
rect 1130 3782 1142 3834
rect 1194 3782 1206 3834
rect 1258 3782 4950 3834
rect 5002 3782 5014 3834
rect 5066 3782 5078 3834
rect 5130 3782 5142 3834
rect 5194 3782 5206 3834
rect 5258 3782 8950 3834
rect 9002 3782 9014 3834
rect 9066 3782 9078 3834
rect 9130 3782 9142 3834
rect 9194 3782 9206 3834
rect 9258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 16836 3834
rect 944 3760 16836 3782
rect 3878 3680 3884 3732
rect 3936 3680 3942 3732
rect 6178 3680 6184 3732
rect 6236 3720 6242 3732
rect 6273 3723 6331 3729
rect 6273 3720 6285 3723
rect 6236 3692 6285 3720
rect 6236 3680 6242 3692
rect 6273 3689 6285 3692
rect 6319 3689 6331 3723
rect 6273 3683 6331 3689
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 7190 3720 7196 3732
rect 6512 3692 7196 3720
rect 6512 3680 6518 3692
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 8110 3680 8116 3732
rect 8168 3680 8174 3732
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 9217 3723 9275 3729
rect 9217 3720 9229 3723
rect 8352 3692 9229 3720
rect 8352 3680 8358 3692
rect 9217 3689 9229 3692
rect 9263 3689 9275 3723
rect 9217 3683 9275 3689
rect 9324 3692 9536 3720
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3516 1823 3519
rect 3326 3516 3332 3528
rect 1811 3488 3332 3516
rect 1811 3485 1823 3488
rect 1765 3479 1823 3485
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3516 3847 3519
rect 3896 3516 3924 3680
rect 9324 3652 9352 3692
rect 5368 3624 9352 3652
rect 9508 3652 9536 3692
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 10870 3720 10876 3732
rect 9732 3692 10876 3720
rect 9732 3680 9738 3692
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 12434 3652 12440 3664
rect 9508 3624 11468 3652
rect 3835 3488 3924 3516
rect 4617 3519 4675 3525
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 5074 3516 5080 3528
rect 4663 3488 5080 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 1397 3451 1455 3457
rect 1397 3448 1409 3451
rect 992 3420 1409 3448
rect 992 3408 998 3420
rect 1397 3417 1409 3420
rect 1443 3417 1455 3451
rect 5368 3448 5396 3624
rect 5534 3544 5540 3596
rect 5592 3584 5598 3596
rect 6638 3584 6644 3596
rect 5592 3556 6040 3584
rect 5592 3544 5598 3556
rect 5442 3476 5448 3528
rect 5500 3476 5506 3528
rect 5644 3525 5672 3556
rect 6012 3525 6040 3556
rect 6104 3556 6644 3584
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3516 5779 3519
rect 5997 3519 6055 3525
rect 5767 3488 5948 3516
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 1397 3411 1455 3417
rect 3712 3420 5396 3448
rect 5460 3448 5488 3476
rect 5813 3451 5871 3457
rect 5813 3448 5825 3451
rect 5460 3420 5825 3448
rect 3712 3392 3740 3420
rect 5813 3417 5825 3420
rect 5859 3417 5871 3451
rect 5920 3448 5948 3488
rect 5997 3485 6009 3519
rect 6043 3485 6055 3519
rect 5997 3479 6055 3485
rect 6104 3448 6132 3556
rect 6638 3544 6644 3556
rect 6696 3584 6702 3596
rect 6696 3556 7696 3584
rect 6696 3544 6702 3556
rect 7668 3525 7696 3556
rect 8386 3544 8392 3596
rect 8444 3544 8450 3596
rect 9585 3587 9643 3593
rect 9585 3553 9597 3587
rect 9631 3584 9643 3587
rect 10686 3584 10692 3596
rect 9631 3556 10692 3584
rect 9631 3553 9643 3556
rect 9585 3547 9643 3553
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 10870 3544 10876 3596
rect 10928 3584 10934 3596
rect 10928 3556 11100 3584
rect 10928 3544 10934 3556
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3516 6239 3519
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 6227 3488 6469 3516
rect 6227 3485 6239 3488
rect 6181 3479 6239 3485
rect 6457 3485 6469 3488
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 7653 3519 7711 3525
rect 7653 3485 7665 3519
rect 7699 3516 7711 3519
rect 8404 3516 8432 3544
rect 9401 3519 9459 3525
rect 9401 3516 9413 3519
rect 7699 3488 8156 3516
rect 8404 3488 9413 3516
rect 7699 3485 7711 3488
rect 7653 3479 7711 3485
rect 5920 3420 6132 3448
rect 7392 3448 7420 3479
rect 7745 3451 7803 3457
rect 7745 3448 7757 3451
rect 7392 3420 7757 3448
rect 5813 3411 5871 3417
rect 7745 3417 7757 3420
rect 7791 3448 7803 3451
rect 7834 3448 7840 3460
rect 7791 3420 7840 3448
rect 7791 3417 7803 3420
rect 7745 3411 7803 3417
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 7929 3451 7987 3457
rect 7929 3417 7941 3451
rect 7975 3448 7987 3451
rect 7975 3420 8064 3448
rect 7975 3417 7987 3420
rect 7929 3411 7987 3417
rect 8036 3392 8064 3420
rect 3694 3340 3700 3392
rect 3752 3340 3758 3392
rect 3973 3383 4031 3389
rect 3973 3349 3985 3383
rect 4019 3380 4031 3383
rect 4062 3380 4068 3392
rect 4019 3352 4068 3380
rect 4019 3349 4031 3352
rect 3973 3343 4031 3349
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 4430 3340 4436 3392
rect 4488 3340 4494 3392
rect 5261 3383 5319 3389
rect 5261 3349 5273 3383
rect 5307 3380 5319 3383
rect 5534 3380 5540 3392
rect 5307 3352 5540 3380
rect 5307 3349 5319 3352
rect 5261 3343 5319 3349
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 7190 3340 7196 3392
rect 7248 3340 7254 3392
rect 7561 3383 7619 3389
rect 7561 3349 7573 3383
rect 7607 3380 7619 3383
rect 8018 3380 8024 3392
rect 7607 3352 8024 3380
rect 7607 3349 7619 3352
rect 7561 3343 7619 3349
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 8128 3380 8156 3488
rect 9401 3485 9413 3488
rect 9447 3485 9459 3519
rect 9401 3479 9459 3485
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3516 9735 3519
rect 10594 3516 10600 3528
rect 9723 3488 10600 3516
rect 9723 3485 9735 3488
rect 9677 3479 9735 3485
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3516 10839 3519
rect 10962 3516 10968 3528
rect 10827 3488 10968 3516
rect 10827 3485 10839 3488
rect 10781 3479 10839 3485
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11072 3525 11100 3556
rect 11057 3519 11115 3525
rect 11057 3485 11069 3519
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 11330 3476 11336 3528
rect 11388 3476 11394 3528
rect 11440 3516 11468 3624
rect 12360 3624 12440 3652
rect 12360 3516 12388 3624
rect 12434 3612 12440 3624
rect 12492 3612 12498 3664
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 11440 3488 14105 3516
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 15930 3476 15936 3528
rect 15988 3476 15994 3528
rect 9490 3408 9496 3460
rect 9548 3448 9554 3460
rect 12802 3448 12808 3460
rect 9548 3420 12808 3448
rect 9548 3408 9554 3420
rect 12802 3408 12808 3420
rect 12860 3408 12866 3460
rect 13354 3408 13360 3460
rect 13412 3448 13418 3460
rect 14277 3451 14335 3457
rect 14277 3448 14289 3451
rect 13412 3420 14289 3448
rect 13412 3408 13418 3420
rect 14277 3417 14289 3420
rect 14323 3417 14335 3451
rect 14277 3411 14335 3417
rect 9674 3380 9680 3392
rect 8128 3352 9680 3380
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 9769 3383 9827 3389
rect 9769 3349 9781 3383
rect 9815 3380 9827 3383
rect 9950 3380 9956 3392
rect 9815 3352 9956 3380
rect 9815 3349 9827 3352
rect 9769 3343 9827 3349
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 10594 3340 10600 3392
rect 10652 3340 10658 3392
rect 10686 3340 10692 3392
rect 10744 3380 10750 3392
rect 10965 3383 11023 3389
rect 10965 3380 10977 3383
rect 10744 3352 10977 3380
rect 10744 3340 10750 3352
rect 10965 3349 10977 3352
rect 11011 3349 11023 3383
rect 10965 3343 11023 3349
rect 11422 3340 11428 3392
rect 11480 3340 11486 3392
rect 14458 3340 14464 3392
rect 14516 3340 14522 3392
rect 16022 3340 16028 3392
rect 16080 3340 16086 3392
rect 1104 3290 16836 3312
rect 1104 3238 1610 3290
rect 1662 3238 1674 3290
rect 1726 3238 1738 3290
rect 1790 3238 1802 3290
rect 1854 3238 1866 3290
rect 1918 3238 5610 3290
rect 5662 3238 5674 3290
rect 5726 3238 5738 3290
rect 5790 3238 5802 3290
rect 5854 3238 5866 3290
rect 5918 3238 9610 3290
rect 9662 3238 9674 3290
rect 9726 3238 9738 3290
rect 9790 3238 9802 3290
rect 9854 3238 9866 3290
rect 9918 3238 13610 3290
rect 13662 3238 13674 3290
rect 13726 3238 13738 3290
rect 13790 3238 13802 3290
rect 13854 3238 13866 3290
rect 13918 3238 16836 3290
rect 1104 3216 16836 3238
rect 2133 3179 2191 3185
rect 2133 3145 2145 3179
rect 2179 3176 2191 3179
rect 3234 3176 3240 3188
rect 2179 3148 3240 3176
rect 2179 3145 2191 3148
rect 2133 3139 2191 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 4430 3136 4436 3188
rect 4488 3136 4494 3188
rect 5074 3136 5080 3188
rect 5132 3176 5138 3188
rect 5132 3148 5396 3176
rect 5132 3136 5138 3148
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3108 1823 3111
rect 3694 3108 3700 3120
rect 1811 3080 3700 3108
rect 1811 3077 1823 3080
rect 1765 3071 1823 3077
rect 3694 3068 3700 3080
rect 3752 3068 3758 3120
rect 4065 3111 4123 3117
rect 4065 3077 4077 3111
rect 4111 3108 4123 3111
rect 4448 3108 4476 3136
rect 4111 3080 4476 3108
rect 4111 3077 4123 3080
rect 4065 3071 4123 3077
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1360 3012 1961 3040
rect 1360 3000 1366 3012
rect 1949 3009 1961 3012
rect 1995 3009 2007 3043
rect 5368 3040 5396 3148
rect 5534 3136 5540 3188
rect 5592 3136 5598 3188
rect 7190 3136 7196 3188
rect 7248 3136 7254 3188
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 8113 3179 8171 3185
rect 8113 3176 8125 3179
rect 8076 3148 8125 3176
rect 8076 3136 8082 3148
rect 8113 3145 8125 3148
rect 8159 3145 8171 3179
rect 8113 3139 8171 3145
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 8628 3148 9260 3176
rect 8628 3136 8634 3148
rect 5552 3108 5580 3136
rect 5552 3080 5948 3108
rect 5920 3049 5948 3080
rect 5629 3043 5687 3049
rect 5629 3040 5641 3043
rect 1949 3003 2007 3009
rect 3786 2932 3792 2984
rect 3844 2932 3850 2984
rect 5184 2972 5212 3026
rect 5368 3012 5641 3040
rect 5629 3009 5641 3012
rect 5675 3009 5687 3043
rect 5629 3003 5687 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 7208 3040 7236 3136
rect 9122 3068 9128 3120
rect 9180 3068 9186 3120
rect 9232 3108 9260 3148
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 10229 3179 10287 3185
rect 9456 3148 9904 3176
rect 9456 3136 9462 3148
rect 9585 3111 9643 3117
rect 9585 3108 9597 3111
rect 9232 3080 9597 3108
rect 9585 3077 9597 3080
rect 9631 3077 9643 3111
rect 9585 3071 9643 3077
rect 9876 3049 9904 3148
rect 10229 3145 10241 3179
rect 10275 3176 10287 3179
rect 10410 3176 10416 3188
rect 10275 3148 10416 3176
rect 10275 3145 10287 3148
rect 10229 3139 10287 3145
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 10594 3136 10600 3188
rect 10652 3136 10658 3188
rect 10686 3136 10692 3188
rect 10744 3136 10750 3188
rect 11517 3179 11575 3185
rect 11517 3145 11529 3179
rect 11563 3145 11575 3179
rect 11517 3139 11575 3145
rect 10318 3068 10324 3120
rect 10376 3068 10382 3120
rect 7055 3012 7236 3040
rect 7469 3043 7527 3049
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 7469 3009 7481 3043
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 5350 2972 5356 2984
rect 5184 2944 5356 2972
rect 5350 2932 5356 2944
rect 5408 2932 5414 2984
rect 5442 2932 5448 2984
rect 5500 2972 5506 2984
rect 5537 2975 5595 2981
rect 5537 2972 5549 2975
rect 5500 2944 5549 2972
rect 5500 2932 5506 2944
rect 5537 2941 5549 2944
rect 5583 2941 5595 2975
rect 5828 2972 5856 3003
rect 6362 2972 6368 2984
rect 5828 2944 6368 2972
rect 5537 2935 5595 2941
rect 6362 2932 6368 2944
rect 6420 2972 6426 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6420 2944 6837 2972
rect 6420 2932 6426 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 7484 2972 7512 3003
rect 10502 3000 10508 3052
rect 10560 3000 10566 3052
rect 10612 3040 10640 3136
rect 10704 3108 10732 3136
rect 10704 3080 10824 3108
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10612 3012 10701 3040
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 10796 3040 10824 3080
rect 10962 3068 10968 3120
rect 11020 3108 11026 3120
rect 11532 3108 11560 3139
rect 14458 3136 14464 3188
rect 14516 3136 14522 3188
rect 15105 3179 15163 3185
rect 15105 3145 15117 3179
rect 15151 3176 15163 3179
rect 15930 3176 15936 3188
rect 15151 3148 15936 3176
rect 15151 3145 15163 3148
rect 15105 3139 15163 3145
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 16022 3136 16028 3188
rect 16080 3176 16086 3188
rect 16080 3148 16160 3176
rect 16080 3136 16086 3148
rect 12710 3108 12716 3120
rect 11020 3080 11560 3108
rect 12558 3080 12716 3108
rect 11020 3068 11026 3080
rect 12710 3068 12716 3080
rect 12768 3068 12774 3120
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 10796 3012 11161 3040
rect 10689 3003 10747 3009
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3040 13323 3043
rect 13446 3040 13452 3052
rect 13311 3012 13452 3040
rect 13311 3009 13323 3012
rect 13265 3003 13323 3009
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 14476 3040 14504 3136
rect 16132 3117 16160 3148
rect 16117 3111 16175 3117
rect 16117 3077 16129 3111
rect 16163 3077 16175 3111
rect 16117 3071 16175 3077
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 14476 3012 14933 3040
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 15654 3000 15660 3052
rect 15712 3000 15718 3052
rect 10520 2972 10548 3000
rect 7239 2944 7512 2972
rect 7576 2944 10548 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 6840 2904 6868 2935
rect 7576 2904 7604 2944
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12492 2944 13001 2972
rect 12492 2932 12498 2944
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 12989 2935 13047 2941
rect 6840 2876 7604 2904
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1489 2839 1547 2845
rect 1489 2836 1501 2839
rect 72 2808 1501 2836
rect 72 2796 78 2808
rect 1489 2805 1501 2808
rect 1535 2805 1547 2839
rect 1489 2799 1547 2805
rect 7282 2796 7288 2848
rect 7340 2796 7346 2848
rect 9122 2796 9128 2848
rect 9180 2836 9186 2848
rect 10410 2836 10416 2848
rect 9180 2808 10416 2836
rect 9180 2796 9186 2808
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 10870 2796 10876 2848
rect 10928 2796 10934 2848
rect 11330 2796 11336 2848
rect 11388 2796 11394 2848
rect 15746 2796 15752 2848
rect 15804 2796 15810 2848
rect 16393 2839 16451 2845
rect 16393 2805 16405 2839
rect 16439 2836 16451 2839
rect 16758 2836 16764 2848
rect 16439 2808 16764 2836
rect 16439 2805 16451 2808
rect 16393 2799 16451 2805
rect 16758 2796 16764 2808
rect 16816 2796 16822 2848
rect 944 2746 16836 2768
rect 944 2694 950 2746
rect 1002 2694 1014 2746
rect 1066 2694 1078 2746
rect 1130 2694 1142 2746
rect 1194 2694 1206 2746
rect 1258 2694 4950 2746
rect 5002 2694 5014 2746
rect 5066 2694 5078 2746
rect 5130 2694 5142 2746
rect 5194 2694 5206 2746
rect 5258 2694 8950 2746
rect 9002 2694 9014 2746
rect 9066 2694 9078 2746
rect 9130 2694 9142 2746
rect 9194 2694 9206 2746
rect 9258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 16836 2746
rect 944 2672 16836 2694
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 7892 2604 8125 2632
rect 7892 2592 7898 2604
rect 8113 2601 8125 2604
rect 8159 2601 8171 2635
rect 8113 2595 8171 2601
rect 11057 2635 11115 2641
rect 11057 2601 11069 2635
rect 11103 2632 11115 2635
rect 12434 2632 12440 2644
rect 11103 2604 12440 2632
rect 11103 2601 11115 2604
rect 11057 2595 11115 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 15930 2592 15936 2644
rect 15988 2592 15994 2644
rect 11146 2564 11152 2576
rect 8680 2536 11152 2564
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 6052 2468 6377 2496
rect 6052 2456 6058 2468
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6365 2459 6423 2465
rect 6641 2499 6699 2505
rect 6641 2465 6653 2499
rect 6687 2496 6699 2499
rect 7282 2496 7288 2508
rect 6687 2468 7288 2496
rect 6687 2465 6699 2468
rect 6641 2459 6699 2465
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2866 2428 2872 2440
rect 2179 2400 2872 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 4062 2428 4068 2440
rect 3559 2400 4068 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2428 6147 2431
rect 6270 2428 6276 2440
rect 6135 2400 6276 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 934 2320 940 2372
rect 992 2360 998 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 992 2332 1777 2360
rect 992 2320 998 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 4801 2363 4859 2369
rect 4801 2329 4813 2363
rect 4847 2360 4859 2363
rect 4847 2332 7052 2360
rect 4847 2329 4859 2332
rect 4801 2323 4859 2329
rect 3234 2252 3240 2304
rect 3292 2252 3298 2304
rect 4522 2252 4528 2304
rect 4580 2252 4586 2304
rect 5997 2295 6055 2301
rect 5997 2261 6009 2295
rect 6043 2292 6055 2295
rect 6454 2292 6460 2304
rect 6043 2264 6460 2292
rect 6043 2261 6055 2264
rect 5997 2255 6055 2261
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 7024 2292 7052 2332
rect 7098 2320 7104 2372
rect 7156 2320 7162 2372
rect 8680 2369 8708 2536
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 15948 2496 15976 2592
rect 15672 2468 15976 2496
rect 9858 2388 9864 2440
rect 9916 2388 9922 2440
rect 10870 2388 10876 2440
rect 10928 2388 10934 2440
rect 11330 2388 11336 2440
rect 11388 2388 11394 2440
rect 11422 2388 11428 2440
rect 11480 2428 11486 2440
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 11480 2400 11805 2428
rect 11480 2388 11486 2400
rect 11793 2397 11805 2400
rect 11839 2397 11851 2431
rect 11793 2391 11851 2397
rect 15102 2388 15108 2440
rect 15160 2388 15166 2440
rect 15672 2437 15700 2468
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 15746 2388 15752 2440
rect 15804 2428 15810 2440
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 15804 2400 16129 2428
rect 15804 2388 15810 2400
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2329 8723 2363
rect 16942 2360 16948 2372
rect 8665 2323 8723 2329
rect 15856 2332 16948 2360
rect 7374 2292 7380 2304
rect 7024 2264 7380 2292
rect 7374 2252 7380 2264
rect 7432 2252 7438 2304
rect 8386 2252 8392 2304
rect 8444 2252 8450 2304
rect 9950 2252 9956 2304
rect 10008 2252 10014 2304
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11885 2295 11943 2301
rect 11885 2292 11897 2295
rect 11664 2264 11897 2292
rect 11664 2252 11670 2264
rect 11885 2261 11897 2264
rect 11931 2261 11943 2295
rect 11885 2255 11943 2261
rect 14826 2252 14832 2304
rect 14884 2252 14890 2304
rect 15856 2301 15884 2332
rect 16942 2320 16948 2332
rect 17000 2320 17006 2372
rect 15841 2295 15899 2301
rect 15841 2261 15853 2295
rect 15887 2261 15899 2295
rect 15841 2255 15899 2261
rect 16390 2252 16396 2304
rect 16448 2252 16454 2304
rect 1104 2202 16836 2224
rect 1104 2150 1610 2202
rect 1662 2150 1674 2202
rect 1726 2150 1738 2202
rect 1790 2150 1802 2202
rect 1854 2150 1866 2202
rect 1918 2150 5610 2202
rect 5662 2150 5674 2202
rect 5726 2150 5738 2202
rect 5790 2150 5802 2202
rect 5854 2150 5866 2202
rect 5918 2150 9610 2202
rect 9662 2150 9674 2202
rect 9726 2150 9738 2202
rect 9790 2150 9802 2202
rect 9854 2150 9866 2202
rect 9918 2150 13610 2202
rect 13662 2150 13674 2202
rect 13726 2150 13738 2202
rect 13790 2150 13802 2202
rect 13854 2150 13866 2202
rect 13918 2150 16836 2202
rect 1104 2128 16836 2150
<< via1 >>
rect 950 15750 1002 15802
rect 1014 15750 1066 15802
rect 1078 15750 1130 15802
rect 1142 15750 1194 15802
rect 1206 15750 1258 15802
rect 4950 15750 5002 15802
rect 5014 15750 5066 15802
rect 5078 15750 5130 15802
rect 5142 15750 5194 15802
rect 5206 15750 5258 15802
rect 8950 15750 9002 15802
rect 9014 15750 9066 15802
rect 9078 15750 9130 15802
rect 9142 15750 9194 15802
rect 9206 15750 9258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 1492 15691 1544 15700
rect 1492 15657 1501 15691
rect 1501 15657 1535 15691
rect 1535 15657 1544 15691
rect 1492 15648 1544 15657
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 2780 15648 2832 15657
rect 5816 15648 5868 15700
rect 7840 15648 7892 15700
rect 9312 15648 9364 15700
rect 11060 15648 11112 15700
rect 12808 15648 12860 15700
rect 14372 15691 14424 15700
rect 14372 15657 14381 15691
rect 14381 15657 14415 15691
rect 14415 15657 14424 15691
rect 14372 15648 14424 15657
rect 16212 15691 16264 15700
rect 16212 15657 16221 15691
rect 16221 15657 16255 15691
rect 16255 15657 16264 15691
rect 16212 15648 16264 15657
rect 17408 15580 17460 15632
rect 664 15444 716 15496
rect 4528 15444 4580 15496
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 2320 15419 2372 15428
rect 2320 15385 2329 15419
rect 2329 15385 2363 15419
rect 2363 15385 2372 15419
rect 2320 15376 2372 15385
rect 3056 15419 3108 15428
rect 3056 15385 3065 15419
rect 3065 15385 3099 15419
rect 3099 15385 3108 15419
rect 3056 15376 3108 15385
rect 6276 15376 6328 15428
rect 6460 15419 6512 15428
rect 6460 15385 6469 15419
rect 6469 15385 6503 15419
rect 6503 15385 6512 15419
rect 6460 15376 6512 15385
rect 8208 15419 8260 15428
rect 8208 15385 8217 15419
rect 8217 15385 8251 15419
rect 8251 15385 8260 15419
rect 8208 15376 8260 15385
rect 11612 15419 11664 15428
rect 11612 15385 11621 15419
rect 11621 15385 11655 15419
rect 11655 15385 11664 15419
rect 11612 15376 11664 15385
rect 12808 15376 12860 15428
rect 14648 15419 14700 15428
rect 14648 15385 14657 15419
rect 14657 15385 14691 15419
rect 14691 15385 14700 15419
rect 14648 15376 14700 15385
rect 15292 15376 15344 15428
rect 15568 15419 15620 15428
rect 15568 15385 15577 15419
rect 15577 15385 15611 15419
rect 15611 15385 15620 15419
rect 15568 15376 15620 15385
rect 6000 15308 6052 15360
rect 1610 15206 1662 15258
rect 1674 15206 1726 15258
rect 1738 15206 1790 15258
rect 1802 15206 1854 15258
rect 1866 15206 1918 15258
rect 5610 15206 5662 15258
rect 5674 15206 5726 15258
rect 5738 15206 5790 15258
rect 5802 15206 5854 15258
rect 5866 15206 5918 15258
rect 9610 15206 9662 15258
rect 9674 15206 9726 15258
rect 9738 15206 9790 15258
rect 9802 15206 9854 15258
rect 9866 15206 9918 15258
rect 13610 15206 13662 15258
rect 13674 15206 13726 15258
rect 13738 15206 13790 15258
rect 13802 15206 13854 15258
rect 13866 15206 13918 15258
rect 2320 15104 2372 15156
rect 6460 15104 6512 15156
rect 8208 15104 8260 15156
rect 14648 15104 14700 15156
rect 16488 15104 16540 15156
rect 1400 15079 1452 15088
rect 1400 15045 1409 15079
rect 1409 15045 1443 15079
rect 1443 15045 1452 15079
rect 1400 15036 1452 15045
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 3148 15011 3200 15020
rect 3148 14977 3157 15011
rect 3157 14977 3191 15011
rect 3191 14977 3200 15011
rect 3148 14968 3200 14977
rect 6184 15011 6236 15020
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 8208 15011 8260 15020
rect 8208 14977 8217 15011
rect 8217 14977 8251 15011
rect 8251 14977 8260 15011
rect 8208 14968 8260 14977
rect 15292 14968 15344 15020
rect 16120 15011 16172 15020
rect 16120 14977 16129 15011
rect 16129 14977 16163 15011
rect 16163 14977 16172 15011
rect 16120 14968 16172 14977
rect 11612 14900 11664 14952
rect 950 14662 1002 14714
rect 1014 14662 1066 14714
rect 1078 14662 1130 14714
rect 1142 14662 1194 14714
rect 1206 14662 1258 14714
rect 4950 14662 5002 14714
rect 5014 14662 5066 14714
rect 5078 14662 5130 14714
rect 5142 14662 5194 14714
rect 5206 14662 5258 14714
rect 8950 14662 9002 14714
rect 9014 14662 9066 14714
rect 9078 14662 9130 14714
rect 9142 14662 9194 14714
rect 9206 14662 9258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 5080 14288 5132 14340
rect 15936 14288 15988 14340
rect 16948 14288 17000 14340
rect 2872 14220 2924 14272
rect 3792 14220 3844 14272
rect 5540 14220 5592 14272
rect 1610 14118 1662 14170
rect 1674 14118 1726 14170
rect 1738 14118 1790 14170
rect 1802 14118 1854 14170
rect 1866 14118 1918 14170
rect 5610 14118 5662 14170
rect 5674 14118 5726 14170
rect 5738 14118 5790 14170
rect 5802 14118 5854 14170
rect 5866 14118 5918 14170
rect 9610 14118 9662 14170
rect 9674 14118 9726 14170
rect 9738 14118 9790 14170
rect 9802 14118 9854 14170
rect 9866 14118 9918 14170
rect 13610 14118 13662 14170
rect 13674 14118 13726 14170
rect 13738 14118 13790 14170
rect 13802 14118 13854 14170
rect 13866 14118 13918 14170
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 1952 13880 2004 13932
rect 2872 13923 2924 13932
rect 2872 13889 2881 13923
rect 2881 13889 2915 13923
rect 2915 13889 2924 13923
rect 2872 13880 2924 13889
rect 3792 14016 3844 14068
rect 4528 14016 4580 14068
rect 5080 14016 5132 14068
rect 4160 13948 4212 14000
rect 4528 13880 4580 13932
rect 4804 13923 4856 13932
rect 4804 13889 4813 13923
rect 4813 13889 4847 13923
rect 4847 13889 4856 13923
rect 4804 13880 4856 13889
rect 4252 13812 4304 13864
rect 4620 13812 4672 13864
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 6736 13880 6788 13932
rect 6920 13880 6972 13932
rect 7472 13880 7524 13932
rect 6828 13812 6880 13864
rect 5356 13744 5408 13796
rect 1676 13719 1728 13728
rect 1676 13685 1685 13719
rect 1685 13685 1719 13719
rect 1719 13685 1728 13719
rect 1676 13676 1728 13685
rect 4712 13719 4764 13728
rect 4712 13685 4721 13719
rect 4721 13685 4755 13719
rect 4755 13685 4764 13719
rect 4712 13676 4764 13685
rect 7104 13719 7156 13728
rect 7104 13685 7113 13719
rect 7113 13685 7147 13719
rect 7147 13685 7156 13719
rect 7104 13676 7156 13685
rect 950 13574 1002 13626
rect 1014 13574 1066 13626
rect 1078 13574 1130 13626
rect 1142 13574 1194 13626
rect 1206 13574 1258 13626
rect 4950 13574 5002 13626
rect 5014 13574 5066 13626
rect 5078 13574 5130 13626
rect 5142 13574 5194 13626
rect 5206 13574 5258 13626
rect 8950 13574 9002 13626
rect 9014 13574 9066 13626
rect 9078 13574 9130 13626
rect 9142 13574 9194 13626
rect 9206 13574 9258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 3056 13472 3108 13524
rect 3332 13472 3384 13524
rect 4620 13515 4672 13524
rect 4620 13481 4629 13515
rect 4629 13481 4663 13515
rect 4663 13481 4672 13515
rect 4620 13472 4672 13481
rect 4804 13404 4856 13456
rect 2964 13336 3016 13388
rect 4160 13379 4212 13388
rect 4160 13345 4169 13379
rect 4169 13345 4203 13379
rect 4203 13345 4212 13379
rect 4160 13336 4212 13345
rect 1676 13243 1728 13252
rect 1676 13209 1685 13243
rect 1685 13209 1719 13243
rect 1719 13209 1728 13243
rect 1676 13200 1728 13209
rect 4068 13200 4120 13252
rect 5356 13404 5408 13456
rect 5540 13404 5592 13456
rect 6828 13336 6880 13388
rect 7104 13336 7156 13388
rect 7380 13336 7432 13388
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 2596 13132 2648 13184
rect 7196 13311 7248 13320
rect 7196 13277 7205 13311
rect 7205 13277 7239 13311
rect 7239 13277 7248 13311
rect 7196 13268 7248 13277
rect 9312 13472 9364 13524
rect 12808 13472 12860 13524
rect 10232 13404 10284 13456
rect 4896 13132 4948 13184
rect 6920 13132 6972 13184
rect 7012 13175 7064 13184
rect 7012 13141 7021 13175
rect 7021 13141 7055 13175
rect 7055 13141 7064 13175
rect 7012 13132 7064 13141
rect 7288 13132 7340 13184
rect 8668 13200 8720 13252
rect 10876 13268 10928 13320
rect 11428 13243 11480 13252
rect 11428 13209 11437 13243
rect 11437 13209 11471 13243
rect 11471 13209 11480 13243
rect 11428 13200 11480 13209
rect 12716 13200 12768 13252
rect 16120 13243 16172 13252
rect 16120 13209 16129 13243
rect 16129 13209 16163 13243
rect 16163 13209 16172 13243
rect 16120 13200 16172 13209
rect 14004 13132 14056 13184
rect 16948 13132 17000 13184
rect 1610 13030 1662 13082
rect 1674 13030 1726 13082
rect 1738 13030 1790 13082
rect 1802 13030 1854 13082
rect 1866 13030 1918 13082
rect 5610 13030 5662 13082
rect 5674 13030 5726 13082
rect 5738 13030 5790 13082
rect 5802 13030 5854 13082
rect 5866 13030 5918 13082
rect 9610 13030 9662 13082
rect 9674 13030 9726 13082
rect 9738 13030 9790 13082
rect 9802 13030 9854 13082
rect 9866 13030 9918 13082
rect 13610 13030 13662 13082
rect 13674 13030 13726 13082
rect 13738 13030 13790 13082
rect 13802 13030 13854 13082
rect 13866 13030 13918 13082
rect 1952 12971 2004 12980
rect 1952 12937 1961 12971
rect 1961 12937 1995 12971
rect 1995 12937 2004 12971
rect 1952 12928 2004 12937
rect 2596 12928 2648 12980
rect 2872 12928 2924 12980
rect 4896 12928 4948 12980
rect 4068 12860 4120 12912
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 2964 12792 3016 12844
rect 4344 12792 4396 12844
rect 2872 12767 2924 12776
rect 2872 12733 2881 12767
rect 2881 12733 2915 12767
rect 2915 12733 2924 12767
rect 2872 12724 2924 12733
rect 3240 12724 3292 12776
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 7196 12928 7248 12980
rect 7288 12971 7340 12980
rect 7288 12937 7297 12971
rect 7297 12937 7331 12971
rect 7331 12937 7340 12971
rect 7288 12928 7340 12937
rect 7380 12928 7432 12980
rect 8668 12928 8720 12980
rect 5080 12792 5132 12844
rect 5540 12792 5592 12844
rect 4252 12656 4304 12708
rect 5356 12656 5408 12708
rect 10600 12903 10652 12912
rect 10600 12869 10609 12903
rect 10609 12869 10643 12903
rect 10643 12869 10652 12903
rect 10600 12860 10652 12869
rect 11428 12928 11480 12980
rect 15292 12971 15344 12980
rect 15292 12937 15301 12971
rect 15301 12937 15335 12971
rect 15335 12937 15344 12971
rect 15292 12928 15344 12937
rect 15568 12928 15620 12980
rect 15936 12971 15988 12980
rect 15936 12937 15945 12971
rect 15945 12937 15979 12971
rect 15979 12937 15988 12971
rect 15936 12928 15988 12937
rect 16120 12971 16172 12980
rect 16120 12937 16129 12971
rect 16129 12937 16163 12971
rect 16163 12937 16172 12971
rect 16120 12928 16172 12937
rect 8576 12835 8628 12844
rect 8576 12801 8585 12835
rect 8585 12801 8619 12835
rect 8619 12801 8628 12835
rect 8576 12792 8628 12801
rect 9312 12792 9364 12844
rect 9496 12792 9548 12844
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 6920 12724 6972 12776
rect 7288 12724 7340 12776
rect 11796 12724 11848 12776
rect 15108 12835 15160 12844
rect 15108 12801 15117 12835
rect 15117 12801 15151 12835
rect 15151 12801 15160 12835
rect 15108 12792 15160 12801
rect 15752 12835 15804 12844
rect 15752 12801 15761 12835
rect 15761 12801 15795 12835
rect 15795 12801 15804 12835
rect 15752 12792 15804 12801
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 2504 12588 2556 12640
rect 5080 12588 5132 12640
rect 5540 12588 5592 12640
rect 6276 12588 6328 12640
rect 9128 12631 9180 12640
rect 9128 12597 9137 12631
rect 9137 12597 9171 12631
rect 9171 12597 9180 12631
rect 9128 12588 9180 12597
rect 9404 12588 9456 12640
rect 11796 12588 11848 12640
rect 13820 12588 13872 12640
rect 950 12486 1002 12538
rect 1014 12486 1066 12538
rect 1078 12486 1130 12538
rect 1142 12486 1194 12538
rect 1206 12486 1258 12538
rect 4950 12486 5002 12538
rect 5014 12486 5066 12538
rect 5078 12486 5130 12538
rect 5142 12486 5194 12538
rect 5206 12486 5258 12538
rect 8950 12486 9002 12538
rect 9014 12486 9066 12538
rect 9078 12486 9130 12538
rect 9142 12486 9194 12538
rect 9206 12486 9258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 2136 12384 2188 12436
rect 7288 12384 7340 12436
rect 8576 12427 8628 12436
rect 8576 12393 8585 12427
rect 8585 12393 8619 12427
rect 8619 12393 8628 12427
rect 8576 12384 8628 12393
rect 11704 12384 11756 12436
rect 2872 12316 2924 12368
rect 7472 12316 7524 12368
rect 12256 12316 12308 12368
rect 14188 12384 14240 12436
rect 12532 12359 12584 12368
rect 12532 12325 12541 12359
rect 12541 12325 12575 12359
rect 12575 12325 12584 12359
rect 12532 12316 12584 12325
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 3332 12223 3384 12232
rect 3332 12189 3341 12223
rect 3341 12189 3375 12223
rect 3375 12189 3384 12223
rect 3332 12180 3384 12189
rect 5540 12291 5592 12300
rect 5540 12257 5549 12291
rect 5549 12257 5583 12291
rect 5583 12257 5592 12291
rect 5540 12248 5592 12257
rect 3884 12180 3936 12232
rect 4068 12180 4120 12232
rect 10876 12248 10928 12300
rect 11336 12248 11388 12300
rect 9312 12180 9364 12232
rect 10968 12180 11020 12232
rect 1952 12044 2004 12096
rect 2320 12044 2372 12096
rect 3608 12044 3660 12096
rect 5448 12044 5500 12096
rect 10140 12112 10192 12164
rect 10416 12087 10468 12096
rect 10416 12053 10425 12087
rect 10425 12053 10459 12087
rect 10459 12053 10468 12087
rect 10416 12044 10468 12053
rect 12256 12223 12308 12232
rect 12256 12189 12265 12223
rect 12265 12189 12299 12223
rect 12299 12189 12308 12223
rect 12256 12180 12308 12189
rect 12808 12180 12860 12232
rect 12624 12112 12676 12164
rect 13820 12223 13872 12232
rect 13820 12189 13829 12223
rect 13829 12189 13863 12223
rect 13863 12189 13872 12223
rect 13820 12180 13872 12189
rect 14280 12112 14332 12164
rect 15384 12112 15436 12164
rect 13452 12044 13504 12096
rect 15016 12044 15068 12096
rect 1610 11942 1662 11994
rect 1674 11942 1726 11994
rect 1738 11942 1790 11994
rect 1802 11942 1854 11994
rect 1866 11942 1918 11994
rect 5610 11942 5662 11994
rect 5674 11942 5726 11994
rect 5738 11942 5790 11994
rect 5802 11942 5854 11994
rect 5866 11942 5918 11994
rect 9610 11942 9662 11994
rect 9674 11942 9726 11994
rect 9738 11942 9790 11994
rect 9802 11942 9854 11994
rect 9866 11942 9918 11994
rect 13610 11942 13662 11994
rect 13674 11942 13726 11994
rect 13738 11942 13790 11994
rect 13802 11942 13854 11994
rect 13866 11942 13918 11994
rect 4528 11840 4580 11892
rect 3240 11747 3292 11756
rect 3240 11713 3249 11747
rect 3249 11713 3283 11747
rect 3283 11713 3292 11747
rect 3240 11704 3292 11713
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 3608 11636 3660 11645
rect 4068 11636 4120 11688
rect 4160 11636 4212 11688
rect 5448 11772 5500 11824
rect 7472 11772 7524 11824
rect 9496 11772 9548 11824
rect 10048 11772 10100 11824
rect 7196 11747 7248 11756
rect 7196 11713 7205 11747
rect 7205 11713 7239 11747
rect 7239 11713 7248 11747
rect 7196 11704 7248 11713
rect 12532 11840 12584 11892
rect 14280 11840 14332 11892
rect 15108 11883 15160 11892
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 14096 11772 14148 11824
rect 11336 11636 11388 11688
rect 11428 11636 11480 11688
rect 12256 11636 12308 11688
rect 6736 11568 6788 11620
rect 6828 11611 6880 11620
rect 6828 11577 6837 11611
rect 6837 11577 6871 11611
rect 6871 11577 6880 11611
rect 6828 11568 6880 11577
rect 12716 11568 12768 11620
rect 13452 11636 13504 11688
rect 15016 11704 15068 11756
rect 14832 11636 14884 11688
rect 3240 11500 3292 11552
rect 8484 11543 8536 11552
rect 8484 11509 8493 11543
rect 8493 11509 8527 11543
rect 8527 11509 8536 11543
rect 8484 11500 8536 11509
rect 13360 11500 13412 11552
rect 14188 11500 14240 11552
rect 950 11398 1002 11450
rect 1014 11398 1066 11450
rect 1078 11398 1130 11450
rect 1142 11398 1194 11450
rect 1206 11398 1258 11450
rect 4950 11398 5002 11450
rect 5014 11398 5066 11450
rect 5078 11398 5130 11450
rect 5142 11398 5194 11450
rect 5206 11398 5258 11450
rect 8950 11398 9002 11450
rect 9014 11398 9066 11450
rect 9078 11398 9130 11450
rect 9142 11398 9194 11450
rect 9206 11398 9258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 2872 11296 2924 11348
rect 3148 11296 3200 11348
rect 3884 11339 3936 11348
rect 3884 11305 3893 11339
rect 3893 11305 3927 11339
rect 3927 11305 3936 11339
rect 3884 11296 3936 11305
rect 6736 11296 6788 11348
rect 8484 11296 8536 11348
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 2780 11135 2832 11144
rect 2780 11101 2789 11135
rect 2789 11101 2823 11135
rect 2823 11101 2832 11135
rect 2780 11092 2832 11101
rect 2964 11024 3016 11076
rect 6368 11228 6420 11280
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 4528 11203 4580 11212
rect 4528 11169 4537 11203
rect 4537 11169 4571 11203
rect 4571 11169 4580 11203
rect 4528 11160 4580 11169
rect 10416 11296 10468 11348
rect 10600 11296 10652 11348
rect 12624 11296 12676 11348
rect 10324 11228 10376 11280
rect 4068 11092 4120 11144
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 3240 11067 3292 11076
rect 3240 11033 3249 11067
rect 3249 11033 3283 11067
rect 3283 11033 3292 11067
rect 3240 11024 3292 11033
rect 3424 11024 3476 11076
rect 5080 11067 5132 11076
rect 5080 11033 5089 11067
rect 5089 11033 5123 11067
rect 5123 11033 5132 11067
rect 5080 11024 5132 11033
rect 6644 11024 6696 11076
rect 1492 10956 1544 11008
rect 4252 10999 4304 11008
rect 4252 10965 4261 10999
rect 4261 10965 4295 10999
rect 4295 10965 4304 10999
rect 4252 10956 4304 10965
rect 8484 11024 8536 11076
rect 9404 11092 9456 11144
rect 11336 11160 11388 11212
rect 14096 11339 14148 11348
rect 14096 11305 14105 11339
rect 14105 11305 14139 11339
rect 14139 11305 14148 11339
rect 14096 11296 14148 11305
rect 16488 11160 16540 11212
rect 14832 11092 14884 11144
rect 7012 10956 7064 11008
rect 11244 11067 11296 11076
rect 11244 11033 11253 11067
rect 11253 11033 11287 11067
rect 11287 11033 11296 11067
rect 11244 11024 11296 11033
rect 15108 11024 15160 11076
rect 9956 10999 10008 11008
rect 9956 10965 9965 10999
rect 9965 10965 9999 10999
rect 9999 10965 10008 10999
rect 9956 10956 10008 10965
rect 10600 10956 10652 11008
rect 11428 10956 11480 11008
rect 12072 10956 12124 11008
rect 12532 10956 12584 11008
rect 12808 10999 12860 11008
rect 12808 10965 12817 10999
rect 12817 10965 12851 10999
rect 12851 10965 12860 10999
rect 12808 10956 12860 10965
rect 12900 10956 12952 11008
rect 1610 10854 1662 10906
rect 1674 10854 1726 10906
rect 1738 10854 1790 10906
rect 1802 10854 1854 10906
rect 1866 10854 1918 10906
rect 5610 10854 5662 10906
rect 5674 10854 5726 10906
rect 5738 10854 5790 10906
rect 5802 10854 5854 10906
rect 5866 10854 5918 10906
rect 9610 10854 9662 10906
rect 9674 10854 9726 10906
rect 9738 10854 9790 10906
rect 9802 10854 9854 10906
rect 9866 10854 9918 10906
rect 13610 10854 13662 10906
rect 13674 10854 13726 10906
rect 13738 10854 13790 10906
rect 13802 10854 13854 10906
rect 13866 10854 13918 10906
rect 1492 10752 1544 10804
rect 4344 10752 4396 10804
rect 5356 10752 5408 10804
rect 9312 10752 9364 10804
rect 3332 10616 3384 10668
rect 4252 10616 4304 10668
rect 8576 10684 8628 10736
rect 9404 10684 9456 10736
rect 10416 10727 10468 10736
rect 10416 10693 10438 10727
rect 10438 10693 10468 10727
rect 11244 10752 11296 10804
rect 12072 10752 12124 10804
rect 12808 10752 12860 10804
rect 14004 10752 14056 10804
rect 15108 10795 15160 10804
rect 15108 10761 15117 10795
rect 15117 10761 15151 10795
rect 15151 10761 15160 10795
rect 15108 10752 15160 10761
rect 10416 10684 10468 10693
rect 6368 10616 6420 10668
rect 6920 10616 6972 10668
rect 8300 10616 8352 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 4804 10548 4856 10600
rect 6828 10548 6880 10600
rect 7012 10591 7064 10600
rect 7012 10557 7021 10591
rect 7021 10557 7055 10591
rect 7055 10557 7064 10591
rect 7012 10548 7064 10557
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 9956 10616 10008 10668
rect 11612 10684 11664 10736
rect 12256 10684 12308 10736
rect 5080 10480 5132 10532
rect 2964 10412 3016 10464
rect 4712 10455 4764 10464
rect 4712 10421 4721 10455
rect 4721 10421 4755 10455
rect 4755 10421 4764 10455
rect 4712 10412 4764 10421
rect 5356 10480 5408 10532
rect 10048 10480 10100 10532
rect 10324 10548 10376 10600
rect 11704 10548 11756 10600
rect 8852 10455 8904 10464
rect 8852 10421 8861 10455
rect 8861 10421 8895 10455
rect 8895 10421 8904 10455
rect 8852 10412 8904 10421
rect 11520 10480 11572 10532
rect 11612 10480 11664 10532
rect 12440 10616 12492 10668
rect 13360 10727 13412 10736
rect 13360 10693 13369 10727
rect 13369 10693 13403 10727
rect 13403 10693 13412 10727
rect 13360 10684 13412 10693
rect 15384 10684 15436 10736
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 12716 10523 12768 10532
rect 12716 10489 12725 10523
rect 12725 10489 12759 10523
rect 12759 10489 12768 10523
rect 12716 10480 12768 10489
rect 10784 10455 10836 10464
rect 10784 10421 10793 10455
rect 10793 10421 10827 10455
rect 10827 10421 10836 10455
rect 10784 10412 10836 10421
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 12624 10412 12676 10464
rect 13544 10412 13596 10464
rect 14832 10455 14884 10464
rect 14832 10421 14841 10455
rect 14841 10421 14875 10455
rect 14875 10421 14884 10455
rect 14832 10412 14884 10421
rect 950 10310 1002 10362
rect 1014 10310 1066 10362
rect 1078 10310 1130 10362
rect 1142 10310 1194 10362
rect 1206 10310 1258 10362
rect 4950 10310 5002 10362
rect 5014 10310 5066 10362
rect 5078 10310 5130 10362
rect 5142 10310 5194 10362
rect 5206 10310 5258 10362
rect 8950 10310 9002 10362
rect 9014 10310 9066 10362
rect 9078 10310 9130 10362
rect 9142 10310 9194 10362
rect 9206 10310 9258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 940 10208 992 10260
rect 6276 10208 6328 10260
rect 6920 10208 6972 10260
rect 8852 10208 8904 10260
rect 9404 10208 9456 10260
rect 10140 10208 10192 10260
rect 10784 10208 10836 10260
rect 11520 10208 11572 10260
rect 14832 10208 14884 10260
rect 14924 10251 14976 10260
rect 14924 10217 14933 10251
rect 14933 10217 14967 10251
rect 14967 10217 14976 10251
rect 14924 10208 14976 10217
rect 4804 10072 4856 10124
rect 6920 10115 6972 10124
rect 6920 10081 6929 10115
rect 6929 10081 6963 10115
rect 6963 10081 6972 10115
rect 6920 10072 6972 10081
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 5356 10004 5408 10056
rect 6828 10004 6880 10056
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 10324 10072 10376 10124
rect 10600 10004 10652 10056
rect 10324 9936 10376 9988
rect 7656 9868 7708 9920
rect 11244 9868 11296 9920
rect 11336 9868 11388 9920
rect 11520 9868 11572 9920
rect 12808 10004 12860 10056
rect 15384 10004 15436 10056
rect 14556 9979 14608 9988
rect 14556 9945 14565 9979
rect 14565 9945 14599 9979
rect 14599 9945 14608 9979
rect 14556 9936 14608 9945
rect 13452 9868 13504 9920
rect 1610 9766 1662 9818
rect 1674 9766 1726 9818
rect 1738 9766 1790 9818
rect 1802 9766 1854 9818
rect 1866 9766 1918 9818
rect 5610 9766 5662 9818
rect 5674 9766 5726 9818
rect 5738 9766 5790 9818
rect 5802 9766 5854 9818
rect 5866 9766 5918 9818
rect 9610 9766 9662 9818
rect 9674 9766 9726 9818
rect 9738 9766 9790 9818
rect 9802 9766 9854 9818
rect 9866 9766 9918 9818
rect 13610 9766 13662 9818
rect 13674 9766 13726 9818
rect 13738 9766 13790 9818
rect 13802 9766 13854 9818
rect 13866 9766 13918 9818
rect 6920 9664 6972 9716
rect 11244 9664 11296 9716
rect 2136 9596 2188 9648
rect 1400 9528 1452 9580
rect 4068 9528 4120 9580
rect 2044 9503 2096 9512
rect 2044 9469 2053 9503
rect 2053 9469 2087 9503
rect 2087 9469 2096 9503
rect 2044 9460 2096 9469
rect 2136 9460 2188 9512
rect 3332 9460 3384 9512
rect 4620 9528 4672 9580
rect 5448 9528 5500 9580
rect 6276 9528 6328 9580
rect 8852 9596 8904 9648
rect 9404 9596 9456 9648
rect 13268 9596 13320 9648
rect 13636 9596 13688 9648
rect 15384 9596 15436 9648
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 6828 9528 6880 9580
rect 7380 9528 7432 9580
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 2688 9324 2740 9376
rect 6368 9392 6420 9444
rect 6552 9392 6604 9444
rect 3516 9367 3568 9376
rect 3516 9333 3525 9367
rect 3525 9333 3559 9367
rect 3559 9333 3568 9367
rect 3516 9324 3568 9333
rect 8300 9392 8352 9444
rect 10048 9392 10100 9444
rect 6920 9324 6972 9376
rect 7564 9324 7616 9376
rect 10232 9324 10284 9376
rect 12808 9460 12860 9512
rect 13360 9528 13412 9580
rect 13544 9460 13596 9512
rect 13636 9503 13688 9512
rect 13636 9469 13645 9503
rect 13645 9469 13679 9503
rect 13679 9469 13688 9503
rect 13636 9460 13688 9469
rect 13820 9503 13872 9512
rect 13820 9469 13829 9503
rect 13829 9469 13863 9503
rect 13863 9469 13872 9503
rect 13820 9460 13872 9469
rect 11796 9324 11848 9376
rect 12256 9324 12308 9376
rect 12808 9324 12860 9376
rect 13728 9324 13780 9376
rect 14372 9503 14424 9512
rect 14372 9469 14381 9503
rect 14381 9469 14415 9503
rect 14415 9469 14424 9503
rect 14372 9460 14424 9469
rect 14556 9324 14608 9376
rect 16120 9324 16172 9376
rect 950 9222 1002 9274
rect 1014 9222 1066 9274
rect 1078 9222 1130 9274
rect 1142 9222 1194 9274
rect 1206 9222 1258 9274
rect 4950 9222 5002 9274
rect 5014 9222 5066 9274
rect 5078 9222 5130 9274
rect 5142 9222 5194 9274
rect 5206 9222 5258 9274
rect 8950 9222 9002 9274
rect 9014 9222 9066 9274
rect 9078 9222 9130 9274
rect 9142 9222 9194 9274
rect 9206 9222 9258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 2044 9120 2096 9172
rect 3516 8984 3568 9036
rect 3884 8984 3936 9036
rect 1952 8916 2004 8968
rect 940 8848 992 8900
rect 4620 8916 4672 8968
rect 5448 9095 5500 9104
rect 5448 9061 5457 9095
rect 5457 9061 5491 9095
rect 5491 9061 5500 9095
rect 5448 9052 5500 9061
rect 6000 9052 6052 9104
rect 7656 9120 7708 9172
rect 9496 9120 9548 9172
rect 4436 8780 4488 8832
rect 6368 8916 6420 8968
rect 6552 9027 6604 9036
rect 6552 8993 6561 9027
rect 6561 8993 6595 9027
rect 6595 8993 6604 9027
rect 6552 8984 6604 8993
rect 9220 9095 9272 9104
rect 9220 9061 9229 9095
rect 9229 9061 9263 9095
rect 9263 9061 9272 9095
rect 9220 9052 9272 9061
rect 12256 9052 12308 9104
rect 7012 8984 7064 9036
rect 7472 8984 7524 9036
rect 8760 8984 8812 9036
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 10048 8984 10100 9036
rect 10140 8984 10192 9036
rect 11520 9027 11572 9036
rect 11520 8993 11529 9027
rect 11529 8993 11563 9027
rect 11563 8993 11572 9027
rect 11520 8984 11572 8993
rect 11612 8984 11664 9036
rect 9404 8916 9456 8968
rect 9772 8916 9824 8968
rect 11336 8916 11388 8968
rect 11704 8959 11756 8968
rect 11704 8925 11713 8959
rect 11713 8925 11747 8959
rect 11747 8925 11756 8959
rect 11704 8916 11756 8925
rect 11888 8959 11940 8968
rect 11888 8925 11897 8959
rect 11897 8925 11931 8959
rect 11931 8925 11940 8959
rect 11888 8916 11940 8925
rect 12624 9120 12676 9172
rect 14004 9120 14056 9172
rect 14372 9120 14424 9172
rect 12532 8984 12584 9036
rect 15568 8984 15620 9036
rect 13728 8916 13780 8968
rect 16120 8959 16172 8968
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 16120 8916 16172 8925
rect 7288 8780 7340 8832
rect 10876 8848 10928 8900
rect 11428 8848 11480 8900
rect 16764 8848 16816 8900
rect 10140 8780 10192 8832
rect 11520 8780 11572 8832
rect 12532 8823 12584 8832
rect 12532 8789 12559 8823
rect 12559 8789 12584 8823
rect 12532 8780 12584 8789
rect 1610 8678 1662 8730
rect 1674 8678 1726 8730
rect 1738 8678 1790 8730
rect 1802 8678 1854 8730
rect 1866 8678 1918 8730
rect 5610 8678 5662 8730
rect 5674 8678 5726 8730
rect 5738 8678 5790 8730
rect 5802 8678 5854 8730
rect 5866 8678 5918 8730
rect 9610 8678 9662 8730
rect 9674 8678 9726 8730
rect 9738 8678 9790 8730
rect 9802 8678 9854 8730
rect 9866 8678 9918 8730
rect 13610 8678 13662 8730
rect 13674 8678 13726 8730
rect 13738 8678 13790 8730
rect 13802 8678 13854 8730
rect 13866 8678 13918 8730
rect 3884 8576 3936 8628
rect 4160 8508 4212 8560
rect 2688 8440 2740 8492
rect 4528 8483 4580 8492
rect 4528 8449 4537 8483
rect 4537 8449 4571 8483
rect 4571 8449 4580 8483
rect 4528 8440 4580 8449
rect 4804 8440 4856 8492
rect 6000 8576 6052 8628
rect 8944 8619 8996 8628
rect 5356 8508 5408 8560
rect 5540 8508 5592 8560
rect 8944 8585 8953 8619
rect 8953 8585 8987 8619
rect 8987 8585 8996 8619
rect 8944 8576 8996 8585
rect 9220 8576 9272 8628
rect 11336 8576 11388 8628
rect 13360 8576 13412 8628
rect 14004 8576 14056 8628
rect 14648 8576 14700 8628
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 2320 8372 2372 8424
rect 6644 8372 6696 8424
rect 8760 8440 8812 8492
rect 8944 8440 8996 8492
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 10140 8508 10192 8560
rect 11428 8508 11480 8560
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 9036 8372 9088 8424
rect 10968 8440 11020 8492
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 15752 8576 15804 8628
rect 16120 8440 16172 8492
rect 10416 8372 10468 8424
rect 13636 8415 13688 8424
rect 13636 8381 13645 8415
rect 13645 8381 13679 8415
rect 13679 8381 13688 8415
rect 13636 8372 13688 8381
rect 13728 8372 13780 8424
rect 4252 8236 4304 8288
rect 5356 8236 5408 8288
rect 8668 8236 8720 8288
rect 9312 8347 9364 8356
rect 9312 8313 9321 8347
rect 9321 8313 9355 8347
rect 9355 8313 9364 8347
rect 9312 8304 9364 8313
rect 10876 8304 10928 8356
rect 11060 8236 11112 8288
rect 11704 8236 11756 8288
rect 14188 8236 14240 8288
rect 15200 8279 15252 8288
rect 15200 8245 15209 8279
rect 15209 8245 15243 8279
rect 15243 8245 15252 8279
rect 15200 8236 15252 8245
rect 950 8134 1002 8186
rect 1014 8134 1066 8186
rect 1078 8134 1130 8186
rect 1142 8134 1194 8186
rect 1206 8134 1258 8186
rect 4950 8134 5002 8186
rect 5014 8134 5066 8186
rect 5078 8134 5130 8186
rect 5142 8134 5194 8186
rect 5206 8134 5258 8186
rect 8950 8134 9002 8186
rect 9014 8134 9066 8186
rect 9078 8134 9130 8186
rect 9142 8134 9194 8186
rect 9206 8134 9258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 4160 8032 4212 8084
rect 4804 8032 4856 8084
rect 5356 8032 5408 8084
rect 6644 8032 6696 8084
rect 11428 8032 11480 8084
rect 11060 7964 11112 8016
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 4436 7896 4488 7948
rect 5448 7896 5500 7948
rect 7288 7896 7340 7948
rect 7380 7896 7432 7948
rect 3884 7871 3936 7880
rect 3884 7837 3893 7871
rect 3893 7837 3927 7871
rect 3927 7837 3936 7871
rect 3884 7828 3936 7837
rect 4160 7828 4212 7880
rect 6000 7828 6052 7880
rect 7564 7871 7616 7880
rect 7564 7837 7573 7871
rect 7573 7837 7607 7871
rect 7607 7837 7616 7871
rect 7564 7828 7616 7837
rect 9956 7828 10008 7880
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 10140 7828 10192 7880
rect 10416 7828 10468 7880
rect 11980 7964 12032 8016
rect 12532 8032 12584 8084
rect 13452 8032 13504 8084
rect 13636 8032 13688 8084
rect 15200 8032 15252 8084
rect 12440 7896 12492 7948
rect 2044 7692 2096 7744
rect 4252 7692 4304 7744
rect 4896 7692 4948 7744
rect 6092 7692 6144 7744
rect 6368 7735 6420 7744
rect 6368 7701 6377 7735
rect 6377 7701 6411 7735
rect 6411 7701 6420 7735
rect 6368 7692 6420 7701
rect 9312 7692 9364 7744
rect 11520 7871 11572 7880
rect 11520 7837 11543 7871
rect 11543 7837 11572 7871
rect 11520 7828 11572 7837
rect 14648 7939 14700 7948
rect 14648 7905 14657 7939
rect 14657 7905 14691 7939
rect 14691 7905 14700 7939
rect 14648 7896 14700 7905
rect 11888 7803 11940 7812
rect 11888 7769 11897 7803
rect 11897 7769 11931 7803
rect 11931 7769 11940 7803
rect 11888 7760 11940 7769
rect 13360 7828 13412 7880
rect 11704 7735 11756 7744
rect 11704 7701 11713 7735
rect 11713 7701 11747 7735
rect 11747 7701 11756 7735
rect 11704 7692 11756 7701
rect 11796 7692 11848 7744
rect 15568 7828 15620 7880
rect 12624 7692 12676 7744
rect 12808 7692 12860 7744
rect 13360 7692 13412 7744
rect 14096 7692 14148 7744
rect 14832 7692 14884 7744
rect 16764 7692 16816 7744
rect 1610 7590 1662 7642
rect 1674 7590 1726 7642
rect 1738 7590 1790 7642
rect 1802 7590 1854 7642
rect 1866 7590 1918 7642
rect 5610 7590 5662 7642
rect 5674 7590 5726 7642
rect 5738 7590 5790 7642
rect 5802 7590 5854 7642
rect 5866 7590 5918 7642
rect 9610 7590 9662 7642
rect 9674 7590 9726 7642
rect 9738 7590 9790 7642
rect 9802 7590 9854 7642
rect 9866 7590 9918 7642
rect 13610 7590 13662 7642
rect 13674 7590 13726 7642
rect 13738 7590 13790 7642
rect 13802 7590 13854 7642
rect 13866 7590 13918 7642
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 4160 7488 4212 7540
rect 4252 7488 4304 7540
rect 2320 7420 2372 7472
rect 3884 7463 3936 7472
rect 3884 7429 3902 7463
rect 3902 7429 3936 7463
rect 3884 7420 3936 7429
rect 3148 7352 3200 7404
rect 7564 7488 7616 7540
rect 11704 7488 11756 7540
rect 9220 7420 9272 7472
rect 10692 7420 10744 7472
rect 11980 7488 12032 7540
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 5356 7352 5408 7404
rect 3976 7284 4028 7336
rect 4160 7216 4212 7268
rect 4436 7284 4488 7336
rect 6092 7352 6144 7404
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7564 7352 7616 7404
rect 9496 7352 9548 7404
rect 10048 7352 10100 7404
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 13452 7420 13504 7472
rect 11152 7284 11204 7336
rect 2320 7191 2372 7200
rect 2320 7157 2329 7191
rect 2329 7157 2363 7191
rect 2363 7157 2372 7191
rect 2320 7148 2372 7157
rect 2872 7148 2924 7200
rect 3332 7148 3384 7200
rect 5540 7148 5592 7200
rect 7564 7148 7616 7200
rect 10968 7148 11020 7200
rect 11244 7259 11296 7268
rect 11244 7225 11253 7259
rect 11253 7225 11287 7259
rect 11287 7225 11296 7259
rect 11888 7284 11940 7336
rect 12440 7284 12492 7336
rect 14004 7284 14056 7336
rect 14832 7284 14884 7336
rect 11244 7216 11296 7225
rect 12532 7148 12584 7200
rect 12808 7148 12860 7200
rect 16120 7148 16172 7200
rect 950 7046 1002 7098
rect 1014 7046 1066 7098
rect 1078 7046 1130 7098
rect 1142 7046 1194 7098
rect 1206 7046 1258 7098
rect 4950 7046 5002 7098
rect 5014 7046 5066 7098
rect 5078 7046 5130 7098
rect 5142 7046 5194 7098
rect 5206 7046 5258 7098
rect 8950 7046 9002 7098
rect 9014 7046 9066 7098
rect 9078 7046 9130 7098
rect 9142 7046 9194 7098
rect 9206 7046 9258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 3148 6987 3200 6996
rect 3148 6953 3157 6987
rect 3157 6953 3191 6987
rect 3191 6953 3200 6987
rect 3148 6944 3200 6953
rect 3884 6944 3936 6996
rect 2412 6808 2464 6860
rect 4160 6851 4212 6860
rect 4160 6817 4169 6851
rect 4169 6817 4203 6851
rect 4203 6817 4212 6851
rect 4160 6808 4212 6817
rect 6276 6944 6328 6996
rect 6368 6944 6420 6996
rect 9312 6944 9364 6996
rect 10692 6987 10744 6996
rect 10692 6953 10701 6987
rect 10701 6953 10735 6987
rect 10735 6953 10744 6987
rect 10692 6944 10744 6953
rect 12440 6944 12492 6996
rect 12624 6944 12676 6996
rect 13544 6944 13596 6996
rect 8116 6876 8168 6928
rect 4620 6808 4672 6860
rect 4988 6808 5040 6860
rect 3608 6783 3660 6792
rect 3608 6749 3617 6783
rect 3617 6749 3651 6783
rect 3651 6749 3660 6783
rect 3608 6740 3660 6749
rect 1952 6672 2004 6724
rect 3148 6672 3200 6724
rect 3976 6740 4028 6792
rect 5632 6808 5684 6860
rect 5356 6672 5408 6724
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 8024 6672 8076 6724
rect 1492 6604 1544 6656
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 3884 6604 3936 6656
rect 4712 6604 4764 6656
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 6736 6604 6788 6656
rect 7288 6604 7340 6656
rect 8116 6647 8168 6656
rect 8116 6613 8125 6647
rect 8125 6613 8159 6647
rect 8159 6613 8168 6647
rect 8116 6604 8168 6613
rect 8208 6604 8260 6656
rect 11060 6876 11112 6928
rect 11980 6876 12032 6928
rect 8760 6740 8812 6792
rect 9956 6808 10008 6860
rect 10416 6808 10468 6860
rect 10876 6851 10928 6860
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 10508 6740 10560 6792
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 12900 6808 12952 6860
rect 14004 6740 14056 6792
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 9404 6604 9456 6656
rect 11152 6672 11204 6724
rect 12624 6604 12676 6656
rect 13452 6604 13504 6656
rect 13544 6604 13596 6656
rect 1610 6502 1662 6554
rect 1674 6502 1726 6554
rect 1738 6502 1790 6554
rect 1802 6502 1854 6554
rect 1866 6502 1918 6554
rect 5610 6502 5662 6554
rect 5674 6502 5726 6554
rect 5738 6502 5790 6554
rect 5802 6502 5854 6554
rect 5866 6502 5918 6554
rect 9610 6502 9662 6554
rect 9674 6502 9726 6554
rect 9738 6502 9790 6554
rect 9802 6502 9854 6554
rect 9866 6502 9918 6554
rect 13610 6502 13662 6554
rect 13674 6502 13726 6554
rect 13738 6502 13790 6554
rect 13802 6502 13854 6554
rect 13866 6502 13918 6554
rect 2320 6400 2372 6452
rect 2412 6443 2464 6452
rect 2412 6409 2421 6443
rect 2421 6409 2455 6443
rect 2455 6409 2464 6443
rect 2412 6400 2464 6409
rect 4804 6400 4856 6452
rect 5356 6400 5408 6452
rect 5816 6400 5868 6452
rect 940 6332 992 6384
rect 4528 6375 4580 6384
rect 4528 6341 4537 6375
rect 4537 6341 4571 6375
rect 4571 6341 4580 6375
rect 4528 6332 4580 6341
rect 6092 6332 6144 6384
rect 4988 6264 5040 6316
rect 7472 6332 7524 6384
rect 4436 6128 4488 6180
rect 5448 6128 5500 6180
rect 5540 6171 5592 6180
rect 5540 6137 5549 6171
rect 5549 6137 5583 6171
rect 5583 6137 5592 6171
rect 5540 6128 5592 6137
rect 5816 6128 5868 6180
rect 6736 6196 6788 6248
rect 7104 6196 7156 6248
rect 8208 6332 8260 6384
rect 8760 6400 8812 6452
rect 9312 6400 9364 6452
rect 10508 6400 10560 6452
rect 10692 6400 10744 6452
rect 8116 6264 8168 6316
rect 16028 6264 16080 6316
rect 12348 6239 12400 6248
rect 12348 6205 12357 6239
rect 12357 6205 12391 6239
rect 12391 6205 12400 6239
rect 12348 6196 12400 6205
rect 3792 6060 3844 6112
rect 4712 6103 4764 6112
rect 4712 6069 4721 6103
rect 4721 6069 4755 6103
rect 4755 6069 4764 6103
rect 4712 6060 4764 6069
rect 7104 6103 7156 6112
rect 7104 6069 7113 6103
rect 7113 6069 7147 6103
rect 7147 6069 7156 6103
rect 7104 6060 7156 6069
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 8300 6060 8352 6112
rect 9588 6060 9640 6112
rect 12440 6060 12492 6112
rect 12716 6060 12768 6112
rect 950 5958 1002 6010
rect 1014 5958 1066 6010
rect 1078 5958 1130 6010
rect 1142 5958 1194 6010
rect 1206 5958 1258 6010
rect 4950 5958 5002 6010
rect 5014 5958 5066 6010
rect 5078 5958 5130 6010
rect 5142 5958 5194 6010
rect 5206 5958 5258 6010
rect 8950 5958 9002 6010
rect 9014 5958 9066 6010
rect 9078 5958 9130 6010
rect 9142 5958 9194 6010
rect 9206 5958 9258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 3608 5856 3660 5908
rect 4712 5856 4764 5908
rect 5264 5856 5316 5908
rect 6000 5856 6052 5908
rect 6828 5856 6880 5908
rect 3884 5788 3936 5840
rect 1492 5763 1544 5772
rect 1492 5729 1501 5763
rect 1501 5729 1535 5763
rect 1535 5729 1544 5763
rect 1492 5720 1544 5729
rect 3792 5720 3844 5772
rect 7104 5788 7156 5840
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 5264 5652 5316 5704
rect 6092 5720 6144 5772
rect 3148 5584 3200 5636
rect 1952 5516 2004 5568
rect 2596 5516 2648 5568
rect 7288 5720 7340 5772
rect 7932 5763 7984 5772
rect 7932 5729 7941 5763
rect 7941 5729 7975 5763
rect 7975 5729 7984 5763
rect 10324 5856 10376 5908
rect 11152 5856 11204 5908
rect 13452 5856 13504 5908
rect 14004 5856 14056 5908
rect 7932 5720 7984 5729
rect 9404 5720 9456 5772
rect 9680 5720 9732 5772
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 7196 5652 7248 5704
rect 10416 5652 10468 5704
rect 10968 5652 11020 5704
rect 6736 5627 6788 5636
rect 6736 5593 6745 5627
rect 6745 5593 6779 5627
rect 6779 5593 6788 5627
rect 6736 5584 6788 5593
rect 4528 5559 4580 5568
rect 4528 5525 4537 5559
rect 4537 5525 4571 5559
rect 4571 5525 4580 5559
rect 4528 5516 4580 5525
rect 6092 5516 6144 5568
rect 6644 5516 6696 5568
rect 8392 5516 8444 5568
rect 9956 5516 10008 5568
rect 10876 5516 10928 5568
rect 16488 5516 16540 5568
rect 1610 5414 1662 5466
rect 1674 5414 1726 5466
rect 1738 5414 1790 5466
rect 1802 5414 1854 5466
rect 1866 5414 1918 5466
rect 5610 5414 5662 5466
rect 5674 5414 5726 5466
rect 5738 5414 5790 5466
rect 5802 5414 5854 5466
rect 5866 5414 5918 5466
rect 9610 5414 9662 5466
rect 9674 5414 9726 5466
rect 9738 5414 9790 5466
rect 9802 5414 9854 5466
rect 9866 5414 9918 5466
rect 13610 5414 13662 5466
rect 13674 5414 13726 5466
rect 13738 5414 13790 5466
rect 13802 5414 13854 5466
rect 13866 5414 13918 5466
rect 1952 5355 2004 5364
rect 1952 5321 1961 5355
rect 1961 5321 1995 5355
rect 1995 5321 2004 5355
rect 1952 5312 2004 5321
rect 2044 5312 2096 5364
rect 2504 5312 2556 5364
rect 2596 5244 2648 5296
rect 756 5176 808 5228
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 2780 5176 2832 5228
rect 3516 5312 3568 5364
rect 3792 5244 3844 5296
rect 4528 5312 4580 5364
rect 5264 5312 5316 5364
rect 6736 5312 6788 5364
rect 8392 5312 8444 5364
rect 3240 5108 3292 5160
rect 3332 5040 3384 5092
rect 3148 5015 3200 5024
rect 3148 4981 3157 5015
rect 3157 4981 3191 5015
rect 3191 4981 3200 5015
rect 5356 5176 5408 5228
rect 7840 5244 7892 5296
rect 8024 5244 8076 5296
rect 9956 5312 10008 5364
rect 12624 5312 12676 5364
rect 12808 5312 12860 5364
rect 6368 5176 6420 5228
rect 6644 5108 6696 5160
rect 6920 5108 6972 5160
rect 7196 5108 7248 5160
rect 10324 5108 10376 5160
rect 10876 5151 10928 5160
rect 10876 5117 10885 5151
rect 10885 5117 10919 5151
rect 10919 5117 10928 5151
rect 10876 5108 10928 5117
rect 3148 4972 3200 4981
rect 5724 4972 5776 5024
rect 6368 4972 6420 5024
rect 8852 4972 8904 5024
rect 9312 4972 9364 5024
rect 11152 5108 11204 5160
rect 12624 5108 12676 5160
rect 13452 5108 13504 5160
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 950 4870 1002 4922
rect 1014 4870 1066 4922
rect 1078 4870 1130 4922
rect 1142 4870 1194 4922
rect 1206 4870 1258 4922
rect 4950 4870 5002 4922
rect 5014 4870 5066 4922
rect 5078 4870 5130 4922
rect 5142 4870 5194 4922
rect 5206 4870 5258 4922
rect 8950 4870 9002 4922
rect 9014 4870 9066 4922
rect 9078 4870 9130 4922
rect 9142 4870 9194 4922
rect 9206 4870 9258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 3424 4768 3476 4820
rect 3516 4811 3568 4820
rect 3516 4777 3525 4811
rect 3525 4777 3559 4811
rect 3559 4777 3568 4811
rect 3516 4768 3568 4777
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 5724 4700 5776 4752
rect 6276 4768 6328 4820
rect 7932 4768 7984 4820
rect 8300 4768 8352 4820
rect 8576 4768 8628 4820
rect 11152 4768 11204 4820
rect 11520 4768 11572 4820
rect 12348 4811 12400 4820
rect 12348 4777 12357 4811
rect 12357 4777 12391 4811
rect 12391 4777 12400 4811
rect 12348 4768 12400 4777
rect 12716 4768 12768 4820
rect 12992 4768 13044 4820
rect 3056 4675 3108 4684
rect 3056 4641 3065 4675
rect 3065 4641 3099 4675
rect 3099 4641 3108 4675
rect 3056 4632 3108 4641
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 6092 4675 6144 4684
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 6828 4632 6880 4684
rect 10324 4700 10376 4752
rect 11428 4700 11480 4752
rect 7288 4632 7340 4684
rect 2780 4496 2832 4548
rect 3240 4564 3292 4616
rect 7196 4564 7248 4616
rect 7748 4564 7800 4616
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 8392 4675 8444 4684
rect 8392 4641 8401 4675
rect 8401 4641 8435 4675
rect 8435 4641 8444 4675
rect 8392 4632 8444 4641
rect 9312 4632 9364 4684
rect 5540 4496 5592 4548
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 1952 4428 2004 4480
rect 3332 4428 3384 4480
rect 8116 4496 8168 4548
rect 9036 4564 9088 4616
rect 11060 4632 11112 4684
rect 12532 4700 12584 4752
rect 10784 4607 10836 4616
rect 10784 4573 10793 4607
rect 10793 4573 10827 4607
rect 10827 4573 10836 4607
rect 10784 4564 10836 4573
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 12992 4675 13044 4684
rect 12992 4641 13001 4675
rect 13001 4641 13035 4675
rect 13035 4641 13044 4675
rect 12992 4632 13044 4641
rect 10508 4496 10560 4548
rect 12440 4564 12492 4616
rect 14188 4700 14240 4752
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 9956 4428 10008 4480
rect 10140 4471 10192 4480
rect 10140 4437 10149 4471
rect 10149 4437 10183 4471
rect 10183 4437 10192 4471
rect 10140 4428 10192 4437
rect 10968 4471 11020 4480
rect 10968 4437 10977 4471
rect 10977 4437 11011 4471
rect 11011 4437 11020 4471
rect 10968 4428 11020 4437
rect 11888 4471 11940 4480
rect 11888 4437 11897 4471
rect 11897 4437 11931 4471
rect 11931 4437 11940 4471
rect 11888 4428 11940 4437
rect 14096 4471 14148 4480
rect 14096 4437 14105 4471
rect 14105 4437 14139 4471
rect 14139 4437 14148 4471
rect 14096 4428 14148 4437
rect 16764 4428 16816 4480
rect 1610 4326 1662 4378
rect 1674 4326 1726 4378
rect 1738 4326 1790 4378
rect 1802 4326 1854 4378
rect 1866 4326 1918 4378
rect 5610 4326 5662 4378
rect 5674 4326 5726 4378
rect 5738 4326 5790 4378
rect 5802 4326 5854 4378
rect 5866 4326 5918 4378
rect 9610 4326 9662 4378
rect 9674 4326 9726 4378
rect 9738 4326 9790 4378
rect 9802 4326 9854 4378
rect 9866 4326 9918 4378
rect 13610 4326 13662 4378
rect 13674 4326 13726 4378
rect 13738 4326 13790 4378
rect 13802 4326 13854 4378
rect 13866 4326 13918 4378
rect 2780 4224 2832 4276
rect 1952 4156 2004 4208
rect 3148 4156 3200 4208
rect 3332 4088 3384 4140
rect 3792 4088 3844 4140
rect 7288 4267 7340 4276
rect 7288 4233 7297 4267
rect 7297 4233 7331 4267
rect 7331 4233 7340 4267
rect 7288 4224 7340 4233
rect 8392 4224 8444 4276
rect 5448 4156 5500 4208
rect 6000 4156 6052 4208
rect 7012 4156 7064 4208
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 6460 4020 6512 4072
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 6736 4063 6788 4072
rect 6736 4029 6745 4063
rect 6745 4029 6779 4063
rect 6779 4029 6788 4063
rect 6736 4020 6788 4029
rect 5540 3952 5592 4004
rect 7380 4088 7432 4140
rect 8392 4088 8444 4140
rect 7196 3952 7248 4004
rect 8576 4020 8628 4072
rect 9956 4224 10008 4276
rect 11888 4224 11940 4276
rect 3332 3927 3384 3936
rect 3332 3893 3341 3927
rect 3341 3893 3375 3927
rect 3375 3893 3384 3927
rect 3332 3884 3384 3893
rect 3884 3884 3936 3936
rect 8024 3884 8076 3936
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 9404 4020 9456 4072
rect 10416 4020 10468 4072
rect 14096 4156 14148 4208
rect 12716 4088 12768 4140
rect 12624 4020 12676 4072
rect 13452 4020 13504 4072
rect 10140 3884 10192 3936
rect 10784 3884 10836 3936
rect 12440 3884 12492 3936
rect 950 3782 1002 3834
rect 1014 3782 1066 3834
rect 1078 3782 1130 3834
rect 1142 3782 1194 3834
rect 1206 3782 1258 3834
rect 4950 3782 5002 3834
rect 5014 3782 5066 3834
rect 5078 3782 5130 3834
rect 5142 3782 5194 3834
rect 5206 3782 5258 3834
rect 8950 3782 9002 3834
rect 9014 3782 9066 3834
rect 9078 3782 9130 3834
rect 9142 3782 9194 3834
rect 9206 3782 9258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 3884 3680 3936 3732
rect 6184 3680 6236 3732
rect 6460 3680 6512 3732
rect 7196 3680 7248 3732
rect 8116 3723 8168 3732
rect 8116 3689 8125 3723
rect 8125 3689 8159 3723
rect 8159 3689 8168 3723
rect 8116 3680 8168 3689
rect 8300 3680 8352 3732
rect 3332 3476 3384 3528
rect 9680 3680 9732 3732
rect 10876 3680 10928 3732
rect 5080 3476 5132 3528
rect 940 3408 992 3460
rect 5540 3544 5592 3596
rect 5448 3519 5500 3528
rect 5448 3485 5457 3519
rect 5457 3485 5491 3519
rect 5491 3485 5500 3519
rect 5448 3476 5500 3485
rect 6644 3544 6696 3596
rect 8392 3544 8444 3596
rect 10692 3544 10744 3596
rect 10876 3544 10928 3596
rect 7840 3408 7892 3460
rect 3700 3340 3752 3392
rect 4068 3340 4120 3392
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 5540 3340 5592 3392
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 8024 3340 8076 3392
rect 10600 3476 10652 3528
rect 10968 3476 11020 3528
rect 11336 3519 11388 3528
rect 11336 3485 11345 3519
rect 11345 3485 11379 3519
rect 11379 3485 11388 3519
rect 11336 3476 11388 3485
rect 12440 3612 12492 3664
rect 15936 3519 15988 3528
rect 15936 3485 15945 3519
rect 15945 3485 15979 3519
rect 15979 3485 15988 3519
rect 15936 3476 15988 3485
rect 9496 3408 9548 3460
rect 12808 3408 12860 3460
rect 13360 3408 13412 3460
rect 9680 3340 9732 3392
rect 9956 3340 10008 3392
rect 10600 3383 10652 3392
rect 10600 3349 10609 3383
rect 10609 3349 10643 3383
rect 10643 3349 10652 3383
rect 10600 3340 10652 3349
rect 10692 3340 10744 3392
rect 11428 3383 11480 3392
rect 11428 3349 11437 3383
rect 11437 3349 11471 3383
rect 11471 3349 11480 3383
rect 11428 3340 11480 3349
rect 14464 3383 14516 3392
rect 14464 3349 14473 3383
rect 14473 3349 14507 3383
rect 14507 3349 14516 3383
rect 14464 3340 14516 3349
rect 16028 3383 16080 3392
rect 16028 3349 16037 3383
rect 16037 3349 16071 3383
rect 16071 3349 16080 3383
rect 16028 3340 16080 3349
rect 1610 3238 1662 3290
rect 1674 3238 1726 3290
rect 1738 3238 1790 3290
rect 1802 3238 1854 3290
rect 1866 3238 1918 3290
rect 5610 3238 5662 3290
rect 5674 3238 5726 3290
rect 5738 3238 5790 3290
rect 5802 3238 5854 3290
rect 5866 3238 5918 3290
rect 9610 3238 9662 3290
rect 9674 3238 9726 3290
rect 9738 3238 9790 3290
rect 9802 3238 9854 3290
rect 9866 3238 9918 3290
rect 13610 3238 13662 3290
rect 13674 3238 13726 3290
rect 13738 3238 13790 3290
rect 13802 3238 13854 3290
rect 13866 3238 13918 3290
rect 3240 3136 3292 3188
rect 4436 3136 4488 3188
rect 5080 3136 5132 3188
rect 3700 3068 3752 3120
rect 1308 3000 1360 3052
rect 5540 3136 5592 3188
rect 7196 3136 7248 3188
rect 8024 3136 8076 3188
rect 8576 3136 8628 3188
rect 3792 2975 3844 2984
rect 3792 2941 3801 2975
rect 3801 2941 3835 2975
rect 3835 2941 3844 2975
rect 3792 2932 3844 2941
rect 9128 3068 9180 3120
rect 9404 3136 9456 3188
rect 10416 3136 10468 3188
rect 10600 3136 10652 3188
rect 10692 3136 10744 3188
rect 10324 3111 10376 3120
rect 10324 3077 10333 3111
rect 10333 3077 10367 3111
rect 10367 3077 10376 3111
rect 10324 3068 10376 3077
rect 5356 2932 5408 2984
rect 5448 2932 5500 2984
rect 6368 2932 6420 2984
rect 10508 3043 10560 3052
rect 10508 3009 10517 3043
rect 10517 3009 10551 3043
rect 10551 3009 10560 3043
rect 10508 3000 10560 3009
rect 10968 3111 11020 3120
rect 10968 3077 10977 3111
rect 10977 3077 11011 3111
rect 11011 3077 11020 3111
rect 14464 3136 14516 3188
rect 15936 3136 15988 3188
rect 16028 3136 16080 3188
rect 10968 3068 11020 3077
rect 12716 3068 12768 3120
rect 13452 3000 13504 3052
rect 15660 3043 15712 3052
rect 15660 3009 15669 3043
rect 15669 3009 15703 3043
rect 15703 3009 15712 3043
rect 15660 3000 15712 3009
rect 12440 2932 12492 2984
rect 20 2796 72 2848
rect 7288 2839 7340 2848
rect 7288 2805 7297 2839
rect 7297 2805 7331 2839
rect 7331 2805 7340 2839
rect 7288 2796 7340 2805
rect 9128 2796 9180 2848
rect 10416 2796 10468 2848
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 11336 2839 11388 2848
rect 11336 2805 11345 2839
rect 11345 2805 11379 2839
rect 11379 2805 11388 2839
rect 11336 2796 11388 2805
rect 15752 2839 15804 2848
rect 15752 2805 15761 2839
rect 15761 2805 15795 2839
rect 15795 2805 15804 2839
rect 15752 2796 15804 2805
rect 16764 2796 16816 2848
rect 950 2694 1002 2746
rect 1014 2694 1066 2746
rect 1078 2694 1130 2746
rect 1142 2694 1194 2746
rect 1206 2694 1258 2746
rect 4950 2694 5002 2746
rect 5014 2694 5066 2746
rect 5078 2694 5130 2746
rect 5142 2694 5194 2746
rect 5206 2694 5258 2746
rect 8950 2694 9002 2746
rect 9014 2694 9066 2746
rect 9078 2694 9130 2746
rect 9142 2694 9194 2746
rect 9206 2694 9258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 7840 2592 7892 2644
rect 12440 2592 12492 2644
rect 15936 2592 15988 2644
rect 11152 2567 11204 2576
rect 6000 2456 6052 2508
rect 7288 2456 7340 2508
rect 2872 2388 2924 2440
rect 4068 2388 4120 2440
rect 6276 2388 6328 2440
rect 940 2320 992 2372
rect 3240 2295 3292 2304
rect 3240 2261 3249 2295
rect 3249 2261 3283 2295
rect 3283 2261 3292 2295
rect 3240 2252 3292 2261
rect 4528 2295 4580 2304
rect 4528 2261 4537 2295
rect 4537 2261 4571 2295
rect 4571 2261 4580 2295
rect 4528 2252 4580 2261
rect 6460 2252 6512 2304
rect 7104 2320 7156 2372
rect 11152 2533 11161 2567
rect 11161 2533 11195 2567
rect 11195 2533 11204 2567
rect 11152 2524 11204 2533
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 10876 2431 10928 2440
rect 10876 2397 10885 2431
rect 10885 2397 10919 2431
rect 10919 2397 10928 2431
rect 10876 2388 10928 2397
rect 11336 2431 11388 2440
rect 11336 2397 11345 2431
rect 11345 2397 11379 2431
rect 11379 2397 11388 2431
rect 11336 2388 11388 2397
rect 11428 2388 11480 2440
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 15752 2388 15804 2440
rect 7380 2252 7432 2304
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 11612 2252 11664 2304
rect 14832 2295 14884 2304
rect 14832 2261 14841 2295
rect 14841 2261 14875 2295
rect 14875 2261 14884 2295
rect 14832 2252 14884 2261
rect 16948 2320 17000 2372
rect 16396 2295 16448 2304
rect 16396 2261 16405 2295
rect 16405 2261 16439 2295
rect 16439 2261 16448 2295
rect 16396 2252 16448 2261
rect 1610 2150 1662 2202
rect 1674 2150 1726 2202
rect 1738 2150 1790 2202
rect 1802 2150 1854 2202
rect 1866 2150 1918 2202
rect 5610 2150 5662 2202
rect 5674 2150 5726 2202
rect 5738 2150 5790 2202
rect 5802 2150 5854 2202
rect 5866 2150 5918 2202
rect 9610 2150 9662 2202
rect 9674 2150 9726 2202
rect 9738 2150 9790 2202
rect 9802 2150 9854 2202
rect 9866 2150 9918 2202
rect 13610 2150 13662 2202
rect 13674 2150 13726 2202
rect 13738 2150 13790 2202
rect 13802 2150 13854 2202
rect 13866 2150 13918 2202
<< metal2 >>
rect 662 17200 718 18000
rect 1490 17776 1546 17785
rect 1490 17711 1546 17720
rect 676 15502 704 17200
rect 1398 16008 1454 16017
rect 1398 15943 1454 15952
rect 950 15804 1258 15813
rect 950 15802 956 15804
rect 1012 15802 1036 15804
rect 1092 15802 1116 15804
rect 1172 15802 1196 15804
rect 1252 15802 1258 15804
rect 1012 15750 1014 15802
rect 1194 15750 1196 15802
rect 950 15748 956 15750
rect 1012 15748 1036 15750
rect 1092 15748 1116 15750
rect 1172 15748 1196 15750
rect 1252 15748 1258 15750
rect 950 15739 1258 15748
rect 664 15496 716 15502
rect 664 15438 716 15444
rect 1412 15094 1440 15943
rect 1504 15706 1532 17711
rect 2594 17200 2650 18000
rect 4526 17200 4582 18000
rect 5814 17200 5870 18000
rect 7746 17354 7802 18000
rect 9034 17354 9090 18000
rect 7746 17326 7880 17354
rect 7746 17200 7802 17326
rect 2608 16574 2636 17200
rect 2608 16546 2820 16574
rect 2792 15706 2820 16546
rect 1492 15700 1544 15706
rect 1492 15642 1544 15648
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 4540 15502 4568 17200
rect 4950 15804 5258 15813
rect 4950 15802 4956 15804
rect 5012 15802 5036 15804
rect 5092 15802 5116 15804
rect 5172 15802 5196 15804
rect 5252 15802 5258 15804
rect 5012 15750 5014 15802
rect 5194 15750 5196 15802
rect 4950 15748 4956 15750
rect 5012 15748 5036 15750
rect 5092 15748 5116 15750
rect 5172 15748 5196 15750
rect 5252 15748 5258 15750
rect 4950 15739 5258 15748
rect 5828 15706 5856 17200
rect 7852 15706 7880 17326
rect 9034 17326 9352 17354
rect 9034 17200 9090 17326
rect 8950 15804 9258 15813
rect 8950 15802 8956 15804
rect 9012 15802 9036 15804
rect 9092 15802 9116 15804
rect 9172 15802 9196 15804
rect 9252 15802 9258 15804
rect 9012 15750 9014 15802
rect 9194 15750 9196 15802
rect 8950 15748 8956 15750
rect 9012 15748 9036 15750
rect 9092 15748 9116 15750
rect 9172 15748 9196 15750
rect 9252 15748 9258 15750
rect 8950 15739 9258 15748
rect 9324 15706 9352 17326
rect 10966 17200 11022 18000
rect 12898 17200 12954 18000
rect 14186 17200 14242 18000
rect 16118 17354 16174 18000
rect 16118 17326 16252 17354
rect 16118 17200 16174 17326
rect 10980 15722 11008 17200
rect 12912 16574 12940 17200
rect 12820 16546 12940 16574
rect 14200 16574 14228 17200
rect 14200 16546 14412 16574
rect 10980 15706 11100 15722
rect 12820 15706 12848 16546
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 14384 15706 14412 16546
rect 16224 15706 16252 17326
rect 17406 17200 17462 18000
rect 16486 16416 16542 16425
rect 16486 16351 16542 16360
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 9312 15700 9364 15706
rect 10980 15700 11112 15706
rect 10980 15694 11060 15700
rect 9312 15642 9364 15648
rect 11060 15642 11112 15648
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 2320 15428 2372 15434
rect 2320 15370 2372 15376
rect 3056 15428 3108 15434
rect 3056 15370 3108 15376
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 8208 15428 8260 15434
rect 8208 15370 8260 15376
rect 1610 15260 1918 15269
rect 1610 15258 1616 15260
rect 1672 15258 1696 15260
rect 1752 15258 1776 15260
rect 1832 15258 1856 15260
rect 1912 15258 1918 15260
rect 1672 15206 1674 15258
rect 1854 15206 1856 15258
rect 1610 15204 1616 15206
rect 1672 15204 1696 15206
rect 1752 15204 1776 15206
rect 1832 15204 1856 15206
rect 1912 15204 1918 15206
rect 1610 15195 1918 15204
rect 2332 15162 2360 15370
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 1400 15088 1452 15094
rect 1400 15030 1452 15036
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 950 14716 1258 14725
rect 950 14714 956 14716
rect 1012 14714 1036 14716
rect 1092 14714 1116 14716
rect 1172 14714 1196 14716
rect 1252 14714 1258 14716
rect 1012 14662 1014 14714
rect 1194 14662 1196 14714
rect 950 14660 956 14662
rect 1012 14660 1036 14662
rect 1092 14660 1116 14662
rect 1172 14660 1196 14662
rect 1252 14660 1258 14662
rect 950 14651 1258 14660
rect 1610 14172 1918 14181
rect 1610 14170 1616 14172
rect 1672 14170 1696 14172
rect 1752 14170 1776 14172
rect 1832 14170 1856 14172
rect 1912 14170 1918 14172
rect 1672 14118 1674 14170
rect 1854 14118 1856 14170
rect 1610 14116 1616 14118
rect 1672 14116 1696 14118
rect 1752 14116 1776 14118
rect 1832 14116 1856 14118
rect 1912 14116 1918 14118
rect 1610 14107 1918 14116
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1412 13705 1440 13874
rect 1676 13728 1728 13734
rect 1398 13696 1454 13705
rect 1676 13670 1728 13676
rect 950 13628 1258 13637
rect 1398 13631 1454 13640
rect 950 13626 956 13628
rect 1012 13626 1036 13628
rect 1092 13626 1116 13628
rect 1172 13626 1196 13628
rect 1252 13626 1258 13628
rect 1012 13574 1014 13626
rect 1194 13574 1196 13626
rect 950 13572 956 13574
rect 1012 13572 1036 13574
rect 1092 13572 1116 13574
rect 1172 13572 1196 13574
rect 1252 13572 1258 13574
rect 950 13563 1258 13572
rect 1688 13258 1716 13670
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 1610 13084 1918 13093
rect 1610 13082 1616 13084
rect 1672 13082 1696 13084
rect 1752 13082 1776 13084
rect 1832 13082 1856 13084
rect 1912 13082 1918 13084
rect 1672 13030 1674 13082
rect 1854 13030 1856 13082
rect 1610 13028 1616 13030
rect 1672 13028 1696 13030
rect 1752 13028 1776 13030
rect 1832 13028 1856 13030
rect 1912 13028 1918 13030
rect 1610 13019 1918 13028
rect 1964 12986 1992 13874
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 950 12540 1258 12549
rect 950 12538 956 12540
rect 1012 12538 1036 12540
rect 1092 12538 1116 12540
rect 1172 12538 1196 12540
rect 1252 12538 1258 12540
rect 1012 12486 1014 12538
rect 1194 12486 1196 12538
rect 950 12484 956 12486
rect 1012 12484 1036 12486
rect 1092 12484 1116 12486
rect 1172 12484 1196 12486
rect 1252 12484 1258 12486
rect 950 12475 1258 12484
rect 1504 12345 1532 12582
rect 2148 12442 2176 12786
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 2332 12102 2360 14962
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2884 13938 2912 14214
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2596 13184 2648 13190
rect 2884 13138 2912 13874
rect 3068 13530 3096 15370
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 5610 15260 5918 15269
rect 5610 15258 5616 15260
rect 5672 15258 5696 15260
rect 5752 15258 5776 15260
rect 5832 15258 5856 15260
rect 5912 15258 5918 15260
rect 5672 15206 5674 15258
rect 5854 15206 5856 15258
rect 5610 15204 5616 15206
rect 5672 15204 5696 15206
rect 5752 15204 5776 15206
rect 5832 15204 5856 15206
rect 5912 15204 5918 15206
rect 5610 15195 5918 15204
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 2596 13126 2648 13132
rect 2608 12986 2636 13126
rect 2792 13110 2912 13138
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 1610 11996 1918 12005
rect 1610 11994 1616 11996
rect 1672 11994 1696 11996
rect 1752 11994 1776 11996
rect 1832 11994 1856 11996
rect 1912 11994 1918 11996
rect 1672 11942 1674 11994
rect 1854 11942 1856 11994
rect 1610 11940 1616 11942
rect 1672 11940 1696 11942
rect 1752 11940 1776 11942
rect 1832 11940 1856 11942
rect 1912 11940 1918 11942
rect 1610 11931 1918 11940
rect 950 11452 1258 11461
rect 950 11450 956 11452
rect 1012 11450 1036 11452
rect 1092 11450 1116 11452
rect 1172 11450 1196 11452
rect 1252 11450 1258 11452
rect 1012 11398 1014 11450
rect 1194 11398 1196 11450
rect 950 11396 956 11398
rect 1012 11396 1036 11398
rect 1092 11396 1116 11398
rect 1172 11396 1196 11398
rect 1252 11396 1258 11398
rect 950 11387 1258 11396
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1504 10810 1532 10950
rect 1610 10908 1918 10917
rect 1610 10906 1616 10908
rect 1672 10906 1696 10908
rect 1752 10906 1776 10908
rect 1832 10906 1856 10908
rect 1912 10906 1918 10908
rect 1672 10854 1674 10906
rect 1854 10854 1856 10906
rect 1610 10852 1616 10854
rect 1672 10852 1696 10854
rect 1752 10852 1776 10854
rect 1832 10852 1856 10854
rect 1912 10852 1918 10854
rect 1610 10843 1918 10852
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 950 10364 1258 10373
rect 950 10362 956 10364
rect 1012 10362 1036 10364
rect 1092 10362 1116 10364
rect 1172 10362 1196 10364
rect 1252 10362 1258 10364
rect 1012 10310 1014 10362
rect 1194 10310 1196 10362
rect 950 10308 956 10310
rect 1012 10308 1036 10310
rect 1092 10308 1116 10310
rect 1172 10308 1196 10310
rect 1252 10308 1258 10310
rect 950 10299 1258 10308
rect 940 10260 992 10266
rect 940 10202 992 10208
rect 952 10169 980 10202
rect 938 10160 994 10169
rect 938 10095 994 10104
rect 1412 9586 1440 10542
rect 1610 9820 1918 9829
rect 1610 9818 1616 9820
rect 1672 9818 1696 9820
rect 1752 9818 1776 9820
rect 1832 9818 1856 9820
rect 1912 9818 1918 9820
rect 1672 9766 1674 9818
rect 1854 9766 1856 9818
rect 1610 9764 1616 9766
rect 1672 9764 1696 9766
rect 1752 9764 1776 9766
rect 1832 9764 1856 9766
rect 1912 9764 1918 9766
rect 1610 9755 1918 9764
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 950 9276 1258 9285
rect 950 9274 956 9276
rect 1012 9274 1036 9276
rect 1092 9274 1116 9276
rect 1172 9274 1196 9276
rect 1252 9274 1258 9276
rect 1012 9222 1014 9274
rect 1194 9222 1196 9274
rect 950 9220 956 9222
rect 1012 9220 1036 9222
rect 1092 9220 1116 9222
rect 1172 9220 1196 9222
rect 1252 9220 1258 9222
rect 950 9211 1258 9220
rect 938 8936 994 8945
rect 938 8871 940 8880
rect 992 8871 994 8880
rect 940 8842 992 8848
rect 950 8188 1258 8197
rect 950 8186 956 8188
rect 1012 8186 1036 8188
rect 1092 8186 1116 8188
rect 1172 8186 1196 8188
rect 1252 8186 1258 8188
rect 1012 8134 1014 8186
rect 1194 8134 1196 8186
rect 950 8132 956 8134
rect 1012 8132 1036 8134
rect 1092 8132 1116 8134
rect 1172 8132 1196 8134
rect 1252 8132 1258 8134
rect 950 8123 1258 8132
rect 1412 7954 1440 9522
rect 1964 8974 1992 12038
rect 2228 11144 2280 11150
rect 2516 11132 2544 12582
rect 2792 12322 2820 13110
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2884 12782 2912 12922
rect 2976 12850 3004 13330
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2700 12294 2820 12322
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2700 12238 2728 12294
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2792 11234 2820 12294
rect 2884 11354 2912 12310
rect 3160 11354 3188 14962
rect 4950 14716 5258 14725
rect 4950 14714 4956 14716
rect 5012 14714 5036 14716
rect 5092 14714 5116 14716
rect 5172 14714 5196 14716
rect 5252 14714 5258 14716
rect 5012 14662 5014 14714
rect 5194 14662 5196 14714
rect 4950 14660 4956 14662
rect 5012 14660 5036 14662
rect 5092 14660 5116 14662
rect 5172 14660 5196 14662
rect 5252 14660 5258 14662
rect 4950 14651 5258 14660
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3804 14074 3832 14214
rect 5092 14074 5120 14282
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3252 11762 3280 12718
rect 3344 12238 3372 13466
rect 4172 13394 4200 13942
rect 4540 13938 4568 14010
rect 5552 13938 5580 14214
rect 5610 14172 5918 14181
rect 5610 14170 5616 14172
rect 5672 14170 5696 14172
rect 5752 14170 5776 14172
rect 5832 14170 5856 14172
rect 5912 14170 5918 14172
rect 5672 14118 5674 14170
rect 5854 14118 5856 14170
rect 5610 14116 5616 14118
rect 5672 14116 5696 14118
rect 5752 14116 5776 14118
rect 5832 14116 5856 14118
rect 5912 14116 5918 14118
rect 5610 14107 5918 14116
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 4080 12918 4108 13194
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 4080 12434 4108 12854
rect 4264 12714 4292 13806
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4080 12406 4200 12434
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3620 11694 3648 12038
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 2792 11206 3096 11234
rect 2792 11150 2820 11206
rect 2280 11104 2544 11132
rect 2780 11144 2832 11150
rect 2228 11086 2280 11092
rect 2780 11086 2832 11092
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2148 9518 2176 9590
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2056 9178 2084 9454
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1610 8732 1918 8741
rect 1610 8730 1616 8732
rect 1672 8730 1696 8732
rect 1752 8730 1776 8732
rect 1832 8730 1856 8732
rect 1912 8730 1918 8732
rect 1672 8678 1674 8730
rect 1854 8678 1856 8730
rect 1610 8676 1616 8678
rect 1672 8676 1696 8678
rect 1752 8676 1776 8678
rect 1832 8676 1856 8678
rect 1912 8676 1918 8678
rect 1610 8667 1918 8676
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 2044 7744 2096 7750
rect 2148 7732 2176 9454
rect 2096 7704 2176 7732
rect 2044 7686 2096 7692
rect 1610 7644 1918 7653
rect 1610 7642 1616 7644
rect 1672 7642 1696 7644
rect 1752 7642 1776 7644
rect 1832 7642 1856 7644
rect 1912 7642 1918 7644
rect 1672 7590 1674 7642
rect 1854 7590 1856 7642
rect 1610 7588 1616 7590
rect 1672 7588 1696 7590
rect 1752 7588 1776 7590
rect 1832 7588 1856 7590
rect 1912 7588 1918 7590
rect 1610 7579 1918 7588
rect 2056 7546 2084 7686
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 950 7100 1258 7109
rect 950 7098 956 7100
rect 1012 7098 1036 7100
rect 1092 7098 1116 7100
rect 1172 7098 1196 7100
rect 1252 7098 1258 7100
rect 1012 7046 1014 7098
rect 1194 7046 1196 7098
rect 950 7044 956 7046
rect 1012 7044 1036 7046
rect 1092 7044 1116 7046
rect 1172 7044 1196 7046
rect 1252 7044 1258 7046
rect 950 7035 1258 7044
rect 938 6896 994 6905
rect 938 6831 994 6840
rect 952 6390 980 6831
rect 1952 6724 2004 6730
rect 2004 6684 2084 6712
rect 1952 6666 2004 6672
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 940 6384 992 6390
rect 940 6326 992 6332
rect 950 6012 1258 6021
rect 950 6010 956 6012
rect 1012 6010 1036 6012
rect 1092 6010 1116 6012
rect 1172 6010 1196 6012
rect 1252 6010 1258 6012
rect 1012 5958 1014 6010
rect 1194 5958 1196 6010
rect 950 5956 956 5958
rect 1012 5956 1036 5958
rect 1092 5956 1116 5958
rect 1172 5956 1196 5958
rect 1252 5956 1258 5958
rect 950 5947 1258 5956
rect 1504 5778 1532 6598
rect 1610 6556 1918 6565
rect 1610 6554 1616 6556
rect 1672 6554 1696 6556
rect 1752 6554 1776 6556
rect 1832 6554 1856 6556
rect 1912 6554 1918 6556
rect 1672 6502 1674 6554
rect 1854 6502 1856 6554
rect 1610 6500 1616 6502
rect 1672 6500 1696 6502
rect 1752 6500 1776 6502
rect 1832 6500 1856 6502
rect 1912 6500 1918 6502
rect 1610 6491 1918 6500
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1610 5468 1918 5477
rect 1610 5466 1616 5468
rect 1672 5466 1696 5468
rect 1752 5466 1776 5468
rect 1832 5466 1856 5468
rect 1912 5466 1918 5468
rect 1672 5414 1674 5466
rect 1854 5414 1856 5466
rect 1610 5412 1616 5414
rect 1672 5412 1696 5414
rect 1752 5412 1776 5414
rect 1832 5412 1856 5414
rect 1912 5412 1918 5414
rect 1610 5403 1918 5412
rect 1964 5370 1992 5510
rect 2056 5370 2084 6684
rect 2240 6338 2268 11086
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2976 10470 3004 11018
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2700 8498 2728 9318
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2332 7478 2360 8366
rect 2320 7472 2372 7478
rect 2372 7432 2544 7460
rect 2320 7414 2372 7420
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2332 6458 2360 7142
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2424 6458 2452 6802
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2240 6310 2360 6338
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 756 5228 808 5234
rect 756 5170 808 5176
rect 768 5137 796 5170
rect 754 5128 810 5137
rect 754 5063 810 5072
rect 950 4924 1258 4933
rect 950 4922 956 4924
rect 1012 4922 1036 4924
rect 1092 4922 1116 4924
rect 1172 4922 1196 4924
rect 1252 4922 1258 4924
rect 1012 4870 1014 4922
rect 1194 4870 1196 4922
rect 950 4868 956 4870
rect 1012 4868 1036 4870
rect 1092 4868 1116 4870
rect 1172 4868 1196 4870
rect 1252 4868 1258 4870
rect 950 4859 1258 4868
rect 2332 4622 2360 6310
rect 2424 5234 2452 6394
rect 2516 5370 2544 7432
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2884 5794 2912 7142
rect 2792 5766 2912 5794
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2608 5302 2636 5510
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2792 5234 2820 5766
rect 2976 5522 3004 10406
rect 2884 5494 3004 5522
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1610 4380 1918 4389
rect 1610 4378 1616 4380
rect 1672 4378 1696 4380
rect 1752 4378 1776 4380
rect 1832 4378 1856 4380
rect 1912 4378 1918 4380
rect 1672 4326 1674 4378
rect 1854 4326 1856 4378
rect 1610 4324 1616 4326
rect 1672 4324 1696 4326
rect 1752 4324 1776 4326
rect 1832 4324 1856 4326
rect 1912 4324 1918 4326
rect 1610 4315 1918 4324
rect 1964 4214 1992 4422
rect 2792 4282 2820 4490
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 950 3836 1258 3845
rect 950 3834 956 3836
rect 1012 3834 1036 3836
rect 1092 3834 1116 3836
rect 1172 3834 1196 3836
rect 1252 3834 1258 3836
rect 1012 3782 1014 3834
rect 1194 3782 1196 3834
rect 950 3780 956 3782
rect 1012 3780 1036 3782
rect 1092 3780 1116 3782
rect 1172 3780 1196 3782
rect 1252 3780 1258 3782
rect 950 3771 1258 3780
rect 938 3496 994 3505
rect 938 3431 940 3440
rect 992 3431 994 3440
rect 940 3402 992 3408
rect 1610 3292 1918 3301
rect 1610 3290 1616 3292
rect 1672 3290 1696 3292
rect 1752 3290 1776 3292
rect 1832 3290 1856 3292
rect 1912 3290 1918 3292
rect 1672 3238 1674 3290
rect 1854 3238 1856 3290
rect 1610 3236 1616 3238
rect 1672 3236 1696 3238
rect 1752 3236 1776 3238
rect 1832 3236 1856 3238
rect 1912 3236 1918 3238
rect 1610 3227 1918 3236
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 32 800 60 2790
rect 950 2748 1258 2757
rect 950 2746 956 2748
rect 1012 2746 1036 2748
rect 1092 2746 1116 2748
rect 1172 2746 1196 2748
rect 1252 2746 1258 2748
rect 1012 2694 1014 2746
rect 1194 2694 1196 2746
rect 950 2692 956 2694
rect 1012 2692 1036 2694
rect 1092 2692 1116 2694
rect 1172 2692 1196 2694
rect 1252 2692 1258 2694
rect 950 2683 1258 2692
rect 940 2372 992 2378
rect 940 2314 992 2320
rect 952 1465 980 2314
rect 938 1456 994 1465
rect 938 1391 994 1400
rect 1320 800 1348 2994
rect 2884 2446 2912 5494
rect 3068 4690 3096 11206
rect 3252 11082 3280 11494
rect 3896 11354 3924 12174
rect 4080 11694 4108 12174
rect 4172 11694 4200 12406
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 4080 11150 4108 11630
rect 4356 11218 4384 12786
rect 4540 11898 4568 13874
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4632 13530 4660 13806
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4724 12850 4752 13670
rect 4816 13462 4844 13874
rect 5368 13802 5396 13874
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 4950 13628 5258 13637
rect 4950 13626 4956 13628
rect 5012 13626 5036 13628
rect 5092 13626 5116 13628
rect 5172 13626 5196 13628
rect 5252 13626 5258 13628
rect 5012 13574 5014 13626
rect 5194 13574 5196 13626
rect 4950 13572 4956 13574
rect 5012 13572 5036 13574
rect 5092 13572 5116 13574
rect 5172 13572 5196 13574
rect 5252 13572 5258 13574
rect 4950 13563 5258 13572
rect 5368 13462 5396 13738
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4908 12986 4936 13126
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 5552 12850 5580 13398
rect 5610 13084 5918 13093
rect 5610 13082 5616 13084
rect 5672 13082 5696 13084
rect 5752 13082 5776 13084
rect 5832 13082 5856 13084
rect 5912 13082 5918 13084
rect 5672 13030 5674 13082
rect 5854 13030 5856 13082
rect 5610 13028 5616 13030
rect 5672 13028 5696 13030
rect 5752 13028 5776 13030
rect 5832 13028 5856 13030
rect 5912 13028 5918 13030
rect 5610 13019 5918 13028
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5092 12646 5120 12786
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 4950 12540 5258 12549
rect 4950 12538 4956 12540
rect 5012 12538 5036 12540
rect 5092 12538 5116 12540
rect 5172 12538 5196 12540
rect 5252 12538 5258 12540
rect 5012 12486 5014 12538
rect 5194 12486 5196 12538
rect 4950 12484 4956 12486
rect 5012 12484 5036 12486
rect 5092 12484 5116 12486
rect 5172 12484 5196 12486
rect 5252 12484 5258 12486
rect 4950 12475 5258 12484
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4540 11218 4568 11834
rect 4950 11452 5258 11461
rect 4950 11450 4956 11452
rect 5012 11450 5036 11452
rect 5092 11450 5116 11452
rect 5172 11450 5196 11452
rect 5252 11450 5258 11452
rect 5012 11398 5014 11450
rect 5194 11398 5196 11450
rect 4950 11396 4956 11398
rect 5012 11396 5036 11398
rect 5092 11396 5116 11398
rect 5172 11396 5196 11398
rect 5252 11396 5258 11398
rect 4950 11387 5258 11396
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3344 9518 3372 10610
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3160 7002 3188 7346
rect 3436 7313 3464 11018
rect 4080 9586 4108 11086
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10674 4292 10950
rect 4356 10810 4384 11154
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3528 9042 3556 9318
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3896 8634 3924 8978
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3896 7886 3924 8570
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 4172 8090 4200 8502
rect 4264 8294 4292 10610
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4632 9586 4660 9998
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4172 7886 4200 8026
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3896 7478 3924 7822
rect 4172 7546 4200 7822
rect 4264 7750 4292 8230
rect 4448 7954 4476 8774
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4264 7546 4292 7686
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3422 7304 3478 7313
rect 3422 7239 3478 7248
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 3160 5642 3188 6666
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3160 5030 3188 5578
rect 3252 5166 3280 6598
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3344 5098 3372 7142
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 3160 4214 3188 4966
rect 3436 4826 3464 7239
rect 3896 7002 3924 7414
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3988 6798 4016 7278
rect 4172 7274 4200 7482
rect 4448 7342 4476 7890
rect 4540 7449 4568 8434
rect 4526 7440 4582 7449
rect 4526 7375 4582 7384
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4172 6866 4200 7210
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3620 5914 3648 6734
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3804 5778 3832 6054
rect 3896 5846 3924 6598
rect 4448 6186 4476 7278
rect 4540 6390 4568 7375
rect 4632 6866 4660 8910
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4724 6662 4752 10406
rect 4816 10130 4844 10542
rect 5092 10538 5120 11018
rect 5368 10810 5396 12650
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 12306 5580 12582
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5460 11830 5488 12038
rect 5610 11996 5918 12005
rect 5610 11994 5616 11996
rect 5672 11994 5696 11996
rect 5752 11994 5776 11996
rect 5832 11994 5856 11996
rect 5912 11994 5918 11996
rect 5672 11942 5674 11994
rect 5854 11942 5856 11994
rect 5610 11940 5616 11942
rect 5672 11940 5696 11942
rect 5752 11940 5776 11942
rect 5832 11940 5856 11942
rect 5912 11940 5918 11942
rect 5610 11931 5918 11940
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5368 10538 5396 10746
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 4950 10364 5258 10373
rect 4950 10362 4956 10364
rect 5012 10362 5036 10364
rect 5092 10362 5116 10364
rect 5172 10362 5196 10364
rect 5252 10362 5258 10364
rect 5012 10310 5014 10362
rect 5194 10310 5196 10362
rect 4950 10308 4956 10310
rect 5012 10308 5036 10310
rect 5092 10308 5116 10310
rect 5172 10308 5196 10310
rect 5252 10308 5258 10310
rect 4950 10299 5258 10308
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 4950 9276 5258 9285
rect 4950 9274 4956 9276
rect 5012 9274 5036 9276
rect 5092 9274 5116 9276
rect 5172 9274 5196 9276
rect 5252 9274 5258 9276
rect 5012 9222 5014 9274
rect 5194 9222 5196 9274
rect 4950 9220 4956 9222
rect 5012 9220 5036 9222
rect 5092 9220 5116 9222
rect 5172 9220 5196 9222
rect 5252 9220 5258 9222
rect 4950 9211 5258 9220
rect 5368 8566 5396 9998
rect 5460 9586 5488 11766
rect 5610 10908 5918 10917
rect 5610 10906 5616 10908
rect 5672 10906 5696 10908
rect 5752 10906 5776 10908
rect 5832 10906 5856 10908
rect 5912 10906 5918 10908
rect 5672 10854 5674 10906
rect 5854 10854 5856 10906
rect 5610 10852 5616 10854
rect 5672 10852 5696 10854
rect 5752 10852 5776 10854
rect 5832 10852 5856 10854
rect 5912 10852 5918 10854
rect 5610 10843 5918 10852
rect 5610 9820 5918 9829
rect 5610 9818 5616 9820
rect 5672 9818 5696 9820
rect 5752 9818 5776 9820
rect 5832 9818 5856 9820
rect 5912 9818 5918 9820
rect 5672 9766 5674 9818
rect 5854 9766 5856 9818
rect 5610 9764 5616 9766
rect 5672 9764 5696 9766
rect 5752 9764 5776 9766
rect 5832 9764 5856 9766
rect 5912 9764 5918 9766
rect 5610 9755 5918 9764
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 6012 9110 6040 15302
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4816 8090 4844 8434
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 4950 8188 5258 8197
rect 4950 8186 4956 8188
rect 5012 8186 5036 8188
rect 5092 8186 5116 8188
rect 5172 8186 5196 8188
rect 5252 8186 5258 8188
rect 5012 8134 5014 8186
rect 5194 8134 5196 8186
rect 4950 8132 4956 8134
rect 5012 8132 5036 8134
rect 5092 8132 5116 8134
rect 5172 8132 5196 8134
rect 5252 8132 5258 8134
rect 4950 8123 5258 8132
rect 5368 8090 5396 8230
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5460 7954 5488 9046
rect 5610 8732 5918 8741
rect 5610 8730 5616 8732
rect 5672 8730 5696 8732
rect 5752 8730 5776 8732
rect 5832 8730 5856 8732
rect 5912 8730 5918 8732
rect 5672 8678 5674 8730
rect 5854 8678 5856 8730
rect 5610 8676 5616 8678
rect 5672 8676 5696 8678
rect 5752 8676 5776 8678
rect 5832 8676 5856 8678
rect 5912 8676 5918 8678
rect 5610 8667 5918 8676
rect 6012 8634 6040 9046
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4908 7410 4936 7686
rect 4896 7404 4948 7410
rect 4816 7364 4896 7392
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4816 6458 4844 7364
rect 4896 7346 4948 7352
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5368 7313 5396 7346
rect 5354 7304 5410 7313
rect 5552 7290 5580 8502
rect 6012 7886 6040 8570
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 5610 7644 5918 7653
rect 5610 7642 5616 7644
rect 5672 7642 5696 7644
rect 5752 7642 5776 7644
rect 5832 7642 5856 7644
rect 5912 7642 5918 7644
rect 5672 7590 5674 7642
rect 5854 7590 5856 7642
rect 5610 7588 5616 7590
rect 5672 7588 5696 7590
rect 5752 7588 5776 7590
rect 5832 7588 5856 7590
rect 5912 7588 5918 7590
rect 5610 7579 5918 7588
rect 6104 7410 6132 7686
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 5552 7262 5672 7290
rect 5354 7239 5410 7248
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 4950 7100 5258 7109
rect 4950 7098 4956 7100
rect 5012 7098 5036 7100
rect 5092 7098 5116 7100
rect 5172 7098 5196 7100
rect 5252 7098 5258 7100
rect 5012 7046 5014 7098
rect 5194 7046 5196 7098
rect 4950 7044 4956 7046
rect 5012 7044 5036 7046
rect 5092 7044 5116 7046
rect 5172 7044 5196 7046
rect 5252 7044 5258 7046
rect 4950 7035 5258 7044
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4724 5914 4752 6054
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 3884 5840 3936 5846
rect 3884 5782 3936 5788
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3528 4826 3556 5306
rect 3804 5302 3832 5714
rect 4712 5704 4764 5710
rect 4816 5692 4844 6394
rect 5000 6322 5028 6802
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5368 6458 5396 6666
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5460 6186 5488 6598
rect 5552 6186 5580 7142
rect 5644 6866 5672 7262
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5610 6556 5918 6565
rect 5610 6554 5616 6556
rect 5672 6554 5696 6556
rect 5752 6554 5776 6556
rect 5832 6554 5856 6556
rect 5912 6554 5918 6556
rect 5672 6502 5674 6554
rect 5854 6502 5856 6554
rect 5610 6500 5616 6502
rect 5672 6500 5696 6502
rect 5752 6500 5776 6502
rect 5832 6500 5856 6502
rect 5912 6500 5918 6502
rect 5610 6491 5918 6500
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5828 6186 5856 6394
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5816 6180 5868 6186
rect 5816 6122 5868 6128
rect 5460 6066 5488 6122
rect 5460 6038 5580 6066
rect 4950 6012 5258 6021
rect 4950 6010 4956 6012
rect 5012 6010 5036 6012
rect 5092 6010 5116 6012
rect 5172 6010 5196 6012
rect 5252 6010 5258 6012
rect 5012 5958 5014 6010
rect 5194 5958 5196 6010
rect 4950 5956 4956 5958
rect 5012 5956 5036 5958
rect 5092 5956 5116 5958
rect 5172 5956 5196 5958
rect 5252 5956 5258 5958
rect 4950 5947 5258 5956
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5276 5710 5304 5850
rect 4764 5664 4844 5692
rect 5264 5704 5316 5710
rect 4712 5646 4764 5652
rect 5264 5646 5316 5652
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4540 5370 4568 5510
rect 5276 5370 5304 5646
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 3252 3194 3280 4558
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4146 3372 4422
rect 3804 4146 3832 5238
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 4950 4924 5258 4933
rect 4950 4922 4956 4924
rect 5012 4922 5036 4924
rect 5092 4922 5116 4924
rect 5172 4922 5196 4924
rect 5252 4922 5258 4924
rect 5012 4870 5014 4922
rect 5194 4870 5196 4922
rect 4950 4868 4956 4870
rect 5012 4868 5036 4870
rect 5092 4868 5116 4870
rect 5172 4868 5196 4870
rect 5252 4868 5258 4870
rect 4950 4859 5258 4868
rect 5368 4196 5396 5170
rect 5552 4554 5580 6038
rect 6012 5914 6040 6734
rect 6104 6390 6132 7346
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6104 5778 6132 6326
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 5610 5468 5918 5477
rect 5610 5466 5616 5468
rect 5672 5466 5696 5468
rect 5752 5466 5776 5468
rect 5832 5466 5856 5468
rect 5912 5466 5918 5468
rect 5672 5414 5674 5466
rect 5854 5414 5856 5466
rect 5610 5412 5616 5414
rect 5672 5412 5696 5414
rect 5752 5412 5776 5414
rect 5832 5412 5856 5414
rect 5912 5412 5918 5414
rect 5610 5403 5918 5412
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4758 5764 4966
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 6104 4690 6132 5510
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 5828 4570 5856 4626
rect 5540 4548 5592 4554
rect 5828 4542 6040 4570
rect 5540 4490 5592 4496
rect 5448 4208 5500 4214
rect 5368 4168 5448 4196
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3344 3942 3372 4082
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3344 3534 3372 3878
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3712 3126 3740 3334
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 3804 2990 3832 4082
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3896 3738 3924 3878
rect 4950 3836 5258 3845
rect 4950 3834 4956 3836
rect 5012 3834 5036 3836
rect 5092 3834 5116 3836
rect 5172 3834 5196 3836
rect 5252 3834 5258 3836
rect 5012 3782 5014 3834
rect 5194 3782 5196 3834
rect 4950 3780 4956 3782
rect 5012 3780 5036 3782
rect 5092 3780 5116 3782
rect 5172 3780 5196 3782
rect 5252 3780 5258 3782
rect 4950 3771 5258 3780
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 5080 3528 5132 3534
rect 4066 3496 4122 3505
rect 5080 3470 5132 3476
rect 4066 3431 4122 3440
rect 4080 3398 4108 3431
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 4080 2446 4108 3334
rect 4448 3194 4476 3334
rect 5092 3194 5120 3470
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5368 2990 5396 4168
rect 5448 4150 5500 4156
rect 5552 4010 5580 4490
rect 5610 4380 5918 4389
rect 5610 4378 5616 4380
rect 5672 4378 5696 4380
rect 5752 4378 5776 4380
rect 5832 4378 5856 4380
rect 5912 4378 5918 4380
rect 5672 4326 5674 4378
rect 5854 4326 5856 4378
rect 5610 4324 5616 4326
rect 5672 4324 5696 4326
rect 5752 4324 5776 4326
rect 5832 4324 5856 4326
rect 5912 4324 5918 4326
rect 5610 4315 5918 4324
rect 6012 4214 6040 4542
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5552 3602 5580 3946
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5460 2990 5488 3470
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5552 3194 5580 3334
rect 5610 3292 5918 3301
rect 5610 3290 5616 3292
rect 5672 3290 5696 3292
rect 5752 3290 5776 3292
rect 5832 3290 5856 3292
rect 5912 3290 5918 3292
rect 5672 3238 5674 3290
rect 5854 3238 5856 3290
rect 5610 3236 5616 3238
rect 5672 3236 5696 3238
rect 5752 3236 5776 3238
rect 5832 3236 5856 3238
rect 5912 3236 5918 3238
rect 5610 3227 5918 3236
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 4950 2748 5258 2757
rect 4950 2746 4956 2748
rect 5012 2746 5036 2748
rect 5092 2746 5116 2748
rect 5172 2746 5196 2748
rect 5252 2746 5258 2748
rect 5012 2694 5014 2746
rect 5194 2694 5196 2746
rect 4950 2692 4956 2694
rect 5012 2692 5036 2694
rect 5092 2692 5116 2694
rect 5172 2692 5196 2694
rect 5252 2692 5258 2694
rect 4950 2683 5258 2692
rect 6012 2514 6040 4150
rect 6196 3738 6224 14962
rect 6288 12646 6316 15370
rect 6472 15162 6500 15370
rect 8220 15162 8248 15370
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 6748 13326 6776 13874
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 13394 6868 13806
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6932 13190 6960 13874
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7116 13394 7144 13670
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 6932 12782 6960 13126
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6288 10266 6316 12582
rect 7024 12434 7052 13126
rect 7208 12986 7236 13262
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12986 7328 13126
rect 7392 12986 7420 13330
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7300 12442 7328 12718
rect 7288 12436 7340 12442
rect 7024 12406 7236 12434
rect 7208 11762 7236 12406
rect 7288 12378 7340 12384
rect 7484 12374 7512 13874
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7484 11830 7512 12310
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 6748 11354 6776 11562
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 6380 10674 6408 11222
rect 6748 11150 6776 11290
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6288 7002 6316 9522
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6380 8974 6408 9386
rect 6564 9042 6592 9386
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6656 8430 6684 11018
rect 6748 9586 6776 11086
rect 6840 10606 6868 11562
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6932 10266 6960 10610
rect 7024 10606 7052 10950
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6840 9586 6868 9998
rect 6932 9722 6960 10066
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6656 8090 6684 8366
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6380 7002 6408 7686
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6288 6882 6316 6938
rect 6288 6854 6592 6882
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6380 5234 6408 6734
rect 6368 5228 6420 5234
rect 6288 5188 6368 5216
rect 6288 4826 6316 5188
rect 6368 5170 6420 5176
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6196 2774 6224 3674
rect 6380 2990 6408 4966
rect 6564 4078 6592 6854
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6748 6254 6776 6598
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6748 5642 6776 6190
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6840 5710 6868 5850
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6656 5250 6684 5510
rect 6748 5370 6776 5578
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6656 5222 6776 5250
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6472 3738 6500 4014
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6656 3602 6684 5102
rect 6748 4078 6776 5222
rect 6932 5166 6960 9318
rect 7024 9042 7052 10542
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7300 8498 7328 8774
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7300 7954 7328 8434
rect 7392 7954 7420 9522
rect 7576 9382 7604 10066
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7668 9178 7696 9862
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7300 6662 7328 7346
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7116 6118 7144 6190
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7116 5846 7144 6054
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 7300 5778 7328 6598
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7208 5166 7236 5646
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7208 4706 7236 5102
rect 7208 4690 7328 4706
rect 6828 4684 6880 4690
rect 7208 4684 7340 4690
rect 7208 4678 7288 4684
rect 6828 4626 6880 4632
rect 7288 4626 7340 4632
rect 6840 4146 6868 4626
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7012 4208 7064 4214
rect 7208 4162 7236 4558
rect 7300 4282 7328 4626
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7064 4156 7236 4162
rect 7012 4150 7236 4156
rect 6828 4140 6880 4146
rect 7024 4134 7236 4150
rect 7392 4146 7420 7890
rect 7484 6390 7512 8978
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7576 7546 7604 7822
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7562 7440 7618 7449
rect 7562 7375 7564 7384
rect 7616 7375 7618 7384
rect 7564 7346 7616 7352
rect 7576 7206 7604 7346
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5302 7880 6054
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7944 4826 7972 5714
rect 8036 5302 8064 6666
rect 8128 6662 8156 6870
rect 8220 6746 8248 14962
rect 8950 14716 9258 14725
rect 8950 14714 8956 14716
rect 9012 14714 9036 14716
rect 9092 14714 9116 14716
rect 9172 14714 9196 14716
rect 9252 14714 9258 14716
rect 9012 14662 9014 14714
rect 9194 14662 9196 14714
rect 8950 14660 8956 14662
rect 9012 14660 9036 14662
rect 9092 14660 9116 14662
rect 9172 14660 9196 14662
rect 9252 14660 9258 14662
rect 8950 14651 9258 14660
rect 8950 13628 9258 13637
rect 8950 13626 8956 13628
rect 9012 13626 9036 13628
rect 9092 13626 9116 13628
rect 9172 13626 9196 13628
rect 9252 13626 9258 13628
rect 9012 13574 9014 13626
rect 9194 13574 9196 13626
rect 8950 13572 8956 13574
rect 9012 13572 9036 13574
rect 9092 13572 9116 13574
rect 9172 13572 9196 13574
rect 9252 13572 9258 13574
rect 8950 13563 9258 13572
rect 9324 13530 9352 15438
rect 11612 15428 11664 15434
rect 11612 15370 11664 15376
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 14648 15428 14700 15434
rect 14648 15370 14700 15376
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 9610 15260 9918 15269
rect 9610 15258 9616 15260
rect 9672 15258 9696 15260
rect 9752 15258 9776 15260
rect 9832 15258 9856 15260
rect 9912 15258 9918 15260
rect 9672 15206 9674 15258
rect 9854 15206 9856 15258
rect 9610 15204 9616 15206
rect 9672 15204 9696 15206
rect 9752 15204 9776 15206
rect 9832 15204 9856 15206
rect 9912 15204 9918 15206
rect 9610 15195 9918 15204
rect 11624 14958 11652 15370
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 9610 14172 9918 14181
rect 9610 14170 9616 14172
rect 9672 14170 9696 14172
rect 9752 14170 9776 14172
rect 9832 14170 9856 14172
rect 9912 14170 9918 14172
rect 9672 14118 9674 14170
rect 9854 14118 9856 14170
rect 9610 14116 9616 14118
rect 9672 14116 9696 14118
rect 9752 14116 9776 14118
rect 9832 14116 9856 14118
rect 9912 14116 9918 14118
rect 9610 14107 9918 14116
rect 12820 13530 12848 15370
rect 13610 15260 13918 15269
rect 13610 15258 13616 15260
rect 13672 15258 13696 15260
rect 13752 15258 13776 15260
rect 13832 15258 13856 15260
rect 13912 15258 13918 15260
rect 13672 15206 13674 15258
rect 13854 15206 13856 15258
rect 13610 15204 13616 15206
rect 13672 15204 13696 15206
rect 13752 15204 13776 15206
rect 13832 15204 13856 15206
rect 13912 15204 13918 15206
rect 13610 15195 13918 15204
rect 14660 15162 14688 15370
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 15304 15026 15332 15370
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13610 14172 13918 14181
rect 13610 14170 13616 14172
rect 13672 14170 13696 14172
rect 13752 14170 13776 14172
rect 13832 14170 13856 14172
rect 13912 14170 13918 14172
rect 13672 14118 13674 14170
rect 13854 14118 13856 14170
rect 13610 14116 13616 14118
rect 13672 14116 13696 14118
rect 13752 14116 13776 14118
rect 13832 14116 13856 14118
rect 13912 14116 13918 14118
rect 13610 14107 13918 14116
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8680 12986 8708 13194
rect 9610 13084 9918 13093
rect 9610 13082 9616 13084
rect 9672 13082 9696 13084
rect 9752 13082 9776 13084
rect 9832 13082 9856 13084
rect 9912 13082 9918 13084
rect 9672 13030 9674 13082
rect 9854 13030 9856 13082
rect 9610 13028 9616 13030
rect 9672 13028 9696 13030
rect 9752 13028 9776 13030
rect 9832 13028 9856 13030
rect 9912 13028 9918 13030
rect 9610 13019 9918 13028
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8588 12442 8616 12786
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 11354 8524 11494
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8496 10724 8524 11018
rect 8576 10736 8628 10742
rect 8496 10696 8576 10724
rect 8576 10678 8628 10684
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8312 9450 8340 10610
rect 8680 9586 8708 12922
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9324 12730 9352 12786
rect 9324 12702 9444 12730
rect 9416 12646 9444 12702
rect 9128 12640 9180 12646
rect 9404 12640 9456 12646
rect 9180 12600 9352 12628
rect 9128 12582 9180 12588
rect 8950 12540 9258 12549
rect 8950 12538 8956 12540
rect 9012 12538 9036 12540
rect 9092 12538 9116 12540
rect 9172 12538 9196 12540
rect 9252 12538 9258 12540
rect 9012 12486 9014 12538
rect 9194 12486 9196 12538
rect 8950 12484 8956 12486
rect 9012 12484 9036 12486
rect 9092 12484 9116 12486
rect 9172 12484 9196 12486
rect 9252 12484 9258 12486
rect 8950 12475 9258 12484
rect 9324 12238 9352 12600
rect 9404 12582 9456 12588
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9508 11830 9536 12786
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 9610 11996 9918 12005
rect 9610 11994 9616 11996
rect 9672 11994 9696 11996
rect 9752 11994 9776 11996
rect 9832 11994 9856 11996
rect 9912 11994 9918 11996
rect 9672 11942 9674 11994
rect 9854 11942 9856 11994
rect 9610 11940 9616 11942
rect 9672 11940 9696 11942
rect 9752 11940 9776 11942
rect 9832 11940 9856 11942
rect 9912 11940 9918 11942
rect 9610 11931 9918 11940
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 8950 11452 9258 11461
rect 8950 11450 8956 11452
rect 9012 11450 9036 11452
rect 9092 11450 9116 11452
rect 9172 11450 9196 11452
rect 9252 11450 9258 11452
rect 9012 11398 9014 11450
rect 9194 11398 9196 11450
rect 8950 11396 8956 11398
rect 9012 11396 9036 11398
rect 9092 11396 9116 11398
rect 9172 11396 9196 11398
rect 9252 11396 9258 11398
rect 8950 11387 9258 11396
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 10266 8892 10406
rect 8950 10364 9258 10373
rect 8950 10362 8956 10364
rect 9012 10362 9036 10364
rect 9092 10362 9116 10364
rect 9172 10362 9196 10364
rect 9252 10362 9258 10364
rect 9012 10310 9014 10362
rect 9194 10310 9196 10362
rect 8950 10308 8956 10310
rect 9012 10308 9036 10310
rect 9092 10308 9116 10310
rect 9172 10308 9196 10310
rect 9252 10308 9258 10310
rect 8950 10299 9258 10308
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8772 8498 8800 8978
rect 8760 8492 8812 8498
rect 8864 8480 8892 9590
rect 8950 9276 9258 9285
rect 8950 9274 8956 9276
rect 9012 9274 9036 9276
rect 9092 9274 9116 9276
rect 9172 9274 9196 9276
rect 9252 9274 9258 9276
rect 9012 9222 9014 9274
rect 9194 9222 9196 9274
rect 8950 9220 8956 9222
rect 9012 9220 9036 9222
rect 9092 9220 9116 9222
rect 9172 9220 9196 9222
rect 9252 9220 9258 9222
rect 8950 9211 9258 9220
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8956 8634 8984 8910
rect 9232 8634 9260 9046
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9324 8514 9352 10746
rect 9416 10742 9444 11086
rect 9404 10736 9456 10742
rect 9404 10678 9456 10684
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9416 10266 9444 10542
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9508 10146 9536 11766
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9610 10908 9918 10917
rect 9610 10906 9616 10908
rect 9672 10906 9696 10908
rect 9752 10906 9776 10908
rect 9832 10906 9856 10908
rect 9912 10906 9918 10908
rect 9672 10854 9674 10906
rect 9854 10854 9856 10906
rect 9610 10852 9616 10854
rect 9672 10852 9696 10854
rect 9752 10852 9776 10854
rect 9832 10852 9856 10854
rect 9912 10852 9918 10854
rect 9610 10843 9918 10852
rect 9968 10674 9996 10950
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10060 10538 10088 11766
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 10152 10266 10180 12106
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 9416 10118 9536 10146
rect 9416 9654 9444 10118
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9416 8974 9444 9590
rect 9508 9178 9536 9998
rect 9610 9820 9918 9829
rect 9610 9818 9616 9820
rect 9672 9818 9696 9820
rect 9752 9818 9776 9820
rect 9832 9818 9856 9820
rect 9912 9818 9918 9820
rect 9672 9766 9674 9818
rect 9854 9766 9856 9818
rect 9610 9764 9616 9766
rect 9672 9764 9696 9766
rect 9752 9764 9776 9766
rect 9832 9764 9856 9766
rect 9912 9764 9918 9766
rect 9610 9755 9918 9764
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 10060 9042 10088 9386
rect 10244 9382 10272 13398
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10428 11354 10456 12038
rect 10612 11354 10640 12854
rect 10888 12850 10916 13262
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 11440 12986 11468 13194
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 10888 12306 10916 12786
rect 11716 12442 11744 12786
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11808 12646 11836 12718
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10324 11280 10376 11286
rect 10324 11222 10376 11228
rect 10336 10606 10364 11222
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10336 10130 10364 10542
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9772 8968 9824 8974
rect 10152 8922 10180 8978
rect 9824 8916 10180 8922
rect 9772 8910 10180 8916
rect 9784 8894 10180 8910
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 9610 8732 9918 8741
rect 9610 8730 9616 8732
rect 9672 8730 9696 8732
rect 9752 8730 9776 8732
rect 9832 8730 9856 8732
rect 9912 8730 9918 8732
rect 9672 8678 9674 8730
rect 9854 8678 9856 8730
rect 9610 8676 9616 8678
rect 9672 8676 9696 8678
rect 9752 8676 9776 8678
rect 9832 8676 9856 8678
rect 9912 8676 9918 8678
rect 9610 8667 9918 8676
rect 10152 8566 10180 8774
rect 9140 8498 9352 8514
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 8944 8492 8996 8498
rect 8864 8452 8944 8480
rect 8760 8434 8812 8440
rect 8944 8434 8996 8440
rect 9128 8492 9352 8498
rect 9180 8486 9352 8492
rect 9404 8492 9456 8498
rect 9128 8434 9180 8440
rect 9404 8434 9456 8440
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 8668 8288 8720 8294
rect 9048 8276 9076 8366
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 8720 8248 9076 8276
rect 8668 8230 8720 8236
rect 8950 8188 9258 8197
rect 8950 8186 8956 8188
rect 9012 8186 9036 8188
rect 9092 8186 9116 8188
rect 9172 8186 9196 8188
rect 9252 8186 9258 8188
rect 9012 8134 9014 8186
rect 9194 8134 9196 8186
rect 8950 8132 8956 8134
rect 9012 8132 9036 8134
rect 9092 8132 9116 8134
rect 9172 8132 9196 8134
rect 9252 8132 9258 8134
rect 8950 8123 9258 8132
rect 9324 7834 9352 8298
rect 9232 7806 9352 7834
rect 9232 7478 9260 7806
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 8950 7100 9258 7109
rect 8950 7098 8956 7100
rect 9012 7098 9036 7100
rect 9092 7098 9116 7100
rect 9172 7098 9196 7100
rect 9252 7098 9258 7100
rect 9012 7046 9014 7098
rect 9194 7046 9196 7098
rect 8950 7044 8956 7046
rect 9012 7044 9036 7046
rect 9092 7044 9116 7046
rect 9172 7044 9196 7046
rect 9252 7044 9258 7046
rect 8950 7035 9258 7044
rect 9324 7002 9352 7686
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9416 6882 9444 8434
rect 10152 7886 10180 8502
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 9610 7644 9918 7653
rect 9610 7642 9616 7644
rect 9672 7642 9696 7644
rect 9752 7642 9776 7644
rect 9832 7642 9856 7644
rect 9912 7642 9918 7644
rect 9672 7590 9674 7642
rect 9854 7590 9856 7642
rect 9610 7588 9616 7590
rect 9672 7588 9696 7590
rect 9752 7588 9776 7590
rect 9832 7588 9856 7590
rect 9912 7588 9918 7590
rect 9610 7579 9918 7588
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9324 6854 9444 6882
rect 8760 6792 8812 6798
rect 8220 6718 8340 6746
rect 8760 6734 8812 6740
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8128 6322 8156 6598
rect 8220 6390 8248 6598
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8312 6118 8340 6718
rect 8772 6458 8800 6734
rect 9324 6458 9352 6854
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8036 4706 8064 5238
rect 8312 4826 8340 6054
rect 8950 6012 9258 6021
rect 8950 6010 8956 6012
rect 9012 6010 9036 6012
rect 9092 6010 9116 6012
rect 9172 6010 9196 6012
rect 9252 6010 9258 6012
rect 9012 5958 9014 6010
rect 9194 5958 9196 6010
rect 8950 5956 8956 5958
rect 9012 5956 9036 5958
rect 9092 5956 9116 5958
rect 9172 5956 9196 5958
rect 9252 5956 9258 5958
rect 8950 5947 9258 5956
rect 9416 5778 9444 6598
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8404 5370 8432 5510
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 7760 4678 8064 4706
rect 8404 4690 8432 5306
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8300 4684 8352 4690
rect 7760 4622 7788 4678
rect 8300 4626 8352 4632
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 7380 4140 7432 4146
rect 6828 4082 6880 4088
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6196 2746 6316 2774
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6288 2446 6316 2746
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 7116 2378 7144 4134
rect 7380 4082 7432 4088
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7208 3738 7236 3946
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7208 3194 7236 3334
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7300 2514 7328 2790
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7392 2310 7420 4082
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7852 2650 7880 3402
rect 8036 3398 8064 3878
rect 8128 3738 8156 4490
rect 8312 3738 8340 4626
rect 8404 4282 8432 4626
rect 8588 4622 8616 4762
rect 8576 4616 8628 4622
rect 8864 4604 8892 4966
rect 8950 4924 9258 4933
rect 8950 4922 8956 4924
rect 9012 4922 9036 4924
rect 9092 4922 9116 4924
rect 9172 4922 9196 4924
rect 9252 4922 9258 4924
rect 9012 4870 9014 4922
rect 9194 4870 9196 4922
rect 8950 4868 8956 4870
rect 9012 4868 9036 4870
rect 9092 4868 9116 4870
rect 9172 4868 9196 4870
rect 9252 4868 9258 4870
rect 8950 4859 9258 4868
rect 9324 4690 9352 4966
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9036 4616 9088 4622
rect 8864 4576 9036 4604
rect 8576 4558 8628 4564
rect 9036 4558 9088 4564
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8404 3602 8432 4082
rect 8588 4078 8616 4558
rect 9416 4078 9444 5714
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 8036 3194 8064 3334
rect 8588 3194 8616 3878
rect 8950 3836 9258 3845
rect 8950 3834 8956 3836
rect 9012 3834 9036 3836
rect 9092 3834 9116 3836
rect 9172 3834 9196 3836
rect 9252 3834 9258 3836
rect 9012 3782 9014 3834
rect 9194 3782 9196 3834
rect 8950 3780 8956 3782
rect 9012 3780 9036 3782
rect 9092 3780 9116 3782
rect 9172 3780 9196 3782
rect 9252 3780 9258 3782
rect 8950 3771 9258 3780
rect 9416 3194 9444 4014
rect 9508 3466 9536 7346
rect 9968 6866 9996 7822
rect 10060 7410 10088 7822
rect 10152 7410 10180 7822
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9610 6556 9918 6565
rect 9610 6554 9616 6556
rect 9672 6554 9696 6556
rect 9752 6554 9776 6556
rect 9832 6554 9856 6556
rect 9912 6554 9918 6556
rect 9672 6502 9674 6554
rect 9854 6502 9856 6554
rect 9610 6500 9616 6502
rect 9672 6500 9696 6502
rect 9752 6500 9776 6502
rect 9832 6500 9856 6502
rect 9912 6500 9918 6502
rect 9610 6491 9918 6500
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9600 5794 9628 6054
rect 10336 5914 10364 9930
rect 10428 8430 10456 10678
rect 10612 10062 10640 10950
rect 10980 10470 11008 12174
rect 11348 11694 11376 12242
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11348 11218 11376 11630
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11256 10810 11284 11018
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10796 10266 10824 10406
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10428 7886 10456 8366
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10428 7410 10456 7822
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 9600 5778 9720 5794
rect 9600 5772 9732 5778
rect 9600 5766 9680 5772
rect 9680 5714 9732 5720
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9610 5468 9918 5477
rect 9610 5466 9616 5468
rect 9672 5466 9696 5468
rect 9752 5466 9776 5468
rect 9832 5466 9856 5468
rect 9912 5466 9918 5468
rect 9672 5414 9674 5466
rect 9854 5414 9856 5466
rect 9610 5412 9616 5414
rect 9672 5412 9696 5414
rect 9752 5412 9776 5414
rect 9832 5412 9856 5414
rect 9912 5412 9918 5414
rect 9610 5403 9918 5412
rect 9968 5370 9996 5510
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10336 5166 10364 5850
rect 10428 5710 10456 6802
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10520 6458 10548 6734
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 9610 4380 9918 4389
rect 9610 4378 9616 4380
rect 9672 4378 9696 4380
rect 9752 4378 9776 4380
rect 9832 4378 9856 4380
rect 9912 4378 9918 4380
rect 9672 4326 9674 4378
rect 9854 4326 9856 4378
rect 9610 4324 9616 4326
rect 9672 4324 9696 4326
rect 9752 4324 9776 4326
rect 9832 4324 9856 4326
rect 9912 4324 9918 4326
rect 9610 4315 9918 4324
rect 9968 4282 9996 4422
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 10152 3942 10180 4422
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9692 3398 9720 3674
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9610 3292 9918 3301
rect 9610 3290 9616 3292
rect 9672 3290 9696 3292
rect 9752 3290 9776 3292
rect 9832 3290 9856 3292
rect 9912 3290 9918 3292
rect 9672 3238 9674 3290
rect 9854 3238 9856 3290
rect 9610 3236 9616 3238
rect 9672 3236 9696 3238
rect 9752 3236 9776 3238
rect 9832 3236 9856 3238
rect 9912 3236 9918 3238
rect 9610 3227 9918 3236
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9128 3120 9180 3126
rect 9128 3062 9180 3068
rect 9140 2854 9168 3062
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9968 2774 9996 3334
rect 10336 3126 10364 4694
rect 10428 4078 10456 5646
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10428 3194 10456 4014
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10428 2854 10456 3130
rect 10520 3058 10548 4490
rect 10612 3534 10640 9998
rect 11348 9926 11376 11154
rect 11440 11014 11468 11630
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11624 10538 11652 10678
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11520 10532 11572 10538
rect 11520 10474 11572 10480
rect 11612 10532 11664 10538
rect 11612 10474 11664 10480
rect 11532 10266 11560 10474
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11256 9722 11284 9862
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11348 8974 11376 9862
rect 11532 9042 11560 9862
rect 11624 9042 11652 10474
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11716 8974 11744 10542
rect 11808 9382 11836 12582
rect 12256 12368 12308 12374
rect 12256 12310 12308 12316
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12268 12238 12296 12310
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12544 11898 12572 12310
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 10810 12112 10950
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 12268 10742 12296 11630
rect 12636 11354 12664 12106
rect 12728 11778 12756 13194
rect 12820 12238 12848 13466
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 13610 13084 13918 13093
rect 13610 13082 13616 13084
rect 13672 13082 13696 13084
rect 13752 13082 13776 13084
rect 13832 13082 13856 13084
rect 13912 13082 13918 13084
rect 13672 13030 13674 13082
rect 13854 13030 13856 13082
rect 13610 13028 13616 13030
rect 13672 13028 13696 13030
rect 13752 13028 13776 13030
rect 13832 13028 13856 13030
rect 13912 13028 13918 13030
rect 13610 13019 13918 13028
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13832 12238 13860 12582
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 12728 11750 12848 11778
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12268 9110 12296 9318
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10888 8362 10916 8842
rect 11348 8634 11376 8910
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11440 8566 11468 8842
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10704 7002 10732 7414
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10704 6458 10732 6938
rect 10888 6866 10916 8298
rect 10980 7206 11008 8434
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11072 8022 11100 8230
rect 11440 8090 11468 8502
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10980 5710 11008 7142
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10888 5166 10916 5510
rect 10876 5160 10928 5166
rect 10928 5120 11008 5148
rect 10876 5102 10928 5108
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10796 3942 10824 4558
rect 10784 3936 10836 3942
rect 10704 3896 10784 3924
rect 10704 3602 10732 3896
rect 10784 3878 10836 3884
rect 10888 3738 10916 4558
rect 10980 4486 11008 5120
rect 11072 4690 11100 6870
rect 11164 6730 11192 7278
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11256 6798 11284 7210
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11164 5914 11192 6666
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11164 4826 11192 5102
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11440 4758 11468 8026
rect 11532 7886 11560 8774
rect 11716 8294 11744 8910
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11716 7834 11744 8230
rect 11716 7806 11836 7834
rect 11900 7818 11928 8910
rect 12452 8820 12480 10610
rect 12544 9042 12572 10950
rect 12636 10470 12664 11290
rect 12728 10538 12756 11562
rect 12820 11234 12848 11750
rect 13464 11694 13492 12038
rect 13610 11996 13918 12005
rect 13610 11994 13616 11996
rect 13672 11994 13696 11996
rect 13752 11994 13776 11996
rect 13832 11994 13856 11996
rect 13912 11994 13918 11996
rect 13672 11942 13674 11994
rect 13854 11942 13856 11994
rect 13610 11940 13616 11942
rect 13672 11940 13696 11942
rect 13752 11940 13776 11942
rect 13832 11940 13856 11942
rect 13912 11940 13918 11942
rect 13610 11931 13918 11940
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12820 11206 12940 11234
rect 12912 11014 12940 11206
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12820 10810 12848 10950
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12912 10690 12940 10950
rect 13372 10742 13400 11494
rect 12820 10662 12940 10690
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 12716 10532 12768 10538
rect 12716 10474 12768 10480
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12820 10062 12848 10662
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13464 10248 13492 11630
rect 13610 10908 13918 10917
rect 13610 10906 13616 10908
rect 13672 10906 13696 10908
rect 13752 10906 13776 10908
rect 13832 10906 13856 10908
rect 13912 10906 13918 10908
rect 13672 10854 13674 10906
rect 13854 10854 13856 10906
rect 13610 10852 13616 10854
rect 13672 10852 13696 10854
rect 13752 10852 13776 10854
rect 13832 10852 13856 10854
rect 13912 10852 13918 10854
rect 13610 10843 13918 10852
rect 14016 10810 14044 13126
rect 15304 12986 15332 14962
rect 15580 12986 15608 15370
rect 16500 15162 16528 16351
rect 17420 15638 17448 17200
rect 17408 15632 17460 15638
rect 17408 15574 17460 15580
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15948 12986 15976 14282
rect 16132 13410 16160 14962
rect 16946 14376 17002 14385
rect 16946 14311 16948 14320
rect 17000 14311 17002 14320
rect 16948 14282 17000 14288
rect 16040 13382 16160 13410
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14108 11354 14136 11766
rect 14200 11558 14228 12378
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14292 11898 14320 12106
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 15028 11762 15056 12038
rect 15120 11898 15148 12786
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13280 10220 13492 10248
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 13280 9654 13308 10220
rect 13556 10010 13584 10406
rect 13372 9982 13584 10010
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13372 9586 13400 9982
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 12636 9178 12664 9522
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12820 9382 12848 9454
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12532 8832 12584 8838
rect 12452 8792 12532 8820
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11808 7750 11836 7806
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11716 7546 11744 7686
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11900 7342 11928 7754
rect 11992 7546 12020 7958
rect 12452 7954 12480 8792
rect 12532 8774 12584 8780
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11992 6934 12020 7482
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12452 7002 12480 7278
rect 12544 7206 12572 8026
rect 12820 7750 12848 9318
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 13372 8634 13400 9522
rect 13464 9500 13492 9862
rect 13610 9820 13918 9829
rect 13610 9818 13616 9820
rect 13672 9818 13696 9820
rect 13752 9818 13776 9820
rect 13832 9818 13856 9820
rect 13912 9818 13918 9820
rect 13672 9766 13674 9818
rect 13854 9766 13856 9818
rect 13610 9764 13616 9766
rect 13672 9764 13696 9766
rect 13752 9764 13776 9766
rect 13832 9764 13856 9766
rect 13912 9764 13918 9766
rect 13610 9755 13918 9764
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13648 9518 13676 9590
rect 13544 9512 13596 9518
rect 13464 9472 13544 9500
rect 13544 9454 13596 9460
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13648 8922 13676 9454
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13832 9330 13860 9454
rect 14200 9330 14228 11494
rect 14844 11150 14872 11630
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14844 10470 14872 11086
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14844 10266 14872 10406
rect 14936 10266 14964 10610
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 13740 8974 13768 9318
rect 13832 9302 14228 9330
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 13464 8894 13676 8922
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13372 8498 13400 8570
rect 13464 8514 13492 8894
rect 13610 8732 13918 8741
rect 13610 8730 13616 8732
rect 13672 8730 13696 8732
rect 13752 8730 13776 8732
rect 13832 8730 13856 8732
rect 13912 8730 13918 8732
rect 13672 8678 13674 8730
rect 13854 8678 13856 8730
rect 13610 8676 13616 8678
rect 13672 8676 13696 8678
rect 13752 8676 13776 8678
rect 13832 8676 13856 8678
rect 13912 8676 13918 8678
rect 13610 8667 13918 8676
rect 14016 8634 14044 9114
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13464 8486 13768 8514
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 13464 8090 13492 8486
rect 13740 8430 13768 8486
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13648 8090 13676 8366
rect 14200 8294 14228 9302
rect 14384 9178 14412 9454
rect 14568 9382 14596 9930
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13372 7750 13400 7822
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4826 11560 4966
rect 12360 4826 12388 6190
rect 12452 6118 12480 6938
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12544 4758 12572 7142
rect 12636 7002 12664 7686
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12820 6882 12848 7142
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12820 6866 12940 6882
rect 12820 6860 12952 6866
rect 12820 6854 12900 6860
rect 12900 6802 12952 6808
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12636 5370 12664 6598
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4282 11928 4422
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 12452 3942 12480 4558
rect 12636 4078 12664 5102
rect 12728 4826 12756 6054
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12820 4706 12848 5306
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 12728 4678 12848 4706
rect 13004 4690 13032 4762
rect 12992 4684 13044 4690
rect 12728 4146 12756 4678
rect 12992 4626 13044 4632
rect 13004 4434 13032 4626
rect 13372 4622 13400 7686
rect 13610 7644 13918 7653
rect 13610 7642 13616 7644
rect 13672 7642 13696 7644
rect 13752 7642 13776 7644
rect 13832 7642 13856 7644
rect 13912 7642 13918 7644
rect 13672 7590 13674 7642
rect 13854 7590 13856 7642
rect 13610 7588 13616 7590
rect 13672 7588 13696 7590
rect 13752 7588 13776 7590
rect 13832 7588 13856 7590
rect 13912 7588 13918 7590
rect 13610 7579 13918 7588
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13464 6662 13492 7414
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13556 6662 13584 6938
rect 14016 6798 14044 7278
rect 14108 6798 14136 7686
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13610 6556 13918 6565
rect 13610 6554 13616 6556
rect 13672 6554 13696 6556
rect 13752 6554 13776 6556
rect 13832 6554 13856 6556
rect 13912 6554 13918 6556
rect 13672 6502 13674 6554
rect 13854 6502 13856 6554
rect 13610 6500 13616 6502
rect 13672 6500 13696 6502
rect 13752 6500 13776 6502
rect 13832 6500 13856 6502
rect 13912 6500 13918 6502
rect 13610 6491 13918 6500
rect 14016 5914 14044 6734
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 13464 5166 13492 5850
rect 13610 5468 13918 5477
rect 13610 5466 13616 5468
rect 13672 5466 13696 5468
rect 13752 5466 13776 5468
rect 13832 5466 13856 5468
rect 13912 5466 13918 5468
rect 13672 5414 13674 5466
rect 13854 5414 13856 5466
rect 13610 5412 13616 5414
rect 13672 5412 13696 5414
rect 13752 5412 13776 5414
rect 13832 5412 13856 5414
rect 13912 5412 13918 5414
rect 13610 5403 13918 5412
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13004 4406 13400 4434
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10888 3602 10916 3674
rect 12452 3670 12480 3878
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10704 3398 10732 3538
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10612 3194 10640 3334
rect 10704 3194 10732 3334
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10980 3126 11008 3470
rect 11348 3176 11376 3470
rect 11428 3392 11480 3398
rect 11428 3334 11480 3340
rect 11164 3148 11376 3176
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 8950 2748 9258 2757
rect 8950 2746 8956 2748
rect 9012 2746 9036 2748
rect 9092 2746 9116 2748
rect 9172 2746 9196 2748
rect 9252 2746 9258 2748
rect 9012 2694 9014 2746
rect 9194 2694 9196 2746
rect 8950 2692 8956 2694
rect 9012 2692 9036 2694
rect 9092 2692 9116 2694
rect 9172 2692 9196 2694
rect 9252 2692 9258 2694
rect 8950 2683 9258 2692
rect 9876 2746 9996 2774
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 9876 2446 9904 2746
rect 10888 2446 10916 2790
rect 11164 2582 11192 3148
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11348 2446 11376 2790
rect 11440 2446 11468 3334
rect 12728 3126 12756 4082
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13372 3466 13400 4406
rect 13464 4078 13492 5102
rect 14200 4758 14228 8230
rect 14660 7954 14688 8570
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14844 7342 14872 7686
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 13610 4380 13918 4389
rect 13610 4378 13616 4380
rect 13672 4378 13696 4380
rect 13752 4378 13776 4380
rect 13832 4378 13856 4380
rect 13912 4378 13918 4380
rect 13672 4326 13674 4378
rect 13854 4326 13856 4378
rect 13610 4324 13616 4326
rect 13672 4324 13696 4326
rect 13752 4324 13776 4326
rect 13832 4324 13856 4326
rect 13912 4324 13918 4326
rect 13610 4315 13918 4324
rect 14108 4214 14136 4422
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12452 2650 12480 2926
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12820 2530 12848 3402
rect 13464 3058 13492 4014
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 13610 3292 13918 3301
rect 13610 3290 13616 3292
rect 13672 3290 13696 3292
rect 13752 3290 13776 3292
rect 13832 3290 13856 3292
rect 13912 3290 13918 3292
rect 13672 3238 13674 3290
rect 13854 3238 13856 3290
rect 13610 3236 13616 3238
rect 13672 3236 13696 3238
rect 13752 3236 13776 3238
rect 13832 3236 13856 3238
rect 13912 3236 13918 3238
rect 13610 3227 13918 3236
rect 14476 3194 14504 3334
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 15028 2774 15056 11698
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15120 10810 15148 11018
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15396 10742 15424 12106
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15396 10062 15424 10678
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15396 9654 15424 9998
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15212 8090 15240 8230
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15580 7886 15608 8978
rect 15764 8634 15792 12786
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 16040 6322 16068 13382
rect 16120 13252 16172 13258
rect 16120 13194 16172 13200
rect 16132 12986 16160 13194
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16960 13025 16988 13126
rect 16946 13016 17002 13025
rect 16120 12980 16172 12986
rect 16946 12951 17002 12960
rect 16120 12922 16172 12928
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16500 10985 16528 11154
rect 16486 10976 16542 10985
rect 16486 10911 16542 10920
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16132 8974 16160 9318
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16762 8936 16818 8945
rect 16762 8871 16764 8880
rect 16816 8871 16818 8880
rect 16764 8842 16816 8848
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16132 7206 16160 8434
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16776 7585 16804 7686
rect 16762 7576 16818 7585
rect 16762 7511 16818 7520
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 16132 4622 16160 7142
rect 16488 5568 16540 5574
rect 16486 5536 16488 5545
rect 16540 5536 16542 5545
rect 16486 5471 16542 5480
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16776 4185 16804 4422
rect 16762 4176 16818 4185
rect 16762 4111 16818 4120
rect 15936 3528 15988 3534
rect 15658 3496 15714 3505
rect 15936 3470 15988 3476
rect 15658 3431 15714 3440
rect 15672 3058 15700 3431
rect 15948 3194 15976 3470
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16040 3194 16068 3334
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 15028 2746 15148 2774
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 12820 2502 12940 2530
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 1610 2204 1918 2213
rect 1610 2202 1616 2204
rect 1672 2202 1696 2204
rect 1752 2202 1776 2204
rect 1832 2202 1856 2204
rect 1912 2202 1918 2204
rect 1672 2150 1674 2202
rect 1854 2150 1856 2202
rect 1610 2148 1616 2150
rect 1672 2148 1696 2150
rect 1752 2148 1776 2150
rect 1832 2148 1856 2150
rect 1912 2148 1918 2150
rect 1610 2139 1918 2148
rect 3252 800 3280 2246
rect 4540 800 4568 2246
rect 5610 2204 5918 2213
rect 5610 2202 5616 2204
rect 5672 2202 5696 2204
rect 5752 2202 5776 2204
rect 5832 2202 5856 2204
rect 5912 2202 5918 2204
rect 5672 2150 5674 2202
rect 5854 2150 5856 2202
rect 5610 2148 5616 2150
rect 5672 2148 5696 2150
rect 5752 2148 5776 2150
rect 5832 2148 5856 2150
rect 5912 2148 5918 2150
rect 5610 2139 5918 2148
rect 6472 800 6500 2246
rect 8404 800 8432 2246
rect 9610 2204 9918 2213
rect 9610 2202 9616 2204
rect 9672 2202 9696 2204
rect 9752 2202 9776 2204
rect 9832 2202 9856 2204
rect 9912 2202 9918 2204
rect 9672 2150 9674 2202
rect 9854 2150 9856 2202
rect 9610 2148 9616 2150
rect 9672 2148 9696 2150
rect 9752 2148 9776 2150
rect 9832 2148 9856 2150
rect 9912 2148 9918 2150
rect 9610 2139 9918 2148
rect 9692 870 9812 898
rect 9692 800 9720 870
rect 18 0 74 800
rect 1306 0 1362 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 9784 762 9812 870
rect 9968 762 9996 2246
rect 11624 800 11652 2246
rect 12912 800 12940 2502
rect 15120 2446 15148 2746
rect 15764 2446 15792 2790
rect 15948 2650 15976 3130
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 13610 2204 13918 2213
rect 13610 2202 13616 2204
rect 13672 2202 13696 2204
rect 13752 2202 13776 2204
rect 13832 2202 13856 2204
rect 13912 2202 13918 2204
rect 13672 2150 13674 2202
rect 13854 2150 13856 2202
rect 13610 2148 13616 2150
rect 13672 2148 13696 2150
rect 13752 2148 13776 2150
rect 13832 2148 13856 2150
rect 13912 2148 13918 2150
rect 13610 2139 13918 2148
rect 14844 800 14872 2246
rect 9784 734 9996 762
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 14830 0 14886 800
rect 16408 105 16436 2246
rect 16776 800 16804 2790
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 16960 2145 16988 2314
rect 16946 2136 17002 2145
rect 16946 2071 17002 2080
rect 16394 96 16450 105
rect 16394 31 16450 40
rect 16762 0 16818 800
<< via2 >>
rect 1490 17720 1546 17776
rect 1398 15952 1454 16008
rect 956 15802 1012 15804
rect 1036 15802 1092 15804
rect 1116 15802 1172 15804
rect 1196 15802 1252 15804
rect 956 15750 1002 15802
rect 1002 15750 1012 15802
rect 1036 15750 1066 15802
rect 1066 15750 1078 15802
rect 1078 15750 1092 15802
rect 1116 15750 1130 15802
rect 1130 15750 1142 15802
rect 1142 15750 1172 15802
rect 1196 15750 1206 15802
rect 1206 15750 1252 15802
rect 956 15748 1012 15750
rect 1036 15748 1092 15750
rect 1116 15748 1172 15750
rect 1196 15748 1252 15750
rect 4956 15802 5012 15804
rect 5036 15802 5092 15804
rect 5116 15802 5172 15804
rect 5196 15802 5252 15804
rect 4956 15750 5002 15802
rect 5002 15750 5012 15802
rect 5036 15750 5066 15802
rect 5066 15750 5078 15802
rect 5078 15750 5092 15802
rect 5116 15750 5130 15802
rect 5130 15750 5142 15802
rect 5142 15750 5172 15802
rect 5196 15750 5206 15802
rect 5206 15750 5252 15802
rect 4956 15748 5012 15750
rect 5036 15748 5092 15750
rect 5116 15748 5172 15750
rect 5196 15748 5252 15750
rect 8956 15802 9012 15804
rect 9036 15802 9092 15804
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 8956 15750 9002 15802
rect 9002 15750 9012 15802
rect 9036 15750 9066 15802
rect 9066 15750 9078 15802
rect 9078 15750 9092 15802
rect 9116 15750 9130 15802
rect 9130 15750 9142 15802
rect 9142 15750 9172 15802
rect 9196 15750 9206 15802
rect 9206 15750 9252 15802
rect 8956 15748 9012 15750
rect 9036 15748 9092 15750
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 16486 16360 16542 16416
rect 1616 15258 1672 15260
rect 1696 15258 1752 15260
rect 1776 15258 1832 15260
rect 1856 15258 1912 15260
rect 1616 15206 1662 15258
rect 1662 15206 1672 15258
rect 1696 15206 1726 15258
rect 1726 15206 1738 15258
rect 1738 15206 1752 15258
rect 1776 15206 1790 15258
rect 1790 15206 1802 15258
rect 1802 15206 1832 15258
rect 1856 15206 1866 15258
rect 1866 15206 1912 15258
rect 1616 15204 1672 15206
rect 1696 15204 1752 15206
rect 1776 15204 1832 15206
rect 1856 15204 1912 15206
rect 956 14714 1012 14716
rect 1036 14714 1092 14716
rect 1116 14714 1172 14716
rect 1196 14714 1252 14716
rect 956 14662 1002 14714
rect 1002 14662 1012 14714
rect 1036 14662 1066 14714
rect 1066 14662 1078 14714
rect 1078 14662 1092 14714
rect 1116 14662 1130 14714
rect 1130 14662 1142 14714
rect 1142 14662 1172 14714
rect 1196 14662 1206 14714
rect 1206 14662 1252 14714
rect 956 14660 1012 14662
rect 1036 14660 1092 14662
rect 1116 14660 1172 14662
rect 1196 14660 1252 14662
rect 1616 14170 1672 14172
rect 1696 14170 1752 14172
rect 1776 14170 1832 14172
rect 1856 14170 1912 14172
rect 1616 14118 1662 14170
rect 1662 14118 1672 14170
rect 1696 14118 1726 14170
rect 1726 14118 1738 14170
rect 1738 14118 1752 14170
rect 1776 14118 1790 14170
rect 1790 14118 1802 14170
rect 1802 14118 1832 14170
rect 1856 14118 1866 14170
rect 1866 14118 1912 14170
rect 1616 14116 1672 14118
rect 1696 14116 1752 14118
rect 1776 14116 1832 14118
rect 1856 14116 1912 14118
rect 1398 13640 1454 13696
rect 956 13626 1012 13628
rect 1036 13626 1092 13628
rect 1116 13626 1172 13628
rect 1196 13626 1252 13628
rect 956 13574 1002 13626
rect 1002 13574 1012 13626
rect 1036 13574 1066 13626
rect 1066 13574 1078 13626
rect 1078 13574 1092 13626
rect 1116 13574 1130 13626
rect 1130 13574 1142 13626
rect 1142 13574 1172 13626
rect 1196 13574 1206 13626
rect 1206 13574 1252 13626
rect 956 13572 1012 13574
rect 1036 13572 1092 13574
rect 1116 13572 1172 13574
rect 1196 13572 1252 13574
rect 1616 13082 1672 13084
rect 1696 13082 1752 13084
rect 1776 13082 1832 13084
rect 1856 13082 1912 13084
rect 1616 13030 1662 13082
rect 1662 13030 1672 13082
rect 1696 13030 1726 13082
rect 1726 13030 1738 13082
rect 1738 13030 1752 13082
rect 1776 13030 1790 13082
rect 1790 13030 1802 13082
rect 1802 13030 1832 13082
rect 1856 13030 1866 13082
rect 1866 13030 1912 13082
rect 1616 13028 1672 13030
rect 1696 13028 1752 13030
rect 1776 13028 1832 13030
rect 1856 13028 1912 13030
rect 956 12538 1012 12540
rect 1036 12538 1092 12540
rect 1116 12538 1172 12540
rect 1196 12538 1252 12540
rect 956 12486 1002 12538
rect 1002 12486 1012 12538
rect 1036 12486 1066 12538
rect 1066 12486 1078 12538
rect 1078 12486 1092 12538
rect 1116 12486 1130 12538
rect 1130 12486 1142 12538
rect 1142 12486 1172 12538
rect 1196 12486 1206 12538
rect 1206 12486 1252 12538
rect 956 12484 1012 12486
rect 1036 12484 1092 12486
rect 1116 12484 1172 12486
rect 1196 12484 1252 12486
rect 1490 12280 1546 12336
rect 5616 15258 5672 15260
rect 5696 15258 5752 15260
rect 5776 15258 5832 15260
rect 5856 15258 5912 15260
rect 5616 15206 5662 15258
rect 5662 15206 5672 15258
rect 5696 15206 5726 15258
rect 5726 15206 5738 15258
rect 5738 15206 5752 15258
rect 5776 15206 5790 15258
rect 5790 15206 5802 15258
rect 5802 15206 5832 15258
rect 5856 15206 5866 15258
rect 5866 15206 5912 15258
rect 5616 15204 5672 15206
rect 5696 15204 5752 15206
rect 5776 15204 5832 15206
rect 5856 15204 5912 15206
rect 1616 11994 1672 11996
rect 1696 11994 1752 11996
rect 1776 11994 1832 11996
rect 1856 11994 1912 11996
rect 1616 11942 1662 11994
rect 1662 11942 1672 11994
rect 1696 11942 1726 11994
rect 1726 11942 1738 11994
rect 1738 11942 1752 11994
rect 1776 11942 1790 11994
rect 1790 11942 1802 11994
rect 1802 11942 1832 11994
rect 1856 11942 1866 11994
rect 1866 11942 1912 11994
rect 1616 11940 1672 11942
rect 1696 11940 1752 11942
rect 1776 11940 1832 11942
rect 1856 11940 1912 11942
rect 956 11450 1012 11452
rect 1036 11450 1092 11452
rect 1116 11450 1172 11452
rect 1196 11450 1252 11452
rect 956 11398 1002 11450
rect 1002 11398 1012 11450
rect 1036 11398 1066 11450
rect 1066 11398 1078 11450
rect 1078 11398 1092 11450
rect 1116 11398 1130 11450
rect 1130 11398 1142 11450
rect 1142 11398 1172 11450
rect 1196 11398 1206 11450
rect 1206 11398 1252 11450
rect 956 11396 1012 11398
rect 1036 11396 1092 11398
rect 1116 11396 1172 11398
rect 1196 11396 1252 11398
rect 1616 10906 1672 10908
rect 1696 10906 1752 10908
rect 1776 10906 1832 10908
rect 1856 10906 1912 10908
rect 1616 10854 1662 10906
rect 1662 10854 1672 10906
rect 1696 10854 1726 10906
rect 1726 10854 1738 10906
rect 1738 10854 1752 10906
rect 1776 10854 1790 10906
rect 1790 10854 1802 10906
rect 1802 10854 1832 10906
rect 1856 10854 1866 10906
rect 1866 10854 1912 10906
rect 1616 10852 1672 10854
rect 1696 10852 1752 10854
rect 1776 10852 1832 10854
rect 1856 10852 1912 10854
rect 956 10362 1012 10364
rect 1036 10362 1092 10364
rect 1116 10362 1172 10364
rect 1196 10362 1252 10364
rect 956 10310 1002 10362
rect 1002 10310 1012 10362
rect 1036 10310 1066 10362
rect 1066 10310 1078 10362
rect 1078 10310 1092 10362
rect 1116 10310 1130 10362
rect 1130 10310 1142 10362
rect 1142 10310 1172 10362
rect 1196 10310 1206 10362
rect 1206 10310 1252 10362
rect 956 10308 1012 10310
rect 1036 10308 1092 10310
rect 1116 10308 1172 10310
rect 1196 10308 1252 10310
rect 938 10104 994 10160
rect 1616 9818 1672 9820
rect 1696 9818 1752 9820
rect 1776 9818 1832 9820
rect 1856 9818 1912 9820
rect 1616 9766 1662 9818
rect 1662 9766 1672 9818
rect 1696 9766 1726 9818
rect 1726 9766 1738 9818
rect 1738 9766 1752 9818
rect 1776 9766 1790 9818
rect 1790 9766 1802 9818
rect 1802 9766 1832 9818
rect 1856 9766 1866 9818
rect 1866 9766 1912 9818
rect 1616 9764 1672 9766
rect 1696 9764 1752 9766
rect 1776 9764 1832 9766
rect 1856 9764 1912 9766
rect 956 9274 1012 9276
rect 1036 9274 1092 9276
rect 1116 9274 1172 9276
rect 1196 9274 1252 9276
rect 956 9222 1002 9274
rect 1002 9222 1012 9274
rect 1036 9222 1066 9274
rect 1066 9222 1078 9274
rect 1078 9222 1092 9274
rect 1116 9222 1130 9274
rect 1130 9222 1142 9274
rect 1142 9222 1172 9274
rect 1196 9222 1206 9274
rect 1206 9222 1252 9274
rect 956 9220 1012 9222
rect 1036 9220 1092 9222
rect 1116 9220 1172 9222
rect 1196 9220 1252 9222
rect 938 8900 994 8936
rect 938 8880 940 8900
rect 940 8880 992 8900
rect 992 8880 994 8900
rect 956 8186 1012 8188
rect 1036 8186 1092 8188
rect 1116 8186 1172 8188
rect 1196 8186 1252 8188
rect 956 8134 1002 8186
rect 1002 8134 1012 8186
rect 1036 8134 1066 8186
rect 1066 8134 1078 8186
rect 1078 8134 1092 8186
rect 1116 8134 1130 8186
rect 1130 8134 1142 8186
rect 1142 8134 1172 8186
rect 1196 8134 1206 8186
rect 1206 8134 1252 8186
rect 956 8132 1012 8134
rect 1036 8132 1092 8134
rect 1116 8132 1172 8134
rect 1196 8132 1252 8134
rect 4956 14714 5012 14716
rect 5036 14714 5092 14716
rect 5116 14714 5172 14716
rect 5196 14714 5252 14716
rect 4956 14662 5002 14714
rect 5002 14662 5012 14714
rect 5036 14662 5066 14714
rect 5066 14662 5078 14714
rect 5078 14662 5092 14714
rect 5116 14662 5130 14714
rect 5130 14662 5142 14714
rect 5142 14662 5172 14714
rect 5196 14662 5206 14714
rect 5206 14662 5252 14714
rect 4956 14660 5012 14662
rect 5036 14660 5092 14662
rect 5116 14660 5172 14662
rect 5196 14660 5252 14662
rect 5616 14170 5672 14172
rect 5696 14170 5752 14172
rect 5776 14170 5832 14172
rect 5856 14170 5912 14172
rect 5616 14118 5662 14170
rect 5662 14118 5672 14170
rect 5696 14118 5726 14170
rect 5726 14118 5738 14170
rect 5738 14118 5752 14170
rect 5776 14118 5790 14170
rect 5790 14118 5802 14170
rect 5802 14118 5832 14170
rect 5856 14118 5866 14170
rect 5866 14118 5912 14170
rect 5616 14116 5672 14118
rect 5696 14116 5752 14118
rect 5776 14116 5832 14118
rect 5856 14116 5912 14118
rect 1616 8730 1672 8732
rect 1696 8730 1752 8732
rect 1776 8730 1832 8732
rect 1856 8730 1912 8732
rect 1616 8678 1662 8730
rect 1662 8678 1672 8730
rect 1696 8678 1726 8730
rect 1726 8678 1738 8730
rect 1738 8678 1752 8730
rect 1776 8678 1790 8730
rect 1790 8678 1802 8730
rect 1802 8678 1832 8730
rect 1856 8678 1866 8730
rect 1866 8678 1912 8730
rect 1616 8676 1672 8678
rect 1696 8676 1752 8678
rect 1776 8676 1832 8678
rect 1856 8676 1912 8678
rect 1616 7642 1672 7644
rect 1696 7642 1752 7644
rect 1776 7642 1832 7644
rect 1856 7642 1912 7644
rect 1616 7590 1662 7642
rect 1662 7590 1672 7642
rect 1696 7590 1726 7642
rect 1726 7590 1738 7642
rect 1738 7590 1752 7642
rect 1776 7590 1790 7642
rect 1790 7590 1802 7642
rect 1802 7590 1832 7642
rect 1856 7590 1866 7642
rect 1866 7590 1912 7642
rect 1616 7588 1672 7590
rect 1696 7588 1752 7590
rect 1776 7588 1832 7590
rect 1856 7588 1912 7590
rect 956 7098 1012 7100
rect 1036 7098 1092 7100
rect 1116 7098 1172 7100
rect 1196 7098 1252 7100
rect 956 7046 1002 7098
rect 1002 7046 1012 7098
rect 1036 7046 1066 7098
rect 1066 7046 1078 7098
rect 1078 7046 1092 7098
rect 1116 7046 1130 7098
rect 1130 7046 1142 7098
rect 1142 7046 1172 7098
rect 1196 7046 1206 7098
rect 1206 7046 1252 7098
rect 956 7044 1012 7046
rect 1036 7044 1092 7046
rect 1116 7044 1172 7046
rect 1196 7044 1252 7046
rect 938 6840 994 6896
rect 956 6010 1012 6012
rect 1036 6010 1092 6012
rect 1116 6010 1172 6012
rect 1196 6010 1252 6012
rect 956 5958 1002 6010
rect 1002 5958 1012 6010
rect 1036 5958 1066 6010
rect 1066 5958 1078 6010
rect 1078 5958 1092 6010
rect 1116 5958 1130 6010
rect 1130 5958 1142 6010
rect 1142 5958 1172 6010
rect 1196 5958 1206 6010
rect 1206 5958 1252 6010
rect 956 5956 1012 5958
rect 1036 5956 1092 5958
rect 1116 5956 1172 5958
rect 1196 5956 1252 5958
rect 1616 6554 1672 6556
rect 1696 6554 1752 6556
rect 1776 6554 1832 6556
rect 1856 6554 1912 6556
rect 1616 6502 1662 6554
rect 1662 6502 1672 6554
rect 1696 6502 1726 6554
rect 1726 6502 1738 6554
rect 1738 6502 1752 6554
rect 1776 6502 1790 6554
rect 1790 6502 1802 6554
rect 1802 6502 1832 6554
rect 1856 6502 1866 6554
rect 1866 6502 1912 6554
rect 1616 6500 1672 6502
rect 1696 6500 1752 6502
rect 1776 6500 1832 6502
rect 1856 6500 1912 6502
rect 1616 5466 1672 5468
rect 1696 5466 1752 5468
rect 1776 5466 1832 5468
rect 1856 5466 1912 5468
rect 1616 5414 1662 5466
rect 1662 5414 1672 5466
rect 1696 5414 1726 5466
rect 1726 5414 1738 5466
rect 1738 5414 1752 5466
rect 1776 5414 1790 5466
rect 1790 5414 1802 5466
rect 1802 5414 1832 5466
rect 1856 5414 1866 5466
rect 1866 5414 1912 5466
rect 1616 5412 1672 5414
rect 1696 5412 1752 5414
rect 1776 5412 1832 5414
rect 1856 5412 1912 5414
rect 754 5072 810 5128
rect 956 4922 1012 4924
rect 1036 4922 1092 4924
rect 1116 4922 1172 4924
rect 1196 4922 1252 4924
rect 956 4870 1002 4922
rect 1002 4870 1012 4922
rect 1036 4870 1066 4922
rect 1066 4870 1078 4922
rect 1078 4870 1092 4922
rect 1116 4870 1130 4922
rect 1130 4870 1142 4922
rect 1142 4870 1172 4922
rect 1196 4870 1206 4922
rect 1206 4870 1252 4922
rect 956 4868 1012 4870
rect 1036 4868 1092 4870
rect 1116 4868 1172 4870
rect 1196 4868 1252 4870
rect 1616 4378 1672 4380
rect 1696 4378 1752 4380
rect 1776 4378 1832 4380
rect 1856 4378 1912 4380
rect 1616 4326 1662 4378
rect 1662 4326 1672 4378
rect 1696 4326 1726 4378
rect 1726 4326 1738 4378
rect 1738 4326 1752 4378
rect 1776 4326 1790 4378
rect 1790 4326 1802 4378
rect 1802 4326 1832 4378
rect 1856 4326 1866 4378
rect 1866 4326 1912 4378
rect 1616 4324 1672 4326
rect 1696 4324 1752 4326
rect 1776 4324 1832 4326
rect 1856 4324 1912 4326
rect 956 3834 1012 3836
rect 1036 3834 1092 3836
rect 1116 3834 1172 3836
rect 1196 3834 1252 3836
rect 956 3782 1002 3834
rect 1002 3782 1012 3834
rect 1036 3782 1066 3834
rect 1066 3782 1078 3834
rect 1078 3782 1092 3834
rect 1116 3782 1130 3834
rect 1130 3782 1142 3834
rect 1142 3782 1172 3834
rect 1196 3782 1206 3834
rect 1206 3782 1252 3834
rect 956 3780 1012 3782
rect 1036 3780 1092 3782
rect 1116 3780 1172 3782
rect 1196 3780 1252 3782
rect 938 3460 994 3496
rect 938 3440 940 3460
rect 940 3440 992 3460
rect 992 3440 994 3460
rect 1616 3290 1672 3292
rect 1696 3290 1752 3292
rect 1776 3290 1832 3292
rect 1856 3290 1912 3292
rect 1616 3238 1662 3290
rect 1662 3238 1672 3290
rect 1696 3238 1726 3290
rect 1726 3238 1738 3290
rect 1738 3238 1752 3290
rect 1776 3238 1790 3290
rect 1790 3238 1802 3290
rect 1802 3238 1832 3290
rect 1856 3238 1866 3290
rect 1866 3238 1912 3290
rect 1616 3236 1672 3238
rect 1696 3236 1752 3238
rect 1776 3236 1832 3238
rect 1856 3236 1912 3238
rect 956 2746 1012 2748
rect 1036 2746 1092 2748
rect 1116 2746 1172 2748
rect 1196 2746 1252 2748
rect 956 2694 1002 2746
rect 1002 2694 1012 2746
rect 1036 2694 1066 2746
rect 1066 2694 1078 2746
rect 1078 2694 1092 2746
rect 1116 2694 1130 2746
rect 1130 2694 1142 2746
rect 1142 2694 1172 2746
rect 1196 2694 1206 2746
rect 1206 2694 1252 2746
rect 956 2692 1012 2694
rect 1036 2692 1092 2694
rect 1116 2692 1172 2694
rect 1196 2692 1252 2694
rect 938 1400 994 1456
rect 4956 13626 5012 13628
rect 5036 13626 5092 13628
rect 5116 13626 5172 13628
rect 5196 13626 5252 13628
rect 4956 13574 5002 13626
rect 5002 13574 5012 13626
rect 5036 13574 5066 13626
rect 5066 13574 5078 13626
rect 5078 13574 5092 13626
rect 5116 13574 5130 13626
rect 5130 13574 5142 13626
rect 5142 13574 5172 13626
rect 5196 13574 5206 13626
rect 5206 13574 5252 13626
rect 4956 13572 5012 13574
rect 5036 13572 5092 13574
rect 5116 13572 5172 13574
rect 5196 13572 5252 13574
rect 5616 13082 5672 13084
rect 5696 13082 5752 13084
rect 5776 13082 5832 13084
rect 5856 13082 5912 13084
rect 5616 13030 5662 13082
rect 5662 13030 5672 13082
rect 5696 13030 5726 13082
rect 5726 13030 5738 13082
rect 5738 13030 5752 13082
rect 5776 13030 5790 13082
rect 5790 13030 5802 13082
rect 5802 13030 5832 13082
rect 5856 13030 5866 13082
rect 5866 13030 5912 13082
rect 5616 13028 5672 13030
rect 5696 13028 5752 13030
rect 5776 13028 5832 13030
rect 5856 13028 5912 13030
rect 4956 12538 5012 12540
rect 5036 12538 5092 12540
rect 5116 12538 5172 12540
rect 5196 12538 5252 12540
rect 4956 12486 5002 12538
rect 5002 12486 5012 12538
rect 5036 12486 5066 12538
rect 5066 12486 5078 12538
rect 5078 12486 5092 12538
rect 5116 12486 5130 12538
rect 5130 12486 5142 12538
rect 5142 12486 5172 12538
rect 5196 12486 5206 12538
rect 5206 12486 5252 12538
rect 4956 12484 5012 12486
rect 5036 12484 5092 12486
rect 5116 12484 5172 12486
rect 5196 12484 5252 12486
rect 4956 11450 5012 11452
rect 5036 11450 5092 11452
rect 5116 11450 5172 11452
rect 5196 11450 5252 11452
rect 4956 11398 5002 11450
rect 5002 11398 5012 11450
rect 5036 11398 5066 11450
rect 5066 11398 5078 11450
rect 5078 11398 5092 11450
rect 5116 11398 5130 11450
rect 5130 11398 5142 11450
rect 5142 11398 5172 11450
rect 5196 11398 5206 11450
rect 5206 11398 5252 11450
rect 4956 11396 5012 11398
rect 5036 11396 5092 11398
rect 5116 11396 5172 11398
rect 5196 11396 5252 11398
rect 3422 7248 3478 7304
rect 4526 7384 4582 7440
rect 5616 11994 5672 11996
rect 5696 11994 5752 11996
rect 5776 11994 5832 11996
rect 5856 11994 5912 11996
rect 5616 11942 5662 11994
rect 5662 11942 5672 11994
rect 5696 11942 5726 11994
rect 5726 11942 5738 11994
rect 5738 11942 5752 11994
rect 5776 11942 5790 11994
rect 5790 11942 5802 11994
rect 5802 11942 5832 11994
rect 5856 11942 5866 11994
rect 5866 11942 5912 11994
rect 5616 11940 5672 11942
rect 5696 11940 5752 11942
rect 5776 11940 5832 11942
rect 5856 11940 5912 11942
rect 4956 10362 5012 10364
rect 5036 10362 5092 10364
rect 5116 10362 5172 10364
rect 5196 10362 5252 10364
rect 4956 10310 5002 10362
rect 5002 10310 5012 10362
rect 5036 10310 5066 10362
rect 5066 10310 5078 10362
rect 5078 10310 5092 10362
rect 5116 10310 5130 10362
rect 5130 10310 5142 10362
rect 5142 10310 5172 10362
rect 5196 10310 5206 10362
rect 5206 10310 5252 10362
rect 4956 10308 5012 10310
rect 5036 10308 5092 10310
rect 5116 10308 5172 10310
rect 5196 10308 5252 10310
rect 4956 9274 5012 9276
rect 5036 9274 5092 9276
rect 5116 9274 5172 9276
rect 5196 9274 5252 9276
rect 4956 9222 5002 9274
rect 5002 9222 5012 9274
rect 5036 9222 5066 9274
rect 5066 9222 5078 9274
rect 5078 9222 5092 9274
rect 5116 9222 5130 9274
rect 5130 9222 5142 9274
rect 5142 9222 5172 9274
rect 5196 9222 5206 9274
rect 5206 9222 5252 9274
rect 4956 9220 5012 9222
rect 5036 9220 5092 9222
rect 5116 9220 5172 9222
rect 5196 9220 5252 9222
rect 5616 10906 5672 10908
rect 5696 10906 5752 10908
rect 5776 10906 5832 10908
rect 5856 10906 5912 10908
rect 5616 10854 5662 10906
rect 5662 10854 5672 10906
rect 5696 10854 5726 10906
rect 5726 10854 5738 10906
rect 5738 10854 5752 10906
rect 5776 10854 5790 10906
rect 5790 10854 5802 10906
rect 5802 10854 5832 10906
rect 5856 10854 5866 10906
rect 5866 10854 5912 10906
rect 5616 10852 5672 10854
rect 5696 10852 5752 10854
rect 5776 10852 5832 10854
rect 5856 10852 5912 10854
rect 5616 9818 5672 9820
rect 5696 9818 5752 9820
rect 5776 9818 5832 9820
rect 5856 9818 5912 9820
rect 5616 9766 5662 9818
rect 5662 9766 5672 9818
rect 5696 9766 5726 9818
rect 5726 9766 5738 9818
rect 5738 9766 5752 9818
rect 5776 9766 5790 9818
rect 5790 9766 5802 9818
rect 5802 9766 5832 9818
rect 5856 9766 5866 9818
rect 5866 9766 5912 9818
rect 5616 9764 5672 9766
rect 5696 9764 5752 9766
rect 5776 9764 5832 9766
rect 5856 9764 5912 9766
rect 4956 8186 5012 8188
rect 5036 8186 5092 8188
rect 5116 8186 5172 8188
rect 5196 8186 5252 8188
rect 4956 8134 5002 8186
rect 5002 8134 5012 8186
rect 5036 8134 5066 8186
rect 5066 8134 5078 8186
rect 5078 8134 5092 8186
rect 5116 8134 5130 8186
rect 5130 8134 5142 8186
rect 5142 8134 5172 8186
rect 5196 8134 5206 8186
rect 5206 8134 5252 8186
rect 4956 8132 5012 8134
rect 5036 8132 5092 8134
rect 5116 8132 5172 8134
rect 5196 8132 5252 8134
rect 5616 8730 5672 8732
rect 5696 8730 5752 8732
rect 5776 8730 5832 8732
rect 5856 8730 5912 8732
rect 5616 8678 5662 8730
rect 5662 8678 5672 8730
rect 5696 8678 5726 8730
rect 5726 8678 5738 8730
rect 5738 8678 5752 8730
rect 5776 8678 5790 8730
rect 5790 8678 5802 8730
rect 5802 8678 5832 8730
rect 5856 8678 5866 8730
rect 5866 8678 5912 8730
rect 5616 8676 5672 8678
rect 5696 8676 5752 8678
rect 5776 8676 5832 8678
rect 5856 8676 5912 8678
rect 5354 7248 5410 7304
rect 5616 7642 5672 7644
rect 5696 7642 5752 7644
rect 5776 7642 5832 7644
rect 5856 7642 5912 7644
rect 5616 7590 5662 7642
rect 5662 7590 5672 7642
rect 5696 7590 5726 7642
rect 5726 7590 5738 7642
rect 5738 7590 5752 7642
rect 5776 7590 5790 7642
rect 5790 7590 5802 7642
rect 5802 7590 5832 7642
rect 5856 7590 5866 7642
rect 5866 7590 5912 7642
rect 5616 7588 5672 7590
rect 5696 7588 5752 7590
rect 5776 7588 5832 7590
rect 5856 7588 5912 7590
rect 4956 7098 5012 7100
rect 5036 7098 5092 7100
rect 5116 7098 5172 7100
rect 5196 7098 5252 7100
rect 4956 7046 5002 7098
rect 5002 7046 5012 7098
rect 5036 7046 5066 7098
rect 5066 7046 5078 7098
rect 5078 7046 5092 7098
rect 5116 7046 5130 7098
rect 5130 7046 5142 7098
rect 5142 7046 5172 7098
rect 5196 7046 5206 7098
rect 5206 7046 5252 7098
rect 4956 7044 5012 7046
rect 5036 7044 5092 7046
rect 5116 7044 5172 7046
rect 5196 7044 5252 7046
rect 5616 6554 5672 6556
rect 5696 6554 5752 6556
rect 5776 6554 5832 6556
rect 5856 6554 5912 6556
rect 5616 6502 5662 6554
rect 5662 6502 5672 6554
rect 5696 6502 5726 6554
rect 5726 6502 5738 6554
rect 5738 6502 5752 6554
rect 5776 6502 5790 6554
rect 5790 6502 5802 6554
rect 5802 6502 5832 6554
rect 5856 6502 5866 6554
rect 5866 6502 5912 6554
rect 5616 6500 5672 6502
rect 5696 6500 5752 6502
rect 5776 6500 5832 6502
rect 5856 6500 5912 6502
rect 4956 6010 5012 6012
rect 5036 6010 5092 6012
rect 5116 6010 5172 6012
rect 5196 6010 5252 6012
rect 4956 5958 5002 6010
rect 5002 5958 5012 6010
rect 5036 5958 5066 6010
rect 5066 5958 5078 6010
rect 5078 5958 5092 6010
rect 5116 5958 5130 6010
rect 5130 5958 5142 6010
rect 5142 5958 5172 6010
rect 5196 5958 5206 6010
rect 5206 5958 5252 6010
rect 4956 5956 5012 5958
rect 5036 5956 5092 5958
rect 5116 5956 5172 5958
rect 5196 5956 5252 5958
rect 4956 4922 5012 4924
rect 5036 4922 5092 4924
rect 5116 4922 5172 4924
rect 5196 4922 5252 4924
rect 4956 4870 5002 4922
rect 5002 4870 5012 4922
rect 5036 4870 5066 4922
rect 5066 4870 5078 4922
rect 5078 4870 5092 4922
rect 5116 4870 5130 4922
rect 5130 4870 5142 4922
rect 5142 4870 5172 4922
rect 5196 4870 5206 4922
rect 5206 4870 5252 4922
rect 4956 4868 5012 4870
rect 5036 4868 5092 4870
rect 5116 4868 5172 4870
rect 5196 4868 5252 4870
rect 5616 5466 5672 5468
rect 5696 5466 5752 5468
rect 5776 5466 5832 5468
rect 5856 5466 5912 5468
rect 5616 5414 5662 5466
rect 5662 5414 5672 5466
rect 5696 5414 5726 5466
rect 5726 5414 5738 5466
rect 5738 5414 5752 5466
rect 5776 5414 5790 5466
rect 5790 5414 5802 5466
rect 5802 5414 5832 5466
rect 5856 5414 5866 5466
rect 5866 5414 5912 5466
rect 5616 5412 5672 5414
rect 5696 5412 5752 5414
rect 5776 5412 5832 5414
rect 5856 5412 5912 5414
rect 4956 3834 5012 3836
rect 5036 3834 5092 3836
rect 5116 3834 5172 3836
rect 5196 3834 5252 3836
rect 4956 3782 5002 3834
rect 5002 3782 5012 3834
rect 5036 3782 5066 3834
rect 5066 3782 5078 3834
rect 5078 3782 5092 3834
rect 5116 3782 5130 3834
rect 5130 3782 5142 3834
rect 5142 3782 5172 3834
rect 5196 3782 5206 3834
rect 5206 3782 5252 3834
rect 4956 3780 5012 3782
rect 5036 3780 5092 3782
rect 5116 3780 5172 3782
rect 5196 3780 5252 3782
rect 4066 3440 4122 3496
rect 5616 4378 5672 4380
rect 5696 4378 5752 4380
rect 5776 4378 5832 4380
rect 5856 4378 5912 4380
rect 5616 4326 5662 4378
rect 5662 4326 5672 4378
rect 5696 4326 5726 4378
rect 5726 4326 5738 4378
rect 5738 4326 5752 4378
rect 5776 4326 5790 4378
rect 5790 4326 5802 4378
rect 5802 4326 5832 4378
rect 5856 4326 5866 4378
rect 5866 4326 5912 4378
rect 5616 4324 5672 4326
rect 5696 4324 5752 4326
rect 5776 4324 5832 4326
rect 5856 4324 5912 4326
rect 5616 3290 5672 3292
rect 5696 3290 5752 3292
rect 5776 3290 5832 3292
rect 5856 3290 5912 3292
rect 5616 3238 5662 3290
rect 5662 3238 5672 3290
rect 5696 3238 5726 3290
rect 5726 3238 5738 3290
rect 5738 3238 5752 3290
rect 5776 3238 5790 3290
rect 5790 3238 5802 3290
rect 5802 3238 5832 3290
rect 5856 3238 5866 3290
rect 5866 3238 5912 3290
rect 5616 3236 5672 3238
rect 5696 3236 5752 3238
rect 5776 3236 5832 3238
rect 5856 3236 5912 3238
rect 4956 2746 5012 2748
rect 5036 2746 5092 2748
rect 5116 2746 5172 2748
rect 5196 2746 5252 2748
rect 4956 2694 5002 2746
rect 5002 2694 5012 2746
rect 5036 2694 5066 2746
rect 5066 2694 5078 2746
rect 5078 2694 5092 2746
rect 5116 2694 5130 2746
rect 5130 2694 5142 2746
rect 5142 2694 5172 2746
rect 5196 2694 5206 2746
rect 5206 2694 5252 2746
rect 4956 2692 5012 2694
rect 5036 2692 5092 2694
rect 5116 2692 5172 2694
rect 5196 2692 5252 2694
rect 7562 7404 7618 7440
rect 7562 7384 7564 7404
rect 7564 7384 7616 7404
rect 7616 7384 7618 7404
rect 8956 14714 9012 14716
rect 9036 14714 9092 14716
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 8956 14662 9002 14714
rect 9002 14662 9012 14714
rect 9036 14662 9066 14714
rect 9066 14662 9078 14714
rect 9078 14662 9092 14714
rect 9116 14662 9130 14714
rect 9130 14662 9142 14714
rect 9142 14662 9172 14714
rect 9196 14662 9206 14714
rect 9206 14662 9252 14714
rect 8956 14660 9012 14662
rect 9036 14660 9092 14662
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 8956 13626 9012 13628
rect 9036 13626 9092 13628
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 8956 13574 9002 13626
rect 9002 13574 9012 13626
rect 9036 13574 9066 13626
rect 9066 13574 9078 13626
rect 9078 13574 9092 13626
rect 9116 13574 9130 13626
rect 9130 13574 9142 13626
rect 9142 13574 9172 13626
rect 9196 13574 9206 13626
rect 9206 13574 9252 13626
rect 8956 13572 9012 13574
rect 9036 13572 9092 13574
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 9616 15258 9672 15260
rect 9696 15258 9752 15260
rect 9776 15258 9832 15260
rect 9856 15258 9912 15260
rect 9616 15206 9662 15258
rect 9662 15206 9672 15258
rect 9696 15206 9726 15258
rect 9726 15206 9738 15258
rect 9738 15206 9752 15258
rect 9776 15206 9790 15258
rect 9790 15206 9802 15258
rect 9802 15206 9832 15258
rect 9856 15206 9866 15258
rect 9866 15206 9912 15258
rect 9616 15204 9672 15206
rect 9696 15204 9752 15206
rect 9776 15204 9832 15206
rect 9856 15204 9912 15206
rect 9616 14170 9672 14172
rect 9696 14170 9752 14172
rect 9776 14170 9832 14172
rect 9856 14170 9912 14172
rect 9616 14118 9662 14170
rect 9662 14118 9672 14170
rect 9696 14118 9726 14170
rect 9726 14118 9738 14170
rect 9738 14118 9752 14170
rect 9776 14118 9790 14170
rect 9790 14118 9802 14170
rect 9802 14118 9832 14170
rect 9856 14118 9866 14170
rect 9866 14118 9912 14170
rect 9616 14116 9672 14118
rect 9696 14116 9752 14118
rect 9776 14116 9832 14118
rect 9856 14116 9912 14118
rect 13616 15258 13672 15260
rect 13696 15258 13752 15260
rect 13776 15258 13832 15260
rect 13856 15258 13912 15260
rect 13616 15206 13662 15258
rect 13662 15206 13672 15258
rect 13696 15206 13726 15258
rect 13726 15206 13738 15258
rect 13738 15206 13752 15258
rect 13776 15206 13790 15258
rect 13790 15206 13802 15258
rect 13802 15206 13832 15258
rect 13856 15206 13866 15258
rect 13866 15206 13912 15258
rect 13616 15204 13672 15206
rect 13696 15204 13752 15206
rect 13776 15204 13832 15206
rect 13856 15204 13912 15206
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 13616 14170 13672 14172
rect 13696 14170 13752 14172
rect 13776 14170 13832 14172
rect 13856 14170 13912 14172
rect 13616 14118 13662 14170
rect 13662 14118 13672 14170
rect 13696 14118 13726 14170
rect 13726 14118 13738 14170
rect 13738 14118 13752 14170
rect 13776 14118 13790 14170
rect 13790 14118 13802 14170
rect 13802 14118 13832 14170
rect 13856 14118 13866 14170
rect 13866 14118 13912 14170
rect 13616 14116 13672 14118
rect 13696 14116 13752 14118
rect 13776 14116 13832 14118
rect 13856 14116 13912 14118
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 9616 13082 9672 13084
rect 9696 13082 9752 13084
rect 9776 13082 9832 13084
rect 9856 13082 9912 13084
rect 9616 13030 9662 13082
rect 9662 13030 9672 13082
rect 9696 13030 9726 13082
rect 9726 13030 9738 13082
rect 9738 13030 9752 13082
rect 9776 13030 9790 13082
rect 9790 13030 9802 13082
rect 9802 13030 9832 13082
rect 9856 13030 9866 13082
rect 9866 13030 9912 13082
rect 9616 13028 9672 13030
rect 9696 13028 9752 13030
rect 9776 13028 9832 13030
rect 9856 13028 9912 13030
rect 8956 12538 9012 12540
rect 9036 12538 9092 12540
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 8956 12486 9002 12538
rect 9002 12486 9012 12538
rect 9036 12486 9066 12538
rect 9066 12486 9078 12538
rect 9078 12486 9092 12538
rect 9116 12486 9130 12538
rect 9130 12486 9142 12538
rect 9142 12486 9172 12538
rect 9196 12486 9206 12538
rect 9206 12486 9252 12538
rect 8956 12484 9012 12486
rect 9036 12484 9092 12486
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 9616 11994 9672 11996
rect 9696 11994 9752 11996
rect 9776 11994 9832 11996
rect 9856 11994 9912 11996
rect 9616 11942 9662 11994
rect 9662 11942 9672 11994
rect 9696 11942 9726 11994
rect 9726 11942 9738 11994
rect 9738 11942 9752 11994
rect 9776 11942 9790 11994
rect 9790 11942 9802 11994
rect 9802 11942 9832 11994
rect 9856 11942 9866 11994
rect 9866 11942 9912 11994
rect 9616 11940 9672 11942
rect 9696 11940 9752 11942
rect 9776 11940 9832 11942
rect 9856 11940 9912 11942
rect 8956 11450 9012 11452
rect 9036 11450 9092 11452
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 8956 11398 9002 11450
rect 9002 11398 9012 11450
rect 9036 11398 9066 11450
rect 9066 11398 9078 11450
rect 9078 11398 9092 11450
rect 9116 11398 9130 11450
rect 9130 11398 9142 11450
rect 9142 11398 9172 11450
rect 9196 11398 9206 11450
rect 9206 11398 9252 11450
rect 8956 11396 9012 11398
rect 9036 11396 9092 11398
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 8956 10362 9012 10364
rect 9036 10362 9092 10364
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 8956 10310 9002 10362
rect 9002 10310 9012 10362
rect 9036 10310 9066 10362
rect 9066 10310 9078 10362
rect 9078 10310 9092 10362
rect 9116 10310 9130 10362
rect 9130 10310 9142 10362
rect 9142 10310 9172 10362
rect 9196 10310 9206 10362
rect 9206 10310 9252 10362
rect 8956 10308 9012 10310
rect 9036 10308 9092 10310
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 8956 9274 9012 9276
rect 9036 9274 9092 9276
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 8956 9222 9002 9274
rect 9002 9222 9012 9274
rect 9036 9222 9066 9274
rect 9066 9222 9078 9274
rect 9078 9222 9092 9274
rect 9116 9222 9130 9274
rect 9130 9222 9142 9274
rect 9142 9222 9172 9274
rect 9196 9222 9206 9274
rect 9206 9222 9252 9274
rect 8956 9220 9012 9222
rect 9036 9220 9092 9222
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 9616 10906 9672 10908
rect 9696 10906 9752 10908
rect 9776 10906 9832 10908
rect 9856 10906 9912 10908
rect 9616 10854 9662 10906
rect 9662 10854 9672 10906
rect 9696 10854 9726 10906
rect 9726 10854 9738 10906
rect 9738 10854 9752 10906
rect 9776 10854 9790 10906
rect 9790 10854 9802 10906
rect 9802 10854 9832 10906
rect 9856 10854 9866 10906
rect 9866 10854 9912 10906
rect 9616 10852 9672 10854
rect 9696 10852 9752 10854
rect 9776 10852 9832 10854
rect 9856 10852 9912 10854
rect 9616 9818 9672 9820
rect 9696 9818 9752 9820
rect 9776 9818 9832 9820
rect 9856 9818 9912 9820
rect 9616 9766 9662 9818
rect 9662 9766 9672 9818
rect 9696 9766 9726 9818
rect 9726 9766 9738 9818
rect 9738 9766 9752 9818
rect 9776 9766 9790 9818
rect 9790 9766 9802 9818
rect 9802 9766 9832 9818
rect 9856 9766 9866 9818
rect 9866 9766 9912 9818
rect 9616 9764 9672 9766
rect 9696 9764 9752 9766
rect 9776 9764 9832 9766
rect 9856 9764 9912 9766
rect 9616 8730 9672 8732
rect 9696 8730 9752 8732
rect 9776 8730 9832 8732
rect 9856 8730 9912 8732
rect 9616 8678 9662 8730
rect 9662 8678 9672 8730
rect 9696 8678 9726 8730
rect 9726 8678 9738 8730
rect 9738 8678 9752 8730
rect 9776 8678 9790 8730
rect 9790 8678 9802 8730
rect 9802 8678 9832 8730
rect 9856 8678 9866 8730
rect 9866 8678 9912 8730
rect 9616 8676 9672 8678
rect 9696 8676 9752 8678
rect 9776 8676 9832 8678
rect 9856 8676 9912 8678
rect 8956 8186 9012 8188
rect 9036 8186 9092 8188
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 8956 8134 9002 8186
rect 9002 8134 9012 8186
rect 9036 8134 9066 8186
rect 9066 8134 9078 8186
rect 9078 8134 9092 8186
rect 9116 8134 9130 8186
rect 9130 8134 9142 8186
rect 9142 8134 9172 8186
rect 9196 8134 9206 8186
rect 9206 8134 9252 8186
rect 8956 8132 9012 8134
rect 9036 8132 9092 8134
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 8956 7098 9012 7100
rect 9036 7098 9092 7100
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 8956 7046 9002 7098
rect 9002 7046 9012 7098
rect 9036 7046 9066 7098
rect 9066 7046 9078 7098
rect 9078 7046 9092 7098
rect 9116 7046 9130 7098
rect 9130 7046 9142 7098
rect 9142 7046 9172 7098
rect 9196 7046 9206 7098
rect 9206 7046 9252 7098
rect 8956 7044 9012 7046
rect 9036 7044 9092 7046
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 9616 7642 9672 7644
rect 9696 7642 9752 7644
rect 9776 7642 9832 7644
rect 9856 7642 9912 7644
rect 9616 7590 9662 7642
rect 9662 7590 9672 7642
rect 9696 7590 9726 7642
rect 9726 7590 9738 7642
rect 9738 7590 9752 7642
rect 9776 7590 9790 7642
rect 9790 7590 9802 7642
rect 9802 7590 9832 7642
rect 9856 7590 9866 7642
rect 9866 7590 9912 7642
rect 9616 7588 9672 7590
rect 9696 7588 9752 7590
rect 9776 7588 9832 7590
rect 9856 7588 9912 7590
rect 8956 6010 9012 6012
rect 9036 6010 9092 6012
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 8956 5958 9002 6010
rect 9002 5958 9012 6010
rect 9036 5958 9066 6010
rect 9066 5958 9078 6010
rect 9078 5958 9092 6010
rect 9116 5958 9130 6010
rect 9130 5958 9142 6010
rect 9142 5958 9172 6010
rect 9196 5958 9206 6010
rect 9206 5958 9252 6010
rect 8956 5956 9012 5958
rect 9036 5956 9092 5958
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 8956 4922 9012 4924
rect 9036 4922 9092 4924
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 8956 4870 9002 4922
rect 9002 4870 9012 4922
rect 9036 4870 9066 4922
rect 9066 4870 9078 4922
rect 9078 4870 9092 4922
rect 9116 4870 9130 4922
rect 9130 4870 9142 4922
rect 9142 4870 9172 4922
rect 9196 4870 9206 4922
rect 9206 4870 9252 4922
rect 8956 4868 9012 4870
rect 9036 4868 9092 4870
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 8956 3834 9012 3836
rect 9036 3834 9092 3836
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 8956 3782 9002 3834
rect 9002 3782 9012 3834
rect 9036 3782 9066 3834
rect 9066 3782 9078 3834
rect 9078 3782 9092 3834
rect 9116 3782 9130 3834
rect 9130 3782 9142 3834
rect 9142 3782 9172 3834
rect 9196 3782 9206 3834
rect 9206 3782 9252 3834
rect 8956 3780 9012 3782
rect 9036 3780 9092 3782
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 9616 6554 9672 6556
rect 9696 6554 9752 6556
rect 9776 6554 9832 6556
rect 9856 6554 9912 6556
rect 9616 6502 9662 6554
rect 9662 6502 9672 6554
rect 9696 6502 9726 6554
rect 9726 6502 9738 6554
rect 9738 6502 9752 6554
rect 9776 6502 9790 6554
rect 9790 6502 9802 6554
rect 9802 6502 9832 6554
rect 9856 6502 9866 6554
rect 9866 6502 9912 6554
rect 9616 6500 9672 6502
rect 9696 6500 9752 6502
rect 9776 6500 9832 6502
rect 9856 6500 9912 6502
rect 9616 5466 9672 5468
rect 9696 5466 9752 5468
rect 9776 5466 9832 5468
rect 9856 5466 9912 5468
rect 9616 5414 9662 5466
rect 9662 5414 9672 5466
rect 9696 5414 9726 5466
rect 9726 5414 9738 5466
rect 9738 5414 9752 5466
rect 9776 5414 9790 5466
rect 9790 5414 9802 5466
rect 9802 5414 9832 5466
rect 9856 5414 9866 5466
rect 9866 5414 9912 5466
rect 9616 5412 9672 5414
rect 9696 5412 9752 5414
rect 9776 5412 9832 5414
rect 9856 5412 9912 5414
rect 9616 4378 9672 4380
rect 9696 4378 9752 4380
rect 9776 4378 9832 4380
rect 9856 4378 9912 4380
rect 9616 4326 9662 4378
rect 9662 4326 9672 4378
rect 9696 4326 9726 4378
rect 9726 4326 9738 4378
rect 9738 4326 9752 4378
rect 9776 4326 9790 4378
rect 9790 4326 9802 4378
rect 9802 4326 9832 4378
rect 9856 4326 9866 4378
rect 9866 4326 9912 4378
rect 9616 4324 9672 4326
rect 9696 4324 9752 4326
rect 9776 4324 9832 4326
rect 9856 4324 9912 4326
rect 9616 3290 9672 3292
rect 9696 3290 9752 3292
rect 9776 3290 9832 3292
rect 9856 3290 9912 3292
rect 9616 3238 9662 3290
rect 9662 3238 9672 3290
rect 9696 3238 9726 3290
rect 9726 3238 9738 3290
rect 9738 3238 9752 3290
rect 9776 3238 9790 3290
rect 9790 3238 9802 3290
rect 9802 3238 9832 3290
rect 9856 3238 9866 3290
rect 9866 3238 9912 3290
rect 9616 3236 9672 3238
rect 9696 3236 9752 3238
rect 9776 3236 9832 3238
rect 9856 3236 9912 3238
rect 13616 13082 13672 13084
rect 13696 13082 13752 13084
rect 13776 13082 13832 13084
rect 13856 13082 13912 13084
rect 13616 13030 13662 13082
rect 13662 13030 13672 13082
rect 13696 13030 13726 13082
rect 13726 13030 13738 13082
rect 13738 13030 13752 13082
rect 13776 13030 13790 13082
rect 13790 13030 13802 13082
rect 13802 13030 13832 13082
rect 13856 13030 13866 13082
rect 13866 13030 13912 13082
rect 13616 13028 13672 13030
rect 13696 13028 13752 13030
rect 13776 13028 13832 13030
rect 13856 13028 13912 13030
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13616 11994 13672 11996
rect 13696 11994 13752 11996
rect 13776 11994 13832 11996
rect 13856 11994 13912 11996
rect 13616 11942 13662 11994
rect 13662 11942 13672 11994
rect 13696 11942 13726 11994
rect 13726 11942 13738 11994
rect 13738 11942 13752 11994
rect 13776 11942 13790 11994
rect 13790 11942 13802 11994
rect 13802 11942 13832 11994
rect 13856 11942 13866 11994
rect 13866 11942 13912 11994
rect 13616 11940 13672 11942
rect 13696 11940 13752 11942
rect 13776 11940 13832 11942
rect 13856 11940 13912 11942
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 13616 10906 13672 10908
rect 13696 10906 13752 10908
rect 13776 10906 13832 10908
rect 13856 10906 13912 10908
rect 13616 10854 13662 10906
rect 13662 10854 13672 10906
rect 13696 10854 13726 10906
rect 13726 10854 13738 10906
rect 13738 10854 13752 10906
rect 13776 10854 13790 10906
rect 13790 10854 13802 10906
rect 13802 10854 13832 10906
rect 13856 10854 13866 10906
rect 13866 10854 13912 10906
rect 13616 10852 13672 10854
rect 13696 10852 13752 10854
rect 13776 10852 13832 10854
rect 13856 10852 13912 10854
rect 16946 14340 17002 14376
rect 16946 14320 16948 14340
rect 16948 14320 17000 14340
rect 17000 14320 17002 14340
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 13616 9818 13672 9820
rect 13696 9818 13752 9820
rect 13776 9818 13832 9820
rect 13856 9818 13912 9820
rect 13616 9766 13662 9818
rect 13662 9766 13672 9818
rect 13696 9766 13726 9818
rect 13726 9766 13738 9818
rect 13738 9766 13752 9818
rect 13776 9766 13790 9818
rect 13790 9766 13802 9818
rect 13802 9766 13832 9818
rect 13856 9766 13866 9818
rect 13866 9766 13912 9818
rect 13616 9764 13672 9766
rect 13696 9764 13752 9766
rect 13776 9764 13832 9766
rect 13856 9764 13912 9766
rect 13616 8730 13672 8732
rect 13696 8730 13752 8732
rect 13776 8730 13832 8732
rect 13856 8730 13912 8732
rect 13616 8678 13662 8730
rect 13662 8678 13672 8730
rect 13696 8678 13726 8730
rect 13726 8678 13738 8730
rect 13738 8678 13752 8730
rect 13776 8678 13790 8730
rect 13790 8678 13802 8730
rect 13802 8678 13832 8730
rect 13856 8678 13866 8730
rect 13866 8678 13912 8730
rect 13616 8676 13672 8678
rect 13696 8676 13752 8678
rect 13776 8676 13832 8678
rect 13856 8676 13912 8678
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 13616 7642 13672 7644
rect 13696 7642 13752 7644
rect 13776 7642 13832 7644
rect 13856 7642 13912 7644
rect 13616 7590 13662 7642
rect 13662 7590 13672 7642
rect 13696 7590 13726 7642
rect 13726 7590 13738 7642
rect 13738 7590 13752 7642
rect 13776 7590 13790 7642
rect 13790 7590 13802 7642
rect 13802 7590 13832 7642
rect 13856 7590 13866 7642
rect 13866 7590 13912 7642
rect 13616 7588 13672 7590
rect 13696 7588 13752 7590
rect 13776 7588 13832 7590
rect 13856 7588 13912 7590
rect 13616 6554 13672 6556
rect 13696 6554 13752 6556
rect 13776 6554 13832 6556
rect 13856 6554 13912 6556
rect 13616 6502 13662 6554
rect 13662 6502 13672 6554
rect 13696 6502 13726 6554
rect 13726 6502 13738 6554
rect 13738 6502 13752 6554
rect 13776 6502 13790 6554
rect 13790 6502 13802 6554
rect 13802 6502 13832 6554
rect 13856 6502 13866 6554
rect 13866 6502 13912 6554
rect 13616 6500 13672 6502
rect 13696 6500 13752 6502
rect 13776 6500 13832 6502
rect 13856 6500 13912 6502
rect 13616 5466 13672 5468
rect 13696 5466 13752 5468
rect 13776 5466 13832 5468
rect 13856 5466 13912 5468
rect 13616 5414 13662 5466
rect 13662 5414 13672 5466
rect 13696 5414 13726 5466
rect 13726 5414 13738 5466
rect 13738 5414 13752 5466
rect 13776 5414 13790 5466
rect 13790 5414 13802 5466
rect 13802 5414 13832 5466
rect 13856 5414 13866 5466
rect 13866 5414 13912 5466
rect 13616 5412 13672 5414
rect 13696 5412 13752 5414
rect 13776 5412 13832 5414
rect 13856 5412 13912 5414
rect 8956 2746 9012 2748
rect 9036 2746 9092 2748
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 8956 2694 9002 2746
rect 9002 2694 9012 2746
rect 9036 2694 9066 2746
rect 9066 2694 9078 2746
rect 9078 2694 9092 2746
rect 9116 2694 9130 2746
rect 9130 2694 9142 2746
rect 9142 2694 9172 2746
rect 9196 2694 9206 2746
rect 9206 2694 9252 2746
rect 8956 2692 9012 2694
rect 9036 2692 9092 2694
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 13616 4378 13672 4380
rect 13696 4378 13752 4380
rect 13776 4378 13832 4380
rect 13856 4378 13912 4380
rect 13616 4326 13662 4378
rect 13662 4326 13672 4378
rect 13696 4326 13726 4378
rect 13726 4326 13738 4378
rect 13738 4326 13752 4378
rect 13776 4326 13790 4378
rect 13790 4326 13802 4378
rect 13802 4326 13832 4378
rect 13856 4326 13866 4378
rect 13866 4326 13912 4378
rect 13616 4324 13672 4326
rect 13696 4324 13752 4326
rect 13776 4324 13832 4326
rect 13856 4324 13912 4326
rect 13616 3290 13672 3292
rect 13696 3290 13752 3292
rect 13776 3290 13832 3292
rect 13856 3290 13912 3292
rect 13616 3238 13662 3290
rect 13662 3238 13672 3290
rect 13696 3238 13726 3290
rect 13726 3238 13738 3290
rect 13738 3238 13752 3290
rect 13776 3238 13790 3290
rect 13790 3238 13802 3290
rect 13802 3238 13832 3290
rect 13856 3238 13866 3290
rect 13866 3238 13912 3290
rect 13616 3236 13672 3238
rect 13696 3236 13752 3238
rect 13776 3236 13832 3238
rect 13856 3236 13912 3238
rect 16946 12960 17002 13016
rect 16486 10920 16542 10976
rect 16762 8900 16818 8936
rect 16762 8880 16764 8900
rect 16764 8880 16816 8900
rect 16816 8880 16818 8900
rect 16762 7520 16818 7576
rect 16486 5516 16488 5536
rect 16488 5516 16540 5536
rect 16540 5516 16542 5536
rect 16486 5480 16542 5516
rect 16762 4120 16818 4176
rect 15658 3440 15714 3496
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 1616 2202 1672 2204
rect 1696 2202 1752 2204
rect 1776 2202 1832 2204
rect 1856 2202 1912 2204
rect 1616 2150 1662 2202
rect 1662 2150 1672 2202
rect 1696 2150 1726 2202
rect 1726 2150 1738 2202
rect 1738 2150 1752 2202
rect 1776 2150 1790 2202
rect 1790 2150 1802 2202
rect 1802 2150 1832 2202
rect 1856 2150 1866 2202
rect 1866 2150 1912 2202
rect 1616 2148 1672 2150
rect 1696 2148 1752 2150
rect 1776 2148 1832 2150
rect 1856 2148 1912 2150
rect 5616 2202 5672 2204
rect 5696 2202 5752 2204
rect 5776 2202 5832 2204
rect 5856 2202 5912 2204
rect 5616 2150 5662 2202
rect 5662 2150 5672 2202
rect 5696 2150 5726 2202
rect 5726 2150 5738 2202
rect 5738 2150 5752 2202
rect 5776 2150 5790 2202
rect 5790 2150 5802 2202
rect 5802 2150 5832 2202
rect 5856 2150 5866 2202
rect 5866 2150 5912 2202
rect 5616 2148 5672 2150
rect 5696 2148 5752 2150
rect 5776 2148 5832 2150
rect 5856 2148 5912 2150
rect 9616 2202 9672 2204
rect 9696 2202 9752 2204
rect 9776 2202 9832 2204
rect 9856 2202 9912 2204
rect 9616 2150 9662 2202
rect 9662 2150 9672 2202
rect 9696 2150 9726 2202
rect 9726 2150 9738 2202
rect 9738 2150 9752 2202
rect 9776 2150 9790 2202
rect 9790 2150 9802 2202
rect 9802 2150 9832 2202
rect 9856 2150 9866 2202
rect 9866 2150 9912 2202
rect 9616 2148 9672 2150
rect 9696 2148 9752 2150
rect 9776 2148 9832 2150
rect 9856 2148 9912 2150
rect 13616 2202 13672 2204
rect 13696 2202 13752 2204
rect 13776 2202 13832 2204
rect 13856 2202 13912 2204
rect 13616 2150 13662 2202
rect 13662 2150 13672 2202
rect 13696 2150 13726 2202
rect 13726 2150 13738 2202
rect 13738 2150 13752 2202
rect 13776 2150 13790 2202
rect 13790 2150 13802 2202
rect 13802 2150 13832 2202
rect 13856 2150 13866 2202
rect 13866 2150 13912 2202
rect 13616 2148 13672 2150
rect 13696 2148 13752 2150
rect 13776 2148 13832 2150
rect 13856 2148 13912 2150
rect 16946 2080 17002 2136
rect 16394 40 16450 96
<< metal3 >>
rect 0 17778 800 17808
rect 1485 17778 1551 17781
rect 0 17776 1551 17778
rect 0 17720 1490 17776
rect 1546 17720 1551 17776
rect 0 17718 1551 17720
rect 0 17688 800 17718
rect 1485 17715 1551 17718
rect 16481 16418 16547 16421
rect 17200 16418 18000 16448
rect 16481 16416 18000 16418
rect 16481 16360 16486 16416
rect 16542 16360 18000 16416
rect 16481 16358 18000 16360
rect 16481 16355 16547 16358
rect 17200 16328 18000 16358
rect 1393 16010 1459 16013
rect 798 16008 1459 16010
rect 798 15952 1398 16008
rect 1454 15952 1459 16008
rect 798 15950 1459 15952
rect 798 15768 858 15950
rect 1393 15947 1459 15950
rect 0 15678 858 15768
rect 946 15808 1262 15809
rect 946 15744 952 15808
rect 1016 15744 1032 15808
rect 1096 15744 1112 15808
rect 1176 15744 1192 15808
rect 1256 15744 1262 15808
rect 946 15743 1262 15744
rect 4946 15808 5262 15809
rect 4946 15744 4952 15808
rect 5016 15744 5032 15808
rect 5096 15744 5112 15808
rect 5176 15744 5192 15808
rect 5256 15744 5262 15808
rect 4946 15743 5262 15744
rect 8946 15808 9262 15809
rect 8946 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9262 15808
rect 8946 15743 9262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 0 15648 800 15678
rect 1606 15264 1922 15265
rect 1606 15200 1612 15264
rect 1676 15200 1692 15264
rect 1756 15200 1772 15264
rect 1836 15200 1852 15264
rect 1916 15200 1922 15264
rect 1606 15199 1922 15200
rect 5606 15264 5922 15265
rect 5606 15200 5612 15264
rect 5676 15200 5692 15264
rect 5756 15200 5772 15264
rect 5836 15200 5852 15264
rect 5916 15200 5922 15264
rect 5606 15199 5922 15200
rect 9606 15264 9922 15265
rect 9606 15200 9612 15264
rect 9676 15200 9692 15264
rect 9756 15200 9772 15264
rect 9836 15200 9852 15264
rect 9916 15200 9922 15264
rect 9606 15199 9922 15200
rect 13606 15264 13922 15265
rect 13606 15200 13612 15264
rect 13676 15200 13692 15264
rect 13756 15200 13772 15264
rect 13836 15200 13852 15264
rect 13916 15200 13922 15264
rect 13606 15199 13922 15200
rect 946 14720 1262 14721
rect 946 14656 952 14720
rect 1016 14656 1032 14720
rect 1096 14656 1112 14720
rect 1176 14656 1192 14720
rect 1256 14656 1262 14720
rect 946 14655 1262 14656
rect 4946 14720 5262 14721
rect 4946 14656 4952 14720
rect 5016 14656 5032 14720
rect 5096 14656 5112 14720
rect 5176 14656 5192 14720
rect 5256 14656 5262 14720
rect 4946 14655 5262 14656
rect 8946 14720 9262 14721
rect 8946 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9262 14720
rect 8946 14655 9262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 16941 14378 17007 14381
rect 17200 14378 18000 14408
rect 16941 14376 18000 14378
rect 16941 14320 16946 14376
rect 17002 14320 18000 14376
rect 16941 14318 18000 14320
rect 16941 14315 17007 14318
rect 17200 14288 18000 14318
rect 1606 14176 1922 14177
rect 1606 14112 1612 14176
rect 1676 14112 1692 14176
rect 1756 14112 1772 14176
rect 1836 14112 1852 14176
rect 1916 14112 1922 14176
rect 1606 14111 1922 14112
rect 5606 14176 5922 14177
rect 5606 14112 5612 14176
rect 5676 14112 5692 14176
rect 5756 14112 5772 14176
rect 5836 14112 5852 14176
rect 5916 14112 5922 14176
rect 5606 14111 5922 14112
rect 9606 14176 9922 14177
rect 9606 14112 9612 14176
rect 9676 14112 9692 14176
rect 9756 14112 9772 14176
rect 9836 14112 9852 14176
rect 9916 14112 9922 14176
rect 9606 14111 9922 14112
rect 13606 14176 13922 14177
rect 13606 14112 13612 14176
rect 13676 14112 13692 14176
rect 13756 14112 13772 14176
rect 13836 14112 13852 14176
rect 13916 14112 13922 14176
rect 13606 14111 13922 14112
rect 798 13774 1410 13834
rect 798 13728 858 13774
rect 0 13638 858 13728
rect 1350 13701 1410 13774
rect 1350 13696 1459 13701
rect 1350 13640 1398 13696
rect 1454 13640 1459 13696
rect 1350 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 946 13632 1262 13633
rect 946 13568 952 13632
rect 1016 13568 1032 13632
rect 1096 13568 1112 13632
rect 1176 13568 1192 13632
rect 1256 13568 1262 13632
rect 946 13567 1262 13568
rect 4946 13632 5262 13633
rect 4946 13568 4952 13632
rect 5016 13568 5032 13632
rect 5096 13568 5112 13632
rect 5176 13568 5192 13632
rect 5256 13568 5262 13632
rect 4946 13567 5262 13568
rect 8946 13632 9262 13633
rect 8946 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9262 13632
rect 8946 13567 9262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 1606 13088 1922 13089
rect 1606 13024 1612 13088
rect 1676 13024 1692 13088
rect 1756 13024 1772 13088
rect 1836 13024 1852 13088
rect 1916 13024 1922 13088
rect 1606 13023 1922 13024
rect 5606 13088 5922 13089
rect 5606 13024 5612 13088
rect 5676 13024 5692 13088
rect 5756 13024 5772 13088
rect 5836 13024 5852 13088
rect 5916 13024 5922 13088
rect 5606 13023 5922 13024
rect 9606 13088 9922 13089
rect 9606 13024 9612 13088
rect 9676 13024 9692 13088
rect 9756 13024 9772 13088
rect 9836 13024 9852 13088
rect 9916 13024 9922 13088
rect 9606 13023 9922 13024
rect 13606 13088 13922 13089
rect 13606 13024 13612 13088
rect 13676 13024 13692 13088
rect 13756 13024 13772 13088
rect 13836 13024 13852 13088
rect 13916 13024 13922 13088
rect 13606 13023 13922 13024
rect 16941 13018 17007 13021
rect 17200 13018 18000 13048
rect 16941 13016 18000 13018
rect 16941 12960 16946 13016
rect 17002 12960 18000 13016
rect 16941 12958 18000 12960
rect 16941 12955 17007 12958
rect 17200 12928 18000 12958
rect 946 12544 1262 12545
rect 946 12480 952 12544
rect 1016 12480 1032 12544
rect 1096 12480 1112 12544
rect 1176 12480 1192 12544
rect 1256 12480 1262 12544
rect 946 12479 1262 12480
rect 4946 12544 5262 12545
rect 4946 12480 4952 12544
rect 5016 12480 5032 12544
rect 5096 12480 5112 12544
rect 5176 12480 5192 12544
rect 5256 12480 5262 12544
rect 4946 12479 5262 12480
rect 8946 12544 9262 12545
rect 8946 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9262 12544
rect 8946 12479 9262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 1606 12000 1922 12001
rect 1606 11936 1612 12000
rect 1676 11936 1692 12000
rect 1756 11936 1772 12000
rect 1836 11936 1852 12000
rect 1916 11936 1922 12000
rect 1606 11935 1922 11936
rect 5606 12000 5922 12001
rect 5606 11936 5612 12000
rect 5676 11936 5692 12000
rect 5756 11936 5772 12000
rect 5836 11936 5852 12000
rect 5916 11936 5922 12000
rect 5606 11935 5922 11936
rect 9606 12000 9922 12001
rect 9606 11936 9612 12000
rect 9676 11936 9692 12000
rect 9756 11936 9772 12000
rect 9836 11936 9852 12000
rect 9916 11936 9922 12000
rect 9606 11935 9922 11936
rect 13606 12000 13922 12001
rect 13606 11936 13612 12000
rect 13676 11936 13692 12000
rect 13756 11936 13772 12000
rect 13836 11936 13852 12000
rect 13916 11936 13922 12000
rect 13606 11935 13922 11936
rect 946 11456 1262 11457
rect 946 11392 952 11456
rect 1016 11392 1032 11456
rect 1096 11392 1112 11456
rect 1176 11392 1192 11456
rect 1256 11392 1262 11456
rect 946 11391 1262 11392
rect 4946 11456 5262 11457
rect 4946 11392 4952 11456
rect 5016 11392 5032 11456
rect 5096 11392 5112 11456
rect 5176 11392 5192 11456
rect 5256 11392 5262 11456
rect 4946 11391 5262 11392
rect 8946 11456 9262 11457
rect 8946 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9262 11456
rect 8946 11391 9262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 16481 10978 16547 10981
rect 17200 10978 18000 11008
rect 16481 10976 18000 10978
rect 16481 10920 16486 10976
rect 16542 10920 18000 10976
rect 16481 10918 18000 10920
rect 16481 10915 16547 10918
rect 1606 10912 1922 10913
rect 1606 10848 1612 10912
rect 1676 10848 1692 10912
rect 1756 10848 1772 10912
rect 1836 10848 1852 10912
rect 1916 10848 1922 10912
rect 1606 10847 1922 10848
rect 5606 10912 5922 10913
rect 5606 10848 5612 10912
rect 5676 10848 5692 10912
rect 5756 10848 5772 10912
rect 5836 10848 5852 10912
rect 5916 10848 5922 10912
rect 5606 10847 5922 10848
rect 9606 10912 9922 10913
rect 9606 10848 9612 10912
rect 9676 10848 9692 10912
rect 9756 10848 9772 10912
rect 9836 10848 9852 10912
rect 9916 10848 9922 10912
rect 9606 10847 9922 10848
rect 13606 10912 13922 10913
rect 13606 10848 13612 10912
rect 13676 10848 13692 10912
rect 13756 10848 13772 10912
rect 13836 10848 13852 10912
rect 13916 10848 13922 10912
rect 17200 10888 18000 10918
rect 13606 10847 13922 10848
rect 946 10368 1262 10369
rect 0 10298 800 10328
rect 946 10304 952 10368
rect 1016 10304 1032 10368
rect 1096 10304 1112 10368
rect 1176 10304 1192 10368
rect 1256 10304 1262 10368
rect 946 10303 1262 10304
rect 4946 10368 5262 10369
rect 4946 10304 4952 10368
rect 5016 10304 5032 10368
rect 5096 10304 5112 10368
rect 5176 10304 5192 10368
rect 5256 10304 5262 10368
rect 4946 10303 5262 10304
rect 8946 10368 9262 10369
rect 8946 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9262 10368
rect 8946 10303 9262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 0 10208 858 10298
rect 798 10162 858 10208
rect 933 10162 999 10165
rect 798 10160 999 10162
rect 798 10104 938 10160
rect 994 10104 999 10160
rect 798 10102 999 10104
rect 933 10099 999 10102
rect 1606 9824 1922 9825
rect 1606 9760 1612 9824
rect 1676 9760 1692 9824
rect 1756 9760 1772 9824
rect 1836 9760 1852 9824
rect 1916 9760 1922 9824
rect 1606 9759 1922 9760
rect 5606 9824 5922 9825
rect 5606 9760 5612 9824
rect 5676 9760 5692 9824
rect 5756 9760 5772 9824
rect 5836 9760 5852 9824
rect 5916 9760 5922 9824
rect 5606 9759 5922 9760
rect 9606 9824 9922 9825
rect 9606 9760 9612 9824
rect 9676 9760 9692 9824
rect 9756 9760 9772 9824
rect 9836 9760 9852 9824
rect 9916 9760 9922 9824
rect 9606 9759 9922 9760
rect 13606 9824 13922 9825
rect 13606 9760 13612 9824
rect 13676 9760 13692 9824
rect 13756 9760 13772 9824
rect 13836 9760 13852 9824
rect 13916 9760 13922 9824
rect 13606 9759 13922 9760
rect 946 9280 1262 9281
rect 946 9216 952 9280
rect 1016 9216 1032 9280
rect 1096 9216 1112 9280
rect 1176 9216 1192 9280
rect 1256 9216 1262 9280
rect 946 9215 1262 9216
rect 4946 9280 5262 9281
rect 4946 9216 4952 9280
rect 5016 9216 5032 9280
rect 5096 9216 5112 9280
rect 5176 9216 5192 9280
rect 5256 9216 5262 9280
rect 4946 9215 5262 9216
rect 8946 9280 9262 9281
rect 8946 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9262 9280
rect 8946 9215 9262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 16757 8938 16823 8941
rect 17200 8938 18000 8968
rect 16757 8936 18000 8938
rect 16757 8880 16762 8936
rect 16818 8880 18000 8936
rect 16757 8878 18000 8880
rect 16757 8875 16823 8878
rect 17200 8848 18000 8878
rect 1606 8736 1922 8737
rect 1606 8672 1612 8736
rect 1676 8672 1692 8736
rect 1756 8672 1772 8736
rect 1836 8672 1852 8736
rect 1916 8672 1922 8736
rect 1606 8671 1922 8672
rect 5606 8736 5922 8737
rect 5606 8672 5612 8736
rect 5676 8672 5692 8736
rect 5756 8672 5772 8736
rect 5836 8672 5852 8736
rect 5916 8672 5922 8736
rect 5606 8671 5922 8672
rect 9606 8736 9922 8737
rect 9606 8672 9612 8736
rect 9676 8672 9692 8736
rect 9756 8672 9772 8736
rect 9836 8672 9852 8736
rect 9916 8672 9922 8736
rect 9606 8671 9922 8672
rect 13606 8736 13922 8737
rect 13606 8672 13612 8736
rect 13676 8672 13692 8736
rect 13756 8672 13772 8736
rect 13836 8672 13852 8736
rect 13916 8672 13922 8736
rect 13606 8671 13922 8672
rect 946 8192 1262 8193
rect 946 8128 952 8192
rect 1016 8128 1032 8192
rect 1096 8128 1112 8192
rect 1176 8128 1192 8192
rect 1256 8128 1262 8192
rect 946 8127 1262 8128
rect 4946 8192 5262 8193
rect 4946 8128 4952 8192
rect 5016 8128 5032 8192
rect 5096 8128 5112 8192
rect 5176 8128 5192 8192
rect 5256 8128 5262 8192
rect 4946 8127 5262 8128
rect 8946 8192 9262 8193
rect 8946 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9262 8192
rect 8946 8127 9262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 1606 7648 1922 7649
rect 1606 7584 1612 7648
rect 1676 7584 1692 7648
rect 1756 7584 1772 7648
rect 1836 7584 1852 7648
rect 1916 7584 1922 7648
rect 1606 7583 1922 7584
rect 5606 7648 5922 7649
rect 5606 7584 5612 7648
rect 5676 7584 5692 7648
rect 5756 7584 5772 7648
rect 5836 7584 5852 7648
rect 5916 7584 5922 7648
rect 5606 7583 5922 7584
rect 9606 7648 9922 7649
rect 9606 7584 9612 7648
rect 9676 7584 9692 7648
rect 9756 7584 9772 7648
rect 9836 7584 9852 7648
rect 9916 7584 9922 7648
rect 9606 7583 9922 7584
rect 13606 7648 13922 7649
rect 13606 7584 13612 7648
rect 13676 7584 13692 7648
rect 13756 7584 13772 7648
rect 13836 7584 13852 7648
rect 13916 7584 13922 7648
rect 13606 7583 13922 7584
rect 16757 7578 16823 7581
rect 17200 7578 18000 7608
rect 16757 7576 18000 7578
rect 16757 7520 16762 7576
rect 16818 7520 18000 7576
rect 16757 7518 18000 7520
rect 16757 7515 16823 7518
rect 17200 7488 18000 7518
rect 4521 7442 4587 7445
rect 7557 7442 7623 7445
rect 4521 7440 7623 7442
rect 4521 7384 4526 7440
rect 4582 7384 7562 7440
rect 7618 7384 7623 7440
rect 4521 7382 7623 7384
rect 4521 7379 4587 7382
rect 7557 7379 7623 7382
rect 3417 7306 3483 7309
rect 5349 7306 5415 7309
rect 3417 7304 5415 7306
rect 3417 7248 3422 7304
rect 3478 7248 5354 7304
rect 5410 7248 5415 7304
rect 3417 7246 5415 7248
rect 3417 7243 3483 7246
rect 5349 7243 5415 7246
rect 946 7104 1262 7105
rect 946 7040 952 7104
rect 1016 7040 1032 7104
rect 1096 7040 1112 7104
rect 1176 7040 1192 7104
rect 1256 7040 1262 7104
rect 946 7039 1262 7040
rect 4946 7104 5262 7105
rect 4946 7040 4952 7104
rect 5016 7040 5032 7104
rect 5096 7040 5112 7104
rect 5176 7040 5192 7104
rect 5256 7040 5262 7104
rect 4946 7039 5262 7040
rect 8946 7104 9262 7105
rect 8946 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9262 7104
rect 8946 7039 9262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 0 6898 800 6928
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6808 800 6838
rect 933 6835 999 6838
rect 1606 6560 1922 6561
rect 1606 6496 1612 6560
rect 1676 6496 1692 6560
rect 1756 6496 1772 6560
rect 1836 6496 1852 6560
rect 1916 6496 1922 6560
rect 1606 6495 1922 6496
rect 5606 6560 5922 6561
rect 5606 6496 5612 6560
rect 5676 6496 5692 6560
rect 5756 6496 5772 6560
rect 5836 6496 5852 6560
rect 5916 6496 5922 6560
rect 5606 6495 5922 6496
rect 9606 6560 9922 6561
rect 9606 6496 9612 6560
rect 9676 6496 9692 6560
rect 9756 6496 9772 6560
rect 9836 6496 9852 6560
rect 9916 6496 9922 6560
rect 9606 6495 9922 6496
rect 13606 6560 13922 6561
rect 13606 6496 13612 6560
rect 13676 6496 13692 6560
rect 13756 6496 13772 6560
rect 13836 6496 13852 6560
rect 13916 6496 13922 6560
rect 13606 6495 13922 6496
rect 946 6016 1262 6017
rect 946 5952 952 6016
rect 1016 5952 1032 6016
rect 1096 5952 1112 6016
rect 1176 5952 1192 6016
rect 1256 5952 1262 6016
rect 946 5951 1262 5952
rect 4946 6016 5262 6017
rect 4946 5952 4952 6016
rect 5016 5952 5032 6016
rect 5096 5952 5112 6016
rect 5176 5952 5192 6016
rect 5256 5952 5262 6016
rect 4946 5951 5262 5952
rect 8946 6016 9262 6017
rect 8946 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9262 6016
rect 8946 5951 9262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 16481 5538 16547 5541
rect 17200 5538 18000 5568
rect 16481 5536 18000 5538
rect 16481 5480 16486 5536
rect 16542 5480 18000 5536
rect 16481 5478 18000 5480
rect 16481 5475 16547 5478
rect 1606 5472 1922 5473
rect 1606 5408 1612 5472
rect 1676 5408 1692 5472
rect 1756 5408 1772 5472
rect 1836 5408 1852 5472
rect 1916 5408 1922 5472
rect 1606 5407 1922 5408
rect 5606 5472 5922 5473
rect 5606 5408 5612 5472
rect 5676 5408 5692 5472
rect 5756 5408 5772 5472
rect 5836 5408 5852 5472
rect 5916 5408 5922 5472
rect 5606 5407 5922 5408
rect 9606 5472 9922 5473
rect 9606 5408 9612 5472
rect 9676 5408 9692 5472
rect 9756 5408 9772 5472
rect 9836 5408 9852 5472
rect 9916 5408 9922 5472
rect 9606 5407 9922 5408
rect 13606 5472 13922 5473
rect 13606 5408 13612 5472
rect 13676 5408 13692 5472
rect 13756 5408 13772 5472
rect 13836 5408 13852 5472
rect 13916 5408 13922 5472
rect 17200 5448 18000 5478
rect 13606 5407 13922 5408
rect 749 5130 815 5133
rect 749 5128 858 5130
rect 749 5072 754 5128
rect 810 5072 858 5128
rect 749 5067 858 5072
rect 798 4888 858 5067
rect 0 4798 858 4888
rect 946 4928 1262 4929
rect 946 4864 952 4928
rect 1016 4864 1032 4928
rect 1096 4864 1112 4928
rect 1176 4864 1192 4928
rect 1256 4864 1262 4928
rect 946 4863 1262 4864
rect 4946 4928 5262 4929
rect 4946 4864 4952 4928
rect 5016 4864 5032 4928
rect 5096 4864 5112 4928
rect 5176 4864 5192 4928
rect 5256 4864 5262 4928
rect 4946 4863 5262 4864
rect 8946 4928 9262 4929
rect 8946 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9262 4928
rect 8946 4863 9262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 0 4768 800 4798
rect 1606 4384 1922 4385
rect 1606 4320 1612 4384
rect 1676 4320 1692 4384
rect 1756 4320 1772 4384
rect 1836 4320 1852 4384
rect 1916 4320 1922 4384
rect 1606 4319 1922 4320
rect 5606 4384 5922 4385
rect 5606 4320 5612 4384
rect 5676 4320 5692 4384
rect 5756 4320 5772 4384
rect 5836 4320 5852 4384
rect 5916 4320 5922 4384
rect 5606 4319 5922 4320
rect 9606 4384 9922 4385
rect 9606 4320 9612 4384
rect 9676 4320 9692 4384
rect 9756 4320 9772 4384
rect 9836 4320 9852 4384
rect 9916 4320 9922 4384
rect 9606 4319 9922 4320
rect 13606 4384 13922 4385
rect 13606 4320 13612 4384
rect 13676 4320 13692 4384
rect 13756 4320 13772 4384
rect 13836 4320 13852 4384
rect 13916 4320 13922 4384
rect 13606 4319 13922 4320
rect 16757 4178 16823 4181
rect 17200 4178 18000 4208
rect 16757 4176 18000 4178
rect 16757 4120 16762 4176
rect 16818 4120 18000 4176
rect 16757 4118 18000 4120
rect 16757 4115 16823 4118
rect 17200 4088 18000 4118
rect 946 3840 1262 3841
rect 946 3776 952 3840
rect 1016 3776 1032 3840
rect 1096 3776 1112 3840
rect 1176 3776 1192 3840
rect 1256 3776 1262 3840
rect 946 3775 1262 3776
rect 4946 3840 5262 3841
rect 4946 3776 4952 3840
rect 5016 3776 5032 3840
rect 5096 3776 5112 3840
rect 5176 3776 5192 3840
rect 5256 3776 5262 3840
rect 4946 3775 5262 3776
rect 8946 3840 9262 3841
rect 8946 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9262 3840
rect 8946 3775 9262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 4061 3498 4127 3501
rect 15653 3498 15719 3501
rect 4061 3496 15719 3498
rect 4061 3440 4066 3496
rect 4122 3440 15658 3496
rect 15714 3440 15719 3496
rect 4061 3438 15719 3440
rect 4061 3435 4127 3438
rect 15653 3435 15719 3438
rect 1606 3296 1922 3297
rect 1606 3232 1612 3296
rect 1676 3232 1692 3296
rect 1756 3232 1772 3296
rect 1836 3232 1852 3296
rect 1916 3232 1922 3296
rect 1606 3231 1922 3232
rect 5606 3296 5922 3297
rect 5606 3232 5612 3296
rect 5676 3232 5692 3296
rect 5756 3232 5772 3296
rect 5836 3232 5852 3296
rect 5916 3232 5922 3296
rect 5606 3231 5922 3232
rect 9606 3296 9922 3297
rect 9606 3232 9612 3296
rect 9676 3232 9692 3296
rect 9756 3232 9772 3296
rect 9836 3232 9852 3296
rect 9916 3232 9922 3296
rect 9606 3231 9922 3232
rect 13606 3296 13922 3297
rect 13606 3232 13612 3296
rect 13676 3232 13692 3296
rect 13756 3232 13772 3296
rect 13836 3232 13852 3296
rect 13916 3232 13922 3296
rect 13606 3231 13922 3232
rect 946 2752 1262 2753
rect 946 2688 952 2752
rect 1016 2688 1032 2752
rect 1096 2688 1112 2752
rect 1176 2688 1192 2752
rect 1256 2688 1262 2752
rect 946 2687 1262 2688
rect 4946 2752 5262 2753
rect 4946 2688 4952 2752
rect 5016 2688 5032 2752
rect 5096 2688 5112 2752
rect 5176 2688 5192 2752
rect 5256 2688 5262 2752
rect 4946 2687 5262 2688
rect 8946 2752 9262 2753
rect 8946 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9262 2752
rect 8946 2687 9262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 1606 2208 1922 2209
rect 1606 2144 1612 2208
rect 1676 2144 1692 2208
rect 1756 2144 1772 2208
rect 1836 2144 1852 2208
rect 1916 2144 1922 2208
rect 1606 2143 1922 2144
rect 5606 2208 5922 2209
rect 5606 2144 5612 2208
rect 5676 2144 5692 2208
rect 5756 2144 5772 2208
rect 5836 2144 5852 2208
rect 5916 2144 5922 2208
rect 5606 2143 5922 2144
rect 9606 2208 9922 2209
rect 9606 2144 9612 2208
rect 9676 2144 9692 2208
rect 9756 2144 9772 2208
rect 9836 2144 9852 2208
rect 9916 2144 9922 2208
rect 9606 2143 9922 2144
rect 13606 2208 13922 2209
rect 13606 2144 13612 2208
rect 13676 2144 13692 2208
rect 13756 2144 13772 2208
rect 13836 2144 13852 2208
rect 13916 2144 13922 2208
rect 13606 2143 13922 2144
rect 16941 2138 17007 2141
rect 17200 2138 18000 2168
rect 16941 2136 18000 2138
rect 16941 2080 16946 2136
rect 17002 2080 18000 2136
rect 16941 2078 18000 2080
rect 16941 2075 17007 2078
rect 17200 2048 18000 2078
rect 0 1458 800 1488
rect 933 1458 999 1461
rect 0 1456 999 1458
rect 0 1400 938 1456
rect 994 1400 999 1456
rect 0 1398 999 1400
rect 0 1368 800 1398
rect 933 1395 999 1398
rect 16389 98 16455 101
rect 17200 98 18000 128
rect 16389 96 18000 98
rect 16389 40 16394 96
rect 16450 40 18000 96
rect 16389 38 18000 40
rect 16389 35 16455 38
rect 17200 8 18000 38
<< via3 >>
rect 952 15804 1016 15808
rect 952 15748 956 15804
rect 956 15748 1012 15804
rect 1012 15748 1016 15804
rect 952 15744 1016 15748
rect 1032 15804 1096 15808
rect 1032 15748 1036 15804
rect 1036 15748 1092 15804
rect 1092 15748 1096 15804
rect 1032 15744 1096 15748
rect 1112 15804 1176 15808
rect 1112 15748 1116 15804
rect 1116 15748 1172 15804
rect 1172 15748 1176 15804
rect 1112 15744 1176 15748
rect 1192 15804 1256 15808
rect 1192 15748 1196 15804
rect 1196 15748 1252 15804
rect 1252 15748 1256 15804
rect 1192 15744 1256 15748
rect 4952 15804 5016 15808
rect 4952 15748 4956 15804
rect 4956 15748 5012 15804
rect 5012 15748 5016 15804
rect 4952 15744 5016 15748
rect 5032 15804 5096 15808
rect 5032 15748 5036 15804
rect 5036 15748 5092 15804
rect 5092 15748 5096 15804
rect 5032 15744 5096 15748
rect 5112 15804 5176 15808
rect 5112 15748 5116 15804
rect 5116 15748 5172 15804
rect 5172 15748 5176 15804
rect 5112 15744 5176 15748
rect 5192 15804 5256 15808
rect 5192 15748 5196 15804
rect 5196 15748 5252 15804
rect 5252 15748 5256 15804
rect 5192 15744 5256 15748
rect 8952 15804 9016 15808
rect 8952 15748 8956 15804
rect 8956 15748 9012 15804
rect 9012 15748 9016 15804
rect 8952 15744 9016 15748
rect 9032 15804 9096 15808
rect 9032 15748 9036 15804
rect 9036 15748 9092 15804
rect 9092 15748 9096 15804
rect 9032 15744 9096 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 1612 15260 1676 15264
rect 1612 15204 1616 15260
rect 1616 15204 1672 15260
rect 1672 15204 1676 15260
rect 1612 15200 1676 15204
rect 1692 15260 1756 15264
rect 1692 15204 1696 15260
rect 1696 15204 1752 15260
rect 1752 15204 1756 15260
rect 1692 15200 1756 15204
rect 1772 15260 1836 15264
rect 1772 15204 1776 15260
rect 1776 15204 1832 15260
rect 1832 15204 1836 15260
rect 1772 15200 1836 15204
rect 1852 15260 1916 15264
rect 1852 15204 1856 15260
rect 1856 15204 1912 15260
rect 1912 15204 1916 15260
rect 1852 15200 1916 15204
rect 5612 15260 5676 15264
rect 5612 15204 5616 15260
rect 5616 15204 5672 15260
rect 5672 15204 5676 15260
rect 5612 15200 5676 15204
rect 5692 15260 5756 15264
rect 5692 15204 5696 15260
rect 5696 15204 5752 15260
rect 5752 15204 5756 15260
rect 5692 15200 5756 15204
rect 5772 15260 5836 15264
rect 5772 15204 5776 15260
rect 5776 15204 5832 15260
rect 5832 15204 5836 15260
rect 5772 15200 5836 15204
rect 5852 15260 5916 15264
rect 5852 15204 5856 15260
rect 5856 15204 5912 15260
rect 5912 15204 5916 15260
rect 5852 15200 5916 15204
rect 9612 15260 9676 15264
rect 9612 15204 9616 15260
rect 9616 15204 9672 15260
rect 9672 15204 9676 15260
rect 9612 15200 9676 15204
rect 9692 15260 9756 15264
rect 9692 15204 9696 15260
rect 9696 15204 9752 15260
rect 9752 15204 9756 15260
rect 9692 15200 9756 15204
rect 9772 15260 9836 15264
rect 9772 15204 9776 15260
rect 9776 15204 9832 15260
rect 9832 15204 9836 15260
rect 9772 15200 9836 15204
rect 9852 15260 9916 15264
rect 9852 15204 9856 15260
rect 9856 15204 9912 15260
rect 9912 15204 9916 15260
rect 9852 15200 9916 15204
rect 13612 15260 13676 15264
rect 13612 15204 13616 15260
rect 13616 15204 13672 15260
rect 13672 15204 13676 15260
rect 13612 15200 13676 15204
rect 13692 15260 13756 15264
rect 13692 15204 13696 15260
rect 13696 15204 13752 15260
rect 13752 15204 13756 15260
rect 13692 15200 13756 15204
rect 13772 15260 13836 15264
rect 13772 15204 13776 15260
rect 13776 15204 13832 15260
rect 13832 15204 13836 15260
rect 13772 15200 13836 15204
rect 13852 15260 13916 15264
rect 13852 15204 13856 15260
rect 13856 15204 13912 15260
rect 13912 15204 13916 15260
rect 13852 15200 13916 15204
rect 952 14716 1016 14720
rect 952 14660 956 14716
rect 956 14660 1012 14716
rect 1012 14660 1016 14716
rect 952 14656 1016 14660
rect 1032 14716 1096 14720
rect 1032 14660 1036 14716
rect 1036 14660 1092 14716
rect 1092 14660 1096 14716
rect 1032 14656 1096 14660
rect 1112 14716 1176 14720
rect 1112 14660 1116 14716
rect 1116 14660 1172 14716
rect 1172 14660 1176 14716
rect 1112 14656 1176 14660
rect 1192 14716 1256 14720
rect 1192 14660 1196 14716
rect 1196 14660 1252 14716
rect 1252 14660 1256 14716
rect 1192 14656 1256 14660
rect 4952 14716 5016 14720
rect 4952 14660 4956 14716
rect 4956 14660 5012 14716
rect 5012 14660 5016 14716
rect 4952 14656 5016 14660
rect 5032 14716 5096 14720
rect 5032 14660 5036 14716
rect 5036 14660 5092 14716
rect 5092 14660 5096 14716
rect 5032 14656 5096 14660
rect 5112 14716 5176 14720
rect 5112 14660 5116 14716
rect 5116 14660 5172 14716
rect 5172 14660 5176 14716
rect 5112 14656 5176 14660
rect 5192 14716 5256 14720
rect 5192 14660 5196 14716
rect 5196 14660 5252 14716
rect 5252 14660 5256 14716
rect 5192 14656 5256 14660
rect 8952 14716 9016 14720
rect 8952 14660 8956 14716
rect 8956 14660 9012 14716
rect 9012 14660 9016 14716
rect 8952 14656 9016 14660
rect 9032 14716 9096 14720
rect 9032 14660 9036 14716
rect 9036 14660 9092 14716
rect 9092 14660 9096 14716
rect 9032 14656 9096 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 1612 14172 1676 14176
rect 1612 14116 1616 14172
rect 1616 14116 1672 14172
rect 1672 14116 1676 14172
rect 1612 14112 1676 14116
rect 1692 14172 1756 14176
rect 1692 14116 1696 14172
rect 1696 14116 1752 14172
rect 1752 14116 1756 14172
rect 1692 14112 1756 14116
rect 1772 14172 1836 14176
rect 1772 14116 1776 14172
rect 1776 14116 1832 14172
rect 1832 14116 1836 14172
rect 1772 14112 1836 14116
rect 1852 14172 1916 14176
rect 1852 14116 1856 14172
rect 1856 14116 1912 14172
rect 1912 14116 1916 14172
rect 1852 14112 1916 14116
rect 5612 14172 5676 14176
rect 5612 14116 5616 14172
rect 5616 14116 5672 14172
rect 5672 14116 5676 14172
rect 5612 14112 5676 14116
rect 5692 14172 5756 14176
rect 5692 14116 5696 14172
rect 5696 14116 5752 14172
rect 5752 14116 5756 14172
rect 5692 14112 5756 14116
rect 5772 14172 5836 14176
rect 5772 14116 5776 14172
rect 5776 14116 5832 14172
rect 5832 14116 5836 14172
rect 5772 14112 5836 14116
rect 5852 14172 5916 14176
rect 5852 14116 5856 14172
rect 5856 14116 5912 14172
rect 5912 14116 5916 14172
rect 5852 14112 5916 14116
rect 9612 14172 9676 14176
rect 9612 14116 9616 14172
rect 9616 14116 9672 14172
rect 9672 14116 9676 14172
rect 9612 14112 9676 14116
rect 9692 14172 9756 14176
rect 9692 14116 9696 14172
rect 9696 14116 9752 14172
rect 9752 14116 9756 14172
rect 9692 14112 9756 14116
rect 9772 14172 9836 14176
rect 9772 14116 9776 14172
rect 9776 14116 9832 14172
rect 9832 14116 9836 14172
rect 9772 14112 9836 14116
rect 9852 14172 9916 14176
rect 9852 14116 9856 14172
rect 9856 14116 9912 14172
rect 9912 14116 9916 14172
rect 9852 14112 9916 14116
rect 13612 14172 13676 14176
rect 13612 14116 13616 14172
rect 13616 14116 13672 14172
rect 13672 14116 13676 14172
rect 13612 14112 13676 14116
rect 13692 14172 13756 14176
rect 13692 14116 13696 14172
rect 13696 14116 13752 14172
rect 13752 14116 13756 14172
rect 13692 14112 13756 14116
rect 13772 14172 13836 14176
rect 13772 14116 13776 14172
rect 13776 14116 13832 14172
rect 13832 14116 13836 14172
rect 13772 14112 13836 14116
rect 13852 14172 13916 14176
rect 13852 14116 13856 14172
rect 13856 14116 13912 14172
rect 13912 14116 13916 14172
rect 13852 14112 13916 14116
rect 952 13628 1016 13632
rect 952 13572 956 13628
rect 956 13572 1012 13628
rect 1012 13572 1016 13628
rect 952 13568 1016 13572
rect 1032 13628 1096 13632
rect 1032 13572 1036 13628
rect 1036 13572 1092 13628
rect 1092 13572 1096 13628
rect 1032 13568 1096 13572
rect 1112 13628 1176 13632
rect 1112 13572 1116 13628
rect 1116 13572 1172 13628
rect 1172 13572 1176 13628
rect 1112 13568 1176 13572
rect 1192 13628 1256 13632
rect 1192 13572 1196 13628
rect 1196 13572 1252 13628
rect 1252 13572 1256 13628
rect 1192 13568 1256 13572
rect 4952 13628 5016 13632
rect 4952 13572 4956 13628
rect 4956 13572 5012 13628
rect 5012 13572 5016 13628
rect 4952 13568 5016 13572
rect 5032 13628 5096 13632
rect 5032 13572 5036 13628
rect 5036 13572 5092 13628
rect 5092 13572 5096 13628
rect 5032 13568 5096 13572
rect 5112 13628 5176 13632
rect 5112 13572 5116 13628
rect 5116 13572 5172 13628
rect 5172 13572 5176 13628
rect 5112 13568 5176 13572
rect 5192 13628 5256 13632
rect 5192 13572 5196 13628
rect 5196 13572 5252 13628
rect 5252 13572 5256 13628
rect 5192 13568 5256 13572
rect 8952 13628 9016 13632
rect 8952 13572 8956 13628
rect 8956 13572 9012 13628
rect 9012 13572 9016 13628
rect 8952 13568 9016 13572
rect 9032 13628 9096 13632
rect 9032 13572 9036 13628
rect 9036 13572 9092 13628
rect 9092 13572 9096 13628
rect 9032 13568 9096 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 1612 13084 1676 13088
rect 1612 13028 1616 13084
rect 1616 13028 1672 13084
rect 1672 13028 1676 13084
rect 1612 13024 1676 13028
rect 1692 13084 1756 13088
rect 1692 13028 1696 13084
rect 1696 13028 1752 13084
rect 1752 13028 1756 13084
rect 1692 13024 1756 13028
rect 1772 13084 1836 13088
rect 1772 13028 1776 13084
rect 1776 13028 1832 13084
rect 1832 13028 1836 13084
rect 1772 13024 1836 13028
rect 1852 13084 1916 13088
rect 1852 13028 1856 13084
rect 1856 13028 1912 13084
rect 1912 13028 1916 13084
rect 1852 13024 1916 13028
rect 5612 13084 5676 13088
rect 5612 13028 5616 13084
rect 5616 13028 5672 13084
rect 5672 13028 5676 13084
rect 5612 13024 5676 13028
rect 5692 13084 5756 13088
rect 5692 13028 5696 13084
rect 5696 13028 5752 13084
rect 5752 13028 5756 13084
rect 5692 13024 5756 13028
rect 5772 13084 5836 13088
rect 5772 13028 5776 13084
rect 5776 13028 5832 13084
rect 5832 13028 5836 13084
rect 5772 13024 5836 13028
rect 5852 13084 5916 13088
rect 5852 13028 5856 13084
rect 5856 13028 5912 13084
rect 5912 13028 5916 13084
rect 5852 13024 5916 13028
rect 9612 13084 9676 13088
rect 9612 13028 9616 13084
rect 9616 13028 9672 13084
rect 9672 13028 9676 13084
rect 9612 13024 9676 13028
rect 9692 13084 9756 13088
rect 9692 13028 9696 13084
rect 9696 13028 9752 13084
rect 9752 13028 9756 13084
rect 9692 13024 9756 13028
rect 9772 13084 9836 13088
rect 9772 13028 9776 13084
rect 9776 13028 9832 13084
rect 9832 13028 9836 13084
rect 9772 13024 9836 13028
rect 9852 13084 9916 13088
rect 9852 13028 9856 13084
rect 9856 13028 9912 13084
rect 9912 13028 9916 13084
rect 9852 13024 9916 13028
rect 13612 13084 13676 13088
rect 13612 13028 13616 13084
rect 13616 13028 13672 13084
rect 13672 13028 13676 13084
rect 13612 13024 13676 13028
rect 13692 13084 13756 13088
rect 13692 13028 13696 13084
rect 13696 13028 13752 13084
rect 13752 13028 13756 13084
rect 13692 13024 13756 13028
rect 13772 13084 13836 13088
rect 13772 13028 13776 13084
rect 13776 13028 13832 13084
rect 13832 13028 13836 13084
rect 13772 13024 13836 13028
rect 13852 13084 13916 13088
rect 13852 13028 13856 13084
rect 13856 13028 13912 13084
rect 13912 13028 13916 13084
rect 13852 13024 13916 13028
rect 952 12540 1016 12544
rect 952 12484 956 12540
rect 956 12484 1012 12540
rect 1012 12484 1016 12540
rect 952 12480 1016 12484
rect 1032 12540 1096 12544
rect 1032 12484 1036 12540
rect 1036 12484 1092 12540
rect 1092 12484 1096 12540
rect 1032 12480 1096 12484
rect 1112 12540 1176 12544
rect 1112 12484 1116 12540
rect 1116 12484 1172 12540
rect 1172 12484 1176 12540
rect 1112 12480 1176 12484
rect 1192 12540 1256 12544
rect 1192 12484 1196 12540
rect 1196 12484 1252 12540
rect 1252 12484 1256 12540
rect 1192 12480 1256 12484
rect 4952 12540 5016 12544
rect 4952 12484 4956 12540
rect 4956 12484 5012 12540
rect 5012 12484 5016 12540
rect 4952 12480 5016 12484
rect 5032 12540 5096 12544
rect 5032 12484 5036 12540
rect 5036 12484 5092 12540
rect 5092 12484 5096 12540
rect 5032 12480 5096 12484
rect 5112 12540 5176 12544
rect 5112 12484 5116 12540
rect 5116 12484 5172 12540
rect 5172 12484 5176 12540
rect 5112 12480 5176 12484
rect 5192 12540 5256 12544
rect 5192 12484 5196 12540
rect 5196 12484 5252 12540
rect 5252 12484 5256 12540
rect 5192 12480 5256 12484
rect 8952 12540 9016 12544
rect 8952 12484 8956 12540
rect 8956 12484 9012 12540
rect 9012 12484 9016 12540
rect 8952 12480 9016 12484
rect 9032 12540 9096 12544
rect 9032 12484 9036 12540
rect 9036 12484 9092 12540
rect 9092 12484 9096 12540
rect 9032 12480 9096 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 1612 11996 1676 12000
rect 1612 11940 1616 11996
rect 1616 11940 1672 11996
rect 1672 11940 1676 11996
rect 1612 11936 1676 11940
rect 1692 11996 1756 12000
rect 1692 11940 1696 11996
rect 1696 11940 1752 11996
rect 1752 11940 1756 11996
rect 1692 11936 1756 11940
rect 1772 11996 1836 12000
rect 1772 11940 1776 11996
rect 1776 11940 1832 11996
rect 1832 11940 1836 11996
rect 1772 11936 1836 11940
rect 1852 11996 1916 12000
rect 1852 11940 1856 11996
rect 1856 11940 1912 11996
rect 1912 11940 1916 11996
rect 1852 11936 1916 11940
rect 5612 11996 5676 12000
rect 5612 11940 5616 11996
rect 5616 11940 5672 11996
rect 5672 11940 5676 11996
rect 5612 11936 5676 11940
rect 5692 11996 5756 12000
rect 5692 11940 5696 11996
rect 5696 11940 5752 11996
rect 5752 11940 5756 11996
rect 5692 11936 5756 11940
rect 5772 11996 5836 12000
rect 5772 11940 5776 11996
rect 5776 11940 5832 11996
rect 5832 11940 5836 11996
rect 5772 11936 5836 11940
rect 5852 11996 5916 12000
rect 5852 11940 5856 11996
rect 5856 11940 5912 11996
rect 5912 11940 5916 11996
rect 5852 11936 5916 11940
rect 9612 11996 9676 12000
rect 9612 11940 9616 11996
rect 9616 11940 9672 11996
rect 9672 11940 9676 11996
rect 9612 11936 9676 11940
rect 9692 11996 9756 12000
rect 9692 11940 9696 11996
rect 9696 11940 9752 11996
rect 9752 11940 9756 11996
rect 9692 11936 9756 11940
rect 9772 11996 9836 12000
rect 9772 11940 9776 11996
rect 9776 11940 9832 11996
rect 9832 11940 9836 11996
rect 9772 11936 9836 11940
rect 9852 11996 9916 12000
rect 9852 11940 9856 11996
rect 9856 11940 9912 11996
rect 9912 11940 9916 11996
rect 9852 11936 9916 11940
rect 13612 11996 13676 12000
rect 13612 11940 13616 11996
rect 13616 11940 13672 11996
rect 13672 11940 13676 11996
rect 13612 11936 13676 11940
rect 13692 11996 13756 12000
rect 13692 11940 13696 11996
rect 13696 11940 13752 11996
rect 13752 11940 13756 11996
rect 13692 11936 13756 11940
rect 13772 11996 13836 12000
rect 13772 11940 13776 11996
rect 13776 11940 13832 11996
rect 13832 11940 13836 11996
rect 13772 11936 13836 11940
rect 13852 11996 13916 12000
rect 13852 11940 13856 11996
rect 13856 11940 13912 11996
rect 13912 11940 13916 11996
rect 13852 11936 13916 11940
rect 952 11452 1016 11456
rect 952 11396 956 11452
rect 956 11396 1012 11452
rect 1012 11396 1016 11452
rect 952 11392 1016 11396
rect 1032 11452 1096 11456
rect 1032 11396 1036 11452
rect 1036 11396 1092 11452
rect 1092 11396 1096 11452
rect 1032 11392 1096 11396
rect 1112 11452 1176 11456
rect 1112 11396 1116 11452
rect 1116 11396 1172 11452
rect 1172 11396 1176 11452
rect 1112 11392 1176 11396
rect 1192 11452 1256 11456
rect 1192 11396 1196 11452
rect 1196 11396 1252 11452
rect 1252 11396 1256 11452
rect 1192 11392 1256 11396
rect 4952 11452 5016 11456
rect 4952 11396 4956 11452
rect 4956 11396 5012 11452
rect 5012 11396 5016 11452
rect 4952 11392 5016 11396
rect 5032 11452 5096 11456
rect 5032 11396 5036 11452
rect 5036 11396 5092 11452
rect 5092 11396 5096 11452
rect 5032 11392 5096 11396
rect 5112 11452 5176 11456
rect 5112 11396 5116 11452
rect 5116 11396 5172 11452
rect 5172 11396 5176 11452
rect 5112 11392 5176 11396
rect 5192 11452 5256 11456
rect 5192 11396 5196 11452
rect 5196 11396 5252 11452
rect 5252 11396 5256 11452
rect 5192 11392 5256 11396
rect 8952 11452 9016 11456
rect 8952 11396 8956 11452
rect 8956 11396 9012 11452
rect 9012 11396 9016 11452
rect 8952 11392 9016 11396
rect 9032 11452 9096 11456
rect 9032 11396 9036 11452
rect 9036 11396 9092 11452
rect 9092 11396 9096 11452
rect 9032 11392 9096 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 1612 10908 1676 10912
rect 1612 10852 1616 10908
rect 1616 10852 1672 10908
rect 1672 10852 1676 10908
rect 1612 10848 1676 10852
rect 1692 10908 1756 10912
rect 1692 10852 1696 10908
rect 1696 10852 1752 10908
rect 1752 10852 1756 10908
rect 1692 10848 1756 10852
rect 1772 10908 1836 10912
rect 1772 10852 1776 10908
rect 1776 10852 1832 10908
rect 1832 10852 1836 10908
rect 1772 10848 1836 10852
rect 1852 10908 1916 10912
rect 1852 10852 1856 10908
rect 1856 10852 1912 10908
rect 1912 10852 1916 10908
rect 1852 10848 1916 10852
rect 5612 10908 5676 10912
rect 5612 10852 5616 10908
rect 5616 10852 5672 10908
rect 5672 10852 5676 10908
rect 5612 10848 5676 10852
rect 5692 10908 5756 10912
rect 5692 10852 5696 10908
rect 5696 10852 5752 10908
rect 5752 10852 5756 10908
rect 5692 10848 5756 10852
rect 5772 10908 5836 10912
rect 5772 10852 5776 10908
rect 5776 10852 5832 10908
rect 5832 10852 5836 10908
rect 5772 10848 5836 10852
rect 5852 10908 5916 10912
rect 5852 10852 5856 10908
rect 5856 10852 5912 10908
rect 5912 10852 5916 10908
rect 5852 10848 5916 10852
rect 9612 10908 9676 10912
rect 9612 10852 9616 10908
rect 9616 10852 9672 10908
rect 9672 10852 9676 10908
rect 9612 10848 9676 10852
rect 9692 10908 9756 10912
rect 9692 10852 9696 10908
rect 9696 10852 9752 10908
rect 9752 10852 9756 10908
rect 9692 10848 9756 10852
rect 9772 10908 9836 10912
rect 9772 10852 9776 10908
rect 9776 10852 9832 10908
rect 9832 10852 9836 10908
rect 9772 10848 9836 10852
rect 9852 10908 9916 10912
rect 9852 10852 9856 10908
rect 9856 10852 9912 10908
rect 9912 10852 9916 10908
rect 9852 10848 9916 10852
rect 13612 10908 13676 10912
rect 13612 10852 13616 10908
rect 13616 10852 13672 10908
rect 13672 10852 13676 10908
rect 13612 10848 13676 10852
rect 13692 10908 13756 10912
rect 13692 10852 13696 10908
rect 13696 10852 13752 10908
rect 13752 10852 13756 10908
rect 13692 10848 13756 10852
rect 13772 10908 13836 10912
rect 13772 10852 13776 10908
rect 13776 10852 13832 10908
rect 13832 10852 13836 10908
rect 13772 10848 13836 10852
rect 13852 10908 13916 10912
rect 13852 10852 13856 10908
rect 13856 10852 13912 10908
rect 13912 10852 13916 10908
rect 13852 10848 13916 10852
rect 952 10364 1016 10368
rect 952 10308 956 10364
rect 956 10308 1012 10364
rect 1012 10308 1016 10364
rect 952 10304 1016 10308
rect 1032 10364 1096 10368
rect 1032 10308 1036 10364
rect 1036 10308 1092 10364
rect 1092 10308 1096 10364
rect 1032 10304 1096 10308
rect 1112 10364 1176 10368
rect 1112 10308 1116 10364
rect 1116 10308 1172 10364
rect 1172 10308 1176 10364
rect 1112 10304 1176 10308
rect 1192 10364 1256 10368
rect 1192 10308 1196 10364
rect 1196 10308 1252 10364
rect 1252 10308 1256 10364
rect 1192 10304 1256 10308
rect 4952 10364 5016 10368
rect 4952 10308 4956 10364
rect 4956 10308 5012 10364
rect 5012 10308 5016 10364
rect 4952 10304 5016 10308
rect 5032 10364 5096 10368
rect 5032 10308 5036 10364
rect 5036 10308 5092 10364
rect 5092 10308 5096 10364
rect 5032 10304 5096 10308
rect 5112 10364 5176 10368
rect 5112 10308 5116 10364
rect 5116 10308 5172 10364
rect 5172 10308 5176 10364
rect 5112 10304 5176 10308
rect 5192 10364 5256 10368
rect 5192 10308 5196 10364
rect 5196 10308 5252 10364
rect 5252 10308 5256 10364
rect 5192 10304 5256 10308
rect 8952 10364 9016 10368
rect 8952 10308 8956 10364
rect 8956 10308 9012 10364
rect 9012 10308 9016 10364
rect 8952 10304 9016 10308
rect 9032 10364 9096 10368
rect 9032 10308 9036 10364
rect 9036 10308 9092 10364
rect 9092 10308 9096 10364
rect 9032 10304 9096 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 1612 9820 1676 9824
rect 1612 9764 1616 9820
rect 1616 9764 1672 9820
rect 1672 9764 1676 9820
rect 1612 9760 1676 9764
rect 1692 9820 1756 9824
rect 1692 9764 1696 9820
rect 1696 9764 1752 9820
rect 1752 9764 1756 9820
rect 1692 9760 1756 9764
rect 1772 9820 1836 9824
rect 1772 9764 1776 9820
rect 1776 9764 1832 9820
rect 1832 9764 1836 9820
rect 1772 9760 1836 9764
rect 1852 9820 1916 9824
rect 1852 9764 1856 9820
rect 1856 9764 1912 9820
rect 1912 9764 1916 9820
rect 1852 9760 1916 9764
rect 5612 9820 5676 9824
rect 5612 9764 5616 9820
rect 5616 9764 5672 9820
rect 5672 9764 5676 9820
rect 5612 9760 5676 9764
rect 5692 9820 5756 9824
rect 5692 9764 5696 9820
rect 5696 9764 5752 9820
rect 5752 9764 5756 9820
rect 5692 9760 5756 9764
rect 5772 9820 5836 9824
rect 5772 9764 5776 9820
rect 5776 9764 5832 9820
rect 5832 9764 5836 9820
rect 5772 9760 5836 9764
rect 5852 9820 5916 9824
rect 5852 9764 5856 9820
rect 5856 9764 5912 9820
rect 5912 9764 5916 9820
rect 5852 9760 5916 9764
rect 9612 9820 9676 9824
rect 9612 9764 9616 9820
rect 9616 9764 9672 9820
rect 9672 9764 9676 9820
rect 9612 9760 9676 9764
rect 9692 9820 9756 9824
rect 9692 9764 9696 9820
rect 9696 9764 9752 9820
rect 9752 9764 9756 9820
rect 9692 9760 9756 9764
rect 9772 9820 9836 9824
rect 9772 9764 9776 9820
rect 9776 9764 9832 9820
rect 9832 9764 9836 9820
rect 9772 9760 9836 9764
rect 9852 9820 9916 9824
rect 9852 9764 9856 9820
rect 9856 9764 9912 9820
rect 9912 9764 9916 9820
rect 9852 9760 9916 9764
rect 13612 9820 13676 9824
rect 13612 9764 13616 9820
rect 13616 9764 13672 9820
rect 13672 9764 13676 9820
rect 13612 9760 13676 9764
rect 13692 9820 13756 9824
rect 13692 9764 13696 9820
rect 13696 9764 13752 9820
rect 13752 9764 13756 9820
rect 13692 9760 13756 9764
rect 13772 9820 13836 9824
rect 13772 9764 13776 9820
rect 13776 9764 13832 9820
rect 13832 9764 13836 9820
rect 13772 9760 13836 9764
rect 13852 9820 13916 9824
rect 13852 9764 13856 9820
rect 13856 9764 13912 9820
rect 13912 9764 13916 9820
rect 13852 9760 13916 9764
rect 952 9276 1016 9280
rect 952 9220 956 9276
rect 956 9220 1012 9276
rect 1012 9220 1016 9276
rect 952 9216 1016 9220
rect 1032 9276 1096 9280
rect 1032 9220 1036 9276
rect 1036 9220 1092 9276
rect 1092 9220 1096 9276
rect 1032 9216 1096 9220
rect 1112 9276 1176 9280
rect 1112 9220 1116 9276
rect 1116 9220 1172 9276
rect 1172 9220 1176 9276
rect 1112 9216 1176 9220
rect 1192 9276 1256 9280
rect 1192 9220 1196 9276
rect 1196 9220 1252 9276
rect 1252 9220 1256 9276
rect 1192 9216 1256 9220
rect 4952 9276 5016 9280
rect 4952 9220 4956 9276
rect 4956 9220 5012 9276
rect 5012 9220 5016 9276
rect 4952 9216 5016 9220
rect 5032 9276 5096 9280
rect 5032 9220 5036 9276
rect 5036 9220 5092 9276
rect 5092 9220 5096 9276
rect 5032 9216 5096 9220
rect 5112 9276 5176 9280
rect 5112 9220 5116 9276
rect 5116 9220 5172 9276
rect 5172 9220 5176 9276
rect 5112 9216 5176 9220
rect 5192 9276 5256 9280
rect 5192 9220 5196 9276
rect 5196 9220 5252 9276
rect 5252 9220 5256 9276
rect 5192 9216 5256 9220
rect 8952 9276 9016 9280
rect 8952 9220 8956 9276
rect 8956 9220 9012 9276
rect 9012 9220 9016 9276
rect 8952 9216 9016 9220
rect 9032 9276 9096 9280
rect 9032 9220 9036 9276
rect 9036 9220 9092 9276
rect 9092 9220 9096 9276
rect 9032 9216 9096 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 1612 8732 1676 8736
rect 1612 8676 1616 8732
rect 1616 8676 1672 8732
rect 1672 8676 1676 8732
rect 1612 8672 1676 8676
rect 1692 8732 1756 8736
rect 1692 8676 1696 8732
rect 1696 8676 1752 8732
rect 1752 8676 1756 8732
rect 1692 8672 1756 8676
rect 1772 8732 1836 8736
rect 1772 8676 1776 8732
rect 1776 8676 1832 8732
rect 1832 8676 1836 8732
rect 1772 8672 1836 8676
rect 1852 8732 1916 8736
rect 1852 8676 1856 8732
rect 1856 8676 1912 8732
rect 1912 8676 1916 8732
rect 1852 8672 1916 8676
rect 5612 8732 5676 8736
rect 5612 8676 5616 8732
rect 5616 8676 5672 8732
rect 5672 8676 5676 8732
rect 5612 8672 5676 8676
rect 5692 8732 5756 8736
rect 5692 8676 5696 8732
rect 5696 8676 5752 8732
rect 5752 8676 5756 8732
rect 5692 8672 5756 8676
rect 5772 8732 5836 8736
rect 5772 8676 5776 8732
rect 5776 8676 5832 8732
rect 5832 8676 5836 8732
rect 5772 8672 5836 8676
rect 5852 8732 5916 8736
rect 5852 8676 5856 8732
rect 5856 8676 5912 8732
rect 5912 8676 5916 8732
rect 5852 8672 5916 8676
rect 9612 8732 9676 8736
rect 9612 8676 9616 8732
rect 9616 8676 9672 8732
rect 9672 8676 9676 8732
rect 9612 8672 9676 8676
rect 9692 8732 9756 8736
rect 9692 8676 9696 8732
rect 9696 8676 9752 8732
rect 9752 8676 9756 8732
rect 9692 8672 9756 8676
rect 9772 8732 9836 8736
rect 9772 8676 9776 8732
rect 9776 8676 9832 8732
rect 9832 8676 9836 8732
rect 9772 8672 9836 8676
rect 9852 8732 9916 8736
rect 9852 8676 9856 8732
rect 9856 8676 9912 8732
rect 9912 8676 9916 8732
rect 9852 8672 9916 8676
rect 13612 8732 13676 8736
rect 13612 8676 13616 8732
rect 13616 8676 13672 8732
rect 13672 8676 13676 8732
rect 13612 8672 13676 8676
rect 13692 8732 13756 8736
rect 13692 8676 13696 8732
rect 13696 8676 13752 8732
rect 13752 8676 13756 8732
rect 13692 8672 13756 8676
rect 13772 8732 13836 8736
rect 13772 8676 13776 8732
rect 13776 8676 13832 8732
rect 13832 8676 13836 8732
rect 13772 8672 13836 8676
rect 13852 8732 13916 8736
rect 13852 8676 13856 8732
rect 13856 8676 13912 8732
rect 13912 8676 13916 8732
rect 13852 8672 13916 8676
rect 952 8188 1016 8192
rect 952 8132 956 8188
rect 956 8132 1012 8188
rect 1012 8132 1016 8188
rect 952 8128 1016 8132
rect 1032 8188 1096 8192
rect 1032 8132 1036 8188
rect 1036 8132 1092 8188
rect 1092 8132 1096 8188
rect 1032 8128 1096 8132
rect 1112 8188 1176 8192
rect 1112 8132 1116 8188
rect 1116 8132 1172 8188
rect 1172 8132 1176 8188
rect 1112 8128 1176 8132
rect 1192 8188 1256 8192
rect 1192 8132 1196 8188
rect 1196 8132 1252 8188
rect 1252 8132 1256 8188
rect 1192 8128 1256 8132
rect 4952 8188 5016 8192
rect 4952 8132 4956 8188
rect 4956 8132 5012 8188
rect 5012 8132 5016 8188
rect 4952 8128 5016 8132
rect 5032 8188 5096 8192
rect 5032 8132 5036 8188
rect 5036 8132 5092 8188
rect 5092 8132 5096 8188
rect 5032 8128 5096 8132
rect 5112 8188 5176 8192
rect 5112 8132 5116 8188
rect 5116 8132 5172 8188
rect 5172 8132 5176 8188
rect 5112 8128 5176 8132
rect 5192 8188 5256 8192
rect 5192 8132 5196 8188
rect 5196 8132 5252 8188
rect 5252 8132 5256 8188
rect 5192 8128 5256 8132
rect 8952 8188 9016 8192
rect 8952 8132 8956 8188
rect 8956 8132 9012 8188
rect 9012 8132 9016 8188
rect 8952 8128 9016 8132
rect 9032 8188 9096 8192
rect 9032 8132 9036 8188
rect 9036 8132 9092 8188
rect 9092 8132 9096 8188
rect 9032 8128 9096 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 1612 7644 1676 7648
rect 1612 7588 1616 7644
rect 1616 7588 1672 7644
rect 1672 7588 1676 7644
rect 1612 7584 1676 7588
rect 1692 7644 1756 7648
rect 1692 7588 1696 7644
rect 1696 7588 1752 7644
rect 1752 7588 1756 7644
rect 1692 7584 1756 7588
rect 1772 7644 1836 7648
rect 1772 7588 1776 7644
rect 1776 7588 1832 7644
rect 1832 7588 1836 7644
rect 1772 7584 1836 7588
rect 1852 7644 1916 7648
rect 1852 7588 1856 7644
rect 1856 7588 1912 7644
rect 1912 7588 1916 7644
rect 1852 7584 1916 7588
rect 5612 7644 5676 7648
rect 5612 7588 5616 7644
rect 5616 7588 5672 7644
rect 5672 7588 5676 7644
rect 5612 7584 5676 7588
rect 5692 7644 5756 7648
rect 5692 7588 5696 7644
rect 5696 7588 5752 7644
rect 5752 7588 5756 7644
rect 5692 7584 5756 7588
rect 5772 7644 5836 7648
rect 5772 7588 5776 7644
rect 5776 7588 5832 7644
rect 5832 7588 5836 7644
rect 5772 7584 5836 7588
rect 5852 7644 5916 7648
rect 5852 7588 5856 7644
rect 5856 7588 5912 7644
rect 5912 7588 5916 7644
rect 5852 7584 5916 7588
rect 9612 7644 9676 7648
rect 9612 7588 9616 7644
rect 9616 7588 9672 7644
rect 9672 7588 9676 7644
rect 9612 7584 9676 7588
rect 9692 7644 9756 7648
rect 9692 7588 9696 7644
rect 9696 7588 9752 7644
rect 9752 7588 9756 7644
rect 9692 7584 9756 7588
rect 9772 7644 9836 7648
rect 9772 7588 9776 7644
rect 9776 7588 9832 7644
rect 9832 7588 9836 7644
rect 9772 7584 9836 7588
rect 9852 7644 9916 7648
rect 9852 7588 9856 7644
rect 9856 7588 9912 7644
rect 9912 7588 9916 7644
rect 9852 7584 9916 7588
rect 13612 7644 13676 7648
rect 13612 7588 13616 7644
rect 13616 7588 13672 7644
rect 13672 7588 13676 7644
rect 13612 7584 13676 7588
rect 13692 7644 13756 7648
rect 13692 7588 13696 7644
rect 13696 7588 13752 7644
rect 13752 7588 13756 7644
rect 13692 7584 13756 7588
rect 13772 7644 13836 7648
rect 13772 7588 13776 7644
rect 13776 7588 13832 7644
rect 13832 7588 13836 7644
rect 13772 7584 13836 7588
rect 13852 7644 13916 7648
rect 13852 7588 13856 7644
rect 13856 7588 13912 7644
rect 13912 7588 13916 7644
rect 13852 7584 13916 7588
rect 952 7100 1016 7104
rect 952 7044 956 7100
rect 956 7044 1012 7100
rect 1012 7044 1016 7100
rect 952 7040 1016 7044
rect 1032 7100 1096 7104
rect 1032 7044 1036 7100
rect 1036 7044 1092 7100
rect 1092 7044 1096 7100
rect 1032 7040 1096 7044
rect 1112 7100 1176 7104
rect 1112 7044 1116 7100
rect 1116 7044 1172 7100
rect 1172 7044 1176 7100
rect 1112 7040 1176 7044
rect 1192 7100 1256 7104
rect 1192 7044 1196 7100
rect 1196 7044 1252 7100
rect 1252 7044 1256 7100
rect 1192 7040 1256 7044
rect 4952 7100 5016 7104
rect 4952 7044 4956 7100
rect 4956 7044 5012 7100
rect 5012 7044 5016 7100
rect 4952 7040 5016 7044
rect 5032 7100 5096 7104
rect 5032 7044 5036 7100
rect 5036 7044 5092 7100
rect 5092 7044 5096 7100
rect 5032 7040 5096 7044
rect 5112 7100 5176 7104
rect 5112 7044 5116 7100
rect 5116 7044 5172 7100
rect 5172 7044 5176 7100
rect 5112 7040 5176 7044
rect 5192 7100 5256 7104
rect 5192 7044 5196 7100
rect 5196 7044 5252 7100
rect 5252 7044 5256 7100
rect 5192 7040 5256 7044
rect 8952 7100 9016 7104
rect 8952 7044 8956 7100
rect 8956 7044 9012 7100
rect 9012 7044 9016 7100
rect 8952 7040 9016 7044
rect 9032 7100 9096 7104
rect 9032 7044 9036 7100
rect 9036 7044 9092 7100
rect 9092 7044 9096 7100
rect 9032 7040 9096 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 1612 6556 1676 6560
rect 1612 6500 1616 6556
rect 1616 6500 1672 6556
rect 1672 6500 1676 6556
rect 1612 6496 1676 6500
rect 1692 6556 1756 6560
rect 1692 6500 1696 6556
rect 1696 6500 1752 6556
rect 1752 6500 1756 6556
rect 1692 6496 1756 6500
rect 1772 6556 1836 6560
rect 1772 6500 1776 6556
rect 1776 6500 1832 6556
rect 1832 6500 1836 6556
rect 1772 6496 1836 6500
rect 1852 6556 1916 6560
rect 1852 6500 1856 6556
rect 1856 6500 1912 6556
rect 1912 6500 1916 6556
rect 1852 6496 1916 6500
rect 5612 6556 5676 6560
rect 5612 6500 5616 6556
rect 5616 6500 5672 6556
rect 5672 6500 5676 6556
rect 5612 6496 5676 6500
rect 5692 6556 5756 6560
rect 5692 6500 5696 6556
rect 5696 6500 5752 6556
rect 5752 6500 5756 6556
rect 5692 6496 5756 6500
rect 5772 6556 5836 6560
rect 5772 6500 5776 6556
rect 5776 6500 5832 6556
rect 5832 6500 5836 6556
rect 5772 6496 5836 6500
rect 5852 6556 5916 6560
rect 5852 6500 5856 6556
rect 5856 6500 5912 6556
rect 5912 6500 5916 6556
rect 5852 6496 5916 6500
rect 9612 6556 9676 6560
rect 9612 6500 9616 6556
rect 9616 6500 9672 6556
rect 9672 6500 9676 6556
rect 9612 6496 9676 6500
rect 9692 6556 9756 6560
rect 9692 6500 9696 6556
rect 9696 6500 9752 6556
rect 9752 6500 9756 6556
rect 9692 6496 9756 6500
rect 9772 6556 9836 6560
rect 9772 6500 9776 6556
rect 9776 6500 9832 6556
rect 9832 6500 9836 6556
rect 9772 6496 9836 6500
rect 9852 6556 9916 6560
rect 9852 6500 9856 6556
rect 9856 6500 9912 6556
rect 9912 6500 9916 6556
rect 9852 6496 9916 6500
rect 13612 6556 13676 6560
rect 13612 6500 13616 6556
rect 13616 6500 13672 6556
rect 13672 6500 13676 6556
rect 13612 6496 13676 6500
rect 13692 6556 13756 6560
rect 13692 6500 13696 6556
rect 13696 6500 13752 6556
rect 13752 6500 13756 6556
rect 13692 6496 13756 6500
rect 13772 6556 13836 6560
rect 13772 6500 13776 6556
rect 13776 6500 13832 6556
rect 13832 6500 13836 6556
rect 13772 6496 13836 6500
rect 13852 6556 13916 6560
rect 13852 6500 13856 6556
rect 13856 6500 13912 6556
rect 13912 6500 13916 6556
rect 13852 6496 13916 6500
rect 952 6012 1016 6016
rect 952 5956 956 6012
rect 956 5956 1012 6012
rect 1012 5956 1016 6012
rect 952 5952 1016 5956
rect 1032 6012 1096 6016
rect 1032 5956 1036 6012
rect 1036 5956 1092 6012
rect 1092 5956 1096 6012
rect 1032 5952 1096 5956
rect 1112 6012 1176 6016
rect 1112 5956 1116 6012
rect 1116 5956 1172 6012
rect 1172 5956 1176 6012
rect 1112 5952 1176 5956
rect 1192 6012 1256 6016
rect 1192 5956 1196 6012
rect 1196 5956 1252 6012
rect 1252 5956 1256 6012
rect 1192 5952 1256 5956
rect 4952 6012 5016 6016
rect 4952 5956 4956 6012
rect 4956 5956 5012 6012
rect 5012 5956 5016 6012
rect 4952 5952 5016 5956
rect 5032 6012 5096 6016
rect 5032 5956 5036 6012
rect 5036 5956 5092 6012
rect 5092 5956 5096 6012
rect 5032 5952 5096 5956
rect 5112 6012 5176 6016
rect 5112 5956 5116 6012
rect 5116 5956 5172 6012
rect 5172 5956 5176 6012
rect 5112 5952 5176 5956
rect 5192 6012 5256 6016
rect 5192 5956 5196 6012
rect 5196 5956 5252 6012
rect 5252 5956 5256 6012
rect 5192 5952 5256 5956
rect 8952 6012 9016 6016
rect 8952 5956 8956 6012
rect 8956 5956 9012 6012
rect 9012 5956 9016 6012
rect 8952 5952 9016 5956
rect 9032 6012 9096 6016
rect 9032 5956 9036 6012
rect 9036 5956 9092 6012
rect 9092 5956 9096 6012
rect 9032 5952 9096 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 1612 5468 1676 5472
rect 1612 5412 1616 5468
rect 1616 5412 1672 5468
rect 1672 5412 1676 5468
rect 1612 5408 1676 5412
rect 1692 5468 1756 5472
rect 1692 5412 1696 5468
rect 1696 5412 1752 5468
rect 1752 5412 1756 5468
rect 1692 5408 1756 5412
rect 1772 5468 1836 5472
rect 1772 5412 1776 5468
rect 1776 5412 1832 5468
rect 1832 5412 1836 5468
rect 1772 5408 1836 5412
rect 1852 5468 1916 5472
rect 1852 5412 1856 5468
rect 1856 5412 1912 5468
rect 1912 5412 1916 5468
rect 1852 5408 1916 5412
rect 5612 5468 5676 5472
rect 5612 5412 5616 5468
rect 5616 5412 5672 5468
rect 5672 5412 5676 5468
rect 5612 5408 5676 5412
rect 5692 5468 5756 5472
rect 5692 5412 5696 5468
rect 5696 5412 5752 5468
rect 5752 5412 5756 5468
rect 5692 5408 5756 5412
rect 5772 5468 5836 5472
rect 5772 5412 5776 5468
rect 5776 5412 5832 5468
rect 5832 5412 5836 5468
rect 5772 5408 5836 5412
rect 5852 5468 5916 5472
rect 5852 5412 5856 5468
rect 5856 5412 5912 5468
rect 5912 5412 5916 5468
rect 5852 5408 5916 5412
rect 9612 5468 9676 5472
rect 9612 5412 9616 5468
rect 9616 5412 9672 5468
rect 9672 5412 9676 5468
rect 9612 5408 9676 5412
rect 9692 5468 9756 5472
rect 9692 5412 9696 5468
rect 9696 5412 9752 5468
rect 9752 5412 9756 5468
rect 9692 5408 9756 5412
rect 9772 5468 9836 5472
rect 9772 5412 9776 5468
rect 9776 5412 9832 5468
rect 9832 5412 9836 5468
rect 9772 5408 9836 5412
rect 9852 5468 9916 5472
rect 9852 5412 9856 5468
rect 9856 5412 9912 5468
rect 9912 5412 9916 5468
rect 9852 5408 9916 5412
rect 13612 5468 13676 5472
rect 13612 5412 13616 5468
rect 13616 5412 13672 5468
rect 13672 5412 13676 5468
rect 13612 5408 13676 5412
rect 13692 5468 13756 5472
rect 13692 5412 13696 5468
rect 13696 5412 13752 5468
rect 13752 5412 13756 5468
rect 13692 5408 13756 5412
rect 13772 5468 13836 5472
rect 13772 5412 13776 5468
rect 13776 5412 13832 5468
rect 13832 5412 13836 5468
rect 13772 5408 13836 5412
rect 13852 5468 13916 5472
rect 13852 5412 13856 5468
rect 13856 5412 13912 5468
rect 13912 5412 13916 5468
rect 13852 5408 13916 5412
rect 952 4924 1016 4928
rect 952 4868 956 4924
rect 956 4868 1012 4924
rect 1012 4868 1016 4924
rect 952 4864 1016 4868
rect 1032 4924 1096 4928
rect 1032 4868 1036 4924
rect 1036 4868 1092 4924
rect 1092 4868 1096 4924
rect 1032 4864 1096 4868
rect 1112 4924 1176 4928
rect 1112 4868 1116 4924
rect 1116 4868 1172 4924
rect 1172 4868 1176 4924
rect 1112 4864 1176 4868
rect 1192 4924 1256 4928
rect 1192 4868 1196 4924
rect 1196 4868 1252 4924
rect 1252 4868 1256 4924
rect 1192 4864 1256 4868
rect 4952 4924 5016 4928
rect 4952 4868 4956 4924
rect 4956 4868 5012 4924
rect 5012 4868 5016 4924
rect 4952 4864 5016 4868
rect 5032 4924 5096 4928
rect 5032 4868 5036 4924
rect 5036 4868 5092 4924
rect 5092 4868 5096 4924
rect 5032 4864 5096 4868
rect 5112 4924 5176 4928
rect 5112 4868 5116 4924
rect 5116 4868 5172 4924
rect 5172 4868 5176 4924
rect 5112 4864 5176 4868
rect 5192 4924 5256 4928
rect 5192 4868 5196 4924
rect 5196 4868 5252 4924
rect 5252 4868 5256 4924
rect 5192 4864 5256 4868
rect 8952 4924 9016 4928
rect 8952 4868 8956 4924
rect 8956 4868 9012 4924
rect 9012 4868 9016 4924
rect 8952 4864 9016 4868
rect 9032 4924 9096 4928
rect 9032 4868 9036 4924
rect 9036 4868 9092 4924
rect 9092 4868 9096 4924
rect 9032 4864 9096 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 1612 4380 1676 4384
rect 1612 4324 1616 4380
rect 1616 4324 1672 4380
rect 1672 4324 1676 4380
rect 1612 4320 1676 4324
rect 1692 4380 1756 4384
rect 1692 4324 1696 4380
rect 1696 4324 1752 4380
rect 1752 4324 1756 4380
rect 1692 4320 1756 4324
rect 1772 4380 1836 4384
rect 1772 4324 1776 4380
rect 1776 4324 1832 4380
rect 1832 4324 1836 4380
rect 1772 4320 1836 4324
rect 1852 4380 1916 4384
rect 1852 4324 1856 4380
rect 1856 4324 1912 4380
rect 1912 4324 1916 4380
rect 1852 4320 1916 4324
rect 5612 4380 5676 4384
rect 5612 4324 5616 4380
rect 5616 4324 5672 4380
rect 5672 4324 5676 4380
rect 5612 4320 5676 4324
rect 5692 4380 5756 4384
rect 5692 4324 5696 4380
rect 5696 4324 5752 4380
rect 5752 4324 5756 4380
rect 5692 4320 5756 4324
rect 5772 4380 5836 4384
rect 5772 4324 5776 4380
rect 5776 4324 5832 4380
rect 5832 4324 5836 4380
rect 5772 4320 5836 4324
rect 5852 4380 5916 4384
rect 5852 4324 5856 4380
rect 5856 4324 5912 4380
rect 5912 4324 5916 4380
rect 5852 4320 5916 4324
rect 9612 4380 9676 4384
rect 9612 4324 9616 4380
rect 9616 4324 9672 4380
rect 9672 4324 9676 4380
rect 9612 4320 9676 4324
rect 9692 4380 9756 4384
rect 9692 4324 9696 4380
rect 9696 4324 9752 4380
rect 9752 4324 9756 4380
rect 9692 4320 9756 4324
rect 9772 4380 9836 4384
rect 9772 4324 9776 4380
rect 9776 4324 9832 4380
rect 9832 4324 9836 4380
rect 9772 4320 9836 4324
rect 9852 4380 9916 4384
rect 9852 4324 9856 4380
rect 9856 4324 9912 4380
rect 9912 4324 9916 4380
rect 9852 4320 9916 4324
rect 13612 4380 13676 4384
rect 13612 4324 13616 4380
rect 13616 4324 13672 4380
rect 13672 4324 13676 4380
rect 13612 4320 13676 4324
rect 13692 4380 13756 4384
rect 13692 4324 13696 4380
rect 13696 4324 13752 4380
rect 13752 4324 13756 4380
rect 13692 4320 13756 4324
rect 13772 4380 13836 4384
rect 13772 4324 13776 4380
rect 13776 4324 13832 4380
rect 13832 4324 13836 4380
rect 13772 4320 13836 4324
rect 13852 4380 13916 4384
rect 13852 4324 13856 4380
rect 13856 4324 13912 4380
rect 13912 4324 13916 4380
rect 13852 4320 13916 4324
rect 952 3836 1016 3840
rect 952 3780 956 3836
rect 956 3780 1012 3836
rect 1012 3780 1016 3836
rect 952 3776 1016 3780
rect 1032 3836 1096 3840
rect 1032 3780 1036 3836
rect 1036 3780 1092 3836
rect 1092 3780 1096 3836
rect 1032 3776 1096 3780
rect 1112 3836 1176 3840
rect 1112 3780 1116 3836
rect 1116 3780 1172 3836
rect 1172 3780 1176 3836
rect 1112 3776 1176 3780
rect 1192 3836 1256 3840
rect 1192 3780 1196 3836
rect 1196 3780 1252 3836
rect 1252 3780 1256 3836
rect 1192 3776 1256 3780
rect 4952 3836 5016 3840
rect 4952 3780 4956 3836
rect 4956 3780 5012 3836
rect 5012 3780 5016 3836
rect 4952 3776 5016 3780
rect 5032 3836 5096 3840
rect 5032 3780 5036 3836
rect 5036 3780 5092 3836
rect 5092 3780 5096 3836
rect 5032 3776 5096 3780
rect 5112 3836 5176 3840
rect 5112 3780 5116 3836
rect 5116 3780 5172 3836
rect 5172 3780 5176 3836
rect 5112 3776 5176 3780
rect 5192 3836 5256 3840
rect 5192 3780 5196 3836
rect 5196 3780 5252 3836
rect 5252 3780 5256 3836
rect 5192 3776 5256 3780
rect 8952 3836 9016 3840
rect 8952 3780 8956 3836
rect 8956 3780 9012 3836
rect 9012 3780 9016 3836
rect 8952 3776 9016 3780
rect 9032 3836 9096 3840
rect 9032 3780 9036 3836
rect 9036 3780 9092 3836
rect 9092 3780 9096 3836
rect 9032 3776 9096 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 1612 3292 1676 3296
rect 1612 3236 1616 3292
rect 1616 3236 1672 3292
rect 1672 3236 1676 3292
rect 1612 3232 1676 3236
rect 1692 3292 1756 3296
rect 1692 3236 1696 3292
rect 1696 3236 1752 3292
rect 1752 3236 1756 3292
rect 1692 3232 1756 3236
rect 1772 3292 1836 3296
rect 1772 3236 1776 3292
rect 1776 3236 1832 3292
rect 1832 3236 1836 3292
rect 1772 3232 1836 3236
rect 1852 3292 1916 3296
rect 1852 3236 1856 3292
rect 1856 3236 1912 3292
rect 1912 3236 1916 3292
rect 1852 3232 1916 3236
rect 5612 3292 5676 3296
rect 5612 3236 5616 3292
rect 5616 3236 5672 3292
rect 5672 3236 5676 3292
rect 5612 3232 5676 3236
rect 5692 3292 5756 3296
rect 5692 3236 5696 3292
rect 5696 3236 5752 3292
rect 5752 3236 5756 3292
rect 5692 3232 5756 3236
rect 5772 3292 5836 3296
rect 5772 3236 5776 3292
rect 5776 3236 5832 3292
rect 5832 3236 5836 3292
rect 5772 3232 5836 3236
rect 5852 3292 5916 3296
rect 5852 3236 5856 3292
rect 5856 3236 5912 3292
rect 5912 3236 5916 3292
rect 5852 3232 5916 3236
rect 9612 3292 9676 3296
rect 9612 3236 9616 3292
rect 9616 3236 9672 3292
rect 9672 3236 9676 3292
rect 9612 3232 9676 3236
rect 9692 3292 9756 3296
rect 9692 3236 9696 3292
rect 9696 3236 9752 3292
rect 9752 3236 9756 3292
rect 9692 3232 9756 3236
rect 9772 3292 9836 3296
rect 9772 3236 9776 3292
rect 9776 3236 9832 3292
rect 9832 3236 9836 3292
rect 9772 3232 9836 3236
rect 9852 3292 9916 3296
rect 9852 3236 9856 3292
rect 9856 3236 9912 3292
rect 9912 3236 9916 3292
rect 9852 3232 9916 3236
rect 13612 3292 13676 3296
rect 13612 3236 13616 3292
rect 13616 3236 13672 3292
rect 13672 3236 13676 3292
rect 13612 3232 13676 3236
rect 13692 3292 13756 3296
rect 13692 3236 13696 3292
rect 13696 3236 13752 3292
rect 13752 3236 13756 3292
rect 13692 3232 13756 3236
rect 13772 3292 13836 3296
rect 13772 3236 13776 3292
rect 13776 3236 13832 3292
rect 13832 3236 13836 3292
rect 13772 3232 13836 3236
rect 13852 3292 13916 3296
rect 13852 3236 13856 3292
rect 13856 3236 13912 3292
rect 13912 3236 13916 3292
rect 13852 3232 13916 3236
rect 952 2748 1016 2752
rect 952 2692 956 2748
rect 956 2692 1012 2748
rect 1012 2692 1016 2748
rect 952 2688 1016 2692
rect 1032 2748 1096 2752
rect 1032 2692 1036 2748
rect 1036 2692 1092 2748
rect 1092 2692 1096 2748
rect 1032 2688 1096 2692
rect 1112 2748 1176 2752
rect 1112 2692 1116 2748
rect 1116 2692 1172 2748
rect 1172 2692 1176 2748
rect 1112 2688 1176 2692
rect 1192 2748 1256 2752
rect 1192 2692 1196 2748
rect 1196 2692 1252 2748
rect 1252 2692 1256 2748
rect 1192 2688 1256 2692
rect 4952 2748 5016 2752
rect 4952 2692 4956 2748
rect 4956 2692 5012 2748
rect 5012 2692 5016 2748
rect 4952 2688 5016 2692
rect 5032 2748 5096 2752
rect 5032 2692 5036 2748
rect 5036 2692 5092 2748
rect 5092 2692 5096 2748
rect 5032 2688 5096 2692
rect 5112 2748 5176 2752
rect 5112 2692 5116 2748
rect 5116 2692 5172 2748
rect 5172 2692 5176 2748
rect 5112 2688 5176 2692
rect 5192 2748 5256 2752
rect 5192 2692 5196 2748
rect 5196 2692 5252 2748
rect 5252 2692 5256 2748
rect 5192 2688 5256 2692
rect 8952 2748 9016 2752
rect 8952 2692 8956 2748
rect 8956 2692 9012 2748
rect 9012 2692 9016 2748
rect 8952 2688 9016 2692
rect 9032 2748 9096 2752
rect 9032 2692 9036 2748
rect 9036 2692 9092 2748
rect 9092 2692 9096 2748
rect 9032 2688 9096 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 1612 2204 1676 2208
rect 1612 2148 1616 2204
rect 1616 2148 1672 2204
rect 1672 2148 1676 2204
rect 1612 2144 1676 2148
rect 1692 2204 1756 2208
rect 1692 2148 1696 2204
rect 1696 2148 1752 2204
rect 1752 2148 1756 2204
rect 1692 2144 1756 2148
rect 1772 2204 1836 2208
rect 1772 2148 1776 2204
rect 1776 2148 1832 2204
rect 1832 2148 1836 2204
rect 1772 2144 1836 2148
rect 1852 2204 1916 2208
rect 1852 2148 1856 2204
rect 1856 2148 1912 2204
rect 1912 2148 1916 2204
rect 1852 2144 1916 2148
rect 5612 2204 5676 2208
rect 5612 2148 5616 2204
rect 5616 2148 5672 2204
rect 5672 2148 5676 2204
rect 5612 2144 5676 2148
rect 5692 2204 5756 2208
rect 5692 2148 5696 2204
rect 5696 2148 5752 2204
rect 5752 2148 5756 2204
rect 5692 2144 5756 2148
rect 5772 2204 5836 2208
rect 5772 2148 5776 2204
rect 5776 2148 5832 2204
rect 5832 2148 5836 2204
rect 5772 2144 5836 2148
rect 5852 2204 5916 2208
rect 5852 2148 5856 2204
rect 5856 2148 5912 2204
rect 5912 2148 5916 2204
rect 5852 2144 5916 2148
rect 9612 2204 9676 2208
rect 9612 2148 9616 2204
rect 9616 2148 9672 2204
rect 9672 2148 9676 2204
rect 9612 2144 9676 2148
rect 9692 2204 9756 2208
rect 9692 2148 9696 2204
rect 9696 2148 9752 2204
rect 9752 2148 9756 2204
rect 9692 2144 9756 2148
rect 9772 2204 9836 2208
rect 9772 2148 9776 2204
rect 9776 2148 9832 2204
rect 9832 2148 9836 2204
rect 9772 2144 9836 2148
rect 9852 2204 9916 2208
rect 9852 2148 9856 2204
rect 9856 2148 9912 2204
rect 9912 2148 9916 2204
rect 9852 2144 9916 2148
rect 13612 2204 13676 2208
rect 13612 2148 13616 2204
rect 13616 2148 13672 2204
rect 13672 2148 13676 2204
rect 13612 2144 13676 2148
rect 13692 2204 13756 2208
rect 13692 2148 13696 2204
rect 13696 2148 13752 2204
rect 13752 2148 13756 2204
rect 13692 2144 13756 2148
rect 13772 2204 13836 2208
rect 13772 2148 13776 2204
rect 13776 2148 13832 2204
rect 13832 2148 13836 2204
rect 13772 2144 13836 2148
rect 13852 2204 13916 2208
rect 13852 2148 13856 2204
rect 13856 2148 13912 2204
rect 13912 2148 13916 2204
rect 13852 2144 13916 2148
<< metal4 >>
rect 944 15808 1264 15824
rect 944 15744 952 15808
rect 1016 15744 1032 15808
rect 1096 15744 1112 15808
rect 1176 15744 1192 15808
rect 1256 15744 1264 15808
rect 944 14720 1264 15744
rect 944 14656 952 14720
rect 1016 14656 1032 14720
rect 1096 14656 1112 14720
rect 1176 14656 1192 14720
rect 1256 14656 1264 14720
rect 944 14294 1264 14656
rect 944 14058 986 14294
rect 1222 14058 1264 14294
rect 944 13632 1264 14058
rect 944 13568 952 13632
rect 1016 13568 1032 13632
rect 1096 13568 1112 13632
rect 1176 13568 1192 13632
rect 1256 13568 1264 13632
rect 944 12544 1264 13568
rect 944 12480 952 12544
rect 1016 12480 1032 12544
rect 1096 12480 1112 12544
rect 1176 12480 1192 12544
rect 1256 12480 1264 12544
rect 944 11456 1264 12480
rect 944 11392 952 11456
rect 1016 11392 1032 11456
rect 1096 11392 1112 11456
rect 1176 11392 1192 11456
rect 1256 11392 1264 11456
rect 944 10368 1264 11392
rect 944 10304 952 10368
rect 1016 10304 1032 10368
rect 1096 10304 1112 10368
rect 1176 10304 1192 10368
rect 1256 10304 1264 10368
rect 944 10294 1264 10304
rect 944 10058 986 10294
rect 1222 10058 1264 10294
rect 944 9280 1264 10058
rect 944 9216 952 9280
rect 1016 9216 1032 9280
rect 1096 9216 1112 9280
rect 1176 9216 1192 9280
rect 1256 9216 1264 9280
rect 944 8192 1264 9216
rect 944 8128 952 8192
rect 1016 8128 1032 8192
rect 1096 8128 1112 8192
rect 1176 8128 1192 8192
rect 1256 8128 1264 8192
rect 944 7104 1264 8128
rect 944 7040 952 7104
rect 1016 7040 1032 7104
rect 1096 7040 1112 7104
rect 1176 7040 1192 7104
rect 1256 7040 1264 7104
rect 944 6294 1264 7040
rect 944 6058 986 6294
rect 1222 6058 1264 6294
rect 944 6016 1264 6058
rect 944 5952 952 6016
rect 1016 5952 1032 6016
rect 1096 5952 1112 6016
rect 1176 5952 1192 6016
rect 1256 5952 1264 6016
rect 944 4928 1264 5952
rect 944 4864 952 4928
rect 1016 4864 1032 4928
rect 1096 4864 1112 4928
rect 1176 4864 1192 4928
rect 1256 4864 1264 4928
rect 944 3840 1264 4864
rect 944 3776 952 3840
rect 1016 3776 1032 3840
rect 1096 3776 1112 3840
rect 1176 3776 1192 3840
rect 1256 3776 1264 3840
rect 944 2752 1264 3776
rect 944 2688 952 2752
rect 1016 2688 1032 2752
rect 1096 2688 1112 2752
rect 1176 2688 1192 2752
rect 1256 2688 1264 2752
rect 944 2294 1264 2688
rect 944 2058 986 2294
rect 1222 2058 1264 2294
rect 1604 15264 1924 15824
rect 1604 15200 1612 15264
rect 1676 15200 1692 15264
rect 1756 15200 1772 15264
rect 1836 15200 1852 15264
rect 1916 15200 1924 15264
rect 1604 14954 1924 15200
rect 1604 14718 1646 14954
rect 1882 14718 1924 14954
rect 1604 14176 1924 14718
rect 1604 14112 1612 14176
rect 1676 14112 1692 14176
rect 1756 14112 1772 14176
rect 1836 14112 1852 14176
rect 1916 14112 1924 14176
rect 1604 13088 1924 14112
rect 1604 13024 1612 13088
rect 1676 13024 1692 13088
rect 1756 13024 1772 13088
rect 1836 13024 1852 13088
rect 1916 13024 1924 13088
rect 1604 12000 1924 13024
rect 1604 11936 1612 12000
rect 1676 11936 1692 12000
rect 1756 11936 1772 12000
rect 1836 11936 1852 12000
rect 1916 11936 1924 12000
rect 1604 10954 1924 11936
rect 1604 10912 1646 10954
rect 1882 10912 1924 10954
rect 1604 10848 1612 10912
rect 1916 10848 1924 10912
rect 1604 10718 1646 10848
rect 1882 10718 1924 10848
rect 1604 9824 1924 10718
rect 1604 9760 1612 9824
rect 1676 9760 1692 9824
rect 1756 9760 1772 9824
rect 1836 9760 1852 9824
rect 1916 9760 1924 9824
rect 1604 8736 1924 9760
rect 1604 8672 1612 8736
rect 1676 8672 1692 8736
rect 1756 8672 1772 8736
rect 1836 8672 1852 8736
rect 1916 8672 1924 8736
rect 1604 7648 1924 8672
rect 1604 7584 1612 7648
rect 1676 7584 1692 7648
rect 1756 7584 1772 7648
rect 1836 7584 1852 7648
rect 1916 7584 1924 7648
rect 1604 6954 1924 7584
rect 1604 6718 1646 6954
rect 1882 6718 1924 6954
rect 1604 6560 1924 6718
rect 1604 6496 1612 6560
rect 1676 6496 1692 6560
rect 1756 6496 1772 6560
rect 1836 6496 1852 6560
rect 1916 6496 1924 6560
rect 1604 5472 1924 6496
rect 1604 5408 1612 5472
rect 1676 5408 1692 5472
rect 1756 5408 1772 5472
rect 1836 5408 1852 5472
rect 1916 5408 1924 5472
rect 1604 4384 1924 5408
rect 1604 4320 1612 4384
rect 1676 4320 1692 4384
rect 1756 4320 1772 4384
rect 1836 4320 1852 4384
rect 1916 4320 1924 4384
rect 1604 3296 1924 4320
rect 1604 3232 1612 3296
rect 1676 3232 1692 3296
rect 1756 3232 1772 3296
rect 1836 3232 1852 3296
rect 1916 3232 1924 3296
rect 1604 2954 1924 3232
rect 1604 2718 1646 2954
rect 1882 2718 1924 2954
rect 1604 2208 1924 2718
rect 1604 2144 1612 2208
rect 1676 2144 1692 2208
rect 1756 2144 1772 2208
rect 1836 2144 1852 2208
rect 1916 2144 1924 2208
rect 1604 2128 1924 2144
rect 4944 15808 5264 15824
rect 4944 15744 4952 15808
rect 5016 15744 5032 15808
rect 5096 15744 5112 15808
rect 5176 15744 5192 15808
rect 5256 15744 5264 15808
rect 4944 14720 5264 15744
rect 4944 14656 4952 14720
rect 5016 14656 5032 14720
rect 5096 14656 5112 14720
rect 5176 14656 5192 14720
rect 5256 14656 5264 14720
rect 4944 14294 5264 14656
rect 4944 14058 4986 14294
rect 5222 14058 5264 14294
rect 4944 13632 5264 14058
rect 4944 13568 4952 13632
rect 5016 13568 5032 13632
rect 5096 13568 5112 13632
rect 5176 13568 5192 13632
rect 5256 13568 5264 13632
rect 4944 12544 5264 13568
rect 4944 12480 4952 12544
rect 5016 12480 5032 12544
rect 5096 12480 5112 12544
rect 5176 12480 5192 12544
rect 5256 12480 5264 12544
rect 4944 11456 5264 12480
rect 4944 11392 4952 11456
rect 5016 11392 5032 11456
rect 5096 11392 5112 11456
rect 5176 11392 5192 11456
rect 5256 11392 5264 11456
rect 4944 10368 5264 11392
rect 4944 10304 4952 10368
rect 5016 10304 5032 10368
rect 5096 10304 5112 10368
rect 5176 10304 5192 10368
rect 5256 10304 5264 10368
rect 4944 10294 5264 10304
rect 4944 10058 4986 10294
rect 5222 10058 5264 10294
rect 4944 9280 5264 10058
rect 4944 9216 4952 9280
rect 5016 9216 5032 9280
rect 5096 9216 5112 9280
rect 5176 9216 5192 9280
rect 5256 9216 5264 9280
rect 4944 8192 5264 9216
rect 4944 8128 4952 8192
rect 5016 8128 5032 8192
rect 5096 8128 5112 8192
rect 5176 8128 5192 8192
rect 5256 8128 5264 8192
rect 4944 7104 5264 8128
rect 4944 7040 4952 7104
rect 5016 7040 5032 7104
rect 5096 7040 5112 7104
rect 5176 7040 5192 7104
rect 5256 7040 5264 7104
rect 4944 6294 5264 7040
rect 4944 6058 4986 6294
rect 5222 6058 5264 6294
rect 4944 6016 5264 6058
rect 4944 5952 4952 6016
rect 5016 5952 5032 6016
rect 5096 5952 5112 6016
rect 5176 5952 5192 6016
rect 5256 5952 5264 6016
rect 4944 4928 5264 5952
rect 4944 4864 4952 4928
rect 5016 4864 5032 4928
rect 5096 4864 5112 4928
rect 5176 4864 5192 4928
rect 5256 4864 5264 4928
rect 4944 3840 5264 4864
rect 4944 3776 4952 3840
rect 5016 3776 5032 3840
rect 5096 3776 5112 3840
rect 5176 3776 5192 3840
rect 5256 3776 5264 3840
rect 4944 2752 5264 3776
rect 4944 2688 4952 2752
rect 5016 2688 5032 2752
rect 5096 2688 5112 2752
rect 5176 2688 5192 2752
rect 5256 2688 5264 2752
rect 4944 2294 5264 2688
rect 944 2016 1264 2058
rect 4944 2058 4986 2294
rect 5222 2058 5264 2294
rect 5604 15264 5924 15824
rect 5604 15200 5612 15264
rect 5676 15200 5692 15264
rect 5756 15200 5772 15264
rect 5836 15200 5852 15264
rect 5916 15200 5924 15264
rect 5604 14954 5924 15200
rect 5604 14718 5646 14954
rect 5882 14718 5924 14954
rect 5604 14176 5924 14718
rect 5604 14112 5612 14176
rect 5676 14112 5692 14176
rect 5756 14112 5772 14176
rect 5836 14112 5852 14176
rect 5916 14112 5924 14176
rect 5604 13088 5924 14112
rect 5604 13024 5612 13088
rect 5676 13024 5692 13088
rect 5756 13024 5772 13088
rect 5836 13024 5852 13088
rect 5916 13024 5924 13088
rect 5604 12000 5924 13024
rect 5604 11936 5612 12000
rect 5676 11936 5692 12000
rect 5756 11936 5772 12000
rect 5836 11936 5852 12000
rect 5916 11936 5924 12000
rect 5604 10954 5924 11936
rect 5604 10912 5646 10954
rect 5882 10912 5924 10954
rect 5604 10848 5612 10912
rect 5916 10848 5924 10912
rect 5604 10718 5646 10848
rect 5882 10718 5924 10848
rect 5604 9824 5924 10718
rect 5604 9760 5612 9824
rect 5676 9760 5692 9824
rect 5756 9760 5772 9824
rect 5836 9760 5852 9824
rect 5916 9760 5924 9824
rect 5604 8736 5924 9760
rect 5604 8672 5612 8736
rect 5676 8672 5692 8736
rect 5756 8672 5772 8736
rect 5836 8672 5852 8736
rect 5916 8672 5924 8736
rect 5604 7648 5924 8672
rect 5604 7584 5612 7648
rect 5676 7584 5692 7648
rect 5756 7584 5772 7648
rect 5836 7584 5852 7648
rect 5916 7584 5924 7648
rect 5604 6954 5924 7584
rect 5604 6718 5646 6954
rect 5882 6718 5924 6954
rect 5604 6560 5924 6718
rect 5604 6496 5612 6560
rect 5676 6496 5692 6560
rect 5756 6496 5772 6560
rect 5836 6496 5852 6560
rect 5916 6496 5924 6560
rect 5604 5472 5924 6496
rect 5604 5408 5612 5472
rect 5676 5408 5692 5472
rect 5756 5408 5772 5472
rect 5836 5408 5852 5472
rect 5916 5408 5924 5472
rect 5604 4384 5924 5408
rect 5604 4320 5612 4384
rect 5676 4320 5692 4384
rect 5756 4320 5772 4384
rect 5836 4320 5852 4384
rect 5916 4320 5924 4384
rect 5604 3296 5924 4320
rect 5604 3232 5612 3296
rect 5676 3232 5692 3296
rect 5756 3232 5772 3296
rect 5836 3232 5852 3296
rect 5916 3232 5924 3296
rect 5604 2954 5924 3232
rect 5604 2718 5646 2954
rect 5882 2718 5924 2954
rect 5604 2208 5924 2718
rect 5604 2144 5612 2208
rect 5676 2144 5692 2208
rect 5756 2144 5772 2208
rect 5836 2144 5852 2208
rect 5916 2144 5924 2208
rect 5604 2128 5924 2144
rect 8944 15808 9264 15824
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 14720 9264 15744
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 14294 9264 14656
rect 8944 14058 8986 14294
rect 9222 14058 9264 14294
rect 8944 13632 9264 14058
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 12544 9264 13568
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 11456 9264 12480
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 10368 9264 11392
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 10294 9264 10304
rect 8944 10058 8986 10294
rect 9222 10058 9264 10294
rect 8944 9280 9264 10058
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 8192 9264 9216
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 7104 9264 8128
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 6294 9264 7040
rect 8944 6058 8986 6294
rect 9222 6058 9264 6294
rect 8944 6016 9264 6058
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 4928 9264 5952
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 3840 9264 4864
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 2752 9264 3776
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2294 9264 2688
rect 4944 2016 5264 2058
rect 8944 2058 8986 2294
rect 9222 2058 9264 2294
rect 9604 15264 9924 15824
rect 9604 15200 9612 15264
rect 9676 15200 9692 15264
rect 9756 15200 9772 15264
rect 9836 15200 9852 15264
rect 9916 15200 9924 15264
rect 9604 14954 9924 15200
rect 9604 14718 9646 14954
rect 9882 14718 9924 14954
rect 9604 14176 9924 14718
rect 9604 14112 9612 14176
rect 9676 14112 9692 14176
rect 9756 14112 9772 14176
rect 9836 14112 9852 14176
rect 9916 14112 9924 14176
rect 9604 13088 9924 14112
rect 9604 13024 9612 13088
rect 9676 13024 9692 13088
rect 9756 13024 9772 13088
rect 9836 13024 9852 13088
rect 9916 13024 9924 13088
rect 9604 12000 9924 13024
rect 9604 11936 9612 12000
rect 9676 11936 9692 12000
rect 9756 11936 9772 12000
rect 9836 11936 9852 12000
rect 9916 11936 9924 12000
rect 9604 10954 9924 11936
rect 9604 10912 9646 10954
rect 9882 10912 9924 10954
rect 9604 10848 9612 10912
rect 9916 10848 9924 10912
rect 9604 10718 9646 10848
rect 9882 10718 9924 10848
rect 9604 9824 9924 10718
rect 9604 9760 9612 9824
rect 9676 9760 9692 9824
rect 9756 9760 9772 9824
rect 9836 9760 9852 9824
rect 9916 9760 9924 9824
rect 9604 8736 9924 9760
rect 9604 8672 9612 8736
rect 9676 8672 9692 8736
rect 9756 8672 9772 8736
rect 9836 8672 9852 8736
rect 9916 8672 9924 8736
rect 9604 7648 9924 8672
rect 9604 7584 9612 7648
rect 9676 7584 9692 7648
rect 9756 7584 9772 7648
rect 9836 7584 9852 7648
rect 9916 7584 9924 7648
rect 9604 6954 9924 7584
rect 9604 6718 9646 6954
rect 9882 6718 9924 6954
rect 9604 6560 9924 6718
rect 9604 6496 9612 6560
rect 9676 6496 9692 6560
rect 9756 6496 9772 6560
rect 9836 6496 9852 6560
rect 9916 6496 9924 6560
rect 9604 5472 9924 6496
rect 9604 5408 9612 5472
rect 9676 5408 9692 5472
rect 9756 5408 9772 5472
rect 9836 5408 9852 5472
rect 9916 5408 9924 5472
rect 9604 4384 9924 5408
rect 9604 4320 9612 4384
rect 9676 4320 9692 4384
rect 9756 4320 9772 4384
rect 9836 4320 9852 4384
rect 9916 4320 9924 4384
rect 9604 3296 9924 4320
rect 9604 3232 9612 3296
rect 9676 3232 9692 3296
rect 9756 3232 9772 3296
rect 9836 3232 9852 3296
rect 9916 3232 9924 3296
rect 9604 2954 9924 3232
rect 9604 2718 9646 2954
rect 9882 2718 9924 2954
rect 9604 2208 9924 2718
rect 9604 2144 9612 2208
rect 9676 2144 9692 2208
rect 9756 2144 9772 2208
rect 9836 2144 9852 2208
rect 9916 2144 9924 2208
rect 9604 2128 9924 2144
rect 12944 15808 13264 15824
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 14294 13264 14656
rect 12944 14058 12986 14294
rect 13222 14058 13264 14294
rect 12944 13632 13264 14058
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 10294 13264 10304
rect 12944 10058 12986 10294
rect 13222 10058 13264 10294
rect 12944 9280 13264 10058
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6294 13264 7040
rect 12944 6058 12986 6294
rect 13222 6058 13264 6294
rect 12944 6016 13264 6058
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2294 13264 2688
rect 8944 2016 9264 2058
rect 12944 2058 12986 2294
rect 13222 2058 13264 2294
rect 13604 15264 13924 15824
rect 13604 15200 13612 15264
rect 13676 15200 13692 15264
rect 13756 15200 13772 15264
rect 13836 15200 13852 15264
rect 13916 15200 13924 15264
rect 13604 14954 13924 15200
rect 13604 14718 13646 14954
rect 13882 14718 13924 14954
rect 13604 14176 13924 14718
rect 13604 14112 13612 14176
rect 13676 14112 13692 14176
rect 13756 14112 13772 14176
rect 13836 14112 13852 14176
rect 13916 14112 13924 14176
rect 13604 13088 13924 14112
rect 13604 13024 13612 13088
rect 13676 13024 13692 13088
rect 13756 13024 13772 13088
rect 13836 13024 13852 13088
rect 13916 13024 13924 13088
rect 13604 12000 13924 13024
rect 13604 11936 13612 12000
rect 13676 11936 13692 12000
rect 13756 11936 13772 12000
rect 13836 11936 13852 12000
rect 13916 11936 13924 12000
rect 13604 10954 13924 11936
rect 13604 10912 13646 10954
rect 13882 10912 13924 10954
rect 13604 10848 13612 10912
rect 13916 10848 13924 10912
rect 13604 10718 13646 10848
rect 13882 10718 13924 10848
rect 13604 9824 13924 10718
rect 13604 9760 13612 9824
rect 13676 9760 13692 9824
rect 13756 9760 13772 9824
rect 13836 9760 13852 9824
rect 13916 9760 13924 9824
rect 13604 8736 13924 9760
rect 13604 8672 13612 8736
rect 13676 8672 13692 8736
rect 13756 8672 13772 8736
rect 13836 8672 13852 8736
rect 13916 8672 13924 8736
rect 13604 7648 13924 8672
rect 13604 7584 13612 7648
rect 13676 7584 13692 7648
rect 13756 7584 13772 7648
rect 13836 7584 13852 7648
rect 13916 7584 13924 7648
rect 13604 6954 13924 7584
rect 13604 6718 13646 6954
rect 13882 6718 13924 6954
rect 13604 6560 13924 6718
rect 13604 6496 13612 6560
rect 13676 6496 13692 6560
rect 13756 6496 13772 6560
rect 13836 6496 13852 6560
rect 13916 6496 13924 6560
rect 13604 5472 13924 6496
rect 13604 5408 13612 5472
rect 13676 5408 13692 5472
rect 13756 5408 13772 5472
rect 13836 5408 13852 5472
rect 13916 5408 13924 5472
rect 13604 4384 13924 5408
rect 13604 4320 13612 4384
rect 13676 4320 13692 4384
rect 13756 4320 13772 4384
rect 13836 4320 13852 4384
rect 13916 4320 13924 4384
rect 13604 3296 13924 4320
rect 13604 3232 13612 3296
rect 13676 3232 13692 3296
rect 13756 3232 13772 3296
rect 13836 3232 13852 3296
rect 13916 3232 13924 3296
rect 13604 2954 13924 3232
rect 13604 2718 13646 2954
rect 13882 2718 13924 2954
rect 13604 2208 13924 2718
rect 13604 2144 13612 2208
rect 13676 2144 13692 2208
rect 13756 2144 13772 2208
rect 13836 2144 13852 2208
rect 13916 2144 13924 2208
rect 13604 2128 13924 2144
rect 12944 2016 13264 2058
<< via4 >>
rect 986 14058 1222 14294
rect 986 10058 1222 10294
rect 986 6058 1222 6294
rect 986 2058 1222 2294
rect 1646 14718 1882 14954
rect 1646 10912 1882 10954
rect 1646 10848 1676 10912
rect 1676 10848 1692 10912
rect 1692 10848 1756 10912
rect 1756 10848 1772 10912
rect 1772 10848 1836 10912
rect 1836 10848 1852 10912
rect 1852 10848 1882 10912
rect 1646 10718 1882 10848
rect 1646 6718 1882 6954
rect 1646 2718 1882 2954
rect 4986 14058 5222 14294
rect 4986 10058 5222 10294
rect 4986 6058 5222 6294
rect 4986 2058 5222 2294
rect 5646 14718 5882 14954
rect 5646 10912 5882 10954
rect 5646 10848 5676 10912
rect 5676 10848 5692 10912
rect 5692 10848 5756 10912
rect 5756 10848 5772 10912
rect 5772 10848 5836 10912
rect 5836 10848 5852 10912
rect 5852 10848 5882 10912
rect 5646 10718 5882 10848
rect 5646 6718 5882 6954
rect 5646 2718 5882 2954
rect 8986 14058 9222 14294
rect 8986 10058 9222 10294
rect 8986 6058 9222 6294
rect 8986 2058 9222 2294
rect 9646 14718 9882 14954
rect 9646 10912 9882 10954
rect 9646 10848 9676 10912
rect 9676 10848 9692 10912
rect 9692 10848 9756 10912
rect 9756 10848 9772 10912
rect 9772 10848 9836 10912
rect 9836 10848 9852 10912
rect 9852 10848 9882 10912
rect 9646 10718 9882 10848
rect 9646 6718 9882 6954
rect 9646 2718 9882 2954
rect 12986 14058 13222 14294
rect 12986 10058 13222 10294
rect 12986 6058 13222 6294
rect 12986 2058 13222 2294
rect 13646 14718 13882 14954
rect 13646 10912 13882 10954
rect 13646 10848 13676 10912
rect 13676 10848 13692 10912
rect 13692 10848 13756 10912
rect 13756 10848 13772 10912
rect 13772 10848 13836 10912
rect 13836 10848 13852 10912
rect 13852 10848 13882 10912
rect 13646 10718 13882 10848
rect 13646 6718 13882 6954
rect 13646 2718 13882 2954
<< metal5 >>
rect 1056 14954 16884 14996
rect 1056 14718 1646 14954
rect 1882 14718 5646 14954
rect 5882 14718 9646 14954
rect 9882 14718 13646 14954
rect 13882 14718 16884 14954
rect 1056 14676 16884 14718
rect 944 14294 16884 14336
rect 944 14058 986 14294
rect 1222 14058 4986 14294
rect 5222 14058 8986 14294
rect 9222 14058 12986 14294
rect 13222 14058 16884 14294
rect 944 14016 16884 14058
rect 1056 10954 16884 10996
rect 1056 10718 1646 10954
rect 1882 10718 5646 10954
rect 5882 10718 9646 10954
rect 9882 10718 13646 10954
rect 13882 10718 16884 10954
rect 1056 10676 16884 10718
rect 944 10294 16884 10336
rect 944 10058 986 10294
rect 1222 10058 4986 10294
rect 5222 10058 8986 10294
rect 9222 10058 12986 10294
rect 13222 10058 16884 10294
rect 944 10016 16884 10058
rect 1056 6954 16884 6996
rect 1056 6718 1646 6954
rect 1882 6718 5646 6954
rect 5882 6718 9646 6954
rect 9882 6718 13646 6954
rect 13882 6718 16884 6954
rect 1056 6676 16884 6718
rect 944 6294 16884 6336
rect 944 6058 986 6294
rect 1222 6058 4986 6294
rect 5222 6058 8986 6294
rect 9222 6058 12986 6294
rect 13222 6058 16884 6294
rect 944 6016 16884 6058
rect 1056 2954 16884 2996
rect 1056 2718 1646 2954
rect 1882 2718 5646 2954
rect 5882 2718 9646 2954
rect 9882 2718 13646 2954
rect 13882 2718 16884 2954
rect 1056 2676 16884 2718
rect 944 2294 16884 2336
rect 944 2058 986 2294
rect 1222 2058 4986 2294
rect 5222 2058 8986 2294
rect 9222 2058 12986 2294
rect 13222 2058 16884 2294
rect 944 2016 16884 2058
use sky130_fd_sc_hd__and4b_1  _142_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _143_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _144_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5060 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 7176 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 7268 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 7544 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _148_
timestamp 1693170804
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 10396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _150_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 5796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 6716 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _153_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 6256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 5980 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _156_
timestamp 1693170804
transform 1 0 10856 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _157_
timestamp 1693170804
transform 1 0 14076 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _159_
timestamp 1693170804
transform 1 0 15916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _160_
timestamp 1693170804
transform 1 0 3404 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _161_
timestamp 1693170804
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1693170804
transform 1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _163_
timestamp 1693170804
transform 1 0 14536 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _164_
timestamp 1693170804
transform 1 0 14904 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1693170804
transform 1 0 15732 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _166_
timestamp 1693170804
transform -1 0 3404 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _167_
timestamp 1693170804
transform -1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1693170804
transform 1 0 2300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _169_
timestamp 1693170804
transform 1 0 3036 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _170_
timestamp 1693170804
transform -1 0 3220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1693170804
transform -1 0 2300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _172_
timestamp 1693170804
transform 1 0 14720 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _173_
timestamp 1693170804
transform 1 0 15088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1693170804
transform -1 0 14996 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _175_
timestamp 1693170804
transform -1 0 12972 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _176_
timestamp 1693170804
transform -1 0 12420 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1693170804
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _178_
timestamp 1693170804
transform -1 0 16284 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _179_
timestamp 1693170804
transform 1 0 15732 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1693170804
transform 1 0 16008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _181_
timestamp 1693170804
transform 1 0 5796 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _182_
timestamp 1693170804
transform -1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1693170804
transform -1 0 6256 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _184_
timestamp 1693170804
transform 1 0 7728 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _185_
timestamp 1693170804
transform 1 0 8924 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1693170804
transform -1 0 8280 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _187_
timestamp 1693170804
transform 1 0 10948 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _188_
timestamp 1693170804
transform -1 0 11408 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1693170804
transform 1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _190_
timestamp 1693170804
transform 1 0 11960 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _191_
timestamp 1693170804
transform -1 0 12420 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1693170804
transform -1 0 2760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _193_
timestamp 1693170804
transform 1 0 9660 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _194_
timestamp 1693170804
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _195_
timestamp 1693170804
transform -1 0 8648 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8924 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _197_
timestamp 1693170804
transform -1 0 9844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5704 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1693170804
transform -1 0 6440 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4876 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _202_
timestamp 1693170804
transform -1 0 4968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _203_
timestamp 1693170804
transform -1 0 4968 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _204_
timestamp 1693170804
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1693170804
transform 1 0 2208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 5336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _207_
timestamp 1693170804
transform -1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _209_
timestamp 1693170804
transform -1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 2300 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _211_
timestamp 1693170804
transform 1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _212_
timestamp 1693170804
transform 1 0 2208 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _213_
timestamp 1693170804
transform -1 0 3680 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1693170804
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 6348 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__o21ai_4  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9936 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 11684 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 3404 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 11040 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _220_
timestamp 1693170804
transform -1 0 13340 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _221_
timestamp 1693170804
transform 1 0 13340 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _222_
timestamp 1693170804
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _223_
timestamp 1693170804
transform 1 0 2668 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _224_
timestamp 1693170804
transform -1 0 2484 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1693170804
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _226_
timestamp 1693170804
transform 1 0 13432 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _227_
timestamp 1693170804
transform 1 0 12972 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp 1693170804
transform -1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _229_
timestamp 1693170804
transform 1 0 2300 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _230_
timestamp 1693170804
transform -1 0 2392 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1693170804
transform 1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _232_
timestamp 1693170804
transform 1 0 2392 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _233_
timestamp 1693170804
transform -1 0 2392 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1693170804
transform 1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _235_
timestamp 1693170804
transform 1 0 13892 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _236_
timestamp 1693170804
transform -1 0 13984 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 1693170804
transform -1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _238_
timestamp 1693170804
transform 1 0 11868 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _239_
timestamp 1693170804
transform 1 0 11500 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1693170804
transform 1 0 11960 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _241_
timestamp 1693170804
transform 1 0 15180 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _242_
timestamp 1693170804
transform 1 0 14812 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1693170804
transform 1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _244_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _246_
timestamp 1693170804
transform 1 0 11868 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _247_
timestamp 1693170804
transform -1 0 14628 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _248_
timestamp 1693170804
transform -1 0 12788 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _249_
timestamp 1693170804
transform -1 0 11776 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _250_
timestamp 1693170804
transform -1 0 11224 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _251_
timestamp 1693170804
transform -1 0 11224 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _252_
timestamp 1693170804
transform 1 0 8372 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _253_
timestamp 1693170804
transform -1 0 10764 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _254_
timestamp 1693170804
transform -1 0 10672 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _255_
timestamp 1693170804
transform 1 0 9660 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _256_
timestamp 1693170804
transform 1 0 12328 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _257_
timestamp 1693170804
transform -1 0 13340 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _258_
timestamp 1693170804
transform -1 0 13248 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _259_
timestamp 1693170804
transform 1 0 11776 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _260_
timestamp 1693170804
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_2  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _262_
timestamp 1693170804
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _263_
timestamp 1693170804
transform -1 0 8096 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _264_
timestamp 1693170804
transform 1 0 6348 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _265_
timestamp 1693170804
transform 1 0 8096 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _266_
timestamp 1693170804
transform 1 0 8556 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _267_
timestamp 1693170804
transform -1 0 9660 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _268_
timestamp 1693170804
transform -1 0 8832 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _269_
timestamp 1693170804
transform -1 0 11408 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _270_
timestamp 1693170804
transform -1 0 9936 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _271_
timestamp 1693170804
transform 1 0 6440 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _273_
timestamp 1693170804
transform 1 0 5244 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _274_
timestamp 1693170804
transform -1 0 6072 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _275_
timestamp 1693170804
transform -1 0 6072 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1693170804
transform 1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _277_
timestamp 1693170804
transform 1 0 7176 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _278_
timestamp 1693170804
transform 1 0 6808 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp 1693170804
transform 1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _280_
timestamp 1693170804
transform 1 0 10580 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _281_
timestamp 1693170804
transform 1 0 10488 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1693170804
transform -1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _283_
timestamp 1693170804
transform -1 0 11408 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _284_
timestamp 1693170804
transform 1 0 11500 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp 1693170804
transform -1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _286_
timestamp 1693170804
transform 1 0 6624 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _287_
timestamp 1693170804
transform 1 0 6992 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1693170804
transform -1 0 6992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _290_
timestamp 1693170804
transform -1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8464 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4324 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _293_
timestamp 1693170804
transform 1 0 3864 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1693170804
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _295_
timestamp 1693170804
transform 1 0 3680 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _296_
timestamp 1693170804
transform 1 0 5336 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _297_
timestamp 1693170804
transform 1 0 4140 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4140 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4416 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _300_
timestamp 1693170804
transform -1 0 5336 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _301_
timestamp 1693170804
transform 1 0 6992 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _302_
timestamp 1693170804
transform 1 0 6532 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 1693170804
transform 1 0 7176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 8372 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _305_
timestamp 1693170804
transform 1 0 5152 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1693170804
transform 1 0 7360 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _307_
timestamp 1693170804
transform -1 0 7728 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _308_
timestamp 1693170804
transform 1 0 5612 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _309_
timestamp 1693170804
transform -1 0 7452 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _310_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4968 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _311__47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4140 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _312_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 11132 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _313_
timestamp 1693170804
transform 1 0 6348 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 6716 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _315_
timestamp 1693170804
transform 1 0 7268 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8924 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _317_
timestamp 1693170804
transform 1 0 1748 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _318_
timestamp 1693170804
transform 1 0 1380 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _319_
timestamp 1693170804
transform 1 0 1380 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _320_
timestamp 1693170804
transform 1 0 1472 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _321_
timestamp 1693170804
transform -1 0 14168 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 1693170804
transform 1 0 1564 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _323_
timestamp 1693170804
transform 1 0 14076 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _324_
timestamp 1693170804
transform 1 0 1380 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _325_
timestamp 1693170804
transform 1 0 1380 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1693170804
transform 1 0 14076 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _327_
timestamp 1693170804
transform 1 0 11132 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _328_
timestamp 1693170804
transform 1 0 14076 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _329_
timestamp 1693170804
transform 1 0 3588 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _330_
timestamp 1693170804
transform -1 0 13984 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _331_
timestamp 1693170804
transform 1 0 11500 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _332_
timestamp 1693170804
transform 1 0 11224 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _333_
timestamp 1693170804
transform -1 0 10948 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _334_
timestamp 1693170804
transform -1 0 10304 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _335_
timestamp 1693170804
transform 1 0 13064 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _336_
timestamp 1693170804
transform 1 0 10948 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _337_
timestamp 1693170804
transform 1 0 13340 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _338_
timestamp 1693170804
transform 1 0 3864 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _339_
timestamp 1693170804
transform -1 0 9936 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _340_
timestamp 1693170804
transform 1 0 9476 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _341_
timestamp 1693170804
transform 1 0 9016 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _342_
timestamp 1693170804
transform 1 0 5796 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _343_
timestamp 1693170804
transform 1 0 3772 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _344_
timestamp 1693170804
transform 1 0 6348 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _345_
timestamp 1693170804
transform -1 0 13340 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _346_
timestamp 1693170804
transform -1 0 13340 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _347_
timestamp 1693170804
transform 1 0 6992 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _348_
timestamp 1693170804
transform 1 0 8648 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _349_
timestamp 1693170804
transform 1 0 3220 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _350_
timestamp 1693170804
transform 1 0 2484 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _351_
timestamp 1693170804
transform 1 0 5152 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _352_
timestamp 1693170804
transform 1 0 4784 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 9660 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1693170804
transform -1 0 4600 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1693170804
transform -1 0 4600 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1693170804
transform 1 0 10856 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1693170804
transform 1 0 11500 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1693170804
transform -1 0 2300 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 1693170804
transform 1 0 2760 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 1693170804
transform 1 0 11132 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1693170804
transform -1 0 10488 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp 1693170804
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 2300 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_35
timestamp 1693170804
transform 1 0 4324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_42
timestamp 1693170804
transform 1 0 4968 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_77
timestamp 1693170804
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1693170804
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1693170804
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_100
timestamp 1693170804
transform 1 0 10304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_121 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_133
timestamp 1693170804
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1693170804
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_141
timestamp 1693170804
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_147
timestamp 1693170804
transform 1 0 14628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_154
timestamp 1693170804
transform 1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_12
timestamp 1693170804
transform 1 0 2208 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_24
timestamp 1693170804
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_28
timestamp 1693170804
transform 1 0 3680 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1693170804
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 1693170804
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_61
timestamp 1693170804
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_70
timestamp 1693170804
transform 1 0 7544 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_133
timestamp 1693170804
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_145
timestamp 1693170804
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_149
timestamp 1693170804
transform 1 0 14812 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_153
timestamp 1693170804
transform 1 0 15180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_157
timestamp 1693170804
transform 1 0 15548 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_161
timestamp 1693170804
transform 1 0 15916 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_9
timestamp 1693170804
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_21
timestamp 1693170804
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1693170804
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_32
timestamp 1693170804
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_39
timestamp 1693170804
transform 1 0 4692 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_59
timestamp 1693170804
transform 1 0 6532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_65
timestamp 1693170804
transform 1 0 7084 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1693170804
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1693170804
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_96
timestamp 1693170804
transform 1 0 9936 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_102
timestamp 1693170804
transform 1 0 10488 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_109
timestamp 1693170804
transform 1 0 11132 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_114
timestamp 1693170804
transform 1 0 11592 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_126
timestamp 1693170804
transform 1 0 12696 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_138
timestamp 1693170804
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_146
timestamp 1693170804
transform 1 0 14536 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_158
timestamp 1693170804
transform 1 0 15640 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_164
timestamp 1693170804
transform 1 0 16192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_3
timestamp 1693170804
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_50
timestamp 1693170804
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_64
timestamp 1693170804
transform 1 0 6992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_88
timestamp 1693170804
transform 1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1693170804
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_116
timestamp 1693170804
transform 1 0 11776 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_142
timestamp 1693170804
transform 1 0 14168 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_154
timestamp 1693170804
transform 1 0 15272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 1693170804
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_3
timestamp 1693170804
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_15
timestamp 1693170804
transform 1 0 2484 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1693170804
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_41
timestamp 1693170804
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_49
timestamp 1693170804
transform 1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_76
timestamp 1693170804
transform 1 0 8096 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_95
timestamp 1693170804
transform 1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_112
timestamp 1693170804
transform 1 0 11408 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_123
timestamp 1693170804
transform 1 0 12420 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1693170804
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_144
timestamp 1693170804
transform 1 0 14352 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_156
timestamp 1693170804
transform 1 0 15456 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_6
timestamp 1693170804
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_24
timestamp 1693170804
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_47
timestamp 1693170804
transform 1 0 5428 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1693170804
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1693170804
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_65
timestamp 1693170804
transform 1 0 7084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_96
timestamp 1693170804
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_133
timestamp 1693170804
transform 1 0 13340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_145
timestamp 1693170804
transform 1 0 14444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_157
timestamp 1693170804
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 1693170804
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1693170804
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_24
timestamp 1693170804
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_45
timestamp 1693170804
transform 1 0 5244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_66
timestamp 1693170804
transform 1 0 7176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_75
timestamp 1693170804
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1693170804
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 1693170804
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_126
timestamp 1693170804
transform 1 0 12696 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1693170804
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1693170804
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_153
timestamp 1693170804
transform 1 0 15180 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_161
timestamp 1693170804
transform 1 0 15916 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_41
timestamp 1693170804
transform 1 0 4876 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_47
timestamp 1693170804
transform 1 0 5428 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1693170804
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 1693170804
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_82
timestamp 1693170804
transform 1 0 8648 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_94
timestamp 1693170804
transform 1 0 9752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_101
timestamp 1693170804
transform 1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 1693170804
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_123
timestamp 1693170804
transform 1 0 12420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_135
timestamp 1693170804
transform 1 0 13524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_147
timestamp 1693170804
transform 1 0 14628 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_159
timestamp 1693170804
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1693170804
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_37
timestamp 1693170804
transform 1 0 4508 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_112
timestamp 1693170804
transform 1 0 11408 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_147
timestamp 1693170804
transform 1 0 14628 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_159
timestamp 1693170804
transform 1 0 15732 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_167
timestamp 1693170804
transform 1 0 16468 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_3
timestamp 1693170804
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_42
timestamp 1693170804
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1693170804
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57
timestamp 1693170804
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_65
timestamp 1693170804
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_72
timestamp 1693170804
transform 1 0 7728 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_93
timestamp 1693170804
transform 1 0 9660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1693170804
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1693170804
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_23
timestamp 1693170804
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1693170804
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_58
timestamp 1693170804
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1693170804
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_85
timestamp 1693170804
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_109
timestamp 1693170804
transform 1 0 11132 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_116
timestamp 1693170804
transform 1 0 11776 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1693170804
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_157
timestamp 1693170804
transform 1 0 15548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_161
timestamp 1693170804
transform 1 0 15916 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1693170804
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_15
timestamp 1693170804
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_46
timestamp 1693170804
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1693170804
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_68
timestamp 1693170804
transform 1 0 7360 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1693170804
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1693170804
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1693170804
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_165
timestamp 1693170804
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_9
timestamp 1693170804
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1693170804
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1693170804
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_38
timestamp 1693170804
transform 1 0 4600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_51
timestamp 1693170804
transform 1 0 5796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_132
timestamp 1693170804
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_144
timestamp 1693170804
transform 1 0 14352 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_156
timestamp 1693170804
transform 1 0 15456 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 1693170804
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_28
timestamp 1693170804
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_32
timestamp 1693170804
transform 1 0 4048 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1693170804
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_66
timestamp 1693170804
transform 1 0 7176 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_78
timestamp 1693170804
transform 1 0 8280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1693170804
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1693170804
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_117
timestamp 1693170804
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_126
timestamp 1693170804
transform 1 0 12696 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1693170804
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1693170804
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_9
timestamp 1693170804
transform 1 0 1932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_21
timestamp 1693170804
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1693170804
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 1693170804
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_37
timestamp 1693170804
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1693170804
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_53
timestamp 1693170804
transform 1 0 5980 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_59
timestamp 1693170804
transform 1 0 6532 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_73
timestamp 1693170804
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1693170804
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_98
timestamp 1693170804
transform 1 0 10120 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_130
timestamp 1693170804
transform 1 0 13064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1693170804
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_141
timestamp 1693170804
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_145
timestamp 1693170804
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_151
timestamp 1693170804
transform 1 0 14996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_163
timestamp 1693170804
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_167
timestamp 1693170804
transform 1 0 16468 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_23
timestamp 1693170804
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_47
timestamp 1693170804
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1693170804
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_57
timestamp 1693170804
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_92
timestamp 1693170804
transform 1 0 9568 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_104
timestamp 1693170804
transform 1 0 10672 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1693170804
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_113
timestamp 1693170804
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_127
timestamp 1693170804
transform 1 0 12788 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_153
timestamp 1693170804
transform 1 0 15180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1693170804
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_3
timestamp 1693170804
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1693170804
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_29
timestamp 1693170804
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_39
timestamp 1693170804
transform 1 0 4692 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_71
timestamp 1693170804
transform 1 0 7636 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_85
timestamp 1693170804
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_97
timestamp 1693170804
transform 1 0 10028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_105
timestamp 1693170804
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_135
timestamp 1693170804
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1693170804
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_149
timestamp 1693170804
transform 1 0 14812 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_157
timestamp 1693170804
transform 1 0 15548 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1693170804
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_15
timestamp 1693170804
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_44
timestamp 1693170804
transform 1 0 5152 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_48
timestamp 1693170804
transform 1 0 5520 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1693170804
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_61
timestamp 1693170804
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_69
timestamp 1693170804
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_77
timestamp 1693170804
transform 1 0 8188 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_100
timestamp 1693170804
transform 1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_123
timestamp 1693170804
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_133
timestamp 1693170804
transform 1 0 13340 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_146
timestamp 1693170804
transform 1 0 14536 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_153
timestamp 1693170804
transform 1 0 15180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 1693170804
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1693170804
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 1693170804
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_11
timestamp 1693170804
transform 1 0 2116 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_25
timestamp 1693170804
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_32
timestamp 1693170804
transform 1 0 4048 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1693170804
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_77
timestamp 1693170804
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1693170804
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_93
timestamp 1693170804
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_102
timestamp 1693170804
transform 1 0 10488 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_114
timestamp 1693170804
transform 1 0 11592 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_129
timestamp 1693170804
transform 1 0 12972 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_161
timestamp 1693170804
transform 1 0 15916 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_167
timestamp 1693170804
transform 1 0 16468 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_14
timestamp 1693170804
transform 1 0 2392 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_43
timestamp 1693170804
transform 1 0 5060 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1693170804
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1693170804
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_65
timestamp 1693170804
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_69
timestamp 1693170804
transform 1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_77
timestamp 1693170804
transform 1 0 8188 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_82
timestamp 1693170804
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_86
timestamp 1693170804
transform 1 0 9016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_107
timestamp 1693170804
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1693170804
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_121
timestamp 1693170804
transform 1 0 12236 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_133
timestamp 1693170804
transform 1 0 13340 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_145
timestamp 1693170804
transform 1 0 14444 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_151
timestamp 1693170804
transform 1 0 14996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_155
timestamp 1693170804
transform 1 0 15364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1693170804
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_23
timestamp 1693170804
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1693170804
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_29
timestamp 1693170804
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_47
timestamp 1693170804
transform 1 0 5428 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_79
timestamp 1693170804
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1693170804
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_95
timestamp 1693170804
transform 1 0 9844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_107
timestamp 1693170804
transform 1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_129
timestamp 1693170804
transform 1 0 12972 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1693170804
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1693170804
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_153
timestamp 1693170804
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_161
timestamp 1693170804
transform 1 0 15916 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_9
timestamp 1693170804
transform 1 0 1932 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_17
timestamp 1693170804
transform 1 0 2668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_25
timestamp 1693170804
transform 1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1693170804
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1693170804
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_57
timestamp 1693170804
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_63
timestamp 1693170804
transform 1 0 6900 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_67
timestamp 1693170804
transform 1 0 7268 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_79
timestamp 1693170804
transform 1 0 8372 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_91
timestamp 1693170804
transform 1 0 9476 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_103
timestamp 1693170804
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1693170804
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1693170804
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1693170804
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1693170804
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1693170804
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1693170804
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1693170804
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1693170804
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1693170804
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1693170804
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1693170804
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1693170804
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1693170804
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1693170804
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1693170804
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1693170804
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1693170804
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1693170804
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1693170804
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1693170804
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1693170804
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1693170804
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1693170804
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_153
timestamp 1693170804
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_161
timestamp 1693170804
transform 1 0 15916 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_9
timestamp 1693170804
transform 1 0 1932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_16
timestamp 1693170804
transform 1 0 2576 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_23
timestamp 1693170804
transform 1 0 3220 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_35
timestamp 1693170804
transform 1 0 4324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_47
timestamp 1693170804
transform 1 0 5428 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1693170804
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_69
timestamp 1693170804
transform 1 0 7452 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_78
timestamp 1693170804
transform 1 0 8280 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_90
timestamp 1693170804
transform 1 0 9384 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_102
timestamp 1693170804
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1693170804
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1693170804
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1693170804
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_137
timestamp 1693170804
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_145
timestamp 1693170804
transform 1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_151
timestamp 1693170804
transform 1 0 14996 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_159
timestamp 1693170804
transform 1 0 15732 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_15
timestamp 1693170804
transform 1 0 2484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_23
timestamp 1693170804
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1693170804
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1693170804
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_37
timestamp 1693170804
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1693170804
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_53
timestamp 1693170804
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_63
timestamp 1693170804
transform 1 0 6900 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_71
timestamp 1693170804
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 1693170804
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1693170804
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 1693170804
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_90
timestamp 1693170804
transform 1 0 9384 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_102
timestamp 1693170804
transform 1 0 10488 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_110
timestamp 1693170804
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_119
timestamp 1693170804
transform 1 0 12052 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_127
timestamp 1693170804
transform 1 0 12788 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_135
timestamp 1693170804
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1693170804
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_141
timestamp 1693170804
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_149
timestamp 1693170804
transform 1 0 14812 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_155
timestamp 1693170804
transform 1 0 15364 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 11224 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1693170804
transform 1 0 6440 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1693170804
transform -1 0 9936 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1693170804
transform -1 0 3680 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1693170804
transform -1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1693170804
transform -1 0 6440 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1693170804
transform -1 0 13524 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1693170804
transform -1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1693170804
transform -1 0 12696 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1693170804
transform -1 0 10948 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1693170804
transform -1 0 8096 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1693170804
transform -1 0 14812 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1693170804
transform 1 0 9292 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1693170804
transform 1 0 9752 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1693170804
transform -1 0 10856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1693170804
transform -1 0 8648 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1693170804
transform -1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1693170804
transform -1 0 14076 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1693170804
transform -1 0 9568 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1693170804
transform -1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1693170804
transform -1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1693170804
transform 1 0 6624 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1693170804
transform -1 0 5428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1693170804
transform -1 0 7084 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1693170804
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1693170804
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1693170804
transform 1 0 4600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1693170804
transform -1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1693170804
transform -1 0 9384 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1693170804
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 1693170804
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 1693170804
transform 1 0 16008 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1693170804
transform -1 0 2484 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 1693170804
transform -1 0 1932 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1693170804
transform -1 0 14812 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 1693170804
transform 1 0 9752 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1693170804
transform 1 0 16008 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1693170804
transform 1 0 15640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1693170804
transform -1 0 3680 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1693170804
transform -1 0 1932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1693170804
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1693170804
transform 1 0 11500 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1693170804
transform 1 0 16008 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1693170804
transform -1 0 1932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1693170804
transform 1 0 16008 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1693170804
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1693170804
transform -1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1693170804
transform 1 0 16008 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 1693170804
transform -1 0 3220 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1693170804
transform -1 0 2300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1693170804
transform -1 0 15272 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1693170804
transform 1 0 12972 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1693170804
transform 1 0 16008 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1693170804
transform -1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1693170804
transform -1 0 6256 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1693170804
transform 1 0 16008 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1693170804
transform -1 0 8832 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1693170804
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1693170804
transform 1 0 15456 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1693170804
transform 1 0 6348 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1693170804
transform -1 0 8372 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1693170804
transform 1 0 11684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1693170804
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1693170804
transform -1 0 1932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1693170804
transform 1 0 16008 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_25
timestamp 1693170804
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1693170804
transform -1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_26
timestamp 1693170804
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1693170804
transform -1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_27
timestamp 1693170804
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1693170804
transform -1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_28
timestamp 1693170804
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1693170804
transform -1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_29
timestamp 1693170804
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1693170804
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_30
timestamp 1693170804
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1693170804
transform -1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_31
timestamp 1693170804
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1693170804
transform -1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_32
timestamp 1693170804
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1693170804
transform -1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_33
timestamp 1693170804
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1693170804
transform -1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_34
timestamp 1693170804
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1693170804
transform -1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_35
timestamp 1693170804
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1693170804
transform -1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_36
timestamp 1693170804
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1693170804
transform -1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_37
timestamp 1693170804
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1693170804
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_38
timestamp 1693170804
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1693170804
transform -1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_39
timestamp 1693170804
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1693170804
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_40
timestamp 1693170804
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1693170804
transform -1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_41
timestamp 1693170804
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1693170804
transform -1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_42
timestamp 1693170804
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1693170804
transform -1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_43
timestamp 1693170804
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1693170804
transform -1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_44
timestamp 1693170804
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1693170804
transform -1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_45
timestamp 1693170804
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1693170804
transform -1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_46
timestamp 1693170804
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1693170804
transform -1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_47
timestamp 1693170804
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1693170804
transform -1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_48
timestamp 1693170804
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1693170804
transform -1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_49
timestamp 1693170804
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1693170804
transform -1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_51
timestamp 1693170804
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_52
timestamp 1693170804
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_53
timestamp 1693170804
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_54
timestamp 1693170804
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_55
timestamp 1693170804
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_56
timestamp 1693170804
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_57
timestamp 1693170804
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_58
timestamp 1693170804
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_59
timestamp 1693170804
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_60
timestamp 1693170804
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_61
timestamp 1693170804
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp 1693170804
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp 1693170804
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp 1693170804
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_65
timestamp 1693170804
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp 1693170804
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_67
timestamp 1693170804
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_68
timestamp 1693170804
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_69
timestamp 1693170804
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_70
timestamp 1693170804
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_71
timestamp 1693170804
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_72
timestamp 1693170804
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_73
timestamp 1693170804
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_74
timestamp 1693170804
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_75
timestamp 1693170804
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_76
timestamp 1693170804
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_77
timestamp 1693170804
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_78
timestamp 1693170804
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_79
timestamp 1693170804
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_80
timestamp 1693170804
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_81
timestamp 1693170804
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_82
timestamp 1693170804
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_83
timestamp 1693170804
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_84
timestamp 1693170804
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_85
timestamp 1693170804
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_86
timestamp 1693170804
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_87
timestamp 1693170804
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_88
timestamp 1693170804
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_89
timestamp 1693170804
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_90
timestamp 1693170804
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_91
timestamp 1693170804
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_92
timestamp 1693170804
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_93
timestamp 1693170804
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_94
timestamp 1693170804
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_95
timestamp 1693170804
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_96
timestamp 1693170804
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_97
timestamp 1693170804
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_98
timestamp 1693170804
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_99
timestamp 1693170804
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_100
timestamp 1693170804
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_101
timestamp 1693170804
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_102
timestamp 1693170804
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_103
timestamp 1693170804
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_104
timestamp 1693170804
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_105
timestamp 1693170804
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_106
timestamp 1693170804
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_107
timestamp 1693170804
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_108
timestamp 1693170804
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_109
timestamp 1693170804
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_110
timestamp 1693170804
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_111
timestamp 1693170804
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_112
timestamp 1693170804
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_113
timestamp 1693170804
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_114
timestamp 1693170804
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_115
timestamp 1693170804
transform 1 0 11408 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_116
timestamp 1693170804
transform 1 0 13984 0 1 15232
box -38 -48 130 592
<< labels >>
flabel metal4 s 1604 2128 1924 15824 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5604 2128 5924 15824 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9604 2128 9924 15824 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 13604 2128 13924 15824 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 2676 16884 2996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6676 16884 6996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 10676 16884 10996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 14676 16884 14996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 944 2016 1264 15824 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4944 2016 5264 15824 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8944 2016 9264 15824 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2016 13264 15824 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 944 2016 16884 2336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 944 6016 16884 6336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 944 10016 16884 10336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 944 14016 16884 14336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 cal
port 2 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 clk
port 3 nsew signal input
flabel metal2 s 9034 17200 9090 18000 0 FreeSans 224 90 0 0 clkc
port 4 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 comp
port 5 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 ctln[0]
port 6 nsew signal tristate
flabel metal3 s 17200 8 18000 128 0 FreeSans 480 0 0 0 ctln[1]
port 7 nsew signal tristate
flabel metal3 s 17200 10888 18000 11008 0 FreeSans 480 0 0 0 ctln[2]
port 8 nsew signal tristate
flabel metal2 s 662 17200 718 18000 0 FreeSans 224 90 0 0 ctln[3]
port 9 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 ctln[4]
port 10 nsew signal tristate
flabel metal2 s 14186 17200 14242 18000 0 FreeSans 224 90 0 0 ctln[5]
port 11 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 ctln[6]
port 12 nsew signal tristate
flabel metal3 s 17200 12928 18000 13048 0 FreeSans 480 0 0 0 ctln[7]
port 13 nsew signal tristate
flabel metal3 s 17200 2048 18000 2168 0 FreeSans 480 0 0 0 ctlp[0]
port 14 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 ctlp[1]
port 15 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 ctlp[2]
port 16 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 ctlp[3]
port 17 nsew signal tristate
flabel metal2 s 10966 17200 11022 18000 0 FreeSans 224 90 0 0 ctlp[4]
port 18 nsew signal tristate
flabel metal2 s 16118 17200 16174 18000 0 FreeSans 224 90 0 0 ctlp[5]
port 19 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 ctlp[6]
port 20 nsew signal tristate
flabel metal3 s 17200 14288 18000 14408 0 FreeSans 480 0 0 0 ctlp[7]
port 21 nsew signal tristate
flabel metal2 s 4526 17200 4582 18000 0 FreeSans 224 90 0 0 en
port 22 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 result[0]
port 23 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 result[1]
port 24 nsew signal tristate
flabel metal3 s 17200 8848 18000 8968 0 FreeSans 480 0 0 0 result[2]
port 25 nsew signal tristate
flabel metal2 s 2594 17200 2650 18000 0 FreeSans 224 90 0 0 result[3]
port 26 nsew signal tristate
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 result[4]
port 27 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 result[5]
port 28 nsew signal tristate
flabel metal2 s 12898 17200 12954 18000 0 FreeSans 224 90 0 0 result[6]
port 29 nsew signal tristate
flabel metal3 s 17200 4088 18000 4208 0 FreeSans 480 0 0 0 result[7]
port 30 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 rstn
port 31 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 sample
port 32 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 trim[0]
port 33 nsew signal tristate
flabel metal3 s 17200 5448 18000 5568 0 FreeSans 480 0 0 0 trim[1]
port 34 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 trim[2]
port 35 nsew signal tristate
flabel metal3 s 17200 16328 18000 16448 0 FreeSans 480 0 0 0 trim[3]
port 36 nsew signal tristate
flabel metal2 s 17406 17200 17462 18000 0 FreeSans 224 90 0 0 trim[4]
port 37 nsew signal tristate
flabel metal2 s 5814 17200 5870 18000 0 FreeSans 224 90 0 0 trimb[0]
port 38 nsew signal tristate
flabel metal2 s 7746 17200 7802 18000 0 FreeSans 224 90 0 0 trimb[1]
port 39 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 trimb[2]
port 40 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 trimb[3]
port 41 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 trimb[4]
port 42 nsew signal tristate
flabel metal3 s 17200 7488 18000 7608 0 FreeSans 480 0 0 0 valid
port 43 nsew signal tristate
rlabel metal1 8970 15232 8970 15232 0 VGND
rlabel metal1 8890 15776 8890 15776 0 VPWR
rlabel metal1 6522 6970 6522 6970 0 _000_
rlabel metal1 10856 8874 10856 8874 0 _001_
rlabel metal1 6762 8874 6762 8874 0 _002_
rlabel metal1 7728 5270 7728 5270 0 _003_
rlabel metal1 8694 6698 8694 6698 0 _004_
rlabel metal2 1978 5440 1978 5440 0 _005_
rlabel metal1 13984 4182 13984 4182 0 _006_
rlabel metal1 1932 4182 1932 4182 0 _007_
rlabel metal1 14352 9146 14352 9146 0 _008_
rlabel metal2 1702 13464 1702 13464 0 _009_
rlabel metal1 1610 10710 1610 10710 0 _010_
rlabel metal1 14306 12274 14306 12274 0 _011_
rlabel metal1 11730 12954 11730 12954 0 _012_
rlabel metal1 14628 7310 14628 7310 0 _013_
rlabel metal1 3910 5304 3910 5304 0 _014_
rlabel metal1 14131 6970 14131 6970 0 _015_
rlabel metal1 11822 7480 11822 7480 0 _016_
rlabel metal1 11362 10098 11362 10098 0 _017_
rlabel metal1 10672 11322 10672 11322 0 _018_
rlabel metal1 9890 10506 9890 10506 0 _019_
rlabel metal2 13386 11118 13386 11118 0 _020_
rlabel metal1 11546 10778 11546 10778 0 _021_
rlabel metal1 13708 8058 13708 8058 0 _022_
rlabel metal1 5290 4046 5290 4046 0 _023_
rlabel metal1 9430 3094 9430 3094 0 _024_
rlabel metal1 9890 4182 9890 4182 0 _025_
rlabel metal1 9936 5338 9936 5338 0 _026_
rlabel metal1 6440 5678 6440 5678 0 _027_
rlabel metal1 4278 3094 4278 3094 0 _028_
rlabel metal1 6992 2482 6992 2482 0 _029_
rlabel metal1 12742 2958 12742 2958 0 _030_
rlabel metal2 12650 4590 12650 4590 0 _031_
rlabel metal1 7130 10710 7130 10710 0 _032_
rlabel metal1 8878 8364 8878 8364 0 _033_
rlabel metal2 3634 11866 3634 11866 0 _034_
rlabel metal2 2898 12852 2898 12852 0 _035_
rlabel metal1 5382 12614 5382 12614 0 _036_
rlabel metal1 5198 10472 5198 10472 0 _037_
rlabel metal1 2162 9146 2162 9146 0 _038_
rlabel metal1 3036 7922 3036 7922 0 _039_
rlabel metal1 2162 5338 2162 5338 0 _040_
rlabel metal1 4600 6630 4600 6630 0 _041_
rlabel metal1 5750 10030 5750 10030 0 _042_
rlabel metal1 8740 8398 8740 8398 0 _043_
rlabel metal1 7636 7514 7636 7514 0 _044_
rlabel metal1 7268 6834 7268 6834 0 _045_
rlabel metal1 8648 6834 8648 6834 0 _046_
rlabel metal1 5796 9146 5796 9146 0 _047_
rlabel metal1 6164 8942 6164 8942 0 _048_
rlabel metal1 10626 10744 10626 10744 0 _049_
rlabel metal1 10534 6392 10534 6392 0 _050_
rlabel metal1 14720 3026 14720 3026 0 _051_
rlabel metal1 3864 3502 3864 3502 0 _052_
rlabel metal2 14950 10438 14950 10438 0 _053_
rlabel metal1 2070 12172 2070 12172 0 _054_
rlabel metal1 3312 11322 3312 11322 0 _055_
rlabel metal2 15134 12342 15134 12342 0 _056_
rlabel metal2 12558 12104 12558 12104 0 _057_
rlabel metal1 15824 8602 15824 8602 0 _058_
rlabel metal1 6348 3502 6348 3502 0 _059_
rlabel metal2 8142 4114 8142 4114 0 _060_
rlabel metal2 11362 2618 11362 2618 0 _061_
rlabel metal2 12374 5508 12374 5508 0 _062_
rlabel metal1 10120 10234 10120 10234 0 _063_
rlabel metal1 9798 13226 9798 13226 0 _064_
rlabel metal1 6164 7854 6164 7854 0 _065_
rlabel metal1 4646 8874 4646 8874 0 _066_
rlabel metal1 4876 8058 4876 8058 0 _067_
rlabel metal1 5290 12682 5290 12682 0 _068_
rlabel metal1 4646 7922 4646 7922 0 _069_
rlabel metal1 2599 8942 2599 8942 0 _070_
rlabel metal1 5060 7990 5060 7990 0 _071_
rlabel metal1 4416 7854 4416 7854 0 _072_
rlabel metal2 3358 6120 3358 6120 0 _073_
rlabel metal1 2162 6290 2162 6290 0 _074_
rlabel metal2 2438 6630 2438 6630 0 _075_
rlabel metal1 2162 5168 2162 5168 0 _076_
rlabel metal1 8656 11050 8656 11050 0 _077_
rlabel metal1 13846 7854 13846 7854 0 _078_
rlabel metal1 2438 12750 2438 12750 0 _079_
rlabel metal2 2714 12257 2714 12257 0 _080_
rlabel metal1 2622 11220 2622 11220 0 _081_
rlabel metal1 13570 4624 13570 4624 0 _082_
rlabel metal1 14030 4590 14030 4590 0 _083_
rlabel metal1 2254 4624 2254 4624 0 _084_
rlabel metal1 2024 4590 2024 4590 0 _085_
rlabel metal1 13202 9520 13202 9520 0 _086_
rlabel metal1 13938 8942 13938 8942 0 _087_
rlabel metal1 2254 12410 2254 12410 0 _088_
rlabel metal2 1978 13430 1978 13430 0 _089_
rlabel metal1 2162 11152 2162 11152 0 _090_
rlabel metal1 1932 11118 1932 11118 0 _091_
rlabel metal1 14122 11866 14122 11866 0 _092_
rlabel metal1 13432 12206 13432 12206 0 _093_
rlabel metal1 11822 12410 11822 12410 0 _094_
rlabel metal1 12052 12818 12052 12818 0 _095_
rlabel metal1 15042 7888 15042 7888 0 _096_
rlabel metal1 15364 7854 15364 7854 0 _097_
rlabel metal1 4981 5678 4981 5678 0 _098_
rlabel metal1 14398 6698 14398 6698 0 _099_
rlabel via1 11536 7854 11536 7854 0 _100_
rlabel metal1 10902 10030 10902 10030 0 _101_
rlabel metal1 10534 11084 10534 11084 0 _102_
rlabel metal1 9890 10608 9890 10608 0 _103_
rlabel metal2 12742 11050 12742 11050 0 _104_
rlabel metal1 12696 9078 12696 9078 0 _105_
rlabel viali 11170 5270 11170 5270 0 _106_
rlabel metal2 7314 4471 7314 4471 0 _107_
rlabel metal2 6854 4386 6854 4386 0 _108_
rlabel metal1 8786 4114 8786 4114 0 _109_
rlabel metal1 8786 3706 8786 3706 0 _110_
rlabel metal1 10350 5202 10350 5202 0 _111_
rlabel metal2 10902 4080 10902 4080 0 _112_
rlabel metal1 5934 3060 5934 3060 0 _113_
rlabel metal2 10534 3774 10534 3774 0 _114_
rlabel metal1 5520 3026 5520 3026 0 _115_
rlabel metal1 7130 3026 7130 3026 0 _116_
rlabel metal1 7498 2992 7498 2992 0 _117_
rlabel metal1 10672 3026 10672 3026 0 _118_
rlabel metal2 10902 2618 10902 2618 0 _119_
rlabel metal1 11730 4556 11730 4556 0 _120_
rlabel metal1 11730 4114 11730 4114 0 _121_
rlabel metal1 7222 9962 7222 9962 0 _122_
rlabel metal1 6992 10234 6992 10234 0 _123_
rlabel metal2 8970 8772 8970 8772 0 _124_
rlabel metal1 8878 8500 8878 8500 0 _125_
rlabel metal1 4508 12818 4508 12818 0 _126_
rlabel metal2 3910 11764 3910 11764 0 _127_
rlabel metal1 4600 13974 4600 13974 0 _128_
rlabel metal1 4922 13906 4922 13906 0 _129_
rlabel metal2 4646 13668 4646 13668 0 _130_
rlabel metal2 4738 13260 4738 13260 0 _131_
rlabel metal1 7314 13260 7314 13260 0 _132_
rlabel via1 7406 13362 7406 13362 0 _133_
rlabel metal1 7084 13294 7084 13294 0 _134_
rlabel metal2 7314 13056 7314 13056 0 _135_
rlabel metal1 5520 12818 5520 12818 0 _136_
rlabel metal1 5888 10642 5888 10642 0 _137_
rlabel metal2 7038 12789 7038 12789 0 _138_
rlabel metal1 6670 11662 6670 11662 0 _139_
rlabel metal1 6026 10574 6026 10574 0 _140_
rlabel metal3 751 4828 751 4828 0 cal
rlabel metal1 4462 13906 4462 13906 0 cal_count\[0\]
rlabel metal1 5336 13362 5336 13362 0 cal_count\[1\]
rlabel metal1 7176 12750 7176 12750 0 cal_count\[2\]
rlabel metal2 6762 10336 6762 10336 0 cal_count\[3\]
rlabel metal1 2438 7378 2438 7378 0 cal_itt\[0\]
rlabel metal1 2714 7276 2714 7276 0 cal_itt\[1\]
rlabel metal2 3174 7174 3174 7174 0 cal_itt\[2\]
rlabel metal1 4370 5780 4370 5780 0 cal_itt\[3\]
rlabel metal2 6762 5474 6762 5474 0 calibrate
rlabel metal2 12926 1639 12926 1639 0 clk
rlabel metal1 9246 15674 9246 15674 0 clkc
rlabel metal1 10948 5678 10948 5678 0 clknet_0_clk
rlabel metal1 1426 6732 1426 6732 0 clknet_2_0__leaf_clk
rlabel metal1 1610 9554 1610 9554 0 clknet_2_1__leaf_clk
rlabel metal1 13800 4046 13800 4046 0 clknet_2_2__leaf_clk
rlabel metal1 13754 9554 13754 9554 0 clknet_2_3__leaf_clk
rlabel metal3 751 13668 751 13668 0 comp
rlabel metal1 16606 2822 16606 2822 0 ctln[0]
rlabel metal2 16422 1173 16422 1173 0 ctln[1]
rlabel metal1 16468 11186 16468 11186 0 ctln[2]
rlabel metal1 1334 15470 1334 15470 0 ctln[3]
rlabel metal3 751 15708 751 15708 0 ctln[4]
rlabel metal2 14214 16943 14214 16943 0 ctln[5]
rlabel metal2 9706 823 9706 823 0 ctln[6]
rlabel metal2 16974 13073 16974 13073 0 ctln[7]
rlabel metal2 16974 2227 16974 2227 0 ctlp[0]
rlabel metal2 3266 1520 3266 1520 0 ctlp[1]
rlabel metal3 1096 12308 1096 12308 0 ctlp[2]
rlabel metal3 820 8908 820 8908 0 ctlp[3]
rlabel metal1 11408 15674 11408 15674 0 ctlp[4]
rlabel metal2 16199 17340 16199 17340 0 ctlp[5]
rlabel metal3 751 10268 751 10268 0 ctlp[6]
rlabel via2 16974 14331 16974 14331 0 ctlp[7]
rlabel metal1 4600 15470 4600 15470 0 en
rlabel metal1 9752 13430 9752 13430 0 en_co_clk
rlabel metal2 13018 4539 13018 4539 0 mask\[0\]
rlabel metal1 12926 7956 12926 7956 0 mask\[1\]
rlabel metal1 13892 9894 13892 9894 0 mask\[2\]
rlabel metal2 9246 12614 9246 12614 0 mask\[3\]
rlabel metal1 3220 11050 3220 11050 0 mask\[4\]
rlabel metal2 14858 10336 14858 10336 0 mask\[5\]
rlabel metal1 12696 11322 12696 11322 0 mask\[6\]
rlabel metal1 14582 8602 14582 8602 0 mask\[7\]
rlabel metal1 1610 5304 1610 5304 0 net1
rlabel metal1 1978 14994 1978 14994 0 net10
rlabel metal1 14766 15130 14766 15130 0 net11
rlabel metal2 9890 2587 9890 2587 0 net12
rlabel metal2 16146 13090 16146 13090 0 net13
rlabel metal1 15686 2448 15686 2448 0 net14
rlabel metal2 15686 3247 15686 3247 0 net15
rlabel metal1 2208 12886 2208 12886 0 net16
rlabel metal1 1932 12070 1932 12070 0 net17
rlabel metal1 2254 14960 2254 14960 0 net18
rlabel metal1 15134 14994 15134 14994 0 net19
rlabel metal1 6164 13906 6164 13906 0 net2
rlabel metal1 2277 10030 2277 10030 0 net20
rlabel metal2 15962 13634 15962 13634 0 net21
rlabel metal2 12466 3774 12466 3774 0 net22
rlabel metal2 3358 3706 3358 3706 0 net23
rlabel metal1 16008 9350 16008 9350 0 net24
rlabel metal1 3128 13498 3128 13498 0 net25
rlabel metal1 2530 2414 2530 2414 0 net26
rlabel metal2 15134 2587 15134 2587 0 net27
rlabel metal1 12880 13498 12880 13498 0 net28
rlabel metal1 16008 7174 16008 7174 0 net29
rlabel metal1 5428 15334 5428 15334 0 net3
rlabel metal2 6946 9894 6946 9894 0 net30
rlabel metal1 6210 2414 6210 2414 0 net31
rlabel metal1 14283 5610 14283 5610 0 net32
rlabel metal1 9936 2550 9936 2550 0 net33
rlabel metal2 16100 13396 16100 13396 0 net34
rlabel metal1 15594 12920 15594 12920 0 net35
rlabel metal1 6302 15130 6302 15130 0 net36
rlabel metal1 8188 15130 8188 15130 0 net37
rlabel metal1 11638 2414 11638 2414 0 net38
rlabel metal1 1794 6256 1794 6256 0 net39
rlabel metal2 3266 3876 3266 3876 0 net4
rlabel metal1 1794 15368 1794 15368 0 net40
rlabel metal1 15870 7854 15870 7854 0 net41
rlabel metal1 4009 12886 4009 12886 0 net42
rlabel metal2 8050 5984 8050 5984 0 net43
rlabel metal1 12703 13226 12703 13226 0 net44
rlabel metal2 9154 2958 9154 2958 0 net45
rlabel metal1 11362 8874 11362 8874 0 net46
rlabel metal1 4600 9554 4600 9554 0 net47
rlabel metal1 9246 8976 9246 8976 0 net48
rlabel metal2 7130 5950 7130 5950 0 net49
rlabel metal1 9476 13498 9476 13498 0 net5
rlabel metal1 9285 6970 9285 6970 0 net50
rlabel metal2 2806 5491 2806 5491 0 net51
rlabel metal1 7153 5610 7153 5610 0 net52
rlabel metal2 6118 5100 6118 5100 0 net53
rlabel metal2 12834 10880 12834 10880 0 net54
rlabel metal1 13800 7922 13800 7922 0 net55
rlabel metal1 12006 9656 12006 9656 0 net56
rlabel metal1 9522 5134 9522 5134 0 net57
rlabel metal1 6578 4114 6578 4114 0 net58
rlabel metal2 14122 11560 14122 11560 0 net59
rlabel metal1 16146 3128 16146 3128 0 net6
rlabel metal1 10028 10642 10028 10642 0 net60
rlabel metal1 10396 11118 10396 11118 0 net61
rlabel metal1 8878 3978 8878 3978 0 net62
rlabel metal1 7820 6222 7820 6222 0 net63
rlabel metal1 11362 7922 11362 7922 0 net64
rlabel metal1 13110 7174 13110 7174 0 net65
rlabel metal1 8142 10030 8142 10030 0 net66
rlabel metal1 3726 5882 3726 5882 0 net67
rlabel metal1 7176 9146 7176 9146 0 net68
rlabel metal1 7360 11118 7360 11118 0 net69
rlabel metal1 15962 2414 15962 2414 0 net7
rlabel metal1 5014 12886 5014 12886 0 net70
rlabel metal1 6072 12818 6072 12818 0 net71
rlabel metal1 16008 11050 16008 11050 0 net8
rlabel metal1 2392 15130 2392 15130 0 net9
rlabel metal1 782 2822 782 2822 0 result[0]
rlabel metal3 820 3468 820 3468 0 result[1]
rlabel metal1 16652 8874 16652 8874 0 result[2]
rlabel metal2 2622 16943 2622 16943 0 result[3]
rlabel metal3 820 1428 820 1428 0 result[4]
rlabel metal2 14858 1520 14858 1520 0 result[5]
rlabel metal2 12926 16943 12926 16943 0 result[6]
rlabel metal1 16606 4454 16606 4454 0 result[7]
rlabel metal1 1656 3026 1656 3026 0 rstn
rlabel metal2 4554 1520 4554 1520 0 sample
rlabel metal1 6325 9486 6325 9486 0 state\[0\]
rlabel metal2 7314 6562 7314 6562 0 state\[2\]
rlabel metal1 9292 8466 9292 8466 0 state\[3\]
rlabel metal1 11362 5304 11362 5304 0 state\[4\]
rlabel metal1 10028 7378 10028 7378 0 state\[5\]
rlabel metal2 6486 1520 6486 1520 0 trim[0]
rlabel metal1 16468 5542 16468 5542 0 trim[1]
rlabel metal2 8418 1520 8418 1520 0 trim[2]
rlabel metal1 16468 15130 16468 15130 0 trim[3]
rlabel metal2 17434 16466 17434 16466 0 trim[4]
rlabel metal1 5612 6086 5612 6086 0 trim_mask\[0\]
rlabel metal1 8004 3434 8004 3434 0 trim_mask\[1\]
rlabel metal1 10856 3366 10856 3366 0 trim_mask\[2\]
rlabel metal1 11408 4454 11408 4454 0 trim_mask\[3\]
rlabel metal1 8464 5746 8464 5746 0 trim_mask\[4\]
rlabel metal2 5474 3230 5474 3230 0 trim_val\[0\]
rlabel metal1 8004 2618 8004 2618 0 trim_val\[1\]
rlabel metal1 11270 3094 11270 3094 0 trim_val\[2\]
rlabel metal1 11178 4624 11178 4624 0 trim_val\[3\]
rlabel metal1 9108 10574 9108 10574 0 trim_val\[4\]
rlabel metal1 6210 15674 6210 15674 0 trimb[0]
rlabel metal1 7912 15674 7912 15674 0 trimb[1]
rlabel metal2 11638 1520 11638 1520 0 trimb[2]
rlabel metal3 820 6868 820 6868 0 trimb[3]
rlabel metal3 1096 17748 1096 17748 0 trimb[4]
rlabel metal1 16606 7718 16606 7718 0 valid
<< properties >>
string FIXED_BBOX 0 0 18000 18000
<< end >>
