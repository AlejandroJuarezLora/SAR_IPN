magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 1142 542
<< pwell >>
rect 1 -19 1027 163
rect 30 -57 64 -19
<< scnmos >>
rect 79 7 109 137
rect 163 7 193 137
rect 247 7 277 137
rect 331 7 361 137
rect 415 7 445 137
rect 499 7 529 137
rect 583 7 613 137
rect 667 7 697 137
rect 751 7 781 137
rect 835 7 865 137
rect 919 7 949 137
<< scpmoshvt >>
rect 79 257 109 457
rect 163 257 193 457
rect 247 257 277 457
rect 331 257 361 457
rect 415 257 445 457
rect 499 257 529 457
rect 583 257 613 457
rect 667 257 697 457
rect 751 257 781 457
rect 835 257 865 457
rect 919 257 949 457
<< ndiff >>
rect 27 89 79 137
rect 27 55 35 89
rect 69 55 79 89
rect 27 7 79 55
rect 109 57 163 137
rect 109 23 119 57
rect 153 23 163 57
rect 109 7 163 23
rect 193 89 247 137
rect 193 55 203 89
rect 237 55 247 89
rect 193 7 247 55
rect 277 57 331 137
rect 277 23 287 57
rect 321 23 331 57
rect 277 7 331 23
rect 361 89 415 137
rect 361 55 371 89
rect 405 55 415 89
rect 361 7 415 55
rect 445 57 499 137
rect 445 23 455 57
rect 489 23 499 57
rect 445 7 499 23
rect 529 89 583 137
rect 529 55 539 89
rect 573 55 583 89
rect 529 7 583 55
rect 613 57 667 137
rect 613 23 623 57
rect 657 23 667 57
rect 613 7 667 23
rect 697 89 751 137
rect 697 55 707 89
rect 741 55 751 89
rect 697 7 751 55
rect 781 57 835 137
rect 781 23 791 57
rect 825 23 835 57
rect 781 7 835 23
rect 865 89 919 137
rect 865 55 875 89
rect 909 55 919 89
rect 865 7 919 55
rect 949 121 1001 137
rect 949 87 959 121
rect 993 87 1001 121
rect 949 53 1001 87
rect 949 19 959 53
rect 993 19 1001 53
rect 949 7 1001 19
<< pdiff >>
rect 27 439 79 457
rect 27 405 35 439
rect 69 405 79 439
rect 27 371 79 405
rect 27 337 35 371
rect 69 337 79 371
rect 27 303 79 337
rect 27 269 35 303
rect 69 269 79 303
rect 27 257 79 269
rect 109 445 163 457
rect 109 411 119 445
rect 153 411 163 445
rect 109 377 163 411
rect 109 343 119 377
rect 153 343 163 377
rect 109 257 163 343
rect 193 439 247 457
rect 193 405 203 439
rect 237 405 247 439
rect 193 371 247 405
rect 193 337 203 371
rect 237 337 247 371
rect 193 303 247 337
rect 193 269 203 303
rect 237 269 247 303
rect 193 257 247 269
rect 277 445 331 457
rect 277 411 287 445
rect 321 411 331 445
rect 277 377 331 411
rect 277 343 287 377
rect 321 343 331 377
rect 277 257 331 343
rect 361 423 415 457
rect 361 389 371 423
rect 405 389 415 423
rect 361 328 415 389
rect 361 294 371 328
rect 405 294 415 328
rect 361 257 415 294
rect 445 445 499 457
rect 445 411 455 445
rect 489 411 499 445
rect 445 377 499 411
rect 445 343 455 377
rect 489 343 499 377
rect 445 257 499 343
rect 529 423 583 457
rect 529 389 539 423
rect 573 389 583 423
rect 529 328 583 389
rect 529 294 539 328
rect 573 294 583 328
rect 529 257 583 294
rect 613 445 667 457
rect 613 411 623 445
rect 657 411 667 445
rect 613 377 667 411
rect 613 343 623 377
rect 657 343 667 377
rect 613 257 667 343
rect 697 423 751 457
rect 697 389 707 423
rect 741 389 751 423
rect 697 328 751 389
rect 697 294 707 328
rect 741 294 751 328
rect 697 257 751 294
rect 781 445 835 457
rect 781 411 791 445
rect 825 411 835 445
rect 781 377 835 411
rect 781 343 791 377
rect 825 343 835 377
rect 781 257 835 343
rect 865 423 919 457
rect 865 389 875 423
rect 909 389 919 423
rect 865 328 919 389
rect 865 294 875 328
rect 909 294 919 328
rect 865 257 919 294
rect 949 445 1001 457
rect 949 411 959 445
rect 993 411 1001 445
rect 949 377 1001 411
rect 949 343 959 377
rect 993 343 1001 377
rect 949 309 1001 343
rect 949 275 959 309
rect 993 275 1001 309
rect 949 257 1001 275
<< ndiffc >>
rect 35 55 69 89
rect 119 23 153 57
rect 203 55 237 89
rect 287 23 321 57
rect 371 55 405 89
rect 455 23 489 57
rect 539 55 573 89
rect 623 23 657 57
rect 707 55 741 89
rect 791 23 825 57
rect 875 55 909 89
rect 959 87 993 121
rect 959 19 993 53
<< pdiffc >>
rect 35 405 69 439
rect 35 337 69 371
rect 35 269 69 303
rect 119 411 153 445
rect 119 343 153 377
rect 203 405 237 439
rect 203 337 237 371
rect 203 269 237 303
rect 287 411 321 445
rect 287 343 321 377
rect 371 389 405 423
rect 371 294 405 328
rect 455 411 489 445
rect 455 343 489 377
rect 539 389 573 423
rect 539 294 573 328
rect 623 411 657 445
rect 623 343 657 377
rect 707 389 741 423
rect 707 294 741 328
rect 791 411 825 445
rect 791 343 825 377
rect 875 389 909 423
rect 875 294 909 328
rect 959 411 993 445
rect 959 343 993 377
rect 959 275 993 309
<< poly >>
rect 79 457 109 483
rect 163 457 193 483
rect 247 457 277 483
rect 331 457 361 483
rect 415 457 445 483
rect 499 457 529 483
rect 583 457 613 483
rect 667 457 697 483
rect 751 457 781 483
rect 835 457 865 483
rect 919 457 949 483
rect 79 221 109 257
rect 28 219 109 221
rect 163 219 193 257
rect 247 219 277 257
rect 28 209 277 219
rect 28 175 44 209
rect 78 175 112 209
rect 146 175 180 209
rect 214 175 277 209
rect 28 165 277 175
rect 28 163 109 165
rect 79 137 109 163
rect 163 137 193 165
rect 247 137 277 165
rect 331 219 361 257
rect 415 219 445 257
rect 499 219 529 257
rect 583 219 613 257
rect 667 219 697 257
rect 751 219 781 257
rect 835 219 865 257
rect 919 219 949 257
rect 331 209 949 219
rect 331 175 351 209
rect 385 175 419 209
rect 453 175 487 209
rect 521 175 555 209
rect 589 175 623 209
rect 657 175 691 209
rect 725 175 759 209
rect 793 175 949 209
rect 331 165 949 175
rect 331 137 361 165
rect 415 137 445 165
rect 499 137 529 165
rect 583 137 613 165
rect 667 137 697 165
rect 751 137 781 165
rect 835 137 865 165
rect 919 137 949 165
rect 79 -19 109 7
rect 163 -19 193 7
rect 247 -19 277 7
rect 331 -19 361 7
rect 415 -19 445 7
rect 499 -19 529 7
rect 583 -19 613 7
rect 667 -19 697 7
rect 751 -19 781 7
rect 835 -19 865 7
rect 919 -19 949 7
<< polycont >>
rect 44 175 78 209
rect 112 175 146 209
rect 180 175 214 209
rect 351 175 385 209
rect 419 175 453 209
rect 487 175 521 209
rect 555 175 589 209
rect 623 175 657 209
rect 691 175 725 209
rect 759 175 793 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1104 521
rect 19 439 85 453
rect 19 405 35 439
rect 69 405 85 439
rect 19 371 85 405
rect 19 337 35 371
rect 69 337 85 371
rect 19 303 85 337
rect 119 445 153 487
rect 119 377 153 411
rect 119 327 153 343
rect 187 439 253 453
rect 187 405 203 439
rect 237 405 253 439
rect 187 371 253 405
rect 187 337 203 371
rect 237 337 253 371
rect 19 269 35 303
rect 69 283 85 303
rect 187 303 253 337
rect 287 445 321 487
rect 287 377 321 411
rect 287 327 321 343
rect 371 423 405 453
rect 371 328 405 389
rect 187 283 203 303
rect 69 269 203 283
rect 237 283 253 303
rect 439 445 505 487
rect 439 411 455 445
rect 489 411 505 445
rect 439 377 505 411
rect 439 343 455 377
rect 489 343 505 377
rect 439 327 505 343
rect 539 423 573 453
rect 539 328 573 389
rect 371 283 405 294
rect 607 445 673 487
rect 607 411 623 445
rect 657 411 673 445
rect 607 377 673 411
rect 607 343 623 377
rect 657 343 673 377
rect 607 327 673 343
rect 707 423 741 453
rect 707 328 741 389
rect 539 283 573 294
rect 775 445 841 487
rect 775 411 791 445
rect 825 411 841 445
rect 775 377 841 411
rect 775 343 791 377
rect 825 343 841 377
rect 775 327 841 343
rect 875 423 909 453
rect 875 328 909 389
rect 707 283 741 294
rect 875 283 909 294
rect 237 269 319 283
rect 19 249 319 269
rect 371 249 909 283
rect 943 445 1009 487
rect 943 411 959 445
rect 993 411 1009 445
rect 943 377 1009 411
rect 943 343 959 377
rect 993 343 1009 377
rect 943 309 1009 343
rect 943 275 959 309
rect 993 275 1009 309
rect 943 257 1009 275
rect 28 209 248 215
rect 28 175 44 209
rect 78 175 112 209
rect 146 175 180 209
rect 214 175 248 209
rect 284 209 319 249
rect 284 175 351 209
rect 385 175 419 209
rect 453 175 487 209
rect 521 175 555 209
rect 589 175 623 209
rect 657 175 691 209
rect 725 175 759 209
rect 793 175 809 209
rect 284 141 319 175
rect 858 141 909 249
rect 35 107 319 141
rect 371 107 909 141
rect 35 89 69 107
rect 203 89 237 107
rect 35 11 69 55
rect 103 57 169 73
rect 103 23 119 57
rect 153 23 169 57
rect 103 -23 169 23
rect 371 89 405 107
rect 203 12 237 55
rect 271 57 337 73
rect 271 23 287 57
rect 321 23 337 57
rect 271 -23 337 23
rect 539 89 573 107
rect 371 11 405 55
rect 439 57 505 73
rect 439 23 455 57
rect 489 23 505 57
rect 439 -23 505 23
rect 707 89 741 107
rect 539 11 573 55
rect 607 57 673 73
rect 607 23 623 57
rect 657 23 673 57
rect 607 -23 673 23
rect 875 89 909 107
rect 707 11 741 55
rect 775 57 841 73
rect 775 23 791 57
rect 825 23 841 57
rect 775 -23 841 23
rect 875 11 909 55
rect 943 121 1009 137
rect 943 87 959 121
rect 993 87 1009 121
rect 943 53 1009 87
rect 943 19 959 53
rect 993 19 1009 53
rect 943 -23 1009 19
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1104 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 857 487 891 521
rect 949 487 983 521
rect 1041 487 1075 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
rect 857 -57 891 -23
rect 949 -57 983 -23
rect 1041 -57 1075 -23
<< metal1 >>
rect 0 521 1104 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1104 521
rect 0 456 1104 487
rect 0 -23 1104 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1104 -23
rect 0 -88 1104 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 buf_8
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 214 181 248 215 0 FreeSans 200 0 0 0 A
port 7 nsew
flabel locali s 858 113 892 147 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel locali s 858 181 892 215 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel locali s 122 181 156 215 0 FreeSans 200 0 0 0 A
port 7 nsew
flabel locali s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel locali s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel locali s 858 249 892 283 0 FreeSans 200 0 0 0 X
port 8 nsew
flabel locali s 30 181 64 215 0 FreeSans 200 0 0 0 A
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 1104 504
string path 0.000 -1.000 27.600 -1.000 
<< end >>
