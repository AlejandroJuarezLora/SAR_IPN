magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_p >>
rect -560 101 -502 107
rect -442 101 -384 107
rect -324 101 -266 107
rect -206 101 -148 107
rect -88 101 -30 107
rect 30 101 88 107
rect 148 101 206 107
rect 266 101 324 107
rect 384 101 442 107
rect 502 101 560 107
rect -560 67 -548 101
rect -442 67 -430 101
rect -324 67 -312 101
rect -206 67 -194 101
rect -88 67 -76 101
rect 30 67 42 101
rect 148 67 160 101
rect 266 67 278 101
rect 384 67 396 101
rect 502 67 514 101
rect -560 61 -502 67
rect -442 61 -384 67
rect -324 61 -266 67
rect -206 61 -148 67
rect -88 61 -30 67
rect 30 61 88 67
rect 148 61 206 67
rect 266 61 324 67
rect 384 61 442 67
rect 502 61 560 67
<< pwell >>
rect -747 -309 747 229
<< nmos >>
rect -561 -171 -501 29
rect -443 -171 -383 29
rect -325 -171 -265 29
rect -207 -171 -147 29
rect -89 -171 -29 29
rect 29 -171 89 29
rect 147 -171 207 29
rect 265 -171 325 29
rect 383 -171 443 29
rect 501 -171 561 29
<< ndiff >>
rect -619 14 -561 29
rect -619 -20 -607 14
rect -573 -20 -561 14
rect -619 -54 -561 -20
rect -619 -88 -607 -54
rect -573 -88 -561 -54
rect -619 -122 -561 -88
rect -619 -156 -607 -122
rect -573 -156 -561 -122
rect -619 -171 -561 -156
rect -501 14 -443 29
rect -501 -20 -489 14
rect -455 -20 -443 14
rect -501 -54 -443 -20
rect -501 -88 -489 -54
rect -455 -88 -443 -54
rect -501 -122 -443 -88
rect -501 -156 -489 -122
rect -455 -156 -443 -122
rect -501 -171 -443 -156
rect -383 14 -325 29
rect -383 -20 -371 14
rect -337 -20 -325 14
rect -383 -54 -325 -20
rect -383 -88 -371 -54
rect -337 -88 -325 -54
rect -383 -122 -325 -88
rect -383 -156 -371 -122
rect -337 -156 -325 -122
rect -383 -171 -325 -156
rect -265 14 -207 29
rect -265 -20 -253 14
rect -219 -20 -207 14
rect -265 -54 -207 -20
rect -265 -88 -253 -54
rect -219 -88 -207 -54
rect -265 -122 -207 -88
rect -265 -156 -253 -122
rect -219 -156 -207 -122
rect -265 -171 -207 -156
rect -147 14 -89 29
rect -147 -20 -135 14
rect -101 -20 -89 14
rect -147 -54 -89 -20
rect -147 -88 -135 -54
rect -101 -88 -89 -54
rect -147 -122 -89 -88
rect -147 -156 -135 -122
rect -101 -156 -89 -122
rect -147 -171 -89 -156
rect -29 14 29 29
rect -29 -20 -17 14
rect 17 -20 29 14
rect -29 -54 29 -20
rect -29 -88 -17 -54
rect 17 -88 29 -54
rect -29 -122 29 -88
rect -29 -156 -17 -122
rect 17 -156 29 -122
rect -29 -171 29 -156
rect 89 14 147 29
rect 89 -20 101 14
rect 135 -20 147 14
rect 89 -54 147 -20
rect 89 -88 101 -54
rect 135 -88 147 -54
rect 89 -122 147 -88
rect 89 -156 101 -122
rect 135 -156 147 -122
rect 89 -171 147 -156
rect 207 14 265 29
rect 207 -20 219 14
rect 253 -20 265 14
rect 207 -54 265 -20
rect 207 -88 219 -54
rect 253 -88 265 -54
rect 207 -122 265 -88
rect 207 -156 219 -122
rect 253 -156 265 -122
rect 207 -171 265 -156
rect 325 14 383 29
rect 325 -20 337 14
rect 371 -20 383 14
rect 325 -54 383 -20
rect 325 -88 337 -54
rect 371 -88 383 -54
rect 325 -122 383 -88
rect 325 -156 337 -122
rect 371 -156 383 -122
rect 325 -171 383 -156
rect 443 14 501 29
rect 443 -20 455 14
rect 489 -20 501 14
rect 443 -54 501 -20
rect 443 -88 455 -54
rect 489 -88 501 -54
rect 443 -122 501 -88
rect 443 -156 455 -122
rect 489 -156 501 -122
rect 443 -171 501 -156
rect 561 14 619 29
rect 561 -20 573 14
rect 607 -20 619 14
rect 561 -54 619 -20
rect 561 -88 573 -54
rect 607 -88 619 -54
rect 561 -122 619 -88
rect 561 -156 573 -122
rect 607 -156 619 -122
rect 561 -171 619 -156
<< ndiffc >>
rect -607 -20 -573 14
rect -607 -88 -573 -54
rect -607 -156 -573 -122
rect -489 -20 -455 14
rect -489 -88 -455 -54
rect -489 -156 -455 -122
rect -371 -20 -337 14
rect -371 -88 -337 -54
rect -371 -156 -337 -122
rect -253 -20 -219 14
rect -253 -88 -219 -54
rect -253 -156 -219 -122
rect -135 -20 -101 14
rect -135 -88 -101 -54
rect -135 -156 -101 -122
rect -17 -20 17 14
rect -17 -88 17 -54
rect -17 -156 17 -122
rect 101 -20 135 14
rect 101 -88 135 -54
rect 101 -156 135 -122
rect 219 -20 253 14
rect 219 -88 253 -54
rect 219 -156 253 -122
rect 337 -20 371 14
rect 337 -88 371 -54
rect 337 -156 371 -122
rect 455 -20 489 14
rect 455 -88 489 -54
rect 455 -156 489 -122
rect 573 -20 607 14
rect 573 -88 607 -54
rect 573 -156 607 -122
<< psubdiff >>
rect -721 169 -595 203
rect -561 169 -527 203
rect -493 169 -459 203
rect -425 169 -391 203
rect -357 169 -323 203
rect -289 169 -255 203
rect -221 169 -187 203
rect -153 169 -119 203
rect -85 169 -51 203
rect -17 169 17 203
rect 51 169 85 203
rect 119 169 153 203
rect 187 169 221 203
rect 255 169 289 203
rect 323 169 357 203
rect 391 169 425 203
rect 459 169 493 203
rect 527 169 561 203
rect 595 169 721 203
rect -721 79 -687 169
rect 687 79 721 169
rect -721 11 -687 45
rect -721 -57 -687 -23
rect -721 -125 -687 -91
rect -721 -249 -687 -159
rect 687 11 721 45
rect 687 -57 721 -23
rect 687 -125 721 -91
rect 687 -249 721 -159
rect -721 -283 -595 -249
rect -561 -283 -527 -249
rect -493 -283 -459 -249
rect -425 -283 -391 -249
rect -357 -283 -323 -249
rect -289 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 289 -249
rect 323 -283 357 -249
rect 391 -283 425 -249
rect 459 -283 493 -249
rect 527 -283 561 -249
rect 595 -283 721 -249
<< psubdiffcont >>
rect -595 169 -561 203
rect -527 169 -493 203
rect -459 169 -425 203
rect -391 169 -357 203
rect -323 169 -289 203
rect -255 169 -221 203
rect -187 169 -153 203
rect -119 169 -85 203
rect -51 169 -17 203
rect 17 169 51 203
rect 85 169 119 203
rect 153 169 187 203
rect 221 169 255 203
rect 289 169 323 203
rect 357 169 391 203
rect 425 169 459 203
rect 493 169 527 203
rect 561 169 595 203
rect -721 45 -687 79
rect 687 45 721 79
rect -721 -23 -687 11
rect -721 -91 -687 -57
rect -721 -159 -687 -125
rect 687 -23 721 11
rect 687 -91 721 -57
rect 687 -159 721 -125
rect -595 -283 -561 -249
rect -527 -283 -493 -249
rect -459 -283 -425 -249
rect -391 -283 -357 -249
rect -323 -283 -289 -249
rect -255 -283 -221 -249
rect -187 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 187 -249
rect 221 -283 255 -249
rect 289 -283 323 -249
rect 357 -283 391 -249
rect 425 -283 459 -249
rect 493 -283 527 -249
rect 561 -283 595 -249
<< poly >>
rect -564 101 -498 117
rect -564 67 -548 101
rect -514 67 -498 101
rect -564 51 -498 67
rect -446 101 -380 117
rect -446 67 -430 101
rect -396 67 -380 101
rect -446 51 -380 67
rect -328 101 -262 117
rect -328 67 -312 101
rect -278 67 -262 101
rect -328 51 -262 67
rect -210 101 -144 117
rect -210 67 -194 101
rect -160 67 -144 101
rect -210 51 -144 67
rect -92 101 -26 117
rect -92 67 -76 101
rect -42 67 -26 101
rect -92 51 -26 67
rect 26 101 92 117
rect 26 67 42 101
rect 76 67 92 101
rect 26 51 92 67
rect 144 101 210 117
rect 144 67 160 101
rect 194 67 210 101
rect 144 51 210 67
rect 262 101 328 117
rect 262 67 278 101
rect 312 67 328 101
rect 262 51 328 67
rect 380 101 446 117
rect 380 67 396 101
rect 430 67 446 101
rect 380 51 446 67
rect 498 101 564 117
rect 498 67 514 101
rect 548 67 564 101
rect 498 51 564 67
rect -561 29 -501 51
rect -443 29 -383 51
rect -325 29 -265 51
rect -207 29 -147 51
rect -89 29 -29 51
rect 29 29 89 51
rect 147 29 207 51
rect 265 29 325 51
rect 383 29 443 51
rect 501 29 561 51
rect -561 -197 -501 -171
rect -443 -197 -383 -171
rect -325 -197 -265 -171
rect -207 -197 -147 -171
rect -89 -197 -29 -171
rect 29 -197 89 -171
rect 147 -197 207 -171
rect 265 -197 325 -171
rect 383 -197 443 -171
rect 501 -197 561 -171
<< polycont >>
rect -548 67 -514 101
rect -430 67 -396 101
rect -312 67 -278 101
rect -194 67 -160 101
rect -76 67 -42 101
rect 42 67 76 101
rect 160 67 194 101
rect 278 67 312 101
rect 396 67 430 101
rect 514 67 548 101
<< locali >>
rect -721 169 -595 203
rect -561 169 -527 203
rect -493 169 -459 203
rect -425 169 -391 203
rect -357 169 -323 203
rect -289 169 -255 203
rect -221 169 -187 203
rect -153 169 -119 203
rect -85 169 -51 203
rect -17 169 17 203
rect 51 169 85 203
rect 119 169 153 203
rect 187 169 221 203
rect 255 169 289 203
rect 323 169 357 203
rect 391 169 425 203
rect 459 169 493 203
rect 527 169 561 203
rect 595 169 721 203
rect -721 79 -687 169
rect -564 67 -548 101
rect -514 67 -498 101
rect -446 67 -430 101
rect -396 67 -380 101
rect -328 67 -312 101
rect -278 67 -262 101
rect -210 67 -194 101
rect -160 67 -144 101
rect -92 67 -76 101
rect -42 67 -26 101
rect 26 67 42 101
rect 76 67 92 101
rect 144 67 160 101
rect 194 67 210 101
rect 262 67 278 101
rect 312 67 328 101
rect 380 67 396 101
rect 430 67 446 101
rect 498 67 514 101
rect 548 67 564 101
rect 687 79 721 169
rect -721 11 -687 45
rect -721 -57 -687 -23
rect -721 -125 -687 -91
rect -721 -249 -687 -159
rect -607 14 -573 33
rect -607 -54 -573 -52
rect -607 -90 -573 -88
rect -607 -175 -573 -156
rect -489 14 -455 33
rect -489 -54 -455 -52
rect -489 -90 -455 -88
rect -489 -175 -455 -156
rect -371 14 -337 33
rect -371 -54 -337 -52
rect -371 -90 -337 -88
rect -371 -175 -337 -156
rect -253 14 -219 33
rect -253 -54 -219 -52
rect -253 -90 -219 -88
rect -253 -175 -219 -156
rect -135 14 -101 33
rect -135 -54 -101 -52
rect -135 -90 -101 -88
rect -135 -175 -101 -156
rect -17 14 17 33
rect -17 -54 17 -52
rect -17 -90 17 -88
rect -17 -175 17 -156
rect 101 14 135 33
rect 101 -54 135 -52
rect 101 -90 135 -88
rect 101 -175 135 -156
rect 219 14 253 33
rect 219 -54 253 -52
rect 219 -90 253 -88
rect 219 -175 253 -156
rect 337 14 371 33
rect 337 -54 371 -52
rect 337 -90 371 -88
rect 337 -175 371 -156
rect 455 14 489 33
rect 455 -54 489 -52
rect 455 -90 489 -88
rect 455 -175 489 -156
rect 573 14 607 33
rect 573 -54 607 -52
rect 573 -90 607 -88
rect 573 -175 607 -156
rect 687 11 721 45
rect 687 -57 721 -23
rect 687 -125 721 -91
rect 687 -249 721 -159
rect -721 -283 -595 -249
rect -561 -283 -527 -249
rect -493 -283 -459 -249
rect -425 -283 -391 -249
rect -357 -283 -323 -249
rect -289 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 289 -249
rect 323 -283 357 -249
rect 391 -283 425 -249
rect 459 -283 493 -249
rect 527 -283 561 -249
rect 595 -283 721 -249
<< viali >>
rect -548 67 -514 101
rect -430 67 -396 101
rect -312 67 -278 101
rect -194 67 -160 101
rect -76 67 -42 101
rect 42 67 76 101
rect 160 67 194 101
rect 278 67 312 101
rect 396 67 430 101
rect 514 67 548 101
rect -607 -20 -573 -18
rect -607 -52 -573 -20
rect -607 -122 -573 -90
rect -607 -124 -573 -122
rect -489 -20 -455 -18
rect -489 -52 -455 -20
rect -489 -122 -455 -90
rect -489 -124 -455 -122
rect -371 -20 -337 -18
rect -371 -52 -337 -20
rect -371 -122 -337 -90
rect -371 -124 -337 -122
rect -253 -20 -219 -18
rect -253 -52 -219 -20
rect -253 -122 -219 -90
rect -253 -124 -219 -122
rect -135 -20 -101 -18
rect -135 -52 -101 -20
rect -135 -122 -101 -90
rect -135 -124 -101 -122
rect -17 -20 17 -18
rect -17 -52 17 -20
rect -17 -122 17 -90
rect -17 -124 17 -122
rect 101 -20 135 -18
rect 101 -52 135 -20
rect 101 -122 135 -90
rect 101 -124 135 -122
rect 219 -20 253 -18
rect 219 -52 253 -20
rect 219 -122 253 -90
rect 219 -124 253 -122
rect 337 -20 371 -18
rect 337 -52 371 -20
rect 337 -122 371 -90
rect 337 -124 371 -122
rect 455 -20 489 -18
rect 455 -52 489 -20
rect 455 -122 489 -90
rect 455 -124 489 -122
rect 573 -20 607 -18
rect 573 -52 607 -20
rect 573 -122 607 -90
rect 573 -124 607 -122
<< metal1 >>
rect -560 101 -502 107
rect -560 67 -548 101
rect -514 67 -502 101
rect -560 61 -502 67
rect -442 101 -384 107
rect -442 67 -430 101
rect -396 67 -384 101
rect -442 61 -384 67
rect -324 101 -266 107
rect -324 67 -312 101
rect -278 67 -266 101
rect -324 61 -266 67
rect -206 101 -148 107
rect -206 67 -194 101
rect -160 67 -148 101
rect -206 61 -148 67
rect -88 101 -30 107
rect -88 67 -76 101
rect -42 67 -30 101
rect -88 61 -30 67
rect 30 101 88 107
rect 30 67 42 101
rect 76 67 88 101
rect 30 61 88 67
rect 148 101 206 107
rect 148 67 160 101
rect 194 67 206 101
rect 148 61 206 67
rect 266 101 324 107
rect 266 67 278 101
rect 312 67 324 101
rect 266 61 324 67
rect 384 101 442 107
rect 384 67 396 101
rect 430 67 442 101
rect 384 61 442 67
rect 502 101 560 107
rect 502 67 514 101
rect 548 67 560 101
rect 502 61 560 67
rect -613 -18 -567 29
rect -613 -52 -607 -18
rect -573 -52 -567 -18
rect -613 -90 -567 -52
rect -613 -124 -607 -90
rect -573 -124 -567 -90
rect -613 -171 -567 -124
rect -495 -18 -449 29
rect -495 -52 -489 -18
rect -455 -52 -449 -18
rect -495 -90 -449 -52
rect -495 -124 -489 -90
rect -455 -124 -449 -90
rect -495 -171 -449 -124
rect -377 -18 -331 29
rect -377 -52 -371 -18
rect -337 -52 -331 -18
rect -377 -90 -331 -52
rect -377 -124 -371 -90
rect -337 -124 -331 -90
rect -377 -171 -331 -124
rect -259 -18 -213 29
rect -259 -52 -253 -18
rect -219 -52 -213 -18
rect -259 -90 -213 -52
rect -259 -124 -253 -90
rect -219 -124 -213 -90
rect -259 -171 -213 -124
rect -141 -18 -95 29
rect -141 -52 -135 -18
rect -101 -52 -95 -18
rect -141 -90 -95 -52
rect -141 -124 -135 -90
rect -101 -124 -95 -90
rect -141 -171 -95 -124
rect -23 -18 23 29
rect -23 -52 -17 -18
rect 17 -52 23 -18
rect -23 -90 23 -52
rect -23 -124 -17 -90
rect 17 -124 23 -90
rect -23 -171 23 -124
rect 95 -18 141 29
rect 95 -52 101 -18
rect 135 -52 141 -18
rect 95 -90 141 -52
rect 95 -124 101 -90
rect 135 -124 141 -90
rect 95 -171 141 -124
rect 213 -18 259 29
rect 213 -52 219 -18
rect 253 -52 259 -18
rect 213 -90 259 -52
rect 213 -124 219 -90
rect 253 -124 259 -90
rect 213 -171 259 -124
rect 331 -18 377 29
rect 331 -52 337 -18
rect 371 -52 377 -18
rect 331 -90 377 -52
rect 331 -124 337 -90
rect 371 -124 377 -90
rect 331 -171 377 -124
rect 449 -18 495 29
rect 449 -52 455 -18
rect 489 -52 495 -18
rect 449 -90 495 -52
rect 449 -124 455 -90
rect 489 -124 495 -90
rect 449 -171 495 -124
rect 567 -18 613 29
rect 567 -52 573 -18
rect 607 -52 613 -18
rect 567 -90 613 -52
rect 567 -124 573 -90
rect 607 -124 613 -90
rect 567 -171 613 -124
<< properties >>
string FIXED_BBOX -704 -266 704 186
<< end >>
