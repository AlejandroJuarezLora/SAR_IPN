magic
tech sky130B
magscale 1 2
timestamp 1696285870
<< psubdiff >>
rect 842 3849 876 3969
<< locali >>
rect 842 3896 878 3932
rect 844 3874 878 3896
rect 2576 3866 2610 3932
rect 3472 3863 3506 3932
rect 4040 3809 4074 3932
rect 854 3750 986 3784
rect 2596 3756 2728 3790
rect 3494 3754 3626 3788
rect 4060 3748 4192 3782
rect 304 3662 436 3696
<< viali >>
rect 841 3932 881 3966
rect 2573 3932 2613 3966
rect 3469 3932 3509 3972
rect 4037 3932 4077 3972
<< metal1 >>
rect -43 4946 1856 4949
rect 2980 4946 4264 4950
rect -43 4921 4264 4946
rect -43 2595 -15 4921
rect 1810 4920 4264 4921
rect 1810 4918 3062 4920
rect 1006 4154 1042 4160
rect 166 4106 1964 4154
rect 2520 4120 3096 4166
rect 835 3978 887 3984
rect 464 3927 516 3933
rect 835 3920 887 3926
rect 1006 3878 1042 4106
rect 2567 3978 2619 3984
rect 2567 3920 2619 3926
rect 2770 3884 2806 4120
rect 3463 3978 3515 3984
rect 3463 3920 3515 3926
rect 3682 3886 3714 4129
rect 4031 3978 4083 3984
rect 4031 3920 4083 3926
rect 4228 3878 4260 4121
rect 4575 3978 4673 3984
rect 4627 3926 4673 3978
rect 4575 3920 4673 3926
rect 464 3869 516 3875
rect 476 3665 504 3869
rect 472 3321 508 3564
rect 645 3470 677 3636
rect 1188 3531 1220 3833
rect 2928 3606 2960 3849
rect 3834 3696 3866 3837
rect 4389 3807 4668 3839
rect 3833 3664 4670 3696
rect 2928 3574 4670 3606
rect 1188 3499 4670 3531
rect 645 3438 4668 3470
rect 204 3292 4274 3321
rect -43 2567 4296 2595
<< via1 >>
rect 835 3966 887 3978
rect 464 3875 516 3927
rect 835 3932 841 3966
rect 841 3932 881 3966
rect 881 3932 887 3966
rect 835 3926 887 3932
rect 2567 3966 2619 3978
rect 2567 3932 2573 3966
rect 2573 3932 2613 3966
rect 2613 3932 2619 3966
rect 2567 3926 2619 3932
rect 3463 3972 3515 3978
rect 3463 3932 3469 3972
rect 3469 3932 3509 3972
rect 3509 3932 3515 3972
rect 3463 3926 3515 3932
rect 4031 3972 4083 3978
rect 4031 3932 4037 3972
rect 4037 3932 4077 3972
rect 4077 3932 4083 3972
rect 4031 3926 4083 3932
rect 4575 3926 4627 3978
<< metal2 >>
rect 829 3966 835 3978
rect 476 3938 835 3966
rect 476 3927 524 3938
rect 458 3875 464 3927
rect 516 3914 524 3927
rect 829 3926 835 3938
rect 887 3966 893 3978
rect 2561 3966 2567 3978
rect 887 3938 2567 3966
rect 887 3926 893 3938
rect 2561 3926 2567 3938
rect 2619 3966 2625 3978
rect 3457 3966 3463 3978
rect 2619 3938 3463 3966
rect 2619 3926 2625 3938
rect 3457 3926 3463 3938
rect 3515 3966 3521 3978
rect 4025 3966 4031 3978
rect 3515 3938 4031 3966
rect 3515 3926 3521 3938
rect 4025 3926 4031 3938
rect 4083 3966 4089 3978
rect 4569 3966 4575 3978
rect 4083 3938 4575 3966
rect 4083 3926 4089 3938
rect 4569 3926 4575 3938
rect 4627 3926 4633 3978
rect 516 3875 522 3914
use sky130_fd_pr__nfet_01v8_lvt  sky130_fd_pr__nfet_01v8_lvt_0
timestamp 1696285444
transform 0 1 2819 -1 0 3832
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8_lvt  sky130_fd_pr__nfet_01v8_lvt_1
timestamp 1696285444
transform 0 1 4283 -1 0 3826
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8_lvt  sky130_fd_pr__nfet_01v8_lvt_2
timestamp 1696285444
transform 0 1 527 1 0 3618
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8_lvt  sky130_fd_pr__nfet_01v8_lvt_3
timestamp 1696285444
transform 0 1 3715 -1 0 3826
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8_lvt  sky130_fd_pr__nfet_01v8_lvt_4
timestamp 1696285444
transform 0 1 1087 -1 0 3826
box -226 -279 226 279
use trimcap  trimcap_0
timestamp 1696109480
transform 1 0 4034 0 1 2088
box 0 376 476 1324
use trimcap  trimcap_1
timestamp 1696109480
transform 1 0 4030 0 1 3698
box 0 376 476 1324
use trimcap  trimcap_2
timestamp 1696109480
transform 1 0 3454 0 1 3710
box 0 376 476 1324
use trimcap  trimcap_3
timestamp 1696109480
transform 1 0 2868 0 1 3692
box 0 376 476 1324
use trimcap  trimcap_4
timestamp 1696109480
transform 1 0 2292 0 1 3702
box 0 376 476 1324
use trimcap  trimcap_5
timestamp 1696109480
transform 1 0 1714 0 1 3674
box 0 376 476 1324
use trimcap  trimcap_6
timestamp 1696109480
transform 1 0 1140 0 1 3674
box 0 376 476 1324
use trimcap  trimcap_7
timestamp 1696109480
transform 1 0 554 0 1 3672
box 0 376 476 1324
use trimcap  trimcap_8
timestamp 1696109480
transform 1 0 -30 0 1 3668
box 0 376 476 1324
use trimcap  trimcap_9
timestamp 1696109480
transform 1 0 -24 0 1 2092
box 0 376 476 1324
use trimcap  trimcap_10
timestamp 1696109480
transform 1 0 549 0 1 2092
box 0 376 476 1324
use trimcap  trimcap_11
timestamp 1696109480
transform 1 0 1126 0 1 2092
box 0 376 476 1324
use trimcap  trimcap_12
timestamp 1696109480
transform 1 0 1695 0 1 2096
box 0 376 476 1324
use trimcap  trimcap_13
timestamp 1696109480
transform 1 0 2288 0 1 2092
box 0 376 476 1324
use trimcap  trimcap_14
timestamp 1696109480
transform 1 0 2868 0 1 2092
box 0 376 476 1324
use trimcap  trimcap_15
timestamp 1696109480
transform 1 0 3453 0 1 2092
box 0 376 476 1324
<< labels >>
flabel metal1 -43 2567 -15 4949 0 FreeSans 480 0 0 0 DRAIN
port 0 nsew
flabel metal1 4627 3920 4673 3984 0 FreeSans 480 0 0 0 VSS
port 1 nsew
flabel metal1 4661 3820 4661 3820 0 FreeSans 480 0 0 0 d0
port 2 nsew
flabel metal1 4664 3679 4664 3679 0 FreeSans 480 0 0 0 d1
port 3 nsew
flabel metal1 4664 3587 4664 3587 0 FreeSans 480 0 0 0 d2
port 4 nsew
flabel metal1 4662 3511 4662 3511 0 FreeSans 480 0 0 0 d3
port 5 nsew
flabel metal1 4664 3453 4664 3453 0 FreeSans 480 0 0 0 d4
port 6 nsew
<< end >>
