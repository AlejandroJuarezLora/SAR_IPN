* NGSPICE file created from DAC_temp.ext - technology: sky130B

.subckt DAC_temp enb en_buf ctl1 ctl0 dum ctl3 ctl4 ctl5 ctl6 ctl7 ctl2 vin out vss
+ vdd sample
X0 vdd.t109 sample.t0 a_44621_2120.t5 vdd.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 vdd.t60 vss.t164 vdd.t59 vdd.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2 out.t80 m2_30325_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 vdd.t63 vss.t165 vdd.t62 vdd.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4 out.t81 m2_34225_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 out.t82 m2_38125_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 out.t83 carray_0.n6.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 out.t84 carray_0.n5.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 out.t32 a_45464_6355# vin.t34 vss.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X9 vdd.t107 sample.t1 enb.t15 vdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 vdd ctl1.t0 carray_0.n1.t5 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 out.t42 a_45464_2123# vin.t46 vss.t62 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X12 vss.t117 sample.t2 enb vss.t116 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 out.t85 m2_43325_6030# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 out.t86 carray_0.n5.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 out.t87 carray_0.n7.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 out.t88 carray_0.n7.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 a_44621_6352.t7 sample.t3 vdd.t105 vdd.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X18 out.t76 a_44621_2120.t8 vin.t76 vdd.t135 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X19 vdd ctl4.t0 carray_0.n4.t3 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 a_44621_2120.t1 sample.t4 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X21 en_buf.t15 enb.t16 vdd.t163 vdd.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 out.t89 m2_43325_6870# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 out.t90 carray_0.n7.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 out.t91 carray_0.n5.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 out.t92 carray_0.n7.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 out.t93 carray_0.n6.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 out.t94 carray_0.n7.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 out.t95 carray_0.n4.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 out.t96 carray_0.n7.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 out.t97 m2_43325_7710# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 out.t98 carray_0.n7.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 out.t99 carray_0.n5.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 out.t100 carray_0.n7.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 out.t101 carray_0.n6.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 out.t102 carray_0.n7.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 out.t103 carray_0.n7.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 out.t104 carray_0.n4.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 out.t7 en_buf vin.t13 vss.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X39 out.t105 carray_0.n6.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 out.t33 a_45464_6355# vin.t33 vss.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X41 out.t106 m2_3025_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 out.t107 m2_6925_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 out.t108 carray_0.n5.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 vdd.t5 enb.t17 en_buf.t14 vdd.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X45 vin.t58 enb out.t52 vdd.t56 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X46 out.t109 carray_0.n4.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 out.t110 m2_40725_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 out.t111 carray_0.n6.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 vss.t31 ctl2.t0 carray_0.n2.t5 vss.t30 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X50 out.t112 carray_0.n6.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 out.t113 carray_0.n6.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 out.t114 carray_0.n5.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X53 vin.t47 a_44621_6352.t8 out.t47 vdd.t38 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X54 en_buf enb vss.t71 vss.t70 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X55 out.t115 carray_0.n6.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 out.t116 carray_0.n6.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 out.t117 carray_0.n6.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 vss.t28 ctl5.t0 carray_0.n5.t2 vss.t27 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X59 vss.t154 a_44621_2120.t9 a_45464_2123# vss.t153 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X60 out.t118 m2_21225_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 out.t119 m2_25125_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 out.t120 m2_29025_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 out.t121 carray_0.n6.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 enb sample.t5 vss.t115 vss.t114 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X65 out.t122 m2_43325_8550# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 out.t123 carray_0.n5.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 out.t124 carray_0.n7.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 out.t125 carray_0.n7.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 out.t126 carray_0.n7.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 out.t127 carray_0.n7.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 out.t128 carray_0.n3.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 out.t129 carray_0.n7.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 out.t130 carray_0.n7.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 out.t131 carray_0.n7.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 vss.t69 enb en_buf vss.t68 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X76 out.t132 m2_43325_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 vss.t146 vdd.t164 vss.t145 vss.t144 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X78 out.t133 carray_0.n7.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 out.t134 m2_10825_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 out.t135 carray_0.n7.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 out.t136 m2_18625_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 out.t137 m2_14725_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 out.t138 carray_0.n3.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 out.t139 carray_0.n7.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 out.t140 carray_0.n7.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 out.t141 carray_0.n7.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 out.t142 carray_0.n4.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 carray_0.n5.t35 ctl5.t1 vss.t79 vss.t78 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X89 out.t143 carray_0.n7.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 vss.t113 sample.t6 enb.t5 vss.t112 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X91 out.t144 carray_0.n7.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 vss.t111 sample.t7 enb vss.t110 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X93 out.t145 carray_0.n7.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 out.t146 m2_19925_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 out.t147 carray_0.n5.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 out.t148 carray_0.n4.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 out.t5 en_buf vin.t12 vss.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X98 enb.t3 sample.t8 vss.t109 vss.t108 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X99 out.t149 carray_0.n6.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 out.t150 carray_0.n6.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 vin.t48 en_buf.t16 out.t48 vss.t63 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X102 vss.t158 dum.t0 carray_0.ndum.t1 vss.t157 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X103 vss.t73 ctl1.t1 carray_0.n1.t3 vss.t72 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X104 out.t151 carray_0.n5.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 out.t152 carray_0.n4.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 out.t65 enb.t18 vin.t65 vdd.t112 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X107 out.t153 carray_0.n6.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 vin.t63 enb.t19 out.t63 vdd.t75 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X109 out.t154 carray_0.n6.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 out.t155 carray_0.n6.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 out.t156 carray_0.n5.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 vin.t57 enb out.t55 vdd.t55 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X113 vss.t1 ctl4.t1 carray_0.n4.t1 vss.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X114 vin.t19 a_44621_6352.t9 out.t19 vdd.t27 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X115 out.t157 carray_0.n4.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 out.t158 carray_0.n5.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 out.t159 carray_0.n6.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 out.t160 carray_0.n5.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 out.t161 carray_0.n2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 out.t162 carray_0.n7.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 vss.t52 ctl0.t0 carray_0.n0.t2 vss.t51 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X122 vdd.t101 sample.t9 enb vdd.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X123 out.t163 carray_0.n7.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 vss.t143 vdd.t165 vss.t142 vss.t141 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X125 vss.t140 vdd.t166 vss.t139 vss.t138 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X126 carray_0.ndum.t0 dum.t1 vss.t81 vss.t80 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X127 out.t164 carray_0.n5.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 out.t165 carray_0.n7.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 out.t166 carray_0.n7.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 out.t4 en_buf vin.t11 vss.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X131 out.t167 carray_0.n1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 out.t168 carray_0.n7.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 out.t169 carray_0.n7.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 out.t170 carray_0.n7.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 vin.t17 en_buf.t17 out.t17 vss.t22 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X136 en_buf.t5 enb.t20 vss.t122 vss.t121 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X137 vin.t10 en_buf out.t13 vss.t11 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X138 en_buf enb vss.t67 vss.t66 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X139 out.t171 m2_5625_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 out.t172 m2_1725_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 out.t14 enb.t21 vin.t14 vdd.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X142 out.t56 enb vin.t56 vdd.t54 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X143 out.t173 m2_9525_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 out.t174 m2_30325_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 out.t175 m2_34225_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 out.t176 m2_38125_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 out.t177 carray_0.n5.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 out.t178 carray_0.n4.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 out.t179 carray_0.n7.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 out.t180 carray_0.n7.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 out.t181 carray_0.n7.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 out.t3 en_buf.t18 vin.t3 vss.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X153 out.t182 m2_27725_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 out.t183 m2_23825_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 out.t184 carray_0.n7.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 out.t185 carray_0.n7.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 out.t186 carray_0.n7.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 vin.t20 enb.t22 out.t20 vdd.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X159 out.t187 carray_0.n5.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 vin.t55 enb out.t51 vdd.t53 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X161 en_buf enb vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X162 carray_0.n0.t4 ctl0.t1 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X163 vdd.t134 a_44621_2120.t10 a_45464_2123# vdd.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X164 out.t188 m2_32925_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 out.t189 carray_0.n6.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 enb sample.t10 vdd.t99 vdd.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X167 out.t190 carray_0.n6.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 out.t41 a_45464_2123# vin.t45 vss.t61 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X169 vin.t32 a_45464_6355# out.t29 vss.t43 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X170 out.t191 carray_0.n7.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 vdd.t50 enb en_buf vdd.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X172 vin.t18 en_buf.t19 out.t18 vss.t23 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X173 out.t192 carray_0.n6.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 out.t193 carray_0.n7.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 out.t77 a_44621_6352.t10 vin.t77 vdd.t136 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X176 out.t194 carray_0.n6.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 vin.t75 a_44621_2120.t11 out.t72 vdd.t132 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X178 out.t195 carray_0.n7.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 vin.t54 enb out.t53 vdd.t48 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X180 out.t196 carray_0.n6.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 out.t197 carray_0.n7.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 out.t198 carray_0.n7.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 out.t21 enb.t23 vin.t21 vdd.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X184 out.t199 carray_0.n7.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 vdd.t97 sample.t11 enb.t12 vdd.t96 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X186 vdd.t95 sample.t12 enb vdd.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X187 out.t200 carray_0.n7.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 vdd ctl7.t0 carray_0.n7.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X189 out.t201 carray_0.n7.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 out.t202 carray_0.n7.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 out.t203 carray_0.n6.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 carray_0.n1.t4 ctl1.t2 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X193 enb.t10 sample.t13 vdd.t93 vdd.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X194 out.t204 carray_0.n7.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 out.t205 carray_0.n7.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 out.t206 carray_0.n7.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 vdd ctl3.t0 carray_0.n3.t9 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X198 out.t8 en_buf vin.t9 vss.t10 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X199 carray_0.n4.t2 ctl4.t2 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X200 vss.t107 sample.t14 a_44621_2120.t4 vss.t106 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X201 out.t207 m2_43325_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 vdd.t153 vss.t166 vdd.t152 vdd.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X203 out.t208 m2_10825_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 out.t75 a_44621_2120.t12 vin.t74 vdd.t131 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X205 out.t209 m2_14725_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 out.t210 m2_18625_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 carray_0.n7.t1 ctl7.t1 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X208 out.t211 carray_0.n6.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 out.t212 m2_43325_2670# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 out.t213 carray_0.n5.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 out.t214 carray_0.n7.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 out.t215 carray_0.n7.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 vss.t16 a_44621_6352.t11 a_45464_6355# vss.t15 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X214 out.t216 m2_19925_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 out.t217 m2_36825_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 out.t218 m2_43325_3510# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 en_buf.t11 enb.t24 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X218 vin.t31 a_45464_6355# out.t25 vss.t42 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X219 out.t219 carray_0.n5.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 out.t220 carray_0.n7.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 out.t221 carray_0.n7.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 en_buf enb vdd.t47 vdd.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X223 out.t222 carray_0.n7.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 vin.t44 a_45464_2123# out.t37 vss.t60 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X225 out.t223 carray_0.n7.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X226 out.t224 carray_0.n7.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 out.t34 a_45464_6355# vin.t30 vss.t41 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X228 out.t39 a_45464_2123# vin.t43 vss.t59 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X229 out.t225 carray_0.n4.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 out.t226 carray_0.n7.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 out.t227 carray_0.n6.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 vin.t73 a_44621_2120.t13 out.t74 vdd.t130 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X233 out.t228 m2_42025_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 out.t229 carray_0.n7.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X235 out.t230 m2_17325_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 out.t231 m2_13425_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 out.t1 a_44621_6352.t12 vin.t1 vdd.t3 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X238 out.t232 carray_0.n4.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 out.t233 carray_0.n7.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 out.t15 enb.t25 vin.t15 vdd.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X241 a_45464_6355# a_44621_6352.t13 vss.t50 vss.t49 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X242 a_45464_2123# a_44621_2120.t14 vss.t152 vss.t151 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X243 out.t234 carray_0.n7.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 out.t235 carray_0.n7.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 out.t236 carray_0.n1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 out.t237 carray_0.n6.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 a_44621_6352.t3 sample.t15 vss.t105 vss.t104 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X248 vin.t29 a_45464_6355# out.t28 vss.t40 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X249 out.t238 carray_0.n6.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 out.t239 carray_0.n2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 vin.t42 a_45464_2123# out.t46 vss.t58 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X252 out.t240 m2_43325_4350# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 vss.t101 sample.t16 a_44621_6352.t2 vss.t100 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X254 out.t241 carray_0.n5.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 out.t242 m2_1725_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 out.t243 m2_5625_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 out.t244 carray_0.n7.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 out.t245 carray_0.n7.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 out.t246 m2_9525_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 vin.t72 a_44621_2120.t15 out.t71 vdd.t129 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X261 out.t247 carray_0.n6.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 out.t248 carray_0.n3.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 enb.t2 sample.t17 vss.t103 vss.t102 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X264 enb sample.t18 vss.t99 vss.t98 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X265 out.t249 m2_43325_5190# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 out.t250 carray_0.n7.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 out.t251 carray_0.n5.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 out.t252 m2_425_6030# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 out.t253 carray_0.n7.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 out.t254 carray_0.n7.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 out.t255 carray_0.n7.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 out.t256 carray_0.n7.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 out.t257 carray_0.n4.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 vss.t77 ctl7.t2 carray_0.n7.t131 vss.t76 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X275 out.t258 carray_0.n7.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 out.t259 m2_425_6870# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 out.t260 carray_0.n7.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 carray_0.n1.t2 ctl1.t3 vss.t83 vss.t82 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X279 out.t261 carray_0.n7.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 out.t262 carray_0.n4.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 out.t263 carray_0.n7.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X282 out.t264 carray_0.n7.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 out.t40 a_45464_2123# vin.t41 vss.t57 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X284 vss.t160 ctl3.t1 carray_0.n3.t10 vss.t159 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X285 out.t265 m2_23825_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 out.t266 m2_27725_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 out.t267 m2_425_7710# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 carray_0.n4.t0 ctl4.t3 vss.t162 vss.t161 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X289 out.t268 m2_4325_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 out.t36 a_44621_6352.t14 vin.t36 vdd.t37 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X291 out.t67 a_44621_2120.t16 vin.t71 vdd.t128 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X292 out.t269 m2_8225_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 out.t270 carray_0.n4.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 out.t271 carray_0.n5.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 vss.t47 a_44621_6352.t15 a_45464_6355# vss.t46 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X296 out.t272 m2_32925_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 carray_0.n0.t1 ctl0.t2 vss.t25 vss.t24 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X298 carray_0.n7.t130 ctl7.t3 vss.t75 vss.t74 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X299 out.t273 carray_0.n4.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 out.t274 carray_0.n5.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 out.t275 carray_0.n3.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 out.t276 carray_0.n6.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 out.t277 carray_0.n5.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 vdd.t91 sample.t19 a_44621_2120.t2 vdd.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X305 vin.t8 en_buf out.t12 vss.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X306 out.t278 m2_22525_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 out.t279 m2_26425_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 out.t280 carray_0.n5.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 vdd.t156 vss.t167 vdd.t155 vdd.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X310 out.t281 carray_0.n7.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 out.t282 carray_0.n7.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 vin.t28 a_45464_6355# out.t27 vss.t39 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X313 a_45464_6355# a_44621_6352.t16 vss.t4 vss.t3 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X314 out.t283 carray_0.n7.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 out.t58 enb vin.t53 vdd.t45 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X316 out.t78 a_44621_6352.t17 vin.t78 vdd.t159 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X317 out.t284 m2_425_8550# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 vdd.t73 a_44621_6352.t18 a_45464_6355# vdd.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X319 out.t285 carray_0.n7.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 out.t286 carray_0.n7.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 out.t287 carray_0.n6.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 out.t288 carray_0.n7.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 out.t289 carray_0.n7.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 out.t290 carray_0.n7.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 vss.t137 vdd.t167 vss.t136 vss.t135 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X326 out.t291 m2_425_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 out.t292 carray_0.n7.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 out.t293 carray_0.n6.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 out.t294 carray_0.n7.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 out.t295 carray_0.n4.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 out.t296 carray_0.n5.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 out.t297 carray_0.n6.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 out.t298 carray_0.n5.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 vdd ctl6.t0 carray_0.n6.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X335 out.t299 carray_0.n7.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 out.t300 carray_0.n6.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 out.t301 carray_0.n7.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 a_45464_6355# a_44621_6352.t19 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X339 out.t302 carray_0.n5.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 out.t303 carray_0.n4.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 a_45464_2123# a_44621_2120.t17 vdd.t127 vdd.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X342 out.t304 carray_0.n5.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 out.t305 carray_0.n6.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 out.t306 carray_0.n5.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 vdd.t139 vss.t168 vdd.t138 vdd.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X346 vdd.t142 vss.t169 vdd.t141 vdd.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X347 out.t307 carray_0.n5.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X348 out.t308 carray_0.n6.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 out.t309 carray_0.n5.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 a_44621_6352.t6 sample.t20 vdd.t89 vdd.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X351 out.t310 m2_36825_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 out.t79 en_buf.t20 vin.t79 vss.t163 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X353 vdd.t87 sample.t21 a_44621_6352.t5 vdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X354 vin.t24 en_buf.t21 out.t24 vss.t29 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X355 vin.t7 en_buf out.t6 vss.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X356 out.t311 carray_0.n6.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 vin.t27 a_45464_6355# out.t31 vss.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X358 out.t312 m2_42025_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 enb.t9 sample.t22 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X360 out.t49 enb vin.t52 vdd.t44 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X361 out.t313 m2_13425_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 enb sample.t23 vdd.t83 vdd.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X363 out.t314 m2_17325_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 vin.t22 enb.t26 out.t22 vdd.t30 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X365 out.t315 carray_0.n6.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 out.t316 carray_0.n6.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 out.t317 carray_0.n7.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 out.t318 carray_0.n7.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 out.t319 carray_0.n7.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 out.t320 carray_0.n7.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 out.t321 carray_0.n6.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 carray_0.n3.t11 ctl3.t2 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X373 out.t322 m2_31625_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 out.t323 m2_39425_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 out.t324 m2_35525_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 out.t325 carray_0.n7.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 a_44621_2120.t0 sample.t24 vss.t97 vss.t96 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X378 out.t326 carray_0.n7.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 out.t327 carray_0.n6.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X380 out.t328 carray_0.n6.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 out.t329 carray_0.n6.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 out.t330 carray_0.n6.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 out.t331 carray_0.n5.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 carray_0.n6.t0 ctl6.t1 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X385 out.t35 en_buf.t22 vin.t35 vss.t48 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X386 out.t11 en_buf vin.t6 vss.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X387 out.t332 carray_0.n6.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 vdd.t36 a_44621_6352.t20 a_45464_6355# vdd.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X389 out.t333 carray_0.n6.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 out.t334 m2_12125_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 carray_0.n2.t7 ctl2.t1 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X392 out.t335 carray_0.n6.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 out.t336 m2_16025_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 vdd.t68 vss.t170 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X395 out.t50 enb vin.t51 vdd.t43 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X396 vin.t59 enb.t27 out.t59 vdd.t57 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X397 vin.t50 enb out.t54 vdd.t42 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X398 out.t337 carray_0.n6.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 out.t338 carray_0.n6.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 out.t339 carray_0.n6.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 out.t340 carray_0.n6.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 out.t341 carray_0.n0.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 vss.t18 enb.t28 en_buf.t3 vss.t17 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X404 out.t342 carray_0.n7.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 out.t343 carray_0.n7.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 vss.t65 enb en_buf vss.t64 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X407 out.t344 carray_0.n6.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 vin.t23 en_buf.t23 out.t23 vss.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X409 vin.t5 en_buf out.t10 vss.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X410 a_45464_6355# a_44621_6352.t21 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X411 out.t345 carray_0.n6.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X412 out.t346 carray_0.n2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 out.t347 carray_0.n7.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 out.t348 carray_0.n7.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 a_45464_2123# a_44621_2120.t18 vss.t150 vss.t149 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X416 out.t349 carray_0.n7.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 out.t350 m2_4325_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 out.t351 carray_0.n7.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 vss.t35 ctl6.t2 carray_0.n6.t2 vss.t34 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X420 out.t352 m2_8225_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 out.t353 carray_0.n6.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 vss.t148 a_44621_2120.t19 a_45464_2123# vss.t147 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X423 out.t354 carray_0.n7.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 out.t355 carray_0.n3.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 out.t2 enb.t29 vin.t2 vdd.t6 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X426 out.t356 carray_0.n7.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 vss.t134 vdd.t168 vss.t133 vss.t132 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X428 out.t357 carray_0.n7.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 out.t358 carray_0.n7.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 out.t359 carray_0.n7.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 out.t360 carray_0.n7.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 out.t361 carray_0.n6.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 vss.t95 sample.t25 a_44621_6352.t1 vss.t94 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X434 vss.t93 sample.t26 a_44621_2120.t7 vss.t92 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X435 out.t362 carray_0.n7.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 out.t363 carray_0.n7.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 out.t364 carray_0.n6.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 out.t365 carray_0.n6.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 out.t30 a_45464_6355# vin.t26 vss.t37 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X440 out.t366 m2_22525_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 out.t367 m2_26425_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 vin.t40 a_45464_2123# out.t38 vss.t56 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X443 vin.t4 en_buf out.t9 vss.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X444 out.t368 carray_0.n6.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 out.t369 m2_6925_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 out.t370 m2_3025_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 out.t64 en_buf.t24 vin.t64 vss.t120 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X448 out.t69 a_44621_2120.t20 vin.t70 vdd.t125 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X449 vss.t91 sample.t27 enb.t0 vss.t90 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X450 out.t371 carray_0.n3.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 out.t372 carray_0.n6.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 vin.t0 a_44621_6352.t22 out.t0 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X453 vin.t66 enb.t30 out.t66 vdd.t117 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X454 out.t373 m2_40725_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 a_44621_6352.t0 sample.t28 vss.t89 vss.t88 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X456 a_44621_2120.t6 sample.t29 vss.t87 vss.t86 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X457 out.t374 carray_0.n3.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 out.t375 carray_0.n6.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 out.t376 carray_0.n3.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 en_buf.t1 enb.t31 vss.t85 vss.t84 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X461 out.t377 carray_0.n7.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 out.t378 m2_425_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 out.t379 carray_0.n7.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 carray_0.n3.t0 ctl3.t3 vss.t20 vss.t19 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X465 vss.t131 vdd.t169 vss.t130 vss.t129 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X466 vss.t128 vdd.t170 vss.t127 vss.t126 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X467 out.t380 m2_21225_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 out.t381 m2_29025_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 out.t382 m2_25125_9390# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 out.t383 m2_425_2670# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 out.t45 a_45464_2123# vin.t39 vss.t55 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X472 out.t384 carray_0.n7.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 out.t385 carray_0.n7.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 carray_0.n6.t67 ctl6.t3 vss.t156 vss.t155 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X475 out.t57 enb vin.t49 vdd.t41 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X476 out.t386 m2_425_3510# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 carray_0.n2.t4 ctl2.t2 vss.t33 vss.t32 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X478 out.t387 carray_0.n7.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 out.t388 carray_0.n7.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 vss.t119 enb.t32 en_buf.t0 vss.t118 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X481 out.t389 carray_0.n7.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 out.t390 carray_0.n7.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 out.t391 carray_0.n7.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 a_44621_2120.t3 sample.t30 vdd.t81 vdd.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X485 out.t392 carray_0.n7.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 out.t393 carray_0.n7.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 out.t394 carray_0.n7.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 out.t395 carray_0.n2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 out.t396 carray_0.n6.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 vdd dum.t2 carray_0.ndum.t3 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X491 vin.t38 a_45464_2123# out.t44 vss.t54 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X492 out.t397 carray_0.n7.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 out.t26 a_45464_6355# vin.t25 vss.t36 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X494 out.t398 carray_0.n7.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 out.t399 carray_0.n7.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 out.t16 en_buf.t25 vin.t16 vss.t21 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X497 vdd.t71 vss.t171 vdd.t70 vdd.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X498 out.t400 carray_0.ndum.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 out.t401 carray_0.n6.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 vin.t62 a_44621_6352.t23 out.t62 vdd.t74 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X501 vin.t69 a_44621_2120.t21 out.t68 vdd.t124 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X502 vdd ctl2.t3 carray_0.n2.t6 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X503 out.t60 a_44621_6352.t24 vin.t60 vdd.t64 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X504 out.t70 a_44621_2120.t22 vin.t68 vdd.t123 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X505 vdd.t77 enb.t33 en_buf.t9 vdd.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X506 vdd.t40 enb en_buf vdd.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X507 vss.t125 vdd.t171 vss.t124 vss.t123 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X508 vdd ctl0.t3 carray_0.n0.t3 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X509 out.t402 m2_425_4350# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 vdd ctl5.t2 carray_0.n5.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X511 out.t403 m2_31625_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 out.t404 m2_35525_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 out.t405 m2_39425_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 carray_0.ndum.t2 dum.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X515 a_45464_2123# a_44621_2120.t23 vdd.t122 vdd.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X516 out.t406 m2_425_5190# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 out.t407 carray_0.n6.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 out.t408 carray_0.n7.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 out.t409 carray_0.n7.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 vdd.t120 a_44621_2120.t24 a_45464_2123# vdd.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X521 vin.t37 a_45464_2123# out.t43 vss.t53 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X522 out.t410 m2_12125_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 out.t411 m2_16025_1830# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 out.t412 carray_0.n6.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 out.t413 carray_0.n7.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 out.t414 carray_0.n7.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 out.t415 carray_0.n7.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 out.t416 carray_0.n7.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 vin.t61 a_44621_6352.t25 out.t61 vdd.t65 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X530 vin.t67 a_44621_2120.t25 out.t73 vdd.t118 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X531 out.t417 carray_0.n7.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 carray_0.n5.t1 ctl5.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X533 out.t418 carray_0.n6.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 vdd.t79 sample.t31 a_44621_6352.t4 vdd.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X535 out.t419 carray_0.n5.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 sample.n20 sample.t4 212.081
R1 sample.n26 sample.t0 212.081
R2 sample.n24 sample.t30 212.081
R3 sample.n22 sample.t19 212.081
R4 sample.n10 sample.t23 212.081
R5 sample.n16 sample.t12 212.081
R6 sample.n14 sample.t10 212.081
R7 sample.n12 sample.t9 212.081
R8 sample.n0 sample.t3 212.081
R9 sample.n6 sample.t31 212.081
R10 sample.n4 sample.t20 212.081
R11 sample.n2 sample.t21 212.081
R12 sample.n35 sample.t22 212.081
R13 sample.n33 sample.t11 212.081
R14 sample.n38 sample.t13 212.081
R15 sample.n36 sample.t1 212.081
R16 sample.n20 sample.t29 139.78
R17 sample.n26 sample.t26 139.78
R18 sample.n24 sample.t24 139.78
R19 sample.n22 sample.t14 139.78
R20 sample.n10 sample.t18 139.78
R21 sample.n16 sample.t7 139.78
R22 sample.n14 sample.t5 139.78
R23 sample.n12 sample.t2 139.78
R24 sample.n0 sample.t28 139.78
R25 sample.n6 sample.t25 139.78
R26 sample.n4 sample.t15 139.78
R27 sample.n2 sample.t16 139.78
R28 sample.n35 sample.t17 139.78
R29 sample.n33 sample.t6 139.78
R30 sample.n38 sample.t8 139.78
R31 sample.n36 sample.t27 139.78
R32 sample.n23 sample.n21 97.5045
R33 sample.n13 sample.n11 97.5045
R34 sample.n3 sample.n1 97.5045
R35 sample.n40 sample.n37 97.5045
R36 sample.n28 sample.n27 76.0005
R37 sample.n25 sample.n21 76.0005
R38 sample.n18 sample.n17 76.0005
R39 sample.n15 sample.n11 76.0005
R40 sample.n8 sample.n7 76.0005
R41 sample.n5 sample.n1 76.0005
R42 sample.n40 sample.n39 76.0005
R43 sample.n29 sample.n20 44.4802
R44 sample.n19 sample.n10 44.4802
R45 sample.n9 sample.n0 44.4802
R46 sample.n42 sample.n35 44.4802
R47 sample.n30 sample 33.6245
R48 sample.n23 sample.n22 30.6732
R49 sample.n24 sample.n23 30.6732
R50 sample.n25 sample.n24 30.6732
R51 sample.n26 sample.n25 30.6732
R52 sample.n27 sample.n26 30.6732
R53 sample.n27 sample.n20 30.6732
R54 sample.n13 sample.n12 30.6732
R55 sample.n14 sample.n13 30.6732
R56 sample.n15 sample.n14 30.6732
R57 sample.n16 sample.n15 30.6732
R58 sample.n17 sample.n16 30.6732
R59 sample.n17 sample.n10 30.6732
R60 sample.n3 sample.n2 30.6732
R61 sample.n4 sample.n3 30.6732
R62 sample.n5 sample.n4 30.6732
R63 sample.n6 sample.n5 30.6732
R64 sample.n7 sample.n6 30.6732
R65 sample.n7 sample.n0 30.6732
R66 sample.n37 sample.n36 30.6732
R67 sample.n39 sample.n38 30.6732
R68 sample.n34 sample.n33 30.6732
R69 sample.n35 sample.n34 30.6732
R70 sample.n29 sample.n28 23.9042
R71 sample.n19 sample.n18 23.9042
R72 sample.n9 sample.n8 23.9042
R73 sample.n42 sample.n41 23.9042
R74 sample.n28 sample.n21 21.5045
R75 sample.n18 sample.n11 21.5045
R76 sample.n8 sample.n1 21.5045
R77 sample.n41 sample.n40 21.5045
R78 sample sample.n29 5.38578
R79 sample sample.n19 5.38578
R80 sample sample.n9 5.38578
R81 sample sample.n42 5.38445
R82 sample sample.n32 3.3673
R83 sample.n32 sample.n31 3.30675
R84 sample.n31 sample.n30 3.30675
R85 sample.n30 sample 0.0610469
R86 sample.n31 sample 0.0610469
R87 sample.n32 sample 0.0610469
R88 a_44621_2120.n11 a_44621_2120.t23 212.081
R89 a_44621_2120.n9 a_44621_2120.t24 212.081
R90 a_44621_2120.n5 a_44621_2120.t17 212.081
R91 a_44621_2120.n3 a_44621_2120.t10 212.081
R92 a_44621_2120.n26 a_44621_2120.n25 146.423
R93 a_44621_2120.n2 a_44621_2120.n0 144.089
R94 a_44621_2120.n13 a_44621_2120.t16 143.071
R95 a_44621_2120.n21 a_44621_2120.t11 142.75
R96 a_44621_2120.n13 a_44621_2120.t21 142.75
R97 a_44621_2120.n14 a_44621_2120.t8 142.75
R98 a_44621_2120.n15 a_44621_2120.t13 142.75
R99 a_44621_2120.n16 a_44621_2120.t20 142.75
R100 a_44621_2120.n17 a_44621_2120.t25 142.75
R101 a_44621_2120.n18 a_44621_2120.t12 142.75
R102 a_44621_2120.n19 a_44621_2120.t15 142.75
R103 a_44621_2120.n20 a_44621_2120.t22 142.75
R104 a_44621_2120.n11 a_44621_2120.t18 139.78
R105 a_44621_2120.n9 a_44621_2120.t19 139.78
R106 a_44621_2120.n5 a_44621_2120.t14 139.78
R107 a_44621_2120.n3 a_44621_2120.t9 139.78
R108 a_44621_2120.n2 a_44621_2120.n1 107.822
R109 a_44621_2120.n25 a_44621_2120.n24 107.249
R110 a_44621_2120.n7 a_44621_2120.n4 97.5045
R111 a_44621_2120.n7 a_44621_2120.n6 76.0005
R112 a_44621_2120.n23 a_44621_2120.n2 46.6252
R113 a_44621_2120.n12 a_44621_2120.n11 39.8685
R114 a_44621_2120.n4 a_44621_2120.n3 30.6732
R115 a_44621_2120.n6 a_44621_2120.n5 30.6732
R116 a_44621_2120.n10 a_44621_2120.n9 30.6732
R117 a_44621_2120.n11 a_44621_2120.n10 30.6732
R118 a_44621_2120.n24 a_44621_2120.t2 26.5955
R119 a_44621_2120.n24 a_44621_2120.t3 26.5955
R120 a_44621_2120.n26 a_44621_2120.t5 26.5955
R121 a_44621_2120.t1 a_44621_2120.n26 26.5955
R122 a_44621_2120.n0 a_44621_2120.t7 24.9236
R123 a_44621_2120.n0 a_44621_2120.t6 24.9236
R124 a_44621_2120.n1 a_44621_2120.t4 24.9236
R125 a_44621_2120.n1 a_44621_2120.t0 24.9236
R126 a_44621_2120.n8 a_44621_2120.n7 21.5045
R127 a_44621_2120.n12 a_44621_2120.n8 19.201
R128 a_44621_2120.n25 a_44621_2120.n23 14.3512
R129 a_44621_2120.n22 a_44621_2120.n21 9.01046
R130 a_44621_2120.n23 a_44621_2120.n22 4.58256
R131 a_44621_2120.n22 a_44621_2120.n12 1.91581
R132 a_44621_2120.n21 a_44621_2120.n20 0.321152
R133 a_44621_2120.n20 a_44621_2120.n19 0.321152
R134 a_44621_2120.n19 a_44621_2120.n18 0.321152
R135 a_44621_2120.n18 a_44621_2120.n17 0.321152
R136 a_44621_2120.n17 a_44621_2120.n16 0.321152
R137 a_44621_2120.n16 a_44621_2120.n15 0.321152
R138 a_44621_2120.n15 a_44621_2120.n14 0.321152
R139 a_44621_2120.n14 a_44621_2120.n13 0.321152
R140 vdd.t66 vdd.t84 1396.88
R141 vdd.t151 vdd.t104 1396.88
R142 vdd.t69 vdd.t82 1396.88
R143 vdd.t102 vdd.t154 1396.88
R144 vdd.n432 vdd.t66 1225.23
R145 vdd.n684 vdd.t151 1225.23
R146 vdd.n745 vdd.t69 1225.23
R147 vdd.t76 vdd.t137 716.199
R148 vdd.t58 vdd.t72 716.199
R149 vdd.t140 vdd.t39 716.199
R150 vdd.t61 vdd.t133 716.199
R151 vdd.t106 vdd.t17 615.577
R152 vdd.t147 vdd.t86 615.577
R153 vdd.t46 vdd.t100 615.577
R154 vdd.t121 vdd.t90 615.577
R155 vdd.n774 vdd.t91 584.644
R156 vdd.n763 vdd.t134 584.644
R157 vdd.n713 vdd.t101 584.644
R158 vdd.n702 vdd.t40 584.644
R159 vdd.n652 vdd.t87 584.644
R160 vdd.n641 vdd.t73 584.644
R161 vdd.n598 vdd.t107 584.644
R162 vdd.n587 vdd.t77 584.644
R163 vdd.n429 vdd.t58 544.548
R164 vdd.n687 vdd.t140 544.548
R165 vdd.n748 vdd.t61 544.548
R166 vdd.t162 vdd.t76 248.599
R167 vdd.t4 vdd.t162 248.599
R168 vdd.t17 vdd.t4 248.599
R169 vdd.t92 vdd.t106 248.599
R170 vdd.t96 vdd.t92 248.599
R171 vdd.t84 vdd.t96 248.599
R172 vdd.t72 vdd.t25 248.599
R173 vdd.t25 vdd.t35 248.599
R174 vdd.t35 vdd.t147 248.599
R175 vdd.t86 vdd.t88 248.599
R176 vdd.t104 vdd.t78 248.599
R177 vdd.t39 vdd.t51 248.599
R178 vdd.t51 vdd.t49 248.599
R179 vdd.t49 vdd.t46 248.599
R180 vdd.t100 vdd.t98 248.599
R181 vdd.t82 vdd.t94 248.599
R182 vdd.t133 vdd.t126 248.599
R183 vdd.t126 vdd.t119 248.599
R184 vdd.t119 vdd.t121 248.599
R185 vdd.t90 vdd.t80 248.599
R186 vdd.t80 vdd.t108 248.599
R187 vdd.t108 vdd.t102 248.599
R188 vdd.n785 vdd.t155 242.135
R189 vdd.n806 vdd.t156 242.135
R190 vdd.n724 vdd.t70 242.135
R191 vdd.n143 vdd.t71 242.135
R192 vdd.n609 vdd.t67 242.135
R193 vdd.n438 vdd.t68 242.135
R194 vdd.n663 vdd.t152 242.135
R195 vdd.n287 vdd.t153 242.135
R196 vdd.n760 vdd.t63 234.554
R197 vdd.n755 vdd.t62 234.554
R198 vdd.n699 vdd.t142 234.554
R199 vdd.n694 vdd.t141 234.554
R200 vdd.n581 vdd.t138 234.554
R201 vdd.n638 vdd.t60 234.554
R202 vdd.n633 vdd.t59 234.554
R203 vdd.n584 vdd.t139 234.554
R204 vdd.n65 vdd.n63 210.739
R205 vdd.n209 vdd.n207 210.739
R206 vdd.n353 vdd.n351 210.739
R207 vdd.n504 vdd.n502 210.739
R208 vdd.n779 vdd.n778 180.994
R209 vdd.n768 vdd.n767 180.994
R210 vdd.n718 vdd.n717 180.994
R211 vdd.n707 vdd.n706 180.994
R212 vdd.n657 vdd.n656 180.994
R213 vdd.n646 vdd.n645 180.994
R214 vdd.n603 vdd.n602 180.994
R215 vdd.n592 vdd.n591 180.994
R216 vdd.n754 vdd.t166 166.282
R217 vdd.n693 vdd.t170 166.282
R218 vdd.n580 vdd.t169 166.282
R219 vdd.n632 vdd.t165 166.282
R220 vdd.n783 vdd.t103 151.123
R221 vdd.n772 vdd.t122 151.123
R222 vdd.n722 vdd.t83 151.123
R223 vdd.n711 vdd.t47 151.123
R224 vdd.n661 vdd.t105 151.123
R225 vdd.n650 vdd.t148 151.123
R226 vdd.n607 vdd.t85 151.123
R227 vdd.n596 vdd.t18 151.123
R228 vdd.n88 vdd.n87 92.5005
R229 vdd.n87 vdd.n86 92.5005
R230 vdd.n91 vdd.n90 92.5005
R231 vdd.n90 vdd.n89 92.5005
R232 vdd.n94 vdd.n93 92.5005
R233 vdd.n93 vdd.n92 92.5005
R234 vdd.n97 vdd.n96 92.5005
R235 vdd.n96 vdd.n95 92.5005
R236 vdd.n100 vdd.n99 92.5005
R237 vdd.n99 vdd.n98 92.5005
R238 vdd.n103 vdd.n102 92.5005
R239 vdd.n102 vdd.n101 92.5005
R240 vdd.n106 vdd.n105 92.5005
R241 vdd.n105 vdd.n104 92.5005
R242 vdd.n109 vdd.n108 92.5005
R243 vdd.n108 vdd.n107 92.5005
R244 vdd.n112 vdd.n111 92.5005
R245 vdd.n111 vdd.n110 92.5005
R246 vdd.n115 vdd.n114 92.5005
R247 vdd.n114 vdd.n113 92.5005
R248 vdd.n118 vdd.n117 92.5005
R249 vdd.n117 vdd.n116 92.5005
R250 vdd.n121 vdd.n120 92.5005
R251 vdd.n120 vdd.n119 92.5005
R252 vdd.n124 vdd.n123 92.5005
R253 vdd.n123 vdd.n122 92.5005
R254 vdd.n127 vdd.n126 92.5005
R255 vdd.n126 vdd.n125 92.5005
R256 vdd.n130 vdd.n129 92.5005
R257 vdd.n129 vdd.n128 92.5005
R258 vdd.n133 vdd.n132 92.5005
R259 vdd.n132 vdd.n131 92.5005
R260 vdd.n136 vdd.n135 92.5005
R261 vdd.n135 vdd.n134 92.5005
R262 vdd.n138 vdd.n137 92.5005
R263 vdd.n4 vdd.n3 92.5005
R264 vdd.n1 vdd.n0 92.5005
R265 vdd.n81 vdd.n80 92.5005
R266 vdd.n85 vdd.n84 92.5005
R267 vdd.n40 vdd.n39 92.5005
R268 vdd.n38 vdd.n37 92.5005
R269 vdd.n36 vdd.n35 92.5005
R270 vdd.n34 vdd.n33 92.5005
R271 vdd.n32 vdd.n31 92.5005
R272 vdd.n30 vdd.n29 92.5005
R273 vdd.n28 vdd.n27 92.5005
R274 vdd.n26 vdd.n25 92.5005
R275 vdd.n24 vdd.n23 92.5005
R276 vdd.n22 vdd.n21 92.5005
R277 vdd.n20 vdd.n19 92.5005
R278 vdd.n18 vdd.n17 92.5005
R279 vdd.n16 vdd.n15 92.5005
R280 vdd.n14 vdd.n13 92.5005
R281 vdd.n12 vdd.n11 92.5005
R282 vdd.n10 vdd.n9 92.5005
R283 vdd.n8 vdd.n7 92.5005
R284 vdd.n6 vdd.n5 92.5005
R285 vdd.n232 vdd.n231 92.5005
R286 vdd.n231 vdd.n230 92.5005
R287 vdd.n235 vdd.n234 92.5005
R288 vdd.n234 vdd.n233 92.5005
R289 vdd.n238 vdd.n237 92.5005
R290 vdd.n237 vdd.n236 92.5005
R291 vdd.n241 vdd.n240 92.5005
R292 vdd.n240 vdd.n239 92.5005
R293 vdd.n244 vdd.n243 92.5005
R294 vdd.n243 vdd.n242 92.5005
R295 vdd.n247 vdd.n246 92.5005
R296 vdd.n246 vdd.n245 92.5005
R297 vdd.n250 vdd.n249 92.5005
R298 vdd.n249 vdd.n248 92.5005
R299 vdd.n253 vdd.n252 92.5005
R300 vdd.n252 vdd.n251 92.5005
R301 vdd.n256 vdd.n255 92.5005
R302 vdd.n255 vdd.n254 92.5005
R303 vdd.n259 vdd.n258 92.5005
R304 vdd.n258 vdd.n257 92.5005
R305 vdd.n262 vdd.n261 92.5005
R306 vdd.n261 vdd.n260 92.5005
R307 vdd.n265 vdd.n264 92.5005
R308 vdd.n264 vdd.n263 92.5005
R309 vdd.n268 vdd.n267 92.5005
R310 vdd.n267 vdd.n266 92.5005
R311 vdd.n271 vdd.n270 92.5005
R312 vdd.n270 vdd.n269 92.5005
R313 vdd.n274 vdd.n273 92.5005
R314 vdd.n273 vdd.n272 92.5005
R315 vdd.n277 vdd.n276 92.5005
R316 vdd.n276 vdd.n275 92.5005
R317 vdd.n280 vdd.n279 92.5005
R318 vdd.n279 vdd.n278 92.5005
R319 vdd.n282 vdd.n281 92.5005
R320 vdd.n148 vdd.n147 92.5005
R321 vdd.n145 vdd.n144 92.5005
R322 vdd.n225 vdd.n224 92.5005
R323 vdd.n229 vdd.n228 92.5005
R324 vdd.n184 vdd.n183 92.5005
R325 vdd.n182 vdd.n181 92.5005
R326 vdd.n180 vdd.n179 92.5005
R327 vdd.n178 vdd.n177 92.5005
R328 vdd.n176 vdd.n175 92.5005
R329 vdd.n174 vdd.n173 92.5005
R330 vdd.n172 vdd.n171 92.5005
R331 vdd.n170 vdd.n169 92.5005
R332 vdd.n168 vdd.n167 92.5005
R333 vdd.n166 vdd.n165 92.5005
R334 vdd.n164 vdd.n163 92.5005
R335 vdd.n162 vdd.n161 92.5005
R336 vdd.n160 vdd.n159 92.5005
R337 vdd.n158 vdd.n157 92.5005
R338 vdd.n156 vdd.n155 92.5005
R339 vdd.n154 vdd.n153 92.5005
R340 vdd.n152 vdd.n151 92.5005
R341 vdd.n150 vdd.n149 92.5005
R342 vdd.n376 vdd.n375 92.5005
R343 vdd.n375 vdd.n374 92.5005
R344 vdd.n379 vdd.n378 92.5005
R345 vdd.n378 vdd.n377 92.5005
R346 vdd.n382 vdd.n381 92.5005
R347 vdd.n381 vdd.n380 92.5005
R348 vdd.n385 vdd.n384 92.5005
R349 vdd.n384 vdd.n383 92.5005
R350 vdd.n388 vdd.n387 92.5005
R351 vdd.n387 vdd.n386 92.5005
R352 vdd.n391 vdd.n390 92.5005
R353 vdd.n390 vdd.n389 92.5005
R354 vdd.n394 vdd.n393 92.5005
R355 vdd.n393 vdd.n392 92.5005
R356 vdd.n397 vdd.n396 92.5005
R357 vdd.n396 vdd.n395 92.5005
R358 vdd.n400 vdd.n399 92.5005
R359 vdd.n399 vdd.n398 92.5005
R360 vdd.n403 vdd.n402 92.5005
R361 vdd.n402 vdd.n401 92.5005
R362 vdd.n406 vdd.n405 92.5005
R363 vdd.n405 vdd.n404 92.5005
R364 vdd.n409 vdd.n408 92.5005
R365 vdd.n408 vdd.n407 92.5005
R366 vdd.n412 vdd.n411 92.5005
R367 vdd.n411 vdd.n410 92.5005
R368 vdd.n415 vdd.n414 92.5005
R369 vdd.n414 vdd.n413 92.5005
R370 vdd.n418 vdd.n417 92.5005
R371 vdd.n417 vdd.n416 92.5005
R372 vdd.n421 vdd.n420 92.5005
R373 vdd.n420 vdd.n419 92.5005
R374 vdd.n424 vdd.n423 92.5005
R375 vdd.n423 vdd.n422 92.5005
R376 vdd.n426 vdd.n425 92.5005
R377 vdd.n292 vdd.n291 92.5005
R378 vdd.n289 vdd.n288 92.5005
R379 vdd.n369 vdd.n368 92.5005
R380 vdd.n373 vdd.n372 92.5005
R381 vdd.n328 vdd.n327 92.5005
R382 vdd.n326 vdd.n325 92.5005
R383 vdd.n324 vdd.n323 92.5005
R384 vdd.n322 vdd.n321 92.5005
R385 vdd.n320 vdd.n319 92.5005
R386 vdd.n318 vdd.n317 92.5005
R387 vdd.n316 vdd.n315 92.5005
R388 vdd.n314 vdd.n313 92.5005
R389 vdd.n312 vdd.n311 92.5005
R390 vdd.n310 vdd.n309 92.5005
R391 vdd.n308 vdd.n307 92.5005
R392 vdd.n306 vdd.n305 92.5005
R393 vdd.n304 vdd.n303 92.5005
R394 vdd.n302 vdd.n301 92.5005
R395 vdd.n300 vdd.n299 92.5005
R396 vdd.n298 vdd.n297 92.5005
R397 vdd.n296 vdd.n295 92.5005
R398 vdd.n294 vdd.n293 92.5005
R399 vdd.n527 vdd.n526 92.5005
R400 vdd.n526 vdd.n525 92.5005
R401 vdd.n530 vdd.n529 92.5005
R402 vdd.n529 vdd.n528 92.5005
R403 vdd.n533 vdd.n532 92.5005
R404 vdd.n532 vdd.n531 92.5005
R405 vdd.n536 vdd.n535 92.5005
R406 vdd.n535 vdd.n534 92.5005
R407 vdd.n539 vdd.n538 92.5005
R408 vdd.n538 vdd.n537 92.5005
R409 vdd.n542 vdd.n541 92.5005
R410 vdd.n541 vdd.n540 92.5005
R411 vdd.n545 vdd.n544 92.5005
R412 vdd.n544 vdd.n543 92.5005
R413 vdd.n548 vdd.n547 92.5005
R414 vdd.n547 vdd.n546 92.5005
R415 vdd.n551 vdd.n550 92.5005
R416 vdd.n550 vdd.n549 92.5005
R417 vdd.n554 vdd.n553 92.5005
R418 vdd.n553 vdd.n552 92.5005
R419 vdd.n557 vdd.n556 92.5005
R420 vdd.n556 vdd.n555 92.5005
R421 vdd.n560 vdd.n559 92.5005
R422 vdd.n559 vdd.n558 92.5005
R423 vdd.n563 vdd.n562 92.5005
R424 vdd.n562 vdd.n561 92.5005
R425 vdd.n566 vdd.n565 92.5005
R426 vdd.n565 vdd.n564 92.5005
R427 vdd.n569 vdd.n568 92.5005
R428 vdd.n568 vdd.n567 92.5005
R429 vdd.n572 vdd.n571 92.5005
R430 vdd.n571 vdd.n570 92.5005
R431 vdd.n575 vdd.n574 92.5005
R432 vdd.n574 vdd.n573 92.5005
R433 vdd.n577 vdd.n576 92.5005
R434 vdd.n443 vdd.n442 92.5005
R435 vdd.n440 vdd.n439 92.5005
R436 vdd.n520 vdd.n519 92.5005
R437 vdd.n524 vdd.n523 92.5005
R438 vdd.n479 vdd.n478 92.5005
R439 vdd.n477 vdd.n476 92.5005
R440 vdd.n475 vdd.n474 92.5005
R441 vdd.n473 vdd.n472 92.5005
R442 vdd.n471 vdd.n470 92.5005
R443 vdd.n469 vdd.n468 92.5005
R444 vdd.n467 vdd.n466 92.5005
R445 vdd.n465 vdd.n464 92.5005
R446 vdd.n463 vdd.n462 92.5005
R447 vdd.n461 vdd.n460 92.5005
R448 vdd.n459 vdd.n458 92.5005
R449 vdd.n457 vdd.n456 92.5005
R450 vdd.n455 vdd.n454 92.5005
R451 vdd.n453 vdd.n452 92.5005
R452 vdd.n451 vdd.n450 92.5005
R453 vdd.n449 vdd.n448 92.5005
R454 vdd.n447 vdd.n446 92.5005
R455 vdd.n445 vdd.n444 92.5005
R456 vdd.n88 vdd.n85 89.6005
R457 vdd.n6 vdd.n4 89.6005
R458 vdd.n232 vdd.n229 89.6005
R459 vdd.n150 vdd.n148 89.6005
R460 vdd.n376 vdd.n373 89.6005
R461 vdd.n294 vdd.n292 89.6005
R462 vdd.n527 vdd.n524 89.6005
R463 vdd.n445 vdd.n443 89.6005
R464 vdd.n48 vdd.n40 85.71
R465 vdd.n192 vdd.n184 85.71
R466 vdd.n336 vdd.n328 85.71
R467 vdd.n487 vdd.n479 85.71
R468 vdd.n139 vdd.n138 83.9635
R469 vdd.n283 vdd.n282 83.9635
R470 vdd.n427 vdd.n426 83.9635
R471 vdd.n578 vdd.n577 83.9635
R472 vdd.n63 vdd.t128 78.6097
R473 vdd.n207 vdd.t41 78.6097
R474 vdd.n351 vdd.t37 78.6097
R475 vdd.n502 vdd.t112 78.6097
R476 vdd.n793 vdd.n792 76.0005
R477 vdd.n732 vdd.n731 76.0005
R478 vdd.n671 vdd.n670 76.0005
R479 vdd.n617 vdd.n616 76.0005
R480 vdd.n80 vdd.n79 72.7879
R481 vdd.n224 vdd.n223 72.7879
R482 vdd.n368 vdd.n367 72.7879
R483 vdd.n519 vdd.n518 72.7879
R484 vdd.n65 vdd.n64 68.856
R485 vdd.n209 vdd.n208 68.856
R486 vdd.n353 vdd.n352 68.856
R487 vdd.n504 vdd.n503 68.856
R488 vdd.n95 vdd.t123 65.2294
R489 vdd.n239 vdd.t45 65.2294
R490 vdd.n383 vdd.t64 65.2294
R491 vdd.n534 vdd.t29 65.2294
R492 vdd.n747 vdd.n746 60.1149
R493 vdd.n686 vdd.n685 60.1149
R494 vdd.n434 vdd.n433 60.1149
R495 vdd.n52 vdd.n51 56.4711
R496 vdd.n44 vdd.n43 56.4711
R497 vdd.n196 vdd.n195 56.4711
R498 vdd.n188 vdd.n187 56.4711
R499 vdd.n340 vdd.n339 56.4711
R500 vdd.n332 vdd.n331 56.4711
R501 vdd.n491 vdd.n490 56.4711
R502 vdd.n483 vdd.n482 56.4711
R503 vdd.n791 vdd.t168 50.5057
R504 vdd.n730 vdd.t164 50.5057
R505 vdd.n615 vdd.t171 50.5057
R506 vdd.n669 vdd.t167 50.5057
R507 vdd.n751 vdd.n750 50.2453
R508 vdd.n690 vdd.n689 50.2453
R509 vdd.n435 vdd.n431 50.2453
R510 vdd.n67 vdd.n66 49.4123
R511 vdd.n211 vdd.n210 49.4123
R512 vdd.n355 vdd.n354 49.4123
R513 vdd.n506 vdd.n505 49.4123
R514 vdd.n131 vdd.t124 48.504
R515 vdd.n275 vdd.t53 48.504
R516 vdd.n419 vdd.t74 48.504
R517 vdd.n570 vdd.t28 48.504
R518 vdd.n749 vdd.n748 46.2505
R519 vdd.n746 vdd.n745 46.2505
R520 vdd.n688 vdd.n687 46.2505
R521 vdd.n685 vdd.n684 46.2505
R522 vdd.n430 vdd.n429 46.2505
R523 vdd.n433 vdd.n432 46.2505
R524 vdd.n84 vdd.n83 42.8997
R525 vdd.n228 vdd.n227 42.8997
R526 vdd.n372 vdd.n371 42.8997
R527 vdd.n523 vdd.n522 42.8997
R528 vdd.n3 vdd.n2 42.8996
R529 vdd.n147 vdd.n146 42.8996
R530 vdd.n291 vdd.n290 42.8996
R531 vdd.n442 vdd.n441 42.8996
R532 vdd.n110 vdd.t118 41.8139
R533 vdd.n113 vdd.t125 41.8139
R534 vdd.n254 vdd.t48 41.8139
R535 vdd.n257 vdd.t54 41.8139
R536 vdd.n398 vdd.t65 41.8139
R537 vdd.n401 vdd.t159 41.8139
R538 vdd.n549 vdd.t30 41.8139
R539 vdd.n552 vdd.t19 41.8139
R540 vdd.n89 vdd.t132 35.1237
R541 vdd.n233 vdd.t42 35.1237
R542 vdd.n377 vdd.t38 35.1237
R543 vdd.n528 vdd.t57 35.1237
R544 vdd.n83 vdd.n82 33.0688
R545 vdd.n227 vdd.n226 33.0688
R546 vdd.n371 vdd.n370 33.0688
R547 vdd.n522 vdd.n521 33.0688
R548 vdd.n778 vdd.t81 26.5955
R549 vdd.n778 vdd.t109 26.5955
R550 vdd.n767 vdd.t127 26.5955
R551 vdd.n767 vdd.t120 26.5955
R552 vdd.n717 vdd.t99 26.5955
R553 vdd.n717 vdd.t95 26.5955
R554 vdd.n706 vdd.t52 26.5955
R555 vdd.n706 vdd.t50 26.5955
R556 vdd.n656 vdd.t89 26.5955
R557 vdd.n656 vdd.t79 26.5955
R558 vdd.n645 vdd.t26 26.5955
R559 vdd.n645 vdd.t36 26.5955
R560 vdd.n602 vdd.t93 26.5955
R561 vdd.n602 vdd.t97 26.5955
R562 vdd.n591 vdd.t163 26.5955
R563 vdd.n591 vdd.t5 26.5955
R564 vdd.n91 vdd.n88 25.6005
R565 vdd.n94 vdd.n91 25.6005
R566 vdd.n97 vdd.n94 25.6005
R567 vdd.n100 vdd.n97 25.6005
R568 vdd.n103 vdd.n100 25.6005
R569 vdd.n106 vdd.n103 25.6005
R570 vdd.n109 vdd.n106 25.6005
R571 vdd.n112 vdd.n109 25.6005
R572 vdd.n115 vdd.n112 25.6005
R573 vdd.n118 vdd.n115 25.6005
R574 vdd.n121 vdd.n118 25.6005
R575 vdd.n124 vdd.n121 25.6005
R576 vdd.n127 vdd.n124 25.6005
R577 vdd.n130 vdd.n127 25.6005
R578 vdd.n133 vdd.n130 25.6005
R579 vdd.n136 vdd.n133 25.6005
R580 vdd.n138 vdd.n136 25.6005
R581 vdd.n85 vdd.n81 25.6005
R582 vdd.n4 vdd.n1 25.6005
R583 vdd.n8 vdd.n6 25.6005
R584 vdd.n10 vdd.n8 25.6005
R585 vdd.n12 vdd.n10 25.6005
R586 vdd.n14 vdd.n12 25.6005
R587 vdd.n16 vdd.n14 25.6005
R588 vdd.n18 vdd.n16 25.6005
R589 vdd.n20 vdd.n18 25.6005
R590 vdd.n22 vdd.n20 25.6005
R591 vdd.n24 vdd.n22 25.6005
R592 vdd.n26 vdd.n24 25.6005
R593 vdd.n28 vdd.n26 25.6005
R594 vdd.n30 vdd.n28 25.6005
R595 vdd.n32 vdd.n30 25.6005
R596 vdd.n34 vdd.n32 25.6005
R597 vdd.n36 vdd.n34 25.6005
R598 vdd.n38 vdd.n36 25.6005
R599 vdd.n40 vdd.n38 25.6005
R600 vdd.n235 vdd.n232 25.6005
R601 vdd.n238 vdd.n235 25.6005
R602 vdd.n241 vdd.n238 25.6005
R603 vdd.n244 vdd.n241 25.6005
R604 vdd.n247 vdd.n244 25.6005
R605 vdd.n250 vdd.n247 25.6005
R606 vdd.n253 vdd.n250 25.6005
R607 vdd.n256 vdd.n253 25.6005
R608 vdd.n259 vdd.n256 25.6005
R609 vdd.n262 vdd.n259 25.6005
R610 vdd.n265 vdd.n262 25.6005
R611 vdd.n268 vdd.n265 25.6005
R612 vdd.n271 vdd.n268 25.6005
R613 vdd.n274 vdd.n271 25.6005
R614 vdd.n277 vdd.n274 25.6005
R615 vdd.n280 vdd.n277 25.6005
R616 vdd.n282 vdd.n280 25.6005
R617 vdd.n229 vdd.n225 25.6005
R618 vdd.n148 vdd.n145 25.6005
R619 vdd.n152 vdd.n150 25.6005
R620 vdd.n154 vdd.n152 25.6005
R621 vdd.n156 vdd.n154 25.6005
R622 vdd.n158 vdd.n156 25.6005
R623 vdd.n160 vdd.n158 25.6005
R624 vdd.n162 vdd.n160 25.6005
R625 vdd.n164 vdd.n162 25.6005
R626 vdd.n166 vdd.n164 25.6005
R627 vdd.n168 vdd.n166 25.6005
R628 vdd.n170 vdd.n168 25.6005
R629 vdd.n172 vdd.n170 25.6005
R630 vdd.n174 vdd.n172 25.6005
R631 vdd.n176 vdd.n174 25.6005
R632 vdd.n178 vdd.n176 25.6005
R633 vdd.n180 vdd.n178 25.6005
R634 vdd.n182 vdd.n180 25.6005
R635 vdd.n184 vdd.n182 25.6005
R636 vdd.n379 vdd.n376 25.6005
R637 vdd.n382 vdd.n379 25.6005
R638 vdd.n385 vdd.n382 25.6005
R639 vdd.n388 vdd.n385 25.6005
R640 vdd.n391 vdd.n388 25.6005
R641 vdd.n394 vdd.n391 25.6005
R642 vdd.n397 vdd.n394 25.6005
R643 vdd.n400 vdd.n397 25.6005
R644 vdd.n403 vdd.n400 25.6005
R645 vdd.n406 vdd.n403 25.6005
R646 vdd.n409 vdd.n406 25.6005
R647 vdd.n412 vdd.n409 25.6005
R648 vdd.n415 vdd.n412 25.6005
R649 vdd.n418 vdd.n415 25.6005
R650 vdd.n421 vdd.n418 25.6005
R651 vdd.n424 vdd.n421 25.6005
R652 vdd.n426 vdd.n424 25.6005
R653 vdd.n373 vdd.n369 25.6005
R654 vdd.n292 vdd.n289 25.6005
R655 vdd.n296 vdd.n294 25.6005
R656 vdd.n298 vdd.n296 25.6005
R657 vdd.n300 vdd.n298 25.6005
R658 vdd.n302 vdd.n300 25.6005
R659 vdd.n304 vdd.n302 25.6005
R660 vdd.n306 vdd.n304 25.6005
R661 vdd.n308 vdd.n306 25.6005
R662 vdd.n310 vdd.n308 25.6005
R663 vdd.n312 vdd.n310 25.6005
R664 vdd.n314 vdd.n312 25.6005
R665 vdd.n316 vdd.n314 25.6005
R666 vdd.n318 vdd.n316 25.6005
R667 vdd.n320 vdd.n318 25.6005
R668 vdd.n322 vdd.n320 25.6005
R669 vdd.n324 vdd.n322 25.6005
R670 vdd.n326 vdd.n324 25.6005
R671 vdd.n328 vdd.n326 25.6005
R672 vdd.n530 vdd.n527 25.6005
R673 vdd.n533 vdd.n530 25.6005
R674 vdd.n536 vdd.n533 25.6005
R675 vdd.n539 vdd.n536 25.6005
R676 vdd.n542 vdd.n539 25.6005
R677 vdd.n545 vdd.n542 25.6005
R678 vdd.n548 vdd.n545 25.6005
R679 vdd.n551 vdd.n548 25.6005
R680 vdd.n554 vdd.n551 25.6005
R681 vdd.n557 vdd.n554 25.6005
R682 vdd.n560 vdd.n557 25.6005
R683 vdd.n563 vdd.n560 25.6005
R684 vdd.n566 vdd.n563 25.6005
R685 vdd.n569 vdd.n566 25.6005
R686 vdd.n572 vdd.n569 25.6005
R687 vdd.n575 vdd.n572 25.6005
R688 vdd.n577 vdd.n575 25.6005
R689 vdd.n524 vdd.n520 25.6005
R690 vdd.n443 vdd.n440 25.6005
R691 vdd.n447 vdd.n445 25.6005
R692 vdd.n449 vdd.n447 25.6005
R693 vdd.n451 vdd.n449 25.6005
R694 vdd.n453 vdd.n451 25.6005
R695 vdd.n455 vdd.n453 25.6005
R696 vdd.n457 vdd.n455 25.6005
R697 vdd.n459 vdd.n457 25.6005
R698 vdd.n461 vdd.n459 25.6005
R699 vdd.n463 vdd.n461 25.6005
R700 vdd.n465 vdd.n463 25.6005
R701 vdd.n467 vdd.n465 25.6005
R702 vdd.n469 vdd.n467 25.6005
R703 vdd.n471 vdd.n469 25.6005
R704 vdd.n473 vdd.n471 25.6005
R705 vdd.n475 vdd.n473 25.6005
R706 vdd.n477 vdd.n475 25.6005
R707 vdd.n479 vdd.n477 25.6005
R708 vdd.n75 vdd.n74 19.0024
R709 vdd.n76 vdd.n75 19.0024
R710 vdd.n219 vdd.n218 19.0024
R711 vdd.n220 vdd.n219 19.0024
R712 vdd.n363 vdd.n362 19.0024
R713 vdd.n364 vdd.n363 19.0024
R714 vdd.n514 vdd.n513 19.0024
R715 vdd.n515 vdd.n514 19.0024
R716 vdd.n98 vdd.t129 18.3984
R717 vdd.n125 vdd.t135 18.3984
R718 vdd.n242 vdd.t55 18.3984
R719 vdd.n269 vdd.t44 18.3984
R720 vdd.n386 vdd.t0 18.3984
R721 vdd.n413 vdd.t136 18.3984
R722 vdd.n537 vdd.t75 18.3984
R723 vdd.n564 vdd.t20 18.3984
R724 vdd.n77 vdd.n76 17.6476
R725 vdd.n221 vdd.n220 17.6476
R726 vdd.n365 vdd.n364 17.6476
R727 vdd.n516 vdd.n515 17.6476
R728 vdd.n689 vdd.n688 17.1345
R729 vdd.n750 vdd.n749 17.1345
R730 vdd.n431 vdd.n430 17.1345
R731 vdd.n752 vdd.n744 14.2735
R732 vdd.n691 vdd.n683 14.2735
R733 vdd.n630 vdd.n629 14.2735
R734 vdd.n104 vdd.t131 11.7082
R735 vdd.n119 vdd.t130 11.7082
R736 vdd.n248 vdd.t43 11.7082
R737 vdd.n263 vdd.t56 11.7082
R738 vdd.n392 vdd.t3 11.7082
R739 vdd.n407 vdd.t27 11.7082
R740 vdd.n543 vdd.t6 11.7082
R741 vdd.n558 vdd.t117 11.7082
R742 vdd.n691 vdd.n690 9.7285
R743 vdd.n752 vdd.n751 9.7285
R744 vdd.n630 vdd.n435 9.7285
R745 vdd.n68 vdd.n67 9.56145
R746 vdd.n212 vdd.n211 9.56145
R747 vdd.n356 vdd.n355 9.56145
R748 vdd.n507 vdd.n506 9.56145
R749 vdd.n58 vdd.n57 9.3005
R750 vdd.n60 vdd.n59 9.3005
R751 vdd.n56 vdd.n55 9.3005
R752 vdd.n55 vdd.n54 9.3005
R753 vdd.n47 vdd.n46 9.3005
R754 vdd.n70 vdd.n69 9.3005
R755 vdd.n78 vdd.n77 9.3005
R756 vdd.n202 vdd.n201 9.3005
R757 vdd.n204 vdd.n203 9.3005
R758 vdd.n200 vdd.n199 9.3005
R759 vdd.n199 vdd.n198 9.3005
R760 vdd.n191 vdd.n190 9.3005
R761 vdd.n214 vdd.n213 9.3005
R762 vdd.n222 vdd.n221 9.3005
R763 vdd.n346 vdd.n345 9.3005
R764 vdd.n348 vdd.n347 9.3005
R765 vdd.n344 vdd.n343 9.3005
R766 vdd.n343 vdd.n342 9.3005
R767 vdd.n335 vdd.n334 9.3005
R768 vdd.n358 vdd.n357 9.3005
R769 vdd.n366 vdd.n365 9.3005
R770 vdd.n497 vdd.n496 9.3005
R771 vdd.n499 vdd.n498 9.3005
R772 vdd.n495 vdd.n494 9.3005
R773 vdd.n494 vdd.n493 9.3005
R774 vdd.n486 vdd.n485 9.3005
R775 vdd.n509 vdd.n508 9.3005
R776 vdd.n517 vdd.n516 9.3005
R777 vdd.n68 vdd.n65 8.39826
R778 vdd.n212 vdd.n209 8.39826
R779 vdd.n356 vdd.n353 8.39826
R780 vdd.n507 vdd.n504 8.39826
R781 vdd.n792 vdd.n791 7.11866
R782 vdd.n731 vdd.n730 7.11866
R783 vdd.n616 vdd.n615 7.11866
R784 vdd.n670 vdd.n669 7.11866
R785 vdd.n50 vdd.n49 6.02403
R786 vdd.n42 vdd.n41 6.02403
R787 vdd.n194 vdd.n193 6.02403
R788 vdd.n186 vdd.n185 6.02403
R789 vdd.n338 vdd.n337 6.02403
R790 vdd.n330 vdd.n329 6.02403
R791 vdd.n489 vdd.n488 6.02403
R792 vdd.n481 vdd.n480 6.02403
R793 vdd.n62 vdd.n61 5.27109
R794 vdd.n206 vdd.n205 5.27109
R795 vdd.n350 vdd.n349 5.27109
R796 vdd.n501 vdd.n500 5.27109
R797 vdd.n583 vdd.n581 5.07505
R798 vdd.n807 vdd.n806 4.95526
R799 vdd.n142 vdd.n141 4.67352
R800 vdd.n286 vdd.n285 4.67352
R801 vdd.n437 vdd.n436 4.67352
R802 vdd.n690 vdd.n686 4.65934
R803 vdd.n751 vdd.n747 4.65934
R804 vdd.n435 vdd.n434 4.65934
R805 vdd.n583 vdd.n582 4.6505
R806 vdd.n586 vdd.n585 4.6505
R807 vdd.n593 vdd.n592 4.6505
R808 vdd.n597 vdd.n596 4.6505
R809 vdd.n599 vdd.n598 4.6505
R810 vdd.n604 vdd.n603 4.6505
R811 vdd.n608 vdd.n607 4.6505
R812 vdd.n642 vdd.n641 4.6505
R813 vdd.n647 vdd.n646 4.6505
R814 vdd.n651 vdd.n650 4.6505
R815 vdd.n653 vdd.n652 4.6505
R816 vdd.n658 vdd.n657 4.6505
R817 vdd.n662 vdd.n661 4.6505
R818 vdd.n696 vdd.n695 4.6505
R819 vdd.n703 vdd.n702 4.6505
R820 vdd.n708 vdd.n707 4.6505
R821 vdd.n712 vdd.n711 4.6505
R822 vdd.n714 vdd.n713 4.6505
R823 vdd.n719 vdd.n718 4.6505
R824 vdd.n723 vdd.n722 4.6505
R825 vdd.n757 vdd.n756 4.6505
R826 vdd.n764 vdd.n763 4.6505
R827 vdd.n769 vdd.n768 4.6505
R828 vdd.n773 vdd.n772 4.6505
R829 vdd.n775 vdd.n774 4.6505
R830 vdd.n780 vdd.n779 4.6505
R831 vdd.n784 vdd.n783 4.6505
R832 vdd.n590 vdd.n589 4.6505
R833 vdd.n595 vdd.n594 4.6505
R834 vdd.n601 vdd.n600 4.6505
R835 vdd.n606 vdd.n605 4.6505
R836 vdd.n611 vdd.n610 4.6505
R837 vdd.n614 vdd.n613 4.6505
R838 vdd.n619 vdd.n618 4.6505
R839 vdd.n622 vdd.n621 4.6505
R840 vdd.n624 vdd.n623 4.6505
R841 vdd.n629 vdd.n628 4.6505
R842 vdd.n635 vdd.n634 4.6505
R843 vdd.n637 vdd.n636 4.6505
R844 vdd.n640 vdd.n639 4.6505
R845 vdd.n644 vdd.n643 4.6505
R846 vdd.n649 vdd.n648 4.6505
R847 vdd.n655 vdd.n654 4.6505
R848 vdd.n660 vdd.n659 4.6505
R849 vdd.n665 vdd.n664 4.6505
R850 vdd.n668 vdd.n667 4.6505
R851 vdd.n673 vdd.n672 4.6505
R852 vdd.n676 vdd.n675 4.6505
R853 vdd.n678 vdd.n677 4.6505
R854 vdd.n683 vdd.n682 4.6505
R855 vdd.n698 vdd.n697 4.6505
R856 vdd.n701 vdd.n700 4.6505
R857 vdd.n705 vdd.n704 4.6505
R858 vdd.n710 vdd.n709 4.6505
R859 vdd.n716 vdd.n715 4.6505
R860 vdd.n721 vdd.n720 4.6505
R861 vdd.n726 vdd.n725 4.6505
R862 vdd.n729 vdd.n728 4.6505
R863 vdd.n734 vdd.n733 4.6505
R864 vdd.n737 vdd.n736 4.6505
R865 vdd.n739 vdd.n738 4.6505
R866 vdd.n744 vdd.n743 4.6505
R867 vdd.n759 vdd.n758 4.6505
R868 vdd.n762 vdd.n761 4.6505
R869 vdd.n766 vdd.n765 4.6505
R870 vdd.n771 vdd.n770 4.6505
R871 vdd.n777 vdd.n776 4.6505
R872 vdd.n782 vdd.n781 4.6505
R873 vdd.n787 vdd.n786 4.6505
R874 vdd.n790 vdd.n789 4.6505
R875 vdd.n795 vdd.n794 4.6505
R876 vdd.n798 vdd.n797 4.6505
R877 vdd.n800 vdd.n799 4.6505
R878 vdd.n802 vdd.n801 4.6505
R879 vdd.n804 vdd.n803 4.6505
R880 vdd.n588 vdd.n587 4.6505
R881 vdd.n54 vdd.n53 4.56271
R882 vdd.n198 vdd.n197 4.56271
R883 vdd.n342 vdd.n341 4.56271
R884 vdd.n493 vdd.n492 4.56271
R885 vdd.n73 vdd.n72 4.51815
R886 vdd.n217 vdd.n216 4.51815
R887 vdd.n361 vdd.n360 4.51815
R888 vdd.n512 vdd.n511 4.51815
R889 vdd.n143 vdd.n142 4.36875
R890 vdd.n287 vdd.n286 4.36875
R891 vdd.n438 vdd.n437 4.36875
R892 vdd.n54 vdd.n52 3.52991
R893 vdd.n198 vdd.n196 3.52991
R894 vdd.n342 vdd.n340 3.52991
R895 vdd.n493 vdd.n491 3.52991
R896 vdd.n45 vdd.n44 3.30153
R897 vdd.n189 vdd.n188 3.30153
R898 vdd.n333 vdd.n332 3.30153
R899 vdd.n484 vdd.n483 3.30153
R900 vdd vdd.n815 3.09555
R901 vdd.n56 vdd.n48 2.31034
R902 vdd.n200 vdd.n192 2.31034
R903 vdd.n344 vdd.n336 2.31034
R904 vdd.n495 vdd.n487 2.31034
R905 vdd.n692 vdd.n691 2.29662
R906 vdd.n753 vdd.n752 2.29662
R907 vdd.n631 vdd.n630 2.29643
R908 vdd.n805 vdd.n140 2.25407
R909 vdd.n742 vdd.n284 2.25407
R910 vdd.n681 vdd.n428 2.25407
R911 vdd.n627 vdd.n579 2.25407
R912 vdd.n140 vdd.n71 2.09332
R913 vdd.n284 vdd.n215 2.09332
R914 vdd.n428 vdd.n359 2.09332
R915 vdd.n579 vdd.n510 2.09332
R916 vdd.n140 vdd.n139 2.07952
R917 vdd.n284 vdd.n283 2.07952
R918 vdd.n428 vdd.n427 2.07952
R919 vdd.n579 vdd.n578 2.07952
R920 vdd.n139 vdd.n78 2.05645
R921 vdd.n283 vdd.n222 2.05645
R922 vdd.n427 vdd.n366 2.05645
R923 vdd.n578 vdd.n517 2.05645
R924 vdd.n78 vdd.n73 1.88285
R925 vdd.n222 vdd.n217 1.88285
R926 vdd.n366 vdd.n361 1.88285
R927 vdd.n517 vdd.n512 1.88285
R928 vdd.n71 vdd.n70 1.83901
R929 vdd.n215 vdd.n214 1.83901
R930 vdd.n359 vdd.n358 1.83901
R931 vdd.n510 vdd.n509 1.83901
R932 vdd.n48 vdd.n47 1.59246
R933 vdd.n192 vdd.n191 1.59246
R934 vdd.n336 vdd.n335 1.59246
R935 vdd.n487 vdd.n486 1.59246
R936 vdd.n70 vdd.n62 1.12991
R937 vdd.n214 vdd.n206 1.12991
R938 vdd.n358 vdd.n350 1.12991
R939 vdd.n509 vdd.n501 1.12991
R940 vdd.n789 vdd.n788 0.935332
R941 vdd.n728 vdd.n727 0.935332
R942 vdd.n667 vdd.n666 0.935332
R943 vdd.n613 vdd.n612 0.935332
R944 vdd.n755 vdd.n754 0.863992
R945 vdd.n694 vdd.n693 0.863992
R946 vdd.n633 vdd.n632 0.863992
R947 vdd.n581 vdd.n580 0.863992
R948 vdd.n815 vdd.n814 0.689957
R949 vdd.n794 vdd.n793 0.539826
R950 vdd.n733 vdd.n732 0.539826
R951 vdd.n672 vdd.n671 0.539826
R952 vdd.n618 vdd.n617 0.539826
R953 vdd.n69 vdd.n68 0.481606
R954 vdd.n213 vdd.n212 0.481606
R955 vdd.n357 vdd.n356 0.481606
R956 vdd.n508 vdd.n507 0.481606
R957 vdd.n55 vdd.n50 0.376971
R958 vdd.n47 vdd.n42 0.376971
R959 vdd.n199 vdd.n194 0.376971
R960 vdd.n191 vdd.n186 0.376971
R961 vdd.n343 vdd.n338 0.376971
R962 vdd.n335 vdd.n330 0.376971
R963 vdd.n494 vdd.n489 0.376971
R964 vdd.n486 vdd.n481 0.376971
R965 vdd.n756 vdd.n755 0.305262
R966 vdd.n761 vdd.n760 0.305262
R967 vdd.n744 vdd.n143 0.305262
R968 vdd.n695 vdd.n694 0.305262
R969 vdd.n700 vdd.n699 0.305262
R970 vdd.n683 vdd.n287 0.305262
R971 vdd.n634 vdd.n633 0.305262
R972 vdd.n639 vdd.n638 0.305262
R973 vdd.n629 vdd.n438 0.305262
R974 vdd.n585 vdd.n584 0.305262
R975 vdd.n786 vdd.n785 0.21623
R976 vdd.n725 vdd.n724 0.21623
R977 vdd.n664 vdd.n663 0.21623
R978 vdd.n610 vdd.n609 0.21623
R979 vdd.n809 vdd 0.191688
R980 vdd.n696 vdd.n692 0.180294
R981 vdd.n757 vdd.n753 0.180294
R982 vdd.n635 vdd.n631 0.179926
R983 vdd.n46 vdd.n45 0.166918
R984 vdd.n190 vdd.n189 0.166918
R985 vdd.n334 vdd.n333 0.166918
R986 vdd.n485 vdd.n484 0.166918
R987 vdd.n797 vdd.n796 0.14432
R988 vdd.n736 vdd.n735 0.14432
R989 vdd.n675 vdd.n674 0.14432
R990 vdd.n621 vdd.n620 0.14432
R991 vdd.n692 vdd 0.120655
R992 vdd.n753 vdd 0.120655
R993 vdd.n586 vdd.n583 0.120292
R994 vdd.n588 vdd.n586 0.120292
R995 vdd.n590 vdd.n588 0.120292
R996 vdd.n593 vdd.n590 0.120292
R997 vdd.n595 vdd.n593 0.120292
R998 vdd.n597 vdd.n595 0.120292
R999 vdd.n599 vdd.n597 0.120292
R1000 vdd.n601 vdd.n599 0.120292
R1001 vdd.n604 vdd.n601 0.120292
R1002 vdd.n606 vdd.n604 0.120292
R1003 vdd.n608 vdd.n606 0.120292
R1004 vdd.n611 vdd.n608 0.120292
R1005 vdd.n614 vdd.n611 0.120292
R1006 vdd.n619 vdd.n614 0.120292
R1007 vdd.n622 vdd.n619 0.120292
R1008 vdd.n624 vdd.n622 0.120292
R1009 vdd.n625 vdd.n624 0.120292
R1010 vdd.n626 vdd.n625 0.120292
R1011 vdd.n637 vdd.n635 0.120292
R1012 vdd.n640 vdd.n637 0.120292
R1013 vdd.n642 vdd.n640 0.120292
R1014 vdd.n644 vdd.n642 0.120292
R1015 vdd.n647 vdd.n644 0.120292
R1016 vdd.n649 vdd.n647 0.120292
R1017 vdd.n651 vdd.n649 0.120292
R1018 vdd.n653 vdd.n651 0.120292
R1019 vdd.n655 vdd.n653 0.120292
R1020 vdd.n658 vdd.n655 0.120292
R1021 vdd.n660 vdd.n658 0.120292
R1022 vdd.n662 vdd.n660 0.120292
R1023 vdd.n665 vdd.n662 0.120292
R1024 vdd.n668 vdd.n665 0.120292
R1025 vdd.n673 vdd.n668 0.120292
R1026 vdd.n676 vdd.n673 0.120292
R1027 vdd.n678 vdd.n676 0.120292
R1028 vdd.n679 vdd.n678 0.120292
R1029 vdd.n680 vdd.n679 0.120292
R1030 vdd.n698 vdd.n696 0.120292
R1031 vdd.n701 vdd.n698 0.120292
R1032 vdd.n703 vdd.n701 0.120292
R1033 vdd.n705 vdd.n703 0.120292
R1034 vdd.n708 vdd.n705 0.120292
R1035 vdd.n710 vdd.n708 0.120292
R1036 vdd.n712 vdd.n710 0.120292
R1037 vdd.n714 vdd.n712 0.120292
R1038 vdd.n716 vdd.n714 0.120292
R1039 vdd.n719 vdd.n716 0.120292
R1040 vdd.n721 vdd.n719 0.120292
R1041 vdd.n723 vdd.n721 0.120292
R1042 vdd.n726 vdd.n723 0.120292
R1043 vdd.n729 vdd.n726 0.120292
R1044 vdd.n734 vdd.n729 0.120292
R1045 vdd.n737 vdd.n734 0.120292
R1046 vdd.n739 vdd.n737 0.120292
R1047 vdd.n740 vdd.n739 0.120292
R1048 vdd.n741 vdd.n740 0.120292
R1049 vdd.n759 vdd.n757 0.120292
R1050 vdd.n762 vdd.n759 0.120292
R1051 vdd.n764 vdd.n762 0.120292
R1052 vdd.n766 vdd.n764 0.120292
R1053 vdd.n769 vdd.n766 0.120292
R1054 vdd.n771 vdd.n769 0.120292
R1055 vdd.n773 vdd.n771 0.120292
R1056 vdd.n775 vdd.n773 0.120292
R1057 vdd.n777 vdd.n775 0.120292
R1058 vdd.n780 vdd.n777 0.120292
R1059 vdd.n782 vdd.n780 0.120292
R1060 vdd.n784 vdd.n782 0.120292
R1061 vdd.n787 vdd.n784 0.120292
R1062 vdd.n790 vdd.n787 0.120292
R1063 vdd.n795 vdd.n790 0.120292
R1064 vdd.n798 vdd.n795 0.120292
R1065 vdd.n800 vdd.n798 0.120292
R1066 vdd.n802 vdd.n800 0.120292
R1067 vdd.n804 vdd.n802 0.120292
R1068 vdd.n631 vdd 0.12003
R1069 vdd.n140 vdd.n60 0.117348
R1070 vdd.n284 vdd.n204 0.117348
R1071 vdd.n428 vdd.n348 0.117348
R1072 vdd.n579 vdd.n499 0.117348
R1073 vdd.n628 vdd.n627 0.0968542
R1074 vdd.n682 vdd.n681 0.0968542
R1075 vdd.n743 vdd.n742 0.0968542
R1076 vdd.n807 vdd.n805 0.0968542
R1077 vdd.n628 vdd 0.0603958
R1078 vdd.n682 vdd 0.0603958
R1079 vdd.n743 vdd 0.0603958
R1080 vdd vdd.n807 0.0603958
R1081 vdd.n60 vdd.n58 0.0439783
R1082 vdd.n204 vdd.n202 0.0439783
R1083 vdd.n348 vdd.n346 0.0439783
R1084 vdd.n499 vdd.n497 0.0439783
R1085 vdd.n815 vdd.n808 0.0290714
R1086 vdd.n814 vdd.n813 0.0240572
R1087 vdd.n627 vdd.n626 0.0239375
R1088 vdd.n681 vdd.n680 0.0239375
R1089 vdd.n742 vdd.n741 0.0239375
R1090 vdd.n805 vdd.n804 0.0239375
R1091 vdd.n812 vdd.n811 0.0205
R1092 vdd.n813 vdd.n812 0.0205
R1093 vdd.n814 vdd.n810 0.0163636
R1094 vdd.n810 vdd.n809 0.011753
R1095 vdd.n58 vdd.n56 0.00321739
R1096 vdd.n202 vdd.n200 0.00321739
R1097 vdd.n346 vdd.n344 0.00321739
R1098 vdd.n497 vdd.n495 0.00321739
R1099 vss.n184 vss.n183 18699.7
R1100 vss.n185 vss.n184 4406.54
R1101 vss.n183 vss.n182 3471.83
R1102 vss.t123 vss.t102 2592.76
R1103 vss.t135 vss.t88 2592.76
R1104 vss.t144 vss.t98 2592.76
R1105 vss.t86 vss.t132 2592.76
R1106 vss.n758 vss.t123 2274.16
R1107 vss.n816 vss.t135 2274.16
R1108 vss.n874 vss.t144 2274.16
R1109 vss.n671 vss.n670 1717.31
R1110 vss.n509 vss.n508 1717.31
R1111 vss.n347 vss.n346 1717.31
R1112 vss.t17 vss.t129 1329.34
R1113 vss.t141 vss.t15 1329.34
R1114 vss.t126 vss.t64 1329.34
R1115 vss.t138 vss.t153 1329.34
R1116 vss.t90 vss.t121 1142.57
R1117 vss.t3 vss.t100 1142.57
R1118 vss.t66 vss.t116 1142.57
R1119 vss.t149 vss.t106 1142.57
R1120 vss.t32 vss.t159 1068.02
R1121 vss.t19 vss.t0 1068.02
R1122 vss.t161 vss.t27 1068.02
R1123 vss.t76 vss.t155 1068.02
R1124 vss.t72 vss.t74 1068.02
R1125 vss.t51 vss.t82 1068.02
R1126 vss.t157 vss.t24 1068.02
R1127 vss.n762 vss.t141 1010.74
R1128 vss.n820 vss.t126 1010.74
R1129 vss.n878 vss.t138 1010.74
R1130 vss.n112 vss.t30 789.886
R1131 vss.n107 vss.t80 789.886
R1132 vss.n671 vss.n669 611.246
R1133 vss.n509 vss.n507 611.246
R1134 vss.n347 vss.n345 611.246
R1135 vss.n185 vss.n106 611.246
R1136 vss.n182 vss.n107 511.757
R1137 vss.t30 vss.t32 467.257
R1138 vss.t159 vss.t19 467.257
R1139 vss.t0 vss.t161 467.257
R1140 vss.t27 vss.t78 467.257
R1141 vss.t155 vss.t34 467.257
R1142 vss.t74 vss.t76 467.257
R1143 vss.t82 vss.t72 467.257
R1144 vss.t24 vss.t51 467.257
R1145 vss.t80 vss.t157 467.257
R1146 vss.t84 vss.t17 461.423
R1147 vss.t118 vss.t84 461.423
R1148 vss.t121 vss.t118 461.423
R1149 vss.t108 vss.t90 461.423
R1150 vss.t112 vss.t108 461.423
R1151 vss.t102 vss.t112 461.423
R1152 vss.t15 vss.t49 461.423
R1153 vss.t49 vss.t46 461.423
R1154 vss.t46 vss.t3 461.423
R1155 vss.t100 vss.t104 461.423
R1156 vss.t88 vss.t94 461.423
R1157 vss.t64 vss.t70 461.423
R1158 vss.t70 vss.t68 461.423
R1159 vss.t68 vss.t66 461.423
R1160 vss.t116 vss.t114 461.423
R1161 vss.t98 vss.t110 461.423
R1162 vss.t153 vss.t151 461.423
R1163 vss.t151 vss.t147 461.423
R1164 vss.t147 vss.t149 461.423
R1165 vss.t106 vss.t96 461.423
R1166 vss.t96 vss.t92 461.423
R1167 vss.t92 vss.t86 461.423
R1168 vss.n115 vss.n111 294.462
R1169 vss.n114 vss.n113 292.5
R1170 vss.n113 vss.n112 292.5
R1171 vss.n181 vss.n180 292.5
R1172 vss.n182 vss.n181 292.5
R1173 vss.n111 vss.n110 292.5
R1174 vss.n664 vss.n663 292.5
R1175 vss.n662 vss.n661 292.5
R1176 vss.n660 vss.n659 292.5
R1177 vss.n658 vss.n657 292.5
R1178 vss.n656 vss.n655 292.5
R1179 vss.n654 vss.n653 292.5
R1180 vss.n652 vss.n651 292.5
R1181 vss.n650 vss.n649 292.5
R1182 vss.n648 vss.n647 292.5
R1183 vss.n646 vss.n645 292.5
R1184 vss.n644 vss.n643 292.5
R1185 vss.n642 vss.n641 292.5
R1186 vss.n640 vss.n639 292.5
R1187 vss.n638 vss.n637 292.5
R1188 vss.n636 vss.n635 292.5
R1189 vss.n634 vss.n633 292.5
R1190 vss.n632 vss.n631 292.5
R1191 vss.n630 vss.n629 292.5
R1192 vss.n628 vss.n627 292.5
R1193 vss.n625 vss.n624 292.5
R1194 vss.n565 vss.n564 292.5
R1195 vss.n569 vss.n568 292.5
R1196 vss.n572 vss.n571 292.5
R1197 vss.n571 vss.n570 292.5
R1198 vss.n575 vss.n574 292.5
R1199 vss.n574 vss.n573 292.5
R1200 vss.n578 vss.n577 292.5
R1201 vss.n577 vss.n576 292.5
R1202 vss.n581 vss.n580 292.5
R1203 vss.n580 vss.n579 292.5
R1204 vss.n584 vss.n583 292.5
R1205 vss.n583 vss.n582 292.5
R1206 vss.n587 vss.n586 292.5
R1207 vss.n586 vss.n585 292.5
R1208 vss.n590 vss.n589 292.5
R1209 vss.n589 vss.n588 292.5
R1210 vss.n593 vss.n592 292.5
R1211 vss.n592 vss.n591 292.5
R1212 vss.n596 vss.n595 292.5
R1213 vss.n595 vss.n594 292.5
R1214 vss.n599 vss.n598 292.5
R1215 vss.n598 vss.n597 292.5
R1216 vss.n602 vss.n601 292.5
R1217 vss.n601 vss.n600 292.5
R1218 vss.n605 vss.n604 292.5
R1219 vss.n604 vss.n603 292.5
R1220 vss.n608 vss.n607 292.5
R1221 vss.n607 vss.n606 292.5
R1222 vss.n611 vss.n610 292.5
R1223 vss.n610 vss.n609 292.5
R1224 vss.n614 vss.n613 292.5
R1225 vss.n613 vss.n612 292.5
R1226 vss.n617 vss.n616 292.5
R1227 vss.n616 vss.n615 292.5
R1228 vss.n620 vss.n619 292.5
R1229 vss.n619 vss.n618 292.5
R1230 vss.n622 vss.n621 292.5
R1231 vss.n502 vss.n501 292.5
R1232 vss.n500 vss.n499 292.5
R1233 vss.n498 vss.n497 292.5
R1234 vss.n496 vss.n495 292.5
R1235 vss.n494 vss.n493 292.5
R1236 vss.n492 vss.n491 292.5
R1237 vss.n490 vss.n489 292.5
R1238 vss.n488 vss.n487 292.5
R1239 vss.n486 vss.n485 292.5
R1240 vss.n484 vss.n483 292.5
R1241 vss.n482 vss.n481 292.5
R1242 vss.n480 vss.n479 292.5
R1243 vss.n478 vss.n477 292.5
R1244 vss.n476 vss.n475 292.5
R1245 vss.n474 vss.n473 292.5
R1246 vss.n472 vss.n471 292.5
R1247 vss.n470 vss.n469 292.5
R1248 vss.n468 vss.n467 292.5
R1249 vss.n466 vss.n465 292.5
R1250 vss.n463 vss.n462 292.5
R1251 vss.n403 vss.n402 292.5
R1252 vss.n407 vss.n406 292.5
R1253 vss.n410 vss.n409 292.5
R1254 vss.n409 vss.n408 292.5
R1255 vss.n413 vss.n412 292.5
R1256 vss.n412 vss.n411 292.5
R1257 vss.n416 vss.n415 292.5
R1258 vss.n415 vss.n414 292.5
R1259 vss.n419 vss.n418 292.5
R1260 vss.n418 vss.n417 292.5
R1261 vss.n422 vss.n421 292.5
R1262 vss.n421 vss.n420 292.5
R1263 vss.n425 vss.n424 292.5
R1264 vss.n424 vss.n423 292.5
R1265 vss.n428 vss.n427 292.5
R1266 vss.n427 vss.n426 292.5
R1267 vss.n431 vss.n430 292.5
R1268 vss.n430 vss.n429 292.5
R1269 vss.n434 vss.n433 292.5
R1270 vss.n433 vss.n432 292.5
R1271 vss.n437 vss.n436 292.5
R1272 vss.n436 vss.n435 292.5
R1273 vss.n440 vss.n439 292.5
R1274 vss.n439 vss.n438 292.5
R1275 vss.n443 vss.n442 292.5
R1276 vss.n442 vss.n441 292.5
R1277 vss.n446 vss.n445 292.5
R1278 vss.n445 vss.n444 292.5
R1279 vss.n449 vss.n448 292.5
R1280 vss.n448 vss.n447 292.5
R1281 vss.n452 vss.n451 292.5
R1282 vss.n451 vss.n450 292.5
R1283 vss.n455 vss.n454 292.5
R1284 vss.n454 vss.n453 292.5
R1285 vss.n458 vss.n457 292.5
R1286 vss.n457 vss.n456 292.5
R1287 vss.n460 vss.n459 292.5
R1288 vss.n340 vss.n339 292.5
R1289 vss.n338 vss.n337 292.5
R1290 vss.n336 vss.n335 292.5
R1291 vss.n334 vss.n333 292.5
R1292 vss.n332 vss.n331 292.5
R1293 vss.n330 vss.n329 292.5
R1294 vss.n328 vss.n327 292.5
R1295 vss.n326 vss.n325 292.5
R1296 vss.n324 vss.n323 292.5
R1297 vss.n322 vss.n321 292.5
R1298 vss.n320 vss.n319 292.5
R1299 vss.n318 vss.n317 292.5
R1300 vss.n316 vss.n315 292.5
R1301 vss.n314 vss.n313 292.5
R1302 vss.n312 vss.n311 292.5
R1303 vss.n310 vss.n309 292.5
R1304 vss.n308 vss.n307 292.5
R1305 vss.n306 vss.n305 292.5
R1306 vss.n304 vss.n303 292.5
R1307 vss.n301 vss.n300 292.5
R1308 vss.n241 vss.n240 292.5
R1309 vss.n245 vss.n244 292.5
R1310 vss.n248 vss.n247 292.5
R1311 vss.n247 vss.n246 292.5
R1312 vss.n251 vss.n250 292.5
R1313 vss.n250 vss.n249 292.5
R1314 vss.n254 vss.n253 292.5
R1315 vss.n253 vss.n252 292.5
R1316 vss.n257 vss.n256 292.5
R1317 vss.n256 vss.n255 292.5
R1318 vss.n260 vss.n259 292.5
R1319 vss.n259 vss.n258 292.5
R1320 vss.n263 vss.n262 292.5
R1321 vss.n262 vss.n261 292.5
R1322 vss.n266 vss.n265 292.5
R1323 vss.n265 vss.n264 292.5
R1324 vss.n269 vss.n268 292.5
R1325 vss.n268 vss.n267 292.5
R1326 vss.n272 vss.n271 292.5
R1327 vss.n271 vss.n270 292.5
R1328 vss.n275 vss.n274 292.5
R1329 vss.n274 vss.n273 292.5
R1330 vss.n278 vss.n277 292.5
R1331 vss.n277 vss.n276 292.5
R1332 vss.n281 vss.n280 292.5
R1333 vss.n280 vss.n279 292.5
R1334 vss.n284 vss.n283 292.5
R1335 vss.n283 vss.n282 292.5
R1336 vss.n287 vss.n286 292.5
R1337 vss.n286 vss.n285 292.5
R1338 vss.n290 vss.n289 292.5
R1339 vss.n289 vss.n288 292.5
R1340 vss.n293 vss.n292 292.5
R1341 vss.n292 vss.n291 292.5
R1342 vss.n296 vss.n295 292.5
R1343 vss.n295 vss.n294 292.5
R1344 vss.n298 vss.n297 292.5
R1345 vss.n101 vss.n100 292.5
R1346 vss.n99 vss.n98 292.5
R1347 vss.n97 vss.n96 292.5
R1348 vss.n95 vss.n94 292.5
R1349 vss.n93 vss.n92 292.5
R1350 vss.n91 vss.n90 292.5
R1351 vss.n89 vss.n88 292.5
R1352 vss.n87 vss.n86 292.5
R1353 vss.n85 vss.n84 292.5
R1354 vss.n83 vss.n82 292.5
R1355 vss.n81 vss.n80 292.5
R1356 vss.n79 vss.n78 292.5
R1357 vss.n77 vss.n76 292.5
R1358 vss.n75 vss.n74 292.5
R1359 vss.n73 vss.n72 292.5
R1360 vss.n71 vss.n70 292.5
R1361 vss.n69 vss.n68 292.5
R1362 vss.n67 vss.n66 292.5
R1363 vss.n65 vss.n64 292.5
R1364 vss.n62 vss.n61 292.5
R1365 vss.n2 vss.n1 292.5
R1366 vss.n6 vss.n5 292.5
R1367 vss.n9 vss.n8 292.5
R1368 vss.n8 vss.n7 292.5
R1369 vss.n12 vss.n11 292.5
R1370 vss.n11 vss.n10 292.5
R1371 vss.n15 vss.n14 292.5
R1372 vss.n14 vss.n13 292.5
R1373 vss.n18 vss.n17 292.5
R1374 vss.n17 vss.n16 292.5
R1375 vss.n21 vss.n20 292.5
R1376 vss.n20 vss.n19 292.5
R1377 vss.n24 vss.n23 292.5
R1378 vss.n23 vss.n22 292.5
R1379 vss.n27 vss.n26 292.5
R1380 vss.n26 vss.n25 292.5
R1381 vss.n30 vss.n29 292.5
R1382 vss.n29 vss.n28 292.5
R1383 vss.n33 vss.n32 292.5
R1384 vss.n32 vss.n31 292.5
R1385 vss.n36 vss.n35 292.5
R1386 vss.n35 vss.n34 292.5
R1387 vss.n39 vss.n38 292.5
R1388 vss.n38 vss.n37 292.5
R1389 vss.n42 vss.n41 292.5
R1390 vss.n41 vss.n40 292.5
R1391 vss.n45 vss.n44 292.5
R1392 vss.n44 vss.n43 292.5
R1393 vss.n48 vss.n47 292.5
R1394 vss.n47 vss.n46 292.5
R1395 vss.n51 vss.n50 292.5
R1396 vss.n50 vss.n49 292.5
R1397 vss.n54 vss.n53 292.5
R1398 vss.n53 vss.n52 292.5
R1399 vss.n57 vss.n56 292.5
R1400 vss.n56 vss.n55 292.5
R1401 vss.n59 vss.n58 292.5
R1402 vss.n880 vss.n879 292.5
R1403 vss.n879 vss.n878 292.5
R1404 vss.n876 vss.n875 292.5
R1405 vss.n875 vss.n874 292.5
R1406 vss.n822 vss.n821 292.5
R1407 vss.n821 vss.n820 292.5
R1408 vss.n818 vss.n817 292.5
R1409 vss.n817 vss.n816 292.5
R1410 vss.n764 vss.n763 292.5
R1411 vss.n763 vss.n762 292.5
R1412 vss.n760 vss.n759 292.5
R1413 vss.n759 vss.n758 292.5
R1414 vss.n911 vss.t87 193.933
R1415 vss.n900 vss.t150 193.933
R1416 vss.n853 vss.t99 193.933
R1417 vss.n842 vss.t67 193.933
R1418 vss.n795 vss.t89 193.933
R1419 vss.n784 vss.t4 193.933
R1420 vss.n737 vss.t103 193.933
R1421 vss.n726 vss.t122 193.933
R1422 vss.n902 vss.t107 192.982
R1423 vss.n891 vss.t154 192.982
R1424 vss.n844 vss.t117 192.982
R1425 vss.n833 vss.t65 192.982
R1426 vss.n786 vss.t101 192.982
R1427 vss.n775 vss.t16 192.982
R1428 vss.n728 vss.t91 192.982
R1429 vss.n717 vss.t18 192.982
R1430 vss.n713 vss.t168 183.082
R1431 vss.n771 vss.t164 183.082
R1432 vss.n829 vss.t169 183.082
R1433 vss.n887 vss.t165 183.082
R1434 vss.n181 vss.n108 172.611
R1435 vss.n564 vss.n563 147.374
R1436 vss.n402 vss.n401 147.374
R1437 vss.n240 vss.n239 147.374
R1438 vss.n1 vss.n0 147.374
R1439 vss.n576 vss.t120 140.685
R1440 vss.n615 vss.t26 140.685
R1441 vss.n414 vss.t41 140.685
R1442 vss.n453 vss.t42 140.685
R1443 vss.n252 vss.t14 140.685
R1444 vss.n291 vss.t6 140.685
R1445 vss.n13 vss.t59 140.685
R1446 vss.n52 vss.t60 140.685
R1447 vss.n567 vss.n566 134.577
R1448 vss.n405 vss.n404 134.577
R1449 vss.n243 vss.n242 134.577
R1450 vss.n4 vss.n3 134.577
R1451 vss.n712 vss.t130 123.918
R1452 vss.n714 vss.t131 121.956
R1453 vss.n739 vss.t124 121.956
R1454 vss.n562 vss.t125 121.956
R1455 vss.n766 vss.t142 121.956
R1456 vss.n772 vss.t143 121.956
R1457 vss.n797 vss.t136 121.956
R1458 vss.n400 vss.t137 121.956
R1459 vss.n824 vss.t127 121.956
R1460 vss.n830 vss.t128 121.956
R1461 vss.n855 vss.t145 121.956
R1462 vss.n238 vss.t146 121.956
R1463 vss.n882 vss.t139 121.956
R1464 vss.n888 vss.t140 121.956
R1465 vss.n913 vss.t133 121.956
R1466 vss.n942 vss.t134 121.956
R1467 vss.n594 vss.t63 121.279
R1468 vss.n597 vss.t48 121.279
R1469 vss.n432 vss.t40 121.279
R1470 vss.n435 vss.t44 121.279
R1471 vss.n270 vss.t5 121.279
R1472 vss.n273 vss.t7 121.279
R1473 vss.n31 vss.t58 121.279
R1474 vss.n34 vss.t61 121.279
R1475 vss.n907 vss.n906 121.112
R1476 vss.n896 vss.n895 121.112
R1477 vss.n849 vss.n848 121.112
R1478 vss.n838 vss.n837 121.112
R1479 vss.n791 vss.n790 121.112
R1480 vss.n780 vss.n779 121.112
R1481 vss.n733 vss.n732 121.112
R1482 vss.n722 vss.n721 121.112
R1483 vss.n168 vss.t81 116.115
R1484 vss.n162 vss.t25 116.115
R1485 vss.n156 vss.t83 116.115
R1486 vss.n150 vss.t75 116.115
R1487 vss.n144 vss.t156 116.115
R1488 vss.n138 vss.t79 116.115
R1489 vss.n132 vss.t162 116.115
R1490 vss.n126 vss.t20 116.115
R1491 vss.n120 vss.t33 116.115
R1492 vss.n164 vss.t158 113.677
R1493 vss.n158 vss.t52 113.677
R1494 vss.n152 vss.t73 113.677
R1495 vss.n146 vss.t77 113.677
R1496 vss.n140 vss.t35 113.677
R1497 vss.n134 vss.t28 113.677
R1498 vss.n128 vss.t1 113.677
R1499 vss.n122 vss.t160 113.677
R1500 vss.n116 vss.t31 113.677
R1501 vss.n573 vss.t22 101.874
R1502 vss.n618 vss.t163 101.874
R1503 vss.n411 vss.t39 101.874
R1504 vss.n456 vss.t45 101.874
R1505 vss.n249 vss.t11 101.874
R1506 vss.n294 vss.t10 101.874
R1507 vss.n10 vss.t56 101.874
R1508 vss.n55 vss.t62 101.874
R1509 vss.n568 vss.n567 90.6382
R1510 vss.n406 vss.n405 90.6382
R1511 vss.n244 vss.n243 90.6382
R1512 vss.n5 vss.n4 90.6382
R1513 vss.n64 vss.n63 90.6381
R1514 vss.n303 vss.n302 90.6381
R1515 vss.n465 vss.n464 90.6381
R1516 vss.n627 vss.n626 90.6381
R1517 vss.n9 vss.n6 87.7181
R1518 vss.n67 vss.n65 87.7181
R1519 vss.n248 vss.n245 87.7181
R1520 vss.n306 vss.n304 87.7181
R1521 vss.n410 vss.n407 87.7181
R1522 vss.n468 vss.n466 87.7181
R1523 vss.n572 vss.n569 87.7181
R1524 vss.n630 vss.n628 87.7181
R1525 vss.n105 vss.n104 86.9123
R1526 vss.n344 vss.n343 86.9123
R1527 vss.n506 vss.n505 86.9123
R1528 vss.n668 vss.n667 86.9123
R1529 vss.n102 vss.n101 82.0711
R1530 vss.n341 vss.n340 82.0711
R1531 vss.n503 vss.n502 82.0711
R1532 vss.n665 vss.n664 82.0711
R1533 vss.n60 vss.n59 78.3064
R1534 vss.n299 vss.n298 78.3064
R1535 vss.n461 vss.n460 78.3064
R1536 vss.n623 vss.n622 78.3064
R1537 vss.n938 vss.n937 76.0005
R1538 vss.n235 vss.n234 76.0005
R1539 vss.n397 vss.n396 76.0005
R1540 vss.n559 vss.n558 76.0005
R1541 vss.n206 vss.n205 63.7358
R1542 vss.n368 vss.n367 63.7358
R1543 vss.n530 vss.n529 63.7358
R1544 vss.n692 vss.n691 63.7358
R1545 vss.n582 vss.t29 53.3632
R1546 vss.n609 vss.t21 53.3632
R1547 vss.n420 vss.t43 53.3632
R1548 vss.n447 vss.t37 53.3632
R1549 vss.n258 vss.t8 53.3632
R1550 vss.n285 vss.t13 53.3632
R1551 vss.n19 vss.t53 53.3632
R1552 vss.n46 vss.t57 53.3632
R1553 vss.n220 vss.n219 46.3534
R1554 vss.n382 vss.n381 46.3534
R1555 vss.n544 vss.n543 46.3534
R1556 vss.n706 vss.n705 46.3534
R1557 vss.n195 vss.n194 35.3848
R1558 vss.n357 vss.n356 35.3848
R1559 vss.n519 vss.n518 35.3848
R1560 vss.n681 vss.n680 35.3848
R1561 vss.n680 vss.n679 35.3848
R1562 vss.n518 vss.n517 35.3848
R1563 vss.n356 vss.n355 35.3848
R1564 vss.n194 vss.n193 35.3848
R1565 vss.n557 vss.t170 34.2973
R1566 vss.n395 vss.t166 34.2973
R1567 vss.n233 vss.t171 34.2973
R1568 vss.n936 vss.t167 34.2973
R1569 vss.n588 vss.t2 33.9586
R1570 vss.n603 vss.t23 33.9586
R1571 vss.n426 vss.t36 33.9586
R1572 vss.n441 vss.t38 33.9586
R1573 vss.n264 vss.t12 33.9586
R1574 vss.n279 vss.t9 33.9586
R1575 vss.n25 vss.t55 33.9586
R1576 vss.n40 vss.t54 33.9586
R1577 vss.n693 vss.n692 32.3305
R1578 vss.n531 vss.n530 32.3305
R1579 vss.n369 vss.n368 32.3305
R1580 vss.n207 vss.n206 32.3305
R1581 vss.n12 vss.n9 25.6005
R1582 vss.n15 vss.n12 25.6005
R1583 vss.n18 vss.n15 25.6005
R1584 vss.n21 vss.n18 25.6005
R1585 vss.n24 vss.n21 25.6005
R1586 vss.n27 vss.n24 25.6005
R1587 vss.n30 vss.n27 25.6005
R1588 vss.n33 vss.n30 25.6005
R1589 vss.n36 vss.n33 25.6005
R1590 vss.n39 vss.n36 25.6005
R1591 vss.n42 vss.n39 25.6005
R1592 vss.n45 vss.n42 25.6005
R1593 vss.n48 vss.n45 25.6005
R1594 vss.n51 vss.n48 25.6005
R1595 vss.n54 vss.n51 25.6005
R1596 vss.n57 vss.n54 25.6005
R1597 vss.n59 vss.n57 25.6005
R1598 vss.n6 vss.n2 25.6005
R1599 vss.n65 vss.n62 25.6005
R1600 vss.n69 vss.n67 25.6005
R1601 vss.n71 vss.n69 25.6005
R1602 vss.n73 vss.n71 25.6005
R1603 vss.n75 vss.n73 25.6005
R1604 vss.n77 vss.n75 25.6005
R1605 vss.n79 vss.n77 25.6005
R1606 vss.n81 vss.n79 25.6005
R1607 vss.n83 vss.n81 25.6005
R1608 vss.n85 vss.n83 25.6005
R1609 vss.n87 vss.n85 25.6005
R1610 vss.n89 vss.n87 25.6005
R1611 vss.n91 vss.n89 25.6005
R1612 vss.n93 vss.n91 25.6005
R1613 vss.n95 vss.n93 25.6005
R1614 vss.n97 vss.n95 25.6005
R1615 vss.n99 vss.n97 25.6005
R1616 vss.n101 vss.n99 25.6005
R1617 vss.n251 vss.n248 25.6005
R1618 vss.n254 vss.n251 25.6005
R1619 vss.n257 vss.n254 25.6005
R1620 vss.n260 vss.n257 25.6005
R1621 vss.n263 vss.n260 25.6005
R1622 vss.n266 vss.n263 25.6005
R1623 vss.n269 vss.n266 25.6005
R1624 vss.n272 vss.n269 25.6005
R1625 vss.n275 vss.n272 25.6005
R1626 vss.n278 vss.n275 25.6005
R1627 vss.n281 vss.n278 25.6005
R1628 vss.n284 vss.n281 25.6005
R1629 vss.n287 vss.n284 25.6005
R1630 vss.n290 vss.n287 25.6005
R1631 vss.n293 vss.n290 25.6005
R1632 vss.n296 vss.n293 25.6005
R1633 vss.n298 vss.n296 25.6005
R1634 vss.n245 vss.n241 25.6005
R1635 vss.n304 vss.n301 25.6005
R1636 vss.n308 vss.n306 25.6005
R1637 vss.n310 vss.n308 25.6005
R1638 vss.n312 vss.n310 25.6005
R1639 vss.n314 vss.n312 25.6005
R1640 vss.n316 vss.n314 25.6005
R1641 vss.n318 vss.n316 25.6005
R1642 vss.n320 vss.n318 25.6005
R1643 vss.n322 vss.n320 25.6005
R1644 vss.n324 vss.n322 25.6005
R1645 vss.n326 vss.n324 25.6005
R1646 vss.n328 vss.n326 25.6005
R1647 vss.n330 vss.n328 25.6005
R1648 vss.n332 vss.n330 25.6005
R1649 vss.n334 vss.n332 25.6005
R1650 vss.n336 vss.n334 25.6005
R1651 vss.n338 vss.n336 25.6005
R1652 vss.n340 vss.n338 25.6005
R1653 vss.n413 vss.n410 25.6005
R1654 vss.n416 vss.n413 25.6005
R1655 vss.n419 vss.n416 25.6005
R1656 vss.n422 vss.n419 25.6005
R1657 vss.n425 vss.n422 25.6005
R1658 vss.n428 vss.n425 25.6005
R1659 vss.n431 vss.n428 25.6005
R1660 vss.n434 vss.n431 25.6005
R1661 vss.n437 vss.n434 25.6005
R1662 vss.n440 vss.n437 25.6005
R1663 vss.n443 vss.n440 25.6005
R1664 vss.n446 vss.n443 25.6005
R1665 vss.n449 vss.n446 25.6005
R1666 vss.n452 vss.n449 25.6005
R1667 vss.n455 vss.n452 25.6005
R1668 vss.n458 vss.n455 25.6005
R1669 vss.n460 vss.n458 25.6005
R1670 vss.n407 vss.n403 25.6005
R1671 vss.n466 vss.n463 25.6005
R1672 vss.n470 vss.n468 25.6005
R1673 vss.n472 vss.n470 25.6005
R1674 vss.n474 vss.n472 25.6005
R1675 vss.n476 vss.n474 25.6005
R1676 vss.n478 vss.n476 25.6005
R1677 vss.n480 vss.n478 25.6005
R1678 vss.n482 vss.n480 25.6005
R1679 vss.n484 vss.n482 25.6005
R1680 vss.n486 vss.n484 25.6005
R1681 vss.n488 vss.n486 25.6005
R1682 vss.n490 vss.n488 25.6005
R1683 vss.n492 vss.n490 25.6005
R1684 vss.n494 vss.n492 25.6005
R1685 vss.n496 vss.n494 25.6005
R1686 vss.n498 vss.n496 25.6005
R1687 vss.n500 vss.n498 25.6005
R1688 vss.n502 vss.n500 25.6005
R1689 vss.n575 vss.n572 25.6005
R1690 vss.n578 vss.n575 25.6005
R1691 vss.n581 vss.n578 25.6005
R1692 vss.n584 vss.n581 25.6005
R1693 vss.n587 vss.n584 25.6005
R1694 vss.n590 vss.n587 25.6005
R1695 vss.n593 vss.n590 25.6005
R1696 vss.n596 vss.n593 25.6005
R1697 vss.n599 vss.n596 25.6005
R1698 vss.n602 vss.n599 25.6005
R1699 vss.n605 vss.n602 25.6005
R1700 vss.n608 vss.n605 25.6005
R1701 vss.n611 vss.n608 25.6005
R1702 vss.n614 vss.n611 25.6005
R1703 vss.n617 vss.n614 25.6005
R1704 vss.n620 vss.n617 25.6005
R1705 vss.n622 vss.n620 25.6005
R1706 vss.n569 vss.n565 25.6005
R1707 vss.n628 vss.n625 25.6005
R1708 vss.n632 vss.n630 25.6005
R1709 vss.n634 vss.n632 25.6005
R1710 vss.n636 vss.n634 25.6005
R1711 vss.n638 vss.n636 25.6005
R1712 vss.n640 vss.n638 25.6005
R1713 vss.n642 vss.n640 25.6005
R1714 vss.n644 vss.n642 25.6005
R1715 vss.n646 vss.n644 25.6005
R1716 vss.n648 vss.n646 25.6005
R1717 vss.n650 vss.n648 25.6005
R1718 vss.n652 vss.n650 25.6005
R1719 vss.n654 vss.n652 25.6005
R1720 vss.n656 vss.n654 25.6005
R1721 vss.n658 vss.n656 25.6005
R1722 vss.n660 vss.n658 25.6005
R1723 vss.n662 vss.n660 25.6005
R1724 vss.n664 vss.n662 25.6005
R1725 vss.n218 vss.n217 24.962
R1726 vss.n380 vss.n379 24.962
R1727 vss.n542 vss.n541 24.962
R1728 vss.n704 vss.n703 24.962
R1729 vss.n705 vss.n704 24.962
R1730 vss.n543 vss.n542 24.962
R1731 vss.n381 vss.n380 24.962
R1732 vss.n219 vss.n218 24.962
R1733 vss.n906 vss.t97 24.9236
R1734 vss.n906 vss.t93 24.9236
R1735 vss.n895 vss.t152 24.9236
R1736 vss.n895 vss.t148 24.9236
R1737 vss.n848 vss.t115 24.9236
R1738 vss.n848 vss.t111 24.9236
R1739 vss.n837 vss.t71 24.9236
R1740 vss.n837 vss.t69 24.9236
R1741 vss.n790 vss.t105 24.9236
R1742 vss.n790 vss.t95 24.9236
R1743 vss.n779 vss.t50 24.9236
R1744 vss.n779 vss.t47 24.9236
R1745 vss.n732 vss.t109 24.9236
R1746 vss.n732 vss.t113 24.9236
R1747 vss.n721 vss.t85 24.9236
R1748 vss.n721 vss.t119 24.9236
R1749 vss.n196 vss.n195 23.177
R1750 vss.n358 vss.n357 23.177
R1751 vss.n520 vss.n519 23.177
R1752 vss.n682 vss.n681 23.177
R1753 vss.n876 vss.n873 16.1455
R1754 vss.n818 vss.n815 16.1455
R1755 vss.n760 vss.n757 16.1455
R1756 vss.n672 vss.n668 11.1897
R1757 vss.n510 vss.n506 11.1897
R1758 vss.n348 vss.n344 11.1897
R1759 vss.n186 vss.n105 11.1897
R1760 vss.n200 vss.n199 9.3005
R1761 vss.n212 vss.n211 9.3005
R1762 vss.n225 vss.n60 9.3005
R1763 vss.n202 vss.n201 9.3005
R1764 vss.n214 vss.n213 9.3005
R1765 vss.n224 vss.n223 9.3005
R1766 vss.n362 vss.n361 9.3005
R1767 vss.n374 vss.n373 9.3005
R1768 vss.n387 vss.n299 9.3005
R1769 vss.n364 vss.n363 9.3005
R1770 vss.n376 vss.n375 9.3005
R1771 vss.n386 vss.n385 9.3005
R1772 vss.n524 vss.n523 9.3005
R1773 vss.n536 vss.n535 9.3005
R1774 vss.n549 vss.n461 9.3005
R1775 vss.n526 vss.n525 9.3005
R1776 vss.n538 vss.n537 9.3005
R1777 vss.n548 vss.n547 9.3005
R1778 vss.n686 vss.n685 9.3005
R1779 vss.n698 vss.n697 9.3005
R1780 vss.n711 vss.n623 9.3005
R1781 vss.n688 vss.n687 9.3005
R1782 vss.n700 vss.n699 9.3005
R1783 vss.n710 vss.n709 9.3005
R1784 vss.n684 vss.n683 9.3005
R1785 vss.n683 vss.n682 9.3005
R1786 vss.n696 vss.n695 9.3005
R1787 vss.n695 vss.n694 9.3005
R1788 vss.n674 vss.n673 9.3005
R1789 vss.n708 vss.n707 9.3005
R1790 vss.n707 vss.n706 9.3005
R1791 vss.n522 vss.n521 9.3005
R1792 vss.n521 vss.n520 9.3005
R1793 vss.n534 vss.n533 9.3005
R1794 vss.n533 vss.n532 9.3005
R1795 vss.n512 vss.n511 9.3005
R1796 vss.n546 vss.n545 9.3005
R1797 vss.n545 vss.n544 9.3005
R1798 vss.n360 vss.n359 9.3005
R1799 vss.n359 vss.n358 9.3005
R1800 vss.n372 vss.n371 9.3005
R1801 vss.n371 vss.n370 9.3005
R1802 vss.n350 vss.n349 9.3005
R1803 vss.n384 vss.n383 9.3005
R1804 vss.n383 vss.n382 9.3005
R1805 vss.n198 vss.n197 9.3005
R1806 vss.n197 vss.n196 9.3005
R1807 vss.n210 vss.n209 9.3005
R1808 vss.n209 vss.n208 9.3005
R1809 vss.n188 vss.n187 9.3005
R1810 vss.n222 vss.n221 9.3005
R1811 vss.n221 vss.n220 9.3005
R1812 vss.n923 vss.n922 9.3005
R1813 vss.n928 vss.n927 9.0005
R1814 vss.n672 vss.n671 8.98038
R1815 vss.n510 vss.n509 8.98038
R1816 vss.n348 vss.n347 8.98038
R1817 vss.n186 vss.n185 8.98038
R1818 vss.n180 vss.n109 6.57927
R1819 vss.n103 vss.n102 5.64756
R1820 vss.n342 vss.n341 5.64756
R1821 vss.n504 vss.n503 5.64756
R1822 vss.n666 vss.n665 5.64756
R1823 vss.n943 vss.n942 4.91351
R1824 vss.n191 vss.n190 4.89462
R1825 vss.n353 vss.n352 4.89462
R1826 vss.n515 vss.n514 4.89462
R1827 vss.n677 vss.n676 4.89462
R1828 vss.n558 vss.n557 4.85762
R1829 vss.n396 vss.n395 4.85762
R1830 vss.n234 vss.n233 4.85762
R1831 vss.n937 vss.n936 4.85762
R1832 vss.n121 vss.n120 4.6505
R1833 vss.n123 vss.n122 4.6505
R1834 vss.n127 vss.n126 4.6505
R1835 vss.n129 vss.n128 4.6505
R1836 vss.n133 vss.n132 4.6505
R1837 vss.n135 vss.n134 4.6505
R1838 vss.n139 vss.n138 4.6505
R1839 vss.n141 vss.n140 4.6505
R1840 vss.n145 vss.n144 4.6505
R1841 vss.n147 vss.n146 4.6505
R1842 vss.n151 vss.n150 4.6505
R1843 vss.n153 vss.n152 4.6505
R1844 vss.n157 vss.n156 4.6505
R1845 vss.n159 vss.n158 4.6505
R1846 vss.n163 vss.n162 4.6505
R1847 vss.n165 vss.n164 4.6505
R1848 vss.n169 vss.n168 4.6505
R1849 vss.n125 vss.n124 4.6505
R1850 vss.n131 vss.n130 4.6505
R1851 vss.n137 vss.n136 4.6505
R1852 vss.n143 vss.n142 4.6505
R1853 vss.n149 vss.n148 4.6505
R1854 vss.n155 vss.n154 4.6505
R1855 vss.n161 vss.n160 4.6505
R1856 vss.n167 vss.n166 4.6505
R1857 vss.n180 vss.n179 4.6505
R1858 vss.n119 vss.n118 4.6505
R1859 vss.n117 vss.n116 4.6505
R1860 vss.n718 vss.n717 4.6505
R1861 vss.n723 vss.n722 4.6505
R1862 vss.n727 vss.n726 4.6505
R1863 vss.n729 vss.n728 4.6505
R1864 vss.n734 vss.n733 4.6505
R1865 vss.n738 vss.n737 4.6505
R1866 vss.n776 vss.n775 4.6505
R1867 vss.n781 vss.n780 4.6505
R1868 vss.n785 vss.n784 4.6505
R1869 vss.n787 vss.n786 4.6505
R1870 vss.n792 vss.n791 4.6505
R1871 vss.n796 vss.n795 4.6505
R1872 vss.n834 vss.n833 4.6505
R1873 vss.n839 vss.n838 4.6505
R1874 vss.n843 vss.n842 4.6505
R1875 vss.n845 vss.n844 4.6505
R1876 vss.n850 vss.n849 4.6505
R1877 vss.n854 vss.n853 4.6505
R1878 vss.n892 vss.n891 4.6505
R1879 vss.n897 vss.n896 4.6505
R1880 vss.n901 vss.n900 4.6505
R1881 vss.n903 vss.n902 4.6505
R1882 vss.n908 vss.n907 4.6505
R1883 vss.n912 vss.n911 4.6505
R1884 vss.n941 vss.n940 4.6505
R1885 vss.n921 vss.n920 4.6505
R1886 vss.n919 vss.n918 4.6505
R1887 vss.n917 vss.n916 4.6505
R1888 vss.n890 vss.n889 4.6505
R1889 vss.n886 vss.n885 4.6505
R1890 vss.n881 vss.n880 4.6505
R1891 vss.n877 vss.n876 4.6505
R1892 vss.n873 vss.n872 4.6505
R1893 vss.n863 vss.n862 4.6505
R1894 vss.n861 vss.n860 4.6505
R1895 vss.n859 vss.n858 4.6505
R1896 vss.n832 vss.n831 4.6505
R1897 vss.n828 vss.n827 4.6505
R1898 vss.n823 vss.n822 4.6505
R1899 vss.n819 vss.n818 4.6505
R1900 vss.n815 vss.n814 4.6505
R1901 vss.n805 vss.n804 4.6505
R1902 vss.n803 vss.n802 4.6505
R1903 vss.n801 vss.n800 4.6505
R1904 vss.n774 vss.n773 4.6505
R1905 vss.n770 vss.n769 4.6505
R1906 vss.n765 vss.n764 4.6505
R1907 vss.n761 vss.n760 4.6505
R1908 vss.n757 vss.n756 4.6505
R1909 vss.n747 vss.n746 4.6505
R1910 vss.n745 vss.n744 4.6505
R1911 vss.n743 vss.n742 4.6505
R1912 vss.n716 vss.n715 4.6505
R1913 vss.n720 vss.n719 4.6505
R1914 vss.n725 vss.n724 4.6505
R1915 vss.n731 vss.n730 4.6505
R1916 vss.n736 vss.n735 4.6505
R1917 vss.n741 vss.n740 4.6505
R1918 vss.n768 vss.n767 4.6505
R1919 vss.n778 vss.n777 4.6505
R1920 vss.n783 vss.n782 4.6505
R1921 vss.n789 vss.n788 4.6505
R1922 vss.n794 vss.n793 4.6505
R1923 vss.n799 vss.n798 4.6505
R1924 vss.n826 vss.n825 4.6505
R1925 vss.n836 vss.n835 4.6505
R1926 vss.n841 vss.n840 4.6505
R1927 vss.n847 vss.n846 4.6505
R1928 vss.n852 vss.n851 4.6505
R1929 vss.n857 vss.n856 4.6505
R1930 vss.n884 vss.n883 4.6505
R1931 vss.n894 vss.n893 4.6505
R1932 vss.n899 vss.n898 4.6505
R1933 vss.n905 vss.n904 4.6505
R1934 vss.n910 vss.n909 4.6505
R1935 vss.n915 vss.n914 4.6505
R1936 vss.n929 vss.n225 4.37578
R1937 vss.n867 vss.n387 4.37578
R1938 vss.n809 vss.n549 4.37578
R1939 vss.n751 vss.n711 4.37578
R1940 vss.n204 vss.n203 4.14168
R1941 vss.n366 vss.n365 4.14168
R1942 vss.n528 vss.n527 4.14168
R1943 vss.n690 vss.n689 4.14168
R1944 vss.n216 vss.n215 3.38874
R1945 vss.n378 vss.n377 3.38874
R1946 vss.n540 vss.n539 3.38874
R1947 vss.n702 vss.n701 3.38874
R1948 vss.n230 vss.n229 3.37584
R1949 vss.n392 vss.n391 3.37584
R1950 vss.n554 vss.n553 3.37584
R1951 vss.n940 vss.n938 3.2005
R1952 vss.n236 vss.n235 3.2005
R1953 vss.n398 vss.n397 3.2005
R1954 vss.n560 vss.n559 3.2005
R1955 vss.n196 vss.n192 3.16936
R1956 vss.n358 vss.n354 3.16936
R1957 vss.n520 vss.n516 3.16936
R1958 vss.n682 vss.n678 3.16936
R1959 vss.n221 vss.n216 3.01226
R1960 vss.n383 vss.n378 3.01226
R1961 vss.n545 vss.n540 3.01226
R1962 vss.n707 vss.n702 3.01226
R1963 vss.n238 vss.n237 2.63064
R1964 vss.n400 vss.n399 2.63064
R1965 vss.n562 vss.n561 2.63064
R1966 vss vss.n951 2.60076
R1967 vss.n198 vss.n189 2.26191
R1968 vss.n360 vss.n351 2.26191
R1969 vss.n522 vss.n513 2.26191
R1970 vss.n684 vss.n675 2.26191
R1971 vss.n209 vss.n204 2.25932
R1972 vss.n371 vss.n366 2.25932
R1973 vss.n533 vss.n528 2.25932
R1974 vss.n695 vss.n690 2.25932
R1975 vss.n115 vss.n114 1.91313
R1976 vss.n189 vss.n188 1.73128
R1977 vss.n351 vss.n350 1.73128
R1978 vss.n513 vss.n512 1.73128
R1979 vss.n675 vss.n674 1.73128
R1980 vss.n716 vss.n712 1.64549
R1981 vss.n117 vss.n115 1.50714
R1982 vss.n197 vss.n191 1.50638
R1983 vss.n359 vss.n353 1.50638
R1984 vss.n521 vss.n515 1.50638
R1985 vss.n683 vss.n677 1.50638
R1986 vss.n888 vss.n887 1.18311
R1987 vss.n830 vss.n829 1.18311
R1988 vss.n772 vss.n771 1.18311
R1989 vss.n714 vss.n713 1.18311
R1990 vss.n940 vss.n939 1.14023
R1991 vss.n237 vss.n236 1.14023
R1992 vss.n399 vss.n398 1.14023
R1993 vss.n561 vss.n560 1.14023
R1994 vss.n188 vss.n103 0.753441
R1995 vss.n350 vss.n342 0.753441
R1996 vss.n512 vss.n504 0.753441
R1997 vss.n674 vss.n666 0.753441
R1998 vss.n179 vss.n178 0.747896
R1999 vss.n178 vss.n176 0.69215
R2000 vss.n951 vss.n950 0.691743
R2001 vss.n227 vss.n226 0.658034
R2002 vss.n389 vss.n388 0.658034
R2003 vss.n551 vss.n550 0.658034
R2004 vss.n935 vss.n934 0.614199
R2005 vss.n232 vss.n231 0.614199
R2006 vss.n394 vss.n393 0.614199
R2007 vss.n556 vss.n555 0.614199
R2008 vss.n208 vss.n207 0.514956
R2009 vss.n370 vss.n369 0.514956
R2010 vss.n532 vss.n531 0.514956
R2011 vss.n694 vss.n693 0.514956
R2012 vss.n927 vss.n926 0.438856
R2013 vss.n229 vss.n228 0.438856
R2014 vss.n391 vss.n390 0.438856
R2015 vss.n553 vss.n552 0.438856
R2016 vss.n883 vss.n882 0.417891
R2017 vss.n889 vss.n888 0.417891
R2018 vss.n825 vss.n824 0.417891
R2019 vss.n831 vss.n830 0.417891
R2020 vss.n767 vss.n766 0.417891
R2021 vss.n773 vss.n772 0.417891
R2022 vss.n715 vss.n714 0.417891
R2023 vss.n914 vss.n913 0.409011
R2024 vss.n856 vss.n855 0.409011
R2025 vss.n798 vss.n797 0.409011
R2026 vss.n740 vss.n739 0.409011
R2027 vss.n873 vss.n238 0.263514
R2028 vss.n815 vss.n400 0.263514
R2029 vss.n757 vss.n562 0.263514
R2030 vss.n938 vss.n935 0.219678
R2031 vss.n235 vss.n232 0.219678
R2032 vss.n397 vss.n394 0.219678
R2033 vss.n559 vss.n556 0.219678
R2034 vss.n187 vss.n186 0.178872
R2035 vss.n349 vss.n348 0.178872
R2036 vss.n511 vss.n510 0.178872
R2037 vss.n673 vss.n672 0.178872
R2038 vss.n222 vss.n214 0.144522
R2039 vss.n210 vss.n202 0.144522
R2040 vss.n384 vss.n376 0.144522
R2041 vss.n372 vss.n364 0.144522
R2042 vss.n546 vss.n538 0.144522
R2043 vss.n534 vss.n526 0.144522
R2044 vss.n708 vss.n700 0.144522
R2045 vss.n696 vss.n688 0.144522
R2046 vss.n934 vss.n933 0.132007
R2047 vss.n231 vss.n230 0.132007
R2048 vss.n393 vss.n392 0.132007
R2049 vss.n555 vss.n554 0.132007
R2050 vss.n119 vss.n117 0.120292
R2051 vss.n121 vss.n119 0.120292
R2052 vss.n123 vss.n121 0.120292
R2053 vss.n125 vss.n123 0.120292
R2054 vss.n127 vss.n125 0.120292
R2055 vss.n129 vss.n127 0.120292
R2056 vss.n131 vss.n129 0.120292
R2057 vss.n133 vss.n131 0.120292
R2058 vss.n135 vss.n133 0.120292
R2059 vss.n137 vss.n135 0.120292
R2060 vss.n139 vss.n137 0.120292
R2061 vss.n141 vss.n139 0.120292
R2062 vss.n143 vss.n141 0.120292
R2063 vss.n145 vss.n143 0.120292
R2064 vss.n147 vss.n145 0.120292
R2065 vss.n149 vss.n147 0.120292
R2066 vss.n151 vss.n149 0.120292
R2067 vss.n153 vss.n151 0.120292
R2068 vss.n155 vss.n153 0.120292
R2069 vss.n157 vss.n155 0.120292
R2070 vss.n159 vss.n157 0.120292
R2071 vss.n161 vss.n159 0.120292
R2072 vss.n163 vss.n161 0.120292
R2073 vss.n165 vss.n163 0.120292
R2074 vss.n167 vss.n165 0.120292
R2075 vss.n169 vss.n167 0.120292
R2076 vss.n170 vss.n169 0.120292
R2077 vss.n179 vss.n170 0.120292
R2078 vss.n718 vss.n716 0.120292
R2079 vss.n720 vss.n718 0.120292
R2080 vss.n723 vss.n720 0.120292
R2081 vss.n725 vss.n723 0.120292
R2082 vss.n727 vss.n725 0.120292
R2083 vss.n729 vss.n727 0.120292
R2084 vss.n731 vss.n729 0.120292
R2085 vss.n734 vss.n731 0.120292
R2086 vss.n736 vss.n734 0.120292
R2087 vss.n738 vss.n736 0.120292
R2088 vss.n741 vss.n738 0.120292
R2089 vss.n743 vss.n741 0.120292
R2090 vss.n745 vss.n743 0.120292
R2091 vss.n747 vss.n745 0.120292
R2092 vss.n756 vss.n755 0.120292
R2093 vss.n765 vss.n761 0.120292
R2094 vss.n768 vss.n765 0.120292
R2095 vss.n770 vss.n768 0.120292
R2096 vss.n774 vss.n770 0.120292
R2097 vss.n776 vss.n774 0.120292
R2098 vss.n778 vss.n776 0.120292
R2099 vss.n781 vss.n778 0.120292
R2100 vss.n783 vss.n781 0.120292
R2101 vss.n785 vss.n783 0.120292
R2102 vss.n787 vss.n785 0.120292
R2103 vss.n789 vss.n787 0.120292
R2104 vss.n792 vss.n789 0.120292
R2105 vss.n794 vss.n792 0.120292
R2106 vss.n796 vss.n794 0.120292
R2107 vss.n799 vss.n796 0.120292
R2108 vss.n801 vss.n799 0.120292
R2109 vss.n803 vss.n801 0.120292
R2110 vss.n805 vss.n803 0.120292
R2111 vss.n814 vss.n813 0.120292
R2112 vss.n823 vss.n819 0.120292
R2113 vss.n826 vss.n823 0.120292
R2114 vss.n828 vss.n826 0.120292
R2115 vss.n832 vss.n828 0.120292
R2116 vss.n834 vss.n832 0.120292
R2117 vss.n836 vss.n834 0.120292
R2118 vss.n839 vss.n836 0.120292
R2119 vss.n841 vss.n839 0.120292
R2120 vss.n843 vss.n841 0.120292
R2121 vss.n845 vss.n843 0.120292
R2122 vss.n847 vss.n845 0.120292
R2123 vss.n850 vss.n847 0.120292
R2124 vss.n852 vss.n850 0.120292
R2125 vss.n854 vss.n852 0.120292
R2126 vss.n857 vss.n854 0.120292
R2127 vss.n859 vss.n857 0.120292
R2128 vss.n861 vss.n859 0.120292
R2129 vss.n863 vss.n861 0.120292
R2130 vss.n872 vss.n871 0.120292
R2131 vss.n881 vss.n877 0.120292
R2132 vss.n884 vss.n881 0.120292
R2133 vss.n886 vss.n884 0.120292
R2134 vss.n890 vss.n886 0.120292
R2135 vss.n892 vss.n890 0.120292
R2136 vss.n894 vss.n892 0.120292
R2137 vss.n897 vss.n894 0.120292
R2138 vss.n899 vss.n897 0.120292
R2139 vss.n901 vss.n899 0.120292
R2140 vss.n903 vss.n901 0.120292
R2141 vss.n905 vss.n903 0.120292
R2142 vss.n908 vss.n905 0.120292
R2143 vss.n910 vss.n908 0.120292
R2144 vss.n912 vss.n910 0.120292
R2145 vss.n915 vss.n912 0.120292
R2146 vss.n917 vss.n915 0.120292
R2147 vss.n919 vss.n917 0.120292
R2148 vss.n921 vss.n919 0.120292
R2149 vss.n943 vss.n941 0.120292
R2150 vss.n755 vss.n754 0.102062
R2151 vss.n813 vss.n812 0.102062
R2152 vss.n871 vss.n870 0.102062
R2153 vss.n941 vss.n932 0.102062
R2154 vss.n748 vss.n747 0.10076
R2155 vss.n806 vss.n805 0.10076
R2156 vss.n864 vss.n863 0.10076
R2157 vss.n923 vss.n921 0.10076
R2158 vss.n174 vss 0.0887192
R2159 vss.n927 vss.n925 0.0881712
R2160 vss.n228 vss.n227 0.0881712
R2161 vss.n390 vss.n389 0.0881712
R2162 vss.n552 vss.n551 0.0881712
R2163 vss.n945 vss 0.075897
R2164 vss.n756 vss 0.0603958
R2165 vss.n761 vss 0.0603958
R2166 vss.n814 vss 0.0603958
R2167 vss.n819 vss 0.0603958
R2168 vss.n872 vss 0.0603958
R2169 vss.n877 vss 0.0603958
R2170 vss vss.n943 0.0603958
R2171 vss.n752 vss.n751 0.0586951
R2172 vss.n810 vss.n809 0.0586951
R2173 vss.n868 vss.n867 0.0586951
R2174 vss.n930 vss.n929 0.0586951
R2175 vss.n751 vss.n750 0.0578925
R2176 vss.n809 vss.n808 0.0578925
R2177 vss.n867 vss.n866 0.0578925
R2178 vss.n929 vss.n928 0.0578925
R2179 vss.n202 vss.n200 0.0358261
R2180 vss.n364 vss.n362 0.0358261
R2181 vss.n526 vss.n524 0.0358261
R2182 vss.n688 vss.n686 0.0358261
R2183 vss.n178 vss.n177 0.0308571
R2184 vss.n214 vss.n212 0.0303913
R2185 vss.n376 vss.n374 0.0303913
R2186 vss.n538 vss.n536 0.0303913
R2187 vss.n700 vss.n698 0.0303913
R2188 vss.n951 vss.n944 0.0272857
R2189 vss.n225 vss.n224 0.0249565
R2190 vss.n387 vss.n386 0.0249565
R2191 vss.n549 vss.n548 0.0249565
R2192 vss.n711 vss.n710 0.0249565
R2193 vss.n950 vss.n949 0.0240572
R2194 vss.n224 vss.n222 0.0222391
R2195 vss.n386 vss.n384 0.0222391
R2196 vss.n548 vss.n546 0.0222391
R2197 vss.n710 vss.n708 0.0222391
R2198 vss.n173 vss.n172 0.0205
R2199 vss.n172 vss.n171 0.0205
R2200 vss.n948 vss.n947 0.0205
R2201 vss.n949 vss.n948 0.0205
R2202 vss.n749 vss.n748 0.0200312
R2203 vss.n807 vss.n806 0.0200312
R2204 vss.n865 vss.n864 0.0200312
R2205 vss.n924 vss.n923 0.0200312
R2206 vss.n176 vss.n173 0.0187452
R2207 vss.n754 vss.n753 0.0187292
R2208 vss.n812 vss.n811 0.0187292
R2209 vss.n870 vss.n869 0.0187292
R2210 vss.n932 vss.n931 0.0187292
R2211 vss.n212 vss.n210 0.0168043
R2212 vss.n374 vss.n372 0.0168043
R2213 vss.n536 vss.n534 0.0168043
R2214 vss.n698 vss.n696 0.0168043
R2215 vss.n950 vss.n946 0.0163636
R2216 vss.n176 vss.n175 0.0142271
R2217 vss.n175 vss.n174 0.0121722
R2218 vss.n946 vss.n945 0.011753
R2219 vss.n200 vss.n198 0.0113696
R2220 vss.n362 vss.n360 0.0113696
R2221 vss.n524 vss.n522 0.0113696
R2222 vss.n686 vss.n684 0.0113696
R2223 vss.n753 vss.n752 0.00440625
R2224 vss.n811 vss.n810 0.00440625
R2225 vss.n869 vss.n868 0.00440625
R2226 vss.n931 vss.n930 0.00440625
R2227 vss.n750 vss.n749 0.00310417
R2228 vss.n808 vss.n807 0.00310417
R2229 vss.n866 vss.n865 0.00310417
R2230 vss.n928 vss.n924 0.00310417
R2231 out.n40 out.t73 28.5655
R2232 out.n40 out.t69 28.5655
R2233 out.n36 out.t71 28.5655
R2234 out.n36 out.t75 28.5655
R2235 out.n33 out.t72 28.5655
R2236 out.n33 out.t70 28.5655
R2237 out.n44 out.t74 28.5655
R2238 out.n44 out.t76 28.5655
R2239 out.n47 out.t68 28.5655
R2240 out.n47 out.t67 28.5655
R2241 out.n85 out.t53 28.5655
R2242 out.n85 out.t56 28.5655
R2243 out.n81 out.t55 28.5655
R2244 out.n81 out.t50 28.5655
R2245 out.n78 out.t54 28.5655
R2246 out.n78 out.t58 28.5655
R2247 out.n89 out.t52 28.5655
R2248 out.n89 out.t49 28.5655
R2249 out.n92 out.t51 28.5655
R2250 out.n92 out.t57 28.5655
R2251 out.n127 out.t61 28.5655
R2252 out.n127 out.t78 28.5655
R2253 out.n123 out.t0 28.5655
R2254 out.n123 out.t1 28.5655
R2255 out.n120 out.t47 28.5655
R2256 out.n120 out.t60 28.5655
R2257 out.n131 out.t19 28.5655
R2258 out.n131 out.t77 28.5655
R2259 out.n134 out.t62 28.5655
R2260 out.n134 out.t36 28.5655
R2261 out.n12 out.t22 28.5655
R2262 out.n12 out.t14 28.5655
R2263 out.n8 out.t63 28.5655
R2264 out.n8 out.t2 28.5655
R2265 out.n5 out.t59 28.5655
R2266 out.n5 out.t21 28.5655
R2267 out.n16 out.t66 28.5655
R2268 out.n16 out.t15 28.5655
R2269 out.n19 out.t20 28.5655
R2270 out.n19 out.t65 28.5655
R2271 out.n39 out.t46 17.4005
R2272 out.n39 out.t41 17.4005
R2273 out.n35 out.t43 17.4005
R2274 out.n35 out.t45 17.4005
R2275 out.n32 out.t38 17.4005
R2276 out.n32 out.t39 17.4005
R2277 out.n43 out.t44 17.4005
R2278 out.n43 out.t40 17.4005
R2279 out.n46 out.t37 17.4005
R2280 out.n46 out.t42 17.4005
R2281 out.n84 out.t9 17.4005
R2282 out.n84 out.t11 17.4005
R2283 out.n80 out.t6 17.4005
R2284 out.n80 out.t4 17.4005
R2285 out.n77 out.t13 17.4005
R2286 out.n77 out.t7 17.4005
R2287 out.n88 out.t12 17.4005
R2288 out.n88 out.t5 17.4005
R2289 out.n91 out.t10 17.4005
R2290 out.n91 out.t8 17.4005
R2291 out.n126 out.t28 17.4005
R2292 out.n126 out.t33 17.4005
R2293 out.n122 out.t29 17.4005
R2294 out.n122 out.t26 17.4005
R2295 out.n119 out.t27 17.4005
R2296 out.n119 out.t34 17.4005
R2297 out.n130 out.t31 17.4005
R2298 out.n130 out.t30 17.4005
R2299 out.n133 out.t25 17.4005
R2300 out.n133 out.t32 17.4005
R2301 out.n11 out.t48 17.4005
R2302 out.n11 out.t35 17.4005
R2303 out.n7 out.t24 17.4005
R2304 out.n7 out.t3 17.4005
R2305 out.n4 out.t17 17.4005
R2306 out.n4 out.t64 17.4005
R2307 out.n15 out.t18 17.4005
R2308 out.n15 out.t16 17.4005
R2309 out.n18 out.t23 17.4005
R2310 out.n18 out.t79 17.4005
R2311 out.n34 out.n32 7.68987
R2312 out.n37 out.n35 7.68987
R2313 out.n79 out.n77 7.68987
R2314 out.n82 out.n80 7.68987
R2315 out.n121 out.n119 7.68987
R2316 out.n124 out.n122 7.68987
R2317 out.n6 out.n4 7.68987
R2318 out.n41 out.n39 7.68961
R2319 out.n45 out.n43 7.68961
R2320 out.n86 out.n84 7.68961
R2321 out.n90 out.n88 7.68961
R2322 out.n128 out.n126 7.68961
R2323 out.n132 out.n130 7.68961
R2324 out.n13 out.n11 7.68961
R2325 out.n9 out.n7 7.68961
R2326 out.n17 out.n15 7.68961
R2327 out.n48 out.n46 7.68881
R2328 out.n93 out.n91 7.68881
R2329 out.n135 out.n133 7.68881
R2330 out.n20 out.n18 7.68881
R2331 out.n45 out.n44 7.52122
R2332 out.n41 out.n40 7.52122
R2333 out.n90 out.n89 7.52122
R2334 out.n86 out.n85 7.52122
R2335 out.n132 out.n131 7.52122
R2336 out.n128 out.n127 7.52122
R2337 out.n9 out.n8 7.52122
R2338 out.n17 out.n16 7.52122
R2339 out.n13 out.n12 7.52122
R2340 out.n48 out.n47 7.52105
R2341 out.n93 out.n92 7.52105
R2342 out.n135 out.n134 7.52105
R2343 out.n20 out.n19 7.52105
R2344 out.n37 out.n36 7.52096
R2345 out.n34 out.n33 7.52096
R2346 out.n82 out.n81 7.52096
R2347 out.n79 out.n78 7.52096
R2348 out.n124 out.n123 7.52096
R2349 out.n121 out.n120 7.52096
R2350 out.n6 out.n5 7.52096
R2351 out.n38 out.n34 2.54543
R2352 out.n83 out.n79 2.54543
R2353 out.n125 out.n121 2.54543
R2354 out.n10 out.n6 2.54543
R2355 out.n49 out.n48 2.52846
R2356 out.n94 out.n93 2.52846
R2357 out.n136 out.n135 2.52846
R2358 out.n21 out.n20 2.52846
R2359 out.n38 out.n37 2.21834
R2360 out.n49 out.n45 2.21834
R2361 out.n42 out.n41 2.21834
R2362 out.n83 out.n82 2.21834
R2363 out.n94 out.n90 2.21834
R2364 out.n87 out.n86 2.21834
R2365 out.n125 out.n124 2.21834
R2366 out.n136 out.n132 2.21834
R2367 out.n129 out.n128 2.21834
R2368 out.n10 out.n9 2.21834
R2369 out.n21 out.n17 2.21834
R2370 out.n14 out.n13 2.21834
R2371 out.n61 out.n51 1.72892
R2372 out.n56 out.n55 1.7055
R2373 out.n105 out.n104 1.7055
R2374 out.n147 out.n146 1.7055
R2375 out.n25 out.n24 1.7055
R2376 out.n28 out.n0 1.7055
R2377 out.n143 out.n139 1.7055
R2378 out.n101 out.n97 1.7055
R2379 out.n60 out.n59 1.7055
R2380 out.n152 out.n151 1.09861
R2381 out.n110 out.n109 1.09651
R2382 out.n68 out.n67 1.09651
R2383 out out.n50 0.86925
R2384 out out.n95 0.86925
R2385 out out.n137 0.86925
R2386 out out.n22 0.86925
R2387 out.n109 out.n108 0.680902
R2388 out.n151 out.n150 0.680902
R2389 out.n161 out.n31 0.680902
R2390 out.n501 out.n500 0.6115
R2391 out.n500 out.n499 0.6115
R2392 out.n499 out.n498 0.6115
R2393 out.n498 out.n497 0.6115
R2394 out.n497 out.n496 0.6115
R2395 out.n496 out.n495 0.6115
R2396 out.n495 out.n494 0.6115
R2397 out.n494 out.n493 0.6115
R2398 out.n493 out.n492 0.6115
R2399 out.n492 out.n491 0.6115
R2400 out.n491 out.n490 0.6115
R2401 out.n490 out.n489 0.6115
R2402 out.n489 out.n488 0.6115
R2403 out.n488 out.n487 0.6115
R2404 out.n487 out.n486 0.6115
R2405 out.n486 out.n485 0.6115
R2406 out.n485 out.n484 0.6115
R2407 out.n484 out.n483 0.6115
R2408 out.n483 out.n482 0.6115
R2409 out.n482 out.n481 0.6115
R2410 out.n481 out.n480 0.6115
R2411 out.n480 out.n479 0.6115
R2412 out.n479 out.n478 0.6115
R2413 out.n478 out.n477 0.6115
R2414 out.n477 out.n476 0.6115
R2415 out.n476 out.n475 0.6115
R2416 out.n475 out.n474 0.6115
R2417 out.n474 out.n473 0.6115
R2418 out.n473 out.n472 0.6115
R2419 out.n472 out.n471 0.6115
R2420 out.n471 out.n470 0.6115
R2421 out.n470 out.n469 0.6115
R2422 out.n469 out.n468 0.6115
R2423 out out.n161 0.512552
R2424 out.n62 out.n61 0.331771
R2425 out.n42 out.n38 0.327583
R2426 out.n87 out.n83 0.327583
R2427 out.n129 out.n125 0.327583
R2428 out.n14 out.n10 0.327583
R2429 out.n459 out.t378 0.301104
R2430 out.n450 out.t242 0.301104
R2431 out.n441 out.t106 0.301104
R2432 out.n432 out.t350 0.301104
R2433 out.n423 out.t243 0.301104
R2434 out.n414 out.t107 0.301104
R2435 out.n405 out.t352 0.301104
R2436 out.n396 out.t246 0.301104
R2437 out.n387 out.t208 0.301104
R2438 out.n378 out.t410 0.301104
R2439 out.n369 out.t313 0.301104
R2440 out.n360 out.t209 0.301104
R2441 out.n351 out.t411 0.301104
R2442 out.n342 out.t314 0.301104
R2443 out.n333 out.t210 0.301104
R2444 out.n324 out.t216 0.301104
R2445 out.n315 out.t118 0.301104
R2446 out.n306 out.t366 0.301104
R2447 out.n297 out.t265 0.301104
R2448 out.n288 out.t119 0.301104
R2449 out.n279 out.t367 0.301104
R2450 out.n270 out.t266 0.301104
R2451 out.n261 out.t120 0.301104
R2452 out.n252 out.t174 0.301104
R2453 out.n243 out.t403 0.301104
R2454 out.n234 out.t272 0.301104
R2455 out.n225 out.t175 0.301104
R2456 out.n216 out.t404 0.301104
R2457 out.n207 out.t310 0.301104
R2458 out.n198 out.t176 0.301104
R2459 out.n189 out.t405 0.301104
R2460 out.n180 out.t110 0.301104
R2461 out.n171 out.t312 0.301104
R2462 out.n162 out.t207 0.301104
R2463 out.n460 out.n459 0.301104
R2464 out.n461 out.n460 0.301104
R2465 out.n462 out.n461 0.301104
R2466 out.n463 out.n462 0.301104
R2467 out.n464 out.n463 0.301104
R2468 out.n465 out.n464 0.301104
R2469 out.n466 out.n465 0.301104
R2470 out.n467 out.n466 0.301104
R2471 out.n451 out.n450 0.301104
R2472 out.n452 out.n451 0.301104
R2473 out.n453 out.n452 0.301104
R2474 out.n454 out.n453 0.301104
R2475 out.n455 out.n454 0.301104
R2476 out.n456 out.n455 0.301104
R2477 out.n457 out.n456 0.301104
R2478 out.n458 out.n457 0.301104
R2479 out.n442 out.n441 0.301104
R2480 out.n443 out.n442 0.301104
R2481 out.n444 out.n443 0.301104
R2482 out.n445 out.n444 0.301104
R2483 out.n446 out.n445 0.301104
R2484 out.n447 out.n446 0.301104
R2485 out.n448 out.n447 0.301104
R2486 out.n449 out.n448 0.301104
R2487 out.n433 out.n432 0.301104
R2488 out.n434 out.n433 0.301104
R2489 out.n435 out.n434 0.301104
R2490 out.n436 out.n435 0.301104
R2491 out.n437 out.n436 0.301104
R2492 out.n438 out.n437 0.301104
R2493 out.n439 out.n438 0.301104
R2494 out.n440 out.n439 0.301104
R2495 out.n424 out.n423 0.301104
R2496 out.n425 out.n424 0.301104
R2497 out.n426 out.n425 0.301104
R2498 out.n427 out.n426 0.301104
R2499 out.n428 out.n427 0.301104
R2500 out.n429 out.n428 0.301104
R2501 out.n430 out.n429 0.301104
R2502 out.n431 out.n430 0.301104
R2503 out.n415 out.n414 0.301104
R2504 out.n416 out.n415 0.301104
R2505 out.n417 out.n416 0.301104
R2506 out.n418 out.n417 0.301104
R2507 out.n419 out.n418 0.301104
R2508 out.n420 out.n419 0.301104
R2509 out.n421 out.n420 0.301104
R2510 out.n422 out.n421 0.301104
R2511 out.n406 out.n405 0.301104
R2512 out.n407 out.n406 0.301104
R2513 out.n408 out.n407 0.301104
R2514 out.n409 out.n408 0.301104
R2515 out.n410 out.n409 0.301104
R2516 out.n411 out.n410 0.301104
R2517 out.n412 out.n411 0.301104
R2518 out.n413 out.n412 0.301104
R2519 out.n397 out.n396 0.301104
R2520 out.n398 out.n397 0.301104
R2521 out.n399 out.n398 0.301104
R2522 out.n400 out.n399 0.301104
R2523 out.n401 out.n400 0.301104
R2524 out.n402 out.n401 0.301104
R2525 out.n403 out.n402 0.301104
R2526 out.n404 out.n403 0.301104
R2527 out.n388 out.n387 0.301104
R2528 out.n389 out.n388 0.301104
R2529 out.n390 out.n389 0.301104
R2530 out.n391 out.n390 0.301104
R2531 out.n392 out.n391 0.301104
R2532 out.n393 out.n392 0.301104
R2533 out.n394 out.n393 0.301104
R2534 out.n395 out.n394 0.301104
R2535 out.n379 out.n378 0.301104
R2536 out.n380 out.n379 0.301104
R2537 out.n381 out.n380 0.301104
R2538 out.n382 out.n381 0.301104
R2539 out.n383 out.n382 0.301104
R2540 out.n384 out.n383 0.301104
R2541 out.n385 out.n384 0.301104
R2542 out.n386 out.n385 0.301104
R2543 out.n370 out.n369 0.301104
R2544 out.n371 out.n370 0.301104
R2545 out.n372 out.n371 0.301104
R2546 out.n373 out.n372 0.301104
R2547 out.n374 out.n373 0.301104
R2548 out.n375 out.n374 0.301104
R2549 out.n376 out.n375 0.301104
R2550 out.n377 out.n376 0.301104
R2551 out.n361 out.n360 0.301104
R2552 out.n362 out.n361 0.301104
R2553 out.n363 out.n362 0.301104
R2554 out.n364 out.n363 0.301104
R2555 out.n365 out.n364 0.301104
R2556 out.n366 out.n365 0.301104
R2557 out.n367 out.n366 0.301104
R2558 out.n368 out.n367 0.301104
R2559 out.n352 out.n351 0.301104
R2560 out.n353 out.n352 0.301104
R2561 out.n354 out.n353 0.301104
R2562 out.n355 out.n354 0.301104
R2563 out.n356 out.n355 0.301104
R2564 out.n357 out.n356 0.301104
R2565 out.n358 out.n357 0.301104
R2566 out.n359 out.n358 0.301104
R2567 out.n343 out.n342 0.301104
R2568 out.n344 out.n343 0.301104
R2569 out.n345 out.n344 0.301104
R2570 out.n346 out.n345 0.301104
R2571 out.n347 out.n346 0.301104
R2572 out.n348 out.n347 0.301104
R2573 out.n349 out.n348 0.301104
R2574 out.n350 out.n349 0.301104
R2575 out.n334 out.n333 0.301104
R2576 out.n335 out.n334 0.301104
R2577 out.n336 out.n335 0.301104
R2578 out.n337 out.n336 0.301104
R2579 out.n338 out.n337 0.301104
R2580 out.n339 out.n338 0.301104
R2581 out.n340 out.n339 0.301104
R2582 out.n341 out.n340 0.301104
R2583 out.n325 out.n324 0.301104
R2584 out.n326 out.n325 0.301104
R2585 out.n327 out.n326 0.301104
R2586 out.n328 out.n327 0.301104
R2587 out.n329 out.n328 0.301104
R2588 out.n330 out.n329 0.301104
R2589 out.n331 out.n330 0.301104
R2590 out.n332 out.n331 0.301104
R2591 out.n316 out.n315 0.301104
R2592 out.n317 out.n316 0.301104
R2593 out.n318 out.n317 0.301104
R2594 out.n319 out.n318 0.301104
R2595 out.n320 out.n319 0.301104
R2596 out.n321 out.n320 0.301104
R2597 out.n322 out.n321 0.301104
R2598 out.n323 out.n322 0.301104
R2599 out.n307 out.n306 0.301104
R2600 out.n308 out.n307 0.301104
R2601 out.n309 out.n308 0.301104
R2602 out.n310 out.n309 0.301104
R2603 out.n311 out.n310 0.301104
R2604 out.n312 out.n311 0.301104
R2605 out.n313 out.n312 0.301104
R2606 out.n314 out.n313 0.301104
R2607 out.n298 out.n297 0.301104
R2608 out.n299 out.n298 0.301104
R2609 out.n300 out.n299 0.301104
R2610 out.n301 out.n300 0.301104
R2611 out.n302 out.n301 0.301104
R2612 out.n303 out.n302 0.301104
R2613 out.n304 out.n303 0.301104
R2614 out.n305 out.n304 0.301104
R2615 out.n289 out.n288 0.301104
R2616 out.n290 out.n289 0.301104
R2617 out.n291 out.n290 0.301104
R2618 out.n292 out.n291 0.301104
R2619 out.n293 out.n292 0.301104
R2620 out.n294 out.n293 0.301104
R2621 out.n295 out.n294 0.301104
R2622 out.n296 out.n295 0.301104
R2623 out.n280 out.n279 0.301104
R2624 out.n281 out.n280 0.301104
R2625 out.n282 out.n281 0.301104
R2626 out.n283 out.n282 0.301104
R2627 out.n284 out.n283 0.301104
R2628 out.n285 out.n284 0.301104
R2629 out.n286 out.n285 0.301104
R2630 out.n287 out.n286 0.301104
R2631 out.n271 out.n270 0.301104
R2632 out.n272 out.n271 0.301104
R2633 out.n273 out.n272 0.301104
R2634 out.n274 out.n273 0.301104
R2635 out.n275 out.n274 0.301104
R2636 out.n276 out.n275 0.301104
R2637 out.n277 out.n276 0.301104
R2638 out.n278 out.n277 0.301104
R2639 out.n262 out.n261 0.301104
R2640 out.n263 out.n262 0.301104
R2641 out.n264 out.n263 0.301104
R2642 out.n265 out.n264 0.301104
R2643 out.n266 out.n265 0.301104
R2644 out.n267 out.n266 0.301104
R2645 out.n268 out.n267 0.301104
R2646 out.n269 out.n268 0.301104
R2647 out.n253 out.n252 0.301104
R2648 out.n254 out.n253 0.301104
R2649 out.n255 out.n254 0.301104
R2650 out.n256 out.n255 0.301104
R2651 out.n257 out.n256 0.301104
R2652 out.n258 out.n257 0.301104
R2653 out.n259 out.n258 0.301104
R2654 out.n260 out.n259 0.301104
R2655 out.n244 out.n243 0.301104
R2656 out.n245 out.n244 0.301104
R2657 out.n246 out.n245 0.301104
R2658 out.n247 out.n246 0.301104
R2659 out.n248 out.n247 0.301104
R2660 out.n249 out.n248 0.301104
R2661 out.n250 out.n249 0.301104
R2662 out.n251 out.n250 0.301104
R2663 out.n235 out.n234 0.301104
R2664 out.n236 out.n235 0.301104
R2665 out.n237 out.n236 0.301104
R2666 out.n238 out.n237 0.301104
R2667 out.n239 out.n238 0.301104
R2668 out.n240 out.n239 0.301104
R2669 out.n241 out.n240 0.301104
R2670 out.n242 out.n241 0.301104
R2671 out.n226 out.n225 0.301104
R2672 out.n227 out.n226 0.301104
R2673 out.n228 out.n227 0.301104
R2674 out.n229 out.n228 0.301104
R2675 out.n230 out.n229 0.301104
R2676 out.n231 out.n230 0.301104
R2677 out.n232 out.n231 0.301104
R2678 out.n233 out.n232 0.301104
R2679 out.n217 out.n216 0.301104
R2680 out.n218 out.n217 0.301104
R2681 out.n219 out.n218 0.301104
R2682 out.n220 out.n219 0.301104
R2683 out.n221 out.n220 0.301104
R2684 out.n222 out.n221 0.301104
R2685 out.n223 out.n222 0.301104
R2686 out.n224 out.n223 0.301104
R2687 out.n208 out.n207 0.301104
R2688 out.n209 out.n208 0.301104
R2689 out.n210 out.n209 0.301104
R2690 out.n211 out.n210 0.301104
R2691 out.n212 out.n211 0.301104
R2692 out.n213 out.n212 0.301104
R2693 out.n214 out.n213 0.301104
R2694 out.n215 out.n214 0.301104
R2695 out.n199 out.n198 0.301104
R2696 out.n200 out.n199 0.301104
R2697 out.n201 out.n200 0.301104
R2698 out.n202 out.n201 0.301104
R2699 out.n203 out.n202 0.301104
R2700 out.n204 out.n203 0.301104
R2701 out.n205 out.n204 0.301104
R2702 out.n206 out.n205 0.301104
R2703 out.n190 out.n189 0.301104
R2704 out.n191 out.n190 0.301104
R2705 out.n192 out.n191 0.301104
R2706 out.n193 out.n192 0.301104
R2707 out.n194 out.n193 0.301104
R2708 out.n195 out.n194 0.301104
R2709 out.n196 out.n195 0.301104
R2710 out.n197 out.n196 0.301104
R2711 out.n181 out.n180 0.301104
R2712 out.n182 out.n181 0.301104
R2713 out.n183 out.n182 0.301104
R2714 out.n184 out.n183 0.301104
R2715 out.n185 out.n184 0.301104
R2716 out.n186 out.n185 0.301104
R2717 out.n187 out.n186 0.301104
R2718 out.n188 out.n187 0.301104
R2719 out.n172 out.n171 0.301104
R2720 out.n173 out.n172 0.301104
R2721 out.n174 out.n173 0.301104
R2722 out.n175 out.n174 0.301104
R2723 out.n176 out.n175 0.301104
R2724 out.n177 out.n176 0.301104
R2725 out.n178 out.n177 0.301104
R2726 out.n179 out.n178 0.301104
R2727 out.n163 out.n162 0.301104
R2728 out.n164 out.n163 0.301104
R2729 out.n165 out.n164 0.301104
R2730 out.n166 out.n165 0.301104
R2731 out.n167 out.n166 0.301104
R2732 out.n168 out.n167 0.301104
R2733 out.n169 out.n168 0.301104
R2734 out.n170 out.n169 0.301104
R2735 out.n50 out.n49 0.297375
R2736 out.n95 out.n94 0.297375
R2737 out.n137 out.n136 0.297375
R2738 out.n22 out.n21 0.297375
R2739 out out.n501 0.165
R2740 out.n468 out.n467 0.14101
R2741 out.n469 out.n458 0.14101
R2742 out.n470 out.n449 0.14101
R2743 out.n471 out.n440 0.14101
R2744 out.n472 out.n431 0.14101
R2745 out.n473 out.n422 0.14101
R2746 out.n474 out.n413 0.14101
R2747 out.n475 out.n404 0.14101
R2748 out.n476 out.n395 0.14101
R2749 out.n477 out.n386 0.14101
R2750 out.n478 out.n377 0.14101
R2751 out.n479 out.n368 0.14101
R2752 out.n480 out.n359 0.14101
R2753 out.n481 out.n350 0.14101
R2754 out.n482 out.n341 0.14101
R2755 out.n483 out.n332 0.14101
R2756 out.n484 out.n323 0.14101
R2757 out.n485 out.n314 0.14101
R2758 out.n486 out.n305 0.14101
R2759 out.n487 out.n296 0.14101
R2760 out.n488 out.n287 0.14101
R2761 out.n489 out.n278 0.14101
R2762 out.n490 out.n269 0.14101
R2763 out.n491 out.n260 0.14101
R2764 out.n492 out.n251 0.14101
R2765 out.n493 out.n242 0.14101
R2766 out.n494 out.n233 0.14101
R2767 out.n495 out.n224 0.14101
R2768 out.n496 out.n215 0.14101
R2769 out.n497 out.n206 0.14101
R2770 out.n498 out.n197 0.14101
R2771 out.n499 out.n188 0.14101
R2772 out.n500 out.n179 0.14101
R2773 out.n501 out.n170 0.14101
R2774 out.n51 out 0.0505
R2775 out.n96 out 0.0505
R2776 out.n138 out 0.0505
R2777 out.n23 out 0.0505
R2778 out.n97 out.n96 0.03175
R2779 out.n139 out.n138 0.03175
R2780 out.n24 out.n23 0.03175
R2781 out.n61 out.n60 0.025645
R2782 out.n468 out 0.02306
R2783 out.n153 out.n152 0.023016
R2784 out.n161 out.n160 0.0221211
R2785 out.n111 out.n110 0.0221211
R2786 out.n69 out.n68 0.0221211
R2787 out.n151 out.n118 0.0221211
R2788 out.n109 out.n76 0.0221211
R2789 out.n67 out.n66 0.0221211
R2790 out.n53 out.n52 0.018125
R2791 out.n56 out.n54 0.018125
R2792 out.n57 out.n56 0.018125
R2793 out.n60 out.n58 0.018125
R2794 out.n108 out.n107 0.018125
R2795 out.n106 out.n105 0.018125
R2796 out.n105 out.n103 0.018125
R2797 out.n102 out.n101 0.018125
R2798 out.n101 out.n100 0.018125
R2799 out.n99 out.n98 0.018125
R2800 out.n150 out.n149 0.018125
R2801 out.n148 out.n147 0.018125
R2802 out.n147 out.n145 0.018125
R2803 out.n144 out.n143 0.018125
R2804 out.n143 out.n142 0.018125
R2805 out.n141 out.n140 0.018125
R2806 out.n31 out.n30 0.018125
R2807 out.n29 out.n28 0.018125
R2808 out.n28 out.n27 0.018125
R2809 out.n26 out.n25 0.018125
R2810 out.n25 out.n3 0.018125
R2811 out.n2 out.n1 0.018125
R2812 out.n159 out.n158 0.018125
R2813 out.n158 out.n157 0.018125
R2814 out.n156 out.n155 0.018125
R2815 out.n155 out.n154 0.018125
R2816 out.n117 out.n116 0.018125
R2817 out.n116 out.n115 0.018125
R2818 out.n114 out.n113 0.018125
R2819 out.n113 out.n112 0.018125
R2820 out.n75 out.n74 0.018125
R2821 out.n74 out.n73 0.018125
R2822 out.n72 out.n71 0.018125
R2823 out.n71 out.n70 0.018125
R2824 out.n65 out.n64 0.018125
R2825 out.n64 out.n63 0.018125
R2826 out.n50 out.n42 0.0171667
R2827 out.n95 out.n87 0.0171667
R2828 out.n137 out.n129 0.0171667
R2829 out.n22 out.n14 0.0171667
R2830 out.n54 out.n53 0.01225
R2831 out.n58 out.n57 0.01225
R2832 out.n107 out.n106 0.01225
R2833 out.n103 out.n102 0.01225
R2834 out.n100 out.n99 0.01225
R2835 out.n149 out.n148 0.01225
R2836 out.n145 out.n144 0.01225
R2837 out.n142 out.n141 0.01225
R2838 out.n30 out.n29 0.01225
R2839 out.n27 out.n26 0.01225
R2840 out.n3 out.n2 0.01225
R2841 out.n160 out.n159 0.01225
R2842 out.n157 out.n156 0.01225
R2843 out.n154 out.n153 0.01225
R2844 out.n118 out.n117 0.01225
R2845 out.n115 out.n114 0.01225
R2846 out.n112 out.n111 0.01225
R2847 out.n76 out.n75 0.01225
R2848 out.n73 out.n72 0.01225
R2849 out.n70 out.n69 0.01225
R2850 out.n66 out.n65 0.01225
R2851 out.n63 out.n62 0.01225
R2852 out.n459 out.t383 0.00050016
R2853 out.n460 out.t386 0.00050016
R2854 out.n461 out.t402 0.00050016
R2855 out.n462 out.t406 0.00050016
R2856 out.n463 out.t252 0.00050016
R2857 out.n464 out.t259 0.00050016
R2858 out.n465 out.t267 0.00050016
R2859 out.n466 out.t284 0.00050016
R2860 out.n467 out.t291 0.00050016
R2861 out.n450 out.t250 0.00050016
R2862 out.n451 out.t258 0.00050016
R2863 out.n452 out.t282 0.00050016
R2864 out.n453 out.t286 0.00050016
R2865 out.n454 out.t125 0.00050016
R2866 out.n455 out.t133 0.00050016
R2867 out.n456 out.t143 0.00050016
R2868 out.n457 out.t166 0.00050016
R2869 out.n458 out.t172 0.00050016
R2870 out.n441 out.t112 0.00050016
R2871 out.n442 out.t116 0.00050016
R2872 out.n443 out.t150 0.00050016
R2873 out.n444 out.t155 0.00050016
R2874 out.n445 out.t330 0.00050016
R2875 out.n446 out.t333 0.00050016
R2876 out.n447 out.t338 0.00050016
R2877 out.n448 out.t365 0.00050016
R2878 out.n449 out.t370 0.00050016
R2879 out.n432 out.t358 0.00050016
R2880 out.n433 out.t362 0.00050016
R2881 out.n434 out.t385 0.00050016
R2882 out.n435 out.t387 0.00050016
R2883 out.n436 out.t223 0.00050016
R2884 out.n437 out.t229 0.00050016
R2885 out.n438 out.t234 0.00050016
R2886 out.n439 out.t264 0.00050016
R2887 out.n440 out.t268 0.00050016
R2888 out.n423 out.t253 0.00050016
R2889 out.n424 out.t260 0.00050016
R2890 out.n425 out.t281 0.00050016
R2891 out.n426 out.t285 0.00050016
R2892 out.n427 out.t124 0.00050016
R2893 out.n428 out.t135 0.00050016
R2894 out.n429 out.t144 0.00050016
R2895 out.n430 out.t165 0.00050016
R2896 out.n431 out.t171 0.00050016
R2897 out.n414 out.t113 0.00050016
R2898 out.n415 out.t117 0.00050016
R2899 out.n416 out.t149 0.00050016
R2900 out.n417 out.t154 0.00050016
R2901 out.n418 out.t329 0.00050016
R2902 out.n419 out.t335 0.00050016
R2903 out.n420 out.t339 0.00050016
R2904 out.n421 out.t364 0.00050016
R2905 out.n422 out.t369 0.00050016
R2906 out.n405 out.t360 0.00050016
R2907 out.n406 out.t363 0.00050016
R2908 out.n407 out.t384 0.00050016
R2909 out.n408 out.t389 0.00050016
R2910 out.n409 out.t226 0.00050016
R2911 out.n410 out.t233 0.00050016
R2912 out.n411 out.t235 0.00050016
R2913 out.n412 out.t263 0.00050016
R2914 out.n413 out.t269 0.00050016
R2915 out.n396 out.t256 0.00050016
R2916 out.n397 out.t261 0.00050016
R2917 out.n398 out.t283 0.00050016
R2918 out.n399 out.t288 0.00050016
R2919 out.n400 out.t129 0.00050016
R2920 out.n401 out.t139 0.00050016
R2921 out.n402 out.t145 0.00050016
R2922 out.n403 out.t168 0.00050016
R2923 out.n404 out.t173 0.00050016
R2924 out.n387 out.t213 0.00050016
R2925 out.n388 out.t219 0.00050016
R2926 out.n389 out.t241 0.00050016
R2927 out.n390 out.t251 0.00050016
R2928 out.n391 out.t86 0.00050016
R2929 out.n392 out.t91 0.00050016
R2930 out.n393 out.t99 0.00050016
R2931 out.n394 out.t123 0.00050016
R2932 out.n395 out.t134 0.00050016
R2933 out.n378 out.t418 0.00050016
R2934 out.n379 out.t83 0.00050016
R2935 out.n380 out.t105 0.00050016
R2936 out.n381 out.t111 0.00050016
R2937 out.n382 out.t297 0.00050016
R2938 out.n383 out.t305 0.00050016
R2939 out.n384 out.t308 0.00050016
R2940 out.n385 out.t328 0.00050016
R2941 out.n386 out.t334 0.00050016
R2942 out.n369 out.t320 0.00050016
R2943 out.n370 out.t326 0.00050016
R2944 out.n371 out.t351 0.00050016
R2945 out.n372 out.t359 0.00050016
R2946 out.n373 out.t193 0.00050016
R2947 out.n374 out.t197 0.00050016
R2948 out.n375 out.t202 0.00050016
R2949 out.n376 out.t224 0.00050016
R2950 out.n377 out.t231 0.00050016
R2951 out.n360 out.t214 0.00050016
R2952 out.n361 out.t220 0.00050016
R2953 out.n362 out.t245 0.00050016
R2954 out.n363 out.t255 0.00050016
R2955 out.n364 out.t88 0.00050016
R2956 out.n365 out.t90 0.00050016
R2957 out.n366 out.t98 0.00050016
R2958 out.n367 out.t127 0.00050016
R2959 out.n368 out.t137 0.00050016
R2960 out.n351 out.t419 0.00050016
R2961 out.n352 out.t84 0.00050016
R2962 out.n353 out.t108 0.00050016
R2963 out.n354 out.t114 0.00050016
R2964 out.n355 out.t298 0.00050016
R2965 out.n356 out.t304 0.00050016
R2966 out.n357 out.t307 0.00050016
R2967 out.n358 out.t331 0.00050016
R2968 out.n359 out.t336 0.00050016
R2969 out.n342 out.t321 0.00050016
R2970 out.n343 out.t327 0.00050016
R2971 out.n344 out.t353 0.00050016
R2972 out.n345 out.t361 0.00050016
R2973 out.n346 out.t192 0.00050016
R2974 out.n347 out.t196 0.00050016
R2975 out.n348 out.t203 0.00050016
R2976 out.n349 out.t227 0.00050016
R2977 out.n350 out.t230 0.00050016
R2978 out.n333 out.t215 0.00050016
R2979 out.n334 out.t222 0.00050016
R2980 out.n335 out.t244 0.00050016
R2981 out.n336 out.t254 0.00050016
R2982 out.n337 out.t87 0.00050016
R2983 out.n338 out.t92 0.00050016
R2984 out.n339 out.t100 0.00050016
R2985 out.n340 out.t126 0.00050016
R2986 out.n341 out.t136 0.00050016
R2987 out.n324 out.t225 0.00050016
R2988 out.n325 out.t232 0.00050016
R2989 out.n326 out.t257 0.00050016
R2990 out.n327 out.t262 0.00050016
R2991 out.n328 out.t95 0.00050016
R2992 out.n329 out.t104 0.00050016
R2993 out.n330 out.t109 0.00050016
R2994 out.n331 out.t142 0.00050016
R2995 out.n332 out.t146 0.00050016
R2996 out.n315 out.t128 0.00050016
R2997 out.n316 out.t138 0.00050016
R2998 out.n317 out.t161 0.00050016
R2999 out.n318 out.t167 0.00050016
R3000 out.n319 out.t341 0.00050016
R3001 out.n320 out.t346 0.00050016
R3002 out.n321 out.t355 0.00050016
R3003 out.n322 out.t376 0.00050016
R3004 out.n323 out.t380 0.00050016
R3005 out.n306 out.t371 0.00050016
R3006 out.n307 out.t374 0.00050016
R3007 out.n308 out.t395 0.00050016
R3008 out.n309 out.t400 0.00050016
R3009 out.n310 out.t236 0.00050016
R3010 out.n311 out.t239 0.00050016
R3011 out.n312 out.t248 0.00050016
R3012 out.n313 out.t275 0.00050016
R3013 out.n314 out.t278 0.00050016
R3014 out.n297 out.t270 0.00050016
R3015 out.n298 out.t273 0.00050016
R3016 out.n299 out.t295 0.00050016
R3017 out.n300 out.t303 0.00050016
R3018 out.n301 out.t148 0.00050016
R3019 out.n302 out.t152 0.00050016
R3020 out.n303 out.t157 0.00050016
R3021 out.n304 out.t178 0.00050016
R3022 out.n305 out.t183 0.00050016
R3023 out.n288 out.t130 0.00050016
R3024 out.n289 out.t140 0.00050016
R3025 out.n290 out.t162 0.00050016
R3026 out.n291 out.t170 0.00050016
R3027 out.n292 out.t343 0.00050016
R3028 out.n293 out.t348 0.00050016
R3029 out.n294 out.t354 0.00050016
R3030 out.n295 out.t377 0.00050016
R3031 out.n296 out.t382 0.00050016
R3032 out.n279 out.t372 0.00050016
R3033 out.n280 out.t375 0.00050016
R3034 out.n281 out.t396 0.00050016
R3035 out.n282 out.t401 0.00050016
R3036 out.n283 out.t237 0.00050016
R3037 out.n284 out.t238 0.00050016
R3038 out.n285 out.t247 0.00050016
R3039 out.n286 out.t276 0.00050016
R3040 out.n287 out.t279 0.00050016
R3041 out.n270 out.t271 0.00050016
R3042 out.n271 out.t274 0.00050016
R3043 out.n272 out.t296 0.00050016
R3044 out.n273 out.t302 0.00050016
R3045 out.n274 out.t147 0.00050016
R3046 out.n275 out.t151 0.00050016
R3047 out.n276 out.t158 0.00050016
R3048 out.n277 out.t177 0.00050016
R3049 out.n278 out.t182 0.00050016
R3050 out.n261 out.t131 0.00050016
R3051 out.n262 out.t141 0.00050016
R3052 out.n263 out.t163 0.00050016
R3053 out.n264 out.t169 0.00050016
R3054 out.n265 out.t342 0.00050016
R3055 out.n266 out.t347 0.00050016
R3056 out.n267 out.t356 0.00050016
R3057 out.n268 out.t379 0.00050016
R3058 out.n269 out.t381 0.00050016
R3059 out.n252 out.t179 0.00050016
R3060 out.n253 out.t184 0.00050016
R3061 out.n254 out.t198 0.00050016
R3062 out.n255 out.t204 0.00050016
R3063 out.n256 out.t388 0.00050016
R3064 out.n257 out.t392 0.00050016
R3065 out.n258 out.t397 0.00050016
R3066 out.n259 out.t415 0.00050016
R3067 out.n260 out.t80 0.00050016
R3068 out.n243 out.t407 0.00050016
R3069 out.n244 out.t412 0.00050016
R3070 out.n245 out.t93 0.00050016
R3071 out.n246 out.t101 0.00050016
R3072 out.n247 out.t287 0.00050016
R3073 out.n248 out.t293 0.00050016
R3074 out.n249 out.t300 0.00050016
R3075 out.n250 out.t316 0.00050016
R3076 out.n251 out.t322 0.00050016
R3077 out.n234 out.t277 0.00050016
R3078 out.n235 out.t280 0.00050016
R3079 out.n236 out.t306 0.00050016
R3080 out.n237 out.t309 0.00050016
R3081 out.n238 out.t156 0.00050016
R3082 out.n239 out.t160 0.00050016
R3083 out.n240 out.t164 0.00050016
R3084 out.n241 out.t187 0.00050016
R3085 out.n242 out.t188 0.00050016
R3086 out.n225 out.t180 0.00050016
R3087 out.n226 out.t185 0.00050016
R3088 out.n227 out.t199 0.00050016
R3089 out.n228 out.t205 0.00050016
R3090 out.n229 out.t391 0.00050016
R3091 out.n230 out.t394 0.00050016
R3092 out.n231 out.t399 0.00050016
R3093 out.n232 out.t416 0.00050016
R3094 out.n233 out.t81 0.00050016
R3095 out.n216 out.t408 0.00050016
R3096 out.n217 out.t413 0.00050016
R3097 out.n218 out.t94 0.00050016
R3098 out.n219 out.t103 0.00050016
R3099 out.n220 out.t290 0.00050016
R3100 out.n221 out.t292 0.00050016
R3101 out.n222 out.t299 0.00050016
R3102 out.n223 out.t318 0.00050016
R3103 out.n224 out.t324 0.00050016
R3104 out.n207 out.t311 0.00050016
R3105 out.n208 out.t315 0.00050016
R3106 out.n209 out.t340 0.00050016
R3107 out.n210 out.t345 0.00050016
R3108 out.n211 out.t189 0.00050016
R3109 out.n212 out.t190 0.00050016
R3110 out.n213 out.t194 0.00050016
R3111 out.n214 out.t211 0.00050016
R3112 out.n215 out.t217 0.00050016
R3113 out.n198 out.t181 0.00050016
R3114 out.n199 out.t186 0.00050016
R3115 out.n200 out.t200 0.00050016
R3116 out.n201 out.t206 0.00050016
R3117 out.n202 out.t390 0.00050016
R3118 out.n203 out.t393 0.00050016
R3119 out.n204 out.t398 0.00050016
R3120 out.n205 out.t417 0.00050016
R3121 out.n206 out.t82 0.00050016
R3122 out.n189 out.t409 0.00050016
R3123 out.n190 out.t414 0.00050016
R3124 out.n191 out.t96 0.00050016
R3125 out.n192 out.t102 0.00050016
R3126 out.n193 out.t289 0.00050016
R3127 out.n194 out.t294 0.00050016
R3128 out.n195 out.t301 0.00050016
R3129 out.n196 out.t317 0.00050016
R3130 out.n197 out.t323 0.00050016
R3131 out.n180 out.t115 0.00050016
R3132 out.n181 out.t121 0.00050016
R3133 out.n182 out.t153 0.00050016
R3134 out.n183 out.t159 0.00050016
R3135 out.n184 out.t332 0.00050016
R3136 out.n185 out.t337 0.00050016
R3137 out.n186 out.t344 0.00050016
R3138 out.n187 out.t368 0.00050016
R3139 out.n188 out.t373 0.00050016
R3140 out.n171 out.t319 0.00050016
R3141 out.n172 out.t325 0.00050016
R3142 out.n173 out.t349 0.00050016
R3143 out.n174 out.t357 0.00050016
R3144 out.n175 out.t191 0.00050016
R3145 out.n176 out.t195 0.00050016
R3146 out.n177 out.t201 0.00050016
R3147 out.n178 out.t221 0.00050016
R3148 out.n179 out.t228 0.00050016
R3149 out.n162 out.t212 0.00050016
R3150 out.n163 out.t218 0.00050016
R3151 out.n164 out.t240 0.00050016
R3152 out.n165 out.t249 0.00050016
R3153 out.n166 out.t85 0.00050016
R3154 out.n167 out.t89 0.00050016
R3155 out.n168 out.t97 0.00050016
R3156 out.n169 out.t122 0.00050016
R3157 out.n170 out.t132 0.00050016
R3158 carray_0.n6.n68 carray_0.n6.n67 92.6295
R3159 carray_0.n6.n73 carray_0.n6.t1 25.6105
R3160 carray_0.n6.n67 carray_0.n6.t2 24.9236
R3161 carray_0.n6.n67 carray_0.n6.t67 24.9236
R3162 carray_0.n6.n71 carray_0.n6.t0 18.6113
R3163 carray_0.n6.n69 carray_0.n6.n68 11.8308
R3164 carray_0.n6.n74 carray_0.n6.n73 9.3005
R3165 carray_0.n6.n72 carray_0.n6.n71 7.77627
R3166 carray_0.n6.n76 carray_0.n6.n75 7.57622
R3167 carray_0.n6.n39 carray_0.n6.n30 5.84104
R3168 carray_0.n6.n14 carray_0.n6.n6 5.75627
R3169 carray_0.n6.n49 carray_0.n6.n48 3.46484
R3170 carray_0.n6.n14 carray_0.n6.n13 3.46465
R3171 carray_0.n6.n22 carray_0.n6.n21 3.46465
R3172 carray_0.n6.n30 carray_0.n6.n29 3.46465
R3173 carray_0.n6.n57 carray_0.n6.n56 3.46465
R3174 carray_0.n6.n65 carray_0.n6.n64 3.46465
R3175 carray_0.n6.n49 carray_0.n6.n39 3.05649
R3176 carray_0.n6.n57 carray_0.n6.n49 3.05623
R3177 carray_0.n6.n22 carray_0.n6.n14 3.05587
R3178 carray_0.n6.n30 carray_0.n6.n22 3.05587
R3179 carray_0.n6 carray_0.n6.n77 2.95985
R3180 carray_0.n6.n38 carray_0.n6.n37 2.6155
R3181 carray_0.n6.n65 carray_0.n6.n57 2.29212
R3182 carray_0.n6.n0 carray_0.n6.t10 2.15593
R3183 carray_0.n6.n7 carray_0.n6.t43 2.15593
R3184 carray_0.n6.n15 carray_0.n6.t29 2.15593
R3185 carray_0.n6.n23 carray_0.n6.t38 2.15593
R3186 carray_0.n6.n31 carray_0.n6.t42 2.15593
R3187 carray_0.n6.n50 carray_0.n6.t12 2.15593
R3188 carray_0.n6.n58 carray_0.n6.t11 2.15593
R3189 carray_0.n6.n40 carray_0.n6.t26 2.15593
R3190 carray_0.n6.n75 carray_0.n6.n74 1.93989
R3191 carray_0.n6.n74 carray_0.n6.n70 1.93989
R3192 carray_0.n6 carray_0.n6.n65 1.51622
R3193 carray_0.n6.n75 carray_0.n6.n66 1.35808
R3194 carray_0.n6.n70 carray_0.n6.n69 1.35808
R3195 carray_0.n6.n50 carray_0.n6.t18 1.16583
R3196 carray_0.n6.n51 carray_0.n6.t21 1.16583
R3197 carray_0.n6.n52 carray_0.n6.t25 1.16583
R3198 carray_0.n6.n53 carray_0.n6.t52 1.16583
R3199 carray_0.n6.n54 carray_0.n6.t55 1.16583
R3200 carray_0.n6.n55 carray_0.n6.t57 1.16583
R3201 carray_0.n6.n56 carray_0.n6.t60 1.16583
R3202 carray_0.n6.n58 carray_0.n6.t19 1.16583
R3203 carray_0.n6.n59 carray_0.n6.t22 1.16583
R3204 carray_0.n6.n60 carray_0.n6.t24 1.16583
R3205 carray_0.n6.n61 carray_0.n6.t51 1.16583
R3206 carray_0.n6.n62 carray_0.n6.t54 1.16583
R3207 carray_0.n6.n63 carray_0.n6.t58 1.16583
R3208 carray_0.n6.n64 carray_0.n6.t61 1.16583
R3209 carray_0.n6.n40 carray_0.n6.t32 1.16583
R3210 carray_0.n6.n41 carray_0.n6.t33 1.16583
R3211 carray_0.n6.n42 carray_0.n6.t35 1.16583
R3212 carray_0.n6.n43 carray_0.n6.t62 1.16583
R3213 carray_0.n6.n44 carray_0.n6.t63 1.16583
R3214 carray_0.n6.n48 carray_0.n6.t3 1.16583
R3215 carray_0.n6.n47 carray_0.n6.n46 1.14596
R3216 carray_0.n6.n46 carray_0.n6.n45 1.12999
R3217 carray_0.n6.n6 carray_0.n6.t59 1.10593
R3218 carray_0.n6.n5 carray_0.n6.t56 1.10593
R3219 carray_0.n6.n4 carray_0.n6.t53 1.10593
R3220 carray_0.n6.n3 carray_0.n6.t50 1.10593
R3221 carray_0.n6.n2 carray_0.n6.t23 1.10593
R3222 carray_0.n6.n1 carray_0.n6.t20 1.10593
R3223 carray_0.n6.n0 carray_0.n6.t16 1.10593
R3224 carray_0.n6.n13 carray_0.n6.t31 1.10593
R3225 carray_0.n6.n12 carray_0.n6.t30 1.10593
R3226 carray_0.n6.n11 carray_0.n6.t17 1.10593
R3227 carray_0.n6.n10 carray_0.n6.t15 1.10593
R3228 carray_0.n6.n9 carray_0.n6.t49 1.10593
R3229 carray_0.n6.n8 carray_0.n6.t48 1.10593
R3230 carray_0.n6.n7 carray_0.n6.t46 1.10593
R3231 carray_0.n6.n21 carray_0.n6.t5 1.10593
R3232 carray_0.n6.n20 carray_0.n6.t4 1.10593
R3233 carray_0.n6.n19 carray_0.n6.t65 1.10593
R3234 carray_0.n6.n18 carray_0.n6.t64 1.10593
R3235 carray_0.n6.n17 carray_0.n6.t37 1.10593
R3236 carray_0.n6.n16 carray_0.n6.t36 1.10593
R3237 carray_0.n6.n15 carray_0.n6.t34 1.10593
R3238 carray_0.n6.n29 carray_0.n6.t9 1.10593
R3239 carray_0.n6.n28 carray_0.n6.t8 1.10593
R3240 carray_0.n6.n27 carray_0.n6.t7 1.10593
R3241 carray_0.n6.n26 carray_0.n6.t6 1.10593
R3242 carray_0.n6.n25 carray_0.n6.t41 1.10593
R3243 carray_0.n6.n24 carray_0.n6.t40 1.10593
R3244 carray_0.n6.n23 carray_0.n6.t39 1.10593
R3245 carray_0.n6.n31 carray_0.n6.t44 1.10593
R3246 carray_0.n6.n32 carray_0.n6.t45 1.10593
R3247 carray_0.n6.n33 carray_0.n6.t47 1.10593
R3248 carray_0.n6.n34 carray_0.n6.t13 1.10593
R3249 carray_0.n6.n35 carray_0.n6.t14 1.10593
R3250 carray_0.n6.n36 carray_0.n6.t27 1.10593
R3251 carray_0.n6.n37 carray_0.n6.t28 1.10593
R3252 carray_0.n6.n1 carray_0.n6.n0 1.0505
R3253 carray_0.n6.n2 carray_0.n6.n1 1.0505
R3254 carray_0.n6.n3 carray_0.n6.n2 1.0505
R3255 carray_0.n6.n4 carray_0.n6.n3 1.0505
R3256 carray_0.n6.n5 carray_0.n6.n4 1.0505
R3257 carray_0.n6.n6 carray_0.n6.n5 1.0505
R3258 carray_0.n6.n8 carray_0.n6.n7 1.0505
R3259 carray_0.n6.n9 carray_0.n6.n8 1.0505
R3260 carray_0.n6.n10 carray_0.n6.n9 1.0505
R3261 carray_0.n6.n11 carray_0.n6.n10 1.0505
R3262 carray_0.n6.n12 carray_0.n6.n11 1.0505
R3263 carray_0.n6.n13 carray_0.n6.n12 1.0505
R3264 carray_0.n6.n16 carray_0.n6.n15 1.0505
R3265 carray_0.n6.n17 carray_0.n6.n16 1.0505
R3266 carray_0.n6.n18 carray_0.n6.n17 1.0505
R3267 carray_0.n6.n19 carray_0.n6.n18 1.0505
R3268 carray_0.n6.n20 carray_0.n6.n19 1.0505
R3269 carray_0.n6.n21 carray_0.n6.n20 1.0505
R3270 carray_0.n6.n24 carray_0.n6.n23 1.0505
R3271 carray_0.n6.n25 carray_0.n6.n24 1.0505
R3272 carray_0.n6.n26 carray_0.n6.n25 1.0505
R3273 carray_0.n6.n27 carray_0.n6.n26 1.0505
R3274 carray_0.n6.n28 carray_0.n6.n27 1.0505
R3275 carray_0.n6.n29 carray_0.n6.n28 1.0505
R3276 carray_0.n6.n32 carray_0.n6.n31 1.0505
R3277 carray_0.n6.n33 carray_0.n6.n32 1.0505
R3278 carray_0.n6.n34 carray_0.n6.n33 1.0505
R3279 carray_0.n6.n35 carray_0.n6.n34 1.0505
R3280 carray_0.n6.n36 carray_0.n6.n35 1.0505
R3281 carray_0.n6.n37 carray_0.n6.n36 1.0505
R3282 carray_0.n6.n51 carray_0.n6.n50 1.0505
R3283 carray_0.n6.n52 carray_0.n6.n51 1.0505
R3284 carray_0.n6.n53 carray_0.n6.n52 1.0505
R3285 carray_0.n6.n54 carray_0.n6.n53 1.0505
R3286 carray_0.n6.n55 carray_0.n6.n54 1.0505
R3287 carray_0.n6.n56 carray_0.n6.n55 1.0505
R3288 carray_0.n6.n59 carray_0.n6.n58 1.0505
R3289 carray_0.n6.n60 carray_0.n6.n59 1.0505
R3290 carray_0.n6.n61 carray_0.n6.n60 1.0505
R3291 carray_0.n6.n62 carray_0.n6.n61 1.0505
R3292 carray_0.n6.n63 carray_0.n6.n62 1.0505
R3293 carray_0.n6.n64 carray_0.n6.n63 1.0505
R3294 carray_0.n6.n41 carray_0.n6.n40 1.0505
R3295 carray_0.n6.n42 carray_0.n6.n41 1.0505
R3296 carray_0.n6.n43 carray_0.n6.n42 1.0505
R3297 carray_0.n6.n44 carray_0.n6.n43 1.0505
R3298 carray_0.n6.n47 carray_0.n6.n44 1.0505
R3299 carray_0.n6.n48 carray_0.n6.n47 1.0505
R3300 carray_0.n6.n73 carray_0.n6.n72 0.9855
R3301 carray_0.n6.n39 carray_0.n6.n38 0.849651
R3302 carray_0.n6.n38 carray_0.n6 0.0505
R3303 carray_0.n6.n77 carray_0.n6.n76 0.0333125
R3304 carray_0.n6.n46 carray_0.n6.t66 0.02118
R3305 carray_0.n5.n35 carray_0.n5.n34 92.6295
R3306 carray_0.n5.n40 carray_0.n5.t0 25.6105
R3307 carray_0.n5.n34 carray_0.n5.t2 24.9236
R3308 carray_0.n5.n34 carray_0.n5.t35 24.9236
R3309 carray_0.n5.n38 carray_0.n5.t1 18.6113
R3310 carray_0.n5.n36 carray_0.n5.n35 11.8308
R3311 carray_0.n5.n41 carray_0.n5.n40 9.3005
R3312 carray_0.n5.n39 carray_0.n5.n38 7.77627
R3313 carray_0.n5 carray_0.n5.n42 10.6365
R3314 carray_0.n5.n24 carray_0.n5.n15 7.36916
R3315 carray_0.n5.n15 carray_0.n5.n6 6.32002
R3316 carray_0.n5 carray_0.n5.n32 6.09872
R3317 carray_0.n5.n24 carray_0.n5.n23 3.26484
R3318 carray_0.n5.n32 carray_0.n5.n31 3.26465
R3319 carray_0.n5.n32 carray_0.n5.n24 3.05623
R3320 carray_0.n5.n14 carray_0.n5.n13 2.4155
R3321 carray_0.n5.n0 carray_0.n5.t20 2.15593
R3322 carray_0.n5.n7 carray_0.n5.t21 2.15593
R3323 carray_0.n5.n25 carray_0.n5.t28 2.15593
R3324 carray_0.n5.n16 carray_0.n5.t4 2.15593
R3325 carray_0.n5.n42 carray_0.n5.n41 1.93989
R3326 carray_0.n5.n41 carray_0.n5.n37 1.93989
R3327 carray_0.n5.t34 carray_0.n5.n21 1.43549
R3328 carray_0.n5.n42 carray_0.n5.n33 1.35808
R3329 carray_0.n5.n37 carray_0.n5.n36 1.35808
R3330 carray_0.n5.n25 carray_0.n5.t31 1.16583
R3331 carray_0.n5.n26 carray_0.n5.t32 1.16583
R3332 carray_0.n5.n27 carray_0.n5.t33 1.16583
R3333 carray_0.n5.n28 carray_0.n5.t16 1.16583
R3334 carray_0.n5.n29 carray_0.n5.t17 1.16583
R3335 carray_0.n5.n30 carray_0.n5.t18 1.16583
R3336 carray_0.n5.n31 carray_0.n5.t19 1.16583
R3337 carray_0.n5.n6 carray_0.n5.t13 1.10593
R3338 carray_0.n5.n5 carray_0.n5.t12 1.10593
R3339 carray_0.n5.n4 carray_0.n5.t7 1.10593
R3340 carray_0.n5.n3 carray_0.n5.t5 1.10593
R3341 carray_0.n5.n2 carray_0.n5.t25 1.10593
R3342 carray_0.n5.n1 carray_0.n5.t23 1.10593
R3343 carray_0.n5.n0 carray_0.n5.t22 1.10593
R3344 carray_0.n5.n13 carray_0.n5.t15 1.10593
R3345 carray_0.n5.n12 carray_0.n5.t14 1.10593
R3346 carray_0.n5.n11 carray_0.n5.t11 1.10593
R3347 carray_0.n5.n10 carray_0.n5.t9 1.10593
R3348 carray_0.n5.n9 carray_0.n5.t27 1.10593
R3349 carray_0.n5.n8 carray_0.n5.t26 1.10593
R3350 carray_0.n5.n7 carray_0.n5.t24 1.10593
R3351 carray_0.n5.n16 carray_0.n5.t6 1.10593
R3352 carray_0.n5.n17 carray_0.n5.t8 1.10593
R3353 carray_0.n5.n18 carray_0.n5.t10 1.10593
R3354 carray_0.n5.n19 carray_0.n5.t29 1.10593
R3355 carray_0.n5.n20 carray_0.n5.t30 1.10593
R3356 carray_0.n5.n23 carray_0.n5.t3 1.10593
R3357 carray_0.n5.n22 carray_0.n5.t34 1.08606
R3358 carray_0.n5.n1 carray_0.n5.n0 1.0505
R3359 carray_0.n5.n2 carray_0.n5.n1 1.0505
R3360 carray_0.n5.n3 carray_0.n5.n2 1.0505
R3361 carray_0.n5.n4 carray_0.n5.n3 1.0505
R3362 carray_0.n5.n5 carray_0.n5.n4 1.0505
R3363 carray_0.n5.n6 carray_0.n5.n5 1.0505
R3364 carray_0.n5.n8 carray_0.n5.n7 1.0505
R3365 carray_0.n5.n9 carray_0.n5.n8 1.0505
R3366 carray_0.n5.n10 carray_0.n5.n9 1.0505
R3367 carray_0.n5.n11 carray_0.n5.n10 1.0505
R3368 carray_0.n5.n12 carray_0.n5.n11 1.0505
R3369 carray_0.n5.n13 carray_0.n5.n12 1.0505
R3370 carray_0.n5.n26 carray_0.n5.n25 1.0505
R3371 carray_0.n5.n27 carray_0.n5.n26 1.0505
R3372 carray_0.n5.n28 carray_0.n5.n27 1.0505
R3373 carray_0.n5.n29 carray_0.n5.n28 1.0505
R3374 carray_0.n5.n30 carray_0.n5.n29 1.0505
R3375 carray_0.n5.n31 carray_0.n5.n30 1.0505
R3376 carray_0.n5.n17 carray_0.n5.n16 1.0505
R3377 carray_0.n5.n18 carray_0.n5.n17 1.0505
R3378 carray_0.n5.n19 carray_0.n5.n18 1.0505
R3379 carray_0.n5.n20 carray_0.n5.n19 1.0505
R3380 carray_0.n5.n22 carray_0.n5.n20 1.0505
R3381 carray_0.n5.n23 carray_0.n5.n22 1.0505
R3382 carray_0.n5.n40 carray_0.n5.n39 0.9855
R3383 carray_0.n5.n15 carray_0.n5.n14 0.849651
R3384 carray_0.n5.n14 carray_0.n5 0.0505
R3385 vin.n77 vin.t75 36.639
R3386 vin.n99 vin.t71 36.639
R3387 vin.n72 vin.t50 36.639
R3388 vin.n112 vin.t49 36.639
R3389 vin.n32 vin.t47 36.639
R3390 vin.n52 vin.t36 36.639
R3391 vin.n6 vin.t59 36.639
R3392 vin.n26 vin.t65 36.6387
R3393 vin.n83 vin.t68 28.5655
R3394 vin.n83 vin.t72 28.5655
R3395 vin.n87 vin.t74 28.5655
R3396 vin.n87 vin.t67 28.5655
R3397 vin.n91 vin.t70 28.5655
R3398 vin.n91 vin.t73 28.5655
R3399 vin.n95 vin.t76 28.5655
R3400 vin.n95 vin.t69 28.5655
R3401 vin.n64 vin.t53 28.5655
R3402 vin.n64 vin.t57 28.5655
R3403 vin.n67 vin.t51 28.5655
R3404 vin.n67 vin.t54 28.5655
R3405 vin.n104 vin.t56 28.5655
R3406 vin.n104 vin.t58 28.5655
R3407 vin.n108 vin.t52 28.5655
R3408 vin.n108 vin.t55 28.5655
R3409 vin.n36 vin.t60 28.5655
R3410 vin.n36 vin.t0 28.5655
R3411 vin.n40 vin.t1 28.5655
R3412 vin.n40 vin.t61 28.5655
R3413 vin.n44 vin.t78 28.5655
R3414 vin.n44 vin.t19 28.5655
R3415 vin.n48 vin.t77 28.5655
R3416 vin.n48 vin.t62 28.5655
R3417 vin.n22 vin.t15 28.5655
R3418 vin.n22 vin.t20 28.5655
R3419 vin.n18 vin.t14 28.5655
R3420 vin.n18 vin.t66 28.5655
R3421 vin.n14 vin.t2 28.5655
R3422 vin.n14 vin.t22 28.5655
R3423 vin.n10 vin.t21 28.5655
R3424 vin.n10 vin.t63 28.5655
R3425 vin.n75 vin.t40 24.4033
R3426 vin.n79 vin.t46 24.4033
R3427 vin.n61 vin.t10 24.4033
R3428 vin.n114 vin.t9 24.4033
R3429 vin.n1 vin.t28 24.4033
R3430 vin.n54 vin.t34 24.4033
R3431 vin.n28 vin.t79 24.4033
R3432 vin.n3 vin.t17 24.4033
R3433 vin.n82 vin.t43 17.4005
R3434 vin.n82 vin.t37 17.4005
R3435 vin.n86 vin.t39 17.4005
R3436 vin.n86 vin.t42 17.4005
R3437 vin.n90 vin.t45 17.4005
R3438 vin.n90 vin.t38 17.4005
R3439 vin.n94 vin.t41 17.4005
R3440 vin.n94 vin.t44 17.4005
R3441 vin.n63 vin.t13 17.4005
R3442 vin.n63 vin.t7 17.4005
R3443 vin.n66 vin.t11 17.4005
R3444 vin.n66 vin.t4 17.4005
R3445 vin.n103 vin.t6 17.4005
R3446 vin.n103 vin.t8 17.4005
R3447 vin.n107 vin.t12 17.4005
R3448 vin.n107 vin.t5 17.4005
R3449 vin.n35 vin.t30 17.4005
R3450 vin.n35 vin.t32 17.4005
R3451 vin.n39 vin.t25 17.4005
R3452 vin.n39 vin.t29 17.4005
R3453 vin.n43 vin.t33 17.4005
R3454 vin.n43 vin.t27 17.4005
R3455 vin.n47 vin.t26 17.4005
R3456 vin.n47 vin.t31 17.4005
R3457 vin.n21 vin.t16 17.4005
R3458 vin.n21 vin.t23 17.4005
R3459 vin.n17 vin.t35 17.4005
R3460 vin.n17 vin.t18 17.4005
R3461 vin.n13 vin.t3 17.4005
R3462 vin.n13 vin.t48 17.4005
R3463 vin.n9 vin.t64 17.4005
R3464 vin.n9 vin.t24 17.4005
R3465 vin.n11 vin.n10 8.14078
R3466 vin.n15 vin.n14 8.14078
R3467 vin.n19 vin.n18 8.14078
R3468 vin.n23 vin.n22 8.14078
R3469 vin.n84 vin.n83 8.14053
R3470 vin.n88 vin.n87 8.14053
R3471 vin.n92 vin.n91 8.14053
R3472 vin.n96 vin.n95 8.14053
R3473 vin.n65 vin.n64 8.14053
R3474 vin.n68 vin.n67 8.14053
R3475 vin.n105 vin.n104 8.14053
R3476 vin.n109 vin.n108 8.14053
R3477 vin.n37 vin.n36 8.14053
R3478 vin.n41 vin.n40 8.14053
R3479 vin.n45 vin.n44 8.14053
R3480 vin.n49 vin.n48 8.14053
R3481 vin.n96 vin.n94 7.07031
R3482 vin.n92 vin.n90 7.07031
R3483 vin.n88 vin.n86 7.07031
R3484 vin.n84 vin.n82 7.07031
R3485 vin.n109 vin.n107 7.07031
R3486 vin.n105 vin.n103 7.07031
R3487 vin.n68 vin.n66 7.07031
R3488 vin.n65 vin.n63 7.07031
R3489 vin.n49 vin.n47 7.07031
R3490 vin.n45 vin.n43 7.07031
R3491 vin.n41 vin.n39 7.07031
R3492 vin.n37 vin.n35 7.07031
R3493 vin.n23 vin.n21 7.07005
R3494 vin.n19 vin.n17 7.07005
R3495 vin.n15 vin.n13 7.07005
R3496 vin.n11 vin.n9 7.07005
R3497 vin.n80 vin.n79 4.5005
R3498 vin.n100 vin.n99 4.5005
R3499 vin.n76 vin.n75 4.5005
R3500 vin.n78 vin.n77 4.5005
R3501 vin.n115 vin.n114 4.5005
R3502 vin.n113 vin.n112 4.5005
R3503 vin.n62 vin.n61 4.5005
R3504 vin.n73 vin.n72 4.5005
R3505 vin.n55 vin.n54 4.5005
R3506 vin.n53 vin.n52 4.5005
R3507 vin.n2 vin.n1 4.5005
R3508 vin.n33 vin.n32 4.5005
R3509 vin.n4 vin.n3 4.5005
R3510 vin.n7 vin.n6 4.5005
R3511 vin.n27 vin.n26 4.5005
R3512 vin.n29 vin.n28 4.5005
R3513 vin.n97 vin.n96 2.21834
R3514 vin.n93 vin.n92 2.21834
R3515 vin.n89 vin.n88 2.21834
R3516 vin.n85 vin.n84 2.21834
R3517 vin.n110 vin.n109 2.21834
R3518 vin.n106 vin.n105 2.21834
R3519 vin.n69 vin.n68 2.21834
R3520 vin.n70 vin.n65 2.21834
R3521 vin.n50 vin.n49 2.21834
R3522 vin.n46 vin.n45 2.21834
R3523 vin.n42 vin.n41 2.21834
R3524 vin.n38 vin.n37 2.21834
R3525 vin.n12 vin.n11 2.21834
R3526 vin.n16 vin.n15 2.21834
R3527 vin.n20 vin.n19 2.21834
R3528 vin.n24 vin.n23 2.21834
R3529 vin.n101 vin.n100 1.71175
R3530 vin.n102 vin.n76 1.71175
R3531 vin.n102 vin.n78 1.71175
R3532 vin.n116 vin.n115 1.71175
R3533 vin.n116 vin.n113 1.71175
R3534 vin.n74 vin.n62 1.71175
R3535 vin.n74 vin.n73 1.71175
R3536 vin.n56 vin.n55 1.71175
R3537 vin.n56 vin.n53 1.71175
R3538 vin.n33 vin.n31 1.71175
R3539 vin.n7 vin.n5 1.71175
R3540 vin.n30 vin.n29 1.71175
R3541 vin.n30 vin.n27 1.71175
R3542 vin.n0 vin 1.62229
R3543 vin.n60 vin.n59 1.13247
R3544 vin.n58 vin.n0 1.13247
R3545 vin.n97 vin.n93 0.327583
R3546 vin.n93 vin.n89 0.327583
R3547 vin.n89 vin.n85 0.327583
R3548 vin.n110 vin.n106 0.327583
R3549 vin.n70 vin.n69 0.327583
R3550 vin.n50 vin.n46 0.327583
R3551 vin.n46 vin.n42 0.327583
R3552 vin.n42 vin.n38 0.327583
R3553 vin.n16 vin.n12 0.327583
R3554 vin.n20 vin.n16 0.327583
R3555 vin.n24 vin.n20 0.327583
R3556 vin.n98 vin.n97 0.285917
R3557 vin.n85 vin.n81 0.285917
R3558 vin.n111 vin.n110 0.285917
R3559 vin.n71 vin.n70 0.285917
R3560 vin.n51 vin.n50 0.285917
R3561 vin.n38 vin.n34 0.285917
R3562 vin.n12 vin.n8 0.285917
R3563 vin.n25 vin.n24 0.285917
R3564 vin.n31 vin.n30 0.22845
R3565 vin.n116 vin.n102 0.22845
R3566 vin.n5 vin 0.203188
R3567 vin.n31 vin 0.203188
R3568 vin vin.n74 0.203188
R3569 vin.n102 vin 0.203188
R3570 vin.n30 vin 0.191438
R3571 vin.n56 vin 0.191438
R3572 vin vin.n116 0.191438
R3573 vin vin.n101 0.191438
R3574 vin.n74 vin.n60 0.105075
R3575 vin.n57 vin.n56 0.100375
R3576 vin.n98 vin.n80 0.041125
R3577 vin.n34 vin.n2 0.041125
R3578 vin.n8 vin.n4 0.041125
R3579 vin.n60 vin.n58 0.016595
R3580 vin.n100 vin.n98 0.009875
R3581 vin.n81 vin.n78 0.009875
R3582 vin.n113 vin.n111 0.009875
R3583 vin.n73 vin.n71 0.009875
R3584 vin.n53 vin.n51 0.009875
R3585 vin.n34 vin.n33 0.009875
R3586 vin.n8 vin.n7 0.009875
R3587 vin.n27 vin.n25 0.009875
R3588 vin.n58 vin.n57 0.00879751
R3589 enb.n24 enb.t24 212.081
R3590 enb.n22 enb.t17 212.081
R3591 enb.n18 enb.t16 212.081
R3592 enb.n16 enb.t33 212.081
R3593 enb.n14 enb.n12 146.424
R3594 enb.n11 enb.n9 144.089
R3595 enb.n0 enb.t18 143.071
R3596 enb.n8 enb.t27 142.75
R3597 enb.n0 enb.t22 142.75
R3598 enb.n1 enb.t25 142.75
R3599 enb.n2 enb.t30 142.75
R3600 enb.n3 enb.t21 142.75
R3601 enb.n4 enb.t26 142.75
R3602 enb.n5 enb.t29 142.75
R3603 enb.n6 enb.t19 142.75
R3604 enb.n7 enb.t23 142.75
R3605 enb.n24 enb.t20 139.78
R3606 enb.n22 enb.t32 139.78
R3607 enb.n18 enb.t31 139.78
R3608 enb.n16 enb.t28 139.78
R3609 enb.n11 enb.n10 107.822
R3610 enb.n14 enb.n13 107.249
R3611 enb.n20 enb.n17 97.5045
R3612 enb.n20 enb.n19 76.0005
R3613 enb.n15 enb.n11 46.6252
R3614 enb.n25 enb.n24 39.8685
R3615 enb.n17 enb.n16 30.6732
R3616 enb.n19 enb.n18 30.6732
R3617 enb.n23 enb.n22 30.6732
R3618 enb.n24 enb.n23 30.6732
R3619 enb.n13 enb.t15 26.5955
R3620 enb.n13 enb.t10 26.5955
R3621 enb.n12 enb.t12 26.5955
R3622 enb.n12 enb.t9 26.5955
R3623 enb.n9 enb.t5 24.9236
R3624 enb.n9 enb.t2 24.9236
R3625 enb.n10 enb.t0 24.9236
R3626 enb.n10 enb.t3 24.9236
R3627 enb.n21 enb.n20 21.5045
R3628 enb.n25 enb.n21 19.201
R3629 enb.n15 enb.n14 14.3512
R3630 enb.n27 enb.n8 6.80862
R3631 enb.n26 enb.n15 4.58314
R3632 enb.n27 enb.n26 2.20245
R3633 enb.n26 enb.n25 1.91723
R3634 enb.n8 enb.n7 0.321152
R3635 enb.n7 enb.n6 0.321152
R3636 enb.n6 enb.n5 0.321152
R3637 enb.n5 enb.n4 0.321152
R3638 enb.n4 enb.n3 0.321152
R3639 enb.n3 enb.n2 0.321152
R3640 enb.n2 enb.n1 0.321152
R3641 enb.n1 enb.n0 0.321152
R3642 enb enb.n27 0.063
R3643 ctl1.n0 ctl1.t2 212.081
R3644 ctl1.n1 ctl1.t0 212.081
R3645 ctl1.n0 ctl1.t3 139.78
R3646 ctl1.n1 ctl1.t1 139.78
R3647 ctl1.n1 ctl1.n0 61.346
R3648 ctl1 ctl1.n1 44.6884
R3649 carray_0.n1.n3 carray_0.n1.n2 92.6295
R3650 carray_0.n1.n8 carray_0.n1.t5 25.6105
R3651 carray_0.n1.n2 carray_0.n1.t3 24.9236
R3652 carray_0.n1.n2 carray_0.n1.t2 24.9236
R3653 carray_0.n1.n6 carray_0.n1.t4 18.6113
R3654 carray_0.n1 carray_0.n1.n0 15.0693
R3655 carray_0.n1.n4 carray_0.n1.n3 11.8308
R3656 carray_0.n1.n9 carray_0.n1.n8 9.3005
R3657 carray_0.n1.n7 carray_0.n1.n6 7.77627
R3658 carray_0.n1 carray_0.n1.n10 10.4321
R3659 carray_0.n1.n0 carray_0.n1.t0 7.07593
R3660 carray_0.n1.n0 carray_0.n1.t1 6.02718
R3661 carray_0.n1.n10 carray_0.n1.n9 1.93989
R3662 carray_0.n1.n9 carray_0.n1.n5 1.93989
R3663 carray_0.n1.n10 carray_0.n1.n1 1.35808
R3664 carray_0.n1.n5 carray_0.n1.n4 1.35808
R3665 carray_0.n1.n8 carray_0.n1.n7 0.9855
R3666 carray_0.n7.n135 carray_0.n7.n134 92.6295
R3667 carray_0.n7.n140 carray_0.n7.t0 25.6105
R3668 carray_0.n7.n134 carray_0.n7.t131 24.9236
R3669 carray_0.n7.n134 carray_0.n7.t130 24.9236
R3670 carray_0.n7.n138 carray_0.n7.t1 18.6113
R3671 carray_0.n7.n136 carray_0.n7.n135 11.8308
R3672 carray_0.n7.n141 carray_0.n7.n140 9.3005
R3673 carray_0.n7.n139 carray_0.n7.n138 7.77627
R3674 carray_0.n7.n15 carray_0.n7.n7 5.19252
R3675 carray_0.n7.n0 carray_0.n7.n142 4.57427
R3676 carray_0.n7.n74 carray_0.n7.n64 4.31395
R3677 carray_0.n7.n74 carray_0.n7.n73 3.66484
R3678 carray_0.n7.n15 carray_0.n7.n14 3.66465
R3679 carray_0.n7.n23 carray_0.n7.n22 3.66465
R3680 carray_0.n7.n31 carray_0.n7.n30 3.66465
R3681 carray_0.n7.n39 carray_0.n7.n38 3.66465
R3682 carray_0.n7.n47 carray_0.n7.n46 3.66465
R3683 carray_0.n7.n55 carray_0.n7.n54 3.66465
R3684 carray_0.n7.n82 carray_0.n7.n81 3.66465
R3685 carray_0.n7.n90 carray_0.n7.n89 3.66465
R3686 carray_0.n7.n98 carray_0.n7.n97 3.66465
R3687 carray_0.n7.n106 carray_0.n7.n105 3.66465
R3688 carray_0.n7.n114 carray_0.n7.n113 3.66465
R3689 carray_0.n7.n122 carray_0.n7.n121 3.66465
R3690 carray_0.n7.n130 carray_0.n7.n129 3.66465
R3691 carray_0.n7.n143 carray_0.n7.n0 3.0005
R3692 carray_0.n7 carray_0.n7.n144 2.8917
R3693 carray_0.n7.n63 carray_0.n7.n62 2.8155
R3694 carray_0.n7.n82 carray_0.n7.n74 2.29248
R3695 carray_0.n7.n64 carray_0.n7.n55 2.29232
R3696 carray_0.n7.n47 carray_0.n7.n39 2.29212
R3697 carray_0.n7.n98 carray_0.n7.n90 2.29212
R3698 carray_0.n7.n1 carray_0.n7.t76 2.15593
R3699 carray_0.n7.n8 carray_0.n7.t43 2.15593
R3700 carray_0.n7.n16 carray_0.n7.t2 2.15593
R3701 carray_0.n7.n24 carray_0.n7.t42 2.15593
R3702 carray_0.n7.n32 carray_0.n7.t3 2.15593
R3703 carray_0.n7.n40 carray_0.n7.t4 2.15593
R3704 carray_0.n7.n48 carray_0.n7.t22 2.15593
R3705 carray_0.n7.n56 carray_0.n7.t23 2.15593
R3706 carray_0.n7.n75 carray_0.n7.t116 2.15593
R3707 carray_0.n7.n83 carray_0.n7.t73 2.15593
R3708 carray_0.n7.n91 carray_0.n7.t100 2.15593
R3709 carray_0.n7.n99 carray_0.n7.t57 2.15593
R3710 carray_0.n7.n107 carray_0.n7.t102 2.15593
R3711 carray_0.n7.n115 carray_0.n7.t56 2.15593
R3712 carray_0.n7.n123 carray_0.n7.t101 2.15593
R3713 carray_0.n7.n65 carray_0.n7.t117 2.15593
R3714 carray_0.n7.n142 carray_0.n7.n141 1.93989
R3715 carray_0.n7.n141 carray_0.n7.n137 1.93989
R3716 carray_0.n7.n68 carray_0.n7.n67 1.63916
R3717 carray_0.n7.n31 carray_0.n7.n23 1.52837
R3718 carray_0.n7.n130 carray_0.n7.n122 1.52837
R3719 carray_0.n7.n114 carray_0.n7.n106 1.52837
R3720 carray_0.n7.n142 carray_0.n7.n133 1.35808
R3721 carray_0.n7.n137 carray_0.n7.n136 1.35808
R3722 carray_0.n7.n75 carray_0.n7.t123 1.16583
R3723 carray_0.n7.n76 carray_0.n7.t127 1.16583
R3724 carray_0.n7.n77 carray_0.n7.t128 1.16583
R3725 carray_0.n7.n78 carray_0.n7.t62 1.16583
R3726 carray_0.n7.n79 carray_0.n7.t66 1.16583
R3727 carray_0.n7.n80 carray_0.n7.t77 1.16583
R3728 carray_0.n7.n81 carray_0.n7.t79 1.16583
R3729 carray_0.n7.n83 carray_0.n7.t83 1.16583
R3730 carray_0.n7.n84 carray_0.n7.t88 1.16583
R3731 carray_0.n7.n85 carray_0.n7.t90 1.16583
R3732 carray_0.n7.n86 carray_0.n7.t27 1.16583
R3733 carray_0.n7.n87 carray_0.n7.t32 1.16583
R3734 carray_0.n7.n88 carray_0.n7.t38 1.16583
R3735 carray_0.n7.n89 carray_0.n7.t40 1.16583
R3736 carray_0.n7.n91 carray_0.n7.t105 1.16583
R3737 carray_0.n7.n92 carray_0.n7.t110 1.16583
R3738 carray_0.n7.n93 carray_0.n7.t115 1.16583
R3739 carray_0.n7.n94 carray_0.n7.t50 1.16583
R3740 carray_0.n7.n95 carray_0.n7.t53 1.16583
R3741 carray_0.n7.n96 carray_0.n7.t58 1.16583
R3742 carray_0.n7.n97 carray_0.n7.t61 1.16583
R3743 carray_0.n7.n99 carray_0.n7.t68 1.16583
R3744 carray_0.n7.n100 carray_0.n7.t70 1.16583
R3745 carray_0.n7.n101 carray_0.n7.t72 1.16583
R3746 carray_0.n7.n102 carray_0.n7.t17 1.16583
R3747 carray_0.n7.n103 carray_0.n7.t21 1.16583
R3748 carray_0.n7.n104 carray_0.n7.t24 1.16583
R3749 carray_0.n7.n105 carray_0.n7.t26 1.16583
R3750 carray_0.n7.n107 carray_0.n7.t106 1.16583
R3751 carray_0.n7.n108 carray_0.n7.t111 1.16583
R3752 carray_0.n7.n109 carray_0.n7.t119 1.16583
R3753 carray_0.n7.n110 carray_0.n7.t52 1.16583
R3754 carray_0.n7.n111 carray_0.n7.t55 1.16583
R3755 carray_0.n7.n112 carray_0.n7.t59 1.16583
R3756 carray_0.n7.n113 carray_0.n7.t64 1.16583
R3757 carray_0.n7.n115 carray_0.n7.t69 1.16583
R3758 carray_0.n7.n116 carray_0.n7.t71 1.16583
R3759 carray_0.n7.n117 carray_0.n7.t74 1.16583
R3760 carray_0.n7.n118 carray_0.n7.t19 1.16583
R3761 carray_0.n7.n119 carray_0.n7.t20 1.16583
R3762 carray_0.n7.n120 carray_0.n7.t25 1.16583
R3763 carray_0.n7.n121 carray_0.n7.t28 1.16583
R3764 carray_0.n7.n123 carray_0.n7.t107 1.16583
R3765 carray_0.n7.n124 carray_0.n7.t112 1.16583
R3766 carray_0.n7.n125 carray_0.n7.t118 1.16583
R3767 carray_0.n7.n126 carray_0.n7.t51 1.16583
R3768 carray_0.n7.n127 carray_0.n7.t54 1.16583
R3769 carray_0.n7.n128 carray_0.n7.t60 1.16583
R3770 carray_0.n7.n129 carray_0.n7.t65 1.16583
R3771 carray_0.n7.n7 carray_0.n7.t41 1.10593
R3772 carray_0.n7.n6 carray_0.n7.t39 1.10593
R3773 carray_0.n7.n5 carray_0.n7.t33 1.10593
R3774 carray_0.n7.n4 carray_0.n7.t29 1.10593
R3775 carray_0.n7.n3 carray_0.n7.t91 1.10593
R3776 carray_0.n7.n2 carray_0.n7.t89 1.10593
R3777 carray_0.n7.n1 carray_0.n7.t84 1.10593
R3778 carray_0.n7.n14 carray_0.n7.t7 1.10593
R3779 carray_0.n7.n13 carray_0.n7.t5 1.10593
R3780 carray_0.n7.n12 carray_0.n7.t124 1.10593
R3781 carray_0.n7.n11 carray_0.n7.t121 1.10593
R3782 carray_0.n7.n10 carray_0.n7.t49 1.10593
R3783 carray_0.n7.n9 carray_0.n7.t46 1.10593
R3784 carray_0.n7.n8 carray_0.n7.t44 1.10593
R3785 carray_0.n7.n22 carray_0.n7.t95 1.10593
R3786 carray_0.n7.n21 carray_0.n7.t92 1.10593
R3787 carray_0.n7.n20 carray_0.n7.t85 1.10593
R3788 carray_0.n7.n19 carray_0.n7.t80 1.10593
R3789 carray_0.n7.n18 carray_0.n7.t16 1.10593
R3790 carray_0.n7.n17 carray_0.n7.t13 1.10593
R3791 carray_0.n7.n16 carray_0.n7.t10 1.10593
R3792 carray_0.n7.n30 carray_0.n7.t8 1.10593
R3793 carray_0.n7.n29 carray_0.n7.t6 1.10593
R3794 carray_0.n7.n28 carray_0.n7.t125 1.10593
R3795 carray_0.n7.n27 carray_0.n7.t120 1.10593
R3796 carray_0.n7.n26 carray_0.n7.t48 1.10593
R3797 carray_0.n7.n25 carray_0.n7.t47 1.10593
R3798 carray_0.n7.n24 carray_0.n7.t45 1.10593
R3799 carray_0.n7.n38 carray_0.n7.t96 1.10593
R3800 carray_0.n7.n37 carray_0.n7.t93 1.10593
R3801 carray_0.n7.n36 carray_0.n7.t86 1.10593
R3802 carray_0.n7.n35 carray_0.n7.t81 1.10593
R3803 carray_0.n7.n34 carray_0.n7.t15 1.10593
R3804 carray_0.n7.n33 carray_0.n7.t12 1.10593
R3805 carray_0.n7.n32 carray_0.n7.t9 1.10593
R3806 carray_0.n7.n46 carray_0.n7.t97 1.10593
R3807 carray_0.n7.n45 carray_0.n7.t94 1.10593
R3808 carray_0.n7.n44 carray_0.n7.t87 1.10593
R3809 carray_0.n7.n43 carray_0.n7.t82 1.10593
R3810 carray_0.n7.n42 carray_0.n7.t18 1.10593
R3811 carray_0.n7.n41 carray_0.n7.t14 1.10593
R3812 carray_0.n7.n40 carray_0.n7.t11 1.10593
R3813 carray_0.n7.n54 carray_0.n7.t113 1.10593
R3814 carray_0.n7.n53 carray_0.n7.t108 1.10593
R3815 carray_0.n7.n52 carray_0.n7.t103 1.10593
R3816 carray_0.n7.n51 carray_0.n7.t99 1.10593
R3817 carray_0.n7.n50 carray_0.n7.t37 1.10593
R3818 carray_0.n7.n49 carray_0.n7.t35 1.10593
R3819 carray_0.n7.n48 carray_0.n7.t30 1.10593
R3820 carray_0.n7.n62 carray_0.n7.t114 1.10593
R3821 carray_0.n7.n61 carray_0.n7.t109 1.10593
R3822 carray_0.n7.n60 carray_0.n7.t104 1.10593
R3823 carray_0.n7.n59 carray_0.n7.t98 1.10593
R3824 carray_0.n7.n58 carray_0.n7.t36 1.10593
R3825 carray_0.n7.n57 carray_0.n7.t34 1.10593
R3826 carray_0.n7.n56 carray_0.n7.t31 1.10593
R3827 carray_0.n7.n65 carray_0.n7.t122 1.10593
R3828 carray_0.n7.n66 carray_0.n7.t126 1.10593
R3829 carray_0.n7.n70 carray_0.n7.t63 1.10593
R3830 carray_0.n7.n71 carray_0.n7.t67 1.10593
R3831 carray_0.n7.n72 carray_0.n7.t75 1.10593
R3832 carray_0.n7.n73 carray_0.n7.t78 1.10593
R3833 carray_0.n7.n69 carray_0.n7.n68 1.08606
R3834 carray_0.n7.n2 carray_0.n7.n1 1.0505
R3835 carray_0.n7.n3 carray_0.n7.n2 1.0505
R3836 carray_0.n7.n4 carray_0.n7.n3 1.0505
R3837 carray_0.n7.n5 carray_0.n7.n4 1.0505
R3838 carray_0.n7.n6 carray_0.n7.n5 1.0505
R3839 carray_0.n7.n7 carray_0.n7.n6 1.0505
R3840 carray_0.n7.n9 carray_0.n7.n8 1.0505
R3841 carray_0.n7.n10 carray_0.n7.n9 1.0505
R3842 carray_0.n7.n11 carray_0.n7.n10 1.0505
R3843 carray_0.n7.n12 carray_0.n7.n11 1.0505
R3844 carray_0.n7.n13 carray_0.n7.n12 1.0505
R3845 carray_0.n7.n14 carray_0.n7.n13 1.0505
R3846 carray_0.n7.n17 carray_0.n7.n16 1.0505
R3847 carray_0.n7.n18 carray_0.n7.n17 1.0505
R3848 carray_0.n7.n19 carray_0.n7.n18 1.0505
R3849 carray_0.n7.n20 carray_0.n7.n19 1.0505
R3850 carray_0.n7.n21 carray_0.n7.n20 1.0505
R3851 carray_0.n7.n22 carray_0.n7.n21 1.0505
R3852 carray_0.n7.n25 carray_0.n7.n24 1.0505
R3853 carray_0.n7.n26 carray_0.n7.n25 1.0505
R3854 carray_0.n7.n27 carray_0.n7.n26 1.0505
R3855 carray_0.n7.n28 carray_0.n7.n27 1.0505
R3856 carray_0.n7.n29 carray_0.n7.n28 1.0505
R3857 carray_0.n7.n30 carray_0.n7.n29 1.0505
R3858 carray_0.n7.n33 carray_0.n7.n32 1.0505
R3859 carray_0.n7.n34 carray_0.n7.n33 1.0505
R3860 carray_0.n7.n35 carray_0.n7.n34 1.0505
R3861 carray_0.n7.n36 carray_0.n7.n35 1.0505
R3862 carray_0.n7.n37 carray_0.n7.n36 1.0505
R3863 carray_0.n7.n38 carray_0.n7.n37 1.0505
R3864 carray_0.n7.n41 carray_0.n7.n40 1.0505
R3865 carray_0.n7.n42 carray_0.n7.n41 1.0505
R3866 carray_0.n7.n43 carray_0.n7.n42 1.0505
R3867 carray_0.n7.n44 carray_0.n7.n43 1.0505
R3868 carray_0.n7.n45 carray_0.n7.n44 1.0505
R3869 carray_0.n7.n46 carray_0.n7.n45 1.0505
R3870 carray_0.n7.n49 carray_0.n7.n48 1.0505
R3871 carray_0.n7.n50 carray_0.n7.n49 1.0505
R3872 carray_0.n7.n51 carray_0.n7.n50 1.0505
R3873 carray_0.n7.n52 carray_0.n7.n51 1.0505
R3874 carray_0.n7.n53 carray_0.n7.n52 1.0505
R3875 carray_0.n7.n54 carray_0.n7.n53 1.0505
R3876 carray_0.n7.n57 carray_0.n7.n56 1.0505
R3877 carray_0.n7.n58 carray_0.n7.n57 1.0505
R3878 carray_0.n7.n59 carray_0.n7.n58 1.0505
R3879 carray_0.n7.n60 carray_0.n7.n59 1.0505
R3880 carray_0.n7.n61 carray_0.n7.n60 1.0505
R3881 carray_0.n7.n62 carray_0.n7.n61 1.0505
R3882 carray_0.n7.n76 carray_0.n7.n75 1.0505
R3883 carray_0.n7.n77 carray_0.n7.n76 1.0505
R3884 carray_0.n7.n78 carray_0.n7.n77 1.0505
R3885 carray_0.n7.n79 carray_0.n7.n78 1.0505
R3886 carray_0.n7.n80 carray_0.n7.n79 1.0505
R3887 carray_0.n7.n81 carray_0.n7.n80 1.0505
R3888 carray_0.n7.n84 carray_0.n7.n83 1.0505
R3889 carray_0.n7.n85 carray_0.n7.n84 1.0505
R3890 carray_0.n7.n86 carray_0.n7.n85 1.0505
R3891 carray_0.n7.n87 carray_0.n7.n86 1.0505
R3892 carray_0.n7.n88 carray_0.n7.n87 1.0505
R3893 carray_0.n7.n89 carray_0.n7.n88 1.0505
R3894 carray_0.n7.n92 carray_0.n7.n91 1.0505
R3895 carray_0.n7.n93 carray_0.n7.n92 1.0505
R3896 carray_0.n7.n94 carray_0.n7.n93 1.0505
R3897 carray_0.n7.n95 carray_0.n7.n94 1.0505
R3898 carray_0.n7.n96 carray_0.n7.n95 1.0505
R3899 carray_0.n7.n97 carray_0.n7.n96 1.0505
R3900 carray_0.n7.n100 carray_0.n7.n99 1.0505
R3901 carray_0.n7.n101 carray_0.n7.n100 1.0505
R3902 carray_0.n7.n102 carray_0.n7.n101 1.0505
R3903 carray_0.n7.n103 carray_0.n7.n102 1.0505
R3904 carray_0.n7.n104 carray_0.n7.n103 1.0505
R3905 carray_0.n7.n105 carray_0.n7.n104 1.0505
R3906 carray_0.n7.n108 carray_0.n7.n107 1.0505
R3907 carray_0.n7.n109 carray_0.n7.n108 1.0505
R3908 carray_0.n7.n110 carray_0.n7.n109 1.0505
R3909 carray_0.n7.n111 carray_0.n7.n110 1.0505
R3910 carray_0.n7.n112 carray_0.n7.n111 1.0505
R3911 carray_0.n7.n113 carray_0.n7.n112 1.0505
R3912 carray_0.n7.n116 carray_0.n7.n115 1.0505
R3913 carray_0.n7.n117 carray_0.n7.n116 1.0505
R3914 carray_0.n7.n118 carray_0.n7.n117 1.0505
R3915 carray_0.n7.n119 carray_0.n7.n118 1.0505
R3916 carray_0.n7.n120 carray_0.n7.n119 1.0505
R3917 carray_0.n7.n121 carray_0.n7.n120 1.0505
R3918 carray_0.n7.n124 carray_0.n7.n123 1.0505
R3919 carray_0.n7.n125 carray_0.n7.n124 1.0505
R3920 carray_0.n7.n126 carray_0.n7.n125 1.0505
R3921 carray_0.n7.n127 carray_0.n7.n126 1.0505
R3922 carray_0.n7.n128 carray_0.n7.n127 1.0505
R3923 carray_0.n7.n129 carray_0.n7.n128 1.0505
R3924 carray_0.n7.n66 carray_0.n7.n65 1.0505
R3925 carray_0.n7.n69 carray_0.n7.n66 1.0505
R3926 carray_0.n7.n70 carray_0.n7.n69 1.0505
R3927 carray_0.n7.n71 carray_0.n7.n70 1.0505
R3928 carray_0.n7.n72 carray_0.n7.n71 1.0505
R3929 carray_0.n7.n73 carray_0.n7.n72 1.0505
R3930 carray_0.n7.n140 carray_0.n7.n139 0.9855
R3931 carray_0.n7.n64 carray_0.n7.n63 0.84191
R3932 carray_0.n7.n23 carray_0.n7.n15 0.764617
R3933 carray_0.n7.n39 carray_0.n7.n31 0.764617
R3934 carray_0.n7.n55 carray_0.n7.n47 0.764617
R3935 carray_0.n7.n122 carray_0.n7.n114 0.764617
R3936 carray_0.n7.n106 carray_0.n7.n98 0.764617
R3937 carray_0.n7.n90 carray_0.n7.n82 0.764617
R3938 carray_0.n7 carray_0.n7.n130 0.752473
R3939 carray_0.n7.n63 carray_0.n7 0.08175
R3940 carray_0.n7.n63 carray_0.n7 0.04925
R3941 carray_0.n7.n144 carray_0.n7.n143 0.0333125
R3942 carray_0.n7.n68 carray_0.n7.t129 0.02118
R3943 carray_0.n7.n0 carray_0.n7.n132 0.0126789
R3944 carray_0.n7.n0 carray_0.n7.n131 0.0122188
R3945 a_44621_6352.n11 a_44621_6352.t21 212.081
R3946 a_44621_6352.n9 a_44621_6352.t20 212.081
R3947 a_44621_6352.n5 a_44621_6352.t19 212.081
R3948 a_44621_6352.n3 a_44621_6352.t18 212.081
R3949 a_44621_6352.n26 a_44621_6352.n25 146.423
R3950 a_44621_6352.n2 a_44621_6352.n0 144.089
R3951 a_44621_6352.n13 a_44621_6352.t14 143.071
R3952 a_44621_6352.n21 a_44621_6352.t8 142.75
R3953 a_44621_6352.n13 a_44621_6352.t23 142.75
R3954 a_44621_6352.n14 a_44621_6352.t10 142.75
R3955 a_44621_6352.n15 a_44621_6352.t9 142.75
R3956 a_44621_6352.n16 a_44621_6352.t17 142.75
R3957 a_44621_6352.n17 a_44621_6352.t25 142.75
R3958 a_44621_6352.n18 a_44621_6352.t12 142.75
R3959 a_44621_6352.n19 a_44621_6352.t22 142.75
R3960 a_44621_6352.n20 a_44621_6352.t24 142.75
R3961 a_44621_6352.n11 a_44621_6352.t16 139.78
R3962 a_44621_6352.n9 a_44621_6352.t15 139.78
R3963 a_44621_6352.n5 a_44621_6352.t13 139.78
R3964 a_44621_6352.n3 a_44621_6352.t11 139.78
R3965 a_44621_6352.n2 a_44621_6352.n1 107.822
R3966 a_44621_6352.n25 a_44621_6352.n24 107.249
R3967 a_44621_6352.n7 a_44621_6352.n4 97.5045
R3968 a_44621_6352.n7 a_44621_6352.n6 76.0005
R3969 a_44621_6352.n23 a_44621_6352.n2 46.6252
R3970 a_44621_6352.n12 a_44621_6352.n11 39.8685
R3971 a_44621_6352.n4 a_44621_6352.n3 30.6732
R3972 a_44621_6352.n6 a_44621_6352.n5 30.6732
R3973 a_44621_6352.n10 a_44621_6352.n9 30.6732
R3974 a_44621_6352.n11 a_44621_6352.n10 30.6732
R3975 a_44621_6352.n24 a_44621_6352.t5 26.5955
R3976 a_44621_6352.n24 a_44621_6352.t6 26.5955
R3977 a_44621_6352.n26 a_44621_6352.t4 26.5955
R3978 a_44621_6352.t7 a_44621_6352.n26 26.5955
R3979 a_44621_6352.n0 a_44621_6352.t1 24.9236
R3980 a_44621_6352.n0 a_44621_6352.t0 24.9236
R3981 a_44621_6352.n1 a_44621_6352.t2 24.9236
R3982 a_44621_6352.n1 a_44621_6352.t3 24.9236
R3983 a_44621_6352.n8 a_44621_6352.n7 21.5045
R3984 a_44621_6352.n12 a_44621_6352.n8 19.201
R3985 a_44621_6352.n25 a_44621_6352.n23 14.3512
R3986 a_44621_6352.n22 a_44621_6352.n21 9.01046
R3987 a_44621_6352.n23 a_44621_6352.n22 4.58256
R3988 a_44621_6352.n22 a_44621_6352.n12 1.91581
R3989 a_44621_6352.n21 a_44621_6352.n20 0.321152
R3990 a_44621_6352.n20 a_44621_6352.n19 0.321152
R3991 a_44621_6352.n19 a_44621_6352.n18 0.321152
R3992 a_44621_6352.n18 a_44621_6352.n17 0.321152
R3993 a_44621_6352.n17 a_44621_6352.n16 0.321152
R3994 a_44621_6352.n16 a_44621_6352.n15 0.321152
R3995 a_44621_6352.n15 a_44621_6352.n14 0.321152
R3996 a_44621_6352.n14 a_44621_6352.n13 0.321152
R3997 ctl4.n0 ctl4.t2 212.081
R3998 ctl4.n1 ctl4.t0 212.081
R3999 ctl4.n0 ctl4.t3 139.78
R4000 ctl4.n1 ctl4.t1 139.78
R4001 ctl4.n1 ctl4.n0 61.346
R4002 ctl4 ctl4.n1 44.6884
R4003 carray_0.n4.n17 carray_0.n4.n16 92.6295
R4004 carray_0.n4.n22 carray_0.n4.t3 25.6105
R4005 carray_0.n4.n16 carray_0.n4.t1 24.9236
R4006 carray_0.n4.n16 carray_0.n4.t0 24.9236
R4007 carray_0.n4.n20 carray_0.n4.t2 18.6113
R4008 carray_0.n4.n18 carray_0.n4.n17 11.8308
R4009 carray_0.n4 carray_0.n4.n14 11.445
R4010 carray_0.n4.n23 carray_0.n4.n22 9.3005
R4011 carray_0.n4.n21 carray_0.n4.n20 7.77627
R4012 carray_0.n4 carray_0.n4.n24 10.7047
R4013 carray_0.n4.n14 carray_0.n4.n6 5.85019
R4014 carray_0.n4.n14 carray_0.n4.n13 3.06465
R4015 carray_0.n4.n0 carray_0.n4.t12 2.15593
R4016 carray_0.n4.n7 carray_0.n4.t16 2.15593
R4017 carray_0.n4.n24 carray_0.n4.n23 1.93989
R4018 carray_0.n4.n23 carray_0.n4.n19 1.93989
R4019 carray_0.n4.n24 carray_0.n4.n15 1.35808
R4020 carray_0.n4.n19 carray_0.n4.n18 1.35808
R4021 carray_0.n4.n6 carray_0.n4.t7 1.10593
R4022 carray_0.n4.n5 carray_0.n4.t6 1.10593
R4023 carray_0.n4.n4 carray_0.n4.t5 1.10593
R4024 carray_0.n4.n3 carray_0.n4.t4 1.10593
R4025 carray_0.n4.n2 carray_0.n4.t15 1.10593
R4026 carray_0.n4.n1 carray_0.n4.t14 1.10593
R4027 carray_0.n4.n0 carray_0.n4.t13 1.10593
R4028 carray_0.n4.n7 carray_0.n4.t17 1.10593
R4029 carray_0.n4.n8 carray_0.n4.t18 1.10593
R4030 carray_0.n4.n9 carray_0.n4.t19 1.10593
R4031 carray_0.n4.n10 carray_0.n4.t8 1.10593
R4032 carray_0.n4.n11 carray_0.n4.t9 1.10593
R4033 carray_0.n4.n12 carray_0.n4.t10 1.10593
R4034 carray_0.n4.n13 carray_0.n4.t11 1.10593
R4035 carray_0.n4.n1 carray_0.n4.n0 1.0505
R4036 carray_0.n4.n2 carray_0.n4.n1 1.0505
R4037 carray_0.n4.n3 carray_0.n4.n2 1.0505
R4038 carray_0.n4.n4 carray_0.n4.n3 1.0505
R4039 carray_0.n4.n5 carray_0.n4.n4 1.0505
R4040 carray_0.n4.n6 carray_0.n4.n5 1.0505
R4041 carray_0.n4.n8 carray_0.n4.n7 1.0505
R4042 carray_0.n4.n9 carray_0.n4.n8 1.0505
R4043 carray_0.n4.n10 carray_0.n4.n9 1.0505
R4044 carray_0.n4.n11 carray_0.n4.n10 1.0505
R4045 carray_0.n4.n12 carray_0.n4.n11 1.0505
R4046 carray_0.n4.n13 carray_0.n4.n12 1.0505
R4047 carray_0.n4.n22 carray_0.n4.n21 0.9855
R4048 en_buf.n5 en_buf.n3 146.424
R4049 en_buf.n2 en_buf.n0 144.089
R4050 en_buf.n7 en_buf.t17 135.841
R4051 en_buf.n11 en_buf.t20 135.841
R4052 en_buf.n9 en_buf.t18 135.52
R4053 en_buf.n8 en_buf.t21 135.52
R4054 en_buf.n7 en_buf.t24 135.52
R4055 en_buf.n11 en_buf.t23 135.52
R4056 en_buf.n12 en_buf.t25 135.52
R4057 en_buf.n13 en_buf.t19 135.52
R4058 en_buf.n14 en_buf.t22 134.576
R4059 en_buf.n10 en_buf.t16 134.576
R4060 en_buf.n2 en_buf.n1 107.822
R4061 en_buf.n5 en_buf.n4 107.249
R4062 en_buf.n6 en_buf.n2 46.6252
R4063 en_buf.n4 en_buf.t9 26.5955
R4064 en_buf.n4 en_buf.t15 26.5955
R4065 en_buf.n3 en_buf.t14 26.5955
R4066 en_buf.n3 en_buf.t11 26.5955
R4067 en_buf.n0 en_buf.t0 24.9236
R4068 en_buf.n0 en_buf.t5 24.9236
R4069 en_buf.n1 en_buf.t3 24.9236
R4070 en_buf.n1 en_buf.t1 24.9236
R4071 en_buf.n6 en_buf.n5 14.3512
R4072 en_buf en_buf.n6 8.71285
R4073 en_buf en_buf.n15 1.05289
R4074 en_buf.n8 en_buf.n7 0.321152
R4075 en_buf.n9 en_buf.n8 0.321152
R4076 en_buf.n13 en_buf.n12 0.321152
R4077 en_buf.n12 en_buf.n11 0.321152
R4078 en_buf.n10 en_buf.n9 0.315896
R4079 en_buf.n14 en_buf.n13 0.315896
R4080 en_buf.n15 en_buf.n10 0.121984
R4081 en_buf.n15 en_buf.n14 0.121984
R4082 ctl2.n0 ctl2.t1 212.081
R4083 ctl2.n1 ctl2.t3 212.081
R4084 ctl2.n0 ctl2.t2 139.78
R4085 ctl2.n1 ctl2.t0 139.78
R4086 ctl2.n1 ctl2.n0 61.346
R4087 ctl2 ctl2.n1 44.6884
R4088 carray_0.n2.n5 carray_0.n2.n4 92.6295
R4089 carray_0.n2.n10 carray_0.n2.t6 25.6105
R4090 carray_0.n2.n4 carray_0.n2.t5 24.9236
R4091 carray_0.n2.n4 carray_0.n2.t4 24.9236
R4092 carray_0.n2.n8 carray_0.n2.t7 18.6113
R4093 carray_0.n2 carray_0.n2.n2 12.103
R4094 carray_0.n2.n6 carray_0.n2.n5 11.8308
R4095 carray_0.n2.n11 carray_0.n2.n10 9.3005
R4096 carray_0.n2.n9 carray_0.n2.n8 7.77627
R4097 carray_0.n2 carray_0.n2.n12 10.841
R4098 carray_0.n2.n0 carray_0.n2.t2 4.59115
R4099 carray_0.n2.n1 carray_0.n2.t1 4.591
R4100 carray_0.n2.n0 carray_0.n2.t0 3.41984
R4101 carray_0.n2.n1 carray_0.n2.t3 3.4197
R4102 carray_0.n2.n2 carray_0.n2.n0 2.81726
R4103 carray_0.n2.n12 carray_0.n2.n11 1.93989
R4104 carray_0.n2.n11 carray_0.n2.n7 1.93989
R4105 carray_0.n2.n2 carray_0.n2.n1 1.46601
R4106 carray_0.n2.n12 carray_0.n2.n3 1.35808
R4107 carray_0.n2.n7 carray_0.n2.n6 1.35808
R4108 carray_0.n2.n10 carray_0.n2.n9 0.9855
R4109 ctl5.n0 ctl5.t3 212.081
R4110 ctl5.n1 ctl5.t2 212.081
R4111 ctl5.n0 ctl5.t1 139.78
R4112 ctl5.n1 ctl5.t0 139.78
R4113 ctl5.n1 ctl5.n0 61.346
R4114 ctl5 ctl5.n1 44.6884
R4115 carray_0.n3.n9 carray_0.n3.n8 92.6295
R4116 carray_0.n3.n14 carray_0.n3.t9 25.6105
R4117 carray_0.n3.n8 carray_0.n3.t10 24.9236
R4118 carray_0.n3.n8 carray_0.n3.t0 24.9236
R4119 carray_0.n3.n12 carray_0.n3.t11 18.6113
R4120 carray_0.n3 carray_0.n3.n6 12.2087
R4121 carray_0.n3.n10 carray_0.n3.n9 11.8308
R4122 carray_0.n3.n15 carray_0.n3.n14 9.3005
R4123 carray_0.n3.n13 carray_0.n3.n12 7.77627
R4124 carray_0.n3.n1 carray_0.n3.n0 5.2505
R4125 carray_0.n3.n4 carray_0.n3.n3 5.2505
R4126 carray_0.n3 carray_0.n3.n16 10.7728
R4127 carray_0.n3.n6 carray_0.n3.n2 4.12269
R4128 carray_0.n3.n6 carray_0.n3.n5 2.86465
R4129 carray_0.n3.n0 carray_0.n3.t5 2.15593
R4130 carray_0.n3.n3 carray_0.n3.t1 2.15593
R4131 carray_0.n3.n16 carray_0.n3.n15 1.93989
R4132 carray_0.n3.n15 carray_0.n3.n11 1.93989
R4133 carray_0.n3.n16 carray_0.n3.n7 1.35808
R4134 carray_0.n3.n11 carray_0.n3.n10 1.35808
R4135 carray_0.n3.n2 carray_0.n3.t3 1.10593
R4136 carray_0.n3.n1 carray_0.n3.t2 1.10593
R4137 carray_0.n3.n0 carray_0.n3.t6 1.10593
R4138 carray_0.n3.n3 carray_0.n3.t4 1.10593
R4139 carray_0.n3.n4 carray_0.n3.t7 1.10593
R4140 carray_0.n3.n5 carray_0.n3.t8 1.10593
R4141 carray_0.n3.n2 carray_0.n3.n1 1.0505
R4142 carray_0.n3.n5 carray_0.n3.n4 1.0505
R4143 carray_0.n3.n14 carray_0.n3.n13 0.9855
R4144 dum.n0 dum.t3 212.081
R4145 dum.n1 dum.t2 212.081
R4146 dum.n0 dum.t1 139.78
R4147 dum.n1 dum.t0 139.78
R4148 dum.n1 dum.n0 61.346
R4149 dum dum.n1 44.6494
R4150 carray_0.ndum.n2 carray_0.ndum.n1 92.6295
R4151 carray_0.ndum.n7 carray_0.ndum.t3 25.6105
R4152 carray_0.ndum.n1 carray_0.ndum.t1 24.9236
R4153 carray_0.ndum.n1 carray_0.ndum.t0 24.9236
R4154 carray_0.ndum carray_0.ndum.t4 22.0057
R4155 carray_0.ndum.n5 carray_0.ndum.t2 18.6113
R4156 carray_0.ndum.n3 carray_0.ndum.n2 11.8308
R4157 carray_0.ndum.n8 carray_0.ndum.n7 9.3005
R4158 carray_0.ndum.n6 carray_0.ndum.n5 7.77627
R4159 carray_0.ndum carray_0.ndum.n9 10.2958
R4160 carray_0.ndum.n9 carray_0.ndum.n8 1.93989
R4161 carray_0.ndum.n8 carray_0.ndum.n4 1.93989
R4162 carray_0.ndum.n9 carray_0.ndum.n0 1.35808
R4163 carray_0.ndum.n4 carray_0.ndum.n3 1.35808
R4164 carray_0.ndum.n7 carray_0.ndum.n6 0.9855
R4165 ctl0.n0 ctl0.t1 212.081
R4166 ctl0.n1 ctl0.t3 212.081
R4167 ctl0.n0 ctl0.t2 139.78
R4168 ctl0.n1 ctl0.t0 139.78
R4169 ctl0.n1 ctl0.n0 61.346
R4170 ctl0 ctl0.n1 44.6884
R4171 carray_0.n0.n2 carray_0.n0.n1 92.6295
R4172 carray_0.n0.n7 carray_0.n0.t3 25.6105
R4173 carray_0.n0.n1 carray_0.n0.t2 24.9236
R4174 carray_0.n0.n1 carray_0.n0.t1 24.9236
R4175 carray_0.n0 carray_0.n0.t0 21.6121
R4176 carray_0.n0.n5 carray_0.n0.t4 18.6113
R4177 carray_0.n0.n3 carray_0.n0.n2 11.8308
R4178 carray_0.n0.n8 carray_0.n0.n7 9.3005
R4179 carray_0.n0.n6 carray_0.n0.n5 7.77627
R4180 carray_0.n0 carray_0.n0.n9 10.3639
R4181 carray_0.n0.n9 carray_0.n0.n8 1.93989
R4182 carray_0.n0.n8 carray_0.n0.n4 1.93989
R4183 carray_0.n0.n9 carray_0.n0.n0 1.35808
R4184 carray_0.n0.n4 carray_0.n0.n3 1.35808
R4185 carray_0.n0.n7 carray_0.n0.n6 0.9855
R4186 ctl7.n0 ctl7.t1 212.081
R4187 ctl7.n1 ctl7.t0 212.081
R4188 ctl7.n0 ctl7.t3 139.78
R4189 ctl7.n1 ctl7.t2 139.78
R4190 ctl7.n1 ctl7.n0 61.346
R4191 ctl7 ctl7.n1 44.6884
R4192 ctl3.n0 ctl3.t2 212.081
R4193 ctl3.n1 ctl3.t0 212.081
R4194 ctl3.n0 ctl3.t3 139.78
R4195 ctl3.n1 ctl3.t1 139.78
R4196 ctl3.n1 ctl3.n0 61.346
R4197 ctl3 ctl3.n1 44.6884
R4198 ctl6.n0 ctl6.t1 212.081
R4199 ctl6.n1 ctl6.t0 212.081
R4200 ctl6.n0 ctl6.t3 139.78
R4201 ctl6.n1 ctl6.t2 139.78
R4202 ctl6.n1 ctl6.n0 61.346
R4203 ctl6 ctl6.n1 44.6884
C0 m2_4325_1830# m2_5029_1610# 0.251f
C1 carray_0.n6 out 48.6f
C2 m3_40429_1610# out 0.187f
C3 carray_0.ndum carray_0.n3 1.36f
C4 carray_0.ndum m2_16729_1610# 3.15e-20
C5 m2_12125_9390# m2_12829_1610# 0.251f
C6 m2_425_5190# out 0.719f
C7 m3_35029_1610# out 0.187f
C8 carray_0.n6 m3_38929_1610# 0.00746f
C9 m3_40229_1610# m3_39129_1610# 0.148f
C10 carray_0.n6 m3_32429_1610# 4.08f
C11 ctl7 sample 0.00169f
C12 carray_0.n7 m2_9525_1830# 0.452f
C13 carray_0.n7 m2_3729_1610# 1.13f
C14 carray_0.n6 m2_26425_9390# 0.452f
C15 out vin 21.5f
C16 carray_0.n7 m3_19429_1610# 1.98f
C17 m2_37929_1610# m2_38125_9390# 0.251f
C18 carray_0.n7 m2_22525_1830# 9.11e-20
C19 carray_0.n0 m2_11529_1610# 6.36e-20
C20 m2_37929_1610# out 0.267f
C21 enb vdd 4.26f
C22 m3_4029_1610# m2_4325_1830# 0.247f
C23 m3_5129_1610# m2_4325_9390# 0.247f
C24 m3_35229_1610# m2_35329_1610# 2.11f
C25 carray_0.n5 m2_23825_1830# 2.03e-19
C26 m2_37929_1610# m3_38929_1610# 0.0061f
C27 carray_0.n6 m2_31429_1610# 2.39f
C28 m2_38125_9390# m3_37829_1610# 0.247f
C29 m2_43325_4350# vin 0.0402f
C30 m3_37829_1610# out 0.187f
C31 ctl0 carray_0.n1 0.0175f
C32 ctl1 carray_0.n0 0.00139f
C33 m3_37829_1610# m3_38929_1610# 0.148f
C34 m2_35329_1610# out 0.267f
C35 m2_26229_1610# out 0.267f
C36 carray_0.n2 m2_425_1830# 0.332f
C37 m2_425_9390# out 0.779f
C38 m2_12829_1610# m3_12929_1610# 2.11f
C39 m2_10229_1610# m3_10529_1610# 0.181f
C40 m2_24929_1610# sample 6.55e-20
C41 m2_34029_1610# m3_33929_1610# 2.11f
C42 m2_30325_1830# out 0.643f
C43 m3_3829_1610# m3_4029_1610# 3.35f
C44 carray_0.n7 m2_8225_9390# 0.452f
C45 carray_0.n2 m2_4325_1830# 0.169f
C46 m2_26229_1610# m2_26425_9390# 0.251f
C47 carray_0.n2 m3_20729_1610# 3.43f
C48 m2_425_9390# m2_425_8550# 0.199f
C49 carray_0.n5 m3_24829_1610# 0.00889f
C50 m3_30029_1610# m3_31129_1610# 0.148f
C51 carray_0.n1 m2_8929_1610# 8.05e-20
C52 m2_425_4350# m2_1129_1610# 0.251f
C53 carray_0.n5 m2_29025_1830# 0.0714f
C54 ctl0 dum 0.193f
C55 m3_29829_1610# m2_28829_1610# 0.0061f
C56 carray_0.n1 m2_22525_9390# 0.251f
C57 m3_28529_1610# m2_28829_1610# 0.181f
C58 m2_15429_1610# m3_15529_1610# 2.11f
C59 carray_0.n6 m2_23629_1610# 1.43e-19
C60 m3_3829_1610# m2_3025_9390# 0.247f
C61 m2_1129_1610# out 0.267f
C62 m2_32925_1830# m3_32629_1610# 0.247f
C63 m2_32925_9390# m3_33729_1610# 0.247f
C64 carray_0.n2 m3_3829_1610# 0.021f
C65 sample m2_30129_1610# 6.55e-20
C66 m2_14129_1610# m3_13129_1610# 0.0061f
C67 carray_0.n7 m3_40229_1610# 4.08f
C68 carray_0.n0 carray_0.n4 0.0773f
C69 m2_425_8550# m2_1129_1610# 0.251f
C70 m3_23529_1610# out 0.187f
C71 m2_5029_1610# out 0.267f
C72 carray_0.n4 m2_17325_1830# 2.85e-19
C73 carray_0.n3 m2_9525_1830# 4.28e-19
C74 m3_9229_1610# m3_10329_1610# 0.148f
C75 carray_0.n1 m2_6925_1830# 9.38e-20
C76 carray_0.n6 m3_31329_1610# 1.98f
C77 carray_0.n2 m3_9229_1610# 0.021f
C78 carray_0.n3 m2_3729_1610# 5.59e-19
C79 carray_0.n2 m2_2429_1610# 0.00855f
C80 carray_0.n3 m2_22525_1830# 0.453f
C81 ctl5 vdd 0.158f
C82 vin m2_43129_1610# 0.00125f
C83 carray_0.n1 sample 0.00244f
C84 carray_0.n6 m2_28829_1610# 1.43e-19
C85 carray_0.n7 m2_36825_1830# 1.18e-19
C86 m2_12125_9390# m3_12929_1610# 0.247f
C87 out m2_42025_1830# 0.643f
C88 m2_40725_1830# carray_0.n6 0.512f
C89 m2_40725_9390# m3_41529_1610# 0.247f
C90 m2_40725_1830# m3_40429_1610# 0.247f
C91 m3_4029_1610# out 0.187f
C92 carray_0.n4 m2_14725_1830# 2.85e-19
C93 m2_20629_1610# carray_0.n2 0.256f
C94 m3_31129_1610# out 0.187f
C95 carray_0.n6 m2_3025_1830# 0.452f
C96 carray_0.n7 m2_34225_1830# 0.452f
C97 m2_18625_9390# m3_18329_1610# 0.247f
C98 m2_35525_1830# sample 9.23e-21
C99 carray_0.n7 m2_25125_1830# 0.452f
C100 carray_0.n1 carray_0.ndum 3.54f
C101 m2_40725_9390# out 0.849f
C102 m2_39229_1610# m2_39425_1830# 0.251f
C103 carray_0.n7 m2_30325_9390# 0.452f
C104 dum sample 0.00816f
C105 m3_10329_1610# out 0.187f
C106 m2_3025_9390# out 0.849f
C107 m2_25125_9390# m3_24829_1610# 0.247f
C108 carray_0.n2 out 3.35f
C109 ctl1 ctl0 0.193f
C110 m3_41529_1610# m3_41729_1610# 3.35f
C111 m3_31129_1610# m2_31429_1610# 0.181f
C112 carray_0.n6 m3_36529_1610# 1.99f
C113 m2_425_4350# m2_425_3510# 0.199f
C114 m3_35229_1610# m3_36329_1610# 0.148f
C115 carray_0.n7 m2_32925_1830# 1.18e-19
C116 carray_0.ndum dum 0.107f
C117 carray_0.n7 m2_425_1830# 1.18e-19
C118 m2_23629_1610# m3_23529_1610# 2.11f
C119 m3_41729_1610# out 0.187f
C120 m3_36329_1610# out 0.187f
C121 m2_425_3510# out 0.719f
C122 carray_0.n6 m3_33729_1610# 0.00746f
C123 carray_0.n6 m2_16025_1830# 1.52e-19
C124 carray_0.n6 m3_16829_1610# 0.181f
C125 carray_0.n7 m2_4325_1830# 0.452f
C126 carray_0.n5 m2_6329_1610# 2.05e-19
C127 m2_38125_1830# out 0.643f
C128 m3_5129_1610# m2_5029_1610# 2.11f
C129 m2_14725_9390# m2_15429_1610# 0.251f
C130 m2_38125_1830# m3_38929_1610# 0.247f
C131 m2_43325_2670# vin 0.0183f
C132 m3_39129_1610# out 0.187f
C133 carray_0.n5 vdd 0.304f
C134 carray_0.n5 m2_10825_1830# 0.452f
C135 m3_32629_1610# out 0.187f
C136 m2_43325_3510# out 0.764f
C137 m3_38929_1610# m3_39129_1610# 3.35f
C138 m2_16025_9390# out 0.849f
C139 m2_425_7710# out 0.719f
C140 m3_32429_1610# m3_32629_1610# 3.35f
C141 m3_43029_1610# vin 9.27e-20
C142 m2_13425_9390# m3_13129_1610# 0.247f
C143 m3_42829_1610# out 0.187f
C144 carray_0.n7 m3_3829_1610# 0.181f
C145 m2_43325_4350# m2_43325_3510# 0.199f
C146 carray_0.ndum m2_14129_1610# 3.15e-20
C147 carray_0.n7 m3_30029_1610# 2.16f
C148 m2_34225_1830# m3_33929_1610# 0.247f
C149 m2_31625_9390# out 0.849f
C150 m3_4029_1610# m3_5129_1610# 0.148f
C151 carray_0.n5 m3_15529_1610# 0.181f
C152 carray_0.n7 m3_28729_1610# 1.98f
C153 m2_31625_9390# m3_32429_1610# 0.247f
C154 m2_425_8550# m2_425_7710# 0.199f
C155 m3_31129_1610# m3_31329_1610# 3.35f
C156 carray_0.n5 m3_26129_1610# 0.00889f
C157 carray_0.n2 m2_23629_1610# 0.247f
C158 ctl1 sample 0.00255f
C159 carray_0.n1 m2_9525_1830# 9.38e-20
C160 carray_0.n5 m3_11629_1610# 1.98f
C161 carray_0.n7 m3_9229_1610# 4.08f
C162 m3_27229_1610# m3_26129_1610# 0.148f
C163 carray_0.n1 m2_3729_1610# 8.05e-20
C164 m3_29829_1610# m2_29025_1830# 0.247f
C165 carray_0.n1 m2_22525_1830# 0.251f
C166 carray_0.n7 m2_2429_1610# 2.39f
C167 carray_0.n4 m2_8929_1610# 3.19e-19
C168 m3_28729_1610# m2_29025_9390# 0.247f
C169 carray_0.ndum m2_11529_1610# 3.15e-20
C170 m2_31429_1610# m2_31625_9390# 0.251f
C171 en_buf vdd 1.53f
C172 carray_0.n6 m2_23825_1830# 1.52e-19
C173 m2_39229_1610# sample 6.55e-20
C174 carray_0.n2 m3_5129_1610# 0.021f
C175 ctl0 carray_0.n0 0.107f
C176 carray_0.n3 m2_425_1830# 0.00133f
C177 carray_0.n7 m2_20629_1610# 1.05e-19
C178 carray_0.n7 m3_41529_1610# 0.00642f
C179 m2_425_6870# m2_1129_1610# 0.251f
C180 carray_0.n7 m3_35229_1610# 2.16f
C181 m3_10329_1610# m3_10529_1610# 3.35f
C182 m2_23825_9390# out 0.849f
C183 carray_0.n2 m3_10529_1610# 0.021f
C184 carray_0.n3 m3_20729_1610# 0.174f
C185 m3_6629_1610# m2_6925_1830# 0.247f
C186 carray_0.n3 m2_4325_1830# 4.28e-19
C187 m3_19429_1610# m3_18329_1610# 0.148f
C188 vin m2_43325_8550# 0.04f
C189 carray_0.n2 m2_3025_1830# 0.169f
C190 carray_0.n4 m2_6925_1830# 2.85e-19
C191 carray_0.n7 m2_38125_9390# 0.452f
C192 carray_0.n6 m2_29025_1830# 1.52e-19
C193 carray_0.n0 m2_8929_1610# 6.36e-20
C194 out m2_43325_9390# 0.932f
C195 carray_0.n7 out 97.1f
C196 m2_24929_1610# m2_25125_1830# 0.251f
C197 m2_41829_1610# m3_41529_1610# 0.181f
C198 m3_5329_1610# out 0.187f
C199 carray_0.n4 sample 5.55e-19
C200 carray_0.n7 m3_38929_1610# 4.08f
C201 m2_43325_3510# m2_43129_1610# 0.251f
C202 carray_0.n5 m2_12829_1610# 2.05e-19
C203 out m3_24629_1610# 0.187f
C204 m3_42829_1610# m2_43129_1610# 0.181f
C205 out m2_29025_9390# 0.849f
C206 m2_41829_1610# out 0.267f
C207 carray_0.n7 m2_31429_1610# 1.13f
C208 carray_0.ndum carray_0.n4 0.0771f
C209 m2_25125_1830# m3_25929_1610# 0.247f
C210 m3_31329_1610# m2_31625_9390# 0.247f
C211 m2_43325_7710# vin 0.0358f
C212 m2_30325_9390# m2_30129_1610# 0.251f
C213 m3_36329_1610# m3_36529_1610# 3.35f
C214 carray_0.n3 m2_2429_1610# 5.59e-19
C215 carray_0.n2 m2_16025_1830# 0.169f
C216 carray_0.n0 sample 0.00854f
C217 carray_0.n2 m3_16829_1610# 0.021f
C218 carray_0.n7 m2_1725_9390# 0.452f
C219 m2_23825_1830# m3_23529_1610# 0.247f
C220 m2_23629_1610# m2_23825_9390# 0.251f
C221 m2_20629_1610# carray_0.n3 1.09f
C222 carray_0.n6 m2_17325_9390# 0.452f
C223 carray_0.n6 m3_18129_1610# 1.98f
C224 carray_0.n0 carray_0.ndum 14.5f
C225 carray_0.n7 m2_23629_1610# 1.05e-19
C226 m3_33929_1610# out 0.187f
C227 m2_35525_9390# m2_35329_1610# 0.251f
C228 carray_0.n3 out 6.38f
C229 m2_16729_1610# out 0.267f
C230 m2_43129_1610# m2_43325_9390# 0.251f
C231 m2_43325_1830# out 0.64f
C232 m3_17029_1610# out 0.187f
C233 carray_0.n7 m2_43129_1610# 1.13f
C234 m2_23629_1610# m3_24629_1610# 0.0061f
C235 m3_32629_1610# m3_33729_1610# 0.148f
C236 m2_43325_3510# m2_43325_2670# 0.199f
C237 carray_0.n7 m3_5129_1610# 2.16f
C238 m2_16025_9390# m3_16829_1610# 0.247f
C239 carray_0.n7 m3_31329_1610# 0.181f
C240 m3_5129_1610# m3_5329_1610# 3.35f
C241 carray_0.n1 m2_425_1830# 9.38e-20
C242 m3_43029_1610# m2_43325_3510# 0.247f
C243 carray_0.n7 m2_28829_1610# 2.39f
C244 m2_425_7710# m2_425_6870# 0.199f
C245 carray_0.n7 m2_40725_1830# 1.18e-19
C246 a_45464_6355# vdd 0.77f
C247 m3_7929_1610# m2_8929_1610# 0.0061f
C248 m3_42829_1610# m3_43029_1610# 3.35f
C249 carray_0.n6 m2_6329_1610# 1.13f
C250 m3_30029_1610# m2_30129_1610# 2.11f
C251 carray_0.n1 m2_4325_1830# 9.38e-20
C252 carray_0.n7 m2_3025_1830# 1.18e-19
C253 carray_0.n4 m2_9525_1830# 2.85e-19
C254 carray_0.n4 m2_3729_1610# 3.19e-19
C255 carray_0.n4 m3_19429_1610# 0.181f
C256 m2_28829_1610# m2_29025_9390# 0.251f
C257 carray_0.n4 m2_22525_1830# 2.21e-19
C258 m2_39425_1830# sample 9.23e-21
C259 carray_0.n6 vdd 0.305f
C260 carray_0.n6 m2_10825_1830# 1.52e-19
C261 carray_0.n2 m3_14229_1610# 0.021f
C262 m2_5625_1830# out 0.643f
C263 carray_0.n2 m3_24829_1610# 3.16e-19
C264 carray_0.n7 m3_36529_1610# 0.181f
C265 vdd vin 3.41f
C266 m2_24929_1610# out 0.267f
C267 m2_10825_9390# out 0.849f
C268 m3_7729_1610# m2_7629_1610# 2.11f
C269 carray_0.n3 m2_23629_1610# 1.09f
C270 m3_1229_1610# m2_425_2670# 0.247f
C271 ctl0 sample 0.00375f
C272 carray_0.n6 m3_26129_1610# 1.98f
C273 m2_39229_1610# m3_40229_1610# 0.0061f
C274 carray_0.n6 m3_11629_1610# 0.181f
C275 carray_0.n0 m2_3729_1610# 6.36e-20
C276 m2_42025_9390# m3_41729_1610# 0.247f
C277 m2_43325_1830# m2_43129_1610# 0.251f
C278 carray_0.n1 m2_2429_1610# 8.05e-20
C279 out m3_14429_1610# 0.187f
C280 carray_0.n7 m2_16025_1830# 1.18e-19
C281 ctl2 vdd 0.162f
C282 carray_0.n5 m2_13425_1830# 2.03e-19
C283 out m3_25929_1610# 0.187f
C284 out m2_30129_1610# 0.267f
C285 m3_43029_1610# m2_43325_9390# 0.247f
C286 carray_0.n7 m3_43029_1610# 0.181f
C287 ctl0 carray_0.ndum 0.00139f
C288 carray_0.n1 m2_20629_1610# 8.05e-20
C289 m2_26425_1830# sample 9.23e-21
C290 carray_0.n6 m3_6429_1610# 0.181f
C291 carray_0.n4 m2_19925_9390# 0.452f
C292 m2_26229_1610# m3_26129_1610# 2.11f
C293 carray_0.n5 m2_18029_1610# 2.05e-19
C294 m2_43325_6030# vin 0.0375f
C295 m2_43325_6870# out 0.871f
C296 carray_0.n3 m2_3025_1830# 4.28e-19
C297 carray_0.n6 m2_36629_1610# 2.39f
C298 m2_42025_9390# m3_42829_1610# 0.247f
C299 carray_0.n1 out 1.99f
C300 carray_0.ndum m2_8929_1610# 3.15e-20
C301 carray_0.n2 m3_18129_1610# 0.021f
C302 m2_35525_1830# m3_35229_1610# 0.247f
C303 m2_35525_9390# m3_36329_1610# 0.247f
C304 a_45464_2123# sample 0.192f
C305 carray_0.n5 m2_15429_1610# 1.13f
C306 carray_0.ndum m2_22525_9390# 0.247f
C307 carray_0.n6 m2_12829_1610# 2.39f
C308 carray_0.n7 m2_5625_9390# 0.452f
C309 m2_35525_1830# out 0.643f
C310 m3_5329_1610# m2_5625_9390# 0.247f
C311 enb en_buf 1.56f
C312 m2_36825_9390# m3_37629_1610# 0.247f
C313 carray_0.n7 m2_23825_1830# 1.18e-19
C314 m2_12125_1830# out 0.643f
C315 m2_43325_9390# m2_43325_8550# 0.199f
C316 m3_18329_1610# out 0.187f
C317 m2_23825_1830# m3_24629_1610# 0.247f
C318 m2_425_5190# m3_1229_1610# 0.247f
C319 m3_33729_1610# m3_33929_1610# 3.35f
C320 m2_43325_2670# m2_43325_1830# 0.199f
C321 carray_0.ndum sample 11.1f
C322 m2_16025_1830# m2_16729_1610# 0.251f
C323 carray_0.n3 m2_16025_1830# 4.28e-19
C324 carray_0.n7 m3_14229_1610# 2.16f
C325 m2_16729_1610# m3_16829_1610# 2.11f
C326 carray_0.n2 m2_6329_1610# 0.00855f
C327 m3_16829_1610# m3_17029_1610# 3.35f
C328 carray_0.n7 m3_24829_1610# 1.98f
C329 m3_43029_1610# m2_43325_1830# 0.247f
C330 m2_10825_9390# m3_10529_1610# 0.247f
C331 carray_0.n7 m2_29025_1830# 0.452f
C332 ctl5 carray_0.n5 0.106f
C333 carray_0.n4 m2_425_1830# 8.3e-19
C334 carray_0.n2 m2_10825_1830# 0.169f
C335 carray_0.n7 m2_42025_9390# 0.452f
C336 carray_0.n2 vdd 0.311f
C337 m2_425_9390# m3_1229_1610# 0.247f
C338 m3_24629_1610# m3_24829_1610# 3.35f
C339 m2_43325_6870# m2_43129_1610# 0.251f
C340 carray_0.n4 m3_20729_1610# 1.98f
C341 m2_14129_1610# out 0.267f
C342 carray_0.n4 m2_4325_1830# 2.85e-19
C343 carray_0.n6 m2_12125_9390# 0.452f
C344 carray_0.n2 m3_15529_1610# 0.021f
C345 m2_6925_9390# out 0.849f
C346 m2_41829_1610# m2_42025_9390# 0.251f
C347 m2_34029_1610# sample 6.55e-20
C348 ctl6 vdd 0.158f
C349 carray_0.n2 m3_11629_1610# 0.021f
C350 m2_11529_1610# out 0.267f
C351 carray_0.n5 m2_31625_1830# 0.0714f
C352 carray_0.n7 m2_35525_9390# 0.452f
C353 m3_7929_1610# m2_8225_9390# 0.247f
C354 m3_1229_1610# m2_1129_1610# 2.11f
C355 m2_39425_1830# m3_40229_1610# 0.247f
C356 m2_43325_3510# vdd 0.00801f
C357 carray_0.n6 m3_12929_1610# 1.98f
C358 carray_0.n0 m3_20729_1610# 3.12e-19
C359 carray_0.n5 m2_27529_1610# 2.39f
C360 m2_32729_1610# sample 6.55e-20
C361 m2_18625_9390# m3_19429_1610# 0.247f
C362 carray_0.n1 m2_3025_1830# 9.38e-20
C363 out m3_15729_1610# 0.187f
C364 carray_0.n7 m3_18129_1610# 0.181f
C365 m3_2729_1610# m2_3729_1610# 0.0061f
C366 carray_0.n2 m3_6429_1610# 0.021f
C367 carray_0.n5 m2_21225_1830# 1.57e-19
C368 carray_0.n4 m2_2429_1610# 3.19e-19
C369 m2_27529_1610# m3_27229_1610# 0.181f
C370 m2_39229_1610# out 0.267f
C371 m2_8929_1610# m2_8225_9390# 0.251f
C372 m3_11829_1610# out 0.187f
C373 m2_39229_1610# m3_38929_1610# 0.181f
C374 carray_0.n4 m2_20629_1610# 2.39f
C375 carray_0.n6 m3_7729_1610# 1.98f
C376 carray_0.n5 m2_18625_1830# 2.03e-19
C377 m2_22525_1830# sample 4.62e-21
C378 m2_43325_5190# out 0.798f
C379 carray_0.n2 m2_12829_1610# 0.00855f
C380 carray_0.n5 m2_7629_1610# 2.05e-19
C381 carray_0.n5 m3_27229_1610# 0.00889f
C382 m2_43325_5190# m2_43325_4350# 0.199f
C383 m2_36629_1610# m3_36329_1610# 0.181f
C384 m3_6629_1610# out 0.187f
C385 carray_0.ndum m2_3729_1610# 3.15e-20
C386 carray_0.n0 m2_2429_1610# 6.36e-20
C387 carray_0.n4 out 12.2f
C388 carray_0.ndum m2_22525_1830# 0.381f
C389 ctl3 vdd 0.158f
C390 carray_0.n6 m2_13425_1830# 1.52e-19
C391 carray_0.n1 m2_16025_1830# 9.38e-20
C392 m2_43325_6870# m3_43029_1610# 0.247f
C393 a_45464_6355# enb 0.00726f
C394 carray_0.n7 m2_6329_1610# 2.39f
C395 m2_36825_9390# out 0.849f
C396 m3_1429_1610# m2_2429_1610# 0.0061f
C397 m3_2529_1610# m2_1725_1830# 0.247f
C398 carray_0.n2 m3_1229_1610# 0.0361f
C399 m3_5329_1610# m2_6329_1610# 0.0061f
C400 carray_0.n0 m2_20629_1610# 1.98e-19
C401 m2_19329_1610# m2_18625_1830# 0.251f
C402 vdd m2_43325_9390# 0.0203f
C403 carray_0.n7 m2_10825_1830# 1.18e-19
C404 carray_0.n7 vdd 0.305f
C405 carray_0.n5 m2_19329_1610# 2.05e-19
C406 carray_0.n6 m2_18029_1610# 2.39f
C407 m2_13425_9390# out 0.849f
C408 carray_0.n6 m3_2529_1610# 0.181f
C409 m2_425_3510# m3_1229_1610# 0.247f
C410 m2_24929_1610# m3_24829_1610# 2.11f
C411 enb vin 1.1f
C412 carray_0.n0 out 0.921f
C413 m2_17325_9390# m3_17029_1610# 0.247f
C414 carray_0.n7 m3_15529_1610# 1.98f
C415 m2_17325_1830# out 0.643f
C416 m3_17029_1610# m3_18129_1610# 0.148f
C417 carray_0.n7 m3_26129_1610# 0.181f
C418 carray_0.n6 m2_15429_1610# 1.43e-19
C419 m3_1429_1610# out 0.187f
C420 m2_11529_1610# m3_10529_1610# 0.0061f
C421 m3_14229_1610# m3_14429_1610# 3.35f
C422 m2_425_7710# m3_1229_1610# 0.247f
C423 m3_24829_1610# m3_25929_1610# 0.148f
C424 m2_36825_1830# sample 9.23e-21
C425 m2_14725_1830# out 0.643f
C426 m2_43325_5190# m2_43129_1610# 0.251f
C427 carray_0.n4 m2_23629_1610# 2.39f
C428 carray_0.n7 m3_6429_1610# 1.98f
C429 m2_25125_1830# sample 9.23e-21
C430 m2_34225_1830# sample 9.23e-21
C431 m2_9525_9390# m2_10229_1610# 0.251f
C432 m2_27529_1610# m2_27725_1830# 0.251f
C433 m3_6429_1610# m3_5329_1610# 0.148f
C434 carray_0.n2 m3_12929_1610# 0.021f
C435 carray_0.n3 m2_6329_1610# 5.59e-19
C436 carray_0.n7 m2_36629_1610# 1.13f
C437 carray_0.n5 m2_32925_9390# 0.452f
C438 ctl5 carray_0.n6 0.00139f
C439 carray_0.n6 m2_40529_1610# 2.39f
C440 m2_40529_1610# m3_40429_1610# 2.11f
C441 m3_1429_1610# m2_1725_9390# 0.247f
C442 carray_0.n3 m2_10825_1830# 4.28e-19
C443 m2_43325_1830# vdd 0.0196f
C444 carray_0.n3 vdd 0.301f
C445 m2_43325_7710# m2_43325_6870# 0.199f
C446 carray_0.n7 m2_12829_1610# 1.13f
C447 carray_0.n5 m2_10229_1610# 1.13f
C448 carray_0.n0 m2_23629_1610# 6.79e-20
C449 carray_0.n5 m2_27725_1830# 0.523f
C450 m2_32925_1830# sample 9.23e-21
C451 carray_0.n2 m3_7729_1610# 0.021f
C452 carray_0.n4 m2_3025_1830# 2.85e-19
C453 m2_27725_9390# m3_27429_1610# 0.247f
C454 m2_27529_1610# m3_28529_1610# 0.0061f
C455 m2_39425_1830# out 0.643f
C456 m2_16025_1830# m3_15729_1610# 0.247f
C457 m3_16829_1610# m3_15729_1610# 0.148f
C458 m3_13129_1610# out 0.187f
C459 m2_39425_9390# m3_39129_1610# 0.247f
C460 ctl7 vdd 0.158f
C461 m2_8929_1610# m3_9229_1610# 0.181f
C462 carray_0.n7 m3_1229_1610# 0.181f
C463 m3_3829_1610# m3_2729_1610# 0.148f
C464 m2_5625_1830# m2_6329_1610# 0.251f
C465 carray_0.n6 m2_31625_1830# 0.452f
C466 m2_34029_1610# m2_34225_1830# 0.251f
C467 carray_0.n5 m3_29829_1610# 0.00889f
C468 carray_0.n2 m2_13425_1830# 0.169f
C469 carray_0.n5 m2_8225_1830# 2.03e-19
C470 carray_0.n2 m2_21225_9390# 0.247f
C471 carray_0.n5 m3_28529_1610# 4.09f
C472 carray_0.ndum m3_20729_1610# 1.58e-19
C473 m2_36825_9390# m3_36529_1610# 0.247f
C474 m3_7929_1610# out 0.187f
C475 carray_0.n7 m2_14725_9390# 0.452f
C476 carray_0.n6 m2_27529_1610# 1.13f
C477 m2_19329_1610# m3_19629_1610# 0.181f
C478 m2_43325_5190# m3_43029_1610# 0.247f
C479 m2_14129_1610# m3_14229_1610# 2.11f
C480 carray_0.n2 m2_18029_1610# 0.00855f
C481 carray_0.n5 m2_1725_1830# 2.03e-19
C482 carray_0.n6 m2_21225_1830# 1.17e-19
C483 m3_2729_1610# m2_2429_1610# 0.181f
C484 carray_0.n2 m3_2529_1610# 0.021f
C485 carray_0.n4 m2_16025_1830# 2.85e-19
C486 m2_26425_1830# out 0.643f
C487 m2_8929_1610# out 0.267f
C488 carray_0.n6 m2_18625_1830# 1.52e-19
C489 carray_0.n5 m2_19925_1830# 2.03e-19
C490 m2_22525_9390# out 0.849f
C491 carray_0.n5 carray_0.n6 17.4f
C492 carray_0.n2 m2_15429_1610# 0.00855f
C493 carray_0.n3 m2_12829_1610# 5.59e-19
C494 carray_0.n6 m3_27229_1610# 4.08f
C495 carray_0.n6 m2_7629_1610# 2.39f
C496 m2_10825_9390# m3_11629_1610# 0.247f
C497 m3_18129_1610# m3_18329_1610# 3.35f
C498 m2_18625_9390# out 0.849f
C499 carray_0.n7 m2_39425_9390# 0.452f
C500 carray_0.ndum m2_2429_1610# 3.15e-20
C501 a_45464_2123# out 0.286f
C502 m3_2729_1610# out 0.187f
C503 carray_0.n7 m3_12929_1610# 0.181f
C504 m2_32729_1610# m2_32925_1830# 0.251f
C505 m3_14429_1610# m3_15529_1610# 0.148f
C506 a_45464_6355# en_buf 0.00369f
C507 ctl4 vdd 0.158f
C508 carray_0.n1 m2_6329_1610# 8.05e-20
C509 m3_6429_1610# m2_5625_1830# 0.247f
C510 m2_6925_1830# out 0.643f
C511 m2_43325_6870# vdd 0.0106f
C512 carray_0.n5 m2_26229_1610# 0.002f
C513 carray_0.ndum m2_20629_1610# 9.94e-20
C514 m3_25929_1610# m3_26129_1610# 3.35f
C515 out sample 0.0106f
C516 carray_0.n1 m2_10825_1830# 9.38e-20
C517 carray_0.n1 vdd 0.306f
C518 m2_40725_9390# m2_40529_1610# 0.251f
C519 carray_0.n5 m2_30325_1830# 0.0714f
C520 carray_0.n4 m2_23825_1830# 0.541f
C521 carray_0.n6 m2_19329_1610# 1.43e-19
C522 m2_26229_1610# m3_27229_1610# 0.0061f
C523 carray_0.n7 m3_7729_1610# 0.181f
C524 en_buf vin 0.797f
C525 carray_0.ndum out 0.917f
C526 m2_31429_1610# sample 6.55e-20
C527 dum vdd 0.165f
C528 carray_0.n5 m2_1129_1610# 3.41e-19
C529 carray_0.n4 m3_24829_1610# 0.181f
C530 m2_43325_6870# m2_43325_6030# 0.199f
C531 ctl5 ctl6 0.193f
C532 carray_0.n7 m2_13425_1830# 0.452f
C533 m3_35029_1610# m2_34225_9390# 0.247f
C534 m3_3829_1610# m2_3729_1610# 2.11f
C535 carray_0.n5 m2_5029_1610# 2.05e-19
C536 m2_27725_1830# m3_28529_1610# 0.247f
C537 m2_13425_9390# m3_14229_1610# 0.247f
C538 m2_36825_1830# m3_37629_1610# 0.247f
C539 enb m2_43325_9390# 0.0244f
C540 m2_34029_1610# out 0.267f
C541 carray_0.n7 m2_18029_1610# 1.13f
C542 m2_9525_9390# m3_10329_1610# 0.247f
C543 m2_9525_1830# m3_9229_1610# 0.247f
C544 carray_0.n7 m3_2529_1610# 1.98f
C545 m2_23629_1610# sample 6.55e-20
C546 carray_0.n5 m3_31129_1610# 0.00889f
C547 carray_0.n2 m2_21225_1830# 0.352f
C548 sample m2_43129_1610# 3.33e-19
C549 carray_0.n7 m2_15429_1610# 2.39f
C550 carray_0.n1 m2_12829_1610# 8.05e-20
C551 m2_19925_9390# m3_20729_1610# 0.247f
C552 carray_0.n6 m2_27725_1830# 1.52e-19
C553 carray_0.n6 m2_10229_1610# 1.43e-19
C554 m2_19925_1830# m3_19629_1610# 0.247f
C555 carray_0.ndum m2_23629_1610# 1.34e-19
C556 m2_32729_1610# out 0.267f
C557 carray_0.n5 m3_10329_1610# 0.181f
C558 carray_0.n2 m2_18625_1830# 0.169f
C559 m2_14725_9390# m3_14429_1610# 0.247f
C560 m3_2729_1610# m2_3025_1830# 0.247f
C561 carray_0.n5 carray_0.n2 0.196f
C562 m2_32729_1610# m3_32429_1610# 0.181f
C563 m2_10825_1830# m2_11529_1610# 0.251f
C564 sample m2_28829_1610# 6.55e-20
C565 m3_9029_1610# m2_8225_1830# 0.247f
C566 m2_40725_1830# sample 9.23e-21
C567 carray_0.n2 m2_7629_1610# 0.00855f
C568 ctl1 vdd 0.158f
C569 m2_27725_9390# out 0.849f
C570 m2_9525_1830# out 0.643f
C571 m3_19429_1610# out 0.187f
C572 m2_3729_1610# out 0.267f
C573 m2_22525_1830# out 0.643f
C574 m2_12125_1830# m2_12829_1610# 0.251f
C575 carray_0.n3 m2_13425_1830# 4.28e-19
C576 ctl6 carray_0.n5 0.0166f
C577 carray_0.n6 m2_8225_1830# 1.52e-19
C578 carray_0.n3 m2_21225_9390# 0.452f
C579 m2_11529_1610# m3_11629_1610# 2.11f
C580 carray_0.n7 m2_40529_1610# 1.13f
C581 m3_15529_1610# m3_15729_1610# 3.35f
C582 m2_19329_1610# carray_0.n2 0.00869f
C583 carray_0.n3 m2_18029_1610# 5.59e-19
C584 m2_8225_9390# out 0.849f
C585 m2_18029_1610# m3_17029_1610# 0.0061f
C586 m3_6629_1610# m2_6329_1610# 0.181f
C587 carray_0.n5 m3_32629_1610# 1.99f
C588 m2_17325_1830# m3_18129_1610# 0.247f
C589 carray_0.n6 m2_1725_1830# 1.52e-19
C590 m3_27429_1610# out 0.187f
C591 carray_0.n5 m2_16025_9390# 0.452f
C592 m2_43325_5190# vdd 0.0208f
C593 m3_13129_1610# m3_14229_1610# 0.148f
C594 m2_425_2670# m2_1129_1610# 0.251f
C595 carray_0.n4 m2_6329_1610# 3.19e-19
C596 m2_19925_9390# m2_20629_1610# 0.251f
C597 a_45464_6355# vin 0.412f
C598 carray_0.n6 m2_19925_1830# 1.52e-19
C599 m3_11629_1610# m3_11829_1610# 3.35f
C600 carray_0.n4 m2_10825_1830# 2.85e-19
C601 carray_0.n4 vdd 0.303f
C602 carray_0.n6 m3_40429_1610# 1.99f
C603 carray_0.n3 m2_15429_1610# 5.59e-19
C604 m3_30029_1610# m2_30325_9390# 0.247f
C605 carray_0.n6 m3_35029_1610# 0.00746f
C606 m3_43029_1610# sample 0.0051f
C607 carray_0.n7 m2_31625_1830# 1.18e-19
C608 m2_19925_9390# out 0.849f
C609 m2_4325_9390# m2_5029_1610# 0.251f
C610 carray_0.n6 m2_37929_1610# 1.13f
C611 m3_40229_1610# out 0.187f
C612 m2_425_6030# out 0.719f
C613 carray_0.n6 m3_37829_1610# 0.188f
C614 carray_0.n0 m2_6329_1610# 6.36e-20
C615 carray_0.n7 m2_9525_9390# 0.452f
C616 carray_0.n7 m2_27529_1610# 1.05e-19
C617 m2_43325_6030# m2_43325_5190# 0.199f
C618 carray_0.n6 m2_26229_1610# 2.39f
C619 carray_0.n6 m2_35329_1610# 0.00135f
C620 m2_36825_1830# out 0.643f
C621 carray_0.n7 m2_21225_1830# 9.11e-20
C622 m3_35029_1610# m2_35329_1610# 0.181f
C623 m3_4029_1610# m2_4325_9390# 0.247f
C624 carray_0.n0 vdd 0.306f
C625 carray_0.n6 m2_30325_1830# 1.52e-19
C626 m2_37929_1610# m3_37829_1610# 2.11f
C627 m3_37629_1610# out 0.187f
C628 carray_0.n2 m2_425_2670# 0.0993f
C629 m2_25125_1830# out 0.643f
C630 carray_0.n7 m2_18625_1830# 0.452f
C631 m2_34225_1830# out 0.643f
C632 carray_0.n7 carray_0.n5 1.06f
C633 m3_6429_1610# m3_6629_1610# 3.35f
C634 m2_12829_1610# m3_11829_1610# 0.0061f
C635 m2_12125_1830# m3_12929_1610# 0.247f
C636 m2_10229_1610# m3_10329_1610# 2.11f
C637 m2_23825_1830# sample 9.23e-21
C638 m2_34029_1610# m3_33729_1610# 0.181f
C639 m2_30325_9390# out 0.849f
C640 carray_0.n2 m2_10229_1610# 0.00855f
C641 m2_3729_1610# m2_3025_1830# 0.251f
C642 carray_0.n7 m2_7629_1610# 1.13f
C643 carray_0.n2 m3_19629_1610# 0.0214f
C644 carray_0.n6 m2_1129_1610# 1.7e-19
C645 carray_0.n5 m3_24629_1610# 0.00889f
C646 m2_425_3510# m2_425_2670# 0.199f
C647 m2_425_5190# m2_1129_1610# 0.251f
C648 carray_0.n1 m2_13425_1830# 9.38e-20
C649 m2_20629_1610# m3_20729_1610# 2.11f
C650 m2_36629_1610# m2_36825_9390# 0.251f
C651 carray_0.n1 m2_21225_9390# 0.251f
C652 m2_32925_1830# out 0.643f
C653 carray_0.n6 m2_5029_1610# 1.43e-19
C654 carray_0.n4 m2_12829_1610# 3.19e-19
C655 m2_14725_1830# m3_15529_1610# 0.247f
C656 m2_15429_1610# m3_14429_1610# 0.0061f
C657 m2_425_1830# out 0.639f
C658 m2_32925_9390# m3_32629_1610# 0.247f
C659 m2_32729_1610# m3_33729_1610# 0.0061f
C660 sample m2_29025_1830# 9.23e-21
C661 carray_0.n7 m2_19329_1610# 2.39f
C662 carray_0.n2 m2_8225_1830# 0.169f
C663 carray_0.n1 m2_18029_1610# 8.05e-20
C664 m2_425_9390# m2_1129_1610# 0.251f
C665 m3_20729_1610# out 0.187f
C666 m2_4325_1830# out 0.643f
C667 carray_0.n2 m3_9029_1610# 0.021f
C668 carray_0.n3 m2_21225_1830# 0.453f
C669 carray_0.n2 m2_1725_1830# 0.169f
C670 m2_12125_9390# m3_11829_1610# 0.247f
C671 carray_0.n1 m2_15429_1610# 8.05e-20
C672 m2_40725_9390# carray_0.n6 0.452f
C673 carray_0.n0 m2_12829_1610# 6.36e-20
C674 m3_3829_1610# out 0.187f
C675 m2_40725_9390# m3_40429_1610# 0.247f
C676 m3_30029_1610# out 0.187f
C677 m2_19925_1830# carray_0.n2 0.169f
C678 carray_0.n6 m2_3025_9390# 0.452f
C679 carray_0.n3 m2_18625_1830# 4.28e-19
C680 carray_0.n5 m3_33929_1610# 0.181f
C681 carray_0.n5 carray_0.n3 0.161f
C682 m2_18029_1610# m3_18329_1610# 0.181f
C683 m3_7729_1610# m2_6925_9390# 0.247f
C684 carray_0.n6 carray_0.n2 0.39f
C685 carray_0.n7 m2_25125_9390# 0.452f
C686 m3_28729_1610# out 0.187f
C687 carray_0.n7 m2_34225_9390# 0.452f
C688 carray_0.n5 m2_16729_1610# 2.39f
C689 m2_39229_1610# m2_39425_9390# 0.251f
C690 ctl0 vdd 0.158f
C691 carray_0.n3 m2_7629_1610# 5.59e-19
C692 m3_9229_1610# out 0.187f
C693 m3_11829_1610# m3_12929_1610# 0.148f
C694 m2_14129_1610# m2_13425_1830# 0.251f
C695 m2_2429_1610# out 0.267f
C696 carray_0.n6 m3_41729_1610# 0.181f
C697 ctl5 ctl4 0.193f
C698 m3_1229_1610# m3_1429_1610# 3.35f
C699 m3_31129_1610# m2_30325_1830# 0.247f
C700 carray_0.n6 m3_36329_1610# 0.00746f
C701 ctl6 carray_0.n6 0.107f
C702 ctl7 carray_0.n5 3.35e-20
C703 m2_20629_1610# out 0.267f
C704 m3_41529_1610# out 0.187f
C705 carray_0.n6 m2_38125_1830# 0.0598f
C706 m2_425_4350# out 0.719f
C707 m2_36825_1830# m3_36529_1610# 0.247f
C708 carray_0.n2 ctl2 0.106f
C709 carray_0.n6 m3_39129_1610# 0.00746f
C710 m3_35229_1610# out 0.187f
C711 m2_19329_1610# carray_0.n3 5.59e-19
C712 carray_0.n6 m3_32629_1610# 0.181f
C713 carray_0.n7 m2_27725_1830# 1.18e-19
C714 carray_0.n7 m2_10229_1610# 2.39f
C715 m3_36529_1610# m3_37629_1610# 0.148f
C716 carray_0.n7 m2_4325_9390# 0.452f
C717 carray_0.n5 m2_5625_1830# 2.03e-19
C718 m2_37929_1610# m2_38125_1830# 0.251f
C719 m2_38125_9390# out 0.849f
C720 m3_36329_1610# m2_35329_1610# 0.0061f
C721 m3_4029_1610# m2_5029_1610# 0.0061f
C722 m3_5129_1610# m2_4325_1830# 0.247f
C723 m2_425_6870# m2_425_6030# 0.199f
C724 m2_38125_1830# m3_37829_1610# 0.247f
C725 carray_0.n6 m2_31625_9390# 0.452f
C726 m2_38125_9390# m3_38929_1610# 0.247f
C727 carray_0.n5 m2_24929_1610# 0.002f
C728 m2_26425_1830# m3_26129_1610# 0.247f
C729 m3_38929_1610# out 0.187f
C730 m2_43325_3510# vin 0.0351f
C731 m3_32429_1610# out 0.187f
C732 a_45464_2123# vdd 0.77f
C733 carray_0.n5 m2_10825_9390# 0.452f
C734 m2_43325_4350# out 0.776f
C735 m2_2429_1610# m2_1725_9390# 0.251f
C736 carray_0.n2 m2_1129_1610# 0.0102f
C737 m2_425_8550# out 0.722f
C738 m2_26425_9390# out 0.849f
C739 m2_12829_1610# m3_13129_1610# 0.181f
C740 m3_6629_1610# m3_7729_1610# 0.148f
C741 m2_34225_9390# m3_33929_1610# 0.247f
C742 carray_0.n7 m3_29829_1610# 4.08f
C743 m2_31429_1610# out 0.267f
C744 sample vdd 1.58f
C745 carray_0.n7 m2_8225_1830# 0.452f
C746 carray_0.n2 m3_23529_1610# 3.4f
C747 carray_0.n2 m2_5029_1610# 0.00855f
C748 m2_31429_1610# m3_32429_1610# 0.0061f
C749 carray_0.ndum m2_6329_1610# 3.15e-20
C750 carray_0.n5 m3_25929_1610# 0.00889f
C751 m2_425_3510# m2_1129_1610# 0.251f
C752 carray_0.n5 m2_30129_1610# 0.002f
C753 carray_0.n7 m3_9029_1610# 2.16f
C754 m3_29829_1610# m2_29025_9390# 0.247f
C755 carray_0.n1 m2_21225_1830# 0.251f
C756 carray_0.n7 m2_1725_1830# 0.452f
C757 m3_28729_1610# m2_28829_1610# 2.11f
C758 carray_0.n5 ctl4 0.00139f
C759 carray_0.n4 m2_13425_1830# 2.85e-19
C760 carray_0.ndum vdd 0.34f
C761 m2_43325_5190# enb 0.0247f
C762 m2_15429_1610# m3_15729_1610# 0.181f
C763 m2_1725_9390# out 0.849f
C764 m3_3829_1610# m2_3025_1830# 0.247f
C765 m2_32925_1830# m3_33729_1610# 0.247f
C766 carray_0.n2 m3_4029_1610# 0.021f
C767 carray_0.n7 m2_19925_1830# 1.18e-19
C768 carray_0.n1 m2_18625_1830# 9.38e-20
C769 carray_0.n7 m3_40429_1610# 0.181f
C770 carray_0.n1 carray_0.n5 0.0772f
C771 m3_41729_1610# m2_42025_1830# 0.247f
C772 carray_0.n7 carray_0.n6 22.1f
C773 m2_425_7710# m2_1129_1610# 0.251f
C774 carray_0.n7 m3_35029_1610# 4.08f
C775 carray_0.n4 m2_18029_1610# 3.19e-19
C776 m2_23629_1610# out 0.267f
C777 carray_0.n3 m2_10229_1610# 5.59e-19
C778 carray_0.n2 m3_10329_1610# 0.021f
C779 carray_0.n1 m2_7629_1610# 8.05e-20
C780 vin m2_43325_9390# 0.0292f
C781 carray_0.n7 m2_37929_1610# 2.39f
C782 out m2_43129_1610# 0.322f
C783 m2_24929_1610# m2_25125_9390# 0.251f
C784 m2_41829_1610# carray_0.n6 1.13f
C785 carray_0.n7 m3_37829_1610# 1.98f
C786 ctl2 ctl3 0.193f
C787 m3_5129_1610# out 0.187f
C788 m2_40725_1830# m3_41529_1610# 0.247f
C789 m2_43325_4350# m2_43129_1610# 0.251f
C790 carray_0.n4 m2_15429_1610# 3.19e-19
C791 carray_0.n0 m2_21225_9390# 0.247f
C792 m3_31329_1610# out 0.187f
C793 carray_0.n5 m2_12125_1830# 2.03e-19
C794 carray_0.n7 m2_26229_1610# 1.13f
C795 carray_0.n7 m2_35329_1610# 3.52f
C796 m2_18625_1830# m3_18329_1610# 0.247f
C797 m2_36629_1610# sample 6.55e-20
C798 m3_42829_1610# m2_42025_1830# 0.247f
C799 m3_31329_1610# m3_32429_1610# 0.148f
C800 out m2_28829_1610# 0.267f
C801 carray_0.n0 m2_18029_1610# 6.36e-20
C802 m2_40725_1830# out 0.643f
C803 carray_0.n1 m2_19329_1610# 8.05e-20
C804 carray_0.n7 m2_30325_1830# 0.452f
C805 carray_0.n3 m2_8225_1830# 4.28e-19
C806 m2_17325_1830# m2_18029_1610# 0.251f
C807 m3_10529_1610# out 0.187f
C808 m3_12929_1610# m3_13129_1610# 3.35f
C809 m2_25125_1830# m3_24829_1610# 0.247f
C810 m2_25125_9390# m3_25929_1610# 0.247f
C811 m2_3025_1830# out 0.643f
C812 m3_31329_1610# m2_31429_1610# 2.11f
C813 m3_1429_1610# m3_2529_1610# 0.148f
C814 carray_0.n3 m2_1725_1830# 4.28e-19
C815 carray_0.n0 m2_15429_1610# 6.36e-20
C816 m2_23825_9390# m3_23529_1610# 0.247f
C817 carray_0.ndum m2_12829_1610# 3.15e-20
C818 carray_0.n7 m2_1129_1610# 1.13f
C819 m3_36529_1610# out 0.187f
C820 carray_0.n5 m2_14129_1610# 2.05e-19
C821 ctl5 carray_0.n4 0.0164f
C822 m2_19925_1830# carray_0.n3 4.28e-19
C823 m2_19329_1610# m3_18329_1610# 0.0061f
C824 carray_0.n6 m3_33929_1610# 0.00746f
C825 carray_0.n6 m2_16729_1610# 1.13f
C826 carray_0.n6 carray_0.n3 0.314f
C827 carray_0.n6 m3_17029_1610# 4.08f
C828 m3_35029_1610# m3_33929_1610# 0.148f
C829 carray_0.n7 m2_5029_1610# 3.52f
C830 m3_5329_1610# m2_5029_1610# 0.181f
C831 m3_42829_1610# m3_41729_1610# 0.148f
C832 m2_14725_1830# m2_15429_1610# 0.251f
C833 m2_7629_1610# m2_6925_9390# 0.251f
C834 m2_43325_1830# vin 0.017f
C835 carray_0.n5 m2_11529_1610# 2.39f
C836 m3_33729_1610# out 0.187f
C837 m2_16025_1830# out 0.643f
C838 m3_23529_1610# m3_24629_1610# 0.148f
C839 m2_43325_2670# out 0.857f
C840 m3_16829_1610# out 0.187f
C841 carray_0.n7 m2_42025_1830# 0.503f
C842 m2_425_6870# out 0.719f
C843 m3_7729_1610# m3_7929_1610# 3.35f
C844 ctl7 carray_0.n6 0.0169f
C845 ctl1 carray_0.n5 3.35e-20
C846 m2_13425_1830# m3_13129_1610# 0.247f
C847 carray_0.n7 m3_4029_1610# 4.08f
C848 m3_43029_1610# out 0.215f
C849 carray_0.n7 m3_31129_1610# 4.08f
C850 carray_0.n5 m3_15729_1610# 4.08f
C851 carray_0.n2 ctl3 0.0164f
C852 carray_0.n3 ctl2 0.00139f
C853 m3_43029_1610# m2_43325_4350# 0.247f
C854 carray_0.n1 m2_10229_1610# 8.05e-20
C855 m2_41829_1610# m2_42025_1830# 0.251f
C856 carray_0.n7 m3_10329_1610# 1.98f
C857 carray_0.n6 m2_5625_1830# 1.52e-19
C858 m3_29829_1610# m2_30129_1610# 0.181f
C859 m3_28729_1610# m2_29025_1830# 0.247f
C860 carray_0.n7 carray_0.n2 0.781f
C861 carray_0.n6 m2_24929_1610# 1.43e-19
C862 carray_0.n4 m2_21225_1830# 2.21e-19
C863 carray_0.n2 m3_5329_1610# 0.021f
C864 carray_0.n3 m2_1129_1610# 0.00153f
C865 carray_0.n2 m3_24629_1610# 4.18e-19
C866 m2_5625_9390# out 0.849f
C867 carray_0.n7 m3_41729_1610# 1.99f
C868 carray_0.n7 m3_36329_1610# 4.08f
C869 carray_0.n4 m2_18625_1830# 2.85e-19
C870 m2_23825_1830# out 0.643f
C871 ctl6 carray_0.n7 0.00139f
C872 carray_0.n4 carray_0.n5 12.7f
C873 carray_0.n3 m3_23529_1610# 0.174f
C874 carray_0.n1 m2_8225_1830# 9.38e-20
C875 m3_7729_1610# m2_6925_1830# 0.247f
C876 carray_0.n3 m2_5029_1610# 5.59e-19
C877 m3_6629_1610# m2_7629_1610# 0.0061f
C878 carray_0.n4 m2_7629_1610# 3.19e-19
C879 carray_0.n6 m2_30129_1610# 1.43e-19
C880 out m2_43325_8550# 0.781f
C881 carray_0.n7 m2_38125_1830# 0.452f
C882 carray_0.n7 m3_39129_1610# 2.16f
C883 m2_41829_1610# m3_41729_1610# 2.11f
C884 carray_0.n0 m2_21225_1830# 0.381f
C885 carray_0.n1 m2_1725_1830# 9.38e-20
C886 m2_43325_2670# m2_43129_1610# 0.251f
C887 out m3_14229_1610# 0.187f
C888 out m3_24829_1610# 0.187f
C889 carray_0.n7 m3_42829_1610# 4.08f
C890 out m2_29025_1830# 0.643f
C891 m3_43029_1610# m2_43129_1610# 2.11f
C892 m2_42025_9390# out 0.849f
C893 carray_0.n1 m2_19925_1830# 9.38e-20
C894 carray_0.n1 carray_0.n6 0.0844f
C895 carray_0.n0 carray_0.n5 0.0775f
C896 a_45464_2123# enb 1e-20
C897 carray_0.n4 m2_19329_1610# 1.13f
C898 carray_0.n5 m2_17325_1830# 2.03e-19
C899 m2_26229_1610# m3_25929_1610# 0.181f
C900 m2_43325_6870# vin 0.0175f
C901 m3_2529_1610# m3_2729_1610# 3.35f
C902 carray_0.n0 m2_7629_1610# 6.36e-20
C903 m2_43325_7710# out 0.765f
C904 m2_30325_1830# m2_30129_1610# 0.251f
C905 carray_0.n2 carray_0.n3 20.7f
C906 m2_41829_1610# m3_42829_1610# 0.0061f
C907 carray_0.n6 m2_35525_1830# 0.0598f
C908 enb sample 0.834f
C909 carray_0.n2 m2_16729_1610# 0.00855f
C910 carray_0.n2 m3_17029_1610# 0.021f
C911 m2_35525_9390# m3_35229_1610# 0.247f
C912 carray_0.n5 m2_14725_1830# 2.03e-19
C913 m2_23629_1610# m2_23825_1830# 0.251f
C914 carray_0.n6 dum 6.25e-20
C915 carray_0.n6 m2_12125_1830# 0.452f
C916 m2_36825_1830# m2_36629_1610# 0.251f
C917 m2_35525_9390# out 0.849f
C918 m2_36629_1610# m3_37629_1610# 0.0061f
C919 carray_0.ndum m2_18029_1610# 3.15e-20
C920 carray_0.n0 m2_19329_1610# 6.36e-20
C921 m2_35525_1830# m2_35329_1610# 0.251f
C922 m2_17325_9390# out 0.849f
C923 m2_43129_1610# m2_43325_8550# 0.251f
C924 m3_18129_1610# out 0.187f
C925 m2_425_6030# m3_1229_1610# 0.247f
C926 m2_23825_9390# m3_24629_1610# 0.247f
C927 carray_0.n7 m3_5329_1610# 4.08f
C928 m2_16025_9390# m2_16729_1610# 0.251f
C929 carray_0.ndum m2_15429_1610# 3.15e-20
C930 m2_16025_1830# m3_16829_1610# 0.247f
C931 carray_0.n2 m2_5625_1830# 0.169f
C932 carray_0.n1 m2_1129_1610# 8.05e-20
C933 ctl6 ctl7 0.193f
C934 carray_0.n6 m2_14129_1610# 1.43e-19
C935 m3_43029_1610# m2_43325_2670# 0.247f
C936 carray_0.n7 m2_29025_9390# 0.452f
C937 carray_0.n2 m2_24929_1610# 1.36e-19
C938 carray_0.n7 m2_41829_1610# 2.39f
C939 m3_31129_1610# m2_30129_1610# 0.0061f
C940 carray_0.n1 m2_5029_1610# 8.05e-20
C941 carray_0.n6 m2_6925_9390# 0.452f
C942 carray_0.n4 m2_10229_1610# 3.19e-19
C943 m2_43325_7710# m2_43129_1610# 0.251f
C944 carray_0.n4 m3_19629_1610# 4.08f
C945 m2_28829_1610# m2_29025_1830# 0.251f
C946 carray_0.n6 m2_11529_1610# 1.13f
C947 m2_40529_1610# sample 6.55e-20
C948 carray_0.n2 m3_14429_1610# 0.021f
C949 m2_6329_1610# out 0.267f
C950 ctl0 carray_0.n5 4.89e-20
C951 ctl1 carray_0.n6 1.31e-19
C952 m2_10825_1830# out 0.643f
C953 out vdd 1.6f
C954 carray_0.n3 ctl3 0.106f
C955 m3_7929_1610# m2_7629_1610# 0.181f
C956 carray_0.n4 m2_8225_1830# 2.85e-19
C957 carray_0.n6 m2_39229_1610# 0.00135f
C958 m3_1229_1610# m2_425_1830# 0.247f
C959 m2_43325_4350# vdd 0.0212f
C960 m2_39425_9390# m3_40229_1610# 0.247f
C961 carray_0.n0 m2_10229_1610# 6.36e-20
C962 carray_0.n6 m3_11829_1610# 4.08f
C963 carray_0.n5 m2_8929_1610# 2.05e-19
C964 carray_0.n7 carray_0.n3 0.623f
C965 m2_31625_1830# sample 9.23e-21
C966 carray_0.n7 m3_33929_1610# 1.98f
C967 carray_0.n1 carray_0.n2 2.02f
C968 carray_0.n5 m2_26425_1830# 0.0714f
C969 carray_0.n7 m2_16729_1610# 1.05e-19
C970 out m3_15529_1610# 0.187f
C971 carray_0.n4 m2_1725_1830# 2.85e-19
C972 out m3_26129_1610# 0.187f
C973 m2_26425_1830# m3_27229_1610# 0.247f
C974 m3_43029_1610# m2_43325_8550# 0.247f
C975 m3_11629_1610# out 0.187f
C976 m2_27529_1610# sample 6.55e-20
C977 carray_0.n6 m3_6629_1610# 4.08f
C978 m2_26425_9390# m3_26129_1610# 0.247f
C979 carray_0.n4 m2_19925_1830# 0.453f
C980 m2_43325_5190# vin 0.0325f
C981 carray_0.n4 carray_0.n6 0.318f
C982 m2_43325_6030# out 0.764f
C983 ctl7 carray_0.n7 0.107f
C984 carray_0.n2 m2_12125_1830# 0.169f
C985 carray_0.n6 m2_36825_9390# 0.452f
C986 carray_0.n5 m2_6925_1830# 2.03e-19
C987 carray_0.n2 m3_18329_1610# 0.021f
C988 m3_6429_1610# out 0.187f
C989 m2_35525_1830# m3_36329_1610# 0.247f
C990 carray_0.n5 sample 0.0017f
C991 m2_6925_1830# m2_7629_1610# 0.251f
C992 m2_43325_7710# m3_43029_1610# 0.247f
C993 carray_0.n7 m2_5625_1830# 0.452f
C994 m3_1429_1610# m2_1725_1830# 0.247f
C995 m2_36629_1610# out 0.267f
C996 m3_5329_1610# m2_5625_1830# 0.247f
C997 carray_0.n7 m2_24929_1610# 2.39f
C998 carray_0.n0 carray_0.n6 0.0803f
C999 vdd m2_43129_1610# 0.0238f
C1000 carray_0.ndum carray_0.n5 0.0767f
C1001 a_45464_2123# en_buf 0.00185f
C1002 m2_19329_1610# m2_18625_9390# 0.251f
C1003 m2_12829_1610# out 0.267f
C1004 carray_0.n6 m2_17325_1830# 0.452f
C1005 carray_0.ndum m2_7629_1610# 3.15e-20
C1006 carray_0.n2 m2_14129_1610# 0.00855f
C1007 m2_425_4350# m3_1229_1610# 0.247f
C1008 m2_24929_1610# m3_24629_1610# 0.181f
C1009 carray_0.n3 m2_16729_1610# 5.59e-19
C1010 en_buf sample 0.264f
C1011 m2_16729_1610# m3_17029_1610# 0.181f
C1012 carray_0.n7 m3_14429_1610# 4.08f
C1013 carray_0.n7 m3_25929_1610# 4.08f
C1014 ctl3 ctl4 0.193f
C1015 m3_1229_1610# out 0.187f
C1016 carray_0.n6 m2_14725_1830# 1.52e-19
C1017 m2_10825_1830# m3_10529_1610# 0.247f
C1018 carray_0.n7 m2_30129_1610# 3.52f
C1019 carray_0.n4 m2_1129_1610# 8.3e-19
C1020 carray_0.n2 m2_11529_1610# 0.00855f
C1021 m2_425_8550# m3_1229_1610# 0.247f
C1022 carray_0.ndum m2_19329_1610# 3.15e-20
C1023 carray_0.n5 m2_34029_1610# 1.13f
C1024 carray_0.n4 m3_23529_1610# 1.99f
C1025 m2_43325_7710# m2_43325_8550# 0.199f
C1026 m2_43325_6030# m2_43129_1610# 0.251f
C1027 carray_0.n4 m2_5029_1610# 3.19e-19
C1028 m2_14725_9390# out 0.849f
C1029 carray_0.n7 carray_0.n1 11.4f
C1030 carray_0.n2 m3_15729_1610# 0.021f
C1031 m3_10529_1610# m3_11629_1610# 0.148f
C1032 m2_27529_1610# m2_27725_9390# 0.251f
C1033 carray_0.n2 m3_11829_1610# 0.021f
C1034 carray_0.n3 m2_5625_1830# 4.28e-19
C1035 carray_0.n0 m2_1129_1610# 6.36e-20
C1036 m2_12125_9390# out 0.849f
C1037 carray_0.n7 m2_35525_1830# 0.452f
C1038 carray_0.n5 m2_32729_1610# 2.39f
C1039 m3_7929_1610# m2_8225_1830# 0.247f
C1040 carray_0.n6 m2_39425_1830# 0.0598f
C1041 m2_40529_1610# m3_40229_1610# 0.181f
C1042 m3_1429_1610# m2_1129_1610# 0.181f
C1043 m2_43325_2670# vdd 0.0108f
C1044 carray_0.n0 m3_23529_1610# 1.58e-19
C1045 carray_0.n0 m2_5029_1610# 6.36e-20
C1046 carray_0.n7 dum 2.59e-19
C1047 carray_0.n7 m2_12125_1830# 1.18e-19
C1048 m3_7929_1610# m3_9029_1610# 0.148f
C1049 carray_0.n5 m2_9525_1830# 2.03e-19
C1050 m2_18625_1830# m3_19429_1610# 0.247f
C1051 carray_0.n5 m2_27725_9390# 0.452f
C1052 m3_43029_1610# vdd 0.00943f
C1053 carray_0.n7 m3_18329_1610# 4.08f
C1054 carray_0.n5 m2_3729_1610# 2.05e-19
C1055 carray_0.n2 m3_6629_1610# 0.021f
C1056 carray_0.n5 m2_22525_1830# 1.57e-19
C1057 m2_27529_1610# m3_27429_1610# 2.11f
C1058 m2_8929_1610# m2_8225_1830# 0.251f
C1059 m2_39425_9390# out 0.849f
C1060 carray_0.n4 carray_0.n2 0.144f
C1061 m2_16025_9390# m3_15729_1610# 0.247f
C1062 m3_12929_1610# out 0.187f
C1063 m2_39229_1610# m3_39129_1610# 2.11f
C1064 m2_27725_1830# sample 9.23e-21
C1065 ctl0 carray_0.n6 1.31e-19
C1066 m2_8929_1610# m3_9029_1610# 2.11f
C1067 m2_5625_9390# m2_6329_1610# 0.251f
C1068 carray_0.n3 ctl4 0.0164f
C1069 m2_34029_1610# m2_34225_9390# 0.251f
C1070 ctl6 carray_0.n4 1.72e-20
C1071 carray_0.n5 m3_27429_1610# 1.99f
C1072 carray_0.ndum m2_10229_1610# 3.15e-20
C1073 carray_0.n7 m2_14129_1610# 3.52f
C1074 m2_36629_1610# m3_36529_1610# 2.11f
C1075 m3_7729_1610# out 0.187f
C1076 carray_0.n6 m2_8929_1610# 1.43e-19
C1077 m2_19329_1610# m3_19429_1610# 2.11f
C1078 carray_0.n6 m2_26425_1830# 0.452f
C1079 m3_27229_1610# m3_27429_1610# 3.35f
C1080 carray_0.n1 carray_0.n3 3.36f
C1081 carray_0.n0 carray_0.n2 1.42f
C1082 m2_43325_6030# m3_43029_1610# 0.247f
C1083 carray_0.n1 m2_16729_1610# 8.05e-20
C1084 carray_0.n2 m2_17325_1830# 0.169f
C1085 m3_2529_1610# m2_2429_1610# 2.11f
C1086 carray_0.n2 m3_1429_1610# 0.021f
C1087 vdd m2_43325_8550# 0.0226f
C1088 carray_0.n7 m2_11529_1610# 1.05e-19
C1089 m2_13425_1830# out 0.643f
C1090 ctl1 carray_0.n7 0.0172f
C1091 carray_0.n6 m3_2729_1610# 4.08f
C1092 ctl7 carray_0.n1 0.00139f
C1093 a_45464_6355# sample 0.192f
C1094 m2_21225_9390# out 0.849f
C1095 carray_0.n2 m2_14725_1830# 0.169f
C1096 m2_24929_1610# m3_25929_1610# 0.0061f
C1097 carray_0.n3 m2_12125_1830# 4.28e-19
C1098 m2_26425_1830# m2_26229_1610# 0.251f
C1099 carray_0.n6 m2_6925_1830# 0.452f
C1100 m2_17325_9390# m3_18129_1610# 0.247f
C1101 enb out 0.978f
C1102 a_45464_2123# vin 0.365f
C1103 m2_18029_1610# out 0.267f
C1104 carray_0.n6 sample 0.0059f
C1105 carray_0.n7 m2_39229_1610# 3.52f
C1106 m3_2529_1610# out 0.187f
C1107 m2_32729_1610# m2_32925_9390# 0.251f
C1108 m2_43325_4350# enb 0.0258f
C1109 carray_0.n1 m2_5625_1830# 9.38e-20
C1110 m3_6429_1610# m2_5625_9390# 0.247f
C1111 m2_43325_7710# vdd 0.00874f
C1112 sample vin 0.346f
C1113 carray_0.n5 m2_25125_1830# 0.0714f
C1114 m2_425_6870# m3_1229_1610# 0.247f
C1115 m2_37929_1610# sample 6.55e-20
C1116 m2_15429_1610# out 0.267f
C1117 carray_0.ndum carray_0.n6 0.0782f
C1118 carray_0.n4 ctl3 0.00139f
C1119 carray_0.n4 m2_23825_9390# 0.452f
C1120 carray_0.n3 m2_14129_1610# 5.59e-19
C1121 m2_35329_1610# sample 6.55e-20
C1122 m2_26229_1610# sample 6.55e-20
C1123 m2_9525_1830# m2_10229_1610# 0.251f
C1124 carray_0.n2 m3_13129_1610# 0.021f
C1125 carray_0.n7 carray_0.n4 0.678f
C1126 m2_30325_1830# sample 9.23e-21
C1127 m3_19429_1610# m3_19629_1610# 3.35f
C1128 carray_0.n5 m2_32925_1830# 0.523f
C1129 carray_0.n5 m2_425_1830# 0.00136f
C1130 m3_2529_1610# m2_1725_9390# 0.247f
C1131 carray_0.n4 m3_24629_1610# 4.08f
C1132 m2_40529_1610# m3_41529_1610# 0.0061f
C1133 carray_0.n3 m2_11529_1610# 5.59e-19
C1134 carray_0.n7 m2_13425_9390# 0.452f
C1135 carray_0.n6 m2_34029_1610# 0.00135f
C1136 carray_0.n2 m3_7929_1610# 0.021f
C1137 m3_35029_1610# m2_34029_1610# 0.0061f
C1138 carray_0.n5 m2_4325_1830# 2.03e-19
C1139 m2_27725_9390# m3_28529_1610# 0.247f
C1140 m2_27725_1830# m3_27429_1610# 0.247f
C1141 m2_40529_1610# out 0.267f
C1142 carray_0.n7 carray_0.n0 0.0953f
C1143 enb m2_43129_1610# 0.00743f
C1144 m2_16729_1610# m3_15729_1610# 0.0061f
C1145 m2_39425_1830# m3_39129_1610# 0.247f
C1146 carray_0.n7 m2_17325_1830# 1.18e-19
C1147 carray_0.n7 m3_1429_1610# 4.08f
C1148 m2_9525_9390# m3_9229_1610# 0.247f
C1149 ctl7 ctl1 0.193f
C1150 carray_0.n2 m2_8929_1610# 0.00855f
C1151 carray_0.ndum m2_1129_1610# 3.15e-20
C1152 carray_0.n6 m2_32729_1610# 1.13f
C1153 carray_0.n5 m3_30029_1610# 0.00889f
C1154 carray_0.n2 m2_22525_9390# 0.247f
C1155 carray_0.n5 m3_28729_1610# 0.19f
C1156 sample m2_42025_1830# 9.23e-21
C1157 carray_0.ndum m3_23529_1610# 3.12e-19
C1158 carray_0.n7 m2_14725_1830# 0.452f
C1159 carray_0.ndum m2_5029_1610# 3.15e-20
C1160 carray_0.n1 dum 1.97e-19
C1161 carray_0.n1 m2_12125_1830# 9.38e-20
C1162 carray_0.n6 m2_9525_1830# 1.52e-19
C1163 m2_19925_9390# m3_19629_1610# 0.247f
C1164 m3_27429_1610# m3_28529_1610# 0.148f
C1165 m2_31625_1830# out 0.643f
C1166 m2_14129_1610# m3_14429_1610# 0.181f
C1167 carray_0.n6 m2_3729_1610# 2.39f
C1168 carray_0.n6 m2_22525_1830# 1.17e-19
C1169 m3_2729_1610# m2_3025_9390# 0.247f
C1170 carray_0.n5 m2_2429_1610# 2.05e-19
C1171 carray_0.n2 m3_2729_1610# 0.021f
C1172 carray_0.n4 m2_16729_1610# 3.19e-19
C1173 m2_10825_9390# m2_11529_1610# 0.251f
C1174 carray_0.n4 carray_0.n3 12.1f
C1175 m2_31625_1830# m3_32429_1610# 0.247f
C1176 m3_9029_1610# m2_8225_9390# 0.247f
C1177 m2_9525_9390# out 0.849f
C1178 m2_27529_1610# out 0.267f
C1179 carray_0.n2 m2_6925_1830# 0.169f
C1180 carray_0.n5 m2_20629_1610# 2.05e-19
C1181 m2_31625_1830# m2_31429_1610# 0.251f
C1182 m2_21225_1830# out 0.643f
C1183 carray_0.n6 m3_27429_1610# 0.181f
C1184 ctl7 carray_0.n4 1.72e-20
C1185 m2_10825_1830# m3_11629_1610# 0.247f
C1186 m2_18625_1830# out 0.643f
C1187 carray_0.n1 m2_14129_1610# 8.05e-20
C1188 carray_0.n7 m2_39425_1830# 0.452f
C1189 carray_0.n5 out 24.3f
C1190 carray_0.n0 m2_16729_1610# 6.36e-20
C1191 carray_0.n7 m3_13129_1610# 4.08f
C1192 carray_0.n0 carray_0.n3 1.36f
C1193 carray_0.ndum carray_0.n2 1.42f
C1194 carray_0.n3 m2_17325_1830# 4.28e-19
C1195 m3_27229_1610# out 0.187f
C1196 carray_0.n5 m3_32429_1610# 0.00889f
C1197 m3_6429_1610# m2_6329_1610# 2.11f
C1198 m2_17325_1830# m3_17029_1610# 0.247f
C1199 m2_7629_1610# out 0.267f
C1200 m2_43325_6030# vdd 0.0178f
C1201 m2_425_2670# m2_425_1830# 0.199f
C1202 m3_43029_1610# enb 0.00364f
C1203 carray_0.n4 m2_5625_1830# 2.85e-19
C1204 m2_38125_1830# sample 9.23e-21
C1205 carray_0.n1 m2_11529_1610# 8.05e-20
C1206 m2_26425_9390# m3_27229_1610# 0.247f
C1207 carray_0.n5 m2_31429_1610# 0.002f
C1208 carray_0.n4 m2_24929_1610# 1.13f
C1209 m2_40725_1830# m2_40529_1610# 0.251f
C1210 carray_0.n6 m3_40229_1610# 0.00746f
C1211 m3_40229_1610# m3_40429_1610# 3.35f
C1212 ctl1 carray_0.n1 0.107f
C1213 ctl0 carray_0.n7 1.64e-19
C1214 carray_0.n3 m2_14725_1830# 4.28e-19
C1215 carray_0.n7 m3_7929_1610# 4.08f
C1216 m2_425_6030# m2_425_5190# 0.199f
C1217 m3_42829_1610# sample 0.0051f
C1218 en_buf out 0.58f
C1219 m2_19329_1610# out 0.267f
C1220 m3_19629_1610# m3_20729_1610# 0.148f
C1221 carray_0.n6 m2_36825_1830# 0.512f
C1222 m2_31625_1830# m3_31329_1610# 0.247f
C1223 carray_0.n6 m3_37629_1610# 4.09f
C1224 carray_0.n7 m2_8929_1610# 3.52f
C1225 carray_0.n7 m2_26425_1830# 1.18e-19
C1226 carray_0.n6 m2_34225_1830# 0.0598f
C1227 carray_0.n6 m2_25125_1830# 1.52e-19
C1228 carray_0.n4 ctl4 0.106f
C1229 m3_35029_1610# m2_34225_1830# 0.247f
C1230 m3_4029_1610# m2_3729_1610# 0.181f
C1231 carray_0.n5 m2_23629_1610# 2.05e-19
C1232 m2_37929_1610# m3_37629_1610# 0.181f
C1233 m2_13425_1830# m3_14229_1610# 0.247f
C1234 enb m2_43325_8550# 0.0236f
C1235 m3_37629_1610# m3_37829_1610# 3.35f
C1236 carray_0.n7 m2_18625_9390# 0.452f
C1237 m2_25125_9390# out 0.849f
C1238 m2_34225_9390# out 0.849f
C1239 carray_0.n1 carray_0.n4 0.0766f
C1240 m2_12125_1830# m3_11829_1610# 0.247f
C1241 m2_9525_1830# m3_10329_1610# 0.247f
C1242 m2_10229_1610# m3_9229_1610# 0.0061f
C1243 carray_0.n2 m2_9525_1830# 0.169f
C1244 carray_0.n7 m2_6925_1830# 1.18e-19
C1245 carray_0.n6 m2_32925_1830# 1.52e-19
C1246 carray_0.n2 m2_3729_1610# 0.00855f
C1247 carray_0.n5 m3_31329_1610# 0.00889f
C1248 carray_0.n2 m3_19429_1610# 0.0213f
C1249 m2_3729_1610# m2_3025_9390# 0.251f
C1250 carray_0.n6 m2_425_1830# 1.52e-19
C1251 carray_0.n2 m2_22525_1830# 0.352f
C1252 m3_29829_1610# m3_30029_1610# 3.35f
C1253 carray_0.n7 sample 4.96f
C1254 m2_425_6030# m2_1129_1610# 0.251f
C1255 carray_0.n5 m2_28829_1610# 1.14f
C1256 m3_29829_1610# m3_28729_1610# 0.148f
C1257 m2_19925_1830# m3_20729_1610# 0.247f
C1258 m3_28529_1610# m3_28729_1610# 3.35f
C1259 m2_20629_1610# m3_19629_1610# 0.0061f
C1260 m2_32925_9390# out 0.849f
C1261 carray_0.n5 m3_10529_1610# 4.08f
C1262 carray_0.n6 m2_4325_1830# 1.52e-19
C1263 carray_0.n4 m2_12125_1830# 2.85e-19
C1264 m2_14725_1830# m3_14429_1610# 0.247f
C1265 m2_14725_9390# m3_15529_1610# 0.247f
C1266 carray_0.n5 m2_3025_1830# 2.03e-19
C1267 m2_425_2670# out 0.719f
C1268 m2_32729_1610# m3_32629_1610# 2.11f
C1269 carray_0.n1 carray_0.n0 14.5f
C1270 carray_0.n7 carray_0.ndum 0.177f
C1271 m2_41829_1610# sample 6.55e-20
C1272 carray_0.n1 m2_17325_1830# 9.38e-20
C1273 m2_10229_1610# out 0.267f
C1274 m2_27725_1830# out 0.643f
C1275 m2_4325_9390# out 0.849f
C1276 m3_19629_1610# out 0.187f
C1277 carray_0.n6 m3_3829_1610# 1.98f
C1278 m3_9029_1610# m3_9229_1610# 3.35f
C1279 carray_0.n3 m2_8929_1610# 5.59e-19
C1280 m2_1725_1830# m2_2429_1610# 0.251f
C1281 carray_0.n3 m2_22525_9390# 0.452f
C1282 m2_11529_1610# m3_11829_1610# 0.181f
C1283 carray_0.n0 dum 0.0178f
C1284 carray_0.n1 m2_14725_1830# 9.38e-20
C1285 carray_0.n4 m2_14129_1610# 3.19e-19
C1286 m3_29829_1610# out 0.187f
C1287 carray_0.n6 m2_2429_1610# 1.13f
C1288 carray_0.n5 m3_33729_1610# 4.08f
C1289 m2_18029_1610# m2_17325_9390# 0.251f
C1290 m3_28529_1610# out 0.187f
C1291 m2_8225_1830# out 0.643f
C1292 carray_0.n7 m2_34029_1610# 2.39f
C1293 m3_6629_1610# m2_6925_9390# 0.247f
C1294 m2_18029_1610# m3_18129_1610# 2.11f
C1295 carray_0.n5 m3_16829_1610# 1.98f
C1296 carray_0.n5 m2_16025_1830# 0.452f
C1297 m2_425_1830# m2_1129_1610# 0.251f
C1298 m2_19925_1830# m2_20629_1610# 0.251f
C1299 carray_0.n3 m2_6925_1830# 4.28e-19
C1300 m3_9029_1610# out 0.187f
C1301 carray_0.n6 m2_20629_1610# 1.43e-19
C1302 m2_1725_1830# out 0.643f
C1303 m2_14129_1610# m2_13425_9390# 0.251f
C1304 carray_0.n4 m2_11529_1610# 3.19e-19
C1305 carray_0.n3 sample 3.92e-19
C1306 m2_43325_1830# sample 0.0408f
C1307 carray_0.n6 m3_41529_1610# 4.08f
C1308 m3_40429_1610# m3_41529_1610# 0.148f
C1309 a_45464_6355# out 0.29f
C1310 m3_31129_1610# m2_30325_9390# 0.247f
C1311 m3_30029_1610# m2_30325_1830# 0.247f
C1312 carray_0.n6 m3_35229_1610# 0.00746f
C1313 m2_425_5190# m2_425_4350# 0.199f
C1314 ctl1 carray_0.n4 1.72e-20
C1315 m3_35029_1610# m3_35229_1610# 3.35f
C1316 carray_0.n7 m2_32729_1610# 1.05e-19
C1317 m2_19925_1830# out 0.643f
C1318 carray_0.n0 m2_14129_1610# 6.36e-20
.ends

