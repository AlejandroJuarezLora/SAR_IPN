magic
tech sky130B
magscale 1 2
timestamp 1696358972
<< nwell >>
rect -226 -284 226 284
<< pmos >>
rect -30 -136 30 64
<< pdiff >>
rect -88 34 -30 64
rect -88 -106 -76 34
rect -42 -106 -30 34
rect -88 -136 -30 -106
rect 30 34 88 64
rect 30 -106 42 34
rect 76 -106 88 34
rect 30 -136 88 -106
<< pdiffc >>
rect -76 -106 -42 34
rect 42 -106 76 34
<< nsubdiff >>
rect -190 214 190 248
rect -190 -214 -156 214
rect 156 -214 190 214
rect -190 -248 -75 -214
rect 75 -248 190 -214
<< nsubdiffcont >>
rect -75 -248 75 -214
<< poly >>
rect -33 145 33 161
rect -33 111 -17 145
rect 17 111 33 145
rect -33 95 33 111
rect -30 64 30 95
rect -30 -162 30 -136
<< polycont >>
rect -17 111 17 145
<< locali >>
rect -33 111 -17 145
rect 17 111 33 145
rect -76 34 -42 50
rect -76 -122 -42 -106
rect 42 34 76 50
rect 42 -122 76 -106
rect -91 -248 -75 -214
rect 75 -248 91 -214
<< viali >>
rect -17 111 17 145
rect -76 -106 -42 34
rect 42 -89 76 17
<< metal1 >>
rect -29 145 29 157
rect -29 111 -17 145
rect 17 111 29 145
rect -29 99 29 111
rect -82 34 -36 46
rect -82 -106 -76 34
rect -42 -106 -36 34
rect 36 17 82 29
rect 36 -89 42 17
rect 76 -89 82 17
rect 36 -101 82 -89
rect -82 -118 -36 -106
<< labels >>
flabel metal1 -29 99 29 157 0 FreeSans 480 0 0 0 G
port 2 nsew
flabel metal1 -82 -118 -76 46 0 FreeSans 480 0 0 0 D
port 0 nsew
flabel metal1 76 -101 82 29 0 FreeSans 480 0 0 0 S
port 1 nsew
flabel locali 2 -232 2 -231 0 FreeSans 480 0 0 0 B
port 3 nsew
<< properties >>
string FIXED_BBOX -173 -231 173 231
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.3 m 1 nf 1 diffcov 80 polycov 80 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 80 rlcov 80 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 60 viadrn 80 viagate 80 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
