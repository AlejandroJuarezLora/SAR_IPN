magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect 0 269 536 590
<< pwell >>
rect 49 29 487 211
<< scnmos >>
rect 127 55 157 185
rect 211 55 241 185
rect 295 55 325 185
rect 379 55 409 185
<< scpmoshvt >>
rect 127 305 157 505
rect 211 305 241 505
rect 295 305 325 505
rect 379 305 409 505
<< ndiff >>
rect 75 101 127 185
rect 75 67 83 101
rect 117 67 127 101
rect 75 55 127 67
rect 157 109 211 185
rect 157 75 167 109
rect 201 75 211 109
rect 157 55 211 75
rect 241 101 295 185
rect 241 67 251 101
rect 285 67 295 101
rect 241 55 295 67
rect 325 109 379 185
rect 325 75 335 109
rect 369 75 379 109
rect 325 55 379 75
rect 409 102 461 185
rect 409 68 419 102
rect 453 68 461 102
rect 409 55 461 68
<< pdiff >>
rect 75 493 127 505
rect 75 459 83 493
rect 117 459 127 493
rect 75 425 127 459
rect 75 391 83 425
rect 117 391 127 425
rect 75 357 127 391
rect 75 323 83 357
rect 117 323 127 357
rect 75 305 127 323
rect 157 493 211 505
rect 157 459 167 493
rect 201 459 211 493
rect 157 425 211 459
rect 157 391 167 425
rect 201 391 211 425
rect 157 357 211 391
rect 157 323 167 357
rect 201 323 211 357
rect 157 305 211 323
rect 241 493 295 505
rect 241 459 251 493
rect 285 459 295 493
rect 241 425 295 459
rect 241 391 251 425
rect 285 391 295 425
rect 241 305 295 391
rect 325 493 379 505
rect 325 459 335 493
rect 369 459 379 493
rect 325 425 379 459
rect 325 391 335 425
rect 369 391 379 425
rect 325 357 379 391
rect 325 323 335 357
rect 369 323 379 357
rect 325 305 379 323
rect 409 493 461 505
rect 409 459 419 493
rect 453 459 461 493
rect 409 305 461 459
<< ndiffc >>
rect 83 67 117 101
rect 167 75 201 109
rect 251 67 285 101
rect 335 75 369 109
rect 419 68 453 102
<< pdiffc >>
rect 83 459 117 493
rect 83 391 117 425
rect 83 323 117 357
rect 167 459 201 493
rect 167 391 201 425
rect 167 323 201 357
rect 251 459 285 493
rect 251 391 285 425
rect 335 459 369 493
rect 335 391 369 425
rect 335 323 369 357
rect 419 459 453 493
<< poly >>
rect 127 505 157 531
rect 211 505 241 531
rect 295 505 325 531
rect 379 505 409 531
rect 127 273 157 305
rect 211 273 241 305
rect 295 273 325 305
rect 379 273 409 305
rect 59 257 409 273
rect 59 223 75 257
rect 109 223 167 257
rect 201 223 251 257
rect 285 223 335 257
rect 369 223 409 257
rect 59 207 409 223
rect 127 185 157 207
rect 211 185 241 207
rect 295 185 325 207
rect 379 185 409 207
rect 127 29 157 55
rect 211 29 241 55
rect 295 29 325 55
rect 379 29 409 55
<< polycont >>
rect 75 223 109 257
rect 167 223 201 257
rect 251 223 285 257
rect 335 223 369 257
<< locali >>
rect 38 535 67 569
rect 101 535 159 569
rect 193 535 251 569
rect 285 535 343 569
rect 377 535 435 569
rect 469 535 498 569
rect 64 493 117 535
rect 64 459 83 493
rect 64 425 117 459
rect 64 391 83 425
rect 64 357 117 391
rect 64 323 83 357
rect 64 307 117 323
rect 151 493 217 501
rect 151 459 167 493
rect 201 459 217 493
rect 151 425 217 459
rect 151 391 167 425
rect 201 391 217 425
rect 151 357 217 391
rect 251 493 285 535
rect 251 425 285 459
rect 251 375 285 391
rect 319 493 385 501
rect 319 459 335 493
rect 369 459 385 493
rect 319 425 385 459
rect 419 493 461 535
rect 453 459 461 493
rect 419 443 461 459
rect 319 391 335 425
rect 369 391 385 425
rect 151 323 167 357
rect 201 341 217 357
rect 319 357 385 391
rect 319 341 335 357
rect 201 323 335 341
rect 369 345 385 357
rect 369 323 472 345
rect 151 307 472 323
rect 59 257 385 273
rect 59 223 75 257
rect 109 223 167 257
rect 201 223 251 257
rect 285 223 335 257
rect 369 223 385 257
rect 419 189 472 307
rect 151 153 472 189
rect 64 101 117 117
rect 64 67 83 101
rect 64 25 117 67
rect 151 109 217 153
rect 151 75 167 109
rect 201 75 217 109
rect 151 59 217 75
rect 251 101 285 117
rect 251 25 285 67
rect 319 109 385 153
rect 319 75 335 109
rect 369 75 385 109
rect 319 59 385 75
rect 419 102 469 118
rect 453 68 469 102
rect 419 25 469 68
rect 38 -9 67 25
rect 101 -9 159 25
rect 193 -9 251 25
rect 285 -9 343 25
rect 377 -9 435 25
rect 469 -9 498 25
<< viali >>
rect 67 535 101 569
rect 159 535 193 569
rect 251 535 285 569
rect 343 535 377 569
rect 435 535 469 569
rect 67 -9 101 25
rect 159 -9 193 25
rect 251 -9 285 25
rect 343 -9 377 25
rect 435 -9 469 25
<< metal1 >>
rect 38 569 498 600
rect 38 535 67 569
rect 101 535 159 569
rect 193 535 251 569
rect 285 535 343 569
rect 377 535 435 569
rect 469 535 498 569
rect 38 504 498 535
rect 38 25 498 56
rect 38 -9 67 25
rect 101 -9 159 25
rect 193 -9 251 25
rect 285 -9 343 25
rect 377 -9 435 25
rect 469 -9 498 25
rect 38 -40 498 -9
<< labels >>
rlabel comment s 38 8 38 8 4 inv_4
flabel comment s 452 178 452 178 0 FreeSans 340 0 0 0 Y
flabel comment s 452 246 452 246 0 FreeSans 340 0 0 0 Y
flabel comment s 452 314 452 314 0 FreeSans 340 0 0 0 Y
flabel comment s 84 246 84 246 0 FreeSans 340 0 0 0 A
flabel comment s 176 246 176 246 0 FreeSans 340 0 0 0 A
flabel comment s 268 246 268 246 0 FreeSans 340 0 0 0 A
flabel comment s 360 246 360 246 0 FreeSans 340 0 0 0 A
<< properties >>
string FIXED_BBOX 38 8 498 552
string path 0.950 0.200 12.450 0.200 
<< end >>
