magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_p >>
rect 15 -25 49 9
<< viali >>
rect 15 -25 49 9
<< metal1 >>
rect 0 -34 6 18
rect 58 -34 64 18
<< via1 >>
rect 6 9 58 18
rect 6 -25 15 9
rect 15 -25 49 9
rect 49 -25 58 9
rect 6 -34 58 -25
<< metal2 >>
rect 6 18 58 24
rect 6 -40 58 -34
<< end >>
