magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 314 542
<< pwell >>
rect 1 -19 275 143
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 197 117
<< scpmoshvt >>
rect 79 283 197 457
<< ndiff >>
rect 27 74 79 117
rect 27 40 35 74
rect 69 40 79 74
rect 27 7 79 40
rect 197 74 249 117
rect 197 40 207 74
rect 241 40 249 74
rect 197 7 249 40
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 350 79 411
rect 27 316 35 350
rect 69 316 79 350
rect 27 283 79 316
rect 197 445 249 457
rect 197 411 207 445
rect 241 411 249 445
rect 197 350 249 411
rect 197 316 207 350
rect 241 316 249 350
rect 197 283 249 316
<< ndiffc >>
rect 35 40 69 74
rect 207 40 241 74
<< pdiffc >>
rect 35 411 69 445
rect 35 316 69 350
rect 207 411 241 445
rect 207 316 241 350
<< poly >>
rect 79 457 197 483
rect 79 253 197 283
rect 79 251 117 253
rect 51 235 117 251
rect 51 201 67 235
rect 101 201 117 235
rect 51 185 117 201
rect 159 195 225 211
rect 159 161 175 195
rect 209 161 225 195
rect 159 145 225 161
rect 159 143 197 145
rect 79 117 197 143
rect 79 -19 197 7
<< polycont >>
rect 67 201 101 235
rect 175 161 209 195
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 276 521
rect 17 445 259 487
rect 17 411 35 445
rect 69 411 207 445
rect 241 411 259 445
rect 17 350 259 411
rect 17 316 35 350
rect 69 316 207 350
rect 241 316 259 350
rect 17 269 259 316
rect 17 201 67 235
rect 101 201 121 235
rect 17 127 121 201
rect 155 195 259 269
rect 155 161 175 195
rect 209 161 259 195
rect 17 74 259 127
rect 17 40 35 74
rect 69 40 207 74
rect 241 40 259 74
rect 17 -23 259 40
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 276 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
<< metal1 >>
rect 0 521 276 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 276 521
rect 0 456 276 487
rect 0 -23 276 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 276 -23
rect 0 -88 276 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 decap_3
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
<< properties >>
string FIXED_BBOX 0 -40 276 504
string path 0.000 -1.000 6.900 -1.000 
<< end >>
