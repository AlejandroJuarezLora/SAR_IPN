magic
tech sky130B
timestamp 1696364841
<< metal2 >>
rect 0 54 40 60
rect 0 26 6 54
rect 34 26 40 54
rect 0 14 40 26
rect 0 -14 6 14
rect 34 -14 40 14
rect 0 -20 40 -14
<< via2 >>
rect 6 26 34 54
rect 6 -14 34 14
<< metal3 >>
rect 0 54 40 60
rect 0 26 6 54
rect 34 26 40 54
rect 0 14 40 26
rect 0 -14 6 14
rect 34 -14 40 14
rect 0 -20 40 -14
<< end >>
