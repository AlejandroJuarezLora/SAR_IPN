magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 498 542
<< pwell >>
rect 182 117 456 163
rect 1 -19 456 117
rect 30 -57 64 -19
<< scnmos >>
rect 79 7 109 91
rect 163 7 193 91
rect 264 7 294 137
rect 348 7 378 137
<< scpmoshvt >>
rect 91 257 121 341
rect 163 257 193 341
rect 264 257 294 457
rect 348 257 378 457
<< ndiff >>
rect 208 91 264 137
rect 27 63 79 91
rect 27 29 35 63
rect 69 29 79 63
rect 27 7 79 29
rect 109 63 163 91
rect 109 29 119 63
rect 153 29 163 63
rect 109 7 163 29
rect 193 63 264 91
rect 193 29 219 63
rect 253 29 264 63
rect 193 7 264 29
rect 294 90 348 137
rect 294 56 304 90
rect 338 56 348 90
rect 294 7 348 56
rect 378 55 430 137
rect 378 21 388 55
rect 422 21 430 55
rect 378 7 430 21
<< pdiff >>
rect 208 447 264 457
rect 208 413 220 447
rect 254 413 264 447
rect 208 379 264 413
rect 208 345 220 379
rect 254 345 264 379
rect 208 341 264 345
rect 39 309 91 341
rect 39 275 47 309
rect 81 275 91 309
rect 39 257 91 275
rect 121 257 163 341
rect 193 257 264 341
rect 294 445 348 457
rect 294 411 304 445
rect 338 411 348 445
rect 294 377 348 411
rect 294 343 304 377
rect 338 343 348 377
rect 294 257 348 343
rect 378 445 430 457
rect 378 411 388 445
rect 422 411 430 445
rect 378 257 430 411
<< ndiffc >>
rect 35 29 69 63
rect 119 29 153 63
rect 219 29 253 63
rect 304 56 338 90
rect 388 21 422 55
<< pdiffc >>
rect 220 413 254 447
rect 220 345 254 379
rect 47 275 81 309
rect 304 411 338 445
rect 304 343 338 377
rect 388 411 422 445
<< poly >>
rect 264 457 294 483
rect 348 457 378 483
rect 91 341 121 367
rect 163 341 193 367
rect 91 225 121 257
rect 25 209 121 225
rect 25 175 35 209
rect 69 175 121 209
rect 25 159 121 175
rect 163 225 193 257
rect 264 225 294 257
rect 348 225 378 257
rect 163 209 217 225
rect 163 175 173 209
rect 207 175 217 209
rect 163 159 217 175
rect 264 209 378 225
rect 264 175 289 209
rect 323 175 378 209
rect 264 159 378 175
rect 79 91 109 159
rect 163 91 193 159
rect 264 137 294 159
rect 348 137 378 159
rect 79 -19 109 7
rect 163 -19 193 7
rect 264 -19 294 7
rect 348 -19 378 7
<< polycont >>
rect 35 175 69 209
rect 173 175 207 209
rect 289 175 323 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 220 447 254 487
rect 220 379 254 413
rect 31 309 103 328
rect 220 327 254 345
rect 288 445 354 453
rect 288 411 304 445
rect 338 411 354 445
rect 288 377 354 411
rect 388 445 422 487
rect 388 395 422 411
rect 288 343 304 377
rect 338 361 354 377
rect 338 343 443 361
rect 288 327 443 343
rect 31 275 47 309
rect 81 293 103 309
rect 81 275 323 293
rect 31 259 323 275
rect 30 209 69 225
rect 30 175 35 209
rect 30 113 69 175
rect 103 79 139 259
rect 173 209 255 225
rect 207 175 255 209
rect 173 113 255 175
rect 289 209 323 259
rect 289 159 323 175
rect 357 125 443 327
rect 304 91 443 125
rect 304 90 338 91
rect 21 63 69 79
rect 21 29 35 63
rect 21 -23 69 29
rect 103 63 161 79
rect 103 29 119 63
rect 153 29 161 63
rect 103 11 161 29
rect 207 63 270 79
rect 207 29 219 63
rect 253 29 270 63
rect 304 37 338 56
rect 372 55 438 57
rect 207 -23 270 29
rect 372 21 388 55
rect 422 21 438 55
rect 372 -23 438 21
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
<< metal1 >>
rect 0 521 460 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 0 456 460 487
rect 0 -23 460 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
rect 0 -88 460 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 or2_2
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 30 181 64 215 0 FreeSans 200 0 0 0 B
port 9 nsew
flabel locali s 398 317 432 351 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 214 181 248 215 0 FreeSans 200 0 0 0 A
port 8 nsew
<< properties >>
string FIXED_BBOX 0 -40 460 504
string path 0.000 12.600 11.500 12.600 
<< end >>
