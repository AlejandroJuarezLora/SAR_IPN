* NGSPICE file created from sw_top_flat.ext - technology: sky130B

.subckt sw_top out en vss in vdd
X0 out.t9 a_456_1956# in.t1 vdd.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 out.t8 a_456_1956# in.t8 vdd.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 out.t19 a_456_865# in.t19 vss.t21 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 vss.t6 vdd.t22 vss.t5 vss sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4 vss.t11 a_456_1956# a_456_865# vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 out.t18 a_456_865# in.t10 vss.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 vss.t4 vdd.t23 vss.t3 vss sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X7 out.t7 a_456_1956# in.t5 vdd.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X8 a_456_865# a_456_1956# vss.t10 vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X9 in.t2 a_456_1956# out.t6 vdd.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X10 vdd.t13 a_456_1956# a_456_865# w_0_349# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 vdd.t21 vss.t22 vdd.t20 w_0_349# sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X12 in.t17 a_456_865# out.t17 vss.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X13 a_456_865# a_456_1956# vdd.t12 w_0_349# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X14 vdd.t19 vss.t23 vdd.t18 w_0_349# sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X15 in.t6 a_456_1956# out.t5 vdd.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X16 out.t16 a_456_865# in.t11 vss.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X17 in.t3 a_456_1956# out.t4 vdd.t10 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X18 out.t15 a_456_865# in.t12 vss.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X19 in.t13 a_456_865# out.t14 vss.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X20 vdd.t0 en.t0 a_456_1956# w_0_349# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X21 vss.t9 a_456_1956# a_456_865# vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 out.t3 a_456_1956# in.t7 vdd.t9 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X23 in.t14 a_456_865# out.t13 vss.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X24 a_456_1956# en.t1 vdd.t3 w_0_349# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 vdd.t1 en.t2 a_456_1956# w_0_349# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 a_456_865# a_456_1956# vss.t8 vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 a_456_1956# en.t3 vdd.t2 w_0_349# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X28 in.t4 a_456_1956# out.t2 vdd.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X29 out.t12 a_456_865# in.t15 vss.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X30 vdd.t7 a_456_1956# a_456_865# w_0_349# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X31 vss.t1 en.t4 a_456_1956# vss sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 in.t0 a_456_1956# out.t1 vdd.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X33 a_456_865# a_456_1956# vdd.t5 w_0_349# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 in.t16 a_456_865# out.t11 vss.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X35 a_456_1956# en.t5 vss.t2 vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 out.t0 a_456_1956# in.t9 vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X37 vss.t0 en.t6 a_456_1956# vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X38 in.t18 a_456_865# out.t10 vss.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X39 a_456_1956# en.t7 vss.t7 vss sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 in.n0 in.t0 36.7058
R1 in.n18 in.t7 36.7048
R2 in.n10 in.t9 28.5655
R3 in.n10 in.t2 28.5655
R4 in.n13 in.t1 28.5655
R5 in.n13 in.t6 28.5655
R6 in.n4 in.t8 28.5655
R7 in.n4 in.t3 28.5655
R8 in.n1 in.t5 28.5655
R9 in.n1 in.t4 28.5655
R10 in.n18 in.t15 24.4699
R11 in.n0 in.t16 24.4699
R12 in.n11 in.t12 17.4005
R13 in.n11 in.t14 17.4005
R14 in.n14 in.t11 17.4005
R15 in.n14 in.t13 17.4005
R16 in.n5 in.t10 17.4005
R17 in.n5 in.t17 17.4005
R18 in.n2 in.t19 17.4005
R19 in.n2 in.t18 17.4005
R20 in.n12 in.n10 8.14039
R21 in.n15 in.n13 8.14039
R22 in.n6 in.n4 8.14039
R23 in.n3 in.n1 8.14039
R24 in.n3 in.n2 7.0705
R25 in.n6 in.n5 7.0705
R26 in.n15 in.n14 7.0705
R27 in.n12 in.n11 7.0705
R28 in.n17 in.n12 2.22302
R29 in.n16 in.n15 2.22302
R30 in.n7 in.n6 2.22302
R31 in.n8 in.n3 2.22302
R32 in.n9 in.n0 2.21834
R33 in.n19 in.n18 2.21834
R34 in in.n9 1.13902
R35 in in.n19 1.12727
R36 in.n8 in.n7 0.36925
R37 in.n17 in.n16 0.36925
R38 in.n9 in.n8 0.348417
R39 in.n19 in.n17 0.348417
R40 out.n7 out.t4 28.5655
R41 out.n7 out.t9 28.5655
R42 out.n11 out.t6 28.5655
R43 out.n11 out.t3 28.5655
R44 out.n14 out.t5 28.5655
R45 out.n14 out.t0 28.5655
R46 out.n3 out.t2 28.5655
R47 out.n3 out.t8 28.5655
R48 out.n0 out.t1 28.5655
R49 out.n0 out.t7 28.5655
R50 out.n8 out.t17 17.4005
R51 out.n8 out.t16 17.4005
R52 out.n12 out.t13 17.4005
R53 out.n12 out.t12 17.4005
R54 out.n15 out.t14 17.4005
R55 out.n15 out.t15 17.4005
R56 out.n4 out.t10 17.4005
R57 out.n4 out.t18 17.4005
R58 out.n1 out.t11 17.4005
R59 out.n1 out.t19 17.4005
R60 out.n9 out.n8 7.68993
R61 out.n13 out.n12 7.68953
R62 out.n16 out.n15 7.68953
R63 out.n5 out.n4 7.68953
R64 out.n2 out.n1 7.68953
R65 out.n16 out.n14 7.52136
R66 out.n2 out.n0 7.52136
R67 out.n5 out.n3 7.52136
R68 out.n13 out.n11 7.5213
R69 out.n9 out.n7 7.52096
R70 out.n17 out.n13 2.59177
R71 out.n6 out.n2 2.59177
R72 out.n17 out.n16 2.22302
R73 out.n6 out.n5 2.22302
R74 out.n10 out.n9 2.21834
R75 out out.n18 0.80675
R76 out.n10 out.n6 0.348417
R77 out.n18 out.n17 0.318208
R78 out.n18 out.n10 0.0171667
R79 vdd.n148 vdd.t7 584.644
R80 vdd.n159 vdd.t0 584.644
R81 vdd.n191 vdd.t21 242.135
R82 vdd.n170 vdd.t20 242.135
R83 vdd.n142 vdd.t18 234.554
R84 vdd.n145 vdd.t19 234.554
R85 vdd.n67 vdd.n66 210.739
R86 vdd.n153 vdd.n152 174.595
R87 vdd.n164 vdd.n163 174.595
R88 vdd.n141 vdd.t23 166.282
R89 vdd.n157 vdd.t12 151.123
R90 vdd.n168 vdd.t2 151.123
R91 vdd.n6 vdd.n5 92.5005
R92 vdd.n8 vdd.n7 92.5005
R93 vdd.n10 vdd.n9 92.5005
R94 vdd.n12 vdd.n11 92.5005
R95 vdd.n14 vdd.n13 92.5005
R96 vdd.n16 vdd.n15 92.5005
R97 vdd.n18 vdd.n17 92.5005
R98 vdd.n20 vdd.n19 92.5005
R99 vdd.n22 vdd.n21 92.5005
R100 vdd.n24 vdd.n23 92.5005
R101 vdd.n26 vdd.n25 92.5005
R102 vdd.n28 vdd.n27 92.5005
R103 vdd.n30 vdd.n29 92.5005
R104 vdd.n32 vdd.n31 92.5005
R105 vdd.n34 vdd.n33 92.5005
R106 vdd.n36 vdd.n35 92.5005
R107 vdd.n38 vdd.n37 92.5005
R108 vdd.n40 vdd.n39 92.5005
R109 vdd.n78 vdd.n77 92.5005
R110 vdd.n74 vdd.n73 92.5005
R111 vdd.n1 vdd.n0 92.5005
R112 vdd.n4 vdd.n3 92.5005
R113 vdd.n131 vdd.n130 92.5005
R114 vdd.n129 vdd.n128 92.5005
R115 vdd.n128 vdd.n127 92.5005
R116 vdd.n126 vdd.n125 92.5005
R117 vdd.n125 vdd.n124 92.5005
R118 vdd.n123 vdd.n122 92.5005
R119 vdd.n122 vdd.n121 92.5005
R120 vdd.n120 vdd.n119 92.5005
R121 vdd.n119 vdd.n118 92.5005
R122 vdd.n117 vdd.n116 92.5005
R123 vdd.n116 vdd.n115 92.5005
R124 vdd.n114 vdd.n113 92.5005
R125 vdd.n113 vdd.n112 92.5005
R126 vdd.n111 vdd.n110 92.5005
R127 vdd.n110 vdd.n109 92.5005
R128 vdd.n108 vdd.n107 92.5005
R129 vdd.n107 vdd.n106 92.5005
R130 vdd.n105 vdd.n104 92.5005
R131 vdd.n104 vdd.n103 92.5005
R132 vdd.n102 vdd.n101 92.5005
R133 vdd.n101 vdd.n100 92.5005
R134 vdd.n99 vdd.n98 92.5005
R135 vdd.n98 vdd.n97 92.5005
R136 vdd.n96 vdd.n95 92.5005
R137 vdd.n95 vdd.n94 92.5005
R138 vdd.n93 vdd.n92 92.5005
R139 vdd.n92 vdd.n91 92.5005
R140 vdd.n90 vdd.n89 92.5005
R141 vdd.n89 vdd.n88 92.5005
R142 vdd.n87 vdd.n86 92.5005
R143 vdd.n86 vdd.n85 92.5005
R144 vdd.n84 vdd.n83 92.5005
R145 vdd.n83 vdd.n82 92.5005
R146 vdd.n80 vdd.n79 92.5005
R147 vdd.n81 vdd.n80 92.5005
R148 vdd.n6 vdd.n4 89.6005
R149 vdd.n81 vdd.n78 89.6005
R150 vdd.n48 vdd.n40 85.71
R151 vdd.n139 vdd.n131 83.9635
R152 vdd.n66 vdd.t9 78.6097
R153 vdd.n178 vdd.n177 76.0005
R154 vdd.n73 vdd.n72 72.7879
R155 vdd.n88 vdd.t15 65.2294
R156 vdd.n176 vdd.t22 50.5057
R157 vdd.n124 vdd.t14 48.504
R158 vdd.n3 vdd.n2 42.8997
R159 vdd.n77 vdd.n76 42.8996
R160 vdd.n135 vdd.n134 42.3534
R161 vdd.n103 vdd.t10 41.8139
R162 vdd.n106 vdd.t17 41.8139
R163 vdd.n82 vdd.t6 35.1237
R164 vdd.n76 vdd.n75 33.0686
R165 vdd.n152 vdd.t5 26.5955
R166 vdd.n152 vdd.t13 26.5955
R167 vdd.n163 vdd.t3 26.5955
R168 vdd.n163 vdd.t1 26.5955
R169 vdd.n8 vdd.n6 25.6005
R170 vdd.n10 vdd.n8 25.6005
R171 vdd.n12 vdd.n10 25.6005
R172 vdd.n14 vdd.n12 25.6005
R173 vdd.n16 vdd.n14 25.6005
R174 vdd.n18 vdd.n16 25.6005
R175 vdd.n20 vdd.n18 25.6005
R176 vdd.n22 vdd.n20 25.6005
R177 vdd.n24 vdd.n22 25.6005
R178 vdd.n26 vdd.n24 25.6005
R179 vdd.n28 vdd.n26 25.6005
R180 vdd.n30 vdd.n28 25.6005
R181 vdd.n32 vdd.n30 25.6005
R182 vdd.n34 vdd.n32 25.6005
R183 vdd.n36 vdd.n34 25.6005
R184 vdd.n38 vdd.n36 25.6005
R185 vdd.n40 vdd.n38 25.6005
R186 vdd.n4 vdd.n1 25.6005
R187 vdd.n78 vdd.n74 25.6005
R188 vdd.n84 vdd.n81 25.6005
R189 vdd.n87 vdd.n84 25.6005
R190 vdd.n90 vdd.n87 25.6005
R191 vdd.n93 vdd.n90 25.6005
R192 vdd.n96 vdd.n93 25.6005
R193 vdd.n99 vdd.n96 25.6005
R194 vdd.n102 vdd.n99 25.6005
R195 vdd.n105 vdd.n102 25.6005
R196 vdd.n108 vdd.n105 25.6005
R197 vdd.n111 vdd.n108 25.6005
R198 vdd.n114 vdd.n111 25.6005
R199 vdd.n117 vdd.n114 25.6005
R200 vdd.n120 vdd.n117 25.6005
R201 vdd.n123 vdd.n120 25.6005
R202 vdd.n126 vdd.n123 25.6005
R203 vdd.n129 vdd.n126 25.6005
R204 vdd.n131 vdd.n129 25.6005
R205 vdd.n44 vdd.n43 24.4976
R206 vdd.n52 vdd.n51 24.4976
R207 vdd.n53 vdd.n52 24.4976
R208 vdd.n45 vdd.n44 24.4976
R209 vdd.n65 vdd.n64 21.7962
R210 vdd.n64 vdd.n63 21.7962
R211 vdd.n91 vdd.t8 18.3984
R212 vdd.n118 vdd.t4 18.3984
R213 vdd.n136 vdd.n135 15.4044
R214 vdd.n97 vdd.t16 11.7082
R215 vdd.n112 vdd.t11 11.7082
R216 vdd.n69 vdd.n65 10.5887
R217 vdd.n58 vdd.n57 9.3005
R218 vdd.n60 vdd.n59 9.3005
R219 vdd.n56 vdd.n55 9.3005
R220 vdd.n55 vdd.n54 9.3005
R221 vdd.n47 vdd.n46 9.3005
R222 vdd.n70 vdd.n69 9.3005
R223 vdd.n138 vdd.n137 9.3005
R224 vdd.n177 vdd.n176 7.11866
R225 vdd.n42 vdd.n41 6.02403
R226 vdd.n50 vdd.n49 6.02403
R227 vdd.n62 vdd.n61 5.27109
R228 vdd.n144 vdd.n142 5.07505
R229 vdd.n192 vdd.n191 4.95526
R230 vdd.n169 vdd.n168 4.6505
R231 vdd.n160 vdd.n159 4.6505
R232 vdd.n158 vdd.n157 4.6505
R233 vdd.n149 vdd.n148 4.6505
R234 vdd.n144 vdd.n143 4.6505
R235 vdd.n147 vdd.n146 4.6505
R236 vdd.n172 vdd.n171 4.6505
R237 vdd.n175 vdd.n174 4.6505
R238 vdd.n180 vdd.n179 4.6505
R239 vdd.n183 vdd.n182 4.6505
R240 vdd.n185 vdd.n184 4.6505
R241 vdd.n187 vdd.n186 4.6505
R242 vdd.n189 vdd.n188 4.6505
R243 vdd.n167 vdd.n166 4.6505
R244 vdd.n165 vdd.n164 4.6505
R245 vdd.n162 vdd.n161 4.6505
R246 vdd.n156 vdd.n155 4.6505
R247 vdd.n154 vdd.n153 4.6505
R248 vdd.n151 vdd.n150 4.6505
R249 vdd.n69 vdd.n68 4.56271
R250 vdd.n133 vdd.n132 4.51815
R251 vdd.n68 vdd.n67 4.5125
R252 vdd.n46 vdd.n45 3.52991
R253 vdd.n54 vdd.n53 3.52991
R254 vdd.n56 vdd.n48 2.31034
R255 vdd.n190 vdd.n140 2.25407
R256 vdd.n140 vdd.n71 2.09329
R257 vdd.n140 vdd.n139 2.07952
R258 vdd.n139 vdd.n138 2.05645
R259 vdd.n138 vdd.n133 1.88285
R260 vdd.n71 vdd.n70 1.83953
R261 vdd.n48 vdd.n47 1.59246
R262 vdd.n70 vdd.n62 1.12991
R263 vdd.n174 vdd.n173 0.935332
R264 vdd.n142 vdd.n141 0.863992
R265 vdd.n137 vdd.n136 0.775333
R266 vdd.n179 vdd.n178 0.539826
R267 vdd.n47 vdd.n42 0.376971
R268 vdd.n55 vdd.n50 0.376971
R269 vdd.n146 vdd.n145 0.305262
R270 vdd.n171 vdd.n170 0.21623
R271 vdd.n182 vdd.n181 0.14432
R272 vdd.n147 vdd.n144 0.120292
R273 vdd.n149 vdd.n147 0.120292
R274 vdd.n151 vdd.n149 0.120292
R275 vdd.n154 vdd.n151 0.120292
R276 vdd.n156 vdd.n154 0.120292
R277 vdd.n158 vdd.n156 0.120292
R278 vdd.n160 vdd.n158 0.120292
R279 vdd.n162 vdd.n160 0.120292
R280 vdd.n165 vdd.n162 0.120292
R281 vdd.n167 vdd.n165 0.120292
R282 vdd.n169 vdd.n167 0.120292
R283 vdd.n172 vdd.n169 0.120292
R284 vdd.n175 vdd.n172 0.120292
R285 vdd.n180 vdd.n175 0.120292
R286 vdd.n183 vdd.n180 0.120292
R287 vdd.n185 vdd.n183 0.120292
R288 vdd.n187 vdd.n185 0.120292
R289 vdd.n189 vdd.n187 0.120292
R290 vdd.n140 vdd.n60 0.117348
R291 vdd.n192 vdd.n190 0.0968542
R292 vdd vdd.n192 0.0603958
R293 vdd.n60 vdd.n58 0.0439783
R294 vdd.n190 vdd.n189 0.0239375
R295 vdd.n58 vdd.n56 0.00321739
R296 vss.n90 vss.n89 611.246
R297 vss.n49 vss.n48 292.5
R298 vss.n51 vss.n50 292.5
R299 vss.n53 vss.n52 292.5
R300 vss.n55 vss.n54 292.5
R301 vss.n57 vss.n56 292.5
R302 vss.n59 vss.n58 292.5
R303 vss.n61 vss.n60 292.5
R304 vss.n63 vss.n62 292.5
R305 vss.n65 vss.n64 292.5
R306 vss.n67 vss.n66 292.5
R307 vss.n69 vss.n68 292.5
R308 vss.n71 vss.n70 292.5
R309 vss.n73 vss.n72 292.5
R310 vss.n75 vss.n74 292.5
R311 vss.n77 vss.n76 292.5
R312 vss.n79 vss.n78 292.5
R313 vss.n81 vss.n80 292.5
R314 vss.n83 vss.n82 292.5
R315 vss.n135 vss.n134 292.5
R316 vss.n131 vss.n130 292.5
R317 vss.n44 vss.n43 292.5
R318 vss.n47 vss.n46 292.5
R319 vss.n188 vss.n187 292.5
R320 vss.n186 vss.n185 292.5
R321 vss.n185 vss.n184 292.5
R322 vss.n183 vss.n182 292.5
R323 vss.n182 vss.n181 292.5
R324 vss.n180 vss.n179 292.5
R325 vss.n179 vss.n178 292.5
R326 vss.n177 vss.n176 292.5
R327 vss.n176 vss.n175 292.5
R328 vss.n174 vss.n173 292.5
R329 vss.n173 vss.n172 292.5
R330 vss.n171 vss.n170 292.5
R331 vss.n170 vss.n169 292.5
R332 vss.n168 vss.n167 292.5
R333 vss.n167 vss.n166 292.5
R334 vss.n165 vss.n164 292.5
R335 vss.n164 vss.n163 292.5
R336 vss.n162 vss.n161 292.5
R337 vss.n161 vss.n160 292.5
R338 vss.n159 vss.n158 292.5
R339 vss.n158 vss.n157 292.5
R340 vss.n156 vss.n155 292.5
R341 vss.n155 vss.n154 292.5
R342 vss.n153 vss.n152 292.5
R343 vss.n152 vss.n151 292.5
R344 vss.n150 vss.n149 292.5
R345 vss.n149 vss.n148 292.5
R346 vss.n147 vss.n146 292.5
R347 vss.n146 vss.n145 292.5
R348 vss.n144 vss.n143 292.5
R349 vss.n143 vss.n142 292.5
R350 vss.n141 vss.n140 292.5
R351 vss.n140 vss.n139 292.5
R352 vss.n137 vss.n136 292.5
R353 vss.n138 vss.n137 292.5
R354 vss.n14 vss.t8 193.933
R355 vss.n25 vss.t7 193.933
R356 vss.n5 vss.t11 192.982
R357 vss.n16 vss.t1 192.982
R358 vss.n1 vss.t23 183.082
R359 vss.n130 vss.n129 147.374
R360 vss.n142 vss.t21 140.685
R361 vss.n181 vss.t15 140.685
R362 vss.n133 vss.n132 134.577
R363 vss.n0 vss.t3 123.918
R364 vss.n204 vss.t6 121.956
R365 vss.n27 vss.t5 121.956
R366 vss.n2 vss.t4 121.956
R367 vss.n160 vss.t19 121.279
R368 vss.n163 vss.t18 121.279
R369 vss.n21 vss.n20 114.713
R370 vss.n10 vss.n9 114.713
R371 vss.n139 vss.t13 101.874
R372 vss.n184 vss.t14 101.874
R373 vss.n46 vss.n45 90.6382
R374 vss.n134 vss.n133 90.6381
R375 vss.n49 vss.n47 87.7181
R376 vss.n138 vss.n135 87.7181
R377 vss.n84 vss.n83 82.0711
R378 vss.n189 vss.n188 78.3064
R379 vss.n200 vss.n199 76.0005
R380 vss.n110 vss.n109 63.7358
R381 vss.n148 vss.t12 53.3632
R382 vss.n175 vss.t17 53.3632
R383 vss.n122 vss.n121 52.1476
R384 vss.n123 vss.n122 42.3273
R385 vss.n87 vss.n86 40.452
R386 vss.n88 vss.n87 40.452
R387 vss.n97 vss.n96 35.3848
R388 vss.n98 vss.n97 35.3848
R389 vss.n112 vss.n110 34.7652
R390 vss.n198 vss.t22 34.2973
R391 vss.n154 vss.t20 33.9586
R392 vss.n169 vss.t16 33.9586
R393 vss.n51 vss.n49 25.6005
R394 vss.n53 vss.n51 25.6005
R395 vss.n55 vss.n53 25.6005
R396 vss.n57 vss.n55 25.6005
R397 vss.n59 vss.n57 25.6005
R398 vss.n61 vss.n59 25.6005
R399 vss.n63 vss.n61 25.6005
R400 vss.n65 vss.n63 25.6005
R401 vss.n67 vss.n65 25.6005
R402 vss.n69 vss.n67 25.6005
R403 vss.n71 vss.n69 25.6005
R404 vss.n73 vss.n71 25.6005
R405 vss.n75 vss.n73 25.6005
R406 vss.n77 vss.n75 25.6005
R407 vss.n79 vss.n77 25.6005
R408 vss.n81 vss.n79 25.6005
R409 vss.n83 vss.n81 25.6005
R410 vss.n47 vss.n44 25.6005
R411 vss.n135 vss.n131 25.6005
R412 vss.n141 vss.n138 25.6005
R413 vss.n144 vss.n141 25.6005
R414 vss.n147 vss.n144 25.6005
R415 vss.n150 vss.n147 25.6005
R416 vss.n153 vss.n150 25.6005
R417 vss.n156 vss.n153 25.6005
R418 vss.n159 vss.n156 25.6005
R419 vss.n162 vss.n159 25.6005
R420 vss.n165 vss.n162 25.6005
R421 vss.n168 vss.n165 25.6005
R422 vss.n171 vss.n168 25.6005
R423 vss.n174 vss.n171 25.6005
R424 vss.n177 vss.n174 25.6005
R425 vss.n180 vss.n177 25.6005
R426 vss.n183 vss.n180 25.6005
R427 vss.n186 vss.n183 25.6005
R428 vss.n188 vss.n186 25.6005
R429 vss.n20 vss.t2 24.9236
R430 vss.n20 vss.t0 24.9236
R431 vss.n9 vss.t10 24.9236
R432 vss.n9 vss.t9 24.9236
R433 vss.n100 vss.n98 23.177
R434 vss.n91 vss.n88 11.5887
R435 vss.n190 vss.n189 9.3005
R436 vss.n116 vss.n115 9.3005
R437 vss.n104 vss.n103 9.3005
R438 vss.n92 vss.n91 9.3005
R439 vss.n91 vss.n90 9.3005
R440 vss.n102 vss.n101 9.3005
R441 vss.n101 vss.n100 9.3005
R442 vss.n106 vss.n105 9.3005
R443 vss.n118 vss.n117 9.3005
R444 vss.n114 vss.n113 9.3005
R445 vss.n113 vss.n112 9.3005
R446 vss.n128 vss.n127 9.3005
R447 vss.n126 vss.n125 9.3005
R448 vss.n125 vss.n124 9.3005
R449 vss.n37 vss.n36 9.3005
R450 vss.n42 vss.n41 9.0005
R451 vss.n85 vss.n84 5.64756
R452 vss.n205 vss.n204 4.91351
R453 vss.n95 vss.n94 4.89462
R454 vss.n199 vss.n198 4.85762
R455 vss.n6 vss.n5 4.6505
R456 vss.n15 vss.n14 4.6505
R457 vss.n17 vss.n16 4.6505
R458 vss.n26 vss.n25 4.6505
R459 vss.n203 vss.n202 4.6505
R460 vss.n4 vss.n3 4.6505
R461 vss.n8 vss.n7 4.6505
R462 vss.n11 vss.n10 4.6505
R463 vss.n13 vss.n12 4.6505
R464 vss.n19 vss.n18 4.6505
R465 vss.n22 vss.n21 4.6505
R466 vss.n24 vss.n23 4.6505
R467 vss.n29 vss.n28 4.6505
R468 vss.n31 vss.n30 4.6505
R469 vss.n33 vss.n32 4.6505
R470 vss.n35 vss.n34 4.6505
R471 vss.n191 vss.n190 4.33251
R472 vss.n108 vss.n107 4.14168
R473 vss.n120 vss.n119 3.38874
R474 vss.n202 vss.n200 3.2005
R475 vss.n100 vss.n99 3.16936
R476 vss.n112 vss.n111 3.16936
R477 vss.n125 vss.n120 3.01226
R478 vss.n102 vss.n93 2.26191
R479 vss.n113 vss.n108 2.25932
R480 vss.n93 vss.n92 1.73128
R481 vss.n4 vss.n0 1.64571
R482 vss.n101 vss.n95 1.50638
R483 vss.n2 vss.n1 1.18311
R484 vss.n202 vss.n201 1.14023
R485 vss.n92 vss.n85 0.753441
R486 vss.n124 vss.n123 0.67388
R487 vss.n197 vss.n196 0.614199
R488 vss.n41 vss.n40 0.438856
R489 vss.n3 vss.n2 0.417891
R490 vss.n28 vss.n27 0.409011
R491 vss.n200 vss.n197 0.219678
R492 vss.n114 vss.n106 0.144522
R493 vss.n126 vss.n118 0.144522
R494 vss.n196 vss.n195 0.132007
R495 vss.n6 vss.n4 0.120292
R496 vss.n8 vss.n6 0.120292
R497 vss.n11 vss.n8 0.120292
R498 vss.n13 vss.n11 0.120292
R499 vss.n15 vss.n13 0.120292
R500 vss.n17 vss.n15 0.120292
R501 vss.n19 vss.n17 0.120292
R502 vss.n22 vss.n19 0.120292
R503 vss.n24 vss.n22 0.120292
R504 vss.n26 vss.n24 0.120292
R505 vss.n29 vss.n26 0.120292
R506 vss.n31 vss.n29 0.120292
R507 vss.n33 vss.n31 0.120292
R508 vss.n35 vss.n33 0.120292
R509 vss.n205 vss.n203 0.120292
R510 vss.n203 vss.n194 0.102062
R511 vss.n37 vss.n35 0.10076
R512 vss.n41 vss.n39 0.0881712
R513 vss vss.n205 0.0603958
R514 vss.n192 vss.n191 0.0599291
R515 vss.n191 vss.n42 0.0583581
R516 vss.n106 vss.n104 0.0358261
R517 vss.n118 vss.n116 0.0303913
R518 vss.n190 vss.n128 0.0249565
R519 vss.n128 vss.n126 0.0222391
R520 vss.n38 vss.n37 0.0200312
R521 vss.n194 vss.n193 0.0187292
R522 vss.n116 vss.n114 0.0168043
R523 vss.n104 vss.n102 0.0113696
R524 vss.n193 vss.n192 0.00440625
R525 vss.n42 vss.n38 0.00310417
R526 en.n5 en.t0 212.081
R527 en.n7 en.t1 212.081
R528 en.n2 en.t2 212.081
R529 en.n4 en.t3 212.081
R530 en.n5 en.t4 139.78
R531 en.n7 en.t5 139.78
R532 en.n2 en.t6 139.78
R533 en.n4 en.t7 139.78
R534 en.n9 en.n6 97.5045
R535 en.n9 en.n8 76.0005
R536 en.n11 en.n4 44.2002
R537 en.n6 en.n5 30.6732
R538 en.n8 en.n7 30.6732
R539 en.n3 en.n2 30.6732
R540 en.n4 en.n3 30.6732
R541 en.n11 en.n10 23.8506
R542 en.n10 en.n9 21.5045
R543 en.n13 en.n12 4.3777
R544 en.n15 en.n14 2.24552
R545 en en.n15 0.704975
R546 en.n12 en.n11 0.61644
R547 en.n15 en.n0 0.011716
R548 en.n14 en.n1 0.0083125
R549 en.n14 en.n13 0.00774115
C0 in a_456_865# 0.365f
C1 a_456_1956# en 0.406f
C2 in a_456_1956# 0.464f
C3 vdd out 0.346f
C4 in en 0.0109f
C5 vdd w_0_349# 0.284f
C6 out a_456_865# 0.281f
C7 w_0_349# a_456_865# 0.0493f
C8 a_456_1956# out 0.423f
C9 a_456_1956# w_0_349# 0.183f
C10 out en 0.00102f
C11 vdd a_456_865# 0.712f
C12 w_0_349# en 0.149f
C13 in out 5.32f
C14 vdd a_456_1956# 1.93f
C15 in w_0_349# 0.00429f
C16 a_456_1956# a_456_865# 0.78f
C17 vdd en 0.171f
C18 in vdd 0.706f
C19 en a_456_865# 0.0721f
.ends

