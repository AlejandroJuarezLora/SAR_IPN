magic
tech sky130B
magscale 1 2
timestamp 1697589538
<< nwell >>
rect 263 1577 1777 2145
rect 0 349 2008 670
<< pwell >>
rect 273 753 1767 1291
rect 39 109 773 271
rect 785 109 1223 291
rect 1245 109 1683 291
rect 1695 109 1969 271
<< nmos >>
rect 459 953 519 1153
rect 577 953 637 1153
rect 695 953 755 1153
rect 813 953 873 1153
rect 931 953 991 1153
rect 1049 953 1109 1153
rect 1167 953 1227 1153
rect 1285 953 1345 1153
rect 1403 953 1463 1153
rect 1521 953 1581 1153
<< scnmos >>
rect 117 135 695 245
rect 863 135 893 265
rect 947 135 977 265
rect 1031 135 1061 265
rect 1115 135 1145 265
rect 1323 135 1353 265
rect 1407 135 1437 265
rect 1491 135 1521 265
rect 1575 135 1605 265
rect 1773 135 1891 245
<< pmos >>
rect 459 1725 519 1925
rect 577 1725 637 1925
rect 695 1725 755 1925
rect 813 1725 873 1925
rect 931 1725 991 1925
rect 1049 1725 1109 1925
rect 1167 1725 1227 1925
rect 1285 1725 1345 1925
rect 1403 1725 1463 1925
rect 1521 1725 1581 1925
<< scpmoshvt >>
rect 117 411 695 585
rect 863 385 893 585
rect 947 385 977 585
rect 1031 385 1061 585
rect 1115 385 1145 585
rect 1323 385 1353 585
rect 1407 385 1437 585
rect 1491 385 1521 585
rect 1575 385 1605 585
rect 1773 411 1891 585
<< ndiff >>
rect 401 1138 459 1153
rect 401 1104 413 1138
rect 447 1104 459 1138
rect 401 1070 459 1104
rect 401 1036 413 1070
rect 447 1036 459 1070
rect 401 1002 459 1036
rect 401 968 413 1002
rect 447 968 459 1002
rect 401 953 459 968
rect 519 1138 577 1153
rect 519 1104 531 1138
rect 565 1104 577 1138
rect 519 1070 577 1104
rect 519 1036 531 1070
rect 565 1036 577 1070
rect 519 1002 577 1036
rect 519 968 531 1002
rect 565 968 577 1002
rect 519 953 577 968
rect 637 1138 695 1153
rect 637 1104 649 1138
rect 683 1104 695 1138
rect 637 1070 695 1104
rect 637 1036 649 1070
rect 683 1036 695 1070
rect 637 1002 695 1036
rect 637 968 649 1002
rect 683 968 695 1002
rect 637 953 695 968
rect 755 1138 813 1153
rect 755 1104 767 1138
rect 801 1104 813 1138
rect 755 1070 813 1104
rect 755 1036 767 1070
rect 801 1036 813 1070
rect 755 1002 813 1036
rect 755 968 767 1002
rect 801 968 813 1002
rect 755 953 813 968
rect 873 1138 931 1153
rect 873 1104 885 1138
rect 919 1104 931 1138
rect 873 1070 931 1104
rect 873 1036 885 1070
rect 919 1036 931 1070
rect 873 1002 931 1036
rect 873 968 885 1002
rect 919 968 931 1002
rect 873 953 931 968
rect 991 1138 1049 1153
rect 991 1104 1003 1138
rect 1037 1104 1049 1138
rect 991 1070 1049 1104
rect 991 1036 1003 1070
rect 1037 1036 1049 1070
rect 991 1002 1049 1036
rect 991 968 1003 1002
rect 1037 968 1049 1002
rect 991 953 1049 968
rect 1109 1138 1167 1153
rect 1109 1104 1121 1138
rect 1155 1104 1167 1138
rect 1109 1070 1167 1104
rect 1109 1036 1121 1070
rect 1155 1036 1167 1070
rect 1109 1002 1167 1036
rect 1109 968 1121 1002
rect 1155 968 1167 1002
rect 1109 953 1167 968
rect 1227 1138 1285 1153
rect 1227 1104 1239 1138
rect 1273 1104 1285 1138
rect 1227 1070 1285 1104
rect 1227 1036 1239 1070
rect 1273 1036 1285 1070
rect 1227 1002 1285 1036
rect 1227 968 1239 1002
rect 1273 968 1285 1002
rect 1227 953 1285 968
rect 1345 1138 1403 1153
rect 1345 1104 1357 1138
rect 1391 1104 1403 1138
rect 1345 1070 1403 1104
rect 1345 1036 1357 1070
rect 1391 1036 1403 1070
rect 1345 1002 1403 1036
rect 1345 968 1357 1002
rect 1391 968 1403 1002
rect 1345 953 1403 968
rect 1463 1138 1521 1153
rect 1463 1104 1475 1138
rect 1509 1104 1521 1138
rect 1463 1070 1521 1104
rect 1463 1036 1475 1070
rect 1509 1036 1521 1070
rect 1463 1002 1521 1036
rect 1463 968 1475 1002
rect 1509 968 1521 1002
rect 1463 953 1521 968
rect 1581 1138 1639 1153
rect 1581 1104 1593 1138
rect 1627 1104 1639 1138
rect 1581 1070 1639 1104
rect 1581 1036 1593 1070
rect 1627 1036 1639 1070
rect 1581 1002 1639 1036
rect 1581 968 1593 1002
rect 1627 968 1639 1002
rect 1581 953 1639 968
rect 65 200 117 245
rect 65 166 73 200
rect 107 166 117 200
rect 65 135 117 166
rect 695 200 747 245
rect 695 166 705 200
rect 739 166 747 200
rect 695 135 747 166
rect 811 181 863 265
rect 811 147 819 181
rect 853 147 863 181
rect 811 135 863 147
rect 893 189 947 265
rect 893 155 903 189
rect 937 155 947 189
rect 893 135 947 155
rect 977 181 1031 265
rect 977 147 987 181
rect 1021 147 1031 181
rect 977 135 1031 147
rect 1061 189 1115 265
rect 1061 155 1071 189
rect 1105 155 1115 189
rect 1061 135 1115 155
rect 1145 182 1197 265
rect 1145 148 1155 182
rect 1189 148 1197 182
rect 1145 135 1197 148
rect 1271 181 1323 265
rect 1271 147 1279 181
rect 1313 147 1323 181
rect 1271 135 1323 147
rect 1353 189 1407 265
rect 1353 155 1363 189
rect 1397 155 1407 189
rect 1353 135 1407 155
rect 1437 181 1491 265
rect 1437 147 1447 181
rect 1481 147 1491 181
rect 1437 135 1491 147
rect 1521 189 1575 265
rect 1521 155 1531 189
rect 1565 155 1575 189
rect 1521 135 1575 155
rect 1605 182 1657 265
rect 1605 148 1615 182
rect 1649 148 1657 182
rect 1605 135 1657 148
rect 1721 202 1773 245
rect 1721 168 1729 202
rect 1763 168 1773 202
rect 1721 135 1773 168
rect 1891 202 1943 245
rect 1891 168 1901 202
rect 1935 168 1943 202
rect 1891 135 1943 168
<< pdiff >>
rect 401 1910 459 1925
rect 401 1876 413 1910
rect 447 1876 459 1910
rect 401 1842 459 1876
rect 401 1808 413 1842
rect 447 1808 459 1842
rect 401 1774 459 1808
rect 401 1740 413 1774
rect 447 1740 459 1774
rect 401 1725 459 1740
rect 519 1910 577 1925
rect 519 1876 531 1910
rect 565 1876 577 1910
rect 519 1842 577 1876
rect 519 1808 531 1842
rect 565 1808 577 1842
rect 519 1774 577 1808
rect 519 1740 531 1774
rect 565 1740 577 1774
rect 519 1725 577 1740
rect 637 1910 695 1925
rect 637 1876 649 1910
rect 683 1876 695 1910
rect 637 1842 695 1876
rect 637 1808 649 1842
rect 683 1808 695 1842
rect 637 1774 695 1808
rect 637 1740 649 1774
rect 683 1740 695 1774
rect 637 1725 695 1740
rect 755 1910 813 1925
rect 755 1876 767 1910
rect 801 1876 813 1910
rect 755 1842 813 1876
rect 755 1808 767 1842
rect 801 1808 813 1842
rect 755 1774 813 1808
rect 755 1740 767 1774
rect 801 1740 813 1774
rect 755 1725 813 1740
rect 873 1910 931 1925
rect 873 1876 885 1910
rect 919 1876 931 1910
rect 873 1842 931 1876
rect 873 1808 885 1842
rect 919 1808 931 1842
rect 873 1774 931 1808
rect 873 1740 885 1774
rect 919 1740 931 1774
rect 873 1725 931 1740
rect 991 1910 1049 1925
rect 991 1876 1003 1910
rect 1037 1876 1049 1910
rect 991 1842 1049 1876
rect 991 1808 1003 1842
rect 1037 1808 1049 1842
rect 991 1774 1049 1808
rect 991 1740 1003 1774
rect 1037 1740 1049 1774
rect 991 1725 1049 1740
rect 1109 1910 1167 1925
rect 1109 1876 1121 1910
rect 1155 1876 1167 1910
rect 1109 1842 1167 1876
rect 1109 1808 1121 1842
rect 1155 1808 1167 1842
rect 1109 1774 1167 1808
rect 1109 1740 1121 1774
rect 1155 1740 1167 1774
rect 1109 1725 1167 1740
rect 1227 1910 1285 1925
rect 1227 1876 1239 1910
rect 1273 1876 1285 1910
rect 1227 1842 1285 1876
rect 1227 1808 1239 1842
rect 1273 1808 1285 1842
rect 1227 1774 1285 1808
rect 1227 1740 1239 1774
rect 1273 1740 1285 1774
rect 1227 1725 1285 1740
rect 1345 1910 1403 1925
rect 1345 1876 1357 1910
rect 1391 1876 1403 1910
rect 1345 1842 1403 1876
rect 1345 1808 1357 1842
rect 1391 1808 1403 1842
rect 1345 1774 1403 1808
rect 1345 1740 1357 1774
rect 1391 1740 1403 1774
rect 1345 1725 1403 1740
rect 1463 1910 1521 1925
rect 1463 1876 1475 1910
rect 1509 1876 1521 1910
rect 1463 1842 1521 1876
rect 1463 1808 1475 1842
rect 1509 1808 1521 1842
rect 1463 1774 1521 1808
rect 1463 1740 1475 1774
rect 1509 1740 1521 1774
rect 1463 1725 1521 1740
rect 1581 1910 1639 1925
rect 1581 1876 1593 1910
rect 1627 1876 1639 1910
rect 1581 1842 1639 1876
rect 1581 1808 1593 1842
rect 1627 1808 1639 1842
rect 1581 1774 1639 1808
rect 1581 1740 1593 1774
rect 1627 1740 1639 1774
rect 1581 1725 1639 1740
rect 65 573 117 585
rect 65 539 73 573
rect 107 539 117 573
rect 65 471 117 539
rect 65 437 73 471
rect 107 437 117 471
rect 65 411 117 437
rect 695 573 747 585
rect 695 539 705 573
rect 739 539 747 573
rect 695 471 747 539
rect 695 437 705 471
rect 739 437 747 471
rect 695 411 747 437
rect 811 573 863 585
rect 811 539 819 573
rect 853 539 863 573
rect 811 505 863 539
rect 811 471 819 505
rect 853 471 863 505
rect 811 437 863 471
rect 811 403 819 437
rect 853 403 863 437
rect 811 385 863 403
rect 893 573 947 585
rect 893 539 903 573
rect 937 539 947 573
rect 893 505 947 539
rect 893 471 903 505
rect 937 471 947 505
rect 893 437 947 471
rect 893 403 903 437
rect 937 403 947 437
rect 893 385 947 403
rect 977 573 1031 585
rect 977 539 987 573
rect 1021 539 1031 573
rect 977 505 1031 539
rect 977 471 987 505
rect 1021 471 1031 505
rect 977 385 1031 471
rect 1061 573 1115 585
rect 1061 539 1071 573
rect 1105 539 1115 573
rect 1061 505 1115 539
rect 1061 471 1071 505
rect 1105 471 1115 505
rect 1061 437 1115 471
rect 1061 403 1071 437
rect 1105 403 1115 437
rect 1061 385 1115 403
rect 1145 573 1197 585
rect 1145 539 1155 573
rect 1189 539 1197 573
rect 1145 385 1197 539
rect 1271 573 1323 585
rect 1271 539 1279 573
rect 1313 539 1323 573
rect 1271 505 1323 539
rect 1271 471 1279 505
rect 1313 471 1323 505
rect 1271 437 1323 471
rect 1271 403 1279 437
rect 1313 403 1323 437
rect 1271 385 1323 403
rect 1353 573 1407 585
rect 1353 539 1363 573
rect 1397 539 1407 573
rect 1353 505 1407 539
rect 1353 471 1363 505
rect 1397 471 1407 505
rect 1353 437 1407 471
rect 1353 403 1363 437
rect 1397 403 1407 437
rect 1353 385 1407 403
rect 1437 573 1491 585
rect 1437 539 1447 573
rect 1481 539 1491 573
rect 1437 505 1491 539
rect 1437 471 1447 505
rect 1481 471 1491 505
rect 1437 385 1491 471
rect 1521 573 1575 585
rect 1521 539 1531 573
rect 1565 539 1575 573
rect 1521 505 1575 539
rect 1521 471 1531 505
rect 1565 471 1575 505
rect 1521 437 1575 471
rect 1521 403 1531 437
rect 1565 403 1575 437
rect 1521 385 1575 403
rect 1605 573 1657 585
rect 1605 539 1615 573
rect 1649 539 1657 573
rect 1605 385 1657 539
rect 1721 573 1773 585
rect 1721 539 1729 573
rect 1763 539 1773 573
rect 1721 478 1773 539
rect 1721 444 1729 478
rect 1763 444 1773 478
rect 1721 411 1773 444
rect 1891 573 1943 585
rect 1891 539 1901 573
rect 1935 539 1943 573
rect 1891 478 1943 539
rect 1891 444 1901 478
rect 1935 444 1943 478
rect 1891 411 1943 444
<< ndiffc >>
rect 413 1104 447 1138
rect 413 1036 447 1070
rect 413 968 447 1002
rect 531 1104 565 1138
rect 531 1036 565 1070
rect 531 968 565 1002
rect 649 1104 683 1138
rect 649 1036 683 1070
rect 649 968 683 1002
rect 767 1104 801 1138
rect 767 1036 801 1070
rect 767 968 801 1002
rect 885 1104 919 1138
rect 885 1036 919 1070
rect 885 968 919 1002
rect 1003 1104 1037 1138
rect 1003 1036 1037 1070
rect 1003 968 1037 1002
rect 1121 1104 1155 1138
rect 1121 1036 1155 1070
rect 1121 968 1155 1002
rect 1239 1104 1273 1138
rect 1239 1036 1273 1070
rect 1239 968 1273 1002
rect 1357 1104 1391 1138
rect 1357 1036 1391 1070
rect 1357 968 1391 1002
rect 1475 1104 1509 1138
rect 1475 1036 1509 1070
rect 1475 968 1509 1002
rect 1593 1104 1627 1138
rect 1593 1036 1627 1070
rect 1593 968 1627 1002
rect 73 166 107 200
rect 705 166 739 200
rect 819 147 853 181
rect 903 155 937 189
rect 987 147 1021 181
rect 1071 155 1105 189
rect 1155 148 1189 182
rect 1279 147 1313 181
rect 1363 155 1397 189
rect 1447 147 1481 181
rect 1531 155 1565 189
rect 1615 148 1649 182
rect 1729 168 1763 202
rect 1901 168 1935 202
<< pdiffc >>
rect 413 1876 447 1910
rect 413 1808 447 1842
rect 413 1740 447 1774
rect 531 1876 565 1910
rect 531 1808 565 1842
rect 531 1740 565 1774
rect 649 1876 683 1910
rect 649 1808 683 1842
rect 649 1740 683 1774
rect 767 1876 801 1910
rect 767 1808 801 1842
rect 767 1740 801 1774
rect 885 1876 919 1910
rect 885 1808 919 1842
rect 885 1740 919 1774
rect 1003 1876 1037 1910
rect 1003 1808 1037 1842
rect 1003 1740 1037 1774
rect 1121 1876 1155 1910
rect 1121 1808 1155 1842
rect 1121 1740 1155 1774
rect 1239 1876 1273 1910
rect 1239 1808 1273 1842
rect 1239 1740 1273 1774
rect 1357 1876 1391 1910
rect 1357 1808 1391 1842
rect 1357 1740 1391 1774
rect 1475 1876 1509 1910
rect 1475 1808 1509 1842
rect 1475 1740 1509 1774
rect 1593 1876 1627 1910
rect 1593 1808 1627 1842
rect 1593 1740 1627 1774
rect 73 539 107 573
rect 73 437 107 471
rect 705 539 739 573
rect 705 437 739 471
rect 819 539 853 573
rect 819 471 853 505
rect 819 403 853 437
rect 903 539 937 573
rect 903 471 937 505
rect 903 403 937 437
rect 987 539 1021 573
rect 987 471 1021 505
rect 1071 539 1105 573
rect 1071 471 1105 505
rect 1071 403 1105 437
rect 1155 539 1189 573
rect 1279 539 1313 573
rect 1279 471 1313 505
rect 1279 403 1313 437
rect 1363 539 1397 573
rect 1363 471 1397 505
rect 1363 403 1397 437
rect 1447 539 1481 573
rect 1447 471 1481 505
rect 1531 539 1565 573
rect 1531 471 1565 505
rect 1531 403 1565 437
rect 1615 539 1649 573
rect 1729 539 1763 573
rect 1729 444 1763 478
rect 1901 539 1935 573
rect 1901 444 1935 478
<< psubdiff >>
rect 299 1231 425 1265
rect 459 1231 493 1265
rect 527 1231 561 1265
rect 595 1231 629 1265
rect 663 1231 697 1265
rect 731 1231 765 1265
rect 799 1231 833 1265
rect 867 1231 901 1265
rect 935 1231 969 1265
rect 1003 1231 1037 1265
rect 1071 1231 1105 1265
rect 1139 1231 1173 1265
rect 1207 1231 1241 1265
rect 1275 1231 1309 1265
rect 1343 1231 1377 1265
rect 1411 1231 1445 1265
rect 1479 1231 1513 1265
rect 1547 1231 1581 1265
rect 1615 1231 1741 1265
rect 299 1141 333 1231
rect 299 1073 333 1107
rect 299 1005 333 1039
rect 299 937 333 971
rect 1707 1141 1741 1231
rect 1707 1073 1741 1107
rect 1707 1005 1741 1039
rect 1707 937 1741 971
rect 299 813 333 903
rect 1707 813 1741 903
rect 299 779 425 813
rect 459 779 493 813
rect 527 779 561 813
rect 595 779 629 813
rect 663 779 697 813
rect 731 779 765 813
rect 799 779 833 813
rect 867 779 901 813
rect 935 779 969 813
rect 1003 779 1037 813
rect 1071 779 1105 813
rect 1139 779 1173 813
rect 1207 779 1241 813
rect 1275 779 1309 813
rect 1343 779 1377 813
rect 1411 779 1445 813
rect 1479 779 1513 813
rect 1547 779 1581 813
rect 1615 779 1741 813
<< nsubdiff >>
rect 299 2075 425 2109
rect 459 2075 493 2109
rect 527 2075 561 2109
rect 595 2075 629 2109
rect 663 2075 697 2109
rect 731 2075 765 2109
rect 799 2075 833 2109
rect 867 2075 901 2109
rect 935 2075 969 2109
rect 1003 2075 1037 2109
rect 1071 2075 1105 2109
rect 1139 2075 1173 2109
rect 1207 2075 1241 2109
rect 1275 2075 1309 2109
rect 1343 2075 1377 2109
rect 1411 2075 1445 2109
rect 1479 2075 1513 2109
rect 1547 2075 1581 2109
rect 1615 2075 1741 2109
rect 299 1980 333 2075
rect 1707 1980 1741 2075
rect 299 1912 333 1946
rect 299 1844 333 1878
rect 299 1776 333 1810
rect 299 1647 333 1742
rect 1707 1912 1741 1946
rect 1707 1844 1741 1878
rect 1707 1776 1741 1810
rect 1707 1647 1741 1742
rect 299 1613 425 1647
rect 459 1613 493 1647
rect 527 1613 561 1647
rect 595 1613 629 1647
rect 663 1613 697 1647
rect 731 1613 765 1647
rect 799 1613 833 1647
rect 867 1613 901 1647
rect 935 1613 969 1647
rect 1003 1613 1037 1647
rect 1071 1613 1105 1647
rect 1139 1613 1173 1647
rect 1207 1613 1241 1647
rect 1275 1613 1309 1647
rect 1343 1613 1377 1647
rect 1411 1613 1445 1647
rect 1479 1613 1513 1647
rect 1547 1613 1581 1647
rect 1615 1613 1741 1647
<< psubdiffcont >>
rect 425 1231 459 1265
rect 493 1231 527 1265
rect 561 1231 595 1265
rect 629 1231 663 1265
rect 697 1231 731 1265
rect 765 1231 799 1265
rect 833 1231 867 1265
rect 901 1231 935 1265
rect 969 1231 1003 1265
rect 1037 1231 1071 1265
rect 1105 1231 1139 1265
rect 1173 1231 1207 1265
rect 1241 1231 1275 1265
rect 1309 1231 1343 1265
rect 1377 1231 1411 1265
rect 1445 1231 1479 1265
rect 1513 1231 1547 1265
rect 1581 1231 1615 1265
rect 299 1107 333 1141
rect 299 1039 333 1073
rect 299 971 333 1005
rect 1707 1107 1741 1141
rect 1707 1039 1741 1073
rect 1707 971 1741 1005
rect 299 903 333 937
rect 1707 903 1741 937
rect 425 779 459 813
rect 493 779 527 813
rect 561 779 595 813
rect 629 779 663 813
rect 697 779 731 813
rect 765 779 799 813
rect 833 779 867 813
rect 901 779 935 813
rect 969 779 1003 813
rect 1037 779 1071 813
rect 1105 779 1139 813
rect 1173 779 1207 813
rect 1241 779 1275 813
rect 1309 779 1343 813
rect 1377 779 1411 813
rect 1445 779 1479 813
rect 1513 779 1547 813
rect 1581 779 1615 813
<< nsubdiffcont >>
rect 425 2075 459 2109
rect 493 2075 527 2109
rect 561 2075 595 2109
rect 629 2075 663 2109
rect 697 2075 731 2109
rect 765 2075 799 2109
rect 833 2075 867 2109
rect 901 2075 935 2109
rect 969 2075 1003 2109
rect 1037 2075 1071 2109
rect 1105 2075 1139 2109
rect 1173 2075 1207 2109
rect 1241 2075 1275 2109
rect 1309 2075 1343 2109
rect 1377 2075 1411 2109
rect 1445 2075 1479 2109
rect 1513 2075 1547 2109
rect 1581 2075 1615 2109
rect 299 1946 333 1980
rect 1707 1946 1741 1980
rect 299 1878 333 1912
rect 299 1810 333 1844
rect 299 1742 333 1776
rect 1707 1878 1741 1912
rect 1707 1810 1741 1844
rect 1707 1742 1741 1776
rect 425 1613 459 1647
rect 493 1613 527 1647
rect 561 1613 595 1647
rect 629 1613 663 1647
rect 697 1613 731 1647
rect 765 1613 799 1647
rect 833 1613 867 1647
rect 901 1613 935 1647
rect 969 1613 1003 1647
rect 1037 1613 1071 1647
rect 1105 1613 1139 1647
rect 1173 1613 1207 1647
rect 1241 1613 1275 1647
rect 1309 1613 1343 1647
rect 1377 1613 1411 1647
rect 1445 1613 1479 1647
rect 1513 1613 1547 1647
rect 1581 1613 1615 1647
<< poly >>
rect 456 2006 522 2022
rect 456 1972 472 2006
rect 506 1972 522 2006
rect 456 1956 522 1972
rect 574 2006 640 2022
rect 574 1972 590 2006
rect 624 1972 640 2006
rect 574 1956 640 1972
rect 692 2006 758 2022
rect 692 1972 708 2006
rect 742 1972 758 2006
rect 692 1956 758 1972
rect 810 2006 876 2022
rect 810 1972 826 2006
rect 860 1972 876 2006
rect 810 1956 876 1972
rect 928 2006 994 2022
rect 928 1972 944 2006
rect 978 1972 994 2006
rect 928 1956 994 1972
rect 1046 2006 1112 2022
rect 1046 1972 1062 2006
rect 1096 1972 1112 2006
rect 1046 1956 1112 1972
rect 1164 2006 1230 2022
rect 1164 1972 1180 2006
rect 1214 1972 1230 2006
rect 1164 1956 1230 1972
rect 1282 2006 1348 2022
rect 1282 1972 1298 2006
rect 1332 1972 1348 2006
rect 1282 1956 1348 1972
rect 1400 2006 1466 2022
rect 1400 1972 1416 2006
rect 1450 1972 1466 2006
rect 1400 1956 1466 1972
rect 1518 2006 1584 2022
rect 1518 1972 1534 2006
rect 1568 1972 1584 2006
rect 1518 1956 1584 1972
rect 459 1925 519 1956
rect 577 1925 637 1956
rect 695 1925 755 1956
rect 813 1925 873 1956
rect 931 1925 991 1956
rect 1049 1925 1109 1956
rect 1167 1925 1227 1956
rect 1285 1925 1345 1956
rect 1403 1925 1463 1956
rect 1521 1925 1581 1956
rect 459 1699 519 1725
rect 577 1699 637 1725
rect 695 1699 755 1725
rect 813 1699 873 1725
rect 931 1699 991 1725
rect 1049 1699 1109 1725
rect 1167 1699 1227 1725
rect 1285 1699 1345 1725
rect 1403 1699 1463 1725
rect 1521 1699 1581 1725
rect 459 1153 519 1179
rect 577 1153 637 1179
rect 695 1153 755 1179
rect 813 1153 873 1179
rect 931 1153 991 1179
rect 1049 1153 1109 1179
rect 1167 1153 1227 1179
rect 1285 1153 1345 1179
rect 1403 1153 1463 1179
rect 1521 1153 1581 1179
rect 459 931 519 953
rect 577 931 637 953
rect 695 931 755 953
rect 813 931 873 953
rect 931 931 991 953
rect 1049 931 1109 953
rect 1167 931 1227 953
rect 1285 931 1345 953
rect 1403 931 1463 953
rect 1521 931 1581 953
rect 456 915 522 931
rect 456 881 472 915
rect 506 881 522 915
rect 456 865 522 881
rect 574 915 640 931
rect 574 881 590 915
rect 624 881 640 915
rect 574 865 640 881
rect 692 915 758 931
rect 692 881 708 915
rect 742 881 758 915
rect 692 865 758 881
rect 810 915 876 931
rect 810 881 826 915
rect 860 881 876 915
rect 810 865 876 881
rect 928 915 994 931
rect 928 881 944 915
rect 978 881 994 915
rect 928 865 994 881
rect 1046 915 1112 931
rect 1046 881 1062 915
rect 1096 881 1112 915
rect 1046 865 1112 881
rect 1164 915 1230 931
rect 1164 881 1180 915
rect 1214 881 1230 915
rect 1164 865 1230 881
rect 1282 915 1348 931
rect 1282 881 1298 915
rect 1332 881 1348 915
rect 1282 865 1348 881
rect 1400 915 1466 931
rect 1400 881 1416 915
rect 1450 881 1466 915
rect 1400 865 1466 881
rect 1518 915 1584 931
rect 1518 881 1534 915
rect 1568 881 1584 915
rect 1518 865 1584 881
rect 117 585 695 611
rect 863 585 893 611
rect 947 585 977 611
rect 1031 585 1061 611
rect 1115 585 1145 611
rect 1323 585 1353 611
rect 1407 585 1437 611
rect 1491 585 1521 611
rect 1575 585 1605 611
rect 1773 585 1891 611
rect 117 385 695 411
rect 117 363 381 385
rect 117 329 133 363
rect 167 329 232 363
rect 266 329 331 363
rect 365 329 381 363
rect 863 353 893 385
rect 947 353 977 385
rect 1031 353 1061 385
rect 1115 353 1145 385
rect 1323 353 1353 385
rect 1407 353 1437 385
rect 1491 353 1521 385
rect 1575 353 1605 385
rect 1773 381 1891 411
rect 1773 379 1811 381
rect 117 313 381 329
rect 423 327 695 343
rect 423 293 439 327
rect 473 293 542 327
rect 576 293 645 327
rect 679 293 695 327
rect 423 271 695 293
rect 795 337 1145 353
rect 795 303 811 337
rect 845 303 903 337
rect 937 303 987 337
rect 1021 303 1071 337
rect 1105 303 1145 337
rect 795 287 1145 303
rect 1255 337 1605 353
rect 1255 303 1271 337
rect 1305 303 1363 337
rect 1397 303 1447 337
rect 1481 303 1531 337
rect 1565 303 1605 337
rect 1745 363 1811 379
rect 1745 329 1761 363
rect 1795 329 1811 363
rect 1745 313 1811 329
rect 1853 323 1919 339
rect 1255 287 1605 303
rect 117 245 695 271
rect 863 265 893 287
rect 947 265 977 287
rect 1031 265 1061 287
rect 1115 265 1145 287
rect 1323 265 1353 287
rect 1407 265 1437 287
rect 1491 265 1521 287
rect 1575 265 1605 287
rect 1853 289 1869 323
rect 1903 289 1919 323
rect 1853 273 1919 289
rect 1853 271 1891 273
rect 1773 245 1891 271
rect 117 109 695 135
rect 863 109 893 135
rect 947 109 977 135
rect 1031 109 1061 135
rect 1115 109 1145 135
rect 1323 109 1353 135
rect 1407 109 1437 135
rect 1491 109 1521 135
rect 1575 109 1605 135
rect 1773 109 1891 135
<< polycont >>
rect 472 1972 506 2006
rect 590 1972 624 2006
rect 708 1972 742 2006
rect 826 1972 860 2006
rect 944 1972 978 2006
rect 1062 1972 1096 2006
rect 1180 1972 1214 2006
rect 1298 1972 1332 2006
rect 1416 1972 1450 2006
rect 1534 1972 1568 2006
rect 472 881 506 915
rect 590 881 624 915
rect 708 881 742 915
rect 826 881 860 915
rect 944 881 978 915
rect 1062 881 1096 915
rect 1180 881 1214 915
rect 1298 881 1332 915
rect 1416 881 1450 915
rect 1534 881 1568 915
rect 133 329 167 363
rect 232 329 266 363
rect 331 329 365 363
rect 439 293 473 327
rect 542 293 576 327
rect 645 293 679 327
rect 811 303 845 337
rect 903 303 937 337
rect 987 303 1021 337
rect 1071 303 1105 337
rect 1271 303 1305 337
rect 1363 303 1397 337
rect 1447 303 1481 337
rect 1531 303 1565 337
rect 1761 329 1795 363
rect 1869 289 1903 323
<< locali >>
rect 299 2075 425 2109
rect 459 2075 493 2109
rect 527 2075 561 2109
rect 595 2075 629 2109
rect 663 2075 697 2109
rect 731 2075 765 2109
rect 799 2075 833 2109
rect 867 2075 901 2109
rect 935 2075 969 2109
rect 1003 2075 1037 2109
rect 1071 2075 1105 2109
rect 1139 2075 1173 2109
rect 1207 2075 1241 2109
rect 1275 2075 1309 2109
rect 1343 2075 1377 2109
rect 1411 2075 1445 2109
rect 1479 2075 1513 2109
rect 1547 2075 1581 2109
rect 1615 2075 1741 2109
rect 299 1982 333 2075
rect 456 1972 472 2006
rect 506 1972 522 2006
rect 574 1972 590 2006
rect 624 1972 640 2006
rect 692 1972 708 2006
rect 742 1972 758 2006
rect 810 1972 826 2006
rect 860 1972 876 2006
rect 928 1972 944 2006
rect 978 1972 994 2006
rect 1046 1972 1062 2006
rect 1096 1972 1112 2006
rect 1164 1972 1180 2006
rect 1214 1972 1230 2006
rect 1282 1972 1298 2006
rect 1332 1972 1348 2006
rect 1400 1972 1416 2006
rect 1450 1972 1466 2006
rect 1518 1972 1534 2006
rect 1568 1972 1584 2006
rect 1707 1980 1741 2075
rect 299 1912 333 1946
rect 299 1844 333 1876
rect 299 1776 333 1804
rect 299 1647 333 1732
rect 413 1910 447 1929
rect 413 1842 447 1844
rect 413 1806 447 1808
rect 413 1721 447 1740
rect 531 1910 565 1929
rect 531 1842 565 1844
rect 531 1806 565 1808
rect 531 1721 565 1740
rect 649 1910 683 1929
rect 649 1842 683 1844
rect 649 1806 683 1808
rect 649 1721 683 1740
rect 767 1910 801 1929
rect 767 1842 801 1844
rect 767 1806 801 1808
rect 767 1721 801 1740
rect 885 1910 919 1929
rect 885 1842 919 1844
rect 885 1806 919 1808
rect 885 1721 919 1740
rect 1003 1910 1037 1929
rect 1003 1842 1037 1844
rect 1003 1806 1037 1808
rect 1003 1721 1037 1740
rect 1121 1910 1155 1929
rect 1121 1842 1155 1844
rect 1121 1806 1155 1808
rect 1121 1721 1155 1740
rect 1239 1910 1273 1929
rect 1239 1842 1273 1844
rect 1239 1806 1273 1808
rect 1239 1721 1273 1740
rect 1357 1910 1391 1929
rect 1357 1842 1391 1844
rect 1357 1806 1391 1808
rect 1357 1721 1391 1740
rect 1475 1910 1509 1929
rect 1475 1842 1509 1844
rect 1475 1806 1509 1808
rect 1475 1721 1509 1740
rect 1593 1910 1627 1929
rect 1593 1842 1627 1844
rect 1593 1806 1627 1808
rect 1593 1721 1627 1740
rect 1707 1912 1741 1946
rect 1707 1844 1741 1878
rect 1707 1776 1741 1810
rect 1707 1647 1741 1742
rect 299 1613 425 1647
rect 459 1613 493 1647
rect 527 1613 561 1647
rect 595 1613 629 1647
rect 663 1613 697 1647
rect 731 1613 765 1647
rect 799 1613 833 1647
rect 867 1613 901 1647
rect 935 1613 969 1647
rect 1003 1613 1037 1647
rect 1071 1613 1105 1647
rect 1139 1613 1173 1647
rect 1207 1613 1241 1647
rect 1275 1613 1309 1647
rect 1343 1613 1377 1647
rect 1411 1613 1445 1647
rect 1479 1613 1513 1647
rect 1547 1613 1581 1647
rect 1615 1613 1741 1647
rect 299 1231 425 1265
rect 459 1231 493 1265
rect 527 1231 561 1265
rect 595 1231 629 1265
rect 663 1231 697 1265
rect 731 1231 765 1265
rect 799 1231 833 1265
rect 867 1231 901 1265
rect 935 1231 969 1265
rect 1003 1231 1037 1265
rect 1071 1231 1105 1265
rect 1139 1231 1173 1265
rect 1207 1231 1241 1265
rect 1275 1231 1309 1265
rect 1343 1231 1377 1265
rect 1411 1231 1445 1265
rect 1479 1231 1513 1265
rect 1547 1231 1581 1265
rect 1615 1231 1741 1265
rect 299 1141 333 1231
rect 299 1073 333 1103
rect 299 1005 333 1031
rect 299 937 333 959
rect 413 1138 447 1157
rect 413 1070 447 1072
rect 413 1034 447 1036
rect 413 949 447 968
rect 531 1138 565 1157
rect 531 1070 565 1072
rect 531 1034 565 1036
rect 531 949 565 968
rect 649 1138 683 1157
rect 649 1070 683 1072
rect 649 1034 683 1036
rect 649 949 683 968
rect 767 1138 801 1157
rect 767 1070 801 1072
rect 767 1034 801 1036
rect 767 949 801 968
rect 885 1138 919 1157
rect 885 1070 919 1072
rect 885 1034 919 1036
rect 885 949 919 968
rect 1003 1138 1037 1157
rect 1003 1070 1037 1072
rect 1003 1034 1037 1036
rect 1003 949 1037 968
rect 1121 1138 1155 1157
rect 1121 1070 1155 1072
rect 1121 1034 1155 1036
rect 1121 949 1155 968
rect 1239 1138 1273 1157
rect 1239 1070 1273 1072
rect 1239 1034 1273 1036
rect 1239 949 1273 968
rect 1357 1138 1391 1157
rect 1357 1070 1391 1072
rect 1357 1034 1391 1036
rect 1357 949 1391 968
rect 1475 1138 1509 1157
rect 1475 1070 1509 1072
rect 1475 1034 1509 1036
rect 1475 949 1509 968
rect 1593 1138 1627 1157
rect 1593 1070 1627 1072
rect 1593 1034 1627 1036
rect 1593 949 1627 968
rect 1707 1141 1741 1231
rect 1707 1073 1741 1107
rect 1707 1005 1741 1039
rect 1707 937 1741 971
rect 299 813 333 887
rect 456 881 472 915
rect 506 881 522 915
rect 574 881 590 915
rect 624 881 640 915
rect 692 881 708 915
rect 742 881 758 915
rect 810 881 826 915
rect 860 881 876 915
rect 928 881 944 915
rect 978 881 994 915
rect 1046 881 1062 915
rect 1096 881 1112 915
rect 1164 881 1180 915
rect 1214 881 1230 915
rect 1282 881 1298 915
rect 1332 881 1348 915
rect 1400 881 1416 915
rect 1450 881 1466 915
rect 1518 881 1534 915
rect 1568 881 1584 915
rect 1707 813 1741 903
rect 299 779 425 813
rect 459 779 493 813
rect 527 779 561 813
rect 595 779 629 813
rect 663 779 697 813
rect 731 779 765 813
rect 799 779 833 813
rect 867 779 901 813
rect 935 779 969 813
rect 1003 779 1037 813
rect 1071 779 1105 813
rect 1139 779 1173 813
rect 1207 779 1241 813
rect 1275 779 1309 813
rect 1343 779 1377 813
rect 1411 779 1445 813
rect 1479 779 1513 813
rect 1547 779 1581 813
rect 1615 779 1741 813
rect 38 615 67 649
rect 101 615 159 649
rect 193 615 251 649
rect 285 615 343 649
rect 377 615 435 649
rect 469 615 527 649
rect 561 615 619 649
rect 653 615 711 649
rect 745 615 803 649
rect 837 615 895 649
rect 929 615 987 649
rect 1021 615 1079 649
rect 1113 615 1171 649
rect 1205 615 1263 649
rect 1297 615 1355 649
rect 1389 615 1447 649
rect 1481 615 1539 649
rect 1573 615 1631 649
rect 1665 615 1723 649
rect 1757 615 1815 649
rect 1849 615 1907 649
rect 1941 615 1970 649
rect 55 573 757 615
rect 55 539 73 573
rect 107 539 705 573
rect 739 539 757 573
rect 55 471 757 539
rect 55 437 73 471
rect 107 437 705 471
rect 739 437 757 471
rect 55 397 757 437
rect 55 329 133 363
rect 167 329 232 363
rect 266 329 331 363
rect 365 329 385 363
rect 55 259 385 329
rect 419 327 757 397
rect 800 573 853 615
rect 800 539 819 573
rect 800 505 853 539
rect 800 471 819 505
rect 800 437 853 471
rect 800 403 819 437
rect 800 387 853 403
rect 887 573 953 581
rect 887 539 903 573
rect 937 539 953 573
rect 887 505 953 539
rect 887 471 903 505
rect 937 471 953 505
rect 887 437 953 471
rect 987 573 1021 615
rect 987 505 1021 539
rect 987 455 1021 471
rect 1055 573 1121 581
rect 1055 539 1071 573
rect 1105 539 1121 573
rect 1055 505 1121 539
rect 1155 573 1197 615
rect 1189 539 1197 573
rect 1155 523 1197 539
rect 1260 573 1313 615
rect 1260 539 1279 573
rect 1055 471 1071 505
rect 1105 471 1121 505
rect 887 403 903 437
rect 937 421 953 437
rect 1055 437 1121 471
rect 1055 421 1071 437
rect 937 403 1071 421
rect 1105 425 1121 437
rect 1260 505 1313 539
rect 1260 471 1279 505
rect 1260 437 1313 471
rect 1105 411 1208 425
rect 1105 403 1171 411
rect 887 387 1171 403
rect 1155 377 1171 387
rect 1205 377 1208 411
rect 1260 403 1279 437
rect 1260 387 1313 403
rect 1347 573 1413 581
rect 1347 539 1363 573
rect 1397 539 1413 573
rect 1347 505 1413 539
rect 1347 471 1363 505
rect 1397 471 1413 505
rect 1347 437 1413 471
rect 1447 573 1481 615
rect 1447 505 1481 539
rect 1447 455 1481 471
rect 1515 573 1581 581
rect 1515 539 1531 573
rect 1565 539 1581 573
rect 1515 505 1581 539
rect 1615 573 1657 615
rect 1649 539 1657 573
rect 1615 523 1657 539
rect 1711 573 1953 615
rect 1711 539 1729 573
rect 1763 539 1901 573
rect 1935 539 1953 573
rect 1515 471 1531 505
rect 1565 471 1581 505
rect 1347 403 1363 437
rect 1397 421 1413 437
rect 1515 437 1581 471
rect 1515 421 1531 437
rect 1397 403 1531 421
rect 1565 425 1581 437
rect 1711 478 1953 539
rect 1711 444 1729 478
rect 1763 444 1901 478
rect 1935 444 1953 478
rect 1565 411 1668 425
rect 1565 403 1631 411
rect 1347 387 1631 403
rect 419 293 439 327
rect 473 293 542 327
rect 576 293 645 327
rect 679 293 757 327
rect 795 343 1121 353
rect 795 309 803 343
rect 837 337 1121 343
rect 795 303 811 309
rect 845 303 903 337
rect 937 303 987 337
rect 1021 303 1071 337
rect 1105 303 1121 337
rect 1155 269 1208 377
rect 1615 377 1631 387
rect 1665 377 1668 411
rect 1711 397 1953 444
rect 1255 345 1581 353
rect 1255 337 1288 345
rect 1322 337 1581 345
rect 1255 303 1271 337
rect 1322 311 1363 337
rect 1305 303 1363 311
rect 1397 303 1447 337
rect 1481 303 1531 337
rect 1565 303 1581 337
rect 1615 269 1668 377
rect 55 200 757 259
rect 55 166 73 200
rect 107 166 705 200
rect 739 166 757 200
rect 887 233 1208 269
rect 1347 233 1668 269
rect 1711 329 1761 363
rect 1795 329 1815 363
rect 1711 255 1815 329
rect 1849 323 1953 397
rect 1849 289 1869 323
rect 1903 289 1953 323
rect 55 105 757 166
rect 800 181 853 197
rect 800 147 819 181
rect 800 105 853 147
rect 887 189 953 233
rect 887 155 903 189
rect 937 155 953 189
rect 887 139 953 155
rect 987 181 1021 197
rect 987 105 1021 147
rect 1055 189 1121 233
rect 1055 155 1071 189
rect 1105 155 1121 189
rect 1055 139 1121 155
rect 1155 182 1205 198
rect 1189 148 1205 182
rect 1155 105 1205 148
rect 1260 181 1313 197
rect 1260 147 1279 181
rect 1260 105 1313 147
rect 1347 189 1413 233
rect 1347 155 1363 189
rect 1397 155 1413 189
rect 1347 139 1413 155
rect 1447 181 1481 197
rect 1447 105 1481 147
rect 1515 189 1581 233
rect 1711 202 1953 255
rect 1515 155 1531 189
rect 1565 155 1581 189
rect 1515 139 1581 155
rect 1615 182 1665 198
rect 1649 148 1665 182
rect 1615 105 1665 148
rect 1711 168 1729 202
rect 1763 168 1901 202
rect 1935 168 1953 202
rect 1711 105 1953 168
rect 38 71 67 105
rect 101 71 159 105
rect 193 71 251 105
rect 285 71 343 105
rect 377 71 435 105
rect 469 71 527 105
rect 561 71 619 105
rect 653 71 711 105
rect 745 71 803 105
rect 837 71 895 105
rect 929 71 987 105
rect 1021 71 1079 105
rect 1113 71 1171 105
rect 1205 71 1263 105
rect 1297 71 1355 105
rect 1389 71 1447 105
rect 1481 71 1539 105
rect 1573 71 1631 105
rect 1665 71 1723 105
rect 1757 71 1815 105
rect 1849 71 1907 105
rect 1941 71 1970 105
<< viali >>
rect 299 1980 333 1982
rect 299 1948 333 1980
rect 472 1972 506 2006
rect 590 1972 624 2006
rect 708 1972 742 2006
rect 826 1972 860 2006
rect 944 1972 978 2006
rect 1062 1972 1096 2006
rect 1180 1972 1214 2006
rect 1298 1972 1332 2006
rect 1416 1972 1450 2006
rect 1534 1972 1568 2006
rect 299 1878 333 1910
rect 299 1876 333 1878
rect 299 1810 333 1838
rect 299 1804 333 1810
rect 299 1742 333 1766
rect 299 1732 333 1742
rect 413 1876 447 1878
rect 413 1844 447 1876
rect 413 1774 447 1806
rect 413 1772 447 1774
rect 531 1876 565 1878
rect 531 1844 565 1876
rect 531 1774 565 1806
rect 531 1772 565 1774
rect 649 1876 683 1878
rect 649 1844 683 1876
rect 649 1774 683 1806
rect 649 1772 683 1774
rect 767 1876 801 1878
rect 767 1844 801 1876
rect 767 1774 801 1806
rect 767 1772 801 1774
rect 885 1876 919 1878
rect 885 1844 919 1876
rect 885 1774 919 1806
rect 885 1772 919 1774
rect 1003 1876 1037 1878
rect 1003 1844 1037 1876
rect 1003 1774 1037 1806
rect 1003 1772 1037 1774
rect 1121 1876 1155 1878
rect 1121 1844 1155 1876
rect 1121 1774 1155 1806
rect 1121 1772 1155 1774
rect 1239 1876 1273 1878
rect 1239 1844 1273 1876
rect 1239 1774 1273 1806
rect 1239 1772 1273 1774
rect 1357 1876 1391 1878
rect 1357 1844 1391 1876
rect 1357 1774 1391 1806
rect 1357 1772 1391 1774
rect 1475 1876 1509 1878
rect 1475 1844 1509 1876
rect 1475 1774 1509 1806
rect 1475 1772 1509 1774
rect 1593 1876 1627 1878
rect 1593 1844 1627 1876
rect 1593 1774 1627 1806
rect 1593 1772 1627 1774
rect 299 1107 333 1137
rect 299 1103 333 1107
rect 299 1039 333 1065
rect 299 1031 333 1039
rect 299 971 333 993
rect 299 959 333 971
rect 413 1104 447 1106
rect 413 1072 447 1104
rect 413 1002 447 1034
rect 413 1000 447 1002
rect 531 1104 565 1106
rect 531 1072 565 1104
rect 531 1002 565 1034
rect 531 1000 565 1002
rect 649 1104 683 1106
rect 649 1072 683 1104
rect 649 1002 683 1034
rect 649 1000 683 1002
rect 767 1104 801 1106
rect 767 1072 801 1104
rect 767 1002 801 1034
rect 767 1000 801 1002
rect 885 1104 919 1106
rect 885 1072 919 1104
rect 885 1002 919 1034
rect 885 1000 919 1002
rect 1003 1104 1037 1106
rect 1003 1072 1037 1104
rect 1003 1002 1037 1034
rect 1003 1000 1037 1002
rect 1121 1104 1155 1106
rect 1121 1072 1155 1104
rect 1121 1002 1155 1034
rect 1121 1000 1155 1002
rect 1239 1104 1273 1106
rect 1239 1072 1273 1104
rect 1239 1002 1273 1034
rect 1239 1000 1273 1002
rect 1357 1104 1391 1106
rect 1357 1072 1391 1104
rect 1357 1002 1391 1034
rect 1357 1000 1391 1002
rect 1475 1104 1509 1106
rect 1475 1072 1509 1104
rect 1475 1002 1509 1034
rect 1475 1000 1509 1002
rect 1593 1104 1627 1106
rect 1593 1072 1627 1104
rect 1593 1002 1627 1034
rect 1593 1000 1627 1002
rect 299 903 333 921
rect 299 887 333 903
rect 472 881 506 915
rect 590 881 624 915
rect 708 881 742 915
rect 826 881 860 915
rect 944 881 978 915
rect 1062 881 1096 915
rect 1180 881 1214 915
rect 1298 881 1332 915
rect 1416 881 1450 915
rect 1534 881 1568 915
rect 67 615 101 649
rect 159 615 193 649
rect 251 615 285 649
rect 343 615 377 649
rect 435 615 469 649
rect 527 615 561 649
rect 619 615 653 649
rect 711 615 745 649
rect 803 615 837 649
rect 895 615 929 649
rect 987 615 1021 649
rect 1079 615 1113 649
rect 1171 615 1205 649
rect 1263 615 1297 649
rect 1355 615 1389 649
rect 1447 615 1481 649
rect 1539 615 1573 649
rect 1631 615 1665 649
rect 1723 615 1757 649
rect 1815 615 1849 649
rect 1907 615 1941 649
rect 1171 377 1205 411
rect 803 337 837 343
rect 803 309 811 337
rect 811 309 837 337
rect 1631 377 1665 411
rect 1288 337 1322 345
rect 1288 311 1305 337
rect 1305 311 1322 337
rect 67 71 101 105
rect 159 71 193 105
rect 251 71 285 105
rect 343 71 377 105
rect 435 71 469 105
rect 527 71 561 105
rect 619 71 653 105
rect 711 71 745 105
rect 803 71 837 105
rect 895 71 929 105
rect 987 71 1021 105
rect 1079 71 1113 105
rect 1171 71 1205 105
rect 1263 71 1297 105
rect 1355 71 1389 105
rect 1447 71 1481 105
rect 1539 71 1573 105
rect 1631 71 1665 105
rect 1723 71 1757 105
rect 1815 71 1849 105
rect 1907 71 1941 105
<< metal1 >>
rect 293 1982 339 2029
rect 293 1948 299 1982
rect 333 1948 339 1982
rect 460 2006 1892 2012
rect 460 1972 472 2006
rect 506 1972 590 2006
rect 624 1972 708 2006
rect 742 1972 826 2006
rect 860 1972 944 2006
rect 978 1972 1062 2006
rect 1096 1972 1180 2006
rect 1214 1972 1298 2006
rect 1332 1972 1416 2006
rect 1450 1972 1534 2006
rect 1568 2000 1892 2006
rect 1568 1972 1836 2000
rect 460 1966 1836 1972
rect 293 1910 339 1948
rect 1832 1948 1836 1966
rect 1888 1948 1892 2000
rect 1832 1936 1892 1948
rect 293 1876 299 1910
rect 333 1876 339 1910
rect 293 1838 339 1876
rect 293 1834 299 1838
rect 128 1804 299 1834
rect 333 1804 339 1838
rect 128 1766 339 1804
rect 128 1732 299 1766
rect 333 1732 339 1766
rect 128 1694 339 1732
rect 407 1878 453 1925
rect 407 1844 413 1878
rect 447 1844 453 1878
rect 407 1806 453 1844
rect 407 1772 413 1806
rect 447 1772 453 1806
rect 128 680 188 1694
rect 407 1395 453 1772
rect 525 1878 571 1925
rect 525 1844 531 1878
rect 565 1844 571 1878
rect 525 1806 571 1844
rect 525 1772 531 1806
rect 565 1772 571 1806
rect 525 1623 571 1772
rect 643 1878 689 1925
rect 643 1844 649 1878
rect 683 1844 689 1878
rect 643 1806 689 1844
rect 643 1772 649 1806
rect 683 1772 689 1806
rect 518 1611 578 1623
rect 518 1559 522 1611
rect 574 1559 578 1611
rect 518 1547 578 1559
rect 518 1495 522 1547
rect 574 1495 578 1547
rect 518 1483 578 1495
rect 400 1383 460 1395
rect 400 1331 404 1383
rect 456 1331 460 1383
rect 400 1319 460 1331
rect 400 1267 404 1319
rect 456 1267 460 1319
rect 400 1255 460 1267
rect 293 1137 339 1184
rect 293 1103 299 1137
rect 333 1103 339 1137
rect 293 1065 339 1103
rect 293 1031 299 1065
rect 333 1031 339 1065
rect 293 993 339 1031
rect 293 959 299 993
rect 333 959 339 993
rect 293 921 339 959
rect 407 1106 453 1255
rect 407 1072 413 1106
rect 447 1072 453 1106
rect 407 1034 453 1072
rect 407 1000 413 1034
rect 447 1000 453 1034
rect 407 953 453 1000
rect 525 1106 571 1483
rect 643 1395 689 1772
rect 761 1878 807 1925
rect 761 1844 767 1878
rect 801 1844 807 1878
rect 761 1806 807 1844
rect 761 1772 767 1806
rect 801 1772 807 1806
rect 761 1623 807 1772
rect 879 1878 925 1925
rect 879 1844 885 1878
rect 919 1844 925 1878
rect 879 1806 925 1844
rect 879 1772 885 1806
rect 919 1772 925 1806
rect 754 1611 814 1623
rect 754 1559 758 1611
rect 810 1559 814 1611
rect 754 1547 814 1559
rect 754 1495 758 1547
rect 810 1495 814 1547
rect 754 1483 814 1495
rect 636 1383 696 1395
rect 636 1331 640 1383
rect 692 1331 696 1383
rect 636 1319 696 1331
rect 636 1267 640 1319
rect 692 1267 696 1319
rect 636 1255 696 1267
rect 525 1072 531 1106
rect 565 1072 571 1106
rect 525 1034 571 1072
rect 525 1000 531 1034
rect 565 1000 571 1034
rect 525 953 571 1000
rect 643 1106 689 1255
rect 643 1072 649 1106
rect 683 1072 689 1106
rect 643 1034 689 1072
rect 643 1000 649 1034
rect 683 1000 689 1034
rect 643 953 689 1000
rect 761 1106 807 1483
rect 879 1395 925 1772
rect 997 1878 1043 1925
rect 997 1844 1003 1878
rect 1037 1844 1043 1878
rect 997 1806 1043 1844
rect 997 1772 1003 1806
rect 1037 1772 1043 1806
rect 997 1623 1043 1772
rect 1115 1878 1161 1925
rect 1115 1844 1121 1878
rect 1155 1844 1161 1878
rect 1115 1806 1161 1844
rect 1115 1772 1121 1806
rect 1155 1772 1161 1806
rect 990 1611 1050 1623
rect 990 1559 994 1611
rect 1046 1559 1050 1611
rect 990 1547 1050 1559
rect 990 1495 994 1547
rect 1046 1495 1050 1547
rect 990 1483 1050 1495
rect 872 1383 932 1395
rect 872 1331 876 1383
rect 928 1331 932 1383
rect 872 1319 932 1331
rect 872 1267 876 1319
rect 928 1267 932 1319
rect 872 1255 932 1267
rect 761 1072 767 1106
rect 801 1072 807 1106
rect 761 1034 807 1072
rect 761 1000 767 1034
rect 801 1000 807 1034
rect 761 953 807 1000
rect 879 1106 925 1255
rect 879 1072 885 1106
rect 919 1072 925 1106
rect 879 1034 925 1072
rect 879 1000 885 1034
rect 919 1000 925 1034
rect 879 953 925 1000
rect 997 1106 1043 1483
rect 1115 1395 1161 1772
rect 1233 1878 1279 1925
rect 1233 1844 1239 1878
rect 1273 1844 1279 1878
rect 1233 1806 1279 1844
rect 1233 1772 1239 1806
rect 1273 1772 1279 1806
rect 1233 1623 1279 1772
rect 1351 1878 1397 1925
rect 1351 1844 1357 1878
rect 1391 1844 1397 1878
rect 1351 1806 1397 1844
rect 1351 1772 1357 1806
rect 1391 1772 1397 1806
rect 1226 1611 1286 1623
rect 1226 1559 1230 1611
rect 1282 1559 1286 1611
rect 1226 1547 1286 1559
rect 1226 1495 1230 1547
rect 1282 1495 1286 1547
rect 1226 1483 1286 1495
rect 1108 1383 1168 1395
rect 1108 1331 1112 1383
rect 1164 1331 1168 1383
rect 1108 1319 1168 1331
rect 1108 1267 1112 1319
rect 1164 1267 1168 1319
rect 1108 1255 1168 1267
rect 997 1072 1003 1106
rect 1037 1072 1043 1106
rect 997 1034 1043 1072
rect 997 1000 1003 1034
rect 1037 1000 1043 1034
rect 997 953 1043 1000
rect 1115 1106 1161 1255
rect 1115 1072 1121 1106
rect 1155 1072 1161 1106
rect 1115 1034 1161 1072
rect 1115 1000 1121 1034
rect 1155 1000 1161 1034
rect 1115 953 1161 1000
rect 1233 1106 1279 1483
rect 1351 1395 1397 1772
rect 1469 1878 1515 1925
rect 1469 1844 1475 1878
rect 1509 1844 1515 1878
rect 1469 1806 1515 1844
rect 1469 1772 1475 1806
rect 1509 1772 1515 1806
rect 1469 1623 1515 1772
rect 1587 1878 1633 1925
rect 1587 1844 1593 1878
rect 1627 1844 1633 1878
rect 1832 1884 1836 1936
rect 1888 1884 1892 1936
rect 1832 1872 1892 1884
rect 1587 1806 1633 1844
rect 1587 1772 1593 1806
rect 1627 1772 1633 1806
rect 1462 1611 1522 1623
rect 1462 1559 1466 1611
rect 1518 1559 1522 1611
rect 1462 1547 1522 1559
rect 1462 1495 1466 1547
rect 1518 1495 1522 1547
rect 1462 1483 1522 1495
rect 1344 1383 1404 1395
rect 1344 1331 1348 1383
rect 1400 1331 1404 1383
rect 1344 1319 1404 1331
rect 1344 1267 1348 1319
rect 1400 1267 1404 1319
rect 1344 1255 1404 1267
rect 1233 1072 1239 1106
rect 1273 1072 1279 1106
rect 1233 1034 1279 1072
rect 1233 1000 1239 1034
rect 1273 1000 1279 1034
rect 1233 953 1279 1000
rect 1351 1106 1397 1255
rect 1351 1072 1357 1106
rect 1391 1072 1397 1106
rect 1351 1034 1397 1072
rect 1351 1000 1357 1034
rect 1391 1000 1397 1034
rect 1351 953 1397 1000
rect 1469 1106 1515 1483
rect 1587 1395 1633 1772
rect 1580 1383 1640 1395
rect 1580 1331 1584 1383
rect 1636 1331 1640 1383
rect 1580 1319 1640 1331
rect 1580 1267 1584 1319
rect 1636 1267 1640 1319
rect 1580 1255 1640 1267
rect 1469 1072 1475 1106
rect 1509 1072 1515 1106
rect 1469 1034 1515 1072
rect 1469 1000 1475 1034
rect 1509 1000 1515 1034
rect 1469 953 1515 1000
rect 1587 1106 1633 1255
rect 1587 1072 1593 1106
rect 1627 1072 1633 1106
rect 1587 1034 1633 1072
rect 1587 1000 1593 1034
rect 1627 1000 1633 1034
rect 1587 953 1633 1000
rect 293 895 299 921
rect 286 887 299 895
rect 333 895 339 921
rect 460 917 1580 921
rect 460 915 962 917
rect 333 887 346 895
rect 286 883 346 887
rect 286 831 290 883
rect 342 831 346 883
rect 460 881 472 915
rect 506 881 590 915
rect 624 881 708 915
rect 742 881 826 915
rect 860 881 944 915
rect 460 875 962 881
rect 950 865 962 875
rect 1014 865 1026 917
rect 1078 915 1580 917
rect 1096 881 1180 915
rect 1214 881 1298 915
rect 1332 881 1416 915
rect 1450 881 1534 915
rect 1568 881 1580 915
rect 1078 875 1580 881
rect 1078 865 1090 875
rect 950 861 1090 865
rect 286 819 346 831
rect 286 767 290 819
rect 342 767 346 819
rect 286 755 346 767
rect 38 649 1970 680
rect 38 615 67 649
rect 101 615 159 649
rect 193 615 251 649
rect 285 615 343 649
rect 377 615 435 649
rect 469 615 527 649
rect 561 615 619 649
rect 653 615 711 649
rect 745 615 803 649
rect 837 615 895 649
rect 929 615 987 649
rect 1021 615 1079 649
rect 1113 615 1171 649
rect 1205 615 1263 649
rect 1297 615 1355 649
rect 1389 615 1447 649
rect 1481 615 1539 649
rect 1573 615 1631 649
rect 1665 615 1723 649
rect 1757 615 1815 649
rect 1849 615 1907 649
rect 1941 615 1970 649
rect 38 584 1970 615
rect 1158 420 1218 426
rect 1158 368 1162 420
rect 1214 368 1218 420
rect 1158 358 1218 368
rect 1622 420 1674 426
rect 1622 362 1674 368
rect 794 352 846 358
rect 794 294 846 300
rect 1158 345 1341 358
rect 1158 311 1288 345
rect 1322 311 1341 345
rect 1158 298 1341 311
rect 38 111 1970 136
rect 38 105 258 111
rect 38 71 67 105
rect 101 71 159 105
rect 193 71 251 105
rect 38 59 258 71
rect 310 59 322 111
rect 374 105 1970 111
rect 377 71 435 105
rect 469 71 527 105
rect 561 71 619 105
rect 653 71 711 105
rect 745 71 803 105
rect 837 71 895 105
rect 929 71 987 105
rect 1021 71 1079 105
rect 1113 71 1171 105
rect 1205 71 1263 105
rect 1297 71 1355 105
rect 1389 71 1447 105
rect 1481 71 1539 105
rect 1573 71 1631 105
rect 1665 71 1723 105
rect 1757 71 1815 105
rect 1849 71 1907 105
rect 1941 71 1970 105
rect 374 59 1970 71
rect 38 40 1970 59
<< via1 >>
rect 1836 1948 1888 2000
rect 522 1559 574 1611
rect 522 1495 574 1547
rect 404 1331 456 1383
rect 404 1267 456 1319
rect 758 1559 810 1611
rect 758 1495 810 1547
rect 640 1331 692 1383
rect 640 1267 692 1319
rect 994 1559 1046 1611
rect 994 1495 1046 1547
rect 876 1331 928 1383
rect 876 1267 928 1319
rect 1230 1559 1282 1611
rect 1230 1495 1282 1547
rect 1112 1331 1164 1383
rect 1112 1267 1164 1319
rect 1836 1884 1888 1936
rect 1466 1559 1518 1611
rect 1466 1495 1518 1547
rect 1348 1331 1400 1383
rect 1348 1267 1400 1319
rect 1584 1331 1636 1383
rect 1584 1267 1636 1319
rect 962 915 1014 917
rect 290 831 342 883
rect 962 881 978 915
rect 978 881 1014 915
rect 962 865 1014 881
rect 1026 915 1078 917
rect 1026 881 1062 915
rect 1062 881 1078 915
rect 1026 865 1078 881
rect 290 767 342 819
rect 1162 411 1214 420
rect 1162 377 1171 411
rect 1171 377 1205 411
rect 1205 377 1214 411
rect 1162 368 1214 377
rect 1622 411 1674 420
rect 1622 377 1631 411
rect 1631 377 1665 411
rect 1665 377 1674 411
rect 1622 368 1674 377
rect 794 343 846 352
rect 794 309 803 343
rect 803 309 837 343
rect 837 309 846 343
rect 794 300 846 309
rect 258 105 310 111
rect 258 71 285 105
rect 285 71 310 105
rect 258 59 310 71
rect 322 105 374 111
rect 322 71 343 105
rect 343 71 374 105
rect 322 59 374 71
<< metal2 >>
rect 954 1613 1054 2308
rect 1822 2000 1902 2002
rect 1822 1948 1836 2000
rect 1888 1948 1902 2000
rect 1822 1936 1902 1948
rect 1822 1884 1836 1936
rect 1888 1884 1902 1936
rect 1822 1882 1902 1884
rect 508 1611 588 1613
rect 508 1559 522 1611
rect 574 1573 588 1611
rect 744 1611 824 1613
rect 744 1573 758 1611
rect 574 1559 758 1573
rect 810 1573 824 1611
rect 954 1611 1060 1613
rect 954 1573 994 1611
rect 810 1559 994 1573
rect 1046 1573 1060 1611
rect 1216 1611 1296 1613
rect 1216 1573 1230 1611
rect 1046 1559 1230 1573
rect 1282 1573 1296 1611
rect 1452 1611 1532 1613
rect 1452 1573 1466 1611
rect 1282 1559 1466 1573
rect 1518 1573 1532 1611
rect 1518 1559 1650 1573
rect 508 1547 1650 1559
rect 508 1495 522 1547
rect 574 1495 758 1547
rect 810 1495 994 1547
rect 1046 1495 1230 1547
rect 1282 1495 1466 1547
rect 1518 1495 1650 1547
rect 508 1493 1650 1495
rect 310 1393 390 1405
rect 310 1337 322 1393
rect 378 1385 390 1393
rect 1650 1393 1730 1405
rect 1650 1385 1662 1393
rect 378 1383 1662 1385
rect 378 1337 404 1383
rect 310 1331 404 1337
rect 456 1331 640 1383
rect 692 1331 876 1383
rect 928 1331 1112 1383
rect 1164 1331 1348 1383
rect 1400 1331 1584 1383
rect 1636 1337 1662 1383
rect 1718 1337 1730 1393
rect 1636 1331 1730 1337
rect 310 1319 1730 1331
rect 310 1313 404 1319
rect 310 1257 322 1313
rect 378 1267 404 1313
rect 456 1305 640 1319
rect 456 1267 470 1305
rect 378 1265 470 1267
rect 626 1267 640 1305
rect 692 1305 876 1319
rect 692 1267 706 1305
rect 626 1265 706 1267
rect 862 1267 876 1305
rect 928 1305 1112 1319
rect 928 1267 942 1305
rect 862 1265 942 1267
rect 1098 1267 1112 1305
rect 1164 1305 1348 1319
rect 1164 1267 1178 1305
rect 1098 1265 1178 1267
rect 1334 1267 1348 1305
rect 1400 1305 1584 1319
rect 1400 1267 1414 1305
rect 1334 1265 1414 1267
rect 1570 1267 1584 1305
rect 1636 1313 1730 1319
rect 1636 1267 1662 1313
rect 1570 1265 1662 1267
rect 378 1257 390 1265
rect 310 1245 390 1257
rect 1650 1257 1662 1265
rect 1718 1257 1730 1313
rect 1650 1245 1730 1257
rect 960 917 1080 931
rect 276 883 356 885
rect 276 831 290 883
rect 342 831 356 883
rect 960 865 962 917
rect 1014 865 1026 917
rect 1078 865 1080 917
rect 960 851 1080 865
rect 276 819 356 831
rect 276 767 290 819
rect 342 767 356 819
rect 276 125 356 767
rect 788 352 852 358
rect 788 300 794 352
rect 846 300 852 352
rect 256 111 376 125
rect 256 59 258 111
rect 310 59 322 111
rect 374 59 376 111
rect 256 45 376 59
rect 788 -40 852 300
rect 990 260 1050 851
rect 1832 769 1892 1882
rect 1158 709 1892 769
rect 1158 420 1218 709
rect 1156 368 1162 420
rect 1214 368 1220 420
rect 1616 368 1622 420
rect 1674 368 1680 420
rect 1158 361 1218 368
rect 1618 260 1678 368
rect 990 200 1678 260
<< via2 >>
rect 322 1337 378 1393
rect 1662 1337 1718 1393
rect 322 1257 378 1313
rect 1662 1257 1718 1313
<< metal3 >>
rect 310 1393 1730 1405
rect 310 1337 322 1393
rect 378 1337 1662 1393
rect 1718 1337 1730 1393
rect 310 1313 1730 1337
rect 310 1257 322 1313
rect 378 1257 1662 1313
rect 1718 1257 1730 1313
rect 310 1245 1730 1257
<< labels >>
flabel metal2 s 954 2258 1054 2308 2 FreeSans 44 0 0 0 out
port 2 nsew
flabel metal2 s 788 -40 852 -9 2 FreeSans 44 0 0 0 en
port 3 nsew
flabel metal1 s 38 584 88 680 2 FreeSans 44 0 0 0 vdd
port 5 nsew
flabel metal1 s 38 40 88 136 2 FreeSans 44 0 0 0 vss
port 6 nsew
flabel metal3 s 1000 1245 1040 1405 2 FreeSans 96 0 0 0 in
port 7 nsew
rlabel comment 1694 88 1694 88 4 decap_3_0.decap_3
rlabel comment 38 88 38 88 4 decap_8_0.decap_8
rlabel comment 1234 88 1234 88 4 inv_4_0.inv_4
flabel comment 1648 258 1648 258 0 FreeSans 340 0 0 0 inv_4_0.Y
flabel comment 1648 326 1648 326 0 FreeSans 340 0 0 0 inv_4_0.Y
flabel comment 1648 394 1648 394 0 FreeSans 340 0 0 0 inv_4_0.Y
flabel comment 1280 326 1280 326 0 FreeSans 340 0 0 0 inv_4_0.A
flabel comment 1372 326 1372 326 0 FreeSans 340 0 0 0 inv_4_0.A
flabel comment 1464 326 1464 326 0 FreeSans 340 0 0 0 inv_4_0.A
flabel comment 1556 326 1556 326 0 FreeSans 340 0 0 0 inv_4_0.A
rlabel comment 774 88 774 88 4 inv_4_1.inv_4
flabel comment 1188 258 1188 258 0 FreeSans 340 0 0 0 inv_4_1.Y
flabel comment 1188 326 1188 326 0 FreeSans 340 0 0 0 inv_4_1.Y
flabel comment 1188 394 1188 394 0 FreeSans 340 0 0 0 inv_4_1.Y
flabel comment 820 326 820 326 0 FreeSans 340 0 0 0 inv_4_1.A
flabel comment 912 326 912 326 0 FreeSans 340 0 0 0 inv_4_1.A
flabel comment 1004 326 1004 326 0 FreeSans 340 0 0 0 inv_4_1.A
flabel comment 1096 326 1096 326 0 FreeSans 340 0 0 0 inv_4_1.A
<< end >>
