magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 590 542
<< pwell >>
rect 1 -19 551 143
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 473 117
<< scpmoshvt >>
rect 79 283 473 457
<< ndiff >>
rect 27 72 79 117
rect 27 38 35 72
rect 69 38 79 72
rect 27 7 79 38
rect 473 72 525 117
rect 473 38 483 72
rect 517 38 525 72
rect 473 7 525 38
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 343 79 411
rect 27 309 35 343
rect 69 309 79 343
rect 27 283 79 309
rect 473 445 525 457
rect 473 411 483 445
rect 517 411 525 445
rect 473 343 525 411
rect 473 309 483 343
rect 517 309 525 343
rect 473 283 525 309
<< ndiffc >>
rect 35 38 69 72
rect 483 38 517 72
<< pdiffc >>
rect 35 411 69 445
rect 35 309 69 343
rect 483 411 517 445
rect 483 309 517 343
<< poly >>
rect 79 457 473 483
rect 79 257 473 283
rect 79 235 255 257
rect 79 201 95 235
rect 129 201 205 235
rect 239 201 255 235
rect 79 185 255 201
rect 297 199 473 215
rect 297 165 313 199
rect 347 165 423 199
rect 457 165 473 199
rect 297 143 473 165
rect 79 117 473 143
rect 79 -19 473 7
<< polycont >>
rect 95 201 129 235
rect 205 201 239 235
rect 313 165 347 199
rect 423 165 457 199
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 552 521
rect 17 445 535 487
rect 17 411 35 445
rect 69 411 483 445
rect 517 411 535 445
rect 17 343 535 411
rect 17 309 35 343
rect 69 309 483 343
rect 517 309 535 343
rect 17 269 535 309
rect 17 201 95 235
rect 129 201 205 235
rect 239 201 259 235
rect 17 131 259 201
rect 293 199 535 269
rect 293 165 313 199
rect 347 165 423 199
rect 457 165 535 199
rect 17 72 535 131
rect 17 38 35 72
rect 69 38 483 72
rect 517 38 535 72
rect 17 -23 535 38
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 552 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
<< metal1 >>
rect 0 521 552 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 552 521
rect 0 456 552 487
rect 0 -23 552 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 552 -23
rect 0 -88 552 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 decap_6
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
<< properties >>
string FIXED_BBOX 0 -40 552 504
string path 0.000 -1.000 13.800 -1.000 
<< end >>
