magic
tech sky130B
magscale 1 2
timestamp 1697571680
<< nwell >>
rect -410 -198 1590 -100
rect -410 -202 -237 -198
rect 878 -519 1590 -198
<< nsubdiff >>
rect -199 -166 78 -165
rect -199 -200 -171 -166
rect -137 -200 78 -166
rect -199 -211 78 -200
<< nsubdiffcont >>
rect -171 -200 -137 -166
<< locali >>
rect 1211 726 1245 823
rect 1210 171 1245 252
rect -200 -166 82 -142
rect -200 -200 -171 -166
rect -137 -200 82 -166
rect -200 -229 82 -200
rect 759 -496 761 -456
rect 795 -496 798 -456
rect 397 -521 560 -520
rect 437 -561 560 -521
rect 759 -616 798 -496
rect 978 -564 1074 -525
rect 1207 -628 1246 -567
<< viali >>
rect 1211 692 1245 726
rect 1207 252 1247 292
rect 761 -496 795 -456
rect 397 -561 437 -521
rect 938 -565 978 -525
rect 1206 -567 1246 -527
<< metal1 >>
rect -32 902 20 908
rect -34 852 -32 891
rect 898 898 950 904
rect 20 891 151 896
rect 20 852 898 891
rect -32 844 20 850
rect 950 852 1080 891
rect 898 840 950 846
rect 1199 726 1257 732
rect -85 477 -49 687
rect 23 622 29 674
rect 81 622 87 674
rect 150 477 186 719
rect 262 676 314 682
rect 256 624 262 676
rect 314 624 320 676
rect 262 618 314 624
rect -85 476 186 477
rect 387 476 423 707
rect 492 624 498 676
rect 550 624 556 676
rect 622 476 658 722
rect 1199 692 1211 726
rect 1245 692 1336 726
rect 1199 686 1257 692
rect 730 624 736 676
rect 788 624 794 676
rect 862 476 898 665
rect 964 624 970 676
rect 1022 624 1028 676
rect 1095 476 1131 668
rect -85 475 1131 476
rect -251 439 1131 475
rect -85 237 -49 439
rect 23 218 29 270
rect 81 218 87 270
rect 150 224 186 439
rect 256 202 262 254
rect 314 202 320 254
rect 387 141 423 439
rect 498 250 550 256
rect 492 198 498 250
rect 550 198 556 250
rect 622 224 658 439
rect 498 192 550 198
rect 730 186 736 238
rect 788 186 794 238
rect 862 232 898 439
rect 964 190 970 242
rect 1022 190 1028 242
rect 1095 201 1131 439
rect 1201 298 1253 304
rect 1201 240 1253 246
rect 1077 73 1083 80
rect -36 34 1083 73
rect 1077 28 1083 34
rect 1135 28 1141 80
rect 1302 -202 1336 692
rect 743 -502 749 -450
rect 801 -502 807 -450
rect 385 -567 391 -515
rect 443 -567 449 -515
rect 932 -519 984 -513
rect 932 -577 984 -571
rect 1194 -573 1200 -521
rect 1252 -573 1258 -521
rect 1418 -807 1424 -755
rect 1476 -807 1482 -755
<< via1 >>
rect -32 850 20 902
rect 898 846 950 898
rect 29 622 81 674
rect 262 624 314 676
rect 498 624 550 676
rect 736 624 788 676
rect 970 624 1022 676
rect 29 218 81 270
rect 262 202 314 254
rect 498 198 550 250
rect 736 186 788 238
rect 970 190 1022 242
rect 1201 292 1253 298
rect 1201 252 1207 292
rect 1207 252 1247 292
rect 1247 252 1253 292
rect 1201 246 1253 252
rect 1083 28 1135 80
rect 749 -456 801 -450
rect 749 -496 761 -456
rect 761 -496 795 -456
rect 795 -496 801 -456
rect 749 -502 801 -496
rect 391 -521 443 -515
rect 391 -561 397 -521
rect 397 -561 437 -521
rect 437 -561 443 -521
rect 391 -567 443 -561
rect 932 -525 984 -519
rect 932 -565 938 -525
rect 938 -565 978 -525
rect 978 -565 984 -525
rect 932 -571 984 -565
rect 1200 -527 1252 -521
rect 1200 -567 1206 -527
rect 1206 -567 1246 -527
rect 1246 -567 1252 -527
rect 1200 -573 1252 -567
rect 1424 -807 1476 -755
<< metal2 >>
rect -38 895 -32 902
rect -147 856 -32 895
rect -147 -347 -108 856
rect -38 850 -32 856
rect 20 850 26 902
rect 892 846 898 898
rect 950 846 956 898
rect 29 674 81 680
rect 262 676 314 682
rect 498 676 550 682
rect 256 624 262 676
rect 314 624 320 676
rect 29 616 81 622
rect 262 618 314 624
rect 498 618 550 624
rect 736 676 788 682
rect 736 618 788 624
rect 970 676 1022 682
rect 970 618 1022 624
rect 36 477 74 616
rect 269 477 307 618
rect 36 475 307 477
rect 505 475 543 618
rect 743 477 781 618
rect 977 479 1015 618
rect 977 477 1375 479
rect 743 475 1375 477
rect 36 441 1375 475
rect 36 439 1015 441
rect 36 276 74 439
rect 269 437 781 439
rect 29 270 81 276
rect 269 260 307 437
rect 29 212 81 218
rect 262 254 314 260
rect 505 256 543 437
rect 498 250 550 256
rect 262 196 314 202
rect 492 198 498 250
rect 550 198 556 250
rect 743 244 781 437
rect 977 248 1015 439
rect 736 238 788 244
rect 498 192 550 198
rect 736 180 788 186
rect 970 242 1022 248
rect 1195 246 1201 298
rect 1253 289 1259 298
rect 1253 254 1467 289
rect 1253 246 1259 254
rect 970 184 1022 190
rect 1083 80 1135 86
rect 1135 35 1245 74
rect 1083 22 1135 28
rect 899 -347 938 -346
rect -147 -386 938 -347
rect 755 -444 794 -386
rect 749 -450 801 -444
rect 749 -508 801 -502
rect 391 -515 443 -509
rect 899 -519 938 -386
rect 1206 -515 1245 35
rect 899 -565 932 -519
rect 391 -573 443 -567
rect 926 -571 932 -565
rect 984 -571 990 -519
rect 1200 -521 1252 -515
rect 396 -892 437 -573
rect 1200 -579 1252 -573
rect 1432 -749 1467 254
rect 1424 -755 1476 -749
rect 1424 -813 1476 -807
use sky130_fd_pr__nfet_01v8_JJRV6Y  sky130_fd_pr__nfet_01v8_JJRV6Y_0
timestamp 1696895721
transform 1 0 523 0 -1 179
box -757 -279 757 279
use sky130_fd_pr__pfet_01v8_VVAZD4  sky130_fd_pr__pfet_01v8_VVAZD4_0
timestamp 1696984848
transform 1 0 525 0 1 743
box -757 -284 757 284
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0
timestamp 1693170804
transform 1 0 1275 0 1 -780
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_0
timestamp 1693170804
transform 1 0 -372 0 1 -780
box -38 -48 774 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1693170804
transform 1 0 815 0 1 -780
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_1
timestamp 1693170804
transform 1 0 362 0 1 -780
box -38 -48 498 592
<< labels >>
flabel metal2 1337 441 1375 479 0 FreeSans 640 0 0 0 out
port 0 nsew
flabel metal1 -251 439 -215 475 0 FreeSans 640 0 0 0 in
port 4 nsew
flabel metal2 396 -892 437 -851 0 FreeSans 640 0 0 0 en
port 1 nsew
flabel metal1 1302 683 1336 717 0 FreeSans 640 0 0 0 vdd
port 3 nsew
flabel metal2 1432 247 1467 286 0 FreeSans 640 0 0 0 vss
port 2 nsew
<< end >>
