magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 498 542
<< pwell >>
rect 1 -19 443 163
rect 30 -57 64 -19
<< scnmos >>
rect 83 7 113 137
rect 167 7 197 137
rect 251 7 281 137
rect 335 7 365 137
<< scpmoshvt >>
rect 83 257 113 457
rect 167 257 197 457
rect 251 257 281 457
rect 335 257 365 457
<< ndiff >>
rect 27 123 83 137
rect 27 89 39 123
rect 73 89 83 123
rect 27 55 83 89
rect 27 21 39 55
rect 73 21 83 55
rect 27 7 83 21
rect 113 123 167 137
rect 113 89 123 123
rect 157 89 167 123
rect 113 55 167 89
rect 113 21 123 55
rect 157 21 167 55
rect 113 7 167 21
rect 197 55 251 137
rect 197 21 207 55
rect 241 21 251 55
rect 197 7 251 21
rect 281 123 335 137
rect 281 89 291 123
rect 325 89 335 123
rect 281 55 335 89
rect 281 21 291 55
rect 325 21 335 55
rect 281 7 335 21
rect 365 55 417 137
rect 365 21 375 55
rect 409 21 417 55
rect 365 7 417 21
<< pdiff >>
rect 27 437 83 457
rect 27 403 39 437
rect 73 403 83 437
rect 27 369 83 403
rect 27 335 39 369
rect 73 335 83 369
rect 27 301 83 335
rect 27 267 39 301
rect 73 267 83 301
rect 27 257 83 267
rect 113 445 167 457
rect 113 411 123 445
rect 157 411 167 445
rect 113 377 167 411
rect 113 343 123 377
rect 157 343 167 377
rect 113 257 167 343
rect 197 437 251 457
rect 197 403 207 437
rect 241 403 251 437
rect 197 369 251 403
rect 197 335 207 369
rect 241 335 251 369
rect 197 301 251 335
rect 197 267 207 301
rect 241 267 251 301
rect 197 257 251 267
rect 281 369 335 457
rect 281 335 291 369
rect 325 335 335 369
rect 281 301 335 335
rect 281 267 291 301
rect 325 267 335 301
rect 281 257 335 267
rect 365 445 417 457
rect 365 411 375 445
rect 409 411 417 445
rect 365 377 417 411
rect 365 343 375 377
rect 409 343 417 377
rect 365 257 417 343
<< ndiffc >>
rect 39 89 73 123
rect 39 21 73 55
rect 123 89 157 123
rect 123 21 157 55
rect 207 21 241 55
rect 291 89 325 123
rect 291 21 325 55
rect 375 21 409 55
<< pdiffc >>
rect 39 403 73 437
rect 39 335 73 369
rect 39 267 73 301
rect 123 411 157 445
rect 123 343 157 377
rect 207 403 241 437
rect 207 335 241 369
rect 207 267 241 301
rect 291 335 325 369
rect 291 267 325 301
rect 375 411 409 445
rect 375 343 409 377
<< poly >>
rect 83 457 113 483
rect 167 457 197 483
rect 251 457 281 483
rect 335 457 365 483
rect 83 225 113 257
rect 167 225 197 257
rect 83 209 197 225
rect 83 175 112 209
rect 146 175 197 209
rect 83 159 197 175
rect 83 137 113 159
rect 167 137 197 159
rect 251 225 281 257
rect 335 225 365 257
rect 251 209 365 225
rect 251 175 291 209
rect 325 175 365 209
rect 251 159 365 175
rect 251 137 281 159
rect 335 137 365 159
rect 83 -19 113 7
rect 167 -19 197 7
rect 251 -19 281 7
rect 335 -19 365 7
<< polycont >>
rect 112 175 146 209
rect 291 175 325 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 18 437 73 453
rect 18 403 39 437
rect 18 369 73 403
rect 18 335 39 369
rect 18 301 73 335
rect 107 445 173 487
rect 107 411 123 445
rect 157 411 173 445
rect 107 377 173 411
rect 107 343 123 377
rect 157 343 173 377
rect 107 327 173 343
rect 207 445 435 453
rect 207 437 375 445
rect 241 419 375 437
rect 207 369 241 403
rect 409 411 435 445
rect 18 267 39 301
rect 207 301 241 335
rect 73 267 207 293
rect 18 251 241 267
rect 275 369 341 385
rect 275 335 291 369
rect 325 335 341 369
rect 275 301 341 335
rect 375 377 435 411
rect 409 343 435 377
rect 375 327 435 343
rect 275 267 291 301
rect 325 293 341 301
rect 325 267 427 293
rect 275 249 427 267
rect 18 209 162 215
rect 18 175 112 209
rect 146 175 162 209
rect 196 209 350 215
rect 196 175 291 209
rect 325 175 350 209
rect 384 141 427 249
rect 18 123 73 141
rect 18 89 39 123
rect 18 55 73 89
rect 18 21 39 55
rect 18 -23 73 21
rect 107 123 427 141
rect 107 89 123 123
rect 157 105 291 123
rect 157 89 173 105
rect 107 55 173 89
rect 275 89 291 105
rect 325 107 427 123
rect 325 89 341 107
rect 107 21 123 55
rect 157 21 173 55
rect 107 11 173 21
rect 207 55 241 71
rect 207 -23 241 21
rect 275 55 341 89
rect 275 21 291 55
rect 325 21 341 55
rect 275 11 341 21
rect 375 55 433 71
rect 409 21 433 55
rect 375 -23 433 21
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
<< metal1 >>
rect 0 521 460 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 0 456 460 487
rect 0 -23 460 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
rect 0 -88 460 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 nor2_2
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 214 181 248 215 0 FreeSans 400 0 0 0 B
port 8 nsew
flabel locali s 306 317 340 351 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel locali s 30 181 64 215 0 FreeSans 400 0 0 0 A
port 10 nsew
<< properties >>
string FIXED_BBOX 0 -40 460 504
string path 0.000 -1.000 11.500 -1.000 
<< end >>
