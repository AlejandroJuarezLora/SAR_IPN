magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< metal1 >>
rect 136 709 654 755
rect 136 409 182 709
rect 254 409 300 619
rect 372 409 418 709
rect 490 409 536 619
rect 608 409 654 709
rect 799 709 1081 755
rect 799 409 845 709
rect 917 409 963 619
rect 1035 409 1081 709
rect 1226 409 1272 755
rect 1344 409 1390 619
rect 1462 409 1508 755
rect 1771 709 2525 755
rect 1653 409 1699 619
rect 1771 409 1817 709
rect 1889 409 1935 619
rect 2007 409 2053 709
rect 2125 409 2171 619
rect 2243 409 2289 709
rect 2361 409 2407 619
rect 2479 409 2525 709
rect 2597 409 2643 619
rect 189 131 601 177
rect 852 131 1028 177
rect 1186 131 1279 177
rect 1455 131 1548 177
rect 1706 131 2590 177
<< metal2 >>
rect 12 519 2768 579
rect 12 359 72 519
rect 2708 359 2768 519
rect 365 -40 425 1
rect 910 -40 970 1
rect 1186 -40 1246 1
rect 1488 -40 1548 1
rect 2118 -40 2178 1
use Guardring_N_2  Guardring_N_2_0
timestamp 1696364841
transform 1 0 -2251 0 1 983
box 2250 -987 5032 -409
use M1_1  M1_1_0
timestamp 1696364841
transform 1 0 1308 0 1 318
box -114 -197 114 117
use M1_1  M1_1_1
timestamp 1696364841
transform 1 0 2561 0 1 318
box -114 -197 114 117
use M1_1  M1_1_2
timestamp 1696364841
transform 1 0 1735 0 1 318
box -114 -197 114 117
use M1_1  M1_1_3
timestamp 1696364841
transform 1 0 1853 0 1 318
box -114 -197 114 117
use M1_1  M1_1_4
timestamp 1696364841
transform 1 0 1971 0 1 318
box -114 -197 114 117
use M1_1  M1_1_5
timestamp 1696364841
transform 1 0 2207 0 1 318
box -114 -197 114 117
use M1_1  M1_1_6
timestamp 1696364841
transform 1 0 2325 0 1 318
box -114 -197 114 117
use M1_1  M1_1_7
timestamp 1696364841
transform 1 0 2089 0 1 318
box -114 -197 114 117
use M1_1  M1_1_8
timestamp 1696364841
transform 1 0 2443 0 1 318
box -114 -197 114 117
use M1_1  M1_1_9
timestamp 1696364841
transform 1 0 1426 0 1 318
box -114 -197 114 117
use M1_1  M1_1_10
timestamp 1696364841
transform 1 0 336 0 1 318
box -114 -197 114 117
use M1_1  M1_1_11
timestamp 1696364841
transform 1 0 454 0 1 318
box -114 -197 114 117
use M1_1  M1_1_12
timestamp 1696364841
transform 1 0 572 0 1 318
box -114 -197 114 117
use M1_1  M1_1_13
timestamp 1696364841
transform 1 0 218 0 1 318
box -114 -197 114 117
use M1_1  M1_1_14
timestamp 1696364841
transform 1 0 881 0 1 318
box -114 -197 114 117
use M1_1  M1_1_15
timestamp 1696364841
transform 1 0 999 0 1 318
box -114 -197 114 117
use via1_1  via1_1_0
timestamp 1696364841
transform 0 -1 25 1 0 269
box -6 -46 124 12
use via1_1  via1_1_1
timestamp 1696364841
transform 0 -1 2721 1 0 269
box -6 -46 124 12
use via2  via2_0
timestamp 1696364841
transform 0 1 2148 -1 0 131
box 0 -40 140 40
use via2  via2_1
timestamp 1696364841
transform 0 1 395 -1 0 131
box 0 -40 140 40
use via2  via2_2
timestamp 1696364841
transform 0 1 940 -1 0 131
box 0 -40 140 40
use via2  via2_3
timestamp 1696364841
transform 0 1 1518 -1 0 131
box 0 -40 140 40
use via2  via2_4
timestamp 1696364841
transform 0 -1 1216 -1 0 131
box 0 -40 140 40
use via2  via2_5
timestamp 1696364841
transform 0 -1 277 -1 0 619
box 0 -40 140 40
use via2  via2_6
timestamp 1696364841
transform 0 -1 1676 -1 0 619
box 0 -40 140 40
use via2  via2_7
timestamp 1696364841
transform 0 -1 513 -1 0 619
box 0 -40 140 40
use via2  via2_8
timestamp 1696364841
transform 0 -1 1912 -1 0 619
box 0 -40 140 40
use via2  via2_9
timestamp 1696364841
transform 0 -1 940 -1 0 619
box 0 -40 140 40
use via2  via2_10
timestamp 1696364841
transform 0 -1 1367 -1 0 619
box 0 -40 140 40
use via2  via2_11
timestamp 1696364841
transform 0 -1 2148 -1 0 619
box 0 -40 140 40
use via2  via2_12
timestamp 1696364841
transform 0 -1 2384 -1 0 619
box 0 -40 140 40
use via2  via2_13
timestamp 1696364841
transform 0 -1 2620 -1 0 619
box 0 -40 140 40
use via2  via2_14
timestamp 1696364841
transform 0 -1 42 -1 0 398
box 0 -40 140 40
use via2  via2_15
timestamp 1696364841
transform 0 -1 2738 -1 0 398
box 0 -40 140 40
<< labels >>
flabel metal2 s 1186 -40 1246 1 3 FreeSans 224 270 0 0 d_0
port 2 nsew
flabel metal2 s 1488 -40 1548 1 3 FreeSans 44 270 0 0 d_1
port 3 nsew
flabel metal2 s 910 -40 970 1 3 FreeSans 44 270 0 0 d_2
port 4 nsew
flabel metal2 s 365 -40 425 1 3 FreeSans 44 270 0 0 d_3
port 5 nsew
flabel metal2 s 2118 -40 2178 1 3 FreeSans 44 270 0 0 d_4
port 6 nsew
flabel metal2 s 12 519 62 579 2 FreeSans 44 0 0 0 vss
port 7 nsew
<< properties >>
string path 7.390 0.770 7.625 0.770 
<< end >>
