* SPICE3 file created from dac_flat.ext - technology: sky130B

.subckt dac ctl0 ctl1 ctl2 ctl3 ctl4 ctl5 ctl6 ctl7 dum vin vdd sample out vss
X0 out.t80 sky130_fd_sc_hd__inv_2_1.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1 out.t81 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X2 out.t82 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 out.t78 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vin.t79 vdd.t138 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X4 vin.t9 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y out.t7 vss.t38 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X5 vss.t121 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y sw_top_1.sky130_fd_sc_hd__inv_4_0.Y vss.t120 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 out.t83 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 vss.t57 sample.t0 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vss.t56 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 vin.t78 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y out.t71 vdd.t137 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X9 vdd.t15 sample.t1 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vdd.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 out.t84 carray_0.unitcap_336.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 out.t85 carray_0.unitcap_151.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 out.t86 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sample.t2 vss.t25 vss.t24 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 out.t87 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 out.t63 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vin.t69 vdd.t120 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X16 out.t19 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y vin.t19 vss.t53 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X17 out.t88 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 out.t89 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 out.t90 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 out.t91 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 out.t92 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 sky130_fd_sc_hd__inv_2_2.Y.t4 ctl7.t0 vdd sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 out.t93 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 out.t94 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 out.t95 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 out.t96 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 vin.t49 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y out.t42 vdd.t79 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X28 vin.t39 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y out.t30 vss.t107 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X29 out.t97 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 out.t98 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 out.t99 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 out.t100 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y sample.t3 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 out.t101 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 out.t102 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 out.t103 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 out.t104 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 out.t105 carray_0.unitcap_47.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 vin.t59 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y out.t53 vdd.t97 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X40 vdd.t140 sample.t4 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vdd.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X41 out.t106 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 vin.t8 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y out.t6 vss.t37 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X43 out.t107 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vss.t129 vss.t128 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X45 out.t108 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 out.t109 carray_0.unitcap_223.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 out.t110 carray_0.unitcap_127.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 out.t111 carray_0.unitcap_16.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 out.t112 sky130_fd_sc_hd__inv_2_2.Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 out.t113 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 out.t68 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vin.t68 vdd.t119 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X52 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vss.t156 vss.t155 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X53 out.t11 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y vin.t18 vss.t52 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X54 vdd.t118 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sw_top_3.sky130_fd_sc_hd__inv_4_0.Y vdd.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X55 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y sample.t5 vdd.t142 vdd.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X56 out.t114 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 out.t115 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 out.t116 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 out.t117 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 vdd ctl2.t0 sky130_fd_sc_hd__inv_2_5.Y.t2 sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X61 vdd ctl5.t0 sky130_fd_sc_hd__inv_2_0.Y.t3 sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X62 vdd.t99 sample.t6 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vdd.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X63 out.t118 carray_0.unitcap_256.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 vdd ctl1.t0 sky130_fd_sc_hd__inv_2_4.Y sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X65 out.t119 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 out.t120 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 out.t121 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 out.t122 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 out.t123 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 vin.t7 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y out.t5 vss.t36 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X71 out.t23 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y vin.t29 vss.t85 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X72 vdd.t55 vss.t182 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X73 out.t124 carray_0.unitcap_0.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 out.t125 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 out.t126 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 out.t127 carray_0.unitcap_328.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X77 out.t128 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 out.t129 carray_0.unitcap_71.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 vdd.t96 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y sw_top_2.sky130_fd_sc_hd__inv_4_0.Y vdd.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X80 out.t130 sky130_fd_sc_hd__inv_2_3.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 out.t131 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 out.t132 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 sky130_fd_sc_hd__inv_2_5.Y.t1 ctl2.t1 vdd sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X84 sky130_fd_sc_hd__inv_2_2.Y.t5 ctl7.t1 vss vss.t41 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X85 out.t133 carray_0.unitcap_167.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 out.t134 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 out.t135 carray_0.unitcap_72.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 vin.t77 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y out.t73 vdd.t136 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X89 out.t136 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 out.t137 carray_0.unitcap_96.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vdd.t116 vdd.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X92 out.t138 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vss.t154 vss.t153 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X94 out.t139 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 vdd.t43 vss.t183 vdd.t42 vdd.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X96 out.t140 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 out.t62 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vin.t67 vdd.t114 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X98 vdd dum.t0 sky130_fd_sc_hd__inv_2_7.Y sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X99 out.t141 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 out.t142 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 out.t143 carray_0.unitcap_152.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 out.t144 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 out.t145 sky130_fd_sc_hd__inv_2_6.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 out.t146 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 out.t147 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 out.t148 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 out.t149 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 out.t40 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vin.t48 vdd.t78 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X109 out.t32 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y vin.t38 vss.t106 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X110 vss dum.t1 sky130_fd_sc_hd__inv_2_7.Y vss.t176 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X111 out.t150 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 out.t151 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 out.t152 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 out.t153 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 sky130_fd_sc_hd__inv_2_6.Y ctl0.t0 vdd sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X116 out.t154 carray_0.unitcap_192.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 vss.t131 sample.t7 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vss.t130 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X118 out.t155 carray_0.unitcap_10.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 out.t156 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 out.t157 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 out.t158 carray_0.unitcap_39.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 vss ctl2.t2 sky130_fd_sc_hd__inv_2_5.Y.t4 vss.t161 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X123 out.t58 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vin.t58 vdd.t94 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X124 out.t159 carray_0.unitcap_224.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 out.t160 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 out.t4 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y vin.t6 vss.t35 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X127 out.t161 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 sky130_fd_sc_hd__inv_2_6.Y ctl0.t1 vss vss.t67 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X129 vss ctl5.t1 sky130_fd_sc_hd__inv_2_0.Y.t4 vss.t179 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X130 vdd.t135 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y sw_top_0.sky130_fd_sc_hd__inv_4_0.Y vdd.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X131 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y sample.t8 vss.t63 vss.t62 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X132 out.t162 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X133 vss ctl1.t1 sky130_fd_sc_hd__inv_2_4.Y vss.t64 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X134 vss.t23 vdd.t146 vss.t22 vss.t21 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X135 vdd.t46 vss.t184 vdd.t45 vdd.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X136 out.t163 carray_0.unitcap_247.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 out.t164 carray_0.unitcap_119.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 vin.t76 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y out.t76 vdd.t133 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X139 out.t165 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 out.t166 sky130_fd_sc_hd__inv_2_3.Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 out.t167 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 out.t168 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X144 vin.t17 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y out.t10 vss.t51 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X145 out.t169 carray_0.unitcap_321.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 out.t170 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 out.t171 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 out.t172 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 sky130_fd_sc_hd__inv_2_5.Y.t3 ctl2.t3 vss vss.t164 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X150 out.t173 carray_0.unitcap_184.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 out.t24 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y vin.t28 vss.t84 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X152 out.t174 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X153 vdd.t77 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y sw_top_1.sky130_fd_sc_hd__inv_4_0.Y vdd.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X154 out.t175 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 out.t176 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 out.t177 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 out.t178 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 out.t179 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 out.t180 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 vss.t20 vdd.t147 vss.t19 vss.t18 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X161 vin.t27 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y out.t29 vss.t83 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X162 vdd.t21 sample.t9 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X163 vss.t59 sample.t10 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vss.t58 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X164 out.t181 carray_0.unitcap_232.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 out.t182 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 out.t183 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X167 out.t184 sky130_fd_sc_hd__inv_2_4.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 out.t185 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 out.t186 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 out.t187 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 out.t3 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y vin.t5 vss.t34 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X172 vin.t75 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y out.t75 vdd.t132 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X173 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y sample.t11 vss.t61 vss.t60 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X174 out.t188 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 out.t189 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 out.t59 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vin.t57 vdd.t93 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X177 out.t190 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 out.t191 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 out.t192 carray_0.unitcap_13.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 out.t193 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 out.t194 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 out.t195 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vss.t127 vss.t126 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X184 vin.t66 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y out.t65 vdd.t111 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X185 out.t196 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 vss.t17 vdd.t148 vss.t16 vss.t15 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X187 out.t197 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 out.t198 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 out.t199 carray_0.unitcap_322.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 out.t200 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 out.t201 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 out.t202 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 out.t203 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 vss.t148 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sw_top_3.sky130_fd_sc_hd__inv_4_0.Y vss.t147 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X195 out.t204 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 out.t205 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 out.t206 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 out.t207 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 vin.t47 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y out.t47 vdd.t75 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X200 vdd ctl3.t0 sky130_fd_sc_hd__inv_2_3.Y.t2 sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X201 vin.t37 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y out.t31 vss.t105 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X202 vdd.t11 sample.t12 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vdd.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X203 out.t208 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 out.t209 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 out.t210 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 out.t211 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 out.t212 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 out.t213 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 out.t214 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 out.t50 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vin.t56 vdd.t92 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X211 out.t215 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X212 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vss.t119 vss.t118 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X213 out.t9 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y vin.t4 vss.t33 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X214 vdd.t91 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y sw_top_2.sky130_fd_sc_hd__inv_4_0.Y vdd.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X215 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sample.t13 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X216 out.t216 carray_0.unitcap_239.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 out.t79 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vin.t74 vdd.t131 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X218 vdd.t49 vss.t185 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X219 out.t217 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 out.t218 sky130_fd_sc_hd__inv_2_5.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 out.t219 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y sample.t14 vss.t91 vss.t90 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X223 out.t220 sky130_fd_sc_hd__inv_2_2.Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X224 out.t221 carray_0.unitcap_95.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X225 out.t15 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y vin.t16 vss.t50 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X226 vdd ctl4.t0 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X227 out.t222 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 out.t223 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 vin.t15 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y out.t14 vss.t49 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X230 out.t224 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 out.t225 carray_0.unitcap_183.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 vss.t152 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y sw_top_0.sky130_fd_sc_hd__inv_4_0.Y vss.t151 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X233 out.t226 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X234 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y sample.t15 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X235 out.t227 sky130_fd_sc_hd__inv_2_7.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 out.t228 carray_0.unitcap_14.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 out.t229 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 out.t230 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 out.t231 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 out.t232 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 out.t233 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 out.t21 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y vin.t26 vss.t82 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X243 sky130_fd_sc_hd__inv_2_0.Y.t1 ctl5.t2 vdd sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X244 out.t234 carray_0.unitcap_56.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 out.t235 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 vdd.t74 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y sw_top_1.sky130_fd_sc_hd__inv_4_0.Y vdd.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X247 sky130_fd_sc_hd__inv_2_4.Y ctl1.t2 vdd sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X248 vin.t25 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y out.t26 vss.t81 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X249 sky130_fd_sc_hd__inv_2_8.Y ctl4.t1 vdd sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X250 out.t236 carray_0.unitcap_326.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 vdd.t17 sample.t16 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vdd.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X252 out.t237 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 out.t238 sky130_fd_sc_hd__inv_2_3.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 out.t239 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 out.t8 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y vin.t3 vss.t32 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X256 vin.t36 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y out.t37 vss.t104 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X257 out.t240 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 vin.t46 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y out.t43 vdd.t72 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X259 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vss.t117 vss.t116 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X260 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sample.t17 vdd.t19 vdd.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X261 out.t241 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 out.t242 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 out.t243 carray_0.unitcap_88.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 out.t244 carray_0.unitcap_136.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 out.t245 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 vdd.t24 vss.t186 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X267 out.t246 carray_0.unitcap_40.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 out.t247 carray_0.unitcap_191.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 out.t72 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vin.t73 vdd.t130 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X270 out.t248 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 out.t249 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 out.t250 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 out.t251 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X274 vin.t55 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y out.t55 vdd.t89 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X275 out.t252 carray_0.unitcap_63.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 vss ctl3.t1 sky130_fd_sc_hd__inv_2_3.Y.t3 vss.t95 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X277 out.t253 carray_0.unitcap_9.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 out.t69 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vin.t65 vdd.t110 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X279 out.t254 carray_0.unitcap_176.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 out.t255 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 vss.t14 vdd.t149 vss.t13 vss.t12 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X282 out.t256 sky130_fd_sc_hd__inv_2_5.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 out.t257 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 out.t258 carray_0.unitcap_80.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 out.t259 carray_0.unitcap_143.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 out.t260 carray_0.unitcap_120.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 vss.t87 sample.t18 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vss.t86 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X288 sky130_fd_sc_hd__inv_2_7.Y dum.t2 vdd sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X289 vin.t35 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y out.t35 vss.t103 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X290 out.t261 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 out.t262 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 out.t263 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 vss ctl4.t2 sky130_fd_sc_hd__inv_2_8.Y vss.t170 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X294 sky130_fd_sc_hd__inv_2_7.Y dum.t3 vss vss.t111 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X295 out.t264 carray_0.unitcap_11.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 vdd.t27 vss.t187 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X297 out.t265 carray_0.unitcap_144.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 out.t266 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vdd.t88 vdd.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X300 out.t267 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 out.t268 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 vin.t45 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y out.t48 vdd.t71 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X303 out.t269 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 out.t270 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 out.t271 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 out.t272 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 out.t273 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 out.t274 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 vin.t54 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y out.t52 vdd.t86 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X310 vin.t2 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y out.t2 vss.t31 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X311 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vdd.t129 vdd.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X312 out.t275 carray_0.unitcap_331.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 out.t276 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 out.t277 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 out.t278 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 sky130_fd_sc_hd__inv_2_0.Y.t2 ctl5.t3 vss vss.t108 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X317 out.t279 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 out.t280 carray_0.unitcap_111.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 out.t281 carray_0.unitcap_200.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 sky130_fd_sc_hd__inv_2_4.Y ctl1.t3 vss vss.t132 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X321 sky130_fd_sc_hd__inv_2_8.Y ctl4.t3 vss vss.t173 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X322 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y sample.t19 vss.t89 vss.t88 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X323 out.t282 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 out.t13 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y vin.t14 vss.t48 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X325 out.t283 carray_0.unitcap_216.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 out.t284 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 out.t285 carray_0.unitcap_175.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 out.t286 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 vdd.t30 vss.t188 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X330 vss.t11 vdd.t150 vss.t10 vss.t9 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X331 out.t287 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 vin.t13 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y out.t12 vss.t47 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X333 vss.t158 sample.t20 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vss.t157 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X334 out.t288 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 out.t289 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 out.t290 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 out.t291 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 out.t292 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 out.t293 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X340 out.t294 carray_0.unitcap_320.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 vin.t44 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y out.t45 vdd.t70 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X342 out.t27 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y vin.t24 vss.t80 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X343 out.t295 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 out.t296 sky130_fd_sc_hd__inv_2_5.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 out.t297 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X346 out.t33 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y vin.t34 vss.t102 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X347 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y sample.t21 vss.t160 vss.t159 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X348 vss.t146 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sw_top_3.sky130_fd_sc_hd__inv_4_0.Y vss.t145 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X349 out.t46 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vin.t43 vdd.t69 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X350 out.t298 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 out.t299 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 out.t300 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X353 vin.t1 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y out.t1 vss.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X354 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vdd.t127 vdd.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X355 out.t301 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 out.t302 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 out.t74 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vin.t72 vdd.t125 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X358 out.t303 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 vss.t40 sample.t22 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vss.t39 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X360 vin.t53 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y out.t56 vdd.t85 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X361 out.t304 carray_0.unitcap_12.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 vss.t8 vdd.t151 vss.t7 vss.t6 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X363 out.t305 sky130_fd_sc_hd__inv_2_0.Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 out.t306 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 out.t307 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 out.t308 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 out.t309 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 out.t310 carray_0.unitcap_55.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X369 out.t311 carray_0.unitcap_23.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 vss.t125 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y sw_top_2.sky130_fd_sc_hd__inv_4_0.Y vss.t124 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X371 out.t64 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vin.t64 vdd.t109 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X372 out.t312 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 out.t313 carray_0.unitcap_337.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 out.t314 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 out.t315 carray_0.unitcap_255.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 out.t316 carray_0.unitcap_135.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 vin.t63 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y out.t61 vdd.t108 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X378 vdd.t52 vss.t189 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X379 vdd.t6 sample.t23 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vdd.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X380 out.t317 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 out.t318 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 out.t319 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 vdd ctl7.t2 sky130_fd_sc_hd__inv_2_2.Y.t0 sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X384 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vss.t144 vss.t143 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X385 vss.t5 vdd.t152 vss.t4 vss.t3 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X386 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y sample.t24 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X387 out.t41 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vin.t42 vdd.t68 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X388 out.t320 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 out.t321 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 out.t34 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y vin.t33 vss.t101 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X391 out.t322 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 out.t323 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 out.t324 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 out.t325 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 out.t326 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 out.t327 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X397 sky130_fd_sc_hd__inv_2_3.Y.t4 ctl3.t2 vdd sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X398 out.t328 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 out.t329 sky130_fd_sc_hd__inv_2_5.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 out.t330 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 vin.t52 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y out.t51 vdd.t84 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X402 out.t331 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 out.t54 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vin.t51 vdd.t83 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X404 out.t332 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 out.t333 carray_0.unitcap_199.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 out.t334 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 out.t335 carray_0.unitcap_31.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 out.t336 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 out.t337 carray_0.unitcap_15.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 vdd ctl6.t0 sky130_fd_sc_hd__inv_2_1.Y.t3 sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X411 out.t338 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X412 out.t339 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 out.t340 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 vdd ctl0.t2 sky130_fd_sc_hd__inv_2_6.Y sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X415 vss.t150 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y sw_top_0.sky130_fd_sc_hd__inv_4_0.Y vss.t149 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X416 vin.t62 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y out.t67 vdd.t107 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X417 vdd.t38 sample.t25 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vdd.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X418 out.t341 carray_0.unitcap_215.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 vin.t12 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y out.t17 vss.t46 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X420 out.t342 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 vin.t23 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y out.t25 vss.t79 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X422 out.t343 carray_0.unitcap_24.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 out.t344 carray_0.unitcap_334.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vss.t142 vss.t141 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X425 out.t345 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y sample.t26 vdd.t102 vdd.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X427 out.t346 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 out.t39 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y vin.t32 vss.t100 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X429 vss.t2 vdd.t153 vss.t1 vss.t0 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X430 out.t347 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 out.t44 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vin.t41 vdd.t67 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X432 out.t348 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 out.t349 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 out.t350 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 out.t351 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 out.t352 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 sky130_fd_sc_hd__inv_2_1.Y.t4 ctl6.t1 vdd sky130_fd_sc_hd__inv_2_7.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X438 out.t353 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 out.t354 carray_0.unitcap_48.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 vss.t115 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y sw_top_1.sky130_fd_sc_hd__inv_4_0.Y vss.t114 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X441 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vdd.t82 vdd.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X442 out.t355 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 vss ctl7.t3 sky130_fd_sc_hd__inv_2_2.Y.t1 vss.t26 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X444 out.t356 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 out.t357 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 out.t358 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 out.t359 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 out.t360 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 out.t361 carray_0.unitcap_79.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X450 vss.t136 sample.t27 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vss.t135 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X451 out.t362 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 out.t363 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 vin.t71 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y out.t77 vdd.t124 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X454 out.t364 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 out.t365 carray_0.unitcap_324.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 vdd.t106 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sw_top_3.sky130_fd_sc_hd__inv_4_0.Y vdd.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X457 out.t366 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 out.t367 carray_0.unitcap_338.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 out.t70 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vin.t70 vdd.t123 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X460 vin.t11 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y out.t16 vss.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X461 out.t368 carray_0.unitcap_104.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 out.t369 carray_0.unitcap_128.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 out.t370 carray_0.unitcap_159.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 sky130_fd_sc_hd__inv_2_3.Y.t5 ctl3.t3 vss vss.t167 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X465 out.t371 carray_0.unitcap_8.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 out.t372 carray_0.unitcap_32.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 out.t373 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 out.t374 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 vin.t61 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y out.t60 vdd.t104 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X470 out.t375 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 out.t38 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y vin.t31 vss.t99 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X472 out.t376 carray_0.unitcap_168.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 vin.t22 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y out.t22 vss.t78 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X474 out.t377 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 out.t378 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X476 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vdd.t66 vdd.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X477 out.t379 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 out.t380 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 out.t381 carray_0.unitcap_64.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 out.t382 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 out.t383 carray_0.unitcap_112.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 out.t384 carray_0.unitcap_208.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 out.t385 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y sample.t28 vdd.t9 vdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X485 out.t49 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vin.t40 vdd.t64 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X486 out.t386 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 vss ctl6.t2 sky130_fd_sc_hd__inv_2_1.Y.t1 vss.t70 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X488 vss ctl0.t3 sky130_fd_sc_hd__inv_2_6.Y vss.t92 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X489 out.t387 carray_0.unitcap_330.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 out.t388 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 out.t0 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y vin.t0 vss.t29 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X492 out.t389 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 out.t390 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 out.t391 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 out.t392 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 vdd.t122 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y sw_top_0.sky130_fd_sc_hd__inv_4_0.Y vdd.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X497 out.t393 carray_0.unitcap_160.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 out.t394 carray_0.unitcap_248.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 out.t395 carray_0.unitcap_288.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 out.t396 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 out.t397 carray_0.unitcap_207.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 out.t398 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 out.t399 carray_0.unitcap_7.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X504 vss.t55 sample.t29 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vss.t54 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X505 out.t57 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vin.t50 vdd.t80 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X506 vin.t60 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y out.t66 vdd.t103 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X507 out.t400 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 sky130_fd_sc_hd__inv_2_1.Y.t2 ctl6.t3 vss vss.t73 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X509 out.t401 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 out.t402 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 out.t403 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 out.t404 carray_0.unitcap_231.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X513 out.t405 carray_0.unitcap_103.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 out.t18 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y vin.t10 vss.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X515 out.t406 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 vss.t123 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y sw_top_2.sky130_fd_sc_hd__inv_4_0.Y vss.t122 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X517 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sample.t30 vss.t138 vss.t137 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X518 out.t407 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 out.t408 carray_0.unitcap_240.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 out.t409 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 vin.t21 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y out.t28 vss.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X522 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X523 vin.t30 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y out.t36 vss.t98 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X524 out.t410 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 out.t411 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 out.t20 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y vin.t20 vss.t76 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X527 out.t412 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 out.t413 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y sample.t31 vss.t140 vss.t139 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X530 out.t414 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 out.t415 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 out.t416 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 out.t417 sky130_fd_sc_hd__inv_2_4.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X534 out.t418 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 out.t419 carray_0.unitcap_87.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 out.n426 out.t52 28.5655
R1 out.n426 out.t57 28.5655
R2 out.n429 out.t56 28.5655
R3 out.n429 out.t58 28.5655
R4 out.n424 out.t51 28.5655
R5 out.n424 out.t59 28.5655
R6 out.n423 out.t53 28.5655
R7 out.n423 out.t50 28.5655
R8 out.n418 out.t55 28.5655
R9 out.n418 out.t54 28.5655
R10 out.n58 out.t66 28.5655
R11 out.n58 out.t69 28.5655
R12 out.n61 out.t65 28.5655
R13 out.n61 out.t64 28.5655
R14 out.n56 out.t61 28.5655
R15 out.n56 out.t63 28.5655
R16 out.n55 out.t67 28.5655
R17 out.n55 out.t68 28.5655
R18 out.n50 out.t60 28.5655
R19 out.n50 out.t62 28.5655
R20 out.n34 out.t45 28.5655
R21 out.n34 out.t40 28.5655
R22 out.n37 out.t42 28.5655
R23 out.n37 out.t46 28.5655
R24 out.n32 out.t47 28.5655
R25 out.n32 out.t41 28.5655
R26 out.n31 out.t43 28.5655
R27 out.n31 out.t44 28.5655
R28 out.n26 out.t48 28.5655
R29 out.n26 out.t49 28.5655
R30 out.n10 out.t75 28.5655
R31 out.n10 out.t74 28.5655
R32 out.n13 out.t71 28.5655
R33 out.n13 out.t78 28.5655
R34 out.n8 out.t77 28.5655
R35 out.n8 out.t79 28.5655
R36 out.n7 out.t73 28.5655
R37 out.n7 out.t72 28.5655
R38 out.n2 out.t76 28.5655
R39 out.n2 out.t70 28.5655
R40 out.n427 out.t25 17.4005
R41 out.n427 out.t23 17.4005
R42 out.n431 out.t22 17.4005
R43 out.n431 out.t21 17.4005
R44 out.n425 out.t28 17.4005
R45 out.n425 out.t24 17.4005
R46 out.n434 out.t29 17.4005
R47 out.n434 out.t27 17.4005
R48 out.n437 out.t26 17.4005
R49 out.n437 out.t20 17.4005
R50 out.n59 out.t5 17.4005
R51 out.n59 out.t8 17.4005
R52 out.n63 out.t2 17.4005
R53 out.n63 out.t0 17.4005
R54 out.n57 out.t1 17.4005
R55 out.n57 out.t4 17.4005
R56 out.n66 out.t7 17.4005
R57 out.n66 out.t3 17.4005
R58 out.n69 out.t6 17.4005
R59 out.n69 out.t9 17.4005
R60 out.n35 out.t16 17.4005
R61 out.n35 out.t15 17.4005
R62 out.n39 out.t10 17.4005
R63 out.n39 out.t13 17.4005
R64 out.n33 out.t12 17.4005
R65 out.n33 out.t18 17.4005
R66 out.n42 out.t14 17.4005
R67 out.n42 out.t19 17.4005
R68 out.n45 out.t17 17.4005
R69 out.n45 out.t11 17.4005
R70 out.n11 out.t35 17.4005
R71 out.n11 out.t38 17.4005
R72 out.n15 out.t36 17.4005
R73 out.n15 out.t32 17.4005
R74 out.n9 out.t30 17.4005
R75 out.n9 out.t33 17.4005
R76 out.n18 out.t31 17.4005
R77 out.n18 out.t34 17.4005
R78 out.n21 out.t37 17.4005
R79 out.n21 out.t39 17.4005
R80 out.n421 out.n420 9.05098
R81 out.n53 out.n52 9.05098
R82 out.n29 out.n28 9.05098
R83 out.n5 out.n4 9.05098
R84 out.n420 out.n419 9.0005
R85 out.n422 out.n421 9.0005
R86 out.n52 out.n51 9.0005
R87 out.n54 out.n53 9.0005
R88 out.n28 out.n27 9.0005
R89 out.n30 out.n29 9.0005
R90 out.n4 out.n3 9.0005
R91 out.n6 out.n5 9.0005
R92 out.n444 out.n443 8.6431
R93 out.n443 out.n442 6.19787
R94 out.n417 out.n416 4.5786
R95 out.n49 out.n48 4.5786
R96 out.n25 out.n24 4.5786
R97 out.n1 out.n0 4.5786
R98 out.n442 out.n441 4.3755
R99 out.n436 out.n423 2.5289
R100 out.n68 out.n55 2.5289
R101 out.n44 out.n31 2.5289
R102 out.n20 out.n7 2.5289
R103 out.n430 out.n429 2.52132
R104 out.n62 out.n61 2.52132
R105 out.n38 out.n37 2.52132
R106 out.n14 out.n13 2.52132
R107 out.n440 out 2.47089
R108 out.n433 out.n424 2.45817
R109 out.n65 out.n56 2.45817
R110 out.n41 out.n32 2.45817
R111 out.n17 out.n8 2.45817
R112 out.n428 out.n426 2.45375
R113 out.n60 out.n58 2.4534
R114 out.n36 out.n34 2.4534
R115 out.n12 out.n10 2.4534
R116 out.n442 out 2.42846
R117 out.n443 out 2.29984
R118 out.n441 out.n440 1.90839
R119 out out.n439 1.05971
R120 out out.n47 1.05971
R121 out out.n23 1.05971
R122 out out.n71 1.05955
R123 out.n435 out.n434 0.750533
R124 out.n67 out.n66 0.750533
R125 out.n43 out.n42 0.750533
R126 out.n19 out.n18 0.750533
R127 out.n438 out.n437 0.747922
R128 out.n70 out.n69 0.747922
R129 out.n46 out.n45 0.747922
R130 out.n22 out.n21 0.747922
R131 out.n433 out.n425 0.729365
R132 out.n65 out.n57 0.729365
R133 out.n41 out.n33 0.729365
R134 out.n17 out.n9 0.729365
R135 out.n432 out.n431 0.725192
R136 out.n64 out.n63 0.725192
R137 out.n40 out.n39 0.725192
R138 out.n16 out.n15 0.725192
R139 out.n435 out.n433 0.720895
R140 out.n67 out.n65 0.720895
R141 out.n43 out.n41 0.720895
R142 out.n19 out.n17 0.720895
R143 out.n433 out.n432 0.714316
R144 out.n65 out.n64 0.714316
R145 out.n41 out.n40 0.714316
R146 out.n17 out.n16 0.714316
R147 out.n430 out.n428 0.704447
R148 out.n62 out.n60 0.704447
R149 out.n38 out.n36 0.704447
R150 out.n14 out.n12 0.704447
R151 out.n428 out.n427 0.66743
R152 out.n60 out.n59 0.66743
R153 out.n36 out.n35 0.66743
R154 out.n12 out.n11 0.66743
R155 out.n438 out.n436 0.645237
R156 out.n70 out.n68 0.645237
R157 out.n46 out.n44 0.645237
R158 out.n22 out.n20 0.645237
R159 out.n439 out.n422 0.57857
R160 out.n71 out.n54 0.57857
R161 out.n47 out.n30 0.57857
R162 out.n23 out.n6 0.57857
R163 out.n441 out.n415 0.438625
R164 out.n101 out 0.400915
R165 out.n102 out 0.400915
R166 out.n103 out 0.400915
R167 out.n104 out 0.400915
R168 out.n105 out 0.400915
R169 out.n106 out 0.400915
R170 out.n107 out 0.400915
R171 out.n108 out 0.400915
R172 out.n109 out 0.400915
R173 out.n110 out 0.400915
R174 out.n111 out 0.400915
R175 out.n112 out 0.400915
R176 out.n113 out 0.400915
R177 out.n114 out 0.400915
R178 out.n115 out 0.400915
R179 out.n116 out 0.400915
R180 out.n117 out 0.400915
R181 out.n118 out 0.400915
R182 out.n119 out 0.400915
R183 out.n120 out 0.400915
R184 out.n121 out 0.400915
R185 out.n122 out 0.400915
R186 out.n123 out 0.400915
R187 out.n124 out 0.400915
R188 out.n125 out 0.400915
R189 out.n126 out 0.400915
R190 out.n127 out 0.400915
R191 out.n128 out 0.400915
R192 out.n129 out 0.400915
R193 out.n130 out 0.400915
R194 out.n131 out 0.400915
R195 out.n132 out 0.400915
R196 out.n133 out 0.400915
R197 out.n134 out 0.400915
R198 out.n135 out 0.400915
R199 out.n136 out 0.400915
R200 out.n137 out 0.400915
R201 out.n138 out 0.400915
R202 out.n139 out 0.400915
R203 out.n140 out 0.400915
R204 out.n141 out 0.400915
R205 out.n142 out 0.400915
R206 out.n143 out 0.400915
R207 out.n144 out 0.400915
R208 out.n145 out 0.400915
R209 out.n146 out 0.400915
R210 out.n147 out 0.400915
R211 out.n148 out 0.400915
R212 out.n149 out 0.400915
R213 out.n150 out 0.400915
R214 out.n151 out 0.400915
R215 out.n152 out 0.400915
R216 out.n153 out 0.400915
R217 out.n154 out 0.400915
R218 out.n155 out 0.400915
R219 out.n156 out 0.400915
R220 out.n157 out 0.400915
R221 out.n158 out 0.400915
R222 out.n159 out 0.400915
R223 out.n160 out 0.400915
R224 out.n161 out 0.400915
R225 out.n162 out 0.400915
R226 out.n163 out 0.400915
R227 out.n164 out 0.400915
R228 out.n165 out 0.400915
R229 out.n166 out 0.400915
R230 out.n167 out 0.400915
R231 out.n168 out 0.400915
R232 out.n169 out 0.400915
R233 out.n170 out 0.400915
R234 out.n171 out 0.400915
R235 out.n172 out 0.400915
R236 out.n173 out 0.400915
R237 out.n174 out 0.400915
R238 out.n175 out 0.400915
R239 out.n176 out 0.400915
R240 out.n177 out 0.400915
R241 out.n178 out 0.400915
R242 out.n179 out 0.400915
R243 out.n180 out 0.400915
R244 out.n181 out 0.400915
R245 out.n182 out 0.400915
R246 out.n183 out 0.400915
R247 out.n184 out 0.400915
R248 out.n185 out 0.400915
R249 out.n186 out 0.400915
R250 out.n187 out 0.400915
R251 out.n188 out 0.400915
R252 out.n189 out 0.400915
R253 out.n190 out 0.400915
R254 out.n191 out 0.400915
R255 out.n192 out 0.400915
R256 out.n193 out 0.400915
R257 out.n194 out 0.400915
R258 out.n195 out 0.400915
R259 out.n196 out 0.400915
R260 out.n197 out 0.400915
R261 out.n198 out 0.400915
R262 out.n199 out 0.400915
R263 out.n200 out 0.400915
R264 out.n201 out 0.400915
R265 out.n202 out 0.400915
R266 out.n203 out 0.400915
R267 out.n204 out 0.400915
R268 out.n205 out 0.400915
R269 out.n206 out 0.400915
R270 out.n207 out 0.400915
R271 out.n208 out 0.400915
R272 out.n209 out 0.400915
R273 out.n210 out 0.400915
R274 out.n211 out 0.400915
R275 out.n212 out 0.400915
R276 out.n213 out 0.400915
R277 out.n214 out 0.400915
R278 out.n215 out 0.400915
R279 out.n216 out 0.400915
R280 out.n217 out 0.400915
R281 out.n218 out 0.400915
R282 out.n219 out 0.400915
R283 out.n220 out 0.400915
R284 out.n221 out 0.400915
R285 out.n222 out 0.400915
R286 out.n223 out 0.400915
R287 out.n224 out 0.400915
R288 out.n225 out 0.400915
R289 out.n226 out 0.400915
R290 out.n227 out 0.400915
R291 out.n228 out 0.400915
R292 out.n229 out 0.400915
R293 out.n230 out 0.400915
R294 out.n231 out 0.400915
R295 out.n232 out 0.400915
R296 out.n233 out 0.400915
R297 out.n234 out 0.400915
R298 out.n235 out 0.400915
R299 out.n236 out 0.400915
R300 out.n237 out 0.400915
R301 out.n238 out 0.400915
R302 out.n239 out 0.400915
R303 out.n240 out 0.400915
R304 out.n241 out 0.400915
R305 out.n242 out 0.400915
R306 out.n243 out 0.400915
R307 out.n244 out 0.400915
R308 out.n245 out 0.400915
R309 out.n246 out 0.400915
R310 out.n247 out 0.400915
R311 out.n248 out 0.400915
R312 out.n249 out 0.400915
R313 out.n250 out 0.400915
R314 out.n251 out 0.400915
R315 out.n252 out 0.400915
R316 out.n253 out 0.400915
R317 out.n254 out 0.400915
R318 out.n255 out 0.400915
R319 out.n256 out 0.400915
R320 out.n257 out 0.400915
R321 out.n258 out 0.400915
R322 out.n259 out 0.400915
R323 out.n260 out 0.400915
R324 out.n261 out 0.400915
R325 out.n262 out 0.400915
R326 out.n263 out 0.400915
R327 out.n264 out 0.400915
R328 out.n265 out 0.400915
R329 out.n266 out 0.400915
R330 out.n267 out 0.400915
R331 out.n268 out 0.400915
R332 out.n269 out 0.400915
R333 out.n270 out 0.400915
R334 out.n271 out 0.400915
R335 out.n272 out 0.400915
R336 out.n273 out 0.400915
R337 out.n274 out 0.400915
R338 out.n275 out 0.400915
R339 out.n276 out 0.400915
R340 out.n277 out 0.400915
R341 out.n278 out 0.400915
R342 out.n279 out 0.400915
R343 out.n280 out 0.400915
R344 out.n281 out 0.400915
R345 out.n282 out 0.400915
R346 out.n283 out 0.400915
R347 out.n284 out 0.400915
R348 out.n285 out 0.400915
R349 out.n286 out 0.400915
R350 out.n287 out 0.400915
R351 out.n288 out 0.400915
R352 out.n289 out 0.400915
R353 out.n290 out 0.400915
R354 out.n291 out 0.400915
R355 out.n292 out 0.400915
R356 out.n293 out 0.400915
R357 out.n294 out 0.400915
R358 out.n295 out 0.400915
R359 out.n296 out 0.400915
R360 out.n297 out 0.400915
R361 out.n298 out 0.400915
R362 out.n299 out 0.400915
R363 out.n300 out 0.400915
R364 out.n301 out 0.400915
R365 out.n302 out 0.400915
R366 out.n303 out 0.400915
R367 out.n304 out 0.400915
R368 out.n305 out 0.400915
R369 out.n306 out 0.400915
R370 out.n307 out 0.400915
R371 out.n308 out 0.400915
R372 out.n309 out 0.400915
R373 out.n310 out 0.400915
R374 out.n311 out 0.400915
R375 out.n312 out 0.400915
R376 out.n313 out 0.400915
R377 out.n314 out 0.400915
R378 out.n315 out 0.400915
R379 out.n316 out 0.400915
R380 out.n317 out 0.400915
R381 out out.n323 0.400915
R382 out out.n324 0.400915
R383 out out.n325 0.400915
R384 out out.n326 0.400915
R385 out out.n327 0.400915
R386 out out.n328 0.400915
R387 out out.n329 0.400915
R388 out out.n330 0.400915
R389 out out.n331 0.400915
R390 out out.n332 0.400915
R391 out out.n333 0.400915
R392 out out.n334 0.400915
R393 out out.n335 0.400915
R394 out out.n336 0.400915
R395 out out.n337 0.400915
R396 out out.n338 0.400915
R397 out out.n339 0.400915
R398 out out.n340 0.400915
R399 out out.n341 0.400915
R400 out out.n342 0.400915
R401 out out.n343 0.400915
R402 out out.n344 0.400915
R403 out out.n345 0.400915
R404 out out.n346 0.400915
R405 out out.n347 0.400915
R406 out out.n348 0.400915
R407 out out.n349 0.400915
R408 out out.n350 0.400915
R409 out out.n351 0.400915
R410 out out.n352 0.400915
R411 out out.n353 0.400915
R412 out out.n354 0.400915
R413 out out.n355 0.400915
R414 out.n368 out 0.400915
R415 out.n369 out 0.400915
R416 out.n370 out 0.400915
R417 out.n371 out 0.400915
R418 out.n372 out 0.400915
R419 out.n373 out 0.400915
R420 out.n374 out 0.400915
R421 out.n375 out 0.400915
R422 out.n376 out 0.400915
R423 out.n377 out 0.400915
R424 out.n378 out 0.400915
R425 out.n379 out 0.400915
R426 out.n380 out 0.400915
R427 out.n381 out 0.400915
R428 out.n382 out 0.400915
R429 out.n383 out 0.400915
R430 out.n384 out 0.400915
R431 out.n385 out 0.400915
R432 out.n386 out 0.400915
R433 out.n387 out 0.400915
R434 out.n388 out 0.400915
R435 out.n389 out 0.400915
R436 out.n390 out 0.400915
R437 out.n391 out 0.400915
R438 out.n392 out 0.400915
R439 out.n393 out 0.400915
R440 out.n394 out 0.400915
R441 out.n395 out 0.400915
R442 out.n396 out 0.400915
R443 out.n397 out 0.400915
R444 out.n398 out 0.400915
R445 out.n399 out 0.400915
R446 out out.n412 0.400915
R447 out out.n413 0.400915
R448 out.n72 out 0.400915
R449 out.n73 out 0.400915
R450 out.n74 out 0.400915
R451 out.n75 out 0.400915
R452 out.n76 out 0.400915
R453 out.n77 out 0.400915
R454 out.n78 out 0.400915
R455 out.n79 out 0.400915
R456 out.n80 out 0.400915
R457 out.n81 out 0.400915
R458 out.n82 out 0.400915
R459 out.n83 out 0.400915
R460 out.n84 out 0.400915
R461 out.n85 out 0.400915
R462 out.n86 out 0.400915
R463 out.n87 out 0.400915
R464 out.n88 out 0.400915
R465 out.n89 out 0.400915
R466 out.n90 out 0.400915
R467 out.n91 out 0.400915
R468 out.n92 out 0.400915
R469 out.n93 out 0.400915
R470 out.n94 out 0.400915
R471 out.n95 out 0.400915
R472 out.n96 out 0.400915
R473 out.n97 out 0.400915
R474 out.n98 out 0.400915
R475 out.n99 out 0.400915
R476 out.n367 out.n366 0.398433
R477 out.n409 out 0.377415
R478 out.n407 out 0.377415
R479 out.n405 out 0.377415
R480 out.n403 out 0.377415
R481 out.n401 out 0.377415
R482 out.n320 out 0.377415
R483 out.n318 out 0.377415
R484 out out.n411 0.377415
R485 out out.n100 0.250087
R486 out out.n319 0.250087
R487 out.n358 out 0.250087
R488 out.n359 out 0.250087
R489 out.n360 out 0.250087
R490 out.n361 out 0.250087
R491 out.n362 out 0.250087
R492 out.n363 out 0.250087
R493 out.n364 out 0.250087
R494 out.n365 out 0.250087
R495 out out.n402 0.250087
R496 out out.n404 0.250087
R497 out out.n406 0.250087
R498 out out.n408 0.250087
R499 out out.n410 0.250087
R500 out.n357 out.n356 0.243372
R501 out.n322 out.n321 0.241767
R502 out out.n400 0.226587
R503 out.n415 out.n414 0.21905
R504 out.n415 out 0.182365
R505 out.n419 out.n418 0.100193
R506 out.n51 out.n50 0.100193
R507 out.n27 out.n26 0.100193
R508 out.n3 out.n2 0.100193
R509 out.n440 out 0.063
R510 out.n420 out.n416 0.0421667
R511 out.n52 out.n48 0.0421667
R512 out.n28 out.n24 0.0421667
R513 out.n4 out.n0 0.0421667
R514 out.n422 out.n416 0.0310556
R515 out.n54 out.n48 0.0310556
R516 out.n30 out.n24 0.0310556
R517 out.n6 out.n0 0.0310556
R518 out out.t296 0.0215188
R519 out out.t184 0.0215188
R520 out out.t417 0.0215188
R521 out out.t145 0.0215188
R522 out out.t227 0.0215188
R523 out out.t256 0.0215188
R524 out out.t329 0.0215188
R525 out out.t218 0.0215188
R526 out out.n101 0.0215186
R527 out out.n102 0.0215186
R528 out out.n103 0.0215186
R529 out out.n104 0.0215186
R530 out out.n105 0.0215186
R531 out out.n106 0.0215186
R532 out out.n107 0.0215186
R533 out out.n108 0.0215186
R534 out out.n109 0.0215186
R535 out out.n110 0.0215186
R536 out out.n111 0.0215186
R537 out out.n112 0.0215186
R538 out out.n113 0.0215186
R539 out out.n114 0.0215186
R540 out out.n115 0.0215186
R541 out out.n116 0.0215186
R542 out out.n117 0.0215186
R543 out out.n118 0.0215186
R544 out out.n119 0.0215186
R545 out out.n120 0.0215186
R546 out out.n121 0.0215186
R547 out out.n122 0.0215186
R548 out out.n123 0.0215186
R549 out out.n124 0.0215186
R550 out out.n125 0.0215186
R551 out out.n126 0.0215186
R552 out out.n127 0.0215186
R553 out out.n128 0.0215186
R554 out out.n129 0.0215186
R555 out out.n130 0.0215186
R556 out out.n131 0.0215186
R557 out out.n132 0.0215186
R558 out out.n133 0.0215186
R559 out out.n134 0.0215186
R560 out out.n135 0.0215186
R561 out out.n136 0.0215186
R562 out out.n137 0.0215186
R563 out out.n138 0.0215186
R564 out out.n139 0.0215186
R565 out out.n140 0.0215186
R566 out out.n141 0.0215186
R567 out out.n142 0.0215186
R568 out out.n143 0.0215186
R569 out out.n144 0.0215186
R570 out out.n145 0.0215186
R571 out out.n146 0.0215186
R572 out out.n147 0.0215186
R573 out out.n148 0.0215186
R574 out out.n149 0.0215186
R575 out out.n150 0.0215186
R576 out out.n151 0.0215186
R577 out out.n152 0.0215186
R578 out out.n153 0.0215186
R579 out out.n154 0.0215186
R580 out out.n155 0.0215186
R581 out out.n156 0.0215186
R582 out out.n157 0.0215186
R583 out out.n158 0.0215186
R584 out out.n159 0.0215186
R585 out out.n160 0.0215186
R586 out out.n161 0.0215186
R587 out out.n162 0.0215186
R588 out out.n163 0.0215186
R589 out out.n164 0.0215186
R590 out out.n165 0.0215186
R591 out out.n166 0.0215186
R592 out out.n167 0.0215186
R593 out out.n168 0.0215186
R594 out out.n169 0.0215186
R595 out out.n170 0.0215186
R596 out out.n171 0.0215186
R597 out out.n172 0.0215186
R598 out out.n173 0.0215186
R599 out out.n174 0.0215186
R600 out out.n175 0.0215186
R601 out out.n176 0.0215186
R602 out out.n177 0.0215186
R603 out out.n178 0.0215186
R604 out out.n179 0.0215186
R605 out out.n180 0.0215186
R606 out out.n181 0.0215186
R607 out out.n182 0.0215186
R608 out out.n183 0.0215186
R609 out out.n184 0.0215186
R610 out out.n185 0.0215186
R611 out out.n186 0.0215186
R612 out out.n187 0.0215186
R613 out out.n188 0.0215186
R614 out out.n189 0.0215186
R615 out out.n190 0.0215186
R616 out out.n191 0.0215186
R617 out out.n192 0.0215186
R618 out out.n193 0.0215186
R619 out out.n194 0.0215186
R620 out out.n195 0.0215186
R621 out out.n196 0.0215186
R622 out out.n197 0.0215186
R623 out out.n198 0.0215186
R624 out out.n199 0.0215186
R625 out out.n200 0.0215186
R626 out out.n201 0.0215186
R627 out out.n202 0.0215186
R628 out out.n203 0.0215186
R629 out out.n204 0.0215186
R630 out out.n205 0.0215186
R631 out out.n206 0.0215186
R632 out out.n207 0.0215186
R633 out out.n208 0.0215186
R634 out out.n209 0.0215186
R635 out out.n210 0.0215186
R636 out out.n211 0.0215186
R637 out out.n212 0.0215186
R638 out out.n213 0.0215186
R639 out out.n214 0.0215186
R640 out out.n215 0.0215186
R641 out out.n216 0.0215186
R642 out out.n217 0.0215186
R643 out out.n218 0.0215186
R644 out out.n219 0.0215186
R645 out out.n220 0.0215186
R646 out out.n221 0.0215186
R647 out out.n222 0.0215186
R648 out out.n223 0.0215186
R649 out out.n224 0.0215186
R650 out out.n225 0.0215186
R651 out out.n226 0.0215186
R652 out out.n227 0.0215186
R653 out out.n228 0.0215186
R654 out out.n229 0.0215186
R655 out out.n230 0.0215186
R656 out out.n231 0.0215186
R657 out out.n232 0.0215186
R658 out out.n233 0.0215186
R659 out out.n234 0.0215186
R660 out out.n235 0.0215186
R661 out out.n236 0.0215186
R662 out out.n237 0.0215186
R663 out out.n238 0.0215186
R664 out out.n239 0.0215186
R665 out out.n240 0.0215186
R666 out out.n241 0.0215186
R667 out out.n242 0.0215186
R668 out out.n243 0.0215186
R669 out out.n244 0.0215186
R670 out out.n245 0.0215186
R671 out out.n246 0.0215186
R672 out out.n247 0.0215186
R673 out out.n248 0.0215186
R674 out out.n249 0.0215186
R675 out out.n250 0.0215186
R676 out out.n251 0.0215186
R677 out out.n252 0.0215186
R678 out out.n253 0.0215186
R679 out out.n254 0.0215186
R680 out out.n255 0.0215186
R681 out out.n256 0.0215186
R682 out out.n257 0.0215186
R683 out out.n258 0.0215186
R684 out out.n259 0.0215186
R685 out out.n260 0.0215186
R686 out out.n261 0.0215186
R687 out out.n262 0.0215186
R688 out out.n263 0.0215186
R689 out out.n264 0.0215186
R690 out out.n265 0.0215186
R691 out out.n266 0.0215186
R692 out out.n267 0.0215186
R693 out out.n268 0.0215186
R694 out out.n269 0.0215186
R695 out out.n270 0.0215186
R696 out out.n271 0.0215186
R697 out out.n272 0.0215186
R698 out out.n273 0.0215186
R699 out out.n274 0.0215186
R700 out out.n275 0.0215186
R701 out out.n276 0.0215186
R702 out out.n277 0.0215186
R703 out out.n278 0.0215186
R704 out out.n279 0.0215186
R705 out out.n280 0.0215186
R706 out out.n281 0.0215186
R707 out out.n282 0.0215186
R708 out out.n283 0.0215186
R709 out out.n284 0.0215186
R710 out out.n285 0.0215186
R711 out out.n286 0.0215186
R712 out out.n287 0.0215186
R713 out out.n288 0.0215186
R714 out out.n289 0.0215186
R715 out out.n290 0.0215186
R716 out out.n291 0.0215186
R717 out out.n292 0.0215186
R718 out out.n293 0.0215186
R719 out out.n294 0.0215186
R720 out out.n295 0.0215186
R721 out out.n296 0.0215186
R722 out out.n297 0.0215186
R723 out out.n298 0.0215186
R724 out out.n299 0.0215186
R725 out out.n300 0.0215186
R726 out out.n301 0.0215186
R727 out out.n302 0.0215186
R728 out out.n303 0.0215186
R729 out out.n304 0.0215186
R730 out out.n305 0.0215186
R731 out out.n306 0.0215186
R732 out out.n307 0.0215186
R733 out out.n308 0.0215186
R734 out out.n309 0.0215186
R735 out out.n310 0.0215186
R736 out out.n311 0.0215186
R737 out out.n312 0.0215186
R738 out out.n313 0.0215186
R739 out out.n314 0.0215186
R740 out out.n315 0.0215186
R741 out out.n316 0.0215186
R742 out out.n317 0.0215186
R743 out.n324 out 0.0215186
R744 out.n325 out 0.0215186
R745 out.n326 out 0.0215186
R746 out.n327 out 0.0215186
R747 out.n328 out 0.0215186
R748 out.n329 out 0.0215186
R749 out.n330 out 0.0215186
R750 out.n331 out 0.0215186
R751 out.n332 out 0.0215186
R752 out.n333 out 0.0215186
R753 out.n334 out 0.0215186
R754 out.n335 out 0.0215186
R755 out.n336 out 0.0215186
R756 out.n337 out 0.0215186
R757 out.n338 out 0.0215186
R758 out.n339 out 0.0215186
R759 out.n340 out 0.0215186
R760 out.n341 out 0.0215186
R761 out.n342 out 0.0215186
R762 out.n343 out 0.0215186
R763 out.n344 out 0.0215186
R764 out.n345 out 0.0215186
R765 out.n346 out 0.0215186
R766 out.n347 out 0.0215186
R767 out.n348 out 0.0215186
R768 out.n349 out 0.0215186
R769 out.n350 out 0.0215186
R770 out.n351 out 0.0215186
R771 out.n352 out 0.0215186
R772 out.n353 out 0.0215186
R773 out.n354 out 0.0215186
R774 out.n355 out 0.0215186
R775 out.n356 out 0.0215186
R776 out out.n367 0.0215186
R777 out out.n368 0.0215186
R778 out out.n369 0.0215186
R779 out out.n370 0.0215186
R780 out out.n371 0.0215186
R781 out out.n372 0.0215186
R782 out out.n373 0.0215186
R783 out out.n374 0.0215186
R784 out out.n375 0.0215186
R785 out out.n376 0.0215186
R786 out out.n377 0.0215186
R787 out out.n378 0.0215186
R788 out out.n379 0.0215186
R789 out out.n380 0.0215186
R790 out out.n381 0.0215186
R791 out out.n382 0.0215186
R792 out out.n383 0.0215186
R793 out out.n384 0.0215186
R794 out out.n385 0.0215186
R795 out out.n386 0.0215186
R796 out out.n387 0.0215186
R797 out out.n388 0.0215186
R798 out out.n389 0.0215186
R799 out out.n390 0.0215186
R800 out out.n391 0.0215186
R801 out out.n392 0.0215186
R802 out out.n393 0.0215186
R803 out out.n394 0.0215186
R804 out out.n395 0.0215186
R805 out out.n396 0.0215186
R806 out out.n397 0.0215186
R807 out out.n398 0.0215186
R808 out.n412 out 0.0215186
R809 out.n413 out 0.0215186
R810 out.n414 out 0.0215186
R811 out out.n72 0.0215186
R812 out out.n73 0.0215186
R813 out out.n74 0.0215186
R814 out out.n75 0.0215186
R815 out out.n76 0.0215186
R816 out out.n77 0.0215186
R817 out out.n78 0.0215186
R818 out out.n79 0.0215186
R819 out out.n80 0.0215186
R820 out out.n81 0.0215186
R821 out out.n82 0.0215186
R822 out out.n83 0.0215186
R823 out out.n84 0.0215186
R824 out out.n85 0.0215186
R825 out out.n86 0.0215186
R826 out out.n87 0.0215186
R827 out out.n88 0.0215186
R828 out out.n89 0.0215186
R829 out out.n90 0.0215186
R830 out out.n91 0.0215186
R831 out out.n92 0.0215186
R832 out out.n93 0.0215186
R833 out out.n94 0.0215186
R834 out out.n95 0.0215186
R835 out out.n96 0.0215186
R836 out out.n97 0.0215186
R837 out out.n98 0.0215186
R838 out out.n99 0.0215186
R839 out.n322 out 0.0193292
R840 out.n400 out 0.0193292
R841 out.n444 out 0.0169474
R842 out out.n444 0.016125
R843 out out.n357 0.0156801
R844 out out.n358 0.0156801
R845 out out.n359 0.0156801
R846 out out.n360 0.0156801
R847 out out.n361 0.0156801
R848 out out.n362 0.0156801
R849 out out.n363 0.0156801
R850 out out.n364 0.0156801
R851 out.n366 out 0.0150963
R852 out.n319 out.n318 0.0139286
R853 out.n408 out.n407 0.012177
R854 out.n410 out.n409 0.012177
R855 out.n321 out.n320 0.0118851
R856 out.n402 out.n401 0.0110093
R857 out.n404 out.n403 0.0110093
R858 out.n406 out.n405 0.00954969
R859 out.n411 out.n100 0.00925776
R860 out.n432 out.n430 0.00707895
R861 out.n436 out.n435 0.00707895
R862 out.n439 out.n438 0.00707895
R863 out.n64 out.n62 0.00707895
R864 out.n68 out.n67 0.00707895
R865 out.n71 out.n70 0.00707895
R866 out.n40 out.n38 0.00707895
R867 out.n44 out.n43 0.00707895
R868 out.n47 out.n46 0.00707895
R869 out.n16 out.n14 0.00707895
R870 out.n20 out.n19 0.00707895
R871 out.n23 out.n22 0.00707895
R872 out.n411 out 0.00692236
R873 out.n405 out 0.00663044
R874 out.n401 out 0.00517081
R875 out.n403 out 0.00517081
R876 out.n320 out 0.00429503
R877 out.n407 out 0.00400311
R878 out.n409 out 0.00400311
R879 out.n323 out.n322 0.00268944
R880 out.n400 out.n399 0.00268944
R881 out.n318 out 0.00225155
R882 out.n419 out.n417 0.00222265
R883 out.n51 out.n49 0.00222265
R884 out.n27 out.n25 0.00222265
R885 out.n3 out.n1 0.00222265
R886 out.n421 out.n417 0.00218088
R887 out.n53 out.n49 0.00218088
R888 out.n29 out.n25 0.00218088
R889 out.n5 out.n1 0.00218088
R890 out.n366 out.n365 0.00108385
R891 out.n101 out.t238 0.000500141
R892 out.n102 out.t141 0.000500141
R893 out.n103 out.t90 0.000500141
R894 out.n104 out.t378 0.000500141
R895 out.n105 out.t322 0.000500141
R896 out.n106 out.t269 0.000500141
R897 out.n107 out.t175 0.000500141
R898 out.n108 out.t317 0.000500141
R899 out.n109 out.t261 0.000500141
R900 out.n110 out.t207 0.000500141
R901 out.n111 out.t152 0.000500141
R902 out.n112 out.t407 0.000500141
R903 out.n113 out.t345 0.000500141
R904 out.n114 out.t297 0.000500141
R905 out.n115 out.t239 0.000500141
R906 out.n116 out.t186 0.000500141
R907 out.n117 out.t91 0.000500141
R908 out.n118 out.t379 0.000500141
R909 out.n119 out.t323 0.000500141
R910 out.n120 out.t201 0.000500141
R911 out.n121 out.t147 0.000500141
R912 out.n122 out.t401 0.000500141
R913 out.n123 out.t338 0.000500141
R914 out.n124 out.t292 0.000500141
R915 out.n125 out.t232 0.000500141
R916 out.n126 out.t180 0.000500141
R917 out.n127 out.t87 0.000500141
R918 out.n128 out.t374 0.000500141
R919 out.n129 out.t319 0.000500141
R920 out.n130 out.t263 0.000500141
R921 out.n131 out.t235 0.000500141
R922 out.n132 out.t130 0.000500141
R923 out.n133 out.t377 0.000500141
R924 out.n134 out.t320 0.000500141
R925 out.n135 out.t267 0.000500141
R926 out.n136 out.t211 0.000500141
R927 out.n137 out.t160 0.000500141
R928 out.n138 out.t411 0.000500141
R929 out.n139 out.t205 0.000500141
R930 out.n140 out.t150 0.000500141
R931 out.n141 out.t100 0.000500141
R932 out.n142 out.t391 0.000500141
R933 out.n143 out.t295 0.000500141
R934 out.n144 out.t237 0.000500141
R935 out.n145 out.t185 0.000500141
R936 out.n146 out.t131 0.000500141
R937 out.n147 out.t81 0.000500141
R938 out.n148 out.t321 0.000500141
R939 out.n149 out.t268 0.000500141
R940 out.n150 out.t212 0.000500141
R941 out.n151 out.t95 0.000500141
R942 out.n152 out.t385 0.000500141
R943 out.n153 out.t290 0.000500141
R944 out.n154 out.t231 0.000500141
R945 out.n155 out.t179 0.000500141
R946 out.n156 out.t122 0.000500141
R947 out.n157 out.t414 0.000500141
R948 out.n158 out.t318 0.000500141
R949 out.n159 out.t262 0.000500141
R950 out.n160 out.t206 0.000500141
R951 out.n161 out.t153 0.000500141
R952 out.n162 out.t123 0.000500141
R953 out.n163 out.t362 0.000500141
R954 out.n164 out.t266 0.000500141
R955 out.n165 out.t209 0.000500141
R956 out.n166 out.t156 0.000500141
R957 out.n167 out.t104 0.000500141
R958 out.n168 out.t398 0.000500141
R959 out.n169 out.t298 0.000500141
R960 out.n170 out.t99 0.000500141
R961 out.n171 out.t389 0.000500141
R962 out.n172 out.t331 0.000500141
R963 out.n173 out.t279 0.000500141
R964 out.n174 out.t183 0.000500141
R965 out.n175 out.t128 0.000500141
R966 out.n176 out.t80 0.000500141
R967 out.n177 out.t363 0.000500141
R968 out.n178 out.t309 0.000500141
R969 out.n179 out.t210 0.000500141
R970 out.n180 out.t157 0.000500141
R971 out.n181 out.t106 0.000500141
R972 out.n182 out.t327 0.000500141
R973 out.n183 out.t272 0.000500141
R974 out.n184 out.t178 0.000500141
R975 out.n185 out.t121 0.000500141
R976 out.n186 out.t413 0.000500141
R977 out.n187 out.t353 0.000500141
R978 out.n188 out.t303 0.000500141
R979 out.n189 out.t204 0.000500141
R980 out.n190 out.t151 0.000500141
R981 out.n191 out.t101 0.000500141
R982 out.n192 out.t390 0.000500141
R983 out.n193 out.t355 0.000500141
R984 out.n194 out.t94 0.000500141
R985 out.n195 out.t336 0.000500141
R986 out.n196 out.t289 0.000500141
R987 out.n197 out.t229 0.000500141
R988 out.n198 out.t176 0.000500141
R989 out.n199 out.t120 0.000500141
R990 out.n200 out.t373 0.000500141
R991 out.n201 out.t170 0.000500141
R992 out.n202 out.t114 0.000500141
R993 out.n203 out.t409 0.000500141
R994 out.n204 out.t346 0.000500141
R995 out.n205 out.t255 0.000500141
R996 out.n206 out.t200 0.000500141
R997 out.n207 out.t144 0.000500141
R998 out.n208 out.t93 0.000500141
R999 out.n209 out.t382 0.000500141
R1000 out.n210 out.t288 0.000500141
R1001 out.n211 out.t230 0.000500141
R1002 out.n212 out.t177 0.000500141
R1003 out.n213 out.t406 0.000500141
R1004 out.n214 out.t342 0.000500141
R1005 out.n215 out.t248 0.000500141
R1006 out.n216 out.t193 0.000500141
R1007 out.n217 out.t139 0.000500141
R1008 out.n218 out.t88 0.000500141
R1009 out.n219 out.t375 0.000500141
R1010 out.n220 out.t284 0.000500141
R1011 out.n221 out.t222 0.000500141
R1012 out.n222 out.t171 0.000500141
R1013 out.n223 out.t117 0.000500141
R1014 out.n224 out.t89 0.000500141
R1015 out.n225 out.t97 0.000500141
R1016 out.n226 out.t83 0.000500141
R1017 out.n227 out.t287 0.000500141
R1018 out.n228 out.t149 0.000500141
R1019 out.n229 out.t350 0.000500141
R1020 out.n230 out.t217 0.000500141
R1021 out.n231 out.t198 0.000500141
R1022 out.n232 out.t103 0.000500141
R1023 out.n233 out.t312 0.000500141
R1024 out.n234 out.t174 0.000500141
R1025 out.n235 out.t386 0.000500141
R1026 out.n236 out.t364 0.000500141
R1027 out.n237 out.t226 0.000500141
R1028 out.n238 out.t96 0.000500141
R1029 out.n239 out.t301 0.000500141
R1030 out.n240 out.t165 0.000500141
R1031 out.n241 out.t142 0.000500141
R1032 out.n242 out.t347 0.000500141
R1033 out.n243 out.t215 0.000500141
R1034 out.n244 out.t146 0.000500141
R1035 out.n245 out.t349 0.000500141
R1036 out.n246 out.t332 0.000500141
R1037 out.n247 out.t197 0.000500141
R1038 out.n248 out.t410 0.000500141
R1039 out.n249 out.t273 0.000500141
R1040 out.n250 out.t136 0.000500141
R1041 out.n251 out.t116 0.000500141
R1042 out.n252 out.t325 0.000500141
R1043 out.n253 out.t188 0.000500141
R1044 out.n254 out.t400 0.000500141
R1045 out.n255 out.t392 0.000500141
R1046 out.n256 out.t202 0.000500141
R1047 out.n257 out.t108 0.000500141
R1048 out.n258 out.t402 0.000500141
R1049 out.n259 out.t339 0.000500141
R1050 out.n260 out.t291 0.000500141
R1051 out.n261 out.t233 0.000500141
R1052 out.n262 out.t138 0.000500141
R1053 out.n263 out.t282 0.000500141
R1054 out.n264 out.t223 0.000500141
R1055 out.n265 out.t172 0.000500141
R1056 out.n266 out.t115 0.000500141
R1057 out.n267 out.t366 0.000500141
R1058 out.n268 out.t314 0.000500141
R1059 out.n269 out.t257 0.000500141
R1060 out.n270 out.t203 0.000500141
R1061 out.n271 out.t148 0.000500141
R1062 out.n272 out.t403 0.000500141
R1063 out.n273 out.t340 0.000500141
R1064 out.n274 out.t293 0.000500141
R1065 out.n275 out.t168 0.000500141
R1066 out.n276 out.t113 0.000500141
R1067 out.n277 out.t360 0.000500141
R1068 out.n278 out.t308 0.000500141
R1069 out.n279 out.t251 0.000500141
R1070 out.n280 out.t195 0.000500141
R1071 out.n281 out.t140 0.000500141
R1072 out.n282 out.t396 0.000500141
R1073 out.n283 out.t334 0.000500141
R1074 out.n284 out.t286 0.000500141
R1075 out.n285 out.t224 0.000500141
R1076 out.n286 out.t196 0.000500141
R1077 out.n287 out.t277 0.000500141
R1078 out.n288 out.t182 0.000500141
R1079 out.n289 out.t125 0.000500141
R1080 out.n290 out.t416 0.000500141
R1081 out.n291 out.t358 0.000500141
R1082 out.n292 out.t307 0.000500141
R1083 out.n293 out.t208 0.000500141
R1084 out.n294 out.t348 0.000500141
R1085 out.n295 out.t299 0.000500141
R1086 out.n296 out.t242 0.000500141
R1087 out.n297 out.t190 0.000500141
R1088 out.n298 out.t98 0.000500141
R1089 out.n299 out.t388 0.000500141
R1090 out.n300 out.t330 0.000500141
R1091 out.n301 out.t278 0.000500141
R1092 out.n302 out.t220 0.000500141
R1093 out.n303 out.t126 0.000500141
R1094 out.n304 out.t418 0.000500141
R1095 out.n305 out.t359 0.000500141
R1096 out.n306 out.t240 0.000500141
R1097 out.n307 out.t187 0.000500141
R1098 out.n308 out.t92 0.000500141
R1099 out.n309 out.t380 0.000500141
R1100 out.n310 out.t326 0.000500141
R1101 out.n311 out.t271 0.000500141
R1102 out.n312 out.t214 0.000500141
R1103 out.n313 out.t119 0.000500141
R1104 out.n314 out.t412 0.000500141
R1105 out.n315 out.t352 0.000500141
R1106 out.n316 out.t302 0.000500141
R1107 out.n317 out.t274 0.000500141
R1108 out.n319 out.t304 0.000500141
R1109 out.n321 out.t228 0.000500141
R1110 out.n323 out.t337 0.000500141
R1111 out.n324 out.t311 0.000500141
R1112 out.n325 out.t335 0.000500141
R1113 out.n326 out.t399 0.000500141
R1114 out.n327 out.t105 0.000500141
R1115 out.n328 out.t158 0.000500141
R1116 out.n329 out.t252 0.000500141
R1117 out.n330 out.t310 0.000500141
R1118 out.n331 out.t361 0.000500141
R1119 out.n332 out.t419 0.000500141
R1120 out.n333 out.t129 0.000500141
R1121 out.n334 out.t221 0.000500141
R1122 out.n335 out.t280 0.000500141
R1123 out.n336 out.t405 0.000500141
R1124 out.n337 out.t110 0.000500141
R1125 out.n338 out.t164 0.000500141
R1126 out.n339 out.t259 0.000500141
R1127 out.n340 out.t316 0.000500141
R1128 out.n341 out.t370 0.000500141
R1129 out.n342 out.t85 0.000500141
R1130 out.n343 out.t133 0.000500141
R1131 out.n344 out.t225 0.000500141
R1132 out.n345 out.t285 0.000500141
R1133 out.n346 out.t333 0.000500141
R1134 out.n347 out.t397 0.000500141
R1135 out.n348 out.t247 0.000500141
R1136 out.n349 out.t341 0.000500141
R1137 out.n350 out.t404 0.000500141
R1138 out.n351 out.t109 0.000500141
R1139 out.n352 out.t163 0.000500141
R1140 out.n353 out.t216 0.000500141
R1141 out.n354 out.t315 0.000500141
R1142 out.n355 out.t367 0.000500141
R1143 out.n356 out.t84 0.000500141
R1144 out.n357 out.t313 0.000500141
R1145 out.n358 out.t387 0.000500141
R1146 out.n359 out.t275 0.000500141
R1147 out.n360 out.t344 0.000500141
R1148 out.n361 out.t236 0.000500141
R1149 out.n362 out.t127 0.000500141
R1150 out.n363 out.t199 0.000500141
R1151 out.n364 out.t365 0.000500141
R1152 out.n365 out.t294 0.000500141
R1153 out.n367 out.t169 0.000500141
R1154 out.n368 out.t394 0.000500141
R1155 out.n369 out.t181 0.000500141
R1156 out.n370 out.t408 0.000500141
R1157 out.n371 out.t283 0.000500141
R1158 out.n372 out.t159 0.000500141
R1159 out.n373 out.t384 0.000500141
R1160 out.n374 out.t173 0.000500141
R1161 out.n375 out.t281 0.000500141
R1162 out.n376 out.t154 0.000500141
R1163 out.n377 out.t376 0.000500141
R1164 out.n378 out.t254 0.000500141
R1165 out.n379 out.t393 0.000500141
R1166 out.n380 out.t265 0.000500141
R1167 out.n381 out.t143 0.000500141
R1168 out.n382 out.t369 0.000500141
R1169 out.n383 out.t244 0.000500141
R1170 out.n384 out.t383 0.000500141
R1171 out.n385 out.t260 0.000500141
R1172 out.n386 out.t137 0.000500141
R1173 out.n387 out.t368 0.000500141
R1174 out.n388 out.t243 0.000500141
R1175 out.n389 out.t381 0.000500141
R1176 out.n390 out.t258 0.000500141
R1177 out.n391 out.t135 0.000500141
R1178 out.n392 out.t354 0.000500141
R1179 out.n393 out.t234 0.000500141
R1180 out.n394 out.t372 0.000500141
R1181 out.n395 out.t246 0.000500141
R1182 out.n396 out.t124 0.000500141
R1183 out.n397 out.t343 0.000500141
R1184 out.n398 out.t111 0.000500141
R1185 out.n399 out.t371 0.000500141
R1186 out.n402 out.t253 0.000500141
R1187 out.n404 out.t118 0.000500141
R1188 out.n406 out.t395 0.000500141
R1189 out.n408 out.t155 0.000500141
R1190 out.n410 out.t264 0.000500141
R1191 out.n100 out.t192 0.000500141
R1192 out.n412 out.t162 0.000500141
R1193 out.n413 out.t191 0.000500141
R1194 out.n414 out.t245 0.000500141
R1195 out.n72 out.t166 0.000500141
R1196 out.n73 out.t415 0.000500141
R1197 out.n74 out.t356 0.000500141
R1198 out.n75 out.t305 0.000500141
R1199 out.n76 out.t249 0.000500141
R1200 out.n77 out.t194 0.000500141
R1201 out.n78 out.t102 0.000500141
R1202 out.n79 out.t241 0.000500141
R1203 out.n80 out.t189 0.000500141
R1204 out.n81 out.t134 0.000500141
R1205 out.n82 out.t86 0.000500141
R1206 out.n83 out.t328 0.000500141
R1207 out.n84 out.t276 0.000500141
R1208 out.n85 out.t219 0.000500141
R1209 out.n86 out.t167 0.000500141
R1210 out.n87 out.t112 0.000500141
R1211 out.n88 out.t357 0.000500141
R1212 out.n89 out.t306 0.000500141
R1213 out.n90 out.t250 0.000500141
R1214 out.n91 out.t132 0.000500141
R1215 out.n92 out.t82 0.000500141
R1216 out.n93 out.t324 0.000500141
R1217 out.n94 out.t270 0.000500141
R1218 out.n95 out.t213 0.000500141
R1219 out.n96 out.t161 0.000500141
R1220 out.n97 out.t107 0.000500141
R1221 out.n98 out.t351 0.000500141
R1222 out.n99 out.t300 0.000500141
R1223 sky130_fd_sc_hd__inv_2_1.Y.n3 sky130_fd_sc_hd__inv_2_1.Y.n2 111.322
R1224 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_sc_hd__inv_2_1.Y.n4 50.4671
R1225 sky130_fd_sc_hd__inv_2_1.Y.n2 sky130_fd_sc_hd__inv_2_1.Y.t3 26.5955
R1226 sky130_fd_sc_hd__inv_2_1.Y.n2 sky130_fd_sc_hd__inv_2_1.Y.t4 26.5955
R1227 sky130_fd_sc_hd__inv_2_1.Y.n4 sky130_fd_sc_hd__inv_2_1.Y.t1 24.9236
R1228 sky130_fd_sc_hd__inv_2_1.Y.n4 sky130_fd_sc_hd__inv_2_1.Y.t2 24.9236
R1229 sky130_fd_sc_hd__inv_2_1.Y.n6 sky130_fd_sc_hd__inv_2_1.Y 13.0565
R1230 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_sc_hd__inv_2_1.Y.n5 11.2645
R1231 sky130_fd_sc_hd__inv_2_1.Y.n5 sky130_fd_sc_hd__inv_2_1.Y 6.1445
R1232 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_sc_hd__inv_2_1.Y.n6 5.55958
R1233 sky130_fd_sc_hd__inv_2_1.Y.n5 sky130_fd_sc_hd__inv_2_1.Y 4.65505
R1234 sky130_fd_sc_hd__inv_2_1.Y.n6 sky130_fd_sc_hd__inv_2_1.Y 4.3525
R1235 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_sc_hd__inv_2_1.Y.n3 2.0485
R1236 sky130_fd_sc_hd__inv_2_1.Y.n3 sky130_fd_sc_hd__inv_2_1.Y 1.55202
R1237 sky130_fd_sc_hd__inv_2_1.Y.t0 sky130_fd_sc_hd__inv_2_1.Y 0.11204
R1238 sky130_fd_sc_hd__inv_2_1.Y.n1 sky130_fd_sc_hd__inv_2_1.Y 0.107011
R1239 sky130_fd_sc_hd__inv_2_1.Y.n1 sky130_fd_sc_hd__inv_2_1.Y.n0 0.0358951
R1240 sky130_fd_sc_hd__inv_2_1.Y.t0 sky130_fd_sc_hd__inv_2_1.Y.n1 0.0237099
R1241 sky130_fd_sc_hd__inv_2_2.Y.n1 sky130_fd_sc_hd__inv_2_2.Y.n0 111.322
R1242 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_sc_hd__inv_2_2.Y.n2 50.4671
R1243 sky130_fd_sc_hd__inv_2_2.Y.n0 sky130_fd_sc_hd__inv_2_2.Y.t0 26.5955
R1244 sky130_fd_sc_hd__inv_2_2.Y.n0 sky130_fd_sc_hd__inv_2_2.Y.t4 26.5955
R1245 sky130_fd_sc_hd__inv_2_2.Y.n2 sky130_fd_sc_hd__inv_2_2.Y.t1 24.9236
R1246 sky130_fd_sc_hd__inv_2_2.Y.n2 sky130_fd_sc_hd__inv_2_2.Y.t5 24.9236
R1247 sky130_fd_sc_hd__inv_2_2.Y.n4 sky130_fd_sc_hd__inv_2_2.Y 13.5685
R1248 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_sc_hd__inv_2_2.Y.n3 11.2645
R1249 sky130_fd_sc_hd__inv_2_2.Y.n3 sky130_fd_sc_hd__inv_2_2.Y 6.1445
R1250 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_sc_hd__inv_2_2.Y.n4 5.17077
R1251 sky130_fd_sc_hd__inv_2_2.Y.n3 sky130_fd_sc_hd__inv_2_2.Y 4.65505
R1252 sky130_fd_sc_hd__inv_2_2.Y.n4 sky130_fd_sc_hd__inv_2_2.Y 3.8405
R1253 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_sc_hd__inv_2_2.Y.n1 2.0485
R1254 sky130_fd_sc_hd__inv_2_2.Y.n1 sky130_fd_sc_hd__inv_2_2.Y 1.55202
R1255 sky130_fd_sc_hd__inv_2_2.Y.t2 sky130_fd_sc_hd__inv_2_2.Y 0.197458
R1256 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_sc_hd__inv_2_2.Y.t2 0.1012
R1257 sky130_fd_sc_hd__inv_2_2.Y.t2 sky130_fd_sc_hd__inv_2_2.Y 0.00959054
R1258 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_sc_hd__inv_2_2.Y.t3 0.00959054
R1259 vin.n8 vin.t55 29.3118
R1260 vin.n22 vin.t61 29.3118
R1261 vin.n37 vin.t45 29.3118
R1262 vin.n52 vin.t76 29.3118
R1263 vin.n13 vin.t50 29.3084
R1264 vin.n27 vin.t65 29.3084
R1265 vin.n42 vin.t48 29.3084
R1266 vin.n57 vin.t72 29.3084
R1267 vin.n6 vin.t51 28.5655
R1268 vin.n6 vin.t59 28.5655
R1269 vin.n4 vin.t56 28.5655
R1270 vin.n4 vin.t52 28.5655
R1271 vin.n2 vin.t57 28.5655
R1272 vin.n2 vin.t53 28.5655
R1273 vin.n0 vin.t58 28.5655
R1274 vin.n0 vin.t54 28.5655
R1275 vin.n20 vin.t67 28.5655
R1276 vin.n20 vin.t62 28.5655
R1277 vin.n18 vin.t68 28.5655
R1278 vin.n18 vin.t63 28.5655
R1279 vin.n16 vin.t69 28.5655
R1280 vin.n16 vin.t66 28.5655
R1281 vin.n14 vin.t64 28.5655
R1282 vin.n14 vin.t60 28.5655
R1283 vin.n35 vin.t40 28.5655
R1284 vin.n35 vin.t46 28.5655
R1285 vin.n33 vin.t41 28.5655
R1286 vin.n33 vin.t47 28.5655
R1287 vin.n31 vin.t42 28.5655
R1288 vin.n31 vin.t49 28.5655
R1289 vin.n29 vin.t43 28.5655
R1290 vin.n29 vin.t44 28.5655
R1291 vin.n50 vin.t70 28.5655
R1292 vin.n50 vin.t77 28.5655
R1293 vin.n48 vin.t73 28.5655
R1294 vin.n48 vin.t71 28.5655
R1295 vin.n46 vin.t74 28.5655
R1296 vin.n46 vin.t78 28.5655
R1297 vin.n44 vin.t79 28.5655
R1298 vin.n44 vin.t75 28.5655
R1299 vin.n8 vin.t25 18.1397
R1300 vin.n13 vin.t29 18.1397
R1301 vin.n22 vin.t8 18.1397
R1302 vin.n27 vin.t3 18.1397
R1303 vin.n37 vin.t12 18.1397
R1304 vin.n42 vin.t16 18.1397
R1305 vin.n52 vin.t36 18.1397
R1306 vin.n57 vin.t31 18.1397
R1307 vin.n7 vin.t20 17.4005
R1308 vin.n7 vin.t27 17.4005
R1309 vin.n5 vin.t24 17.4005
R1310 vin.n5 vin.t21 17.4005
R1311 vin.n3 vin.t28 17.4005
R1312 vin.n3 vin.t22 17.4005
R1313 vin.n1 vin.t26 17.4005
R1314 vin.n1 vin.t23 17.4005
R1315 vin.n21 vin.t4 17.4005
R1316 vin.n21 vin.t9 17.4005
R1317 vin.n19 vin.t5 17.4005
R1318 vin.n19 vin.t1 17.4005
R1319 vin.n17 vin.t6 17.4005
R1320 vin.n17 vin.t2 17.4005
R1321 vin.n15 vin.t0 17.4005
R1322 vin.n15 vin.t7 17.4005
R1323 vin.n36 vin.t18 17.4005
R1324 vin.n36 vin.t15 17.4005
R1325 vin.n34 vin.t19 17.4005
R1326 vin.n34 vin.t13 17.4005
R1327 vin.n32 vin.t10 17.4005
R1328 vin.n32 vin.t17 17.4005
R1329 vin.n30 vin.t14 17.4005
R1330 vin.n30 vin.t11 17.4005
R1331 vin.n51 vin.t32 17.4005
R1332 vin.n51 vin.t37 17.4005
R1333 vin.n49 vin.t33 17.4005
R1334 vin.n49 vin.t39 17.4005
R1335 vin.n47 vin.t34 17.4005
R1336 vin.n47 vin.t30 17.4005
R1337 vin.n45 vin.t38 17.4005
R1338 vin.n45 vin.t35 17.4005
R1339 vin.n61 vin.n60 8.92094
R1340 vin.n59 vin.n58 8.59648
R1341 vin.n60 vin.n59 6.6802
R1342 vin.n61 vin 3.04911
R1343 vin.n59 vin.n43 1.91314
R1344 vin.n60 vin.n28 1.91178
R1345 vin.n10 vin.n9 0.811311
R1346 vin.n24 vin.n23 0.811311
R1347 vin.n39 vin.n38 0.811311
R1348 vin.n54 vin.n53 0.811311
R1349 vin.n12 vin.n11 0.799575
R1350 vin.n26 vin.n25 0.799575
R1351 vin.n41 vin.n40 0.799575
R1352 vin.n56 vin.n55 0.799575
R1353 vin.n11 vin.n10 0.794419
R1354 vin.n25 vin.n24 0.794419
R1355 vin.n40 vin.n39 0.794419
R1356 vin.n55 vin.n54 0.794419
R1357 vin.n9 vin.n8 0.787662
R1358 vin.n23 vin.n22 0.787662
R1359 vin.n38 vin.n37 0.787662
R1360 vin.n53 vin.n52 0.787662
R1361 vin.n13 vin.n12 0.773526
R1362 vin.n27 vin.n26 0.773526
R1363 vin.n42 vin.n41 0.773526
R1364 vin.n57 vin.n56 0.773526
R1365 vin.n9 vin.n6 0.746823
R1366 vin.n10 vin.n4 0.746823
R1367 vin.n11 vin.n2 0.746823
R1368 vin.n23 vin.n20 0.746823
R1369 vin.n24 vin.n18 0.746823
R1370 vin.n25 vin.n16 0.746823
R1371 vin.n38 vin.n35 0.746823
R1372 vin.n39 vin.n33 0.746823
R1373 vin.n40 vin.n31 0.746823
R1374 vin.n53 vin.n50 0.746823
R1375 vin.n54 vin.n48 0.746823
R1376 vin.n55 vin.n46 0.746823
R1377 vin.n12 vin.n0 0.743351
R1378 vin.n26 vin.n14 0.743351
R1379 vin.n41 vin.n29 0.743351
R1380 vin.n56 vin.n44 0.743351
R1381 vin.n9 vin.n7 0.739748
R1382 vin.n10 vin.n5 0.739748
R1383 vin.n11 vin.n3 0.739748
R1384 vin.n12 vin.n1 0.739748
R1385 vin.n23 vin.n21 0.739748
R1386 vin.n24 vin.n19 0.739748
R1387 vin.n25 vin.n17 0.739748
R1388 vin.n26 vin.n15 0.739748
R1389 vin.n38 vin.n36 0.739748
R1390 vin.n39 vin.n34 0.739748
R1391 vin.n40 vin.n32 0.739748
R1392 vin.n41 vin.n30 0.739748
R1393 vin.n53 vin.n51 0.739748
R1394 vin.n54 vin.n49 0.739748
R1395 vin.n55 vin.n47 0.739748
R1396 vin.n56 vin.n45 0.739748
R1397 vin vin.n13 0.636099
R1398 vin.n28 vin.n27 0.580651
R1399 vin.n43 vin.n42 0.579111
R1400 vin.n58 vin.n57 0.573599
R1401 vin vin.n61 0.274806
R1402 vin.n58 vin 0.063
R1403 vin.n43 vin 0.0583961
R1404 vin.n28 vin 0.056769
R1405 vdd.n46 vdd.n42 6176.47
R1406 vdd.n93 vdd.n89 6176.47
R1407 vdd.n18 vdd.n14 6176.47
R1408 vdd.n186 vdd.n179 6176.47
R1409 vdd.n47 vdd.n46 3240
R1410 vdd.n94 vdd.n93 3240
R1411 vdd.n19 vdd.n18 3240
R1412 vdd.n183 vdd.n179 3240
R1413 vdd.n47 vdd.n45 3056.47
R1414 vdd.n94 vdd.n92 3056.47
R1415 vdd.n19 vdd.n17 3056.47
R1416 vdd.n184 vdd.n183 3056.47
R1417 vdd.t53 vdd 895.586
R1418 vdd.t41 vdd 895.586
R1419 vdd vdd.t22 895.586
R1420 vdd.t47 vdd 895.586
R1421 vdd.n40 vdd.t122 584.644
R1422 vdd.n71 vdd.t11 584.644
R1423 vdd.n127 vdd.t74 584.644
R1424 vdd.n120 vdd.t6 584.644
R1425 vdd.n12 vdd.t118 584.644
R1426 vdd.n160 vdd.t15 584.644
R1427 vdd.n216 vdd.t91 584.644
R1428 vdd.n209 vdd.t21 584.644
R1429 vdd.t23 vdd.n168 512.547
R1430 vdd.n111 vdd.t42 512.547
R1431 vdd.t54 vdd.n79 512.547
R1432 vdd.n200 vdd.t48 512.547
R1433 vdd.t50 vdd.n30 489.178
R1434 vdd.n169 vdd.t23 459.192
R1435 vdd.n109 vdd.t42 459.192
R1436 vdd.n80 vdd.t54 459.192
R1437 vdd.n198 vdd.t48 459.192
R1438 vdd vdd.n137 428.521
R1439 vdd.n138 vdd 428.521
R1440 vdd vdd.n226 428.521
R1441 vdd.n228 vdd 428.521
R1442 vdd.t44 vdd 378.64
R1443 vdd vdd.t25 378.64
R1444 vdd.t28 vdd 378.64
R1445 vdd.n137 vdd.t53 340.096
R1446 vdd.n138 vdd.t41 340.096
R1447 vdd.n226 vdd.t22 340.096
R1448 vdd.n228 vdd.t47 340.096
R1449 vdd.t121 vdd 301.551
R1450 vdd.t73 vdd 301.551
R1451 vdd vdd.t117 301.551
R1452 vdd.t90 vdd 301.551
R1453 vdd.n46 vdd.t125 289.37
R1454 vdd.n93 vdd.t78 289.37
R1455 vdd.n18 vdd.t110 289.37
R1456 vdd.t80 vdd.n179 289.37
R1457 vdd.n49 vdd.t133 287.676
R1458 vdd.n96 vdd.t71 287.676
R1459 vdd.n21 vdd.t104 287.676
R1460 vdd.t89 vdd.n181 287.676
R1461 vdd.t10 vdd 285.68
R1462 vdd.t5 vdd 285.68
R1463 vdd vdd.t14 285.68
R1464 vdd.t20 vdd 285.68
R1465 vdd vdd.t50 247.137
R1466 vdd vdd.t44 247.137
R1467 vdd.t25 vdd 247.137
R1468 vdd vdd.t28 247.137
R1469 vdd.n229 vdd.t49 243.03
R1470 vdd.n224 vdd.t24 243.03
R1471 vdd.n29 vdd.t43 243.03
R1472 vdd.n135 vdd.t55 243.03
R1473 vdd vdd.n227 242.905
R1474 vdd.n56 vdd.t51 234.554
R1475 vdd.n59 vdd.t52 234.554
R1476 vdd.n86 vdd.t45 234.554
R1477 vdd.n129 vdd.t46 234.554
R1478 vdd.n145 vdd.t26 234.554
R1479 vdd.n148 vdd.t27 234.554
R1480 vdd.n175 vdd.t29 234.554
R1481 vdd.n218 vdd.t30 234.554
R1482 vdd.t133 vdd.t123 197.359
R1483 vdd.t123 vdd.t136 197.359
R1484 vdd.t136 vdd.t130 197.359
R1485 vdd.t130 vdd.t124 197.359
R1486 vdd.t137 vdd.t131 197.359
R1487 vdd.t138 vdd.t137 197.359
R1488 vdd.t132 vdd.t138 197.359
R1489 vdd.t125 vdd.t132 197.359
R1490 vdd.t71 vdd.t64 197.359
R1491 vdd.t64 vdd.t72 197.359
R1492 vdd.t72 vdd.t67 197.359
R1493 vdd.t67 vdd.t75 197.359
R1494 vdd.t79 vdd.t68 197.359
R1495 vdd.t69 vdd.t79 197.359
R1496 vdd.t70 vdd.t69 197.359
R1497 vdd.t78 vdd.t70 197.359
R1498 vdd.t104 vdd.t114 197.359
R1499 vdd.t114 vdd.t107 197.359
R1500 vdd.t107 vdd.t119 197.359
R1501 vdd.t119 vdd.t108 197.359
R1502 vdd.t111 vdd.t120 197.359
R1503 vdd.t109 vdd.t111 197.359
R1504 vdd.t103 vdd.t109 197.359
R1505 vdd.t110 vdd.t103 197.359
R1506 vdd.t83 vdd.t89 197.359
R1507 vdd.t97 vdd.t83 197.359
R1508 vdd.t92 vdd.t97 197.359
R1509 vdd.t84 vdd.t92 197.359
R1510 vdd.t93 vdd.t85 197.359
R1511 vdd.t85 vdd.t94 197.359
R1512 vdd.t94 vdd.t86 197.359
R1513 vdd.t86 vdd.t80 197.359
R1514 vdd.t128 vdd.t121 190.453
R1515 vdd.t134 vdd.t128 190.453
R1516 vdd.t126 vdd.t134 190.453
R1517 vdd.t2 vdd.t10 190.453
R1518 vdd.t16 vdd.t2 190.453
R1519 vdd.t8 vdd.t16 190.453
R1520 vdd.t65 vdd.t73 190.453
R1521 vdd.t76 vdd.t65 190.453
R1522 vdd.t62 vdd.t76 190.453
R1523 vdd.t141 vdd.t5 190.453
R1524 vdd.t37 vdd.t141 190.453
R1525 vdd.t33 vdd.t37 190.453
R1526 vdd.t117 vdd.t115 190.453
R1527 vdd.t115 vdd.t105 190.453
R1528 vdd.t105 vdd.t112 190.453
R1529 vdd.t14 vdd.t12 190.453
R1530 vdd.t12 vdd.t139 190.453
R1531 vdd.t139 vdd.t18 190.453
R1532 vdd.t81 vdd.t90 190.453
R1533 vdd.t95 vdd.t81 190.453
R1534 vdd.t87 vdd.t95 190.453
R1535 vdd.t35 vdd.t20 190.453
R1536 vdd.t98 vdd.t35 190.453
R1537 vdd.t101 vdd.t98 190.453
R1538 vdd.n137 vdd.n136 185
R1539 vdd.n139 vdd.n138 185
R1540 vdd.n226 vdd.n225 185
R1541 vdd.n230 vdd.n228 185
R1542 vdd.n66 vdd.n39 174.595
R1543 vdd.n73 vdd.n36 174.595
R1544 vdd.n103 vdd.n102 174.595
R1545 vdd.n107 vdd.n106 174.595
R1546 vdd.n155 vdd.n11 174.595
R1547 vdd.n162 vdd.n8 174.595
R1548 vdd.n192 vdd.n191 174.595
R1549 vdd.n196 vdd.n195 174.595
R1550 vdd vdd.t126 170.048
R1551 vdd vdd.t8 170.048
R1552 vdd vdd.t62 170.048
R1553 vdd vdd.t33 170.048
R1554 vdd.t112 vdd 170.048
R1555 vdd.t18 vdd 170.048
R1556 vdd vdd.t87 170.048
R1557 vdd vdd.t101 170.048
R1558 vdd.n57 vdd.t153 166.282
R1559 vdd.n87 vdd.t148 166.282
R1560 vdd.n146 vdd.t151 166.282
R1561 vdd.n176 vdd.t152 166.282
R1562 vdd.n37 vdd.t127 151.123
R1563 vdd.n77 vdd.t9 151.123
R1564 vdd.n121 vdd.t63 151.123
R1565 vdd.n114 vdd.t34 151.123
R1566 vdd.n9 vdd.t113 151.123
R1567 vdd.n166 vdd.t19 151.123
R1568 vdd.n210 vdd.t88 151.123
R1569 vdd.n203 vdd.t102 151.123
R1570 vdd.t124 vdd.n48 98.6801
R1571 vdd.n48 vdd.t131 98.6801
R1572 vdd.t75 vdd.n95 98.6801
R1573 vdd.n95 vdd.t68 98.6801
R1574 vdd.t108 vdd.n20 98.6801
R1575 vdd.n20 vdd.t120 98.6801
R1576 vdd.n182 vdd.t84 98.6801
R1577 vdd.n182 vdd.t93 98.6801
R1578 vdd.n169 vdd.t150 92.9047
R1579 vdd.n109 vdd.t147 92.9047
R1580 vdd.n80 vdd.t146 92.9047
R1581 vdd.n198 vdd.t149 92.9047
R1582 vdd.n50 vdd.n43 76.5867
R1583 vdd.n97 vdd.n90 76.5867
R1584 vdd.n22 vdd.n15 76.5867
R1585 vdd.n180 vdd.n178 76.5867
R1586 vdd.n66 vdd.n65 34.6358
R1587 vdd.n67 vdd.n66 34.6358
R1588 vdd.n73 vdd.n72 34.6358
R1589 vdd.n73 vdd.n34 34.6358
R1590 vdd.n126 vdd.n103 34.6358
R1591 vdd.n122 vdd.n103 34.6358
R1592 vdd.n119 vdd.n107 34.6358
R1593 vdd.n115 vdd.n107 34.6358
R1594 vdd.n155 vdd.n154 34.6358
R1595 vdd.n156 vdd.n155 34.6358
R1596 vdd.n162 vdd.n161 34.6358
R1597 vdd.n162 vdd.n6 34.6358
R1598 vdd.n215 vdd.n192 34.6358
R1599 vdd.n211 vdd.n192 34.6358
R1600 vdd.n208 vdd.n196 34.6358
R1601 vdd.n204 vdd.n196 34.6358
R1602 vdd.n55 vdd 29.3839
R1603 vdd.n235 vdd.n0 27.8654
R1604 vdd.n39 vdd.t129 26.5955
R1605 vdd.n39 vdd.t135 26.5955
R1606 vdd.n36 vdd.t3 26.5955
R1607 vdd.n36 vdd.t17 26.5955
R1608 vdd.n102 vdd.t66 26.5955
R1609 vdd.n102 vdd.t77 26.5955
R1610 vdd.n106 vdd.t142 26.5955
R1611 vdd.n106 vdd.t38 26.5955
R1612 vdd.n11 vdd.t116 26.5955
R1613 vdd.n11 vdd.t106 26.5955
R1614 vdd.n8 vdd.t13 26.5955
R1615 vdd.n8 vdd.t140 26.5955
R1616 vdd.n191 vdd.t82 26.5955
R1617 vdd.n191 vdd.t96 26.5955
R1618 vdd.n195 vdd.t36 26.5955
R1619 vdd.n195 vdd.t99 26.5955
R1620 vdd.n65 vdd.n40 22.2123
R1621 vdd.n67 vdd.n37 22.2123
R1622 vdd.n72 vdd.n71 22.2123
R1623 vdd.n77 vdd.n34 22.2123
R1624 vdd.n127 vdd.n126 22.2123
R1625 vdd.n122 vdd.n121 22.2123
R1626 vdd.n120 vdd.n119 22.2123
R1627 vdd.n115 vdd.n114 22.2123
R1628 vdd.n154 vdd.n12 22.2123
R1629 vdd.n156 vdd.n9 22.2123
R1630 vdd.n161 vdd.n160 22.2123
R1631 vdd.n166 vdd.n6 22.2123
R1632 vdd.n216 vdd.n215 22.2123
R1633 vdd.n211 vdd.n210 22.2123
R1634 vdd.n209 vdd.n208 22.2123
R1635 vdd.n204 vdd.n203 22.2123
R1636 vdd.n60 vdd.n40 21.8029
R1637 vdd.n128 vdd.n127 21.8029
R1638 vdd.n149 vdd.n12 21.8029
R1639 vdd.n217 vdd.n216 21.8029
R1640 vdd.n71 vdd.n37 21.0829
R1641 vdd.n121 vdd.n120 21.0829
R1642 vdd.n160 vdd.n9 21.0829
R1643 vdd.n210 vdd.n209 21.0829
R1644 vdd.n45 vdd.n41 17.2966
R1645 vdd.n92 vdd.n88 17.2966
R1646 vdd.n17 vdd.n13 17.2966
R1647 vdd.n184 vdd.n177 17.2966
R1648 vdd.n51 vdd.n42 16.9954
R1649 vdd.n98 vdd.n89 16.9954
R1650 vdd.n23 vdd.n14 16.9954
R1651 vdd.n187 vdd.n186 16.9954
R1652 vdd.n78 vdd.n77 15.4358
R1653 vdd.n114 vdd.n113 15.4358
R1654 vdd.n167 vdd.n166 15.4358
R1655 vdd.n203 vdd.n202 15.4358
R1656 vdd.n134 vdd.n32 14.2735
R1657 vdd.n144 vdd.n26 14.2735
R1658 vdd.n223 vdd.n4 14.2735
R1659 vdd.n52 vdd.n41 12.4392
R1660 vdd.n99 vdd.n88 12.4392
R1661 vdd.n24 vdd.n13 12.4392
R1662 vdd.n188 vdd.n177 12.4392
R1663 vdd.n50 vdd.n49 9.3005
R1664 vdd.n97 vdd.n96 9.3005
R1665 vdd.n22 vdd.n21 9.3005
R1666 vdd.n181 vdd.n178 9.3005
R1667 vdd.n224 vdd.n223 7.70175
R1668 vdd.n29 vdd.n26 7.70175
R1669 vdd.n135 vdd.n134 7.70175
R1670 vdd.n229 vdd.n0 7.70175
R1671 vdd.n51 vdd.n50 7.66611
R1672 vdd.n98 vdd.n97 7.66611
R1673 vdd.n23 vdd.n22 7.66611
R1674 vdd.n187 vdd.n178 7.66611
R1675 vdd.n203 vdd.n197 4.6505
R1676 vdd.n209 vdd.n194 4.6505
R1677 vdd.n210 vdd.n193 4.6505
R1678 vdd.n216 vdd.n190 4.6505
R1679 vdd.n166 vdd.n165 4.6505
R1680 vdd.n160 vdd.n159 4.6505
R1681 vdd.n158 vdd.n9 4.6505
R1682 vdd.n152 vdd.n12 4.6505
R1683 vdd.n114 vdd.n108 4.6505
R1684 vdd.n120 vdd.n105 4.6505
R1685 vdd.n121 vdd.n104 4.6505
R1686 vdd.n127 vdd.n101 4.6505
R1687 vdd.n77 vdd.n76 4.6505
R1688 vdd.n71 vdd.n70 4.6505
R1689 vdd.n69 vdd.n37 4.6505
R1690 vdd.n63 vdd.n40 4.6505
R1691 vdd.n55 vdd.n54 4.6505
R1692 vdd.n58 vdd.n53 4.6505
R1693 vdd.n61 vdd.n60 4.6505
R1694 vdd.n83 vdd.n82 4.6505
R1695 vdd.n84 vdd.n31 4.6505
R1696 vdd.n132 vdd.n32 4.6505
R1697 vdd.n131 vdd.n130 4.6505
R1698 vdd.n128 vdd.n85 4.6505
R1699 vdd.n28 vdd.n27 4.6505
R1700 vdd.n141 vdd.n140 4.6505
R1701 vdd.n144 vdd.n143 4.6505
R1702 vdd.n147 vdd.n25 4.6505
R1703 vdd.n150 vdd.n149 4.6505
R1704 vdd.n172 vdd.n171 4.6505
R1705 vdd.n173 vdd.n3 4.6505
R1706 vdd.n221 vdd.n4 4.6505
R1707 vdd.n220 vdd.n219 4.6505
R1708 vdd.n217 vdd.n174 4.6505
R1709 vdd.n2 vdd.n1 4.6505
R1710 vdd.n232 vdd.n231 4.6505
R1711 vdd.n205 vdd.n204 4.6505
R1712 vdd.n206 vdd.n196 4.6505
R1713 vdd.n208 vdd.n207 4.6505
R1714 vdd.n212 vdd.n211 4.6505
R1715 vdd.n213 vdd.n192 4.6505
R1716 vdd.n215 vdd.n214 4.6505
R1717 vdd.n164 vdd.n6 4.6505
R1718 vdd.n163 vdd.n162 4.6505
R1719 vdd.n161 vdd.n7 4.6505
R1720 vdd.n157 vdd.n156 4.6505
R1721 vdd.n155 vdd.n10 4.6505
R1722 vdd.n154 vdd.n153 4.6505
R1723 vdd.n116 vdd.n115 4.6505
R1724 vdd.n117 vdd.n107 4.6505
R1725 vdd.n119 vdd.n118 4.6505
R1726 vdd.n123 vdd.n122 4.6505
R1727 vdd.n124 vdd.n103 4.6505
R1728 vdd.n126 vdd.n125 4.6505
R1729 vdd.n75 vdd.n34 4.6505
R1730 vdd.n74 vdd.n73 4.6505
R1731 vdd.n72 vdd.n35 4.6505
R1732 vdd.n68 vdd.n67 4.6505
R1733 vdd.n66 vdd.n38 4.6505
R1734 vdd.n65 vdd.n64 4.6505
R1735 vdd.n59 vdd.n58 4.36875
R1736 vdd.n130 vdd.n129 4.36875
R1737 vdd.n148 vdd.n147 4.36875
R1738 vdd.n219 vdd.n218 4.36875
R1739 vdd.n227 vdd 3.97747
R1740 vdd.n171 vdd.n3 3.57983
R1741 vdd.n140 vdd.n28 3.57983
R1742 vdd.n82 vdd.n31 3.57983
R1743 vdd.n231 vdd.n2 3.57983
R1744 vdd.n58 vdd.n57 3.50526
R1745 vdd.n130 vdd.n87 3.50526
R1746 vdd.n147 vdd.n146 3.50526
R1747 vdd.n219 vdd.n176 3.50526
R1748 vdd vdd.n52 3.35086
R1749 vdd vdd.n99 3.35086
R1750 vdd vdd.n24 3.35086
R1751 vdd vdd.n188 3.34986
R1752 vdd.n30 vdd 3.28549
R1753 vdd.n62 vdd 3.20271
R1754 vdd.n100 vdd 3.20271
R1755 vdd.n151 vdd 3.20271
R1756 vdd.n189 vdd 3.20271
R1757 vdd.n225 vdd.n224 3.08362
R1758 vdd.n139 vdd.n29 3.08362
R1759 vdd.n136 vdd.n135 3.08362
R1760 vdd.n230 vdd.n229 3.08362
R1761 vdd.n170 vdd.n169 2.61352
R1762 vdd.n110 vdd.n109 2.61352
R1763 vdd.n81 vdd.n80 2.61352
R1764 vdd.n199 vdd.n198 2.61352
R1765 vdd.n30 vdd 2.57272
R1766 vdd.n134 vdd.n133 2.29662
R1767 vdd.n142 vdd.n26 2.29662
R1768 vdd.n223 vdd.n222 2.29662
R1769 vdd.n233 vdd.n0 2.29643
R1770 vdd.n171 vdd.n170 2.29594
R1771 vdd.n110 vdd.n28 2.29594
R1772 vdd.n82 vdd.n81 2.29594
R1773 vdd.n199 vdd.n2 2.29594
R1774 vdd.n227 vdd 1.88073
R1775 vdd.n168 vdd.n167 1.84013
R1776 vdd.n113 vdd.n111 1.84013
R1777 vdd.n79 vdd.n78 1.84013
R1778 vdd.n202 vdd.n200 1.84013
R1779 vdd.n49 vdd.n44 1.67304
R1780 vdd.n96 vdd.n91 1.67304
R1781 vdd.n21 vdd.n16 1.67304
R1782 vdd.n185 vdd.n181 1.67304
R1783 vdd.n78 vdd.n33 1.09272
R1784 vdd.n113 vdd.n112 1.09272
R1785 vdd.n167 vdd.n5 1.09272
R1786 vdd.n202 vdd.n201 1.09272
R1787 vdd.n57 vdd.n56 0.863992
R1788 vdd.n87 vdd.n86 0.863992
R1789 vdd.n146 vdd.n145 0.863992
R1790 vdd.n176 vdd.n175 0.863992
R1791 vdd.n52 vdd.n51 0.820933
R1792 vdd.n99 vdd.n98 0.820933
R1793 vdd.n24 vdd.n23 0.820933
R1794 vdd.n188 vdd.n187 0.820933
R1795 vdd.n170 vdd.n168 0.79957
R1796 vdd.n111 vdd.n110 0.79957
R1797 vdd.n81 vdd.n79 0.79957
R1798 vdd.n200 vdd.n199 0.79957
R1799 vdd.n225 vdd.n3 0.467369
R1800 vdd.n140 vdd.n139 0.467369
R1801 vdd.n136 vdd.n31 0.467369
R1802 vdd.n231 vdd.n230 0.467369
R1803 vdd.n56 vdd.n55 0.305262
R1804 vdd.n60 vdd.n59 0.305262
R1805 vdd.n86 vdd.n32 0.305262
R1806 vdd.n129 vdd.n128 0.305262
R1807 vdd.n145 vdd.n144 0.305262
R1808 vdd.n149 vdd.n148 0.305262
R1809 vdd.n175 vdd.n4 0.305262
R1810 vdd.n218 vdd.n217 0.305262
R1811 vdd.n201 vdd.n1 0.294492
R1812 vdd.n172 vdd.n5 0.294492
R1813 vdd.n112 vdd.n27 0.294492
R1814 vdd.n83 vdd.n33 0.294492
R1815 vdd.n44 vdd.n42 0.237984
R1816 vdd.n91 vdd.n89 0.237984
R1817 vdd.n16 vdd.n14 0.237984
R1818 vdd.n186 vdd.n185 0.237984
R1819 vdd.n201 vdd 0.234
R1820 vdd vdd.n5 0.234
R1821 vdd.n112 vdd 0.234
R1822 vdd vdd.n33 0.234
R1823 vdd.n133 vdd.n84 0.180551
R1824 vdd.n142 vdd.n141 0.180551
R1825 vdd.n222 vdd.n173 0.180551
R1826 vdd.n233 vdd.n232 0.179926
R1827 vdd vdd.n235 0.137535
R1828 vdd.n54 vdd.n53 0.120292
R1829 vdd.n61 vdd.n53 0.120292
R1830 vdd.n64 vdd.n63 0.120292
R1831 vdd.n64 vdd.n38 0.120292
R1832 vdd.n68 vdd.n38 0.120292
R1833 vdd.n69 vdd.n68 0.120292
R1834 vdd.n70 vdd.n35 0.120292
R1835 vdd.n74 vdd.n35 0.120292
R1836 vdd.n75 vdd.n74 0.120292
R1837 vdd.n76 vdd.n75 0.120292
R1838 vdd.n84 vdd.n83 0.120292
R1839 vdd.n132 vdd.n131 0.120292
R1840 vdd.n131 vdd.n85 0.120292
R1841 vdd.n125 vdd.n101 0.120292
R1842 vdd.n125 vdd.n124 0.120292
R1843 vdd.n124 vdd.n123 0.120292
R1844 vdd.n123 vdd.n104 0.120292
R1845 vdd.n118 vdd.n105 0.120292
R1846 vdd.n118 vdd.n117 0.120292
R1847 vdd.n117 vdd.n116 0.120292
R1848 vdd.n116 vdd.n108 0.120292
R1849 vdd.n141 vdd.n27 0.120292
R1850 vdd.n143 vdd.n25 0.120292
R1851 vdd.n150 vdd.n25 0.120292
R1852 vdd.n153 vdd.n152 0.120292
R1853 vdd.n153 vdd.n10 0.120292
R1854 vdd.n157 vdd.n10 0.120292
R1855 vdd.n158 vdd.n157 0.120292
R1856 vdd.n159 vdd.n7 0.120292
R1857 vdd.n163 vdd.n7 0.120292
R1858 vdd.n164 vdd.n163 0.120292
R1859 vdd.n165 vdd.n164 0.120292
R1860 vdd.n173 vdd.n172 0.120292
R1861 vdd.n221 vdd.n220 0.120292
R1862 vdd.n220 vdd.n174 0.120292
R1863 vdd.n214 vdd.n190 0.120292
R1864 vdd.n214 vdd.n213 0.120292
R1865 vdd.n213 vdd.n212 0.120292
R1866 vdd.n212 vdd.n193 0.120292
R1867 vdd.n207 vdd.n194 0.120292
R1868 vdd.n207 vdd.n206 0.120292
R1869 vdd.n206 vdd.n205 0.120292
R1870 vdd.n205 vdd.n197 0.120292
R1871 vdd.n232 vdd.n1 0.120292
R1872 vdd.n45 vdd.n44 0.0827222
R1873 vdd.n92 vdd.n91 0.0827222
R1874 vdd.n17 vdd.n16 0.0827222
R1875 vdd.n185 vdd.n184 0.0827222
R1876 vdd.n222 vdd 0.0826382
R1877 vdd vdd.n142 0.0826382
R1878 vdd.n133 vdd 0.0826382
R1879 vdd vdd.n233 0.0822696
R1880 vdd.n235 vdd 0.0720601
R1881 vdd.n54 vdd 0.0603958
R1882 vdd.n63 vdd 0.0603958
R1883 vdd vdd.n132 0.0603958
R1884 vdd.n101 vdd 0.0603958
R1885 vdd.n143 vdd 0.0603958
R1886 vdd.n152 vdd 0.0603958
R1887 vdd vdd.n221 0.0603958
R1888 vdd.n190 vdd 0.0603958
R1889 vdd.n43 vdd.n41 0.0536084
R1890 vdd.n90 vdd.n88 0.0536084
R1891 vdd.n15 vdd.n13 0.0536084
R1892 vdd.n180 vdd.n177 0.0536084
R1893 vdd.n70 vdd 0.0512812
R1894 vdd.n105 vdd 0.0512812
R1895 vdd.n159 vdd 0.0512812
R1896 vdd.n194 vdd 0.0512812
R1897 vdd.n44 vdd.n43 0.0272435
R1898 vdd.n91 vdd.n90 0.0272435
R1899 vdd.n16 vdd.n15 0.0272435
R1900 vdd.n185 vdd.n180 0.0272435
R1901 vdd vdd.n69 0.0226354
R1902 vdd.n76 vdd 0.0226354
R1903 vdd vdd.n104 0.0226354
R1904 vdd vdd.n108 0.0226354
R1905 vdd vdd.n158 0.0226354
R1906 vdd.n165 vdd 0.0226354
R1907 vdd vdd.n193 0.0226354
R1908 vdd vdd.n197 0.0226354
R1909 vdd vdd.n62 0.0200312
R1910 vdd vdd.n100 0.0200312
R1911 vdd vdd.n151 0.0200312
R1912 vdd vdd.n189 0.0200312
R1913 vdd.n234 vdd 0.0200312
R1914 vdd.n234 vdd 0.0187292
R1915 vdd vdd.n234 0.0183571
R1916 vdd.n48 vdd.n47 0.00492753
R1917 vdd.n95 vdd.n94 0.00492753
R1918 vdd.n20 vdd.n19 0.00492753
R1919 vdd.n183 vdd.n182 0.00492753
R1920 vdd.n62 vdd.n61 0.00310417
R1921 vdd.n100 vdd.n85 0.00310417
R1922 vdd.n151 vdd.n150 0.00310417
R1923 vdd.n189 vdd.n174 0.00310417
R1924 vss.n89 vss.n88 125981
R1925 vss.n123 vss.n71 22047.2
R1926 vss.n73 vss.n71 11121.2
R1927 vss.n109 vss.n105 9913.74
R1928 vss.n117 vss.n113 9913.74
R1929 vss.n122 vss.n121 9913.74
R1930 vss.n100 vss.n97 9913.74
R1931 vss.n93 vss.n83 7616.15
R1932 vss.n111 vss.n78 6110.51
R1933 vss.n119 vss.n73 6110.51
R1934 vss.n103 vss.n83 6110.51
R1935 vss.n105 vss.n81 5290.03
R1936 vss.n113 vss.n76 5290.03
R1937 vss.n121 vss.n70 5290.03
R1938 vss.n97 vss.n96 5290.03
R1939 vss.n81 vss.n80 5156.76
R1940 vss.n76 vss.n75 5156.76
R1941 vss.n124 vss.n70 5156.76
R1942 vss.n96 vss.n84 5156.76
R1943 vss.n93 vss.n92 4867.84
R1944 vss.n78 vss.n73 3443.71
R1945 vss.n83 vss.n78 3443.71
R1946 vss.n119 vss.n118 2038.64
R1947 vss.n111 vss.n110 2038.64
R1948 vss.n103 vss.n102 2038.64
R1949 vss.n120 vss.n119 2015.03
R1950 vss.n112 vss.n111 2015.03
R1951 vss.n104 vss.n103 2015.03
R1952 vss.n123 vss.t104 1361.72
R1953 vss.n120 vss.t99 1361.72
R1954 vss.n118 vss.t46 1361.72
R1955 vss.n112 vss.t50 1361.72
R1956 vss.n110 vss.t37 1361.72
R1957 vss.n104 vss.t32 1361.72
R1958 vss.n102 vss.t81 1361.72
R1959 vss.t85 vss.n94 1361.72
R1960 vss.t100 vss.t104 928.802
R1961 vss.t105 vss.t100 928.802
R1962 vss.t101 vss.t105 928.802
R1963 vss.t107 vss.t101 928.802
R1964 vss.t98 vss.t102 928.802
R1965 vss.t106 vss.t98 928.802
R1966 vss.t103 vss.t106 928.802
R1967 vss.t99 vss.t103 928.802
R1968 vss.t52 vss.t46 928.802
R1969 vss.t49 vss.t52 928.802
R1970 vss.t53 vss.t49 928.802
R1971 vss.t47 vss.t53 928.802
R1972 vss.t51 vss.t44 928.802
R1973 vss.t48 vss.t51 928.802
R1974 vss.t45 vss.t48 928.802
R1975 vss.t50 vss.t45 928.802
R1976 vss.t33 vss.t37 928.802
R1977 vss.t38 vss.t33 928.802
R1978 vss.t34 vss.t38 928.802
R1979 vss.t30 vss.t34 928.802
R1980 vss.t31 vss.t35 928.802
R1981 vss.t29 vss.t31 928.802
R1982 vss.t36 vss.t29 928.802
R1983 vss.t32 vss.t36 928.802
R1984 vss.t76 vss.t81 928.802
R1985 vss.t83 vss.t76 928.802
R1986 vss.t80 vss.t83 928.802
R1987 vss.t77 vss.t80 928.802
R1988 vss.t84 vss.t78 928.802
R1989 vss.t78 vss.t82 928.802
R1990 vss.t82 vss.t79 928.802
R1991 vss.t79 vss.t85 928.802
R1992 vss.t21 vss 925.947
R1993 vss.t18 vss 925.947
R1994 vss.t9 vss 925.947
R1995 vss.t12 vss 925.947
R1996 vss vss.t21 794.673
R1997 vss vss.t18 794.673
R1998 vss vss.t9 794.673
R1999 vss vss.t12 794.673
R2000 vss.n100 vss.n99 592.154
R2001 vss.n123 vss.n122 585
R2002 vss.n118 vss.n117 585
R2003 vss.n110 vss.n109 585
R2004 vss.n86 vss.n85 538.854
R2005 vss.t0 vss.n91 514.444
R2006 vss.n72 vss.t107 464.401
R2007 vss.t102 vss.n72 464.401
R2008 vss.n77 vss.t47 464.401
R2009 vss.t44 vss.n77 464.401
R2010 vss.n82 vss.t30 464.401
R2011 vss.t35 vss.n82 464.401
R2012 vss.n95 vss.t77 464.401
R2013 vss.n95 vss.t84 464.401
R2014 vss.n94 vss.n93 401.432
R2015 vss.t15 vss 391.476
R2016 vss.t6 vss 391.476
R2017 vss.t3 vss 391.476
R2018 vss.t151 vss 311.774
R2019 vss.t120 vss 311.774
R2020 vss.t145 vss 311.774
R2021 vss.t122 vss 311.774
R2022 vss.t54 vss 295.365
R2023 vss.t130 vss 295.365
R2024 vss.t86 vss 295.365
R2025 vss.t135 vss 295.365
R2026 vss.n87 vss 292.164
R2027 vss.n89 vss 292.164
R2028 vss.n91 vss.n90 279.687
R2029 vss.n92 vss 258.589
R2030 vss vss.t0 255.514
R2031 vss vss.t15 255.514
R2032 vss vss.t6 255.514
R2033 vss vss.t3 255.514
R2034 vss.n92 vss 253.714
R2035 vss.n91 vss 253.714
R2036 vss.n88 vss.n71 218.686
R2037 vss.t155 vss.t151 196.911
R2038 vss.t149 vss.t155 196.911
R2039 vss.t153 vss.t149 196.911
R2040 vss.t88 vss.t54 196.911
R2041 vss.t56 vss.t88 196.911
R2042 vss.t90 vss.t56 196.911
R2043 vss.t118 vss.t120 196.911
R2044 vss.t114 vss.t118 196.911
R2045 vss.t116 vss.t114 196.911
R2046 vss.t159 vss.t130 196.911
R2047 vss.t58 vss.t159 196.911
R2048 vss.t139 vss.t58 196.911
R2049 vss.t143 vss.t145 196.911
R2050 vss.t147 vss.t143 196.911
R2051 vss.t141 vss.t147 196.911
R2052 vss.t137 vss.t86 196.911
R2053 vss.t157 vss.t137 196.911
R2054 vss.t24 vss.t157 196.911
R2055 vss.t126 vss.t122 196.911
R2056 vss.t124 vss.t126 196.911
R2057 vss.t128 vss.t124 196.911
R2058 vss.t62 vss.t135 196.911
R2059 vss.t39 vss.t62 196.911
R2060 vss.t60 vss.t39 196.911
R2061 vss.n6 vss.t61 193.933
R2062 vss.n281 vss.t129 193.933
R2063 vss.n146 vss.t154 193.933
R2064 vss.n57 vss.t91 193.933
R2065 vss.n191 vss.t117 193.933
R2066 vss.n40 vss.t140 193.933
R2067 vss.n236 vss.t142 193.933
R2068 vss.n23 vss.t25 193.933
R2069 vss.n9 vss.t136 192.982
R2070 vss.n275 vss.t123 192.982
R2071 vss.n140 vss.t152 192.982
R2072 vss.n60 vss.t55 192.982
R2073 vss.n185 vss.t121 192.982
R2074 vss.n43 vss.t131 192.982
R2075 vss.n230 vss.t146 192.982
R2076 vss.n26 vss.t87 192.982
R2077 vss.n88 vss.n87 192.744
R2078 vss.n135 vss.t189 183.082
R2079 vss.n180 vss.t184 183.082
R2080 vss.n225 vss.t187 183.082
R2081 vss.n270 vss.t188 183.082
R2082 vss vss.t153 175.812
R2083 vss vss.t90 175.812
R2084 vss vss.t116 175.812
R2085 vss vss.t139 175.812
R2086 vss vss.t141 175.812
R2087 vss vss.t24 175.812
R2088 vss vss.t128 175.812
R2089 vss vss.t60 175.812
R2090 vss.n303 vss.n302 124.692
R2091 vss.n258 vss.n257 124.692
R2092 vss.n213 vss.n212 124.692
R2093 vss.n168 vss.n167 124.692
R2094 vss.n13 vss.t5 121.956
R2095 vss.n15 vss.t4 121.956
R2096 vss.n292 vss.t13 121.956
R2097 vss.n3 vss.t14 121.956
R2098 vss.n18 vss.t11 121.956
R2099 vss.n247 vss.t10 121.956
R2100 vss.n30 vss.t8 121.956
R2101 vss.n32 vss.t7 121.956
R2102 vss.n35 vss.t20 121.956
R2103 vss.n202 vss.t19 121.956
R2104 vss.n47 vss.t17 121.956
R2105 vss.n49 vss.t16 121.956
R2106 vss.n52 vss.t23 121.956
R2107 vss.n157 vss.t22 121.956
R2108 vss.n64 vss.t2 121.956
R2109 vss.n66 vss.t1 121.956
R2110 vss.n241 vss.n25 114.713
R2111 vss.n234 vss.n28 114.713
R2112 vss.n196 vss.n42 114.713
R2113 vss.n189 vss.n45 114.713
R2114 vss.n151 vss.n59 114.713
R2115 vss.n144 vss.n62 114.713
R2116 vss.n279 vss.n11 114.713
R2117 vss.n286 vss.n8 114.713
R2118 vss.n301 vss.n300 114.398
R2119 vss.n256 vss.n255 114.398
R2120 vss.n211 vss.n210 114.398
R2121 vss.n166 vss.n165 114.398
R2122 vss.n109 vss.n108 104.882
R2123 vss.n117 vss.n116 104.882
R2124 vss.n122 vss.n68 104.882
R2125 vss.n101 vss.n100 104.654
R2126 vss.n302 vss.n2 76.0005
R2127 vss.n167 vss.n54 76.0005
R2128 vss.n212 vss.n37 76.0005
R2129 vss.n257 vss.n20 76.0005
R2130 vss.n87 vss.t26 41.0057
R2131 vss.n286 vss.n285 34.6358
R2132 vss.n287 vss.n286 34.6358
R2133 vss.n279 vss.n12 34.6358
R2134 vss.n280 vss.n279 34.6358
R2135 vss.n144 vss.n63 34.6358
R2136 vss.n145 vss.n144 34.6358
R2137 vss.n151 vss.n150 34.6358
R2138 vss.n152 vss.n151 34.6358
R2139 vss.n189 vss.n46 34.6358
R2140 vss.n190 vss.n189 34.6358
R2141 vss.n196 vss.n195 34.6358
R2142 vss.n197 vss.n196 34.6358
R2143 vss.n234 vss.n29 34.6358
R2144 vss.n235 vss.n234 34.6358
R2145 vss.n241 vss.n240 34.6358
R2146 vss.n242 vss.n241 34.6358
R2147 vss.n301 vss.t185 34.2973
R2148 vss.n256 vss.t186 34.2973
R2149 vss.n211 vss.t183 34.2973
R2150 vss.n166 vss.t182 34.2973
R2151 vss.n107 vss.n106 33.1064
R2152 vss.n115 vss.n114 33.1064
R2153 vss.n126 vss.n125 33.1064
R2154 vss.n99 vss.n98 33.1064
R2155 vss.n128 vss 29.9299
R2156 vss.n308 vss.n0 29.1367
R2157 vss vss.t161 27.9221
R2158 vss vss.t70 27.6987
R2159 vss vss.t170 27.6987
R2160 vss vss.t95 27.6987
R2161 vss vss.t64 27.6987
R2162 vss vss.t176 27.6987
R2163 vss vss.t179 27.4754
R2164 vss vss.t92 27.4754
R2165 vss vss.n89 26.1071
R2166 vss.n25 vss.t138 24.9236
R2167 vss.n25 vss.t158 24.9236
R2168 vss.n28 vss.t144 24.9236
R2169 vss.n28 vss.t148 24.9236
R2170 vss.n42 vss.t160 24.9236
R2171 vss.n42 vss.t59 24.9236
R2172 vss.n45 vss.t119 24.9236
R2173 vss.n45 vss.t115 24.9236
R2174 vss.n59 vss.t89 24.9236
R2175 vss.n59 vss.t57 24.9236
R2176 vss.n62 vss.t156 24.9236
R2177 vss.n62 vss.t150 24.9236
R2178 vss.n11 vss.t127 24.9236
R2179 vss.n11 vss.t125 24.9236
R2180 vss.n8 vss.t63 24.9236
R2181 vss.n8 vss.t40 24.9236
R2182 vss.n285 vss.n9 22.2123
R2183 vss.n287 vss.n6 22.2123
R2184 vss.n275 vss.n12 22.2123
R2185 vss.n281 vss.n280 22.2123
R2186 vss.n140 vss.n63 22.2123
R2187 vss.n146 vss.n145 22.2123
R2188 vss.n150 vss.n60 22.2123
R2189 vss.n152 vss.n57 22.2123
R2190 vss.n185 vss.n46 22.2123
R2191 vss.n191 vss.n190 22.2123
R2192 vss.n195 vss.n43 22.2123
R2193 vss.n197 vss.n40 22.2123
R2194 vss.n230 vss.n29 22.2123
R2195 vss.n236 vss.n235 22.2123
R2196 vss.n240 vss.n26 22.2123
R2197 vss.n242 vss.n23 22.2123
R2198 vss.n275 vss.n274 19.3355
R2199 vss.n140 vss.n139 19.3355
R2200 vss.n185 vss.n184 19.3355
R2201 vss.n230 vss.n229 19.3355
R2202 vss.t26 vss.t41 18.7638
R2203 vss.t70 vss.t73 18.7638
R2204 vss.t179 vss.t108 18.7638
R2205 vss.t170 vss.t173 18.7638
R2206 vss.t95 vss.t167 18.7638
R2207 vss.t161 vss.t164 18.7638
R2208 vss.t64 vss.t132 18.7638
R2209 vss.t92 vss.t67 18.7638
R2210 vss.t176 vss.t111 18.7638
R2211 vss.n281 vss.n9 18.0711
R2212 vss.n146 vss.n60 18.0711
R2213 vss.n191 vss.n43 18.0711
R2214 vss.n236 vss.n26 18.0711
R2215 vss.n291 vss.n6 17.4103
R2216 vss.n156 vss.n57 17.4103
R2217 vss.n201 vss.n40 17.4103
R2218 vss.n246 vss.n23 17.4103
R2219 vss.n173 vss.n172 16.0891
R2220 vss.n218 vss.n217 16.0891
R2221 vss.n263 vss.n262 16.0891
R2222 vss.t41 vss 14.9665
R2223 vss.t73 vss 14.9665
R2224 vss.t108 vss 14.9665
R2225 vss.t173 vss 14.9665
R2226 vss.t167 vss 14.9665
R2227 vss.t164 vss 14.9665
R2228 vss.t132 vss 14.9665
R2229 vss.t111 vss 14.9665
R2230 vss.n90 vss.t67 9.82891
R2231 vss.n227 vss.n226 9.3005
R2232 vss.n182 vss.n181 9.3005
R2233 vss.n137 vss.n136 9.3005
R2234 vss.n134 vss.n65 9.3005
R2235 vss.n179 vss.n48 9.3005
R2236 vss.n224 vss.n31 9.3005
R2237 vss.n269 vss.n14 9.3005
R2238 vss.n272 vss.n271 9.3005
R2239 vss.n266 vss.n265 9.0005
R2240 vss.n267 vss.n266 9.0005
R2241 vss.n268 vss.n267 9.0005
R2242 vss.n222 vss.n221 9.0005
R2243 vss.n223 vss.n222 9.0005
R2244 vss.n177 vss.n176 9.0005
R2245 vss.n178 vss.n177 9.0005
R2246 vss.n132 vss.n131 9.0005
R2247 vss.n133 vss.n132 9.0005
R2248 vss.n34 vss.n33 9.0005
R2249 vss.n51 vss.n50 9.0005
R2250 vss.n127 vss.n67 9.0005
R2251 vss.n106 vss.n80 8.19978
R2252 vss.n114 vss.n75 8.19978
R2253 vss.n125 vss.n124 8.19978
R2254 vss.n98 vss.n84 8.19978
R2255 vss.n294 vss.n293 6.26433
R2256 vss.n294 vss.n4 6.26433
R2257 vss.n159 vss.n158 6.26433
R2258 vss.n159 vss.n55 6.26433
R2259 vss.n204 vss.n203 6.26433
R2260 vss.n204 vss.n38 6.26433
R2261 vss.n249 vss.n248 6.26433
R2262 vss.n249 vss.n21 6.26433
R2263 vss.n293 vss.n292 5.85582
R2264 vss.n158 vss.n157 5.85582
R2265 vss.n203 vss.n202 5.85582
R2266 vss.n248 vss.n247 5.85582
R2267 vss.n298 vss.n4 5.65809
R2268 vss.n163 vss.n55 5.65809
R2269 vss.n208 vss.n38 5.65809
R2270 vss.n253 vss.n21 5.65809
R2271 vss.n90 vss 5.13808
R2272 vss.n133 vss.n66 5.0092
R2273 vss.n178 vss.n49 5.0092
R2274 vss.n223 vss.n32 5.0092
R2275 vss.n268 vss.n15 5.0092
R2276 vss.n302 vss.n301 4.85762
R2277 vss.n257 vss.n256 4.85762
R2278 vss.n212 vss.n211 4.85762
R2279 vss.n167 vss.n166 4.85762
R2280 vss.n231 vss.n230 4.6505
R2281 vss.n237 vss.n236 4.6505
R2282 vss.n238 vss.n26 4.6505
R2283 vss.n244 vss.n23 4.6505
R2284 vss.n186 vss.n185 4.6505
R2285 vss.n192 vss.n191 4.6505
R2286 vss.n193 vss.n43 4.6505
R2287 vss.n199 vss.n40 4.6505
R2288 vss.n141 vss.n140 4.6505
R2289 vss.n147 vss.n146 4.6505
R2290 vss.n148 vss.n60 4.6505
R2291 vss.n154 vss.n57 4.6505
R2292 vss.n289 vss.n6 4.6505
R2293 vss.n283 vss.n9 4.6505
R2294 vss.n282 vss.n281 4.6505
R2295 vss.n276 vss.n275 4.6505
R2296 vss.n306 vss.n0 4.6505
R2297 vss.n305 vss.n304 4.6505
R2298 vss.n299 vss.n1 4.6505
R2299 vss.n298 vss.n297 4.6505
R2300 vss.n296 vss.n4 4.6505
R2301 vss.n295 vss.n294 4.6505
R2302 vss.n293 vss.n5 4.6505
R2303 vss.n291 vss.n290 4.6505
R2304 vss.n288 vss.n287 4.6505
R2305 vss.n286 vss.n7 4.6505
R2306 vss.n285 vss.n284 4.6505
R2307 vss.n280 vss.n10 4.6505
R2308 vss.n279 vss.n278 4.6505
R2309 vss.n277 vss.n12 4.6505
R2310 vss.n274 vss.n273 4.6505
R2311 vss.n129 vss.n128 4.6505
R2312 vss.n139 vss.n138 4.6505
R2313 vss.n142 vss.n63 4.6505
R2314 vss.n144 vss.n143 4.6505
R2315 vss.n145 vss.n61 4.6505
R2316 vss.n150 vss.n149 4.6505
R2317 vss.n151 vss.n58 4.6505
R2318 vss.n153 vss.n152 4.6505
R2319 vss.n156 vss.n155 4.6505
R2320 vss.n158 vss.n56 4.6505
R2321 vss.n160 vss.n159 4.6505
R2322 vss.n161 vss.n55 4.6505
R2323 vss.n163 vss.n162 4.6505
R2324 vss.n164 vss.n53 4.6505
R2325 vss.n170 vss.n169 4.6505
R2326 vss.n172 vss.n171 4.6505
R2327 vss.n174 vss.n173 4.6505
R2328 vss.n184 vss.n183 4.6505
R2329 vss.n187 vss.n46 4.6505
R2330 vss.n189 vss.n188 4.6505
R2331 vss.n190 vss.n44 4.6505
R2332 vss.n195 vss.n194 4.6505
R2333 vss.n196 vss.n41 4.6505
R2334 vss.n198 vss.n197 4.6505
R2335 vss.n201 vss.n200 4.6505
R2336 vss.n203 vss.n39 4.6505
R2337 vss.n205 vss.n204 4.6505
R2338 vss.n206 vss.n38 4.6505
R2339 vss.n208 vss.n207 4.6505
R2340 vss.n209 vss.n36 4.6505
R2341 vss.n215 vss.n214 4.6505
R2342 vss.n217 vss.n216 4.6505
R2343 vss.n219 vss.n218 4.6505
R2344 vss.n229 vss.n228 4.6505
R2345 vss.n232 vss.n29 4.6505
R2346 vss.n234 vss.n233 4.6505
R2347 vss.n235 vss.n27 4.6505
R2348 vss.n240 vss.n239 4.6505
R2349 vss.n241 vss.n24 4.6505
R2350 vss.n243 vss.n242 4.6505
R2351 vss.n246 vss.n245 4.6505
R2352 vss.n248 vss.n22 4.6505
R2353 vss.n250 vss.n249 4.6505
R2354 vss.n251 vss.n21 4.6505
R2355 vss.n253 vss.n252 4.6505
R2356 vss.n254 vss.n19 4.6505
R2357 vss.n260 vss.n259 4.6505
R2358 vss.n262 vss.n261 4.6505
R2359 vss.n264 vss.n263 4.6505
R2360 vss.n136 vss.n135 4.5918
R2361 vss.n181 vss.n180 4.5918
R2362 vss.n226 vss.n225 4.5918
R2363 vss.n271 vss.n270 4.5918
R2364 vss vss.n17 3.61567
R2365 vss vss.n34 3.58168
R2366 vss vss.n51 3.58168
R2367 vss.n127 vss 3.58168
R2368 vss.n300 vss.n299 3.50735
R2369 vss.n165 vss.n164 3.50735
R2370 vss.n210 vss.n209 3.50735
R2371 vss.n255 vss.n254 3.50735
R2372 vss.n304 vss.n2 3.2005
R2373 vss.n169 vss.n54 3.2005
R2374 vss.n214 vss.n37 3.2005
R2375 vss.n259 vss.n20 3.2005
R2376 vss.n131 vss.n130 3.00723
R2377 vss.n176 vss.n175 3.00723
R2378 vss.n221 vss.n220 3.00723
R2379 vss.n17 vss.n16 2.99647
R2380 vss.n303 vss.n3 2.63064
R2381 vss.n168 vss.n52 2.63064
R2382 vss.n213 vss.n35 2.63064
R2383 vss.n258 vss.n18 2.63064
R2384 vss.n135 vss.n64 1.18311
R2385 vss.n180 vss.n47 1.18311
R2386 vss.n225 vss.n30 1.18311
R2387 vss.n270 vss.n13 1.18311
R2388 vss.n304 vss.n303 1.14023
R2389 vss.n169 vss.n168 1.14023
R2390 vss.n214 vss.n213 1.14023
R2391 vss.n259 vss.n258 1.14023
R2392 vss.n134 vss.n133 0.974413
R2393 vss.n179 vss.n178 0.974413
R2394 vss.n224 vss.n223 0.974413
R2395 vss.n269 vss.n268 0.974413
R2396 vss.n299 vss.n2 0.833377
R2397 vss.n164 vss.n54 0.833377
R2398 vss.n209 vss.n37 0.833377
R2399 vss.n254 vss.n20 0.833377
R2400 vss.n107 vss 0.704167
R2401 vss.n115 vss 0.704167
R2402 vss vss.n126 0.704167
R2403 vss.n99 vss 0.700242
R2404 vss.n300 vss.n298 0.526527
R2405 vss.n165 vss.n163 0.526527
R2406 vss.n210 vss.n208 0.526527
R2407 vss.n255 vss.n253 0.526527
R2408 vss.n128 vss.n66 0.417891
R2409 vss.n139 vss.n64 0.417891
R2410 vss.n173 vss.n49 0.417891
R2411 vss.n184 vss.n47 0.417891
R2412 vss.n218 vss.n32 0.417891
R2413 vss.n229 vss.n30 0.417891
R2414 vss.n263 vss.n15 0.417891
R2415 vss.n274 vss.n13 0.417891
R2416 vss.n292 vss.n291 0.409011
R2417 vss.n157 vss.n156 0.409011
R2418 vss.n202 vss.n201 0.409011
R2419 vss.n247 vss.n246 0.409011
R2420 vss.n3 vss.n0 0.263514
R2421 vss.n172 vss.n52 0.263514
R2422 vss.n217 vss.n35 0.263514
R2423 vss.n262 vss.n18 0.263514
R2424 vss.n125 vss.n69 0.260881
R2425 vss.n114 vss.n74 0.260881
R2426 vss.n106 vss.n79 0.260881
R2427 vss.n136 vss.n134 0.209196
R2428 vss.n181 vss.n179 0.209196
R2429 vss.n226 vss.n224 0.209196
R2430 vss.n271 vss.n269 0.209196
R2431 vss.n307 vss 0.195812
R2432 vss.n124 vss.n123 0.172761
R2433 vss.n118 vss.n75 0.172761
R2434 vss.n110 vss.n80 0.172761
R2435 vss.n102 vss.n84 0.172761
R2436 vss vss.n308 0.140087
R2437 vss.n102 vss.n85 0.134398
R2438 vss.n98 vss.n85 0.126534
R2439 vss.n142 vss.n141 0.120292
R2440 vss.n143 vss.n142 0.120292
R2441 vss.n143 vss.n61 0.120292
R2442 vss.n147 vss.n61 0.120292
R2443 vss.n149 vss.n148 0.120292
R2444 vss.n149 vss.n58 0.120292
R2445 vss.n153 vss.n58 0.120292
R2446 vss.n154 vss.n153 0.120292
R2447 vss.n155 vss.n56 0.120292
R2448 vss.n160 vss.n56 0.120292
R2449 vss.n161 vss.n160 0.120292
R2450 vss.n162 vss.n161 0.120292
R2451 vss.n162 vss.n53 0.120292
R2452 vss.n170 vss.n53 0.120292
R2453 vss.n171 vss.n170 0.120292
R2454 vss.n187 vss.n186 0.120292
R2455 vss.n188 vss.n187 0.120292
R2456 vss.n188 vss.n44 0.120292
R2457 vss.n192 vss.n44 0.120292
R2458 vss.n194 vss.n193 0.120292
R2459 vss.n194 vss.n41 0.120292
R2460 vss.n198 vss.n41 0.120292
R2461 vss.n199 vss.n198 0.120292
R2462 vss.n200 vss.n39 0.120292
R2463 vss.n205 vss.n39 0.120292
R2464 vss.n206 vss.n205 0.120292
R2465 vss.n207 vss.n206 0.120292
R2466 vss.n207 vss.n36 0.120292
R2467 vss.n215 vss.n36 0.120292
R2468 vss.n216 vss.n215 0.120292
R2469 vss.n232 vss.n231 0.120292
R2470 vss.n233 vss.n232 0.120292
R2471 vss.n233 vss.n27 0.120292
R2472 vss.n237 vss.n27 0.120292
R2473 vss.n239 vss.n238 0.120292
R2474 vss.n239 vss.n24 0.120292
R2475 vss.n243 vss.n24 0.120292
R2476 vss.n244 vss.n243 0.120292
R2477 vss.n245 vss.n22 0.120292
R2478 vss.n250 vss.n22 0.120292
R2479 vss.n251 vss.n250 0.120292
R2480 vss.n252 vss.n251 0.120292
R2481 vss.n252 vss.n19 0.120292
R2482 vss.n260 vss.n19 0.120292
R2483 vss.n261 vss.n260 0.120292
R2484 vss.n277 vss.n276 0.120292
R2485 vss.n278 vss.n277 0.120292
R2486 vss.n278 vss.n10 0.120292
R2487 vss.n282 vss.n10 0.120292
R2488 vss.n284 vss.n283 0.120292
R2489 vss.n284 vss.n7 0.120292
R2490 vss.n288 vss.n7 0.120292
R2491 vss.n289 vss.n288 0.120292
R2492 vss.n290 vss.n5 0.120292
R2493 vss.n295 vss.n5 0.120292
R2494 vss.n296 vss.n295 0.120292
R2495 vss.n297 vss.n296 0.120292
R2496 vss.n297 vss.n1 0.120292
R2497 vss.n305 vss.n1 0.120292
R2498 vss.n306 vss.n305 0.120292
R2499 vss.n138 vss.n137 0.116385
R2500 vss.n183 vss.n182 0.116385
R2501 vss.n228 vss.n227 0.116385
R2502 vss.n273 vss.n272 0.116385
R2503 vss.n108 vss.n79 0.0856819
R2504 vss.n116 vss.n74 0.0856819
R2505 vss.n69 vss.n68 0.0856819
R2506 vss.n99 vss.n86 0.0720385
R2507 vss.n130 vss.n129 0.0713087
R2508 vss.n175 vss.n174 0.0713087
R2509 vss.n220 vss.n219 0.0713087
R2510 vss.n265 vss.n264 0.0682083
R2511 vss.n121 vss.n120 0.067449
R2512 vss.n113 vss.n112 0.067449
R2513 vss.n105 vss.n104 0.067449
R2514 vss.n97 vss.n94 0.067449
R2515 vss.n129 vss 0.0603958
R2516 vss.n141 vss 0.0603958
R2517 vss.n174 vss 0.0603958
R2518 vss.n186 vss 0.0603958
R2519 vss.n219 vss 0.0603958
R2520 vss.n231 vss 0.0603958
R2521 vss.n264 vss 0.0603958
R2522 vss.n276 vss 0.0603958
R2523 vss.n108 vss.n107 0.0598606
R2524 vss.n116 vss.n115 0.0598606
R2525 vss.n126 vss.n68 0.0598606
R2526 vss.n102 vss.n101 0.0597334
R2527 vss.n155 vss 0.0577917
R2528 vss.n200 vss 0.0577917
R2529 vss.n245 vss 0.0577917
R2530 vss.n290 vss 0.0577917
R2531 vss.n148 vss 0.0512812
R2532 vss.n193 vss 0.0512812
R2533 vss.n238 vss 0.0512812
R2534 vss.n283 vss 0.0512812
R2535 vss.n221 vss.n34 0.0509808
R2536 vss.n176 vss.n51 0.0509808
R2537 vss.n131 vss.n127 0.0509808
R2538 vss.n307 vss 0.0447708
R2539 vss.n132 vss.n67 0.0304479
R2540 vss.n177 vss.n50 0.0304479
R2541 vss.n222 vss.n33 0.0304479
R2542 vss.n267 vss.n16 0.0304479
R2543 vss.n308 vss.n307 0.0286927
R2544 vss.n138 vss 0.0226354
R2545 vss vss.n147 0.0226354
R2546 vss vss.n154 0.0226354
R2547 vss.n171 vss 0.0226354
R2548 vss.n183 vss 0.0226354
R2549 vss vss.n192 0.0226354
R2550 vss vss.n199 0.0226354
R2551 vss.n216 vss 0.0226354
R2552 vss.n228 vss 0.0226354
R2553 vss vss.n237 0.0226354
R2554 vss vss.n244 0.0226354
R2555 vss.n261 vss 0.0226354
R2556 vss.n273 vss 0.0226354
R2557 vss vss.n282 0.0226354
R2558 vss vss.n289 0.0226354
R2559 vss vss.n306 0.0226354
R2560 vss.n132 vss.n65 0.0187292
R2561 vss.n177 vss.n48 0.0187292
R2562 vss.n222 vss.n31 0.0187292
R2563 vss.n267 vss.n14 0.0187292
R2564 vss.n266 vss.n17 0.0178015
R2565 vss.n72 vss.n70 0.0145006
R2566 vss.n77 vss.n76 0.0145006
R2567 vss.n82 vss.n81 0.0145006
R2568 vss.n96 vss.n95 0.0145006
R2569 vss.n101 vss.n86 0.0137979
R2570 vss.n137 vss.n65 0.00440625
R2571 vss.n182 vss.n48 0.00440625
R2572 vss.n227 vss.n31 0.00440625
R2573 vss.n265 vss.n16 0.00440625
R2574 vss.n272 vss.n14 0.00440625
R2575 vss.n130 vss.n67 0.00230479
R2576 vss.n175 vss.n50 0.00230479
R2577 vss.n220 vss.n33 0.00230479
R2578 vss.n123 vss.n69 0.00101777
R2579 vss.n118 vss.n74 0.00101777
R2580 vss.n110 vss.n79 0.00101777
R2581 sample.n64 sample.t12 212.081
R2582 sample.n66 sample.t3 212.081
R2583 sample.n63 sample.t16 212.081
R2584 sample.n71 sample.t28 212.081
R2585 sample.n45 sample.t23 212.081
R2586 sample.n47 sample.t5 212.081
R2587 sample.n44 sample.t25 212.081
R2588 sample.n52 sample.t15 212.081
R2589 sample.n26 sample.t1 212.081
R2590 sample.n28 sample.t13 212.081
R2591 sample.n25 sample.t4 212.081
R2592 sample.n33 sample.t17 212.081
R2593 sample.n5 sample.t9 212.081
R2594 sample.n7 sample.t24 212.081
R2595 sample.n4 sample.t6 212.081
R2596 sample.n12 sample.t26 212.081
R2597 sample.n64 sample.t29 139.78
R2598 sample.n66 sample.t19 139.78
R2599 sample.n63 sample.t0 139.78
R2600 sample.n71 sample.t14 139.78
R2601 sample.n45 sample.t7 139.78
R2602 sample.n47 sample.t21 139.78
R2603 sample.n44 sample.t10 139.78
R2604 sample.n52 sample.t31 139.78
R2605 sample.n26 sample.t18 139.78
R2606 sample.n28 sample.t30 139.78
R2607 sample.n25 sample.t20 139.78
R2608 sample.n33 sample.t2 139.78
R2609 sample.n5 sample.t27 139.78
R2610 sample.n7 sample.t8 139.78
R2611 sample.n4 sample.t22 139.78
R2612 sample.n12 sample.t11 139.78
R2613 sample.n65 sample 78.3045
R2614 sample.n46 sample 78.3045
R2615 sample.n27 sample 78.3045
R2616 sample.n6 sample 78.3045
R2617 sample.n68 sample.n67 76.0005
R2618 sample.n70 sample.n69 76.0005
R2619 sample.n49 sample.n48 76.0005
R2620 sample.n51 sample.n50 76.0005
R2621 sample.n30 sample.n29 76.0005
R2622 sample.n32 sample.n31 76.0005
R2623 sample.n9 sample.n8 76.0005
R2624 sample.n11 sample.n10 76.0005
R2625 sample.n72 sample.n71 44.8017
R2626 sample.n53 sample.n52 44.8017
R2627 sample.n34 sample.n33 44.8017
R2628 sample.n13 sample.n12 44.8017
R2629 sample.n65 sample.n64 30.6732
R2630 sample.n66 sample.n65 30.6732
R2631 sample.n67 sample.n66 30.6732
R2632 sample.n67 sample.n63 30.6732
R2633 sample.n70 sample.n63 30.6732
R2634 sample.n71 sample.n70 30.6732
R2635 sample.n46 sample.n45 30.6732
R2636 sample.n47 sample.n46 30.6732
R2637 sample.n48 sample.n47 30.6732
R2638 sample.n48 sample.n44 30.6732
R2639 sample.n51 sample.n44 30.6732
R2640 sample.n52 sample.n51 30.6732
R2641 sample.n27 sample.n26 30.6732
R2642 sample.n28 sample.n27 30.6732
R2643 sample.n29 sample.n28 30.6732
R2644 sample.n29 sample.n25 30.6732
R2645 sample.n32 sample.n25 30.6732
R2646 sample.n33 sample.n32 30.6732
R2647 sample.n6 sample.n5 30.6732
R2648 sample.n7 sample.n6 30.6732
R2649 sample.n8 sample.n7 30.6732
R2650 sample.n8 sample.n4 30.6732
R2651 sample.n11 sample.n4 30.6732
R2652 sample.n12 sample.n11 30.6732
R2653 sample.n68 sample 19.2005
R2654 sample.n49 sample 19.2005
R2655 sample.n30 sample 19.2005
R2656 sample.n9 sample 19.2005
R2657 sample.n69 sample 17.1525
R2658 sample.n50 sample 17.1525
R2659 sample.n31 sample 17.1525
R2660 sample.n10 sample 17.1525
R2661 sample sample.n60 12.2885
R2662 sample sample.n41 12.2885
R2663 sample sample.n22 12.2885
R2664 sample sample.n2 12.2885
R2665 sample.n60 sample.n58 9.34456
R2666 sample.n41 sample.n39 9.34456
R2667 sample.n22 sample.n20 9.34456
R2668 sample.n72 sample.n59 9.3005
R2669 sample.n62 sample.n61 9.3005
R2670 sample.n53 sample.n40 9.3005
R2671 sample.n43 sample.n42 9.3005
R2672 sample.n34 sample.n21 9.3005
R2673 sample.n24 sample.n23 9.3005
R2674 sample.n61 sample.n57 9.01011
R2675 sample.n42 sample.n38 9.01011
R2676 sample.n23 sample.n19 9.01011
R2677 sample.n69 sample 6.4005
R2678 sample.n50 sample 6.4005
R2679 sample.n31 sample 6.4005
R2680 sample.n10 sample 6.4005
R2681 sample.n76 sample 5.80233
R2682 sample.n77 sample 5.80233
R2683 sample.n78 sample 5.80233
R2684 sample.n73 sample.n60 4.6085
R2685 sample.n72 sample.n62 4.6085
R2686 sample.n54 sample.n41 4.6085
R2687 sample.n53 sample.n43 4.6085
R2688 sample.n35 sample.n22 4.6085
R2689 sample.n34 sample.n24 4.6085
R2690 sample.n14 sample.n2 4.6085
R2691 sample.n13 sample.n3 4.6085
R2692 sample.n75 sample.n74 4.501
R2693 sample.n56 sample.n55 4.501
R2694 sample.n37 sample.n36 4.501
R2695 sample sample.n68 4.3525
R2696 sample sample.n49 4.3525
R2697 sample sample.n30 4.3525
R2698 sample sample.n9 4.3525
R2699 sample.n62 sample 1.7925
R2700 sample.n43 sample 1.7925
R2701 sample.n24 sample 1.7925
R2702 sample.n3 sample 1.7925
R2703 sample sample.n75 0.958647
R2704 sample.n78 sample.n18 0.925142
R2705 sample.n76 sample.n56 0.897671
R2706 sample.n77 sample.n37 0.897671
R2707 sample.n73 sample.n72 0.2565
R2708 sample.n54 sample.n53 0.2565
R2709 sample.n35 sample.n34 0.2565
R2710 sample.n14 sample.n13 0.2565
R2711 sample sample.n76 0.0614756
R2712 sample sample.n77 0.0614756
R2713 sample sample.n78 0.0614756
R2714 sample.n61 sample.n59 0.0437692
R2715 sample.n42 sample.n40 0.0437692
R2716 sample.n23 sample.n21 0.0437692
R2717 sample.n17 sample.n1 0.0437692
R2718 sample.n16 sample.n15 0.0437692
R2719 sample.n75 sample.n57 0.0286442
R2720 sample.n56 sample.n38 0.0286442
R2721 sample.n37 sample.n19 0.0286442
R2722 sample.n74 sample.n59 0.00290385
R2723 sample.n55 sample.n40 0.00290385
R2724 sample.n36 sample.n21 0.00290385
R2725 sample.n17 sample.n16 0.00290385
R2726 sample.n58 sample.n57 0.00216539
R2727 sample.n39 sample.n38 0.00216539
R2728 sample.n20 sample.n19 0.00216539
R2729 sample.n18 sample.n17 0.00166462
R2730 sample.n74 sample.n58 0.0015031
R2731 sample.n55 sample.n39 0.0015031
R2732 sample.n36 sample.n20 0.0015031
R2733 sample.n74 sample.n73 0.0011688
R2734 sample.n55 sample.n54 0.0011688
R2735 sample.n36 sample.n35 0.0011688
R2736 sample.n17 sample.n14 0.0011688
R2737 sample.n18 sample.n0 0.00100408
R2738 ctl7.n3 ctl7.t0 212.081
R2739 ctl7.n2 ctl7.t2 212.081
R2740 ctl7.n3 ctl7.t1 139.78
R2741 ctl7.n2 ctl7.t3 139.78
R2742 ctl7.n3 ctl7.n2 61.346
R2743 ctl7.n5 ctl7.n3 38.5428
R2744 ctl7.n5 ctl7.n0 9.30881
R2745 ctl7.n6 ctl7.n5 9.3005
R2746 ctl7.n7 ctl7.n6 9.01417
R2747 ctl7.n4 ctl7 3.23067
R2748 ctl7.n5 ctl7.n4 1.2812
R2749 ctl7.n7 ctl7.n0 0.0569565
R2750 ctl7.n6 ctl7.n1 0.03175
R2751 ctl7 ctl7.n7 0.00771154
R2752 ctl7.n4 ctl7.n1 0.00147336
R2753 ctl7.n1 ctl7.n0 0.00100057
R2754 sky130_fd_sc_hd__inv_2_3.Y.n4 sky130_fd_sc_hd__inv_2_3.Y.n3 111.32
R2755 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_sc_hd__inv_2_3.Y.n0 50.4671
R2756 sky130_fd_sc_hd__inv_2_3.Y.n3 sky130_fd_sc_hd__inv_2_3.Y.t2 26.5955
R2757 sky130_fd_sc_hd__inv_2_3.Y.n3 sky130_fd_sc_hd__inv_2_3.Y.t4 26.5955
R2758 sky130_fd_sc_hd__inv_2_3.Y.n0 sky130_fd_sc_hd__inv_2_3.Y.t3 24.9236
R2759 sky130_fd_sc_hd__inv_2_3.Y.n0 sky130_fd_sc_hd__inv_2_3.Y.t5 24.9236
R2760 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_sc_hd__inv_2_3.Y.n2 13.3125
R2761 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_sc_hd__inv_2_3.Y.n1 11.2645
R2762 sky130_fd_sc_hd__inv_2_3.Y.n1 sky130_fd_sc_hd__inv_2_3.Y 6.1445
R2763 sky130_fd_sc_hd__inv_2_3.Y.n1 sky130_fd_sc_hd__inv_2_3.Y 4.65505
R2764 sky130_fd_sc_hd__inv_2_3.Y.n2 sky130_fd_sc_hd__inv_2_3.Y 4.0965
R2765 sky130_fd_sc_hd__inv_2_3.Y.n2 sky130_fd_sc_hd__inv_2_3.Y 4.01239
R2766 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_sc_hd__inv_2_3.Y.t0 3.02296
R2767 sky130_fd_sc_hd__inv_2_3.Y.n4 sky130_fd_sc_hd__inv_2_3.Y 2.0485
R2768 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_sc_hd__inv_2_3.Y.n4 1.55202
R2769 sky130_fd_sc_hd__inv_2_3.Y.t1 sky130_fd_sc_hd__inv_2_3.Y 0.227625
R2770 sky130_fd_sc_hd__inv_2_3.Y.t0 sky130_fd_sc_hd__inv_2_3.Y.t1 0.174201
R2771 sky130_fd_sc_hd__inv_2_3.Y.t0 sky130_fd_sc_hd__inv_2_3.Y 0.158396
R2772 sky130_fd_sc_hd__inv_2_0.Y.n1 sky130_fd_sc_hd__inv_2_0.Y.n0 111.322
R2773 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_sc_hd__inv_2_0.Y.n2 50.4671
R2774 sky130_fd_sc_hd__inv_2_0.Y.n0 sky130_fd_sc_hd__inv_2_0.Y.t3 26.5955
R2775 sky130_fd_sc_hd__inv_2_0.Y.n0 sky130_fd_sc_hd__inv_2_0.Y.t1 26.5955
R2776 sky130_fd_sc_hd__inv_2_0.Y.n2 sky130_fd_sc_hd__inv_2_0.Y.t4 24.9236
R2777 sky130_fd_sc_hd__inv_2_0.Y.n2 sky130_fd_sc_hd__inv_2_0.Y.t2 24.9236
R2778 sky130_fd_sc_hd__inv_2_0.Y.n4 sky130_fd_sc_hd__inv_2_0.Y 12.0325
R2779 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_sc_hd__inv_2_0.Y.n3 11.2645
R2780 sky130_fd_sc_hd__inv_2_0.Y.n5 sky130_fd_sc_hd__inv_2_0.Y 8.80626
R2781 sky130_fd_sc_hd__inv_2_0.Y.n3 sky130_fd_sc_hd__inv_2_0.Y 6.1445
R2782 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_sc_hd__inv_2_0.Y.n4 6.0197
R2783 sky130_fd_sc_hd__inv_2_0.Y.n4 sky130_fd_sc_hd__inv_2_0.Y 5.3765
R2784 sky130_fd_sc_hd__inv_2_0.Y.n3 sky130_fd_sc_hd__inv_2_0.Y 4.65505
R2785 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_sc_hd__inv_2_0.Y.n1 2.0485
R2786 sky130_fd_sc_hd__inv_2_0.Y.n1 sky130_fd_sc_hd__inv_2_0.Y 1.55202
R2787 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_sc_hd__inv_2_0.Y.t0 0.127353
R2788 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_sc_hd__inv_2_0.Y.n6 0.119257
R2789 sky130_fd_sc_hd__inv_2_0.Y.n5 sky130_fd_sc_hd__inv_2_0.Y 0.0465389
R2790 sky130_fd_sc_hd__inv_2_0.Y.t0 sky130_fd_sc_hd__inv_2_0.Y.n5 0.0388945
R2791 ctl2.n3 ctl2.t1 212.081
R2792 ctl2.n2 ctl2.t0 212.081
R2793 ctl2.n3 ctl2.t3 139.78
R2794 ctl2.n2 ctl2.t2 139.78
R2795 ctl2.n3 ctl2.n2 61.346
R2796 ctl2.n5 ctl2.n3 37.8794
R2797 ctl2.n5 ctl2.n0 9.30881
R2798 ctl2.n6 ctl2.n5 9.3005
R2799 ctl2.n7 ctl2.n6 9.01417
R2800 ctl2.n4 ctl2 3.48667
R2801 ctl2.n5 ctl2.n4 1.2812
R2802 ctl2.n7 ctl2.n0 0.0569565
R2803 ctl2.n6 ctl2.n1 0.03175
R2804 ctl2 ctl2.n7 0.00771154
R2805 ctl2.n4 ctl2.n1 0.00147336
R2806 ctl2.n1 ctl2.n0 0.00100057
R2807 sky130_fd_sc_hd__inv_2_5.Y.n4 sky130_fd_sc_hd__inv_2_5.Y.n3 111.32
R2808 sky130_fd_sc_hd__inv_2_5.Y sky130_fd_sc_hd__inv_2_5.Y.n0 50.4671
R2809 sky130_fd_sc_hd__inv_2_5.Y.n3 sky130_fd_sc_hd__inv_2_5.Y.t2 26.5955
R2810 sky130_fd_sc_hd__inv_2_5.Y.n3 sky130_fd_sc_hd__inv_2_5.Y.t1 26.5955
R2811 sky130_fd_sc_hd__inv_2_5.Y.n0 sky130_fd_sc_hd__inv_2_5.Y.t4 24.9236
R2812 sky130_fd_sc_hd__inv_2_5.Y.n0 sky130_fd_sc_hd__inv_2_5.Y.t3 24.9236
R2813 sky130_fd_sc_hd__inv_2_5.Y sky130_fd_sc_hd__inv_2_5.Y.n2 13.5685
R2814 sky130_fd_sc_hd__inv_2_5.Y sky130_fd_sc_hd__inv_2_5.Y.n1 11.2645
R2815 sky130_fd_sc_hd__inv_2_5.Y.n1 sky130_fd_sc_hd__inv_2_5.Y 6.1445
R2816 sky130_fd_sc_hd__inv_2_5.Y.n1 sky130_fd_sc_hd__inv_2_5.Y 4.65505
R2817 sky130_fd_sc_hd__inv_2_5.Y.n2 sky130_fd_sc_hd__inv_2_5.Y 3.8405
R2818 sky130_fd_sc_hd__inv_2_5.Y.n2 sky130_fd_sc_hd__inv_2_5.Y 3.68286
R2819 sky130_fd_sc_hd__inv_2_5.Y sky130_fd_sc_hd__inv_2_5.Y.t0 3.62224
R2820 sky130_fd_sc_hd__inv_2_5.Y.n4 sky130_fd_sc_hd__inv_2_5.Y 2.0485
R2821 sky130_fd_sc_hd__inv_2_5.Y sky130_fd_sc_hd__inv_2_5.Y.n4 1.55202
R2822 sky130_fd_sc_hd__inv_2_5.Y.t0 sky130_fd_sc_hd__inv_2_5.Y 0.0722572
R2823 ctl5.n3 ctl5.t2 212.081
R2824 ctl5.n2 ctl5.t0 212.081
R2825 ctl5.n3 ctl5.t3 139.78
R2826 ctl5.n2 ctl5.t1 139.78
R2827 ctl5.n3 ctl5.n2 61.346
R2828 ctl5.n5 ctl5.n3 38.5428
R2829 ctl5.n5 ctl5.n0 9.30881
R2830 ctl5.n6 ctl5.n5 9.3005
R2831 ctl5.n7 ctl5.n6 9.01417
R2832 ctl5.n4 ctl5 3.23067
R2833 ctl5.n5 ctl5.n4 1.2812
R2834 ctl5.n7 ctl5.n0 0.0569565
R2835 ctl5.n6 ctl5.n1 0.03175
R2836 ctl5 ctl5.n7 0.00771154
R2837 ctl5.n4 ctl5.n1 0.00147336
R2838 ctl5.n1 ctl5.n0 0.00100057
R2839 ctl1.n3 ctl1.t2 212.081
R2840 ctl1.n2 ctl1.t0 212.081
R2841 ctl1.n3 ctl1.t3 139.78
R2842 ctl1.n2 ctl1.t1 139.78
R2843 ctl1.n3 ctl1.n2 61.346
R2844 ctl1.n5 ctl1.n3 38.5428
R2845 ctl1.n5 ctl1.n0 9.30881
R2846 ctl1.n6 ctl1.n5 9.3005
R2847 ctl1.n7 ctl1.n6 9.01417
R2848 ctl1.n4 ctl1 3.09989
R2849 ctl1.n5 ctl1.n4 1.53719
R2850 ctl1.n7 ctl1.n0 0.0569565
R2851 ctl1.n6 ctl1.n1 0.03175
R2852 ctl1 ctl1.n7 0.00771154
R2853 ctl1.n4 ctl1.n1 0.00148276
R2854 ctl1.n1 ctl1.n0 0.00100057
R2855 dum.n3 dum.t2 212.081
R2856 dum.n2 dum.t0 212.081
R2857 dum.n3 dum.t3 139.78
R2858 dum.n2 dum.t1 139.78
R2859 dum.n3 dum.n2 61.346
R2860 dum.n5 dum.n3 38.5428
R2861 dum.n5 dum.n0 9.3127
R2862 dum.n6 dum.n5 9.3005
R2863 dum.n7 dum.n6 9.01808
R2864 dum.n4 dum 3.09989
R2865 dum.n5 dum.n4 1.53719
R2866 dum.n7 dum.n0 0.0569562
R2867 dum.n6 dum.n1 0.0278438
R2868 dum dum.n7 0.00771154
R2869 dum.n4 dum.n1 0.00148276
R2870 dum.n1 dum.n0 0.00100086
R2871 ctl0.n3 ctl0.t0 212.081
R2872 ctl0.n2 ctl0.t2 212.081
R2873 ctl0.n3 ctl0.t1 139.78
R2874 ctl0.n2 ctl0.t3 139.78
R2875 ctl0.n3 ctl0.n2 61.346
R2876 ctl0.n5 ctl0.n3 37.8794
R2877 ctl0.n5 ctl0.n0 9.3127
R2878 ctl0.n6 ctl0.n5 9.3005
R2879 ctl0.n7 ctl0.n6 9.01808
R2880 ctl0.n4 ctl0 3.61245
R2881 ctl0.n5 ctl0.n4 1.0252
R2882 ctl0.n7 ctl0.n0 0.0569562
R2883 ctl0.n6 ctl0.n1 0.0278438
R2884 ctl0 ctl0.n7 0.00771154
R2885 ctl0.n4 ctl0.n1 0.00146432
R2886 ctl0.n1 ctl0.n0 0.00100086
R2887 ctl3.n3 ctl3.t2 212.081
R2888 ctl3.n2 ctl3.t0 212.081
R2889 ctl3.n3 ctl3.t3 139.78
R2890 ctl3.n2 ctl3.t1 139.78
R2891 ctl3.n3 ctl3.n2 61.346
R2892 ctl3.n5 ctl3.n3 38.5428
R2893 ctl3.n5 ctl3.n0 9.30881
R2894 ctl3.n6 ctl3.n5 9.3005
R2895 ctl3.n7 ctl3.n6 9.01417
R2896 ctl3.n4 ctl3 3.09989
R2897 ctl3.n5 ctl3.n4 1.53719
R2898 ctl3.n7 ctl3.n0 0.0569565
R2899 ctl3.n6 ctl3.n1 0.03175
R2900 ctl3 ctl3.n7 0.00771154
R2901 ctl3.n4 ctl3.n1 0.00148276
R2902 ctl3.n1 ctl3.n0 0.00100057
R2903 ctl4.n3 ctl4.t1 212.081
R2904 ctl4.n2 ctl4.t0 212.081
R2905 ctl4.n3 ctl4.t3 139.78
R2906 ctl4.n2 ctl4.t2 139.78
R2907 ctl4.n3 ctl4.n2 61.346
R2908 ctl4.n5 ctl4.n3 38.5428
R2909 ctl4.n5 ctl4.n0 9.30881
R2910 ctl4.n6 ctl4.n5 9.3005
R2911 ctl4.n7 ctl4.n6 9.01417
R2912 ctl4.n4 ctl4 3.09989
R2913 ctl4.n5 ctl4.n4 1.53719
R2914 ctl4.n7 ctl4.n0 0.0569565
R2915 ctl4.n6 ctl4.n1 0.03175
R2916 ctl4 ctl4.n7 0.00771154
R2917 ctl4.n4 ctl4.n1 0.00148276
R2918 ctl4.n1 ctl4.n0 0.00100057
R2919 ctl6.n3 ctl6.t1 212.081
R2920 ctl6.n2 ctl6.t0 212.081
R2921 ctl6.n3 ctl6.t3 139.78
R2922 ctl6.n2 ctl6.t2 139.78
R2923 ctl6.n3 ctl6.n2 61.346
R2924 ctl6.n5 ctl6.n3 37.8794
R2925 ctl6.n5 ctl6.n0 9.31076
R2926 ctl6.n6 ctl6.n5 9.3005
R2927 ctl6.n7 ctl6.n6 9.01612
R2928 ctl6.n4 ctl6 3.48667
R2929 ctl6.n5 ctl6.n4 1.2812
R2930 ctl6.n7 ctl6.n0 0.0569564
R2931 ctl6.n6 ctl6.n1 0.0297969
R2932 ctl6 ctl6.n7 0.00771154
R2933 ctl6.n4 ctl6.n1 0.00147336
R2934 ctl6.n1 ctl6.n0 0.00100072
C0 carray_0.unitcap_324.cn sky130_fd_sc_hd__inv_2_7.VPB 8.98e-19
C1 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_sc_hd__inv_2_4.Y 3.2e-19
C2 sky130_fd_sc_hd__inv_2_2.Y carray_0.unitcap_119.cn 0.18f
C3 sky130_fd_sc_hd__inv_2_1.Y carray_0.unitcap_152.cn 0.18f
C4 sky130_fd_sc_hd__inv_2_8.Y ctl6 3.66e-19
C5 sky130_fd_sc_hd__inv_2_4.Y ctl1 0.159f
C6 carray_0.unitcap_8.cn carray_0.unitcap_9.cn 0.18f
C7 vin carray_0.unitcap_12.cn 0.00143f
C8 out carray_0.unitcap_160.cn 0.514f
C9 carray_0.unitcap_322.cn ctl2 0.00222f
C10 carray_0.unitcap_136.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C11 carray_0.unitcap_0.cn carray_0.unitcap_40.cn 0.0902f
C12 out carray_0.unitcap_119.cn 0.51f
C13 dum vdd 0.113f
C14 carray_0.unitcap_32.cn sample 0.00246f
C15 sky130_fd_sc_hd__inv_2_8.Y ctl1 5.89e-21
C16 carray_0.unitcap_216.cn carray_0.unitcap_240.cn 0.0902f
C17 carray_0.unitcap_11.cn sky130_fd_sc_hd__inv_2_2.Y 0.0902f
C18 out carray_0.unitcap_136.cn 0.514f
C19 carray_0.unitcap_331.cn sky130_fd_sc_hd__inv_2_0.Y 0.0445f
C20 carray_0.unitcap_247.cn sky130_fd_sc_hd__inv_2_0.Y 0.00213f
C21 carray_0.unitcap_135.cn sky130_fd_sc_hd__inv_2_1.Y 0.18f
C22 carray_0.unitcap_326.cn ctl7 2.83e-19
C23 vdd sky130_fd_sc_hd__inv_2_2.Y 3.06f
C24 carray_0.unitcap_8.cn out 0.503f
C25 sky130_fd_sc_hd__inv_2_7.Y sky130_fd_sc_hd__inv_2_5.Y 2.23e-21
C26 carray_0.unitcap_11.cn out 0.556f
C27 carray_0.unitcap_322.cn sky130_fd_sc_hd__inv_2_4.Y 0.155f
C28 vdd out 1.69f
C29 carray_0.unitcap_328.cn sky130_fd_sc_hd__inv_2_5.Y 0.131f
C30 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sw_top_1.sky130_fd_sc_hd__inv_4_1.Y 0.00289f
C31 sky130_fd_sc_hd__inv_2_1.Y carray_0.unitcap_192.cn 0.18f
C32 sky130_fd_sc_hd__inv_2_7.VPB carray_0.unitcap_320.cn 7.06e-19
C33 sky130_fd_sc_hd__inv_2_6.Y sky130_fd_sc_hd__inv_2_3.Y 0.0961f
C34 carray_0.unitcap_224.cn sky130_fd_sc_hd__inv_2_0.Y 0.18f
C35 carray_0.unitcap_334.cn sky130_fd_sc_hd__inv_2_7.VPB 0.00202f
C36 ctl2 sky130_fd_sc_hd__inv_2_7.VPB 0.0828f
C37 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_sc_hd__inv_2_7.VPB 0.00865f
C38 carray_0.unitcap_151.cn carray_0.unitcap_167.cn 0.0902f
C39 carray_0.unitcap_322.cn ctl1 0.00219f
C40 ctl5 sky130_fd_sc_hd__inv_2_0.Y 0.16f
C41 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_sc_hd__inv_2_0.Y 0.105f
C42 out carray_0.unitcap_168.cn 0.514f
C43 vdd ctl0 0.116f
C44 vin sw_top_2.sky130_fd_sc_hd__inv_4_1.Y 0.697f
C45 carray_0.unitcap_55.cn carray_0.unitcap_79.cn 0.0902f
C46 carray_0.unitcap_47.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C47 carray_0.unitcap_48.cn sample 0.00246f
C48 carray_0.unitcap_199.cn sky130_fd_sc_hd__inv_2_1.Y 0.18f
C49 carray_0.unitcap_338.cn sky130_fd_sc_hd__inv_2_0.Y 0.00213f
C50 ctl4 sky130_fd_sc_hd__inv_2_7.VPB 0.0827f
C51 carray_0.unitcap_10.cn sky130_fd_sc_hd__inv_2_2.Y 0.0902f
C52 out carray_0.unitcap_47.cn 0.51f
C53 carray_0.unitcap_247.cn carray_0.unitcap_239.cn 0.0902f
C54 carray_0.unitcap_10.cn out 0.557f
C55 sky130_fd_sc_hd__inv_2_4.Y sky130_fd_sc_hd__inv_2_7.VPB 0.00878f
C56 sky130_fd_sc_hd__inv_2_7.VPB ctl6 0.0828f
C57 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y sw_top_0.sky130_fd_sc_hd__inv_4_1.Y 0.585f
C58 out carray_0.unitcap_15.cn 0.501f
C59 carray_0.unitcap_256.cn carray_0.unitcap_9.cn 0.18f
C60 ctl5 carray_0.unitcap_326.cn 9.11e-19
C61 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_sc_hd__inv_2_7.VPB 0.00888f
C62 carray_0.unitcap_326.cn sky130_fd_sc_hd__inv_2_3.Y 0.0467f
C63 carray_0.unitcap_334.cn sky130_fd_sc_hd__inv_2_5.Y 0.348f
C64 ctl1 sky130_fd_sc_hd__inv_2_7.VPB 0.0826f
C65 ctl2 sky130_fd_sc_hd__inv_2_5.Y 0.16f
C66 sky130_fd_sc_hd__inv_2_2.Y carray_0.unitcap_88.cn 0.18f
C67 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_sc_hd__inv_2_5.Y 0.357f
C68 carray_0.unitcap_56.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C69 carray_0.unitcap_80.cn carray_0.unitcap_64.cn 0.0902f
C70 vin sw_top_0.sky130_fd_sc_hd__inv_4_0.Y 0.368f
C71 carray_0.unitcap_256.cn sky130_fd_sc_hd__inv_2_2.Y 0.0902f
C72 carray_0.unitcap_167.cn carray_0.unitcap_183.cn 0.0902f
C73 sky130_fd_sc_hd__inv_2_3.Y carray_0.unitcap_255.cn 0.18f
C74 vin sw_top_2.sky130_fd_sc_hd__inv_4_0.Y 0.368f
C75 out carray_0.unitcap_128.cn 0.514f
C76 sky130_fd_sc_hd__inv_2_7.Y carray_0.unitcap_321.cn 0.18f
C77 out carray_0.unitcap_88.cn 0.514f
C78 carray_0.unitcap_14.cn carray_0.unitcap_12.cn 0.18f
C79 vdd sky130_fd_sc_hd__inv_2_6.Y 0.219f
C80 carray_0.unitcap_79.cn carray_0.unitcap_87.cn 0.0902f
C81 carray_0.unitcap_56.cn out 0.514f
C82 carray_0.unitcap_256.cn out 0.557f
C83 carray_0.unitcap_255.cn carray_0.unitcap_338.cn 0.0902f
C84 vdd sw_top_1.sky130_fd_sc_hd__inv_4_1.Y 1.98f
C85 ctl4 sky130_fd_sc_hd__inv_2_5.Y 3.33e-19
C86 vin sw_top_3.sky130_fd_sc_hd__inv_4_1.Y 0.705f
C87 carray_0.unitcap_103.cn carray_0.unitcap_127.cn 0.0902f
C88 carray_0.unitcap_11.cn carray_0.unitcap_13.cn 0.18f
C89 carray_0.unitcap_31.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C90 carray_0.unitcap_143.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C91 carray_0.unitcap_330.cn sky130_fd_sc_hd__inv_2_1.Y 0.145f
C92 vdd sky130_fd_sc_hd__inv_2_0.Y 0.22f
C93 carray_0.unitcap_224.cn carray_0.unitcap_216.cn 0.0902f
C94 vin carray_0.unitcap_288.cn 0.00185f
C95 vdd carray_0.unitcap_13.cn 4.57e-20
C96 carray_0.unitcap_328.cn ctl3 0.00161f
C97 out carray_0.unitcap_31.cn 0.51f
C98 sky130_fd_sc_hd__inv_2_4.Y sky130_fd_sc_hd__inv_2_5.Y 0.59f
C99 out carray_0.unitcap_143.cn 0.51f
C100 sky130_fd_sc_hd__inv_2_8.Y carray_0.unitcap_240.cn 0.18f
C101 sky130_fd_sc_hd__inv_2_5.Y ctl6 2.94e-20
C102 carray_0.unitcap_322.cn sky130_fd_sc_hd__inv_2_7.VPB 6.68e-19
C103 sample carray_0.unitcap_72.cn 0.00246f
C104 carray_0.unitcap_334.cn ctl7 1.73e-19
C105 sky130_fd_sc_hd__inv_2_7.Y sky130_fd_sc_hd__inv_2_3.Y 0.0925f
C106 carray_0.unitcap_120.cn carray_0.unitcap_112.cn 0.0902f
C107 sky130_fd_sc_hd__inv_2_1.Y ctl7 0.0541f
C108 carray_0.unitcap_191.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C109 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_sc_hd__inv_2_5.Y 0.248f
C110 ctl5 carray_0.unitcap_328.cn 7.05e-21
C111 carray_0.unitcap_328.cn sky130_fd_sc_hd__inv_2_3.Y 0.0124f
C112 ctl1 sky130_fd_sc_hd__inv_2_5.Y 0.00126f
C113 sky130_fd_sc_hd__inv_2_2.Y carray_0.unitcap_96.cn 0.18f
C114 carray_0.unitcap_24.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C115 out carray_0.unitcap_191.cn 0.51f
C116 ctl4 ctl7 1.76e-19
C117 carray_0.unitcap_9.cn sky130_fd_sc_hd__inv_2_2.Y 0.0902f
C118 carray_0.unitcap_48.cn carray_0.unitcap_72.cn 0.0902f
C119 out carray_0.unitcap_144.cn 0.514f
C120 carray_0.unitcap_175.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C121 out carray_0.unitcap_96.cn 0.514f
C122 vdd carray_0.unitcap_326.cn 0.00104f
C123 carray_0.unitcap_24.cn out 0.514f
C124 dum out 9.4e-19
C125 carray_0.unitcap_9.cn out 0.557f
C126 carray_0.unitcap_338.cn carray_0.unitcap_336.cn 0.0902f
C127 sky130_fd_sc_hd__inv_2_4.Y ctl7 5.61e-22
C128 carray_0.unitcap_334.cn carray_0.unitcap_331.cn 0.18f
C129 carray_0.unitcap_127.cn carray_0.unitcap_119.cn 0.0902f
C130 ctl7 ctl6 0.0959f
C131 carray_0.unitcap_321.cn carray_0.unitcap_320.cn 0.0902f
C132 out carray_0.unitcap_175.cn 0.51f
C133 carray_0.unitcap_159.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C134 vdd sw_top_0.sky130_fd_sc_hd__inv_4_1.Y 1.98f
C135 carray_0.unitcap_331.cn sky130_fd_sc_hd__inv_2_1.Y 0.0069f
C136 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y sw_top_1.sky130_fd_sc_hd__inv_4_0.Y 0.00267f
C137 dum ctl0 0.0951f
C138 sky130_fd_sc_hd__inv_2_8.Y ctl7 3.69e-19
C139 carray_0.unitcap_337.cn sky130_fd_sc_hd__inv_2_2.Y 0.138f
C140 out sky130_fd_sc_hd__inv_2_2.Y 84.2f
C141 out carray_0.unitcap_159.cn 0.51f
C142 carray_0.unitcap_11.cn vin 0.0484f
C143 carray_0.unitcap_322.cn sky130_fd_sc_hd__inv_2_5.Y 0.00397f
C144 carray_0.unitcap_191.cn carray_0.unitcap_207.cn 0.0902f
C145 ctl3 ctl2 0.0964f
C146 carray_0.unitcap_167.cn sky130_fd_sc_hd__inv_2_1.Y 0.18f
C147 carray_0.unitcap_223.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C148 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y sw_top_3.sky130_fd_sc_hd__inv_4_0.Y 0.00267f
C149 carray_0.unitcap_112.cn carray_0.unitcap_136.cn 0.0902f
C150 out carray_0.unitcap_337.cn 0.505f
C151 vdd vin 3.04f
C152 carray_0.unitcap_231.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C153 carray_0.unitcap_63.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C154 sample carray_0.unitcap_0.cn 0.00246f
C155 sample sw_top_2.sky130_fd_sc_hd__inv_4_1.Y 0.561f
C156 out carray_0.unitcap_223.cn 0.51f
C157 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sw_top_3.sky130_fd_sc_hd__inv_4_0.Y 0.585f
C158 out carray_0.unitcap_200.cn 0.514f
C159 vdd sky130_fd_sc_hd__inv_2_7.Y 0.219f
C160 ctl4 ctl3 0.0964f
C161 out carray_0.unitcap_231.cn 0.51f
C162 carray_0.unitcap_334.cn sky130_fd_sc_hd__inv_2_3.Y 0.0355f
C163 ctl2 sky130_fd_sc_hd__inv_2_3.Y 0.00122f
C164 ctl5 sky130_fd_sc_hd__inv_2_1.Y 0.00139f
C165 out carray_0.unitcap_63.cn 0.51f
C166 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_sc_hd__inv_2_1.Y 0.325f
C167 out ctl0 9.46e-19
C168 carray_0.unitcap_160.cn carray_0.unitcap_176.cn 0.0902f
C169 carray_0.unitcap_231.cn carray_0.unitcap_223.cn 0.0902f
C170 carray_0.unitcap_207.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C171 vdd carray_0.unitcap_328.cn 9.92e-19
C172 carray_0.unitcap_331.cn sky130_fd_sc_hd__inv_2_8.Y 0.0404f
C173 sky130_fd_sc_hd__inv_2_8.Y carray_0.unitcap_247.cn 0.18f
C174 carray_0.unitcap_324.cn vdd 8.02e-19
C175 sky130_fd_sc_hd__inv_2_4.Y ctl3 4.22e-19
C176 out carray_0.unitcap_208.cn 0.514f
C177 ctl5 ctl4 0.0958f
C178 ctl4 sky130_fd_sc_hd__inv_2_3.Y 0.0504f
C179 out carray_0.unitcap_207.cn 0.51f
C180 carray_0.unitcap_32.cn sw_top_3.sky130_fd_sc_hd__inv_4_1.Y 2.32e-19
C181 sky130_fd_sc_hd__inv_2_5.Y sky130_fd_sc_hd__inv_2_7.VPB 0.00795f
C182 sky130_fd_sc_hd__inv_2_8.Y ctl3 0.00135f
C183 carray_0.unitcap_10.cn vin 0.0542f
C184 carray_0.unitcap_191.cn sky130_fd_sc_hd__inv_2_0.Y 0.18f
C185 dum sky130_fd_sc_hd__inv_2_6.Y 0.00123f
C186 ctl5 sky130_fd_sc_hd__inv_2_4.Y 2.14e-21
C187 sky130_fd_sc_hd__inv_2_4.Y sky130_fd_sc_hd__inv_2_3.Y 0.251f
C188 ctl5 ctl6 0.0958f
C189 sky130_fd_sc_hd__inv_2_3.Y ctl6 2.94e-19
C190 sky130_fd_sc_hd__inv_2_1.Y carray_0.unitcap_160.cn 0.18f
C191 sample sw_top_0.sky130_fd_sc_hd__inv_4_0.Y 0.0117f
C192 carray_0.unitcap_95.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C193 sample sw_top_2.sky130_fd_sc_hd__inv_4_0.Y 0.037f
C194 out carray_0.unitcap_232.cn 0.514f
C195 sky130_fd_sc_hd__inv_2_8.Y ctl5 0.0518f
C196 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_sc_hd__inv_2_3.Y 1.73f
C197 out carray_0.unitcap_95.cn 0.51f
C198 sample sw_top_3.sky130_fd_sc_hd__inv_4_1.Y 0.561f
C199 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_2_2.Y 1.04f
C200 carray_0.unitcap_8.cn carray_0.unitcap_16.cn 0.0902f
C201 carray_0.unitcap_176.cn carray_0.unitcap_168.cn 0.0902f
C202 vdd sw_top_1.sky130_fd_sc_hd__inv_4_0.Y 0.849f
C203 sky130_fd_sc_hd__inv_2_7.VPB ctl7 0.0932f
C204 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_sc_hd__inv_2_2.Y 0.554f
C205 sample carray_0.unitcap_288.cn 0.0193f
C206 out sky130_fd_sc_hd__inv_2_6.Y 0.536f
C207 vdd carray_0.unitcap_320.cn 7.24e-20
C208 carray_0.unitcap_16.cn vdd 0.0016f
C209 carray_0.unitcap_13.cn sky130_fd_sc_hd__inv_2_2.Y 0.0902f
C210 out sw_top_1.sky130_fd_sc_hd__inv_4_1.Y 0.696f
C211 carray_0.unitcap_334.cn vdd 4.49e-19
C212 vdd ctl2 0.116f
C213 vdd sky130_fd_sc_hd__inv_2_1.Y 0.22f
C214 out sky130_fd_sc_hd__inv_2_0.Y 17.5f
C215 vdd sw_top_3.sky130_fd_sc_hd__inv_4_0.Y 0.849f
C216 carray_0.unitcap_337.cn sky130_fd_sc_hd__inv_2_0.Y 0.00682f
C217 out carray_0.unitcap_13.cn 0.558f
C218 sky130_fd_sc_hd__inv_2_6.Y ctl0 0.16f
C219 carray_0.unitcap_223.cn sky130_fd_sc_hd__inv_2_0.Y 0.181f
C220 carray_0.unitcap_23.cn carray_0.unitcap_15.cn 0.0902f
C221 carray_0.unitcap_151.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C222 carray_0.unitcap_159.cn carray_0.unitcap_151.cn 0.0902f
C223 carray_0.unitcap_40.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C224 carray_0.unitcap_231.cn sky130_fd_sc_hd__inv_2_0.Y 0.18f
C225 carray_0.unitcap_322.cn sky130_fd_sc_hd__inv_2_3.Y 0.00223f
C226 vdd ctl4 0.116f
C227 sky130_fd_sc_hd__inv_2_1.Y carray_0.unitcap_168.cn 0.18f
C228 out carray_0.unitcap_151.cn 0.51f
C229 carray_0.unitcap_330.cn sky130_fd_sc_hd__inv_2_5.Y 0.0919f
C230 carray_0.unitcap_40.cn out 0.514f
C231 carray_0.unitcap_32.cn vdd 4.58e-19
C232 carray_0.unitcap_71.cn carray_0.unitcap_87.cn 0.0902f
C233 vdd sky130_fd_sc_hd__inv_2_4.Y 0.219f
C234 carray_0.unitcap_208.cn sky130_fd_sc_hd__inv_2_0.Y 0.18f
C235 vdd ctl6 0.116f
C236 carray_0.unitcap_80.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C237 ctl3 sky130_fd_sc_hd__inv_2_7.VPB 0.0829f
C238 carray_0.unitcap_79.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C239 sky130_fd_sc_hd__inv_2_5.Y ctl7 1.47e-20
C240 carray_0.unitcap_255.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C241 out carray_0.unitcap_326.cn 0.501f
C242 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_2_2.Y 1.27f
C243 vdd sky130_fd_sc_hd__inv_2_8.Y 0.219f
C244 out carray_0.unitcap_80.cn 0.514f
C245 vdd ctl1 0.116f
C246 carray_0.unitcap_8.cn sample 0.00246f
C247 carray_0.unitcap_11.cn sample 4.94e-19
C248 carray_0.unitcap_239.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C249 out carray_0.unitcap_79.cn 0.51f
C250 carray_0.unitcap_183.cn carray_0.unitcap_175.cn 0.0902f
C251 out carray_0.unitcap_255.cn 0.51f
C252 carray_0.unitcap_23.cn carray_0.unitcap_31.cn 0.0902f
C253 out sw_top_0.sky130_fd_sc_hd__inv_4_1.Y 0.678f
C254 dum sky130_fd_sc_hd__inv_2_7.Y 0.162f
C255 sample vdd 1.46f
C256 ctl5 sky130_fd_sc_hd__inv_2_7.VPB 0.0826f
C257 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_sc_hd__inv_2_7.VPB 0.00809f
C258 out carray_0.unitcap_239.cn 0.51f
C259 vin sky130_fd_sc_hd__inv_2_2.Y 1.86f
C260 carray_0.unitcap_183.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C261 sky130_fd_sc_hd__inv_2_1.Y carray_0.unitcap_128.cn 0.18f
C262 sky130_fd_sc_hd__inv_2_2.Y carray_0.unitcap_127.cn 0.18f
C263 carray_0.unitcap_324.cn dum 0.00223f
C264 out vin 9.61f
C265 out carray_0.unitcap_183.cn 0.51f
C266 carray_0.unitcap_15.cn carray_0.unitcap_14.cn 0.18f
C267 carray_0.unitcap_331.cn sky130_fd_sc_hd__inv_2_5.Y 0.135f
C268 carray_0.unitcap_112.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C269 out carray_0.unitcap_127.cn 0.51f
C270 out carray_0.unitcap_216.cn 0.514f
C271 carray_0.unitcap_322.cn vdd 0.00109f
C272 out sky130_fd_sc_hd__inv_2_7.Y 0.542f
C273 out carray_0.unitcap_112.cn 0.514f
C274 ctl3 sky130_fd_sc_hd__inv_2_5.Y 0.0494f
C275 carray_0.unitcap_336.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C276 out carray_0.unitcap_328.cn 0.501f
C277 carray_0.unitcap_330.cn carray_0.unitcap_331.cn 0.18f
C278 carray_0.unitcap_324.cn out 0.505f
C279 ctl0 sky130_fd_sc_hd__inv_2_7.Y 0.0456f
C280 carray_0.unitcap_10.cn sample 0.00331f
C281 carray_0.unitcap_32.cn carray_0.unitcap_56.cn 0.0902f
C282 out carray_0.unitcap_336.cn 0.496f
C283 carray_0.unitcap_337.cn carray_0.unitcap_336.cn 0.18f
C284 carray_0.unitcap_23.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C285 ctl5 sky130_fd_sc_hd__inv_2_5.Y 7e-19
C286 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_sc_hd__inv_2_5.Y 1.03f
C287 carray_0.unitcap_324.cn ctl0 0.00232f
C288 out carray_0.unitcap_23.cn 0.512f
C289 carray_0.unitcap_16.cn carray_0.unitcap_24.cn 0.0902f
C290 sky130_fd_sc_hd__inv_2_1.Y carray_0.unitcap_144.cn 0.18f
C291 carray_0.unitcap_321.cn carray_0.unitcap_248.cn 0.0902f
C292 carray_0.unitcap_338.cn sky130_fd_sc_hd__inv_2_5.Y 0.18f
C293 out carray_0.unitcap_176.cn 0.514f
C294 carray_0.unitcap_326.cn sky130_fd_sc_hd__inv_2_0.Y 0.00206f
C295 vdd sky130_fd_sc_hd__inv_2_7.VPB 0.801f
C296 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y sky130_fd_sc_hd__inv_2_2.Y 0.424f
C297 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y sw_top_2.sky130_fd_sc_hd__inv_4_0.Y 0.585f
C298 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y sw_top_0.sky130_fd_sc_hd__inv_4_1.Y 0.00289f
C299 carray_0.unitcap_7.cn carray_0.unitcap_47.cn 0.0902f
C300 carray_0.unitcap_56.cn sample 0.0026f
C301 carray_0.unitcap_192.cn carray_0.unitcap_168.cn 0.0902f
C302 carray_0.unitcap_175.cn sky130_fd_sc_hd__inv_2_1.Y 0.18f
C303 carray_0.unitcap_256.cn sample 0.207f
C304 carray_0.unitcap_255.cn sky130_fd_sc_hd__inv_2_0.Y 0.00213f
C305 carray_0.unitcap_16.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C306 carray_0.unitcap_111.cn carray_0.unitcap_103.cn 0.0902f
C307 carray_0.unitcap_334.cn sky130_fd_sc_hd__inv_2_2.Y 0.00122f
C308 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y sw_top_3.sky130_fd_sc_hd__inv_4_1.Y 0.00289f
C309 carray_0.unitcap_128.cn carray_0.unitcap_152.cn 0.0902f
C310 out sw_top_1.sky130_fd_sc_hd__inv_4_0.Y 0.302f
C311 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_sc_hd__inv_2_2.Y 4.15f
C312 carray_0.unitcap_239.cn sky130_fd_sc_hd__inv_2_0.Y 0.00213f
C313 carray_0.unitcap_88.cn carray_0.unitcap_104.cn 0.0902f
C314 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y sky130_fd_sc_hd__inv_2_2.Y 0.461f
C315 ctl5 ctl7 1.96e-19
C316 carray_0.unitcap_159.cn sky130_fd_sc_hd__inv_2_1.Y 0.18f
C317 sky130_fd_sc_hd__inv_2_3.Y ctl7 9.34e-19
C318 out carray_0.unitcap_320.cn 0.496f
C319 sky130_fd_sc_hd__inv_2_3.Y carray_0.unitcap_248.cn 0.18f
C320 carray_0.unitcap_16.cn out 0.515f
C321 vin sw_top_1.sky130_fd_sc_hd__inv_4_1.Y 0.705f
C322 carray_0.unitcap_288.cn sw_top_2.sky130_fd_sc_hd__inv_4_1.Y 0.00736f
C323 carray_0.unitcap_334.cn out 0.501f
C324 out ctl2 9.44e-19
C325 vdd carray_0.unitcap_72.cn 0.00146f
C326 out sky130_fd_sc_hd__inv_2_1.Y 35.4f
C327 carray_0.unitcap_337.cn sky130_fd_sc_hd__inv_2_1.Y 0.13f
C328 carray_0.unitcap_56.cn carray_0.unitcap_48.cn 0.0902f
C329 dum sky130_fd_sc_hd__inv_2_4.Y 1.2e-20
C330 sky130_fd_sc_hd__inv_2_6.Y sky130_fd_sc_hd__inv_2_7.Y 0.503f
C331 out sw_top_3.sky130_fd_sc_hd__inv_4_0.Y 0.322f
C332 carray_0.unitcap_47.cn carray_0.unitcap_39.cn 0.0902f
C333 vin carray_0.unitcap_13.cn 0.00557f
C334 sky130_fd_sc_hd__inv_2_1.Y carray_0.unitcap_200.cn 0.18f
C335 carray_0.unitcap_216.cn sky130_fd_sc_hd__inv_2_0.Y 0.18f
C336 carray_0.unitcap_14.cn sky130_fd_sc_hd__inv_2_2.Y 0.0902f
C337 carray_0.unitcap_324.cn sky130_fd_sc_hd__inv_2_6.Y 0.15f
C338 out ctl4 0.00107f
C339 carray_0.unitcap_32.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C340 dum ctl1 5.3e-20
C341 sky130_fd_sc_hd__inv_2_4.Y sky130_fd_sc_hd__inv_2_2.Y 1.29e-23
C342 sky130_fd_sc_hd__inv_2_2.Y ctl6 0.00123f
C343 vdd sky130_fd_sc_hd__inv_2_5.Y 0.219f
C344 out carray_0.unitcap_14.cn 0.556f
C345 carray_0.unitcap_80.cn sw_top_0.sky130_fd_sc_hd__inv_4_1.Y 5.45e-19
C346 sample carray_0.unitcap_24.cn 0.00277f
C347 carray_0.unitcap_32.cn out 0.514f
C348 out sky130_fd_sc_hd__inv_2_4.Y 1.03f
C349 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_sc_hd__inv_2_2.Y 0.291f
C350 out ctl6 0.00107f
C351 carray_0.unitcap_9.cn sample 0.00958f
C352 carray_0.unitcap_207.cn sky130_fd_sc_hd__inv_2_1.Y 0.18f
C353 carray_0.unitcap_31.cn carray_0.unitcap_7.cn 0.0902f
C354 carray_0.unitcap_336.cn sky130_fd_sc_hd__inv_2_0.Y 0.00213f
C355 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sw_top_2.sky130_fd_sc_hd__inv_4_0.Y 4.9e-19
C356 carray_0.unitcap_143.cn carray_0.unitcap_135.cn 0.0902f
C357 carray_0.unitcap_152.cn carray_0.unitcap_144.cn 0.0902f
C358 carray_0.unitcap_255.cn carray_0.unitcap_239.cn 0.0902f
C359 ctl3 sky130_fd_sc_hd__inv_2_3.Y 0.161f
C360 out sky130_fd_sc_hd__inv_2_8.Y 8.84f
C361 carray_0.unitcap_104.cn carray_0.unitcap_96.cn 0.0902f
C362 carray_0.unitcap_64.cn sw_top_0.sky130_fd_sc_hd__inv_4_0.Y 1e-20
C363 out ctl1 8.28e-19
C364 sample sky130_fd_sc_hd__inv_2_2.Y 2.52f
C365 sky130_fd_sc_hd__inv_2_4.Y ctl0 0.00131f
C366 vin sw_top_0.sky130_fd_sc_hd__inv_4_1.Y 0.417f
C367 carray_0.unitcap_11.cn sw_top_2.sky130_fd_sc_hd__inv_4_1.Y 0.00862f
C368 sample out 0.122f
C369 vdd ctl7 0.117f
C370 vdd carray_0.unitcap_0.cn 0.00118f
C371 ctl5 sky130_fd_sc_hd__inv_2_3.Y 2.94e-19
C372 vdd sw_top_2.sky130_fd_sc_hd__inv_4_1.Y 1.99f
C373 carray_0.unitcap_326.cn carray_0.unitcap_328.cn 0.18f
C374 ctl1 ctl0 0.0967f
C375 sky130_fd_sc_hd__inv_2_2.Y carray_0.unitcap_104.cn 0.18f
C376 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y sw_top_1.sky130_fd_sc_hd__inv_4_1.Y 0.585f
C377 carray_0.unitcap_48.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C378 out carray_0.unitcap_152.cn 0.514f
C379 carray_0.unitcap_71.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C380 out carray_0.unitcap_104.cn 0.514f
C381 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y sw_top_1.sky130_fd_sc_hd__inv_4_1.Y 4.9e-19
C382 carray_0.unitcap_191.cn carray_0.unitcap_215.cn 0.0902f
C383 carray_0.unitcap_48.cn out 0.514f
C384 carray_0.unitcap_334.cn sky130_fd_sc_hd__inv_2_0.Y 0.00144f
C385 carray_0.unitcap_322.cn out 0.502f
C386 sky130_fd_sc_hd__inv_2_1.Y sky130_fd_sc_hd__inv_2_0.Y 3.17f
C387 carray_0.unitcap_7.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C388 out carray_0.unitcap_71.cn 0.51f
C389 carray_0.unitcap_135.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C390 carray_0.unitcap_135.cn carray_0.unitcap_159.cn 0.0902f
C391 out carray_0.unitcap_7.cn 0.51f
C392 dum sky130_fd_sc_hd__inv_2_7.VPB 0.0962f
C393 sky130_fd_sc_hd__inv_2_8.Y carray_0.unitcap_232.cn 0.18f
C394 out carray_0.unitcap_135.cn 0.51f
C395 ctl4 sky130_fd_sc_hd__inv_2_0.Y 0.00127f
C396 carray_0.unitcap_151.cn sky130_fd_sc_hd__inv_2_1.Y 0.18f
C397 sky130_fd_sc_hd__inv_2_4.Y sky130_fd_sc_hd__inv_2_6.Y 0.504f
C398 carray_0.unitcap_10.cn sw_top_2.sky130_fd_sc_hd__inv_4_1.Y 0.0123f
C399 vdd sw_top_0.sky130_fd_sc_hd__inv_4_0.Y 0.848f
C400 carray_0.unitcap_324.cn sky130_fd_sc_hd__inv_2_7.Y 0.307f
C401 carray_0.unitcap_215.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C402 vdd sw_top_2.sky130_fd_sc_hd__inv_4_0.Y 0.844f
C403 vdd ctl3 0.116f
C404 carray_0.unitcap_39.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C405 sky130_fd_sc_hd__inv_2_4.Y sky130_fd_sc_hd__inv_2_0.Y 1.23e-21
C406 sky130_fd_sc_hd__inv_2_0.Y ctl6 0.0517f
C407 sky130_fd_sc_hd__inv_2_2.Y sky130_fd_sc_hd__inv_2_7.VPB 0.0164f
C408 out carray_0.unitcap_192.cn 0.514f
C409 carray_0.unitcap_175.cn carray_0.unitcap_199.cn 0.0902f
C410 out carray_0.unitcap_215.cn 0.51f
C411 sky130_fd_sc_hd__inv_2_6.Y ctl1 0.047f
C412 carray_0.unitcap_334.cn carray_0.unitcap_326.cn 0.18f
C413 vdd sw_top_3.sky130_fd_sc_hd__inv_4_1.Y 1.98f
C414 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y sw_top_0.sky130_fd_sc_hd__inv_4_1.Y 4.9e-19
C415 out carray_0.unitcap_39.cn 0.51f
C416 carray_0.unitcap_326.cn sky130_fd_sc_hd__inv_2_1.Y 0.00168f
C417 carray_0.unitcap_192.cn carray_0.unitcap_200.cn 0.0902f
C418 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_sc_hd__inv_2_0.Y 2.06f
C419 out sky130_fd_sc_hd__inv_2_7.VPB 0.00464f
C420 carray_0.unitcap_199.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C421 vdd ctl5 0.116f
C422 vdd sky130_fd_sc_hd__inv_2_3.Y 0.219f
C423 vdd carray_0.unitcap_288.cn 0.107f
C424 carray_0.unitcap_215.cn carray_0.unitcap_231.cn 0.0902f
C425 vdd carray_0.unitcap_64.cn 4.58e-19
C426 sample sw_top_1.sky130_fd_sc_hd__inv_4_1.Y 0.561f
C427 carray_0.unitcap_32.cn carray_0.unitcap_40.cn 0.0902f
C428 carray_0.unitcap_39.cn carray_0.unitcap_63.cn 0.0902f
C429 out carray_0.unitcap_199.cn 0.51f
C430 carray_0.unitcap_72.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C431 vin sw_top_1.sky130_fd_sc_hd__inv_4_0.Y 0.368f
C432 ctl0 sky130_fd_sc_hd__inv_2_7.VPB 0.0827f
C433 dum sky130_fd_sc_hd__inv_2_5.Y 6.19e-21
C434 carray_0.unitcap_71.cn carray_0.unitcap_95.cn 0.0902f
C435 carray_0.unitcap_12.cn sky130_fd_sc_hd__inv_2_2.Y 0.0902f
C436 out carray_0.unitcap_72.cn 0.514f
C437 carray_0.unitcap_10.cn sw_top_2.sky130_fd_sc_hd__inv_4_0.Y 0.00207f
C438 sky130_fd_sc_hd__inv_2_4.Y carray_0.unitcap_326.cn 0.091f
C439 carray_0.unitcap_183.cn sky130_fd_sc_hd__inv_2_1.Y 0.18f
C440 carray_0.unitcap_326.cn ctl6 0.00219f
C441 carray_0.unitcap_322.cn sky130_fd_sc_hd__inv_2_6.Y 0.275f
C442 vin sw_top_3.sky130_fd_sc_hd__inv_4_0.Y 0.368f
C443 carray_0.unitcap_48.cn sw_top_1.sky130_fd_sc_hd__inv_4_1.Y 8.31e-19
C444 sky130_fd_sc_hd__inv_2_7.Y carray_0.unitcap_320.cn 0.109f
C445 out carray_0.unitcap_12.cn 0.556f
C446 sample carray_0.unitcap_40.cn 0.00329f
C447 out carray_0.unitcap_240.cn 0.514f
C448 sky130_fd_sc_hd__inv_2_5.Y sky130_fd_sc_hd__inv_2_2.Y 0.134f
C449 sky130_fd_sc_hd__inv_2_8.Y carray_0.unitcap_326.cn 0.00261f
C450 out carray_0.unitcap_184.cn 0.514f
C451 carray_0.unitcap_199.cn carray_0.unitcap_207.cn 0.0902f
C452 carray_0.unitcap_324.cn carray_0.unitcap_320.cn 0.18f
C453 carray_0.unitcap_10.cn carray_0.unitcap_288.cn 0.18f
C454 out sky130_fd_sc_hd__inv_2_5.Y 2.02f
C455 carray_0.unitcap_337.cn sky130_fd_sc_hd__inv_2_5.Y 0.0902f
C456 carray_0.unitcap_200.cn carray_0.unitcap_184.cn 0.0902f
C457 sample carray_0.unitcap_80.cn 7.14e-19
C458 carray_0.unitcap_24.cn carray_0.unitcap_0.cn 0.0902f
C459 sky130_fd_sc_hd__inv_2_8.Y carray_0.unitcap_239.cn 0.18f
C460 carray_0.unitcap_330.cn sky130_fd_sc_hd__inv_2_2.Y 0.00122f
C461 carray_0.unitcap_11.cn vdd 0.0039f
C462 carray_0.unitcap_24.cn sw_top_2.sky130_fd_sc_hd__inv_4_1.Y 6.3e-19
C463 ctl4 carray_0.unitcap_328.cn 0.00222f
C464 sample sw_top_0.sky130_fd_sc_hd__inv_4_1.Y 0.485f
C465 ctl0 sky130_fd_sc_hd__inv_2_5.Y 1.27e-20
C466 sky130_fd_sc_hd__inv_2_4.Y sky130_fd_sc_hd__inv_2_7.Y 0.00132f
C467 out carray_0.unitcap_330.cn 0.502f
C468 carray_0.unitcap_330.cn carray_0.unitcap_337.cn 0.18f
C469 carray_0.unitcap_208.cn carray_0.unitcap_184.cn 0.0902f
C470 sky130_fd_sc_hd__inv_2_6.Y sky130_fd_sc_hd__inv_2_7.VPB 0.00782f
C471 sky130_fd_sc_hd__inv_2_2.Y ctl7 0.16f
C472 carray_0.unitcap_64.cn carray_0.unitcap_88.cn 0.0902f
C473 carray_0.unitcap_0.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C474 carray_0.unitcap_215.cn sky130_fd_sc_hd__inv_2_0.Y 0.18f
C475 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_2_2.Y 1.16f
C476 sky130_fd_sc_hd__inv_2_4.Y carray_0.unitcap_328.cn 0.317f
C477 carray_0.unitcap_256.cn carray_0.unitcap_288.cn 0.18f
C478 sky130_fd_sc_hd__inv_2_1.Y carray_0.unitcap_176.cn 0.18f
C479 carray_0.unitcap_111.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C480 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_sc_hd__inv_2_7.VPB 0.00896f
C481 ctl1 sky130_fd_sc_hd__inv_2_7.Y 3.56e-20
C482 sample vin 0.00448f
C483 out ctl7 6.9e-19
C484 carray_0.unitcap_0.cn out 0.514f
C485 out carray_0.unitcap_248.cn 0.514f
C486 out sw_top_2.sky130_fd_sc_hd__inv_4_1.Y 0.516f
C487 sky130_fd_sc_hd__inv_2_8.Y carray_0.unitcap_328.cn 0.00246f
C488 carray_0.unitcap_240.cn carray_0.unitcap_232.cn 0.0902f
C489 out carray_0.unitcap_111.cn 0.51f
C490 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y sw_top_1.sky130_fd_sc_hd__inv_4_0.Y 0.00267f
C491 carray_0.unitcap_55.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C492 carray_0.unitcap_11.cn carray_0.unitcap_10.cn 0.18f
C493 carray_0.unitcap_334.cn sky130_fd_sc_hd__inv_2_1.Y 0.00242f
C494 carray_0.unitcap_331.cn sky130_fd_sc_hd__inv_2_2.Y 0.00122f
C495 carray_0.unitcap_247.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C496 carray_0.unitcap_10.cn vdd 0.0185f
C497 out carray_0.unitcap_55.cn 0.51f
C498 carray_0.unitcap_136.cn carray_0.unitcap_128.cn 0.0902f
C499 carray_0.unitcap_120.cn carray_0.unitcap_96.cn 0.0902f
C500 out carray_0.unitcap_331.cn 0.501f
C501 carray_0.unitcap_13.cn carray_0.unitcap_12.cn 0.18f
C502 ctl4 ctl2 3.27e-21
C503 sky130_fd_sc_hd__inv_2_6.Y sky130_fd_sc_hd__inv_2_5.Y 5.1e-21
C504 out carray_0.unitcap_247.cn 0.51f
C505 carray_0.unitcap_326.cn sky130_fd_sc_hd__inv_2_7.VPB 0.00109f
C506 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y sky130_fd_sc_hd__inv_2_2.Y 0.402f
C507 carray_0.unitcap_167.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C508 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y sky130_fd_sc_hd__inv_2_2.Y 0.358f
C509 ctl4 sky130_fd_sc_hd__inv_2_1.Y 3.6e-21
C510 out carray_0.unitcap_321.cn 0.512f
C511 sky130_fd_sc_hd__inv_2_0.Y carray_0.unitcap_184.cn 0.18f
C512 carray_0.unitcap_55.cn carray_0.unitcap_63.cn 0.0902f
C513 carray_0.unitcap_223.cn carray_0.unitcap_247.cn 0.0902f
C514 sky130_fd_sc_hd__inv_2_2.Y carray_0.unitcap_103.cn 0.18f
C515 carray_0.unitcap_322.cn carray_0.unitcap_328.cn 0.18f
C516 carray_0.unitcap_143.cn carray_0.unitcap_119.cn 0.0902f
C517 sky130_fd_sc_hd__inv_2_0.Y sky130_fd_sc_hd__inv_2_5.Y 0.108f
C518 out sw_top_0.sky130_fd_sc_hd__inv_4_0.Y 0.333f
C519 carray_0.unitcap_324.cn carray_0.unitcap_322.cn 0.18f
C520 out carray_0.unitcap_167.cn 0.51f
C521 out ctl3 8.03e-19
C522 carray_0.unitcap_334.cn sky130_fd_sc_hd__inv_2_4.Y 2.28e-19
C523 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y sky130_fd_sc_hd__inv_2_2.Y 1.15f
C524 sky130_fd_sc_hd__inv_2_4.Y ctl2 0.0488f
C525 out sw_top_2.sky130_fd_sc_hd__inv_4_0.Y 0.324f
C526 sky130_fd_sc_hd__inv_2_4.Y sky130_fd_sc_hd__inv_2_1.Y 7.78e-22
C527 sky130_fd_sc_hd__inv_2_1.Y ctl6 0.159f
C528 carray_0.unitcap_120.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C529 out carray_0.unitcap_103.cn 0.51f
C530 carray_0.unitcap_56.cn vdd 0.00108f
C531 carray_0.unitcap_232.cn carray_0.unitcap_248.cn 0.0902f
C532 sky130_fd_sc_hd__inv_2_3.Y sky130_fd_sc_hd__inv_2_2.Y 0.134f
C533 out carray_0.unitcap_224.cn 0.514f
C534 carray_0.unitcap_256.cn vdd 5.2e-19
C535 carray_0.unitcap_288.cn sky130_fd_sc_hd__inv_2_2.Y 0.0902f
C536 out sw_top_3.sky130_fd_sc_hd__inv_4_1.Y 0.692f
C537 sky130_fd_sc_hd__inv_2_8.Y ctl2 4.16e-20
C538 carray_0.unitcap_334.cn sky130_fd_sc_hd__inv_2_8.Y 0.0414f
C539 carray_0.unitcap_64.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C540 out carray_0.unitcap_120.cn 0.514f
C541 carray_0.unitcap_72.cn carray_0.unitcap_80.cn 0.0902f
C542 sky130_fd_sc_hd__inv_2_8.Y sky130_fd_sc_hd__inv_2_1.Y 0.663f
C543 ctl0 ctl3 1.18e-19
C544 carray_0.unitcap_160.cn carray_0.unitcap_144.cn 0.0902f
C545 ctl1 ctl2 0.0956f
C546 sample sw_top_1.sky130_fd_sc_hd__inv_4_0.Y 0.037f
C547 carray_0.unitcap_330.cn sky130_fd_sc_hd__inv_2_0.Y 0.039f
C548 carray_0.unitcap_87.cn sky130_fd_sc_hd__inv_2_2.Y 0.18f
C549 out ctl5 6.9e-19
C550 ctl4 sky130_fd_sc_hd__inv_2_4.Y 2.13e-20
C551 out sky130_fd_sc_hd__inv_2_3.Y 4.38f
C552 carray_0.unitcap_338.cn sky130_fd_sc_hd__inv_2_2.Y 0.161f
C553 carray_0.unitcap_95.cn carray_0.unitcap_111.cn 0.0902f
C554 out carray_0.unitcap_288.cn 0.558f
C555 ctl4 ctl6 1.34e-20
C556 out carray_0.unitcap_64.cn 0.514f
C557 carray_0.unitcap_16.cn sample 0.00246f
C558 sky130_fd_sc_hd__inv_2_7.Y sky130_fd_sc_hd__inv_2_7.VPB 0.0103f
C559 out carray_0.unitcap_87.cn 0.51f
C560 out carray_0.unitcap_338.cn 0.51f
C561 sky130_fd_sc_hd__inv_2_8.Y ctl4 0.16f
C562 sample sw_top_3.sky130_fd_sc_hd__inv_4_0.Y 0.037f
C563 sky130_fd_sc_hd__inv_2_4.Y ctl6 1.36e-21
C564 sky130_fd_sc_hd__inv_2_0.Y ctl7 3.81e-19
C565 carray_0.unitcap_326.cn sky130_fd_sc_hd__inv_2_5.Y 0.34f
C566 carray_0.unitcap_208.cn carray_0.unitcap_224.cn 0.0902f
C567 carray_0.unitcap_328.cn sky130_fd_sc_hd__inv_2_7.VPB 0.00105f
C568 dum vss 0.421f
C569 ctl0 vss 0.328f
C570 ctl1 vss 0.329f
C571 ctl2 vss 0.325f
C572 ctl3 vss 0.325f
C573 sample vss 5.61f
C574 ctl4 vss 0.325f
C575 ctl5 vss 0.324f
C576 ctl6 vss 0.323f
C577 ctl7 vss 0.387f
C578 vdd vss 39.6f
C579 out vss 52.7f
C580 vin vss 4.49f
C581 carray_0.unitcap_320.cn vss 0.267f
C582 carray_0.unitcap_321.cn vss 0.201f
C583 carray_0.unitcap_248.cn vss 0.201f
C584 carray_0.unitcap_232.cn vss 0.201f
C585 carray_0.unitcap_240.cn vss 0.201f
C586 carray_0.unitcap_216.cn vss 0.201f
C587 carray_0.unitcap_224.cn vss 0.201f
C588 carray_0.unitcap_208.cn vss 0.201f
C589 carray_0.unitcap_184.cn vss 0.201f
C590 carray_0.unitcap_200.cn vss 0.201f
C591 carray_0.unitcap_192.cn vss 0.201f
C592 carray_0.unitcap_168.cn vss 0.201f
C593 carray_0.unitcap_176.cn vss 0.201f
C594 carray_0.unitcap_160.cn vss 0.201f
C595 carray_0.unitcap_144.cn vss 0.201f
C596 carray_0.unitcap_152.cn vss 0.201f
C597 carray_0.unitcap_128.cn vss 0.201f
C598 carray_0.unitcap_136.cn vss 0.201f
C599 carray_0.unitcap_112.cn vss 0.201f
C600 carray_0.unitcap_120.cn vss 0.201f
C601 carray_0.unitcap_96.cn vss 0.201f
C602 carray_0.unitcap_104.cn vss 0.201f
C603 carray_0.unitcap_88.cn vss 0.201f
C604 carray_0.unitcap_64.cn vss 0.206f
C605 carray_0.unitcap_80.cn vss 0.206f
C606 carray_0.unitcap_72.cn vss 0.206f
C607 carray_0.unitcap_48.cn vss 0.206f
C608 carray_0.unitcap_56.cn vss 0.206f
C609 carray_0.unitcap_32.cn vss 0.206f
C610 carray_0.unitcap_40.cn vss 0.206f
C611 carray_0.unitcap_0.cn vss 0.206f
C612 carray_0.unitcap_24.cn vss 0.206f
C613 carray_0.unitcap_16.cn vss 0.206f
C614 carray_0.unitcap_8.cn vss 0.274f
C615 carray_0.unitcap_324.cn vss 0.165f
C616 carray_0.unitcap_9.cn vss 0.198f
C617 carray_0.unitcap_322.cn vss 0.161f
C618 carray_0.unitcap_256.cn vss 0.234f
C619 carray_0.unitcap_328.cn vss 0.159f
C620 carray_0.unitcap_288.cn vss 0.177f
C621 carray_0.unitcap_326.cn vss 0.152f
C622 carray_0.unitcap_10.cn vss 0.182f
C623 carray_0.unitcap_334.cn vss 0.154f
C624 carray_0.unitcap_11.cn vss 0.184f
C625 carray_0.unitcap_331.cn vss 0.171f
C626 carray_0.unitcap_13.cn vss 0.189f
C627 carray_0.unitcap_330.cn vss 0.175f
C628 carray_0.unitcap_12.cn vss 0.189f
C629 carray_0.unitcap_337.cn vss 0.175f
C630 carray_0.unitcap_14.cn vss 0.189f
C631 carray_0.unitcap_336.cn vss 0.265f
C632 carray_0.unitcap_338.cn vss 0.196f
C633 carray_0.unitcap_255.cn vss 0.196f
C634 carray_0.unitcap_239.cn vss 0.196f
C635 carray_0.unitcap_247.cn vss 0.196f
C636 carray_0.unitcap_223.cn vss 0.196f
C637 carray_0.unitcap_231.cn vss 0.196f
C638 carray_0.unitcap_215.cn vss 0.196f
C639 carray_0.unitcap_191.cn vss 0.196f
C640 carray_0.unitcap_207.cn vss 0.196f
C641 carray_0.unitcap_199.cn vss 0.196f
C642 carray_0.unitcap_175.cn vss 0.196f
C643 carray_0.unitcap_183.cn vss 0.196f
C644 carray_0.unitcap_167.cn vss 0.196f
C645 carray_0.unitcap_151.cn vss 0.196f
C646 carray_0.unitcap_159.cn vss 0.196f
C647 carray_0.unitcap_135.cn vss 0.196f
C648 carray_0.unitcap_143.cn vss 0.201f
C649 carray_0.unitcap_119.cn vss 0.201f
C650 carray_0.unitcap_127.cn vss 0.201f
C651 carray_0.unitcap_103.cn vss 0.201f
C652 carray_0.unitcap_111.cn vss 0.201f
C653 carray_0.unitcap_95.cn vss 0.201f
C654 carray_0.unitcap_71.cn vss 0.201f
C655 carray_0.unitcap_87.cn vss 0.201f
C656 carray_0.unitcap_79.cn vss 0.201f
C657 carray_0.unitcap_55.cn vss 0.201f
C658 carray_0.unitcap_63.cn vss 0.201f
C659 carray_0.unitcap_39.cn vss 0.201f
C660 carray_0.unitcap_47.cn vss 0.201f
C661 carray_0.unitcap_7.cn vss 0.201f
C662 carray_0.unitcap_31.cn vss 0.201f
C663 carray_0.unitcap_23.cn vss 0.201f
C664 carray_0.unitcap_15.cn vss 0.271f
C665 sky130_fd_sc_hd__inv_2_7.Y vss 1.02f
C666 sky130_fd_sc_hd__inv_2_6.Y vss 0.775f
C667 sky130_fd_sc_hd__inv_2_4.Y vss 1.12f
C668 sky130_fd_sc_hd__inv_2_5.Y vss 2.83f
C669 sky130_fd_sc_hd__inv_2_3.Y vss 4.97f
C670 sky130_fd_sc_hd__inv_2_8.Y vss 3.82f
C671 sky130_fd_sc_hd__inv_2_0.Y vss 29.1f
C672 sky130_fd_sc_hd__inv_2_1.Y vss 55.1f
C673 sw_top_0.sky130_fd_sc_hd__inv_4_0.Y vss 1.99f
C674 sw_top_1.sky130_fd_sc_hd__inv_4_0.Y vss 1.97f
C675 sw_top_3.sky130_fd_sc_hd__inv_4_0.Y vss 1.97f
C676 sw_top_2.sky130_fd_sc_hd__inv_4_0.Y vss 1.97f
C677 sky130_fd_sc_hd__inv_2_2.Y vss 0.119p
C678 sw_top_0.sky130_fd_sc_hd__inv_4_1.Y vss 1.86f
C679 sw_top_1.sky130_fd_sc_hd__inv_4_1.Y vss 1.61f
C680 sw_top_3.sky130_fd_sc_hd__inv_4_1.Y vss 1.61f
C681 sw_top_2.sky130_fd_sc_hd__inv_4_1.Y vss 1.7f
C682 sky130_fd_sc_hd__inv_2_7.VPB vss 3.01f
C683 sky130_fd_sc_hd__inv_2_5.Y.t0 vss 0.567f
C684 sky130_fd_sc_hd__inv_2_5.Y.t4 vss 0.00262f
C685 sky130_fd_sc_hd__inv_2_5.Y.t3 vss 0.00262f
C686 sky130_fd_sc_hd__inv_2_5.Y.n0 vss 0.00621f
C687 sky130_fd_sc_hd__inv_2_5.Y.n1 vss 0.00372f
C688 sky130_fd_sc_hd__inv_2_5.Y.n2 vss 0.0769f
C689 sky130_fd_sc_hd__inv_2_5.Y.t2 vss 0.00404f
C690 sky130_fd_sc_hd__inv_2_5.Y.t1 vss 0.00404f
C691 sky130_fd_sc_hd__inv_2_5.Y.n3 vss 0.0103f
C692 sky130_fd_sc_hd__inv_2_5.Y.n4 vss 0.0178f
C693 sky130_fd_sc_hd__inv_2_0.Y.t3 vss 0.00743f
C694 sky130_fd_sc_hd__inv_2_0.Y.t1 vss 0.00743f
C695 sky130_fd_sc_hd__inv_2_0.Y.n0 vss 0.019f
C696 sky130_fd_sc_hd__inv_2_0.Y.n1 vss 0.0328f
C697 sky130_fd_sc_hd__inv_2_0.Y.t4 vss 0.00483f
C698 sky130_fd_sc_hd__inv_2_0.Y.t2 vss 0.00483f
C699 sky130_fd_sc_hd__inv_2_0.Y.n2 vss 0.0114f
C700 sky130_fd_sc_hd__inv_2_0.Y.n3 vss 0.00686f
C701 sky130_fd_sc_hd__inv_2_0.Y.n4 vss 0.225f
C702 sky130_fd_sc_hd__inv_2_0.Y.n5 vss 0.708f
C703 sky130_fd_sc_hd__inv_2_0.Y.t0 vss 0.543f
C704 sky130_fd_sc_hd__inv_2_0.Y.n6 vss -0.821f
C705 sky130_fd_sc_hd__inv_2_3.Y.t1 vss 0.831f
C706 sky130_fd_sc_hd__inv_2_3.Y.t0 vss 0.809f
C707 sky130_fd_sc_hd__inv_2_3.Y.t3 vss 0.00331f
C708 sky130_fd_sc_hd__inv_2_3.Y.t5 vss 0.00331f
C709 sky130_fd_sc_hd__inv_2_3.Y.n0 vss 0.00784f
C710 sky130_fd_sc_hd__inv_2_3.Y.n1 vss 0.0047f
C711 sky130_fd_sc_hd__inv_2_3.Y.n2 vss 0.123f
C712 sky130_fd_sc_hd__inv_2_3.Y.t2 vss 0.0051f
C713 sky130_fd_sc_hd__inv_2_3.Y.t4 vss 0.0051f
C714 sky130_fd_sc_hd__inv_2_3.Y.n3 vss 0.013f
C715 sky130_fd_sc_hd__inv_2_3.Y.n4 vss 0.0225f
C716 sample.n0 vss 0.00813f
C717 sample.n1 vss 0.00431f
C718 sample.n2 vss 0.00595f
C719 sample.n3 vss 0.00225f
C720 sample.t26 vss 0.0151f
C721 sample.t11 vss 0.00892f
C722 sample.t6 vss 0.0151f
C723 sample.t22 vss 0.00892f
C724 sample.n4 vss 0.0218f
C725 sample.t24 vss 0.0151f
C726 sample.t8 vss 0.00892f
C727 sample.t9 vss 0.0151f
C728 sample.t27 vss 0.00892f
C729 sample.n5 vss 0.0204f
C730 sample.n6 vss 0.0102f
C731 sample.n7 vss 0.0218f
C732 sample.n8 vss 0.00999f
C733 sample.n9 vss 0.00829f
C734 sample.n10 vss 0.00829f
C735 sample.n11 vss 0.00999f
C736 sample.n12 vss 0.0253f
C737 sample.n13 vss 0.013f
C738 sample.n14 vss 0.00171f
C739 sample.n15 vss 0.00412f
C740 sample.n16 vss 0.00178f
C741 sample.n17 vss 0.0018f
C742 sample.n18 vss 0.0224f
C743 sample.n19 vss 0.00813f
C744 sample.n20 vss 0.00429f
C745 sample.n21 vss 0.00178f
C746 sample.n22 vss 0.00597f
C747 sample.n23 vss 0.00412f
C748 sample.n24 vss 0.00225f
C749 sample.t17 vss 0.0151f
C750 sample.t2 vss 0.00892f
C751 sample.t4 vss 0.0151f
C752 sample.t20 vss 0.00892f
C753 sample.n25 vss 0.0218f
C754 sample.t13 vss 0.0151f
C755 sample.t30 vss 0.00892f
C756 sample.t1 vss 0.0151f
C757 sample.t18 vss 0.00892f
C758 sample.n26 vss 0.0204f
C759 sample.n27 vss 0.0102f
C760 sample.n28 vss 0.0218f
C761 sample.n29 vss 0.00999f
C762 sample.n30 vss 0.00829f
C763 sample.n31 vss 0.00829f
C764 sample.n32 vss 0.00999f
C765 sample.n33 vss 0.0253f
C766 sample.n34 vss 0.013f
C767 sample.n35 vss 0.00171f
C768 sample.n36 vss 0.0018f
C769 sample.n37 vss 0.0231f
C770 sample.n38 vss 0.00813f
C771 sample.n39 vss 0.00429f
C772 sample.n40 vss 0.00178f
C773 sample.n41 vss 0.00597f
C774 sample.n42 vss 0.00412f
C775 sample.n43 vss 0.00225f
C776 sample.t15 vss 0.0151f
C777 sample.t31 vss 0.00892f
C778 sample.t25 vss 0.0151f
C779 sample.t10 vss 0.00892f
C780 sample.n44 vss 0.0218f
C781 sample.t5 vss 0.0151f
C782 sample.t21 vss 0.00892f
C783 sample.t23 vss 0.0151f
C784 sample.t7 vss 0.00892f
C785 sample.n45 vss 0.0204f
C786 sample.n46 vss 0.0102f
C787 sample.n47 vss 0.0218f
C788 sample.n48 vss 0.00999f
C789 sample.n49 vss 0.00829f
C790 sample.n50 vss 0.00829f
C791 sample.n51 vss 0.00999f
C792 sample.n52 vss 0.0253f
C793 sample.n53 vss 0.013f
C794 sample.n54 vss 0.00171f
C795 sample.n55 vss 0.0018f
C796 sample.n56 vss 0.0231f
C797 sample.n57 vss 0.00813f
C798 sample.n58 vss 0.00429f
C799 sample.n59 vss 0.00178f
C800 sample.n60 vss 0.00597f
C801 sample.n61 vss 0.00412f
C802 sample.n62 vss 0.00225f
C803 sample.t28 vss 0.0151f
C804 sample.t14 vss 0.00892f
C805 sample.t16 vss 0.0151f
C806 sample.t0 vss 0.00892f
C807 sample.n63 vss 0.0218f
C808 sample.t3 vss 0.0151f
C809 sample.t19 vss 0.00892f
C810 sample.t12 vss 0.0151f
C811 sample.t29 vss 0.00892f
C812 sample.n64 vss 0.0204f
C813 sample.n65 vss 0.0102f
C814 sample.n66 vss 0.0218f
C815 sample.n67 vss 0.00999f
C816 sample.n68 vss 0.00829f
C817 sample.n69 vss 0.00829f
C818 sample.n70 vss 0.00999f
C819 sample.n71 vss 0.0253f
C820 sample.n72 vss 0.013f
C821 sample.n73 vss 0.00171f
C822 sample.n74 vss 0.0018f
C823 sample.n75 vss 0.0248f
C824 sample.n76 vss 0.164f
C825 sample.n77 vss 0.164f
C826 sample.n78 vss 0.165f
C827 vdd.n0 vss 0.00657f
C828 vdd.n1 vss 0.00973f
C829 vdd.n2 vss 0.0138f
C830 vdd.t22 vss 0.0634f
C831 vdd.n3 vss 0.00949f
C832 vdd.n4 vss 0.00455f
C833 vdd.n5 vss 0.00834f
C834 vdd.n6 vss 0.00142f
C835 vdd.t19 vss 0.0061f
C836 vdd.n7 vss 0.0049f
C837 vdd.t13 vss 0.0015f
C838 vdd.t140 vss 0.0015f
C839 vdd.n8 vss 0.0034f
C840 vdd.t113 vss 0.0061f
C841 vdd.n9 vss 0.00846f
C842 vdd.n10 vss 0.0049f
C843 vdd.t116 vss 0.0015f
C844 vdd.t106 vss 0.0015f
C845 vdd.n11 vss 0.0034f
C846 vdd.t118 vss 0.00498f
C847 vdd.n12 vss 0.00496f
C848 vdd.n13 vss 0.00107f
C849 vdd.n14 vss 0.0188f
C850 vdd.n15 vss 5.76e-19
C851 vdd.n16 vss 0.0151f
C852 vdd.t120 vss 0.0279f
C853 vdd.n17 vss 0.00889f
C854 vdd.t111 vss 0.0372f
C855 vdd.t109 vss 0.0372f
C856 vdd.t103 vss 0.0372f
C857 vdd.t110 vss 0.0459f
C858 vdd.n18 vss 0.0749f
C859 vdd.n19 vss 0.0364f
C860 vdd.n20 vss 0.0186f
C861 vdd.t108 vss 0.0279f
C862 vdd.t119 vss 0.0372f
C863 vdd.t107 vss 0.0372f
C864 vdd.t114 vss 0.0372f
C865 vdd.t104 vss 0.0457f
C866 vdd.n21 vss 0.0273f
C867 vdd.n22 vss 0.0026f
C868 vdd.n24 vss 9.72e-19
C869 vdd.n25 vss 0.0049f
C870 vdd.t151 vss 0.00829f
C871 vdd.n26 vss 0.00629f
C872 vdd.n27 vss 0.00973f
C873 vdd.n28 vss 0.0138f
C874 vdd.t43 vss 0.00373f
C875 vdd.n29 vss 0.0143f
C876 vdd.n30 vss 0.0466f
C877 vdd.t50 vss 0.0399f
C878 vdd.t121 vss 0.0252f
C879 vdd.t128 vss 0.0195f
C880 vdd.t134 vss 0.0195f
C881 vdd.t126 vss 0.0185f
C882 vdd.t10 vss 0.0244f
C883 vdd.t2 vss 0.0195f
C884 vdd.t16 vss 0.0195f
C885 vdd.t8 vss 0.0185f
C886 vdd.t53 vss 0.0634f
C887 vdd.n31 vss 0.00949f
C888 vdd.n32 vss 0.00455f
C889 vdd.n33 vss 0.00834f
C890 vdd.n34 vss 0.00142f
C891 vdd.t9 vss 0.0061f
C892 vdd.n35 vss 0.0049f
C893 vdd.t3 vss 0.0015f
C894 vdd.t17 vss 0.0015f
C895 vdd.n36 vss 0.0034f
C896 vdd.t127 vss 0.0061f
C897 vdd.n37 vss 0.00846f
C898 vdd.n38 vss 0.0049f
C899 vdd.t129 vss 0.0015f
C900 vdd.t135 vss 0.0015f
C901 vdd.n39 vss 0.0034f
C902 vdd.t122 vss 0.00498f
C903 vdd.n40 vss 0.00496f
C904 vdd.n41 vss 0.00107f
C905 vdd.n42 vss 0.0188f
C906 vdd.n43 vss 5.76e-19
C907 vdd.n44 vss 0.0151f
C908 vdd.t131 vss 0.0279f
C909 vdd.n45 vss 0.00889f
C910 vdd.t137 vss 0.0372f
C911 vdd.t138 vss 0.0372f
C912 vdd.t132 vss 0.0372f
C913 vdd.t125 vss 0.0459f
C914 vdd.n46 vss 0.0749f
C915 vdd.n47 vss 0.0364f
C916 vdd.n48 vss 0.0186f
C917 vdd.t124 vss 0.0279f
C918 vdd.t130 vss 0.0372f
C919 vdd.t136 vss 0.0372f
C920 vdd.t123 vss 0.0372f
C921 vdd.t133 vss 0.0457f
C922 vdd.n49 vss 0.0273f
C923 vdd.n50 vss 0.0026f
C924 vdd.n52 vss 9.72e-19
C925 vdd.n53 vss 0.0049f
C926 vdd.t153 vss 0.00829f
C927 vdd.n54 vss 0.00368f
C928 vdd.n55 vss 0.00519f
C929 vdd.t51 vss 0.00366f
C930 vdd.n56 vss 0.00297f
C931 vdd.n57 vss 0.0136f
C932 vdd.n58 vss 0.0108f
C933 vdd.t52 vss 0.00366f
C934 vdd.n59 vss 0.00779f
C935 vdd.n60 vss 0.00481f
C936 vdd.n61 vss 0.0025f
C937 vdd.n62 vss 0.00867f
C938 vdd.n63 vss 0.00368f
C939 vdd.n64 vss 0.0049f
C940 vdd.n65 vss 0.00142f
C941 vdd.n66 vss 0.00435f
C942 vdd.n67 vss 0.00142f
C943 vdd.n68 vss 0.0049f
C944 vdd.n69 vss 0.0029f
C945 vdd.n70 vss 0.00349f
C946 vdd.t11 vss 0.00498f
C947 vdd.n71 vss 0.00481f
C948 vdd.n72 vss 0.00142f
C949 vdd.n73 vss 0.00435f
C950 vdd.n74 vss 0.0049f
C951 vdd.n75 vss 0.0049f
C952 vdd.n76 vss 0.0029f
C953 vdd.n77 vss 0.00832f
C954 vdd.n78 vss 0.0113f
C955 vdd.n79 vss 0.0109f
C956 vdd.t146 vss 0.027f
C957 vdd.t54 vss 0.00363f
C958 vdd.n80 vss 0.0565f
C959 vdd.n81 vss 0.0175f
C960 vdd.n82 vss 0.0138f
C961 vdd.n83 vss 0.00973f
C962 vdd.n84 vss 0.00654f
C963 vdd.n85 vss 0.0025f
C964 vdd.t148 vss 0.00829f
C965 vdd.t45 vss 0.00366f
C966 vdd.n86 vss 0.00297f
C967 vdd.n87 vss 0.0136f
C968 vdd.t46 vss 0.00366f
C969 vdd.n88 vss 0.00107f
C970 vdd.n89 vss 0.0188f
C971 vdd.n90 vss 5.76e-19
C972 vdd.n91 vss 0.0151f
C973 vdd.t68 vss 0.0279f
C974 vdd.n92 vss 0.00889f
C975 vdd.t79 vss 0.0372f
C976 vdd.t69 vss 0.0372f
C977 vdd.t70 vss 0.0372f
C978 vdd.t78 vss 0.0459f
C979 vdd.n93 vss 0.0749f
C980 vdd.n94 vss 0.0364f
C981 vdd.n95 vss 0.0186f
C982 vdd.t75 vss 0.0279f
C983 vdd.t67 vss 0.0372f
C984 vdd.t72 vss 0.0372f
C985 vdd.t64 vss 0.0372f
C986 vdd.t71 vss 0.0457f
C987 vdd.n96 vss 0.0273f
C988 vdd.n97 vss 0.0026f
C989 vdd.n99 vss 9.72e-19
C990 vdd.n100 vss 0.00867f
C991 vdd.n101 vss 0.00368f
C992 vdd.t74 vss 0.00498f
C993 vdd.t66 vss 0.0015f
C994 vdd.t77 vss 0.0015f
C995 vdd.n102 vss 0.0034f
C996 vdd.n103 vss 0.00435f
C997 vdd.n104 vss 0.0029f
C998 vdd.t63 vss 0.0061f
C999 vdd.n105 vss 0.00349f
C1000 vdd.t6 vss 0.00498f
C1001 vdd.t142 vss 0.0015f
C1002 vdd.t38 vss 0.0015f
C1003 vdd.n106 vss 0.0034f
C1004 vdd.n107 vss 0.00435f
C1005 vdd.n108 vss 0.0029f
C1006 vdd.t42 vss 0.00363f
C1007 vdd.t147 vss 0.027f
C1008 vdd.n109 vss 0.0565f
C1009 vdd.n110 vss 0.0175f
C1010 vdd.n111 vss 0.0109f
C1011 vdd.n112 vss 0.00834f
C1012 vdd.n113 vss 0.0113f
C1013 vdd.t34 vss 0.0061f
C1014 vdd.n114 vss 0.00832f
C1015 vdd.n115 vss 0.00142f
C1016 vdd.n116 vss 0.0049f
C1017 vdd.n117 vss 0.0049f
C1018 vdd.n118 vss 0.0049f
C1019 vdd.n119 vss 0.00142f
C1020 vdd.n120 vss 0.00481f
C1021 vdd.n121 vss 0.00846f
C1022 vdd.n122 vss 0.00142f
C1023 vdd.n123 vss 0.0049f
C1024 vdd.n124 vss 0.0049f
C1025 vdd.n125 vss 0.0049f
C1026 vdd.n126 vss 0.00142f
C1027 vdd.n127 vss 0.00496f
C1028 vdd.n128 vss 0.00481f
C1029 vdd.n129 vss 0.00779f
C1030 vdd.n130 vss 0.0108f
C1031 vdd.n131 vss 0.0049f
C1032 vdd.n132 vss 0.00368f
C1033 vdd.n133 vss 0.00404f
C1034 vdd.n134 vss 0.00629f
C1035 vdd.t55 vss 0.00373f
C1036 vdd.n135 vss 0.0143f
C1037 vdd.n136 vss 0.016f
C1038 vdd.n137 vss 0.0429f
C1039 vdd.t44 vss 0.0321f
C1040 vdd.t73 vss 0.0252f
C1041 vdd.t65 vss 0.0195f
C1042 vdd.t76 vss 0.0195f
C1043 vdd.t62 vss 0.0185f
C1044 vdd.t5 vss 0.0244f
C1045 vdd.t141 vss 0.0195f
C1046 vdd.t37 vss 0.0195f
C1047 vdd.t33 vss 0.0185f
C1048 vdd.t41 vss 0.0634f
C1049 vdd.t18 vss 0.0185f
C1050 vdd.t139 vss 0.0195f
C1051 vdd.t12 vss 0.0195f
C1052 vdd.t14 vss 0.0244f
C1053 vdd.t112 vss 0.0185f
C1054 vdd.t105 vss 0.0195f
C1055 vdd.t115 vss 0.0195f
C1056 vdd.t117 vss 0.0252f
C1057 vdd.t25 vss 0.0321f
C1058 vdd.n138 vss 0.0429f
C1059 vdd.n139 vss 0.016f
C1060 vdd.n140 vss 0.00949f
C1061 vdd.n141 vss 0.00654f
C1062 vdd.n142 vss 0.00404f
C1063 vdd.n143 vss 0.00368f
C1064 vdd.n144 vss 0.00455f
C1065 vdd.t26 vss 0.00366f
C1066 vdd.n145 vss 0.00297f
C1067 vdd.n146 vss 0.0136f
C1068 vdd.n147 vss 0.0108f
C1069 vdd.t27 vss 0.00366f
C1070 vdd.n148 vss 0.00779f
C1071 vdd.n149 vss 0.00481f
C1072 vdd.n150 vss 0.0025f
C1073 vdd.n151 vss 0.00867f
C1074 vdd.n152 vss 0.00368f
C1075 vdd.n153 vss 0.0049f
C1076 vdd.n154 vss 0.00142f
C1077 vdd.n155 vss 0.00435f
C1078 vdd.n156 vss 0.00142f
C1079 vdd.n157 vss 0.0049f
C1080 vdd.n158 vss 0.0029f
C1081 vdd.n159 vss 0.00349f
C1082 vdd.t15 vss 0.00498f
C1083 vdd.n160 vss 0.00481f
C1084 vdd.n161 vss 0.00142f
C1085 vdd.n162 vss 0.00435f
C1086 vdd.n163 vss 0.0049f
C1087 vdd.n164 vss 0.0049f
C1088 vdd.n165 vss 0.0029f
C1089 vdd.n166 vss 0.00832f
C1090 vdd.n167 vss 0.0113f
C1091 vdd.n168 vss 0.0109f
C1092 vdd.t150 vss 0.027f
C1093 vdd.t23 vss 0.00363f
C1094 vdd.n169 vss 0.0565f
C1095 vdd.n170 vss 0.0175f
C1096 vdd.n171 vss 0.0138f
C1097 vdd.n172 vss 0.00973f
C1098 vdd.n173 vss 0.00654f
C1099 vdd.n174 vss 0.0025f
C1100 vdd.t152 vss 0.00829f
C1101 vdd.t29 vss 0.00366f
C1102 vdd.n175 vss 0.00297f
C1103 vdd.n176 vss 0.0136f
C1104 vdd.t30 vss 0.00366f
C1105 vdd.n177 vss 0.00107f
C1106 vdd.n178 vss 0.0026f
C1107 vdd.n179 vss 0.0749f
C1108 vdd.n180 vss 5.76e-19
C1109 vdd.n181 vss 0.0273f
C1110 vdd.t89 vss 0.0457f
C1111 vdd.t83 vss 0.0372f
C1112 vdd.t97 vss 0.0372f
C1113 vdd.t92 vss 0.0372f
C1114 vdd.t84 vss 0.0279f
C1115 vdd.t80 vss 0.0459f
C1116 vdd.t86 vss 0.0372f
C1117 vdd.t94 vss 0.0372f
C1118 vdd.t85 vss 0.0372f
C1119 vdd.t93 vss 0.0279f
C1120 vdd.n182 vss 0.0186f
C1121 vdd.n183 vss 0.0364f
C1122 vdd.n184 vss 0.00889f
C1123 vdd.n185 vss 0.0151f
C1124 vdd.n186 vss 0.0188f
C1125 vdd.n188 vss 9.72e-19
C1126 vdd.n189 vss 0.00867f
C1127 vdd.n190 vss 0.00368f
C1128 vdd.t91 vss 0.00498f
C1129 vdd.t82 vss 0.0015f
C1130 vdd.t96 vss 0.0015f
C1131 vdd.n191 vss 0.0034f
C1132 vdd.n192 vss 0.00435f
C1133 vdd.n193 vss 0.0029f
C1134 vdd.t88 vss 0.0061f
C1135 vdd.n194 vss 0.00349f
C1136 vdd.t21 vss 0.00498f
C1137 vdd.t36 vss 0.0015f
C1138 vdd.t99 vss 0.0015f
C1139 vdd.n195 vss 0.0034f
C1140 vdd.n196 vss 0.00435f
C1141 vdd.n197 vss 0.0029f
C1142 vdd.t48 vss 0.00363f
C1143 vdd.t149 vss 0.027f
C1144 vdd.n198 vss 0.0565f
C1145 vdd.n199 vss 0.0175f
C1146 vdd.n200 vss 0.0109f
C1147 vdd.n201 vss 0.00834f
C1148 vdd.n202 vss 0.0113f
C1149 vdd.t102 vss 0.0061f
C1150 vdd.n203 vss 0.00832f
C1151 vdd.n204 vss 0.00142f
C1152 vdd.n205 vss 0.0049f
C1153 vdd.n206 vss 0.0049f
C1154 vdd.n207 vss 0.0049f
C1155 vdd.n208 vss 0.00142f
C1156 vdd.n209 vss 0.00481f
C1157 vdd.n210 vss 0.00846f
C1158 vdd.n211 vss 0.00142f
C1159 vdd.n212 vss 0.0049f
C1160 vdd.n213 vss 0.0049f
C1161 vdd.n214 vss 0.0049f
C1162 vdd.n215 vss 0.00142f
C1163 vdd.n216 vss 0.00496f
C1164 vdd.n217 vss 0.00481f
C1165 vdd.n218 vss 0.00779f
C1166 vdd.n219 vss 0.0108f
C1167 vdd.n220 vss 0.0049f
C1168 vdd.n221 vss 0.00368f
C1169 vdd.n222 vss 0.00404f
C1170 vdd.n223 vss 0.00629f
C1171 vdd.t24 vss 0.00373f
C1172 vdd.n224 vss 0.0143f
C1173 vdd.n225 vss 0.016f
C1174 vdd.n226 vss 0.0429f
C1175 vdd.t28 vss 0.0321f
C1176 vdd.t90 vss 0.0252f
C1177 vdd.t81 vss 0.0195f
C1178 vdd.t95 vss 0.0195f
C1179 vdd.t87 vss 0.0185f
C1180 vdd.t20 vss 0.0244f
C1181 vdd.t35 vss 0.0195f
C1182 vdd.t98 vss 0.0195f
C1183 vdd.t101 vss 0.0185f
C1184 vdd.t47 vss 0.0634f
C1185 vdd.n227 vss 0.0332f
C1186 vdd.n228 vss 0.0429f
C1187 vdd.t49 vss 0.00373f
C1188 vdd.n229 vss 0.0143f
C1189 vdd.n230 vss 0.016f
C1190 vdd.n231 vss 0.00949f
C1191 vdd.n232 vss 0.00653f
C1192 vdd.n233 vss 0.00406f
C1193 vdd.n234 vss 0.00115f
C1194 vdd.n235 vss 0.00559f
C1195 vin.t50 vss 0.0221f
C1196 vin.t29 vss 0.0244f
C1197 vin.t58 vss 0.0184f
C1198 vin.t54 vss 0.0184f
C1199 vin.n0 vss 0.129f
C1200 vin.t26 vss 0.0184f
C1201 vin.t23 vss 0.0184f
C1202 vin.n1 vss 0.129f
C1203 vin.t57 vss 0.0184f
C1204 vin.t53 vss 0.0184f
C1205 vin.n2 vss 0.129f
C1206 vin.t28 vss 0.0184f
C1207 vin.t22 vss 0.0184f
C1208 vin.n3 vss 0.129f
C1209 vin.t56 vss 0.0184f
C1210 vin.t52 vss 0.0184f
C1211 vin.n4 vss 0.129f
C1212 vin.t24 vss 0.0184f
C1213 vin.t21 vss 0.0184f
C1214 vin.n5 vss 0.129f
C1215 vin.t51 vss 0.0184f
C1216 vin.t59 vss 0.0184f
C1217 vin.n6 vss 0.129f
C1218 vin.t20 vss 0.0184f
C1219 vin.t27 vss 0.0184f
C1220 vin.n7 vss 0.129f
C1221 vin.t55 vss 0.0222f
C1222 vin.t25 vss 0.0244f
C1223 vin.n8 vss 0.37f
C1224 vin.n9 vss 0.108f
C1225 vin.n10 vss 0.108f
C1226 vin.n11 vss 0.108f
C1227 vin.n12 vss 0.109f
C1228 vin.n13 vss 0.387f
C1229 vin.t65 vss 0.0221f
C1230 vin.t3 vss 0.0244f
C1231 vin.t64 vss 0.0184f
C1232 vin.t60 vss 0.0184f
C1233 vin.n14 vss 0.129f
C1234 vin.t0 vss 0.0184f
C1235 vin.t7 vss 0.0184f
C1236 vin.n15 vss 0.129f
C1237 vin.t69 vss 0.0184f
C1238 vin.t66 vss 0.0184f
C1239 vin.n16 vss 0.129f
C1240 vin.t6 vss 0.0184f
C1241 vin.t2 vss 0.0184f
C1242 vin.n17 vss 0.129f
C1243 vin.t68 vss 0.0184f
C1244 vin.t63 vss 0.0184f
C1245 vin.n18 vss 0.129f
C1246 vin.t5 vss 0.0184f
C1247 vin.t1 vss 0.0184f
C1248 vin.n19 vss 0.129f
C1249 vin.t67 vss 0.0184f
C1250 vin.t62 vss 0.0184f
C1251 vin.n20 vss 0.129f
C1252 vin.t4 vss 0.0184f
C1253 vin.t9 vss 0.0184f
C1254 vin.n21 vss 0.129f
C1255 vin.t61 vss 0.0222f
C1256 vin.t8 vss 0.0244f
C1257 vin.n22 vss 0.37f
C1258 vin.n23 vss 0.108f
C1259 vin.n24 vss 0.108f
C1260 vin.n25 vss 0.108f
C1261 vin.n26 vss 0.109f
C1262 vin.n27 vss 0.386f
C1263 vin.n28 vss 0.0818f
C1264 vin.t48 vss 0.0221f
C1265 vin.t16 vss 0.0244f
C1266 vin.t43 vss 0.0184f
C1267 vin.t44 vss 0.0184f
C1268 vin.n29 vss 0.129f
C1269 vin.t14 vss 0.0184f
C1270 vin.t11 vss 0.0184f
C1271 vin.n30 vss 0.129f
C1272 vin.t42 vss 0.0184f
C1273 vin.t49 vss 0.0184f
C1274 vin.n31 vss 0.129f
C1275 vin.t10 vss 0.0184f
C1276 vin.t17 vss 0.0184f
C1277 vin.n32 vss 0.129f
C1278 vin.t41 vss 0.0184f
C1279 vin.t47 vss 0.0184f
C1280 vin.n33 vss 0.129f
C1281 vin.t19 vss 0.0184f
C1282 vin.t13 vss 0.0184f
C1283 vin.n34 vss 0.129f
C1284 vin.t40 vss 0.0184f
C1285 vin.t46 vss 0.0184f
C1286 vin.n35 vss 0.129f
C1287 vin.t18 vss 0.0184f
C1288 vin.t15 vss 0.0184f
C1289 vin.n36 vss 0.129f
C1290 vin.t45 vss 0.0222f
C1291 vin.t12 vss 0.0244f
C1292 vin.n37 vss 0.37f
C1293 vin.n38 vss 0.108f
C1294 vin.n39 vss 0.108f
C1295 vin.n40 vss 0.108f
C1296 vin.n41 vss 0.109f
C1297 vin.n42 vss 0.386f
C1298 vin.n43 vss 0.0828f
C1299 vin.t72 vss 0.0221f
C1300 vin.t31 vss 0.0244f
C1301 vin.t79 vss 0.0184f
C1302 vin.t75 vss 0.0184f
C1303 vin.n44 vss 0.129f
C1304 vin.t38 vss 0.0184f
C1305 vin.t35 vss 0.0184f
C1306 vin.n45 vss 0.129f
C1307 vin.t74 vss 0.0184f
C1308 vin.t78 vss 0.0184f
C1309 vin.n46 vss 0.129f
C1310 vin.t34 vss 0.0184f
C1311 vin.t30 vss 0.0184f
C1312 vin.n47 vss 0.129f
C1313 vin.t73 vss 0.0184f
C1314 vin.t71 vss 0.0184f
C1315 vin.n48 vss 0.129f
C1316 vin.t33 vss 0.0184f
C1317 vin.t39 vss 0.0184f
C1318 vin.n49 vss 0.129f
C1319 vin.t70 vss 0.0184f
C1320 vin.t77 vss 0.0184f
C1321 vin.n50 vss 0.129f
C1322 vin.t32 vss 0.0184f
C1323 vin.t37 vss 0.0184f
C1324 vin.n51 vss 0.129f
C1325 vin.t76 vss 0.0222f
C1326 vin.t36 vss 0.0244f
C1327 vin.n52 vss 0.37f
C1328 vin.n53 vss 0.108f
C1329 vin.n54 vss 0.108f
C1330 vin.n55 vss 0.108f
C1331 vin.n56 vss 0.109f
C1332 vin.n57 vss 0.385f
C1333 vin.n58 vss 0.307f
C1334 vin.n59 vss 0.566f
C1335 vin.n60 vss 0.577f
C1336 vin.n61 vss 0.406f
C1337 sky130_fd_sc_hd__inv_2_2.Y.t3 vss 0.346f
C1338 sky130_fd_sc_hd__inv_2_2.Y.t2 vss 0.455f
C1339 sky130_fd_sc_hd__inv_2_2.Y.t0 vss 0.00726f
C1340 sky130_fd_sc_hd__inv_2_2.Y.t4 vss 0.00726f
C1341 sky130_fd_sc_hd__inv_2_2.Y.n0 vss 0.0186f
C1342 sky130_fd_sc_hd__inv_2_2.Y.n1 vss 0.032f
C1343 sky130_fd_sc_hd__inv_2_2.Y.t1 vss 0.00472f
C1344 sky130_fd_sc_hd__inv_2_2.Y.t5 vss 0.00472f
C1345 sky130_fd_sc_hd__inv_2_2.Y.n2 vss 0.0112f
C1346 sky130_fd_sc_hd__inv_2_2.Y.n3 vss 0.0067f
C1347 sky130_fd_sc_hd__inv_2_2.Y.n4 vss 0.382f
C1348 sky130_fd_sc_hd__inv_2_1.Y.n0 vss -0.225f
C1349 sky130_fd_sc_hd__inv_2_1.Y.n1 vss 0.421f
C1350 sky130_fd_sc_hd__inv_2_1.Y.t3 vss 0.00682f
C1351 sky130_fd_sc_hd__inv_2_1.Y.t4 vss 0.00682f
C1352 sky130_fd_sc_hd__inv_2_1.Y.n2 vss 0.0174f
C1353 sky130_fd_sc_hd__inv_2_1.Y.n3 vss 0.03f
C1354 sky130_fd_sc_hd__inv_2_1.Y.t1 vss 0.00443f
C1355 sky130_fd_sc_hd__inv_2_1.Y.t2 vss 0.00443f
C1356 sky130_fd_sc_hd__inv_2_1.Y.n4 vss 0.0105f
C1357 sky130_fd_sc_hd__inv_2_1.Y.n5 vss 0.00629f
C1358 sky130_fd_sc_hd__inv_2_1.Y.n6 vss 0.27f
C1359 sky130_fd_sc_hd__inv_2_1.Y.t0 vss 0.433f
C1360 out.n0 vss 0.00165f
C1361 out.t76 vss 0.00464f
C1362 out.t70 vss 0.00464f
C1363 out.n2 vss 0.0207f
C1364 out.n3 vss 0.0076f
C1365 out.n4 vss 0.00177f
C1366 out.n5 vss 0.0027f
C1367 out.n6 vss 0.00615f
C1368 out.t73 vss 0.00464f
C1369 out.t72 vss 0.00464f
C1370 out.n7 vss 0.0329f
C1371 out.t77 vss 0.00464f
C1372 out.t79 vss 0.00464f
C1373 out.n8 vss 0.0326f
C1374 out.t30 vss 0.00464f
C1375 out.t33 vss 0.00464f
C1376 out.n9 vss 0.0383f
C1377 out.t75 vss 0.00464f
C1378 out.t74 vss 0.00464f
C1379 out.n10 vss 0.0327f
C1380 out.t35 vss 0.00464f
C1381 out.t38 vss 0.00464f
C1382 out.n11 vss 0.0361f
C1383 out.n12 vss 0.0281f
C1384 out.t71 vss 0.00464f
C1385 out.t78 vss 0.00464f
C1386 out.n13 vss 0.0324f
C1387 out.n14 vss 0.0199f
C1388 out.t36 vss 0.00464f
C1389 out.t32 vss 0.00464f
C1390 out.n15 vss 0.0389f
C1391 out.n16 vss 0.0147f
C1392 out.n17 vss 0.0336f
C1393 out.t31 vss 0.00464f
C1394 out.t34 vss 0.00464f
C1395 out.n18 vss 0.0403f
C1396 out.n19 vss 0.0144f
C1397 out.n20 vss 0.0192f
C1398 out.t37 vss 0.00464f
C1399 out.t39 vss 0.00464f
C1400 out.n21 vss 0.04f
C1401 out.n22 vss 0.0138f
C1402 out.n23 vss 0.0152f
C1403 out.n24 vss 0.00165f
C1404 out.t48 vss 0.00464f
C1405 out.t49 vss 0.00464f
C1406 out.n26 vss 0.0207f
C1407 out.n27 vss 0.0076f
C1408 out.n28 vss 0.00177f
C1409 out.n29 vss 0.0027f
C1410 out.n30 vss 0.00615f
C1411 out.t43 vss 0.00464f
C1412 out.t44 vss 0.00464f
C1413 out.n31 vss 0.0329f
C1414 out.t47 vss 0.00464f
C1415 out.t41 vss 0.00464f
C1416 out.n32 vss 0.0326f
C1417 out.t12 vss 0.00464f
C1418 out.t18 vss 0.00464f
C1419 out.n33 vss 0.0383f
C1420 out.t45 vss 0.00464f
C1421 out.t40 vss 0.00464f
C1422 out.n34 vss 0.0327f
C1423 out.t16 vss 0.00464f
C1424 out.t15 vss 0.00464f
C1425 out.n35 vss 0.0361f
C1426 out.n36 vss 0.0281f
C1427 out.t42 vss 0.00464f
C1428 out.t46 vss 0.00464f
C1429 out.n37 vss 0.0324f
C1430 out.n38 vss 0.0199f
C1431 out.t10 vss 0.00464f
C1432 out.t13 vss 0.00464f
C1433 out.n39 vss 0.0389f
C1434 out.n40 vss 0.0147f
C1435 out.n41 vss 0.0336f
C1436 out.t14 vss 0.00464f
C1437 out.t19 vss 0.00464f
C1438 out.n42 vss 0.0403f
C1439 out.n43 vss 0.0144f
C1440 out.n44 vss 0.0192f
C1441 out.t17 vss 0.00464f
C1442 out.t11 vss 0.00464f
C1443 out.n45 vss 0.04f
C1444 out.n46 vss 0.0138f
C1445 out.n47 vss 0.0152f
C1446 out.n48 vss 0.00165f
C1447 out.t60 vss 0.00464f
C1448 out.t62 vss 0.00464f
C1449 out.n50 vss 0.0207f
C1450 out.n51 vss 0.0076f
C1451 out.n52 vss 0.00177f
C1452 out.n53 vss 0.0027f
C1453 out.n54 vss 0.00615f
C1454 out.t67 vss 0.00464f
C1455 out.t68 vss 0.00464f
C1456 out.n55 vss 0.0329f
C1457 out.t61 vss 0.00464f
C1458 out.t63 vss 0.00464f
C1459 out.n56 vss 0.0326f
C1460 out.t1 vss 0.00464f
C1461 out.t4 vss 0.00464f
C1462 out.n57 vss 0.0383f
C1463 out.t66 vss 0.00464f
C1464 out.t69 vss 0.00464f
C1465 out.n58 vss 0.0327f
C1466 out.t5 vss 0.00464f
C1467 out.t8 vss 0.00464f
C1468 out.n59 vss 0.0361f
C1469 out.n60 vss 0.0281f
C1470 out.t65 vss 0.00464f
C1471 out.t64 vss 0.00464f
C1472 out.n61 vss 0.0324f
C1473 out.n62 vss 0.0199f
C1474 out.t2 vss 0.00464f
C1475 out.t0 vss 0.00464f
C1476 out.n63 vss 0.0389f
C1477 out.n64 vss 0.0147f
C1478 out.n65 vss 0.0336f
C1479 out.t7 vss 0.00464f
C1480 out.t3 vss 0.00464f
C1481 out.n66 vss 0.0403f
C1482 out.n67 vss 0.0144f
C1483 out.n68 vss 0.0192f
C1484 out.t6 vss 0.00464f
C1485 out.t9 vss 0.00464f
C1486 out.n69 vss 0.04f
C1487 out.n70 vss 0.0138f
C1488 out.n71 vss 0.0152f
C1489 out.t218 vss 0.376f
C1490 out.t166 vss 0.256f
C1491 out.n72 vss 0.139f
C1492 out.t415 vss 0.256f
C1493 out.n73 vss 0.139f
C1494 out.t356 vss 0.256f
C1495 out.n74 vss 0.139f
C1496 out.t305 vss 0.256f
C1497 out.n75 vss 0.139f
C1498 out.t249 vss 0.256f
C1499 out.n76 vss 0.139f
C1500 out.t194 vss 0.256f
C1501 out.n77 vss 0.139f
C1502 out.t102 vss 0.256f
C1503 out.n78 vss 0.139f
C1504 out.t241 vss 0.256f
C1505 out.n79 vss 0.139f
C1506 out.t189 vss 0.256f
C1507 out.n80 vss 0.139f
C1508 out.t134 vss 0.256f
C1509 out.n81 vss 0.139f
C1510 out.t86 vss 0.256f
C1511 out.n82 vss 0.139f
C1512 out.t328 vss 0.256f
C1513 out.n83 vss 0.139f
C1514 out.t276 vss 0.256f
C1515 out.n84 vss 0.139f
C1516 out.t219 vss 0.256f
C1517 out.n85 vss 0.139f
C1518 out.t167 vss 0.256f
C1519 out.n86 vss 0.139f
C1520 out.t112 vss 0.256f
C1521 out.n87 vss 0.139f
C1522 out.t357 vss 0.256f
C1523 out.n88 vss 0.139f
C1524 out.t306 vss 0.256f
C1525 out.n89 vss 0.139f
C1526 out.t250 vss 0.256f
C1527 out.n90 vss 0.139f
C1528 out.t132 vss 0.256f
C1529 out.n91 vss 0.139f
C1530 out.t82 vss 0.256f
C1531 out.n92 vss 0.139f
C1532 out.t324 vss 0.256f
C1533 out.n93 vss 0.139f
C1534 out.t270 vss 0.256f
C1535 out.n94 vss 0.139f
C1536 out.t213 vss 0.256f
C1537 out.n95 vss 0.139f
C1538 out.t161 vss 0.256f
C1539 out.n96 vss 0.139f
C1540 out.t107 vss 0.256f
C1541 out.n97 vss 0.139f
C1542 out.t351 vss 0.256f
C1543 out.n98 vss 0.139f
C1544 out.t300 vss 0.256f
C1545 out.n99 vss 0.139f
C1546 out.t245 vss 0.256f
C1547 out.t191 vss 0.256f
C1548 out.t162 vss 0.256f
C1549 out.t192 vss 0.256f
C1550 out.n100 vss 0.108f
C1551 out.t264 vss 0.256f
C1552 out.t296 vss 0.376f
C1553 out.t238 vss 0.256f
C1554 out.n101 vss 0.139f
C1555 out.t141 vss 0.256f
C1556 out.n102 vss 0.139f
C1557 out.t90 vss 0.256f
C1558 out.n103 vss 0.139f
C1559 out.t378 vss 0.256f
C1560 out.n104 vss 0.139f
C1561 out.t322 vss 0.256f
C1562 out.n105 vss 0.139f
C1563 out.t269 vss 0.256f
C1564 out.n106 vss 0.139f
C1565 out.t175 vss 0.256f
C1566 out.n107 vss 0.139f
C1567 out.t317 vss 0.256f
C1568 out.n108 vss 0.139f
C1569 out.t261 vss 0.256f
C1570 out.n109 vss 0.139f
C1571 out.t207 vss 0.256f
C1572 out.n110 vss 0.139f
C1573 out.t152 vss 0.256f
C1574 out.n111 vss 0.139f
C1575 out.t407 vss 0.256f
C1576 out.n112 vss 0.139f
C1577 out.t345 vss 0.256f
C1578 out.n113 vss 0.139f
C1579 out.t297 vss 0.256f
C1580 out.n114 vss 0.139f
C1581 out.t239 vss 0.256f
C1582 out.n115 vss 0.139f
C1583 out.t186 vss 0.256f
C1584 out.n116 vss 0.139f
C1585 out.t91 vss 0.256f
C1586 out.n117 vss 0.139f
C1587 out.t379 vss 0.256f
C1588 out.n118 vss 0.139f
C1589 out.t323 vss 0.256f
C1590 out.n119 vss 0.139f
C1591 out.t201 vss 0.256f
C1592 out.n120 vss 0.139f
C1593 out.t147 vss 0.256f
C1594 out.n121 vss 0.139f
C1595 out.t401 vss 0.256f
C1596 out.n122 vss 0.139f
C1597 out.t338 vss 0.256f
C1598 out.n123 vss 0.139f
C1599 out.t292 vss 0.256f
C1600 out.n124 vss 0.139f
C1601 out.t232 vss 0.256f
C1602 out.n125 vss 0.139f
C1603 out.t180 vss 0.256f
C1604 out.n126 vss 0.139f
C1605 out.t87 vss 0.256f
C1606 out.n127 vss 0.139f
C1607 out.t374 vss 0.256f
C1608 out.n128 vss 0.139f
C1609 out.t319 vss 0.256f
C1610 out.n129 vss 0.139f
C1611 out.t263 vss 0.256f
C1612 out.n130 vss 0.139f
C1613 out.t235 vss 0.256f
C1614 out.n131 vss 0.139f
C1615 out.t155 vss 0.256f
C1616 out.t184 vss 0.376f
C1617 out.t130 vss 0.256f
C1618 out.n132 vss 0.139f
C1619 out.t377 vss 0.256f
C1620 out.n133 vss 0.139f
C1621 out.t320 vss 0.256f
C1622 out.n134 vss 0.139f
C1623 out.t267 vss 0.256f
C1624 out.n135 vss 0.139f
C1625 out.t211 vss 0.256f
C1626 out.n136 vss 0.139f
C1627 out.t160 vss 0.256f
C1628 out.n137 vss 0.139f
C1629 out.t411 vss 0.256f
C1630 out.n138 vss 0.139f
C1631 out.t205 vss 0.256f
C1632 out.n139 vss 0.139f
C1633 out.t150 vss 0.256f
C1634 out.n140 vss 0.139f
C1635 out.t100 vss 0.256f
C1636 out.n141 vss 0.139f
C1637 out.t391 vss 0.256f
C1638 out.n142 vss 0.139f
C1639 out.t295 vss 0.256f
C1640 out.n143 vss 0.139f
C1641 out.t237 vss 0.256f
C1642 out.n144 vss 0.139f
C1643 out.t185 vss 0.256f
C1644 out.n145 vss 0.139f
C1645 out.t131 vss 0.256f
C1646 out.n146 vss 0.139f
C1647 out.t81 vss 0.256f
C1648 out.n147 vss 0.139f
C1649 out.t321 vss 0.256f
C1650 out.n148 vss 0.139f
C1651 out.t268 vss 0.256f
C1652 out.n149 vss 0.139f
C1653 out.t212 vss 0.256f
C1654 out.n150 vss 0.139f
C1655 out.t95 vss 0.256f
C1656 out.n151 vss 0.139f
C1657 out.t385 vss 0.256f
C1658 out.n152 vss 0.139f
C1659 out.t290 vss 0.256f
C1660 out.n153 vss 0.139f
C1661 out.t231 vss 0.256f
C1662 out.n154 vss 0.139f
C1663 out.t179 vss 0.256f
C1664 out.n155 vss 0.139f
C1665 out.t122 vss 0.256f
C1666 out.n156 vss 0.139f
C1667 out.t414 vss 0.256f
C1668 out.n157 vss 0.139f
C1669 out.t318 vss 0.256f
C1670 out.n158 vss 0.139f
C1671 out.t262 vss 0.256f
C1672 out.n159 vss 0.139f
C1673 out.t206 vss 0.256f
C1674 out.n160 vss 0.139f
C1675 out.t153 vss 0.256f
C1676 out.n161 vss 0.139f
C1677 out.t123 vss 0.256f
C1678 out.n162 vss 0.139f
C1679 out.t395 vss 0.256f
C1680 out.t417 vss 0.376f
C1681 out.t362 vss 0.256f
C1682 out.n163 vss 0.139f
C1683 out.t266 vss 0.256f
C1684 out.n164 vss 0.139f
C1685 out.t209 vss 0.256f
C1686 out.n165 vss 0.139f
C1687 out.t156 vss 0.256f
C1688 out.n166 vss 0.139f
C1689 out.t104 vss 0.256f
C1690 out.n167 vss 0.139f
C1691 out.t398 vss 0.256f
C1692 out.n168 vss 0.139f
C1693 out.t298 vss 0.256f
C1694 out.n169 vss 0.139f
C1695 out.t99 vss 0.256f
C1696 out.n170 vss 0.139f
C1697 out.t389 vss 0.256f
C1698 out.n171 vss 0.139f
C1699 out.t331 vss 0.256f
C1700 out.n172 vss 0.139f
C1701 out.t279 vss 0.256f
C1702 out.n173 vss 0.139f
C1703 out.t183 vss 0.256f
C1704 out.n174 vss 0.139f
C1705 out.t128 vss 0.256f
C1706 out.n175 vss 0.139f
C1707 out.t80 vss 0.256f
C1708 out.n176 vss 0.139f
C1709 out.t363 vss 0.256f
C1710 out.n177 vss 0.139f
C1711 out.t309 vss 0.256f
C1712 out.n178 vss 0.139f
C1713 out.t210 vss 0.256f
C1714 out.n179 vss 0.139f
C1715 out.t157 vss 0.256f
C1716 out.n180 vss 0.139f
C1717 out.t106 vss 0.256f
C1718 out.n181 vss 0.139f
C1719 out.t327 vss 0.256f
C1720 out.n182 vss 0.139f
C1721 out.t272 vss 0.256f
C1722 out.n183 vss 0.139f
C1723 out.t178 vss 0.256f
C1724 out.n184 vss 0.139f
C1725 out.t121 vss 0.256f
C1726 out.n185 vss 0.139f
C1727 out.t413 vss 0.256f
C1728 out.n186 vss 0.139f
C1729 out.t353 vss 0.256f
C1730 out.n187 vss 0.139f
C1731 out.t303 vss 0.256f
C1732 out.n188 vss 0.139f
C1733 out.t204 vss 0.256f
C1734 out.n189 vss 0.139f
C1735 out.t151 vss 0.256f
C1736 out.n190 vss 0.139f
C1737 out.t101 vss 0.256f
C1738 out.n191 vss 0.139f
C1739 out.t390 vss 0.256f
C1740 out.n192 vss 0.139f
C1741 out.t355 vss 0.256f
C1742 out.n193 vss 0.139f
C1743 out.t118 vss 0.256f
C1744 out.t145 vss 0.376f
C1745 out.t94 vss 0.256f
C1746 out.n194 vss 0.139f
C1747 out.t336 vss 0.256f
C1748 out.n195 vss 0.139f
C1749 out.t289 vss 0.256f
C1750 out.n196 vss 0.139f
C1751 out.t229 vss 0.256f
C1752 out.n197 vss 0.139f
C1753 out.t176 vss 0.256f
C1754 out.n198 vss 0.139f
C1755 out.t120 vss 0.256f
C1756 out.n199 vss 0.139f
C1757 out.t373 vss 0.256f
C1758 out.n200 vss 0.139f
C1759 out.t170 vss 0.256f
C1760 out.n201 vss 0.139f
C1761 out.t114 vss 0.256f
C1762 out.n202 vss 0.139f
C1763 out.t409 vss 0.256f
C1764 out.n203 vss 0.139f
C1765 out.t346 vss 0.256f
C1766 out.n204 vss 0.139f
C1767 out.t255 vss 0.256f
C1768 out.n205 vss 0.139f
C1769 out.t200 vss 0.256f
C1770 out.n206 vss 0.139f
C1771 out.t144 vss 0.256f
C1772 out.n207 vss 0.139f
C1773 out.t93 vss 0.256f
C1774 out.n208 vss 0.139f
C1775 out.t382 vss 0.256f
C1776 out.n209 vss 0.139f
C1777 out.t288 vss 0.256f
C1778 out.n210 vss 0.139f
C1779 out.t230 vss 0.256f
C1780 out.n211 vss 0.139f
C1781 out.t177 vss 0.256f
C1782 out.n212 vss 0.139f
C1783 out.t406 vss 0.256f
C1784 out.n213 vss 0.139f
C1785 out.t342 vss 0.256f
C1786 out.n214 vss 0.139f
C1787 out.t248 vss 0.256f
C1788 out.n215 vss 0.139f
C1789 out.t193 vss 0.256f
C1790 out.n216 vss 0.139f
C1791 out.t139 vss 0.256f
C1792 out.n217 vss 0.139f
C1793 out.t88 vss 0.256f
C1794 out.n218 vss 0.139f
C1795 out.t375 vss 0.256f
C1796 out.n219 vss 0.139f
C1797 out.t284 vss 0.256f
C1798 out.n220 vss 0.139f
C1799 out.t222 vss 0.256f
C1800 out.n221 vss 0.139f
C1801 out.t171 vss 0.256f
C1802 out.n222 vss 0.139f
C1803 out.t117 vss 0.256f
C1804 out.n223 vss 0.139f
C1805 out.t89 vss 0.256f
C1806 out.n224 vss 0.139f
C1807 out.t253 vss 0.256f
C1808 out.t227 vss 0.376f
C1809 out.t97 vss 0.256f
C1810 out.n225 vss 0.139f
C1811 out.t83 vss 0.256f
C1812 out.n226 vss 0.139f
C1813 out.t287 vss 0.256f
C1814 out.n227 vss 0.139f
C1815 out.t149 vss 0.256f
C1816 out.n228 vss 0.139f
C1817 out.t350 vss 0.256f
C1818 out.n229 vss 0.139f
C1819 out.t217 vss 0.256f
C1820 out.n230 vss 0.139f
C1821 out.t198 vss 0.256f
C1822 out.n231 vss 0.139f
C1823 out.t103 vss 0.256f
C1824 out.n232 vss 0.139f
C1825 out.t312 vss 0.256f
C1826 out.n233 vss 0.139f
C1827 out.t174 vss 0.256f
C1828 out.n234 vss 0.139f
C1829 out.t386 vss 0.256f
C1830 out.n235 vss 0.139f
C1831 out.t364 vss 0.256f
C1832 out.n236 vss 0.139f
C1833 out.t226 vss 0.256f
C1834 out.n237 vss 0.139f
C1835 out.t96 vss 0.256f
C1836 out.n238 vss 0.139f
C1837 out.t301 vss 0.256f
C1838 out.n239 vss 0.139f
C1839 out.t165 vss 0.256f
C1840 out.n240 vss 0.139f
C1841 out.t142 vss 0.256f
C1842 out.n241 vss 0.139f
C1843 out.t347 vss 0.256f
C1844 out.n242 vss 0.139f
C1845 out.t215 vss 0.256f
C1846 out.n243 vss 0.139f
C1847 out.t146 vss 0.256f
C1848 out.n244 vss 0.139f
C1849 out.t349 vss 0.256f
C1850 out.n245 vss 0.139f
C1851 out.t332 vss 0.256f
C1852 out.n246 vss 0.139f
C1853 out.t197 vss 0.256f
C1854 out.n247 vss 0.139f
C1855 out.t410 vss 0.256f
C1856 out.n248 vss 0.139f
C1857 out.t273 vss 0.256f
C1858 out.n249 vss 0.139f
C1859 out.t136 vss 0.256f
C1860 out.n250 vss 0.139f
C1861 out.t116 vss 0.256f
C1862 out.n251 vss 0.139f
C1863 out.t325 vss 0.256f
C1864 out.n252 vss 0.139f
C1865 out.t188 vss 0.256f
C1866 out.n253 vss 0.139f
C1867 out.t400 vss 0.256f
C1868 out.n254 vss 0.139f
C1869 out.t392 vss 0.256f
C1870 out.n255 vss 0.139f
C1871 out.t84 vss 0.256f
C1872 out.t367 vss 0.256f
C1873 out.t315 vss 0.256f
C1874 out.t216 vss 0.256f
C1875 out.t163 vss 0.256f
C1876 out.t109 vss 0.256f
C1877 out.t404 vss 0.256f
C1878 out.t341 vss 0.256f
C1879 out.t247 vss 0.256f
C1880 out.t397 vss 0.256f
C1881 out.t333 vss 0.256f
C1882 out.t285 vss 0.256f
C1883 out.t225 vss 0.256f
C1884 out.t133 vss 0.256f
C1885 out.t85 vss 0.256f
C1886 out.t370 vss 0.256f
C1887 out.t316 vss 0.256f
C1888 out.t259 vss 0.256f
C1889 out.t164 vss 0.256f
C1890 out.t110 vss 0.256f
C1891 out.t405 vss 0.256f
C1892 out.t280 vss 0.256f
C1893 out.t221 vss 0.256f
C1894 out.t129 vss 0.256f
C1895 out.t419 vss 0.256f
C1896 out.t361 vss 0.256f
C1897 out.t310 vss 0.256f
C1898 out.t252 vss 0.256f
C1899 out.t158 vss 0.256f
C1900 out.t105 vss 0.256f
C1901 out.t399 vss 0.256f
C1902 out.t335 vss 0.256f
C1903 out.t311 vss 0.256f
C1904 out.t337 vss 0.256f
C1905 out.t228 vss 0.256f
C1906 out.t256 vss 0.376f
C1907 out.t202 vss 0.256f
C1908 out.n256 vss 0.139f
C1909 out.t108 vss 0.256f
C1910 out.n257 vss 0.139f
C1911 out.t402 vss 0.256f
C1912 out.n258 vss 0.139f
C1913 out.t339 vss 0.256f
C1914 out.n259 vss 0.139f
C1915 out.t291 vss 0.256f
C1916 out.n260 vss 0.139f
C1917 out.t233 vss 0.256f
C1918 out.n261 vss 0.139f
C1919 out.t138 vss 0.256f
C1920 out.n262 vss 0.139f
C1921 out.t282 vss 0.256f
C1922 out.n263 vss 0.139f
C1923 out.t223 vss 0.256f
C1924 out.n264 vss 0.139f
C1925 out.t172 vss 0.256f
C1926 out.n265 vss 0.139f
C1927 out.t115 vss 0.256f
C1928 out.n266 vss 0.139f
C1929 out.t366 vss 0.256f
C1930 out.n267 vss 0.139f
C1931 out.t314 vss 0.256f
C1932 out.n268 vss 0.139f
C1933 out.t257 vss 0.256f
C1934 out.n269 vss 0.139f
C1935 out.t203 vss 0.256f
C1936 out.n270 vss 0.139f
C1937 out.t148 vss 0.256f
C1938 out.n271 vss 0.139f
C1939 out.t403 vss 0.256f
C1940 out.n272 vss 0.139f
C1941 out.t340 vss 0.256f
C1942 out.n273 vss 0.139f
C1943 out.t293 vss 0.256f
C1944 out.n274 vss 0.139f
C1945 out.t168 vss 0.256f
C1946 out.n275 vss 0.139f
C1947 out.t113 vss 0.256f
C1948 out.n276 vss 0.139f
C1949 out.t360 vss 0.256f
C1950 out.n277 vss 0.139f
C1951 out.t308 vss 0.256f
C1952 out.n278 vss 0.139f
C1953 out.t251 vss 0.256f
C1954 out.n279 vss 0.139f
C1955 out.t195 vss 0.256f
C1956 out.n280 vss 0.139f
C1957 out.t140 vss 0.256f
C1958 out.n281 vss 0.139f
C1959 out.t396 vss 0.256f
C1960 out.n282 vss 0.139f
C1961 out.t334 vss 0.256f
C1962 out.n283 vss 0.139f
C1963 out.t286 vss 0.256f
C1964 out.n284 vss 0.139f
C1965 out.t224 vss 0.256f
C1966 out.n285 vss 0.139f
C1967 out.t196 vss 0.256f
C1968 out.n286 vss 0.139f
C1969 out.t304 vss 0.256f
C1970 out.t329 vss 0.376f
C1971 out.t277 vss 0.256f
C1972 out.n287 vss 0.139f
C1973 out.t182 vss 0.256f
C1974 out.n288 vss 0.139f
C1975 out.t125 vss 0.256f
C1976 out.n289 vss 0.139f
C1977 out.t416 vss 0.256f
C1978 out.n290 vss 0.139f
C1979 out.t358 vss 0.256f
C1980 out.n291 vss 0.139f
C1981 out.t307 vss 0.256f
C1982 out.n292 vss 0.139f
C1983 out.t208 vss 0.256f
C1984 out.n293 vss 0.139f
C1985 out.t348 vss 0.256f
C1986 out.n294 vss 0.139f
C1987 out.t299 vss 0.256f
C1988 out.n295 vss 0.139f
C1989 out.t242 vss 0.256f
C1990 out.n296 vss 0.139f
C1991 out.t190 vss 0.256f
C1992 out.n297 vss 0.139f
C1993 out.t98 vss 0.256f
C1994 out.n298 vss 0.139f
C1995 out.t388 vss 0.256f
C1996 out.n299 vss 0.139f
C1997 out.t330 vss 0.256f
C1998 out.n300 vss 0.139f
C1999 out.t278 vss 0.256f
C2000 out.n301 vss 0.139f
C2001 out.t220 vss 0.256f
C2002 out.n302 vss 0.139f
C2003 out.t126 vss 0.256f
C2004 out.n303 vss 0.139f
C2005 out.t418 vss 0.256f
C2006 out.n304 vss 0.139f
C2007 out.t359 vss 0.256f
C2008 out.n305 vss 0.139f
C2009 out.t240 vss 0.256f
C2010 out.n306 vss 0.139f
C2011 out.t187 vss 0.256f
C2012 out.n307 vss 0.139f
C2013 out.t92 vss 0.256f
C2014 out.n308 vss 0.139f
C2015 out.t380 vss 0.256f
C2016 out.n309 vss 0.139f
C2017 out.t326 vss 0.256f
C2018 out.n310 vss 0.139f
C2019 out.t271 vss 0.256f
C2020 out.n311 vss 0.139f
C2021 out.t214 vss 0.256f
C2022 out.n312 vss 0.139f
C2023 out.t119 vss 0.256f
C2024 out.n313 vss 0.139f
C2025 out.t412 vss 0.256f
C2026 out.n314 vss 0.139f
C2027 out.t352 vss 0.256f
C2028 out.n315 vss 0.139f
C2029 out.t302 vss 0.256f
C2030 out.n316 vss 0.139f
C2031 out.t274 vss 0.256f
C2032 out.n317 vss 0.139f
C2033 out.n318 vss 0.05f
C2034 out.n319 vss 0.116f
C2035 out.n320 vss 0.05f
C2036 out.n321 vss 0.111f
C2037 out.n322 vss 0.0558f
C2038 out.n323 vss 0.106f
C2039 out.n324 vss 0.139f
C2040 out.n325 vss 0.139f
C2041 out.n326 vss 0.139f
C2042 out.n327 vss 0.139f
C2043 out.n328 vss 0.139f
C2044 out.n329 vss 0.139f
C2045 out.n330 vss 0.139f
C2046 out.n331 vss 0.139f
C2047 out.n332 vss 0.139f
C2048 out.n333 vss 0.139f
C2049 out.n334 vss 0.139f
C2050 out.n335 vss 0.139f
C2051 out.n336 vss 0.139f
C2052 out.n337 vss 0.139f
C2053 out.n338 vss 0.139f
C2054 out.n339 vss 0.139f
C2055 out.n340 vss 0.139f
C2056 out.n341 vss 0.139f
C2057 out.n342 vss 0.139f
C2058 out.n343 vss 0.139f
C2059 out.n344 vss 0.139f
C2060 out.n345 vss 0.139f
C2061 out.n346 vss 0.139f
C2062 out.n347 vss 0.139f
C2063 out.n348 vss 0.139f
C2064 out.n349 vss 0.139f
C2065 out.n350 vss 0.139f
C2066 out.n351 vss 0.139f
C2067 out.n352 vss 0.139f
C2068 out.n353 vss 0.139f
C2069 out.n354 vss 0.139f
C2070 out.n355 vss 0.139f
C2071 out.n356 vss 0.138f
C2072 out.t313 vss 0.256f
C2073 out.n357 vss 0.118f
C2074 out.t387 vss 0.256f
C2075 out.n358 vss 0.119f
C2076 out.t275 vss 0.256f
C2077 out.n359 vss 0.119f
C2078 out.t344 vss 0.256f
C2079 out.n360 vss 0.119f
C2080 out.t236 vss 0.256f
C2081 out.n361 vss 0.119f
C2082 out.t127 vss 0.256f
C2083 out.n362 vss 0.119f
C2084 out.t199 vss 0.256f
C2085 out.n363 vss 0.119f
C2086 out.t365 vss 0.256f
C2087 out.n364 vss 0.119f
C2088 out.t294 vss 0.256f
C2089 out.n365 vss 0.0932f
C2090 out.n366 vss 0.0536f
C2091 out.t169 vss 0.256f
C2092 out.n367 vss 0.139f
C2093 out.t394 vss 0.256f
C2094 out.n368 vss 0.139f
C2095 out.t181 vss 0.256f
C2096 out.n369 vss 0.139f
C2097 out.t408 vss 0.256f
C2098 out.n370 vss 0.139f
C2099 out.t283 vss 0.256f
C2100 out.n371 vss 0.139f
C2101 out.t159 vss 0.256f
C2102 out.n372 vss 0.139f
C2103 out.t384 vss 0.256f
C2104 out.n373 vss 0.139f
C2105 out.t173 vss 0.256f
C2106 out.n374 vss 0.139f
C2107 out.t281 vss 0.256f
C2108 out.n375 vss 0.139f
C2109 out.t154 vss 0.256f
C2110 out.n376 vss 0.139f
C2111 out.t376 vss 0.256f
C2112 out.n377 vss 0.139f
C2113 out.t254 vss 0.256f
C2114 out.n378 vss 0.139f
C2115 out.t393 vss 0.256f
C2116 out.n379 vss 0.139f
C2117 out.t265 vss 0.256f
C2118 out.n380 vss 0.139f
C2119 out.t143 vss 0.256f
C2120 out.n381 vss 0.139f
C2121 out.t369 vss 0.256f
C2122 out.n382 vss 0.139f
C2123 out.t244 vss 0.256f
C2124 out.n383 vss 0.139f
C2125 out.t383 vss 0.256f
C2126 out.n384 vss 0.139f
C2127 out.t260 vss 0.256f
C2128 out.n385 vss 0.139f
C2129 out.t137 vss 0.256f
C2130 out.n386 vss 0.139f
C2131 out.t368 vss 0.256f
C2132 out.n387 vss 0.139f
C2133 out.t243 vss 0.256f
C2134 out.n388 vss 0.139f
C2135 out.t381 vss 0.256f
C2136 out.n389 vss 0.139f
C2137 out.t258 vss 0.256f
C2138 out.n390 vss 0.139f
C2139 out.t135 vss 0.256f
C2140 out.n391 vss 0.139f
C2141 out.t354 vss 0.256f
C2142 out.n392 vss 0.139f
C2143 out.t234 vss 0.256f
C2144 out.n393 vss 0.139f
C2145 out.t372 vss 0.256f
C2146 out.n394 vss 0.139f
C2147 out.t246 vss 0.256f
C2148 out.n395 vss 0.139f
C2149 out.t124 vss 0.256f
C2150 out.n396 vss 0.139f
C2151 out.t343 vss 0.256f
C2152 out.n397 vss 0.139f
C2153 out.t111 vss 0.256f
C2154 out.n398 vss 0.139f
C2155 out.t371 vss 0.256f
C2156 out.n399 vss 0.106f
C2157 out.n400 vss 0.0515f
C2158 out.n401 vss 0.05f
C2159 out.n402 vss 0.111f
C2160 out.n403 vss 0.05f
C2161 out.n404 vss 0.111f
C2162 out.n405 vss 0.05f
C2163 out.n406 vss 0.108f
C2164 out.n407 vss 0.05f
C2165 out.n408 vss 0.113f
C2166 out.n409 vss 0.05f
C2167 out.n410 vss 0.113f
C2168 out.n411 vss 0.05f
C2169 out.n412 vss 0.139f
C2170 out.n413 vss 0.139f
C2171 out.n414 vss 0.126f
C2172 out.n415 vss 0.0633f
C2173 out.n416 vss 0.00165f
C2174 out.t55 vss 0.00464f
C2175 out.t54 vss 0.00464f
C2176 out.n418 vss 0.0207f
C2177 out.n419 vss 0.0076f
C2178 out.n420 vss 0.00177f
C2179 out.n421 vss 0.0027f
C2180 out.n422 vss 0.00615f
C2181 out.t53 vss 0.00464f
C2182 out.t50 vss 0.00464f
C2183 out.n423 vss 0.0329f
C2184 out.t51 vss 0.00464f
C2185 out.t59 vss 0.00464f
C2186 out.n424 vss 0.0326f
C2187 out.t28 vss 0.00464f
C2188 out.t24 vss 0.00464f
C2189 out.n425 vss 0.0383f
C2190 out.t52 vss 0.00464f
C2191 out.t57 vss 0.00464f
C2192 out.n426 vss 0.0327f
C2193 out.t25 vss 0.00464f
C2194 out.t23 vss 0.00464f
C2195 out.n427 vss 0.0361f
C2196 out.n428 vss 0.0281f
C2197 out.t56 vss 0.00464f
C2198 out.t58 vss 0.00464f
C2199 out.n429 vss 0.0324f
C2200 out.n430 vss 0.0199f
C2201 out.t22 vss 0.00464f
C2202 out.t21 vss 0.00464f
C2203 out.n431 vss 0.0389f
C2204 out.n432 vss 0.0147f
C2205 out.n433 vss 0.0336f
C2206 out.t29 vss 0.00464f
C2207 out.t27 vss 0.00464f
C2208 out.n434 vss 0.0403f
C2209 out.n435 vss 0.0144f
C2210 out.n436 vss 0.0192f
C2211 out.t26 vss 0.00464f
C2212 out.t20 vss 0.00464f
C2213 out.n437 vss 0.04f
C2214 out.n438 vss 0.0138f
C2215 out.n439 vss 0.0152f
C2216 out.n440 vss 0.0413f
C2217 out.n441 vss 0.0687f
C2218 out.n442 vss 0.12f
C2219 out.n443 vss 0.159f
C2220 out.n444 vss 0.0824f
.ends

