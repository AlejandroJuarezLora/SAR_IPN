magic
tech sky130B
magscale 1 2
timestamp 1696029713
<< metal1 >>
rect 1769 1271 4811 1301
rect 1749 521 4849 551
use nfet_4mimcap_combo  nfet_4mimcap_combo_1
timestamp 1696029615
transform 1 0 0 0 1 0
box 0 0 2196 1334
use trimcap  trimcap_0
timestamp 1695926252
transform 1 0 4574 0 1 58
box 0 426 476 1274
use trimcap  trimcap_1
timestamp 1695926252
transform 1 0 2294 0 1 58
box 0 426 476 1274
use trimcap  trimcap_2
timestamp 1695926252
transform 1 0 2864 0 1 58
box 0 426 476 1274
use trimcap  trimcap_3
timestamp 1695926252
transform 1 0 3432 0 1 58
box 0 426 476 1274
use trimcap  trimcap_4
timestamp 1695926252
transform 1 0 4000 0 1 58
box 0 426 476 1274
<< end >>
