magic
tech sky130B
magscale 1 2
timestamp 1697130564
<< nwell >>
rect 0 657 2306 1331
<< pwell >>
rect 10 527 2296 613
rect 10 45 96 527
rect 165 189 413 441
rect 479 189 727 441
rect 793 189 1041 441
rect 1265 189 1513 441
rect 1579 189 1827 441
rect 1893 189 2141 441
rect 2210 45 2296 527
rect 10 -41 2296 45
<< pmoslvt >>
rect 249 900 329 1100
rect 877 900 957 1100
rect 1349 900 1429 1100
rect 1977 900 2057 1100
<< nmoslvt >>
rect 249 215 329 415
rect 563 215 643 415
rect 877 215 957 415
rect 1349 215 1429 415
rect 1663 215 1743 415
rect 1977 215 2057 415
<< ndiff >>
rect 191 400 249 415
rect 191 366 203 400
rect 237 366 249 400
rect 191 332 249 366
rect 191 298 203 332
rect 237 298 249 332
rect 191 264 249 298
rect 191 230 203 264
rect 237 230 249 264
rect 191 215 249 230
rect 329 400 387 415
rect 329 366 341 400
rect 375 366 387 400
rect 329 332 387 366
rect 329 298 341 332
rect 375 298 387 332
rect 329 264 387 298
rect 329 230 341 264
rect 375 230 387 264
rect 329 215 387 230
rect 505 400 563 415
rect 505 366 517 400
rect 551 366 563 400
rect 505 332 563 366
rect 505 298 517 332
rect 551 298 563 332
rect 505 264 563 298
rect 505 230 517 264
rect 551 230 563 264
rect 505 215 563 230
rect 643 400 701 415
rect 643 366 655 400
rect 689 366 701 400
rect 643 332 701 366
rect 643 298 655 332
rect 689 298 701 332
rect 643 264 701 298
rect 643 230 655 264
rect 689 230 701 264
rect 643 215 701 230
rect 819 400 877 415
rect 819 366 831 400
rect 865 366 877 400
rect 819 332 877 366
rect 819 298 831 332
rect 865 298 877 332
rect 819 264 877 298
rect 819 230 831 264
rect 865 230 877 264
rect 819 215 877 230
rect 957 400 1015 415
rect 957 366 969 400
rect 1003 366 1015 400
rect 957 332 1015 366
rect 957 298 969 332
rect 1003 298 1015 332
rect 957 264 1015 298
rect 957 230 969 264
rect 1003 230 1015 264
rect 957 215 1015 230
rect 1291 400 1349 415
rect 1291 366 1303 400
rect 1337 366 1349 400
rect 1291 332 1349 366
rect 1291 298 1303 332
rect 1337 298 1349 332
rect 1291 264 1349 298
rect 1291 230 1303 264
rect 1337 230 1349 264
rect 1291 215 1349 230
rect 1429 400 1487 415
rect 1429 366 1441 400
rect 1475 366 1487 400
rect 1429 332 1487 366
rect 1429 298 1441 332
rect 1475 298 1487 332
rect 1429 264 1487 298
rect 1429 230 1441 264
rect 1475 230 1487 264
rect 1429 215 1487 230
rect 1605 400 1663 415
rect 1605 366 1617 400
rect 1651 366 1663 400
rect 1605 332 1663 366
rect 1605 298 1617 332
rect 1651 298 1663 332
rect 1605 264 1663 298
rect 1605 230 1617 264
rect 1651 230 1663 264
rect 1605 215 1663 230
rect 1743 400 1801 415
rect 1743 366 1755 400
rect 1789 366 1801 400
rect 1743 332 1801 366
rect 1743 298 1755 332
rect 1789 298 1801 332
rect 1743 264 1801 298
rect 1743 230 1755 264
rect 1789 230 1801 264
rect 1743 215 1801 230
rect 1919 400 1977 415
rect 1919 366 1931 400
rect 1965 366 1977 400
rect 1919 332 1977 366
rect 1919 298 1931 332
rect 1965 298 1977 332
rect 1919 264 1977 298
rect 1919 230 1931 264
rect 1965 230 1977 264
rect 1919 215 1977 230
rect 2057 400 2115 415
rect 2057 366 2069 400
rect 2103 366 2115 400
rect 2057 332 2115 366
rect 2057 298 2069 332
rect 2103 298 2115 332
rect 2057 264 2115 298
rect 2057 230 2069 264
rect 2103 230 2115 264
rect 2057 215 2115 230
<< pdiff >>
rect 191 1085 249 1100
rect 191 1051 203 1085
rect 237 1051 249 1085
rect 191 1017 249 1051
rect 191 983 203 1017
rect 237 983 249 1017
rect 191 949 249 983
rect 191 915 203 949
rect 237 915 249 949
rect 191 900 249 915
rect 329 1085 387 1100
rect 329 1051 341 1085
rect 375 1051 387 1085
rect 329 1017 387 1051
rect 329 983 341 1017
rect 375 983 387 1017
rect 329 949 387 983
rect 329 915 341 949
rect 375 915 387 949
rect 329 900 387 915
rect 819 1085 877 1100
rect 819 1051 831 1085
rect 865 1051 877 1085
rect 819 1017 877 1051
rect 819 983 831 1017
rect 865 983 877 1017
rect 819 949 877 983
rect 819 915 831 949
rect 865 915 877 949
rect 819 900 877 915
rect 957 1085 1015 1100
rect 957 1051 969 1085
rect 1003 1051 1015 1085
rect 957 1017 1015 1051
rect 957 983 969 1017
rect 1003 983 1015 1017
rect 957 949 1015 983
rect 957 915 969 949
rect 1003 915 1015 949
rect 957 900 1015 915
rect 1291 1085 1349 1100
rect 1291 1051 1303 1085
rect 1337 1051 1349 1085
rect 1291 1017 1349 1051
rect 1291 983 1303 1017
rect 1337 983 1349 1017
rect 1291 949 1349 983
rect 1291 915 1303 949
rect 1337 915 1349 949
rect 1291 900 1349 915
rect 1429 1085 1487 1100
rect 1429 1051 1441 1085
rect 1475 1051 1487 1085
rect 1429 1017 1487 1051
rect 1429 983 1441 1017
rect 1475 983 1487 1017
rect 1429 949 1487 983
rect 1429 915 1441 949
rect 1475 915 1487 949
rect 1429 900 1487 915
rect 1919 1085 1977 1100
rect 1919 1051 1931 1085
rect 1965 1051 1977 1085
rect 1919 1017 1977 1051
rect 1919 983 1931 1017
rect 1965 983 1977 1017
rect 1919 949 1977 983
rect 1919 915 1931 949
rect 1965 915 1977 949
rect 1919 900 1977 915
rect 2057 1085 2115 1100
rect 2057 1051 2069 1085
rect 2103 1051 2115 1085
rect 2057 1017 2115 1051
rect 2057 983 2069 1017
rect 2103 983 2115 1017
rect 2057 949 2115 983
rect 2057 915 2069 949
rect 2103 915 2115 949
rect 2057 900 2115 915
<< ndiffc >>
rect 203 366 237 400
rect 203 298 237 332
rect 203 230 237 264
rect 341 366 375 400
rect 341 298 375 332
rect 341 230 375 264
rect 517 366 551 400
rect 517 298 551 332
rect 517 230 551 264
rect 655 366 689 400
rect 655 298 689 332
rect 655 230 689 264
rect 831 366 865 400
rect 831 298 865 332
rect 831 230 865 264
rect 969 366 1003 400
rect 969 298 1003 332
rect 969 230 1003 264
rect 1303 366 1337 400
rect 1303 298 1337 332
rect 1303 230 1337 264
rect 1441 366 1475 400
rect 1441 298 1475 332
rect 1441 230 1475 264
rect 1617 366 1651 400
rect 1617 298 1651 332
rect 1617 230 1651 264
rect 1755 366 1789 400
rect 1755 298 1789 332
rect 1755 230 1789 264
rect 1931 366 1965 400
rect 1931 298 1965 332
rect 1931 230 1965 264
rect 2069 366 2103 400
rect 2069 298 2103 332
rect 2069 230 2103 264
<< pdiffc >>
rect 203 1051 237 1085
rect 203 983 237 1017
rect 203 915 237 949
rect 341 1051 375 1085
rect 341 983 375 1017
rect 341 915 375 949
rect 831 1051 865 1085
rect 831 983 865 1017
rect 831 915 865 949
rect 969 1051 1003 1085
rect 969 983 1003 1017
rect 969 915 1003 949
rect 1303 1051 1337 1085
rect 1303 983 1337 1017
rect 1303 915 1337 949
rect 1441 1051 1475 1085
rect 1441 983 1475 1017
rect 1441 915 1475 949
rect 1931 1051 1965 1085
rect 1931 983 1965 1017
rect 1931 915 1965 949
rect 2069 1051 2103 1085
rect 2069 983 2103 1017
rect 2069 915 2103 949
<< psubdiff >>
rect 36 553 200 587
rect 234 553 268 587
rect 302 553 336 587
rect 370 553 404 587
rect 438 553 472 587
rect 506 553 540 587
rect 574 553 608 587
rect 642 553 676 587
rect 710 553 744 587
rect 778 553 812 587
rect 846 553 880 587
rect 914 553 948 587
rect 982 553 1016 587
rect 1050 553 1084 587
rect 1118 553 1152 587
rect 1186 553 1220 587
rect 1254 553 1288 587
rect 1322 553 1356 587
rect 1390 553 1424 587
rect 1458 553 1492 587
rect 1526 553 1560 587
rect 1594 553 1628 587
rect 1662 553 1696 587
rect 1730 553 1764 587
rect 1798 553 1832 587
rect 1866 553 1900 587
rect 1934 553 1968 587
rect 2002 553 2036 587
rect 2070 553 2270 587
rect 36 355 70 553
rect 36 287 70 321
rect 36 219 70 253
rect 2236 355 2270 553
rect 2236 287 2270 321
rect 2236 219 2270 253
rect 36 19 70 185
rect 2236 19 2270 185
rect 36 -15 268 19
rect 302 -15 336 19
rect 370 -15 404 19
rect 438 -15 472 19
rect 506 -15 540 19
rect 574 -15 608 19
rect 642 -15 676 19
rect 710 -15 744 19
rect 778 -15 812 19
rect 846 -15 880 19
rect 914 -15 948 19
rect 982 -15 1016 19
rect 1050 -15 1084 19
rect 1118 -15 1152 19
rect 1186 -15 1220 19
rect 1254 -15 1288 19
rect 1322 -15 1356 19
rect 1390 -15 1424 19
rect 1458 -15 1492 19
rect 1526 -15 1560 19
rect 1594 -15 1628 19
rect 1662 -15 1696 19
rect 1730 -15 1764 19
rect 1798 -15 1832 19
rect 1866 -15 1900 19
rect 1934 -15 1968 19
rect 2002 -15 2036 19
rect 2070 -15 2270 19
<< nsubdiff >>
rect 36 1261 124 1295
rect 158 1261 192 1295
rect 226 1261 260 1295
rect 294 1261 328 1295
rect 362 1261 396 1295
rect 430 1261 464 1295
rect 498 1261 532 1295
rect 566 1261 600 1295
rect 634 1261 668 1295
rect 702 1261 736 1295
rect 770 1261 804 1295
rect 838 1261 872 1295
rect 906 1261 940 1295
rect 974 1261 1008 1295
rect 1042 1261 1076 1295
rect 1110 1261 1144 1295
rect 1178 1261 1212 1295
rect 1246 1261 1280 1295
rect 1314 1261 1348 1295
rect 1382 1261 1416 1295
rect 1450 1261 1484 1295
rect 1518 1261 1552 1295
rect 1586 1261 1620 1295
rect 1654 1261 1688 1295
rect 1722 1261 1756 1295
rect 1790 1261 1824 1295
rect 1858 1261 1892 1295
rect 1926 1261 1960 1295
rect 1994 1261 2028 1295
rect 2062 1261 2096 1295
rect 2130 1261 2270 1295
rect 36 1155 70 1261
rect 2236 1155 2270 1261
rect 36 1087 70 1121
rect 36 1019 70 1053
rect 36 951 70 985
rect 36 883 70 917
rect 2236 1087 2270 1121
rect 2236 1019 2270 1053
rect 2236 951 2270 985
rect 36 727 70 849
rect 2236 883 2270 917
rect 2236 727 2270 849
rect 36 693 192 727
rect 226 693 260 727
rect 294 693 328 727
rect 362 693 396 727
rect 430 693 464 727
rect 498 693 532 727
rect 566 693 600 727
rect 634 693 668 727
rect 702 693 736 727
rect 770 693 804 727
rect 838 693 872 727
rect 906 693 940 727
rect 974 693 1008 727
rect 1042 693 1076 727
rect 1110 693 1144 727
rect 1178 693 1212 727
rect 1246 693 1280 727
rect 1314 693 1348 727
rect 1382 693 1416 727
rect 1450 693 1484 727
rect 1518 693 1552 727
rect 1586 693 1620 727
rect 1654 693 1688 727
rect 1722 693 1756 727
rect 1790 693 1824 727
rect 1858 693 1892 727
rect 1926 693 1960 727
rect 1994 693 2028 727
rect 2062 693 2096 727
rect 2130 693 2270 727
<< psubdiffcont >>
rect 200 553 234 587
rect 268 553 302 587
rect 336 553 370 587
rect 404 553 438 587
rect 472 553 506 587
rect 540 553 574 587
rect 608 553 642 587
rect 676 553 710 587
rect 744 553 778 587
rect 812 553 846 587
rect 880 553 914 587
rect 948 553 982 587
rect 1016 553 1050 587
rect 1084 553 1118 587
rect 1152 553 1186 587
rect 1220 553 1254 587
rect 1288 553 1322 587
rect 1356 553 1390 587
rect 1424 553 1458 587
rect 1492 553 1526 587
rect 1560 553 1594 587
rect 1628 553 1662 587
rect 1696 553 1730 587
rect 1764 553 1798 587
rect 1832 553 1866 587
rect 1900 553 1934 587
rect 1968 553 2002 587
rect 2036 553 2070 587
rect 36 321 70 355
rect 36 253 70 287
rect 36 185 70 219
rect 2236 321 2270 355
rect 2236 253 2270 287
rect 2236 185 2270 219
rect 268 -15 302 19
rect 336 -15 370 19
rect 404 -15 438 19
rect 472 -15 506 19
rect 540 -15 574 19
rect 608 -15 642 19
rect 676 -15 710 19
rect 744 -15 778 19
rect 812 -15 846 19
rect 880 -15 914 19
rect 948 -15 982 19
rect 1016 -15 1050 19
rect 1084 -15 1118 19
rect 1152 -15 1186 19
rect 1220 -15 1254 19
rect 1288 -15 1322 19
rect 1356 -15 1390 19
rect 1424 -15 1458 19
rect 1492 -15 1526 19
rect 1560 -15 1594 19
rect 1628 -15 1662 19
rect 1696 -15 1730 19
rect 1764 -15 1798 19
rect 1832 -15 1866 19
rect 1900 -15 1934 19
rect 1968 -15 2002 19
rect 2036 -15 2070 19
<< nsubdiffcont >>
rect 124 1261 158 1295
rect 192 1261 226 1295
rect 260 1261 294 1295
rect 328 1261 362 1295
rect 396 1261 430 1295
rect 464 1261 498 1295
rect 532 1261 566 1295
rect 600 1261 634 1295
rect 668 1261 702 1295
rect 736 1261 770 1295
rect 804 1261 838 1295
rect 872 1261 906 1295
rect 940 1261 974 1295
rect 1008 1261 1042 1295
rect 1076 1261 1110 1295
rect 1144 1261 1178 1295
rect 1212 1261 1246 1295
rect 1280 1261 1314 1295
rect 1348 1261 1382 1295
rect 1416 1261 1450 1295
rect 1484 1261 1518 1295
rect 1552 1261 1586 1295
rect 1620 1261 1654 1295
rect 1688 1261 1722 1295
rect 1756 1261 1790 1295
rect 1824 1261 1858 1295
rect 1892 1261 1926 1295
rect 1960 1261 1994 1295
rect 2028 1261 2062 1295
rect 2096 1261 2130 1295
rect 36 1121 70 1155
rect 2236 1121 2270 1155
rect 36 1053 70 1087
rect 36 985 70 1019
rect 36 917 70 951
rect 2236 1053 2270 1087
rect 2236 985 2270 1019
rect 2236 917 2270 951
rect 36 849 70 883
rect 2236 849 2270 883
rect 192 693 226 727
rect 260 693 294 727
rect 328 693 362 727
rect 396 693 430 727
rect 464 693 498 727
rect 532 693 566 727
rect 600 693 634 727
rect 668 693 702 727
rect 736 693 770 727
rect 804 693 838 727
rect 872 693 906 727
rect 940 693 974 727
rect 1008 693 1042 727
rect 1076 693 1110 727
rect 1144 693 1178 727
rect 1212 693 1246 727
rect 1280 693 1314 727
rect 1348 693 1382 727
rect 1416 693 1450 727
rect 1484 693 1518 727
rect 1552 693 1586 727
rect 1620 693 1654 727
rect 1688 693 1722 727
rect 1756 693 1790 727
rect 1824 693 1858 727
rect 1892 693 1926 727
rect 1960 693 1994 727
rect 2028 693 2062 727
rect 2096 693 2130 727
<< poly >>
rect 249 1100 329 1126
rect 877 1100 957 1126
rect 1349 1100 1429 1126
rect 1977 1100 2057 1126
rect 249 853 329 900
rect 249 819 272 853
rect 306 819 329 853
rect 249 803 329 819
rect 877 853 957 900
rect 877 819 900 853
rect 934 819 957 853
rect 877 803 957 819
rect 1349 853 1429 900
rect 1349 819 1372 853
rect 1406 819 1429 853
rect 1349 803 1429 819
rect 1977 853 2057 900
rect 1977 819 2000 853
rect 2034 819 2057 853
rect 1977 803 2057 819
rect 249 487 329 503
rect 249 453 272 487
rect 306 453 329 487
rect 249 415 329 453
rect 563 487 643 503
rect 563 453 586 487
rect 620 453 643 487
rect 563 415 643 453
rect 877 487 957 503
rect 877 453 900 487
rect 934 453 957 487
rect 877 415 957 453
rect 1349 487 1429 503
rect 1349 453 1372 487
rect 1406 453 1429 487
rect 1349 415 1429 453
rect 1663 487 1743 503
rect 1663 453 1686 487
rect 1720 453 1743 487
rect 1663 415 1743 453
rect 1977 487 2057 503
rect 1977 453 2000 487
rect 2034 453 2057 487
rect 1977 415 2057 453
rect 249 189 329 215
rect 563 189 643 215
rect 877 189 957 215
rect 1349 189 1429 215
rect 1663 189 1743 215
rect 1977 189 2057 215
<< polycont >>
rect 272 819 306 853
rect 900 819 934 853
rect 1372 819 1406 853
rect 2000 819 2034 853
rect 272 453 306 487
rect 586 453 620 487
rect 900 453 934 487
rect 1372 453 1406 487
rect 1686 453 1720 487
rect 2000 453 2034 487
<< locali >>
rect 36 1261 124 1295
rect 158 1261 192 1295
rect 226 1261 260 1295
rect 294 1261 328 1295
rect 362 1261 367 1295
rect 430 1261 439 1295
rect 498 1261 532 1295
rect 566 1261 567 1295
rect 634 1261 639 1295
rect 702 1261 736 1295
rect 770 1261 804 1295
rect 838 1261 872 1295
rect 906 1261 940 1295
rect 974 1261 1008 1295
rect 1042 1261 1076 1295
rect 1110 1261 1144 1295
rect 1178 1261 1212 1295
rect 1246 1261 1280 1295
rect 1314 1261 1348 1295
rect 1382 1261 1416 1295
rect 1450 1261 1484 1295
rect 1518 1261 1552 1295
rect 1601 1261 1620 1295
rect 1673 1261 1688 1295
rect 1722 1261 1756 1295
rect 1801 1261 1824 1295
rect 1873 1261 1892 1295
rect 1926 1261 1960 1295
rect 1994 1261 2028 1295
rect 2062 1261 2096 1295
rect 2130 1261 2270 1295
rect 36 1155 70 1261
rect 36 1087 70 1121
rect 2236 1155 2270 1261
rect 36 1019 70 1053
rect 36 951 70 985
rect 36 883 70 917
rect 203 1085 237 1104
rect 203 1017 237 1019
rect 203 981 237 983
rect 203 896 237 915
rect 341 1085 375 1104
rect 341 1017 375 1019
rect 341 981 375 983
rect 341 896 375 915
rect 831 1085 865 1104
rect 831 1017 865 1019
rect 831 981 865 983
rect 831 896 865 915
rect 969 1085 1003 1104
rect 969 1017 1003 1019
rect 969 981 1003 983
rect 969 896 1003 915
rect 1303 1085 1337 1104
rect 1303 1017 1337 1019
rect 1303 981 1337 983
rect 1303 896 1337 915
rect 1441 1085 1475 1104
rect 1441 1017 1475 1019
rect 1441 981 1475 983
rect 1441 896 1475 915
rect 1931 1085 1965 1104
rect 1931 1017 1965 1019
rect 1931 981 1965 983
rect 1931 896 1965 915
rect 2069 1085 2103 1104
rect 2069 1017 2103 1019
rect 2069 981 2103 983
rect 2069 896 2103 915
rect 2236 1087 2270 1121
rect 2236 1019 2270 1053
rect 2236 951 2270 985
rect 2236 883 2270 917
rect 36 727 70 849
rect 249 819 272 853
rect 306 819 329 853
rect 877 819 900 853
rect 934 819 957 853
rect 1349 819 1372 853
rect 1406 819 1429 853
rect 1977 819 2000 853
rect 2034 819 2057 853
rect 2236 727 2270 849
rect 36 693 192 727
rect 226 693 260 727
rect 294 693 328 727
rect 362 693 396 727
rect 430 693 464 727
rect 498 693 532 727
rect 566 693 600 727
rect 634 693 668 727
rect 702 693 736 727
rect 770 693 804 727
rect 838 693 872 727
rect 906 693 940 727
rect 974 693 1008 727
rect 1042 693 1076 727
rect 1110 693 1144 727
rect 1178 693 1212 727
rect 1246 693 1280 727
rect 1314 693 1348 727
rect 1382 693 1416 727
rect 1450 693 1484 727
rect 1518 693 1552 727
rect 1586 693 1620 727
rect 1654 693 1688 727
rect 1722 693 1756 727
rect 1790 693 1824 727
rect 1858 693 1892 727
rect 1926 693 1960 727
rect 1994 693 2028 727
rect 2062 693 2096 727
rect 2130 693 2270 727
rect 36 553 200 587
rect 234 553 268 587
rect 302 553 336 587
rect 370 553 404 587
rect 438 553 472 587
rect 506 553 540 587
rect 574 553 608 587
rect 642 553 676 587
rect 710 553 744 587
rect 778 553 812 587
rect 846 553 880 587
rect 914 553 948 587
rect 982 553 1016 587
rect 1050 553 1084 587
rect 1118 553 1152 587
rect 1186 553 1220 587
rect 1254 553 1288 587
rect 1322 553 1356 587
rect 1390 553 1424 587
rect 1458 553 1492 587
rect 1526 553 1560 587
rect 1594 553 1628 587
rect 1662 553 1696 587
rect 1730 553 1764 587
rect 1798 553 1832 587
rect 1866 553 1900 587
rect 1934 553 1968 587
rect 2002 553 2036 587
rect 2070 553 2270 587
rect 36 355 70 553
rect 249 453 272 487
rect 306 453 329 487
rect 563 453 586 487
rect 620 453 643 487
rect 877 453 900 487
rect 934 453 957 487
rect 1349 453 1372 487
rect 1406 453 1429 487
rect 1663 453 1686 487
rect 1720 453 1743 487
rect 1977 453 2000 487
rect 2034 453 2057 487
rect 36 287 70 321
rect 36 219 70 253
rect 203 400 237 419
rect 203 332 237 334
rect 203 296 237 298
rect 203 211 237 230
rect 341 400 375 419
rect 341 332 375 334
rect 341 296 375 298
rect 341 211 375 230
rect 517 400 551 419
rect 517 332 551 334
rect 517 296 551 298
rect 517 211 551 230
rect 655 400 689 419
rect 655 332 689 334
rect 655 296 689 298
rect 655 211 689 230
rect 831 400 865 419
rect 831 332 865 334
rect 831 296 865 298
rect 831 211 865 230
rect 969 400 1003 419
rect 969 332 1003 334
rect 969 296 1003 298
rect 969 211 1003 230
rect 1303 400 1337 419
rect 1303 332 1337 334
rect 1303 296 1337 298
rect 1303 211 1337 230
rect 1441 400 1475 419
rect 1441 332 1475 334
rect 1441 296 1475 298
rect 1441 211 1475 230
rect 1617 400 1651 419
rect 1617 332 1651 334
rect 1617 296 1651 298
rect 1617 211 1651 230
rect 1755 400 1789 419
rect 1755 332 1789 334
rect 1755 296 1789 298
rect 1755 211 1789 230
rect 1931 400 1965 419
rect 1931 332 1965 334
rect 1931 296 1965 298
rect 1931 211 1965 230
rect 2069 400 2103 419
rect 2069 332 2103 334
rect 2069 296 2103 298
rect 2069 211 2103 230
rect 2236 355 2270 553
rect 2236 287 2270 321
rect 2236 219 2270 253
rect 36 19 70 185
rect 2236 19 2270 185
rect 36 -15 268 19
rect 302 -15 336 19
rect 370 -15 404 19
rect 438 -15 454 19
rect 506 -15 526 19
rect 574 -15 608 19
rect 642 -15 654 19
rect 710 -15 726 19
rect 778 -15 812 19
rect 846 -15 854 19
rect 914 -15 926 19
rect 982 -15 1016 19
rect 1050 -15 1054 19
rect 1118 -15 1126 19
rect 1186 -15 1220 19
rect 1322 -15 1326 19
rect 1390 -15 1424 19
rect 1488 -15 1492 19
rect 1594 -15 1628 19
rect 1688 -15 1696 19
rect 1760 -15 1764 19
rect 1798 -15 1832 19
rect 1866 -15 1900 19
rect 1934 -15 1968 19
rect 2002 -15 2036 19
rect 2070 -15 2270 19
<< viali >>
rect 367 1261 396 1295
rect 396 1261 401 1295
rect 439 1261 464 1295
rect 464 1261 473 1295
rect 567 1261 600 1295
rect 600 1261 601 1295
rect 639 1261 668 1295
rect 668 1261 673 1295
rect 1567 1261 1586 1295
rect 1586 1261 1601 1295
rect 1639 1261 1654 1295
rect 1654 1261 1673 1295
rect 1767 1261 1790 1295
rect 1790 1261 1801 1295
rect 1839 1261 1858 1295
rect 1858 1261 1873 1295
rect 203 1051 237 1053
rect 203 1019 237 1051
rect 203 949 237 981
rect 203 947 237 949
rect 341 1051 375 1053
rect 341 1019 375 1051
rect 341 949 375 981
rect 341 947 375 949
rect 831 1051 865 1053
rect 831 1019 865 1051
rect 831 949 865 981
rect 831 947 865 949
rect 969 1051 1003 1053
rect 969 1019 1003 1051
rect 969 949 1003 981
rect 969 947 1003 949
rect 1303 1051 1337 1053
rect 1303 1019 1337 1051
rect 1303 949 1337 981
rect 1303 947 1337 949
rect 1441 1051 1475 1053
rect 1441 1019 1475 1051
rect 1441 949 1475 981
rect 1441 947 1475 949
rect 1931 1051 1965 1053
rect 1931 1019 1965 1051
rect 1931 949 1965 981
rect 1931 947 1965 949
rect 2069 1051 2103 1053
rect 2069 1019 2103 1051
rect 2069 949 2103 981
rect 2069 947 2103 949
rect 272 819 306 853
rect 900 819 934 853
rect 1372 819 1406 853
rect 2000 819 2034 853
rect 272 453 306 487
rect 586 453 620 487
rect 900 453 934 487
rect 1372 453 1406 487
rect 1686 453 1720 487
rect 2000 453 2034 487
rect 203 366 237 368
rect 203 334 237 366
rect 203 264 237 296
rect 203 262 237 264
rect 341 366 375 368
rect 341 334 375 366
rect 341 264 375 296
rect 341 262 375 264
rect 517 366 551 368
rect 517 334 551 366
rect 517 264 551 296
rect 517 262 551 264
rect 655 366 689 368
rect 655 334 689 366
rect 655 264 689 296
rect 655 262 689 264
rect 831 366 865 368
rect 831 334 865 366
rect 831 264 865 296
rect 831 262 865 264
rect 969 366 1003 368
rect 969 334 1003 366
rect 969 264 1003 296
rect 969 262 1003 264
rect 1303 366 1337 368
rect 1303 334 1337 366
rect 1303 264 1337 296
rect 1303 262 1337 264
rect 1441 366 1475 368
rect 1441 334 1475 366
rect 1441 264 1475 296
rect 1441 262 1475 264
rect 1617 366 1651 368
rect 1617 334 1651 366
rect 1617 264 1651 296
rect 1617 262 1651 264
rect 1755 366 1789 368
rect 1755 334 1789 366
rect 1755 264 1789 296
rect 1755 262 1789 264
rect 1931 366 1965 368
rect 1931 334 1965 366
rect 1931 264 1965 296
rect 1931 262 1965 264
rect 2069 366 2103 368
rect 2069 334 2103 366
rect 2069 264 2103 296
rect 2069 262 2103 264
rect 454 -15 472 19
rect 472 -15 488 19
rect 526 -15 540 19
rect 540 -15 560 19
rect 654 -15 676 19
rect 676 -15 688 19
rect 726 -15 744 19
rect 744 -15 760 19
rect 854 -15 880 19
rect 880 -15 888 19
rect 926 -15 948 19
rect 948 -15 960 19
rect 1054 -15 1084 19
rect 1084 -15 1088 19
rect 1126 -15 1152 19
rect 1152 -15 1160 19
rect 1254 -15 1288 19
rect 1326 -15 1356 19
rect 1356 -15 1360 19
rect 1454 -15 1458 19
rect 1458 -15 1488 19
rect 1526 -15 1560 19
rect 1654 -15 1662 19
rect 1662 -15 1688 19
rect 1726 -15 1730 19
rect 1730 -15 1760 19
<< metal1 >>
rect 150 1304 918 1308
rect 150 1252 162 1304
rect 214 1252 226 1304
rect 278 1295 790 1304
rect 278 1261 367 1295
rect 401 1261 439 1295
rect 473 1261 567 1295
rect 601 1261 639 1295
rect 673 1261 790 1295
rect 278 1252 790 1261
rect 842 1252 854 1304
rect 906 1252 918 1304
rect 150 1248 918 1252
rect 197 1053 243 1248
rect 197 1019 203 1053
rect 237 1019 243 1053
rect 197 981 243 1019
rect 197 947 203 981
rect 237 947 243 981
rect 197 900 243 947
rect 335 1070 381 1100
rect 335 1058 395 1070
rect 335 1006 339 1058
rect 391 1006 395 1058
rect 335 994 395 1006
rect 335 942 339 994
rect 391 942 395 994
rect 335 930 395 942
rect 825 1053 871 1248
rect 825 1019 831 1053
rect 865 1019 871 1053
rect 825 981 871 1019
rect 825 947 831 981
rect 865 947 871 981
rect 335 900 381 930
rect 825 900 871 947
rect 963 1070 1009 1100
rect 963 1058 1023 1070
rect 963 1006 967 1058
rect 1019 1006 1023 1058
rect 963 994 1023 1006
rect 963 942 967 994
rect 1019 942 1023 994
rect 963 930 1023 942
rect 963 900 1009 930
rect 1123 859 1183 1348
rect 1361 1304 2156 1308
rect 1361 1252 1400 1304
rect 1452 1252 1464 1304
rect 1516 1295 2028 1304
rect 1516 1261 1567 1295
rect 1601 1261 1639 1295
rect 1673 1261 1767 1295
rect 1801 1261 1839 1295
rect 1873 1261 2028 1295
rect 1516 1252 2028 1261
rect 2080 1252 2092 1304
rect 2144 1252 2156 1304
rect 1361 1248 2156 1252
rect 1297 1070 1343 1100
rect 1283 1058 1343 1070
rect 1283 1006 1287 1058
rect 1339 1006 1343 1058
rect 1283 994 1343 1006
rect 1283 942 1287 994
rect 1339 942 1343 994
rect 1283 930 1343 942
rect 1297 900 1343 930
rect 1435 1053 1481 1248
rect 1925 1070 1971 1100
rect 1435 1019 1441 1053
rect 1475 1019 1481 1053
rect 1435 981 1481 1019
rect 1435 947 1441 981
rect 1475 947 1481 981
rect 1435 900 1481 947
rect 1911 1058 1971 1070
rect 1911 1006 1915 1058
rect 1967 1006 1971 1058
rect 1911 994 1971 1006
rect 1911 942 1915 994
rect 1967 942 1971 994
rect 1911 930 1971 942
rect 1925 900 1971 930
rect 2063 1053 2109 1248
rect 2063 1019 2069 1053
rect 2103 1019 2109 1053
rect 2063 981 2109 1019
rect 2063 947 2069 981
rect 2103 947 2109 981
rect 2063 900 2109 947
rect 253 853 325 859
rect 253 819 272 853
rect 306 819 325 853
rect 253 683 325 819
rect 881 853 953 859
rect 881 819 900 853
rect 934 819 953 853
rect 53 623 325 683
rect 253 487 325 623
rect 398 711 458 723
rect 398 659 402 711
rect 454 683 458 711
rect 881 683 953 819
rect 1033 853 1425 859
rect 1033 819 1372 853
rect 1406 819 1425 853
rect 1033 813 1425 819
rect 1033 723 1079 813
rect 454 659 633 683
rect 398 647 633 659
rect 398 595 402 647
rect 454 623 633 647
rect 454 595 458 623
rect 398 583 458 595
rect 573 493 633 623
rect 725 623 953 683
rect 253 453 272 487
rect 306 453 325 487
rect 253 447 325 453
rect 567 487 639 493
rect 567 453 586 487
rect 620 453 639 487
rect 567 447 639 453
rect 725 415 785 623
rect 881 493 953 623
rect 1026 711 1086 723
rect 1026 659 1030 711
rect 1082 659 1086 711
rect 1026 647 1086 659
rect 1026 595 1030 647
rect 1082 595 1086 647
rect 1026 583 1086 595
rect 1220 711 1280 723
rect 1220 659 1224 711
rect 1276 659 1280 711
rect 1220 647 1280 659
rect 1220 595 1224 647
rect 1276 595 1280 647
rect 1220 583 1280 595
rect 1353 683 1425 813
rect 1981 853 2053 859
rect 1981 819 2000 853
rect 2034 819 2053 853
rect 1848 711 1908 723
rect 1848 683 1852 711
rect 1353 623 1581 683
rect 1226 493 1272 583
rect 881 487 1272 493
rect 881 453 900 487
rect 934 453 1272 487
rect 881 447 1272 453
rect 1353 487 1425 623
rect 1353 453 1372 487
rect 1406 453 1425 487
rect 1353 447 1425 453
rect 1521 415 1581 623
rect 1673 659 1852 683
rect 1904 659 1908 711
rect 1673 647 1908 659
rect 1673 623 1852 647
rect 1673 493 1733 623
rect 1848 595 1852 623
rect 1904 595 1908 647
rect 1848 583 1908 595
rect 1981 683 2053 819
rect 1981 623 2253 683
rect 1667 487 1739 493
rect 1667 453 1686 487
rect 1720 453 1739 487
rect 1667 447 1739 453
rect 1981 487 2053 623
rect 1981 453 2000 487
rect 2034 453 2053 487
rect 1981 447 2053 453
rect 197 368 243 415
rect 197 334 203 368
rect 237 334 243 368
rect 197 296 243 334
rect 197 262 203 296
rect 237 262 243 296
rect 197 32 243 262
rect 335 385 381 415
rect 335 373 395 385
rect 335 321 339 373
rect 391 321 395 373
rect 335 309 395 321
rect 335 257 339 309
rect 391 257 395 309
rect 335 245 395 257
rect 511 368 557 415
rect 511 334 517 368
rect 551 334 557 368
rect 511 296 557 334
rect 511 262 517 296
rect 551 262 557 296
rect 335 215 381 245
rect 511 32 557 262
rect 649 368 785 415
rect 649 334 655 368
rect 689 355 785 368
rect 825 368 871 415
rect 689 334 695 355
rect 649 296 695 334
rect 649 262 655 296
rect 689 262 695 296
rect 649 215 695 262
rect 825 334 831 368
rect 865 334 871 368
rect 825 296 871 334
rect 825 262 831 296
rect 865 262 871 296
rect 825 32 871 262
rect 963 385 1009 415
rect 1297 385 1343 415
rect 963 373 1023 385
rect 963 321 967 373
rect 1019 321 1023 373
rect 963 309 1023 321
rect 963 257 967 309
rect 1019 257 1023 309
rect 963 245 1023 257
rect 1283 373 1343 385
rect 1283 321 1287 373
rect 1339 321 1343 373
rect 1283 309 1343 321
rect 1283 257 1287 309
rect 1339 257 1343 309
rect 1283 245 1343 257
rect 963 215 1009 245
rect 1297 215 1343 245
rect 1435 368 1481 415
rect 1435 334 1441 368
rect 1475 334 1481 368
rect 1521 368 1657 415
rect 1521 355 1617 368
rect 1435 296 1481 334
rect 1435 262 1441 296
rect 1475 262 1481 296
rect 1435 32 1481 262
rect 1611 334 1617 355
rect 1651 334 1657 368
rect 1611 296 1657 334
rect 1611 262 1617 296
rect 1651 262 1657 296
rect 1611 215 1657 262
rect 1749 368 1795 415
rect 1925 385 1971 415
rect 1749 334 1755 368
rect 1789 334 1795 368
rect 1749 296 1795 334
rect 1749 262 1755 296
rect 1789 262 1795 296
rect 1749 32 1795 262
rect 1911 373 1971 385
rect 1911 321 1915 373
rect 1967 321 1971 373
rect 1911 309 1971 321
rect 1911 257 1915 309
rect 1967 257 1971 309
rect 1911 245 1971 257
rect 1925 215 1971 245
rect 2063 368 2109 415
rect 2063 334 2069 368
rect 2103 334 2109 368
rect 2063 296 2109 334
rect 2063 262 2069 296
rect 2103 262 2109 296
rect 2063 32 2109 262
rect 150 28 2156 32
rect 150 -24 162 28
rect 214 -24 226 28
rect 278 19 476 28
rect 528 19 540 28
rect 592 19 790 28
rect 278 -15 454 19
rect 592 -15 654 19
rect 688 -15 726 19
rect 760 -15 790 19
rect 278 -24 476 -15
rect 528 -24 540 -15
rect 592 -24 790 -15
rect 842 -24 854 28
rect 906 19 1400 28
rect 906 -15 926 19
rect 960 -15 1054 19
rect 1088 -15 1126 19
rect 1160 -15 1254 19
rect 1288 -15 1326 19
rect 1360 -15 1400 19
rect 906 -24 1400 -15
rect 1452 19 1464 28
rect 1516 19 1714 28
rect 1452 -15 1454 19
rect 1516 -15 1526 19
rect 1560 -15 1654 19
rect 1688 -15 1714 19
rect 1452 -24 1464 -15
rect 1516 -24 1714 -15
rect 1766 -24 1778 28
rect 1830 -24 2028 28
rect 2080 -24 2092 28
rect 2144 -24 2156 28
rect 150 -28 2156 -24
<< via1 >>
rect 162 1252 214 1304
rect 226 1252 278 1304
rect 790 1252 842 1304
rect 854 1252 906 1304
rect 339 1053 391 1058
rect 339 1019 341 1053
rect 341 1019 375 1053
rect 375 1019 391 1053
rect 339 1006 391 1019
rect 339 981 391 994
rect 339 947 341 981
rect 341 947 375 981
rect 375 947 391 981
rect 339 942 391 947
rect 967 1053 1019 1058
rect 967 1019 969 1053
rect 969 1019 1003 1053
rect 1003 1019 1019 1053
rect 967 1006 1019 1019
rect 967 981 1019 994
rect 967 947 969 981
rect 969 947 1003 981
rect 1003 947 1019 981
rect 967 942 1019 947
rect 1400 1252 1452 1304
rect 1464 1252 1516 1304
rect 2028 1252 2080 1304
rect 2092 1252 2144 1304
rect 1287 1053 1339 1058
rect 1287 1019 1303 1053
rect 1303 1019 1337 1053
rect 1337 1019 1339 1053
rect 1287 1006 1339 1019
rect 1287 981 1339 994
rect 1287 947 1303 981
rect 1303 947 1337 981
rect 1337 947 1339 981
rect 1287 942 1339 947
rect 1915 1053 1967 1058
rect 1915 1019 1931 1053
rect 1931 1019 1965 1053
rect 1965 1019 1967 1053
rect 1915 1006 1967 1019
rect 1915 981 1967 994
rect 1915 947 1931 981
rect 1931 947 1965 981
rect 1965 947 1967 981
rect 1915 942 1967 947
rect 402 659 454 711
rect 402 595 454 647
rect 1030 659 1082 711
rect 1030 595 1082 647
rect 1224 659 1276 711
rect 1224 595 1276 647
rect 1852 659 1904 711
rect 1852 595 1904 647
rect 339 368 391 373
rect 339 334 341 368
rect 341 334 375 368
rect 375 334 391 368
rect 339 321 391 334
rect 339 296 391 309
rect 339 262 341 296
rect 341 262 375 296
rect 375 262 391 296
rect 339 257 391 262
rect 967 368 1019 373
rect 967 334 969 368
rect 969 334 1003 368
rect 1003 334 1019 368
rect 967 321 1019 334
rect 967 296 1019 309
rect 967 262 969 296
rect 969 262 1003 296
rect 1003 262 1019 296
rect 967 257 1019 262
rect 1287 368 1339 373
rect 1287 334 1303 368
rect 1303 334 1337 368
rect 1337 334 1339 368
rect 1287 321 1339 334
rect 1287 296 1339 309
rect 1287 262 1303 296
rect 1303 262 1337 296
rect 1337 262 1339 296
rect 1287 257 1339 262
rect 1915 368 1967 373
rect 1915 334 1931 368
rect 1931 334 1965 368
rect 1965 334 1967 368
rect 1915 321 1967 334
rect 1915 296 1967 309
rect 1915 262 1931 296
rect 1931 262 1965 296
rect 1965 262 1967 296
rect 1915 257 1967 262
rect 162 -24 214 28
rect 226 -24 278 28
rect 476 19 528 28
rect 540 19 592 28
rect 476 -15 488 19
rect 488 -15 526 19
rect 526 -15 528 19
rect 540 -15 560 19
rect 560 -15 592 19
rect 476 -24 528 -15
rect 540 -24 592 -15
rect 790 -24 842 28
rect 854 19 906 28
rect 854 -15 888 19
rect 888 -15 906 19
rect 854 -24 906 -15
rect 1400 -24 1452 28
rect 1464 19 1516 28
rect 1714 19 1766 28
rect 1464 -15 1488 19
rect 1488 -15 1516 19
rect 1714 -15 1726 19
rect 1726 -15 1760 19
rect 1760 -15 1766 19
rect 1464 -24 1516 -15
rect 1714 -24 1766 -15
rect 1778 -24 1830 28
rect 2028 -24 2080 28
rect 2092 -24 2144 28
<< metal2 >>
rect 160 1304 2146 1318
rect 160 1252 162 1304
rect 214 1252 226 1304
rect 278 1252 790 1304
rect 842 1252 854 1304
rect 906 1252 1400 1304
rect 1452 1252 1464 1304
rect 1516 1252 2028 1304
rect 2080 1252 2092 1304
rect 2144 1252 2146 1304
rect 160 1238 2146 1252
rect 325 1058 405 1060
rect 325 1006 339 1058
rect 391 1006 405 1058
rect 325 994 405 1006
rect 325 942 339 994
rect 391 942 405 994
rect 325 940 405 942
rect 953 1058 1033 1060
rect 953 1006 967 1058
rect 1019 1006 1033 1058
rect 953 994 1033 1006
rect 953 942 967 994
rect 1019 942 1033 994
rect 953 940 1033 942
rect 1273 1058 1353 1060
rect 1273 1006 1287 1058
rect 1339 1006 1353 1058
rect 1273 994 1353 1006
rect 1273 942 1287 994
rect 1339 942 1353 994
rect 1273 940 1353 942
rect 1901 1058 1981 1060
rect 1901 1006 1915 1058
rect 1967 1006 1981 1058
rect 1901 994 1981 1006
rect 1901 942 1915 994
rect 1967 942 1981 994
rect 1901 940 1981 942
rect 342 713 388 940
rect 970 713 1016 940
rect 1290 713 1336 940
rect 1918 713 1964 940
rect 342 711 468 713
rect 342 659 402 711
rect 454 659 468 711
rect 342 647 468 659
rect 342 595 402 647
rect 454 595 468 647
rect 342 593 468 595
rect 970 711 1096 713
rect 970 659 1030 711
rect 1082 659 1096 711
rect 970 647 1096 659
rect 970 595 1030 647
rect 1082 595 1096 647
rect 970 593 1096 595
rect 1210 711 1336 713
rect 1210 659 1224 711
rect 1276 659 1336 711
rect 1210 647 1336 659
rect 1210 595 1224 647
rect 1276 595 1336 647
rect 1210 593 1336 595
rect 1838 711 1964 713
rect 1838 659 1852 711
rect 1904 659 1964 711
rect 1838 647 1964 659
rect 1838 595 1852 647
rect 1904 595 1964 647
rect 1838 593 1964 595
rect 342 375 388 593
rect 970 375 1016 593
rect 1290 375 1336 593
rect 1918 375 1964 593
rect 325 373 405 375
rect 325 321 339 373
rect 391 321 405 373
rect 325 309 405 321
rect 325 257 339 309
rect 391 257 405 309
rect 325 255 405 257
rect 953 373 1033 375
rect 953 321 967 373
rect 1019 321 1033 373
rect 953 309 1033 321
rect 953 257 967 309
rect 1019 257 1033 309
rect 953 255 1033 257
rect 1273 373 1353 375
rect 1273 321 1287 373
rect 1339 321 1353 373
rect 1273 309 1353 321
rect 1273 257 1287 309
rect 1339 257 1353 309
rect 1273 255 1353 257
rect 1901 373 1981 375
rect 1901 321 1915 373
rect 1967 321 1981 373
rect 1901 309 1981 321
rect 1901 257 1915 309
rect 1967 257 1981 309
rect 1901 255 1981 257
rect 160 28 2146 42
rect 160 -24 162 28
rect 214 -24 226 28
rect 278 -24 476 28
rect 528 -24 540 28
rect 592 -24 790 28
rect 842 -24 854 28
rect 906 -24 1400 28
rect 1452 -24 1464 28
rect 1516 -24 1714 28
rect 1766 -24 1778 28
rect 1830 -24 2028 28
rect 2080 -24 2092 28
rect 2144 -24 2146 28
rect 160 -38 2146 -24
<< labels >>
flabel metal2 s 160 1238 203 1318 2 FreeSans 44 0 0 0 vdd
port 2 nsew
flabel metal2 s 160 -38 203 42 2 FreeSans 44 0 0 0 vss
port 3 nsew
flabel metal1 s 1104 447 1178 493 1 FreeSans 44 0 0 0 Qn
port 5 nsew
flabel metal1 s 53 623 83 683 1 FreeSans 44 0 0 0 S
port 6 nsew
flabel metal1 s 2223 623 2253 683 1 FreeSans 44 0 0 0 R
port 7 nsew
flabel metal1 s 1123 1318 1183 1348 1 FreeSans 44 0 0 0 Q
port 8 nsew
<< end >>
