* NGSPICE file created from comparator.ext - technology: sky130B

.subckt sky130_fd_pr__cap_mim_m3_1_FJFAMD m3_n386_n240# c1_n346_n200#
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt trimcap cp cn
XXC2 cn cp sky130_fd_pr__cap_mim_m3_1_FJFAMD
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_E33R59 G D S
X0 D G S S sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.32 ps=2.64 w=1 l=0.3
.ends

.subckt nfet_mimcap_combo sky130_fd_pr__nfet_01v8_lvt_E33R59_0/G trimcap_1/cn trimcap_1/cp
+ VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_E33R59_0 sky130_fd_pr__nfet_01v8_lvt_E33R59_0/G trimcap_1/cn
+ VSUBS sky130_fd_pr__nfet_01v8_lvt_E33R59
Xtrimcap_1 trimcap_1/cp trimcap_1/cn trimcap
.ends

.subckt nfet_2mimcap_combo VSUBS nfet_mimcap_combo_0/sky130_fd_pr__nfet_01v8_lvt_E33R59_0/G
+ trimcap_0/cn trimcap_0/cp
Xtrimcap_0 trimcap_0/cp trimcap_0/cn trimcap
Xnfet_mimcap_combo_0 nfet_mimcap_combo_0/sky130_fd_pr__nfet_01v8_lvt_E33R59_0/G trimcap_0/cn
+ trimcap_0/cp VSUBS nfet_mimcap_combo
.ends

.subckt nfet_4mimcap_combo VSUBS trimcap_1/cn trimcap_1/cp nfet_2mimcap_combo_1/nfet_mimcap_combo_0/sky130_fd_pr__nfet_01v8_lvt_E33R59_0/G
Xtrimcap_0 trimcap_1/cp trimcap_1/cn trimcap
Xtrimcap_1 trimcap_1/cp trimcap_1/cn trimcap
Xnfet_2mimcap_combo_1 VSUBS nfet_2mimcap_combo_1/nfet_mimcap_combo_0/sky130_fd_pr__nfet_01v8_lvt_E33R59_0/G
+ trimcap_1/cn trimcap_1/cp nfet_2mimcap_combo
.ends

.subckt nfet_8mimcap_combo nfet_4mimcap_combo_1/nfet_2mimcap_combo_1/nfet_mimcap_combo_0/sky130_fd_pr__nfet_01v8_lvt_E33R59_0/G
+ trimcap_4/cp VSUBS
Xnfet_4mimcap_combo_1 VSUBS trimcap_4/cn trimcap_4/cp nfet_4mimcap_combo_1/nfet_2mimcap_combo_1/nfet_mimcap_combo_0/sky130_fd_pr__nfet_01v8_lvt_E33R59_0/G
+ nfet_4mimcap_combo
Xtrimcap_0 trimcap_4/cp trimcap_4/cn trimcap
Xtrimcap_1 trimcap_4/cp trimcap_4/cn trimcap
Xtrimcap_2 trimcap_4/cp trimcap_4/cn trimcap
Xtrimcap_3 trimcap_4/cp trimcap_4/cn trimcap
Xtrimcap_4 trimcap_4/cp trimcap_4/cn trimcap
.ends

.subckt trim VSS d0 d1 d2 d3 d4 drain
Xnfet_4mimcap_combo_0 VSS nfet_4mimcap_combo_0/trimcap_1/cn drain d3 nfet_4mimcap_combo
Xnfet_8mimcap_combo_0 d4 drain VSS nfet_8mimcap_combo
Xnfet_2mimcap_combo_0 VSS d2 nfet_2mimcap_combo_0/trimcap_0/cn drain nfet_2mimcap_combo
Xnfet_mimcap_combo_0 d0 nfet_mimcap_combo_0/trimcap_1/cn drain VSS nfet_mimcap_combo
Xnfet_mimcap_combo_1 d1 nfet_mimcap_combo_1/trimcap_1/cn drain VSS nfet_mimcap_combo
.ends

.subckt sky130_fd_pr__nfet_01v8_96AECY G D B S
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt sky130_fd_pr__pfet_01v8_7G6J3C G D B S
X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt comparator vss clk trim0 trim1 trim2 trim3 trim4 trimb0 trimb1 trimb2 trimb3
+ trimb4 vdd
Xtrim_0 vss trim0 trim1 trim2 trim3 trim4 IN trim
Xtrim_1 vss trimb0 trimb1 trimb2 trimb3 trimb4 vdd trim
Xsky130_fd_pr__nfet_01v8_96AECY_0 vdd clk vss IN sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__nfet_01v8_96AECY_1 sky130_fd_pr__nfet_01v8_96AECY_1/G vdd vss vss sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__nfet_01v8_96AECY_2 clk vdd vss vdd sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__nfet_01v8_96AECY_3 sky130_fd_pr__nfet_01v8_96AECY_3/G IN vss vss sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__nfet_01v8_96AECY_5 sky130_fd_pr__nfet_01v8_96AECY_5/G vss vss vss sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__nfet_01v8_96AECY_4 sky130_fd_pr__nfet_01v8_96AECY_4/G vss vss vss sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__pfet_01v8_7G6J3C_0 clk IN vdd vdd sky130_fd_pr__pfet_01v8_7G6J3C
Xsky130_fd_pr__pfet_01v8_7G6J3C_1 vdd clk vdd vdd sky130_fd_pr__pfet_01v8_7G6J3C
Xsky130_fd_pr__pfet_01v8_7G6J3C_2 clk clk vdd vdd sky130_fd_pr__pfet_01v8_7G6J3C
X0 vdd clk vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X1 vdd clk vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=2.61 ps=23.2 w=1 l=0.3
X2 vdd clk vdd vdd sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.3
.ends

