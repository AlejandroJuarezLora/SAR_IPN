magic
tech sky130B
magscale 1 2
timestamp 1696984848
<< error_p >>
rect -560 145 -502 151
rect -442 145 -384 151
rect -324 145 -266 151
rect -206 145 -148 151
rect -88 145 -30 151
rect 30 145 88 151
rect 148 145 206 151
rect 266 145 324 151
rect 384 145 442 151
rect 502 145 560 151
rect -560 111 -548 145
rect -442 111 -430 145
rect -324 111 -312 145
rect -206 111 -194 145
rect -88 111 -76 145
rect 30 111 42 145
rect 148 111 160 145
rect 266 111 278 145
rect 384 111 396 145
rect 502 111 514 145
rect -560 105 -502 111
rect -442 105 -384 111
rect -324 105 -266 111
rect -206 105 -148 111
rect -88 105 -30 111
rect 30 105 88 111
rect 148 105 206 111
rect 266 105 324 111
rect 384 105 442 111
rect 502 105 560 111
<< nwell >>
rect -757 -284 757 284
<< pmos >>
rect -561 -136 -501 64
rect -443 -136 -383 64
rect -325 -136 -265 64
rect -207 -136 -147 64
rect -89 -136 -29 64
rect 29 -136 89 64
rect 147 -136 207 64
rect 265 -136 325 64
rect 383 -136 443 64
rect 501 -136 561 64
<< pdiff >>
rect -619 34 -561 64
rect -619 -106 -607 34
rect -573 -106 -561 34
rect -619 -136 -561 -106
rect -501 34 -443 64
rect -501 -106 -489 34
rect -455 -106 -443 34
rect -501 -136 -443 -106
rect -383 34 -325 64
rect -383 -106 -371 34
rect -337 -106 -325 34
rect -383 -136 -325 -106
rect -265 34 -207 64
rect -265 -106 -253 34
rect -219 -106 -207 34
rect -265 -136 -207 -106
rect -147 34 -89 64
rect -147 -106 -135 34
rect -101 -106 -89 34
rect -147 -136 -89 -106
rect -29 34 29 64
rect -29 -106 -17 34
rect 17 -106 29 34
rect -29 -136 29 -106
rect 89 34 147 64
rect 89 -106 101 34
rect 135 -106 147 34
rect 89 -136 147 -106
rect 207 34 265 64
rect 207 -106 219 34
rect 253 -106 265 34
rect 207 -136 265 -106
rect 325 34 383 64
rect 325 -106 337 34
rect 371 -106 383 34
rect 325 -136 383 -106
rect 443 34 501 64
rect 443 -106 455 34
rect 489 -106 501 34
rect 443 -136 501 -106
rect 561 34 619 64
rect 561 -106 573 34
rect 607 -106 619 34
rect 561 -136 619 -106
<< pdiffc >>
rect -607 -106 -573 34
rect -489 -106 -455 34
rect -371 -106 -337 34
rect -253 -106 -219 34
rect -135 -106 -101 34
rect -17 -106 17 34
rect 101 -106 135 34
rect 219 -106 253 34
rect 337 -106 371 34
rect 455 -106 489 34
rect 573 -106 607 34
<< nsubdiff >>
rect -721 214 -500 248
rect 500 214 721 248
rect -721 121 -687 214
rect 687 121 721 214
rect -721 -214 -687 -121
rect 687 -214 721 -121
rect -721 -248 721 -214
<< nsubdiffcont >>
rect -500 214 500 248
rect -721 -121 -687 121
rect 687 -121 721 121
<< poly >>
rect -564 145 -498 161
rect -564 111 -548 145
rect -514 111 -498 145
rect -564 95 -498 111
rect -446 145 -380 161
rect -446 111 -430 145
rect -396 111 -380 145
rect -446 95 -380 111
rect -328 145 -262 161
rect -328 111 -312 145
rect -278 111 -262 145
rect -328 95 -262 111
rect -210 145 -144 161
rect -210 111 -194 145
rect -160 111 -144 145
rect -210 95 -144 111
rect -92 145 -26 161
rect -92 111 -76 145
rect -42 111 -26 145
rect -92 95 -26 111
rect 26 145 92 161
rect 26 111 42 145
rect 76 111 92 145
rect 26 95 92 111
rect 144 145 210 161
rect 144 111 160 145
rect 194 111 210 145
rect 144 95 210 111
rect 262 145 328 161
rect 262 111 278 145
rect 312 111 328 145
rect 262 95 328 111
rect 380 145 446 161
rect 380 111 396 145
rect 430 111 446 145
rect 380 95 446 111
rect 498 145 564 161
rect 498 111 514 145
rect 548 111 564 145
rect 498 95 564 111
rect -561 64 -501 95
rect -443 64 -383 95
rect -325 64 -265 95
rect -207 64 -147 95
rect -89 64 -29 95
rect 29 64 89 95
rect 147 64 207 95
rect 265 64 325 95
rect 383 64 443 95
rect 501 64 561 95
rect -561 -162 -501 -136
rect -443 -162 -383 -136
rect -325 -162 -265 -136
rect -207 -162 -147 -136
rect -89 -162 -29 -136
rect 29 -162 89 -136
rect 147 -162 207 -136
rect 265 -162 325 -136
rect 383 -162 443 -136
rect 501 -162 561 -136
<< polycont >>
rect -548 111 -514 145
rect -430 111 -396 145
rect -312 111 -278 145
rect -194 111 -160 145
rect -76 111 -42 145
rect 42 111 76 145
rect 160 111 194 145
rect 278 111 312 145
rect 396 111 430 145
rect 514 111 548 145
<< locali >>
rect -516 214 -500 248
rect 500 214 516 248
rect -721 121 -687 137
rect -564 111 -548 145
rect -514 111 -498 145
rect -446 111 -430 145
rect -396 111 -380 145
rect -328 111 -312 145
rect -278 111 -262 145
rect -210 111 -194 145
rect -160 111 -144 145
rect -92 111 -76 145
rect -42 111 -26 145
rect 26 111 42 145
rect 76 111 92 145
rect 144 111 160 145
rect 194 111 210 145
rect 262 111 278 145
rect 312 111 328 145
rect 380 111 396 145
rect 430 111 446 145
rect 498 111 514 145
rect 548 111 564 145
rect 687 121 721 137
rect -721 -137 -687 -121
rect -607 34 -573 50
rect -607 -122 -573 -106
rect -489 34 -455 50
rect -489 -122 -455 -106
rect -371 34 -337 50
rect -371 -122 -337 -106
rect -253 34 -219 50
rect -253 -122 -219 -106
rect -135 34 -101 50
rect -135 -122 -101 -106
rect -17 34 17 50
rect -17 -122 17 -106
rect 101 34 135 50
rect 101 -122 135 -106
rect 219 34 253 50
rect 219 -122 253 -106
rect 337 34 371 50
rect 337 -122 371 -106
rect 455 34 489 50
rect 455 -122 489 -106
rect 573 34 607 50
rect 573 -122 607 -106
rect 687 -137 721 -121
<< viali >>
rect -548 111 -514 145
rect -430 111 -396 145
rect -312 111 -278 145
rect -194 111 -160 145
rect -76 111 -42 145
rect 42 111 76 145
rect 160 111 194 145
rect 278 111 312 145
rect 396 111 430 145
rect 514 111 548 145
rect -607 -106 -573 34
rect -489 -89 -455 17
rect -371 -106 -337 34
rect -253 -89 -219 17
rect -135 -106 -101 34
rect -17 -89 17 17
rect 101 -106 135 34
rect 219 -89 253 17
rect 337 -106 371 34
rect 455 -89 489 17
rect 573 -106 607 34
<< metal1 >>
rect -560 145 -502 151
rect -560 111 -548 145
rect -514 111 -502 145
rect -560 105 -502 111
rect -442 145 -384 151
rect -442 111 -430 145
rect -396 111 -384 145
rect -442 105 -384 111
rect -324 145 -266 151
rect -324 111 -312 145
rect -278 111 -266 145
rect -324 105 -266 111
rect -206 145 -148 151
rect -206 111 -194 145
rect -160 111 -148 145
rect -206 105 -148 111
rect -88 145 -30 151
rect -88 111 -76 145
rect -42 111 -30 145
rect -88 105 -30 111
rect 30 145 88 151
rect 30 111 42 145
rect 76 111 88 145
rect 30 105 88 111
rect 148 145 206 151
rect 148 111 160 145
rect 194 111 206 145
rect 148 105 206 111
rect 266 145 324 151
rect 266 111 278 145
rect 312 111 324 145
rect 266 105 324 111
rect 384 145 442 151
rect 384 111 396 145
rect 430 111 442 145
rect 384 105 442 111
rect 502 145 560 151
rect 502 111 514 145
rect 548 111 560 145
rect 502 105 560 111
rect -613 34 -567 46
rect -613 -106 -607 34
rect -573 -106 -567 34
rect -377 34 -331 46
rect -495 17 -449 29
rect -495 -89 -489 17
rect -455 -89 -449 17
rect -495 -101 -449 -89
rect -613 -118 -567 -106
rect -377 -106 -371 34
rect -337 -106 -331 34
rect -141 34 -95 46
rect -259 17 -213 29
rect -259 -89 -253 17
rect -219 -89 -213 17
rect -259 -101 -213 -89
rect -377 -118 -331 -106
rect -141 -106 -135 34
rect -101 -106 -95 34
rect 95 34 141 46
rect -23 17 23 29
rect -23 -89 -17 17
rect 17 -89 23 17
rect -23 -101 23 -89
rect -141 -118 -95 -106
rect 95 -106 101 34
rect 135 -106 141 34
rect 331 34 377 46
rect 213 17 259 29
rect 213 -89 219 17
rect 253 -89 259 17
rect 213 -101 259 -89
rect 95 -118 141 -106
rect 331 -106 337 34
rect 371 -106 377 34
rect 567 34 613 46
rect 449 17 495 29
rect 449 -89 455 17
rect 489 -89 495 17
rect 449 -101 495 -89
rect 331 -118 377 -106
rect 567 -106 573 34
rect 607 -106 613 34
rect 567 -118 613 -106
<< labels >>
flabel metal1 s -536 126 -532 128 0 FreeSans 480 0 0 0 G0
<< properties >>
string FIXED_BBOX -704 -231 704 231
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.3 m 1 nf 10 diffcov 80 polycov 80 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 80 rlcov 80 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 60 viadrn 80 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
