magic
tech sky130B
magscale 1 2
timestamp 1697762684
<< viali >>
rect 28221 2573 28261 2613
rect 28221 2474 28261 2514
rect 28223 2299 28263 2339
rect 28224 2200 28264 2240
rect 28227 2020 28267 2060
rect 28222 1925 28262 1965
rect 28227 1749 28267 1789
rect 28221 1649 28261 1689
rect 28222 1471 28262 1511
rect 28222 1374 28262 1414
rect 28221 1197 28261 1237
rect 28222 1100 28262 1140
rect 28228 919 28268 959
rect 28222 823 28262 863
rect 28225 649 28265 689
rect 28225 552 28265 592
rect 28227 372 28267 412
rect 28225 274 28265 314
<< metal1 >>
rect 27084 4168 27136 4174
rect 27084 4110 27136 4116
rect 27093 3572 27145 3578
rect 27093 3514 27145 3520
rect -195 3422 6538 3458
rect 636 2869 672 3422
rect 636 2833 778 2869
rect 2654 2836 2690 3422
rect 4578 2836 4614 3422
rect 6502 2836 6538 3422
rect 27076 2958 27128 2964
rect 27076 2900 27128 2906
rect 28215 2619 28267 2625
rect 28215 2561 28267 2567
rect 28215 2520 28267 2526
rect 28215 2462 28267 2468
rect 28217 2345 28269 2351
rect 28217 2287 28269 2293
rect 28218 2246 28270 2252
rect -232 2110 626 2204
rect 8228 2112 8230 2200
rect 28218 2188 28270 2194
rect 28221 2066 28273 2072
rect 28221 2008 28273 2014
rect 28216 1971 28268 1977
rect 28216 1913 28268 1919
rect 28221 1795 28273 1801
rect 28221 1737 28273 1743
rect 28215 1695 28267 1701
rect -280 1572 578 1666
rect 28215 1637 28267 1643
rect 28216 1517 28268 1523
rect 28216 1459 28268 1465
rect 28216 1420 28268 1426
rect 28216 1362 28268 1368
rect 28215 1243 28267 1249
rect 28215 1185 28267 1191
rect 28216 1146 28268 1152
rect 28216 1088 28268 1094
rect 28222 965 28274 971
rect 28222 907 28274 913
rect 28216 869 28268 875
rect 28216 811 28268 817
rect 28219 695 28271 701
rect 28219 637 28271 643
rect 28219 598 28271 604
rect 28219 540 28271 546
rect 28221 418 28273 424
rect 28221 360 28273 366
rect 28219 320 28271 326
rect 28219 262 28271 268
rect 27955 -20 28050 130
rect 28501 -22 28596 128
<< via1 >>
rect 27084 4116 27136 4168
rect 27093 3520 27145 3572
rect 27076 2906 27128 2958
rect 28215 2613 28267 2619
rect 28215 2573 28221 2613
rect 28221 2573 28261 2613
rect 28261 2573 28267 2613
rect 28215 2567 28267 2573
rect 28215 2514 28267 2520
rect 28215 2474 28221 2514
rect 28221 2474 28261 2514
rect 28261 2474 28267 2514
rect 28215 2468 28267 2474
rect 28217 2339 28269 2345
rect 28217 2299 28223 2339
rect 28223 2299 28263 2339
rect 28263 2299 28269 2339
rect 28217 2293 28269 2299
rect 28218 2240 28270 2246
rect 28218 2200 28224 2240
rect 28224 2200 28264 2240
rect 28264 2200 28270 2240
rect 28218 2194 28270 2200
rect 28221 2060 28273 2066
rect 28221 2020 28227 2060
rect 28227 2020 28267 2060
rect 28267 2020 28273 2060
rect 28221 2014 28273 2020
rect 28216 1965 28268 1971
rect 28216 1925 28222 1965
rect 28222 1925 28262 1965
rect 28262 1925 28268 1965
rect 28216 1919 28268 1925
rect 28221 1789 28273 1795
rect 28221 1749 28227 1789
rect 28227 1749 28267 1789
rect 28267 1749 28273 1789
rect 28221 1743 28273 1749
rect 28215 1689 28267 1695
rect 28215 1649 28221 1689
rect 28221 1649 28261 1689
rect 28261 1649 28267 1689
rect 28215 1643 28267 1649
rect 28216 1511 28268 1517
rect 28216 1471 28222 1511
rect 28222 1471 28262 1511
rect 28262 1471 28268 1511
rect 28216 1465 28268 1471
rect 28216 1414 28268 1420
rect 28216 1374 28222 1414
rect 28222 1374 28262 1414
rect 28262 1374 28268 1414
rect 28216 1368 28268 1374
rect 28215 1237 28267 1243
rect 28215 1197 28221 1237
rect 28221 1197 28261 1237
rect 28261 1197 28267 1237
rect 28215 1191 28267 1197
rect 28216 1140 28268 1146
rect 28216 1100 28222 1140
rect 28222 1100 28262 1140
rect 28262 1100 28268 1140
rect 28216 1094 28268 1100
rect 28222 959 28274 965
rect 28222 919 28228 959
rect 28228 919 28268 959
rect 28268 919 28274 959
rect 28222 913 28274 919
rect 28216 863 28268 869
rect 28216 823 28222 863
rect 28222 823 28262 863
rect 28262 823 28268 863
rect 28216 817 28268 823
rect 28219 689 28271 695
rect 28219 649 28225 689
rect 28225 649 28265 689
rect 28265 649 28271 689
rect 28219 643 28271 649
rect 28219 592 28271 598
rect 28219 552 28225 592
rect 28225 552 28265 592
rect 28265 552 28271 592
rect 28219 546 28271 552
rect 28221 412 28273 418
rect 28221 372 28227 412
rect 28227 372 28267 412
rect 28267 372 28273 412
rect 28221 366 28273 372
rect 28219 314 28271 320
rect 28219 274 28225 314
rect 28225 274 28265 314
rect 28265 274 28271 314
rect 28219 268 28271 274
<< metal2 >>
rect 27063 5326 27826 5377
rect 27081 4708 27728 4755
rect 27078 4116 27084 4168
rect 27136 4164 27142 4168
rect 27136 4120 27648 4164
rect 27136 4116 27142 4120
rect 3020 3666 3080 3675
rect 3020 3597 3080 3606
rect 3031 3515 3069 3597
rect 27087 3520 27093 3572
rect 27145 3571 27151 3572
rect 27145 3520 27576 3571
rect 2451 3477 8211 3515
rect 2451 2875 2489 3477
rect 2321 2837 2489 2875
rect 4361 2873 4399 3477
rect 6245 2875 6283 3477
rect 4243 2835 4399 2873
rect 6163 2837 6283 2875
rect 8173 2873 8211 3477
rect 27070 2906 27076 2958
rect 27128 2956 27134 2958
rect 27128 2908 27492 2956
rect 27128 2906 27134 2908
rect 8095 2835 8211 2873
rect 27104 2322 27396 2370
rect 27122 1734 27288 1782
rect -232 1504 7194 1545
rect 27093 690 27136 1137
rect 27240 963 27288 1734
rect 27348 1241 27396 2322
rect 27444 1515 27492 2908
rect 27525 1794 27576 3520
rect 27604 2062 27648 4120
rect 27681 2342 27728 4708
rect 27775 2618 27826 5326
rect 28209 2618 28215 2619
rect 27775 2567 28215 2618
rect 28267 2567 28273 2619
rect 28209 2468 28215 2520
rect 28267 2511 28273 2520
rect 28267 2477 28704 2511
rect 28267 2468 28273 2477
rect 28211 2342 28217 2345
rect 27681 2295 28217 2342
rect 28211 2293 28217 2295
rect 28269 2293 28275 2345
rect 28212 2194 28218 2246
rect 28270 2237 28276 2246
rect 28270 2203 28701 2237
rect 28270 2194 28276 2203
rect 28215 2062 28221 2066
rect 27604 2018 28221 2062
rect 28215 2014 28221 2018
rect 28273 2014 28279 2066
rect 28210 1919 28216 1971
rect 28268 1962 28274 1971
rect 28268 1928 28702 1962
rect 28268 1919 28274 1928
rect 28215 1794 28221 1795
rect 27525 1743 28221 1794
rect 28273 1743 28279 1795
rect 28209 1643 28215 1695
rect 28267 1686 28273 1695
rect 28267 1652 28704 1686
rect 28267 1643 28273 1652
rect 28210 1515 28216 1517
rect 27444 1467 28216 1515
rect 28210 1465 28216 1467
rect 28268 1465 28274 1517
rect 28210 1368 28216 1420
rect 28268 1411 28274 1420
rect 28268 1377 28705 1411
rect 28268 1368 28274 1377
rect 28209 1241 28215 1243
rect 27348 1193 28215 1241
rect 28209 1191 28215 1193
rect 28267 1191 28273 1243
rect 28210 1094 28216 1146
rect 28268 1137 28274 1146
rect 28268 1103 28702 1137
rect 28268 1094 28274 1103
rect 28216 963 28222 965
rect 27240 915 28222 963
rect 28216 913 28222 915
rect 28274 913 28280 965
rect 28210 817 28216 869
rect 28268 860 28274 869
rect 28268 826 28702 860
rect 28268 817 28274 826
rect 28213 690 28219 695
rect 27093 647 28219 690
rect 28213 643 28219 647
rect 28271 643 28277 695
rect 27097 413 27139 571
rect 28213 546 28219 598
rect 28271 589 28277 598
rect 28271 555 28704 589
rect 28271 546 28277 555
rect 28215 413 28221 418
rect 27097 371 28221 413
rect 28215 366 28221 371
rect 28273 366 28279 418
rect 28213 268 28219 320
rect 28271 311 28277 320
rect 28271 277 28704 311
rect 28271 268 28277 277
<< via2 >>
rect 3020 3606 3080 3666
<< metal3 >>
rect 2998 3671 3098 3686
rect 2998 3601 3015 3671
rect 3085 3601 3098 3671
rect 2998 3582 3098 3601
<< via3 >>
rect 3015 3666 3085 3671
rect 3015 3606 3020 3666
rect 3020 3606 3080 3666
rect 3080 3606 3085 3666
rect 3015 3601 3085 3606
<< metal4 >>
rect 3020 3672 3080 3794
rect 3014 3671 3086 3672
rect 3014 3601 3015 3671
rect 3085 3601 3086 3671
rect 3014 3600 3086 3601
use carray  carray_0
timestamp 1697663729
transform 1 0 -62 0 1 5400
box 62 -5400 27238 480
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1693170804
transform 0 1 28005 1 0 1899
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1693170804
transform 0 1 28005 1 0 2173
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_2
timestamp 1693170804
transform 0 1 28005 1 0 2448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_3
timestamp 1693170804
transform 0 1 28005 1 0 1349
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_4
timestamp 1693170804
transform 0 1 28005 1 0 798
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_5
timestamp 1693170804
transform 0 1 28005 1 0 1073
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_6
timestamp 1693170804
transform 0 1 28005 1 0 524
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_7
timestamp 1693170804
transform 0 1 28005 1 0 249
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_8
timestamp 1693170804
transform 0 1 28005 1 0 1624
box -38 -48 314 592
use sky130_fd_sc_hd__tap_2  sky130_fd_sc_hd__tap_2_0
timestamp 1693170804
transform 0 1 28005 -1 0 252
box -38 -48 222 592
use sky130_fd_sc_hd__tap_2  sky130_fd_sc_hd__tap_2_1
timestamp 1693170804
transform 0 1 28005 -1 0 2905
box -38 -48 222 592
use sky130_fd_sc_hd__tap_2  sky130_fd_sc_hd__tap_2_2
timestamp 1693170804
transform 1 0 428 0 1 1616
box -38 -48 222 592
use sky130_fd_sc_hd__tap_2  sky130_fd_sc_hd__tap_2_3
timestamp 1693170804
transform 1 0 8304 0 1 1616
box -38 -48 222 592
use sw_top  sw_top_0
timestamp 1697661741
transform 1 0 6753 0 1 2396
box -410 -892 1590 1027
use sw_top  sw_top_1
timestamp 1697661741
transform 1 0 4830 0 1 2396
box -410 -892 1590 1027
use sw_top  sw_top_2
timestamp 1697661741
transform 1 0 984 0 1 2396
box -410 -892 1590 1027
use sw_top  sw_top_3
timestamp 1697661741
transform 1 0 2907 0 1 2396
box -410 -892 1590 1027
<< labels >>
flabel metal2 -232 1504 -191 1545 0 FreeSans 800 0 0 0 sample
port 11 nsew
flabel metal2 2451 3477 8211 3515 0 FreeSans 1600 0 0 0 out
port 12 nsew
flabel metal1 s -232 2110 -138 2204 0 FreeSans 640 0 0 0 vdd
port 10 nsew
flabel metal1 -280 1572 578 1666 0 FreeSans 800 0 0 0 vss
port 13 nsew
flabel metal1 -185 3422 -149 3458 0 FreeSans 800 0 0 0 vin
port 9 nsew
flabel metal2 28271 277 28704 311 0 FreeSans 800 0 0 0 dum
port 8 nsew
flabel metal2 28271 555 28704 589 0 FreeSans 800 0 0 0 ctl0
port 0 nsew
flabel metal2 28268 826 28702 860 0 FreeSans 800 0 0 0 ctl1
port 1 nsew
flabel metal2 28268 1103 28702 1137 0 FreeSans 800 0 0 0 ctl2
port 2 nsew
flabel metal2 28268 1377 28705 1411 0 FreeSans 800 0 0 0 ctl3
port 3 nsew
flabel metal2 28267 1652 28704 1686 0 FreeSans 800 0 0 0 ctl4
port 4 nsew
flabel metal2 28268 1928 28702 1962 0 FreeSans 800 0 0 0 ctl5
port 5 nsew
flabel metal2 28270 2203 28701 2237 0 FreeSans 800 0 0 0 ctl6
port 6 nsew
flabel metal2 28267 2477 28704 2511 0 FreeSans 800 0 0 0 ctl7
port 7 nsew
flabel metal1 28501 -22 28596 128 0 FreeSans 800 0 0 0 vdd
port 10 nsew
flabel metal1 27955 -20 28050 130 0 FreeSans 800 0 0 0 vss
port 13 nsew
<< end >>
