magic
tech sky130B
magscale 1 2
timestamp 1694808442
<< viali >>
rect 1133 12937 1167 12971
rect 3157 12937 3191 12971
rect 5549 12937 5583 12971
rect 7113 12937 7147 12971
rect 8861 12937 8895 12971
rect 10793 12937 10827 12971
rect 12817 12937 12851 12971
rect 14657 12937 14691 12971
rect 15393 12937 15427 12971
rect 1685 12869 1719 12903
rect 1869 12733 1903 12767
rect 3341 12733 3375 12767
rect 3433 12733 3467 12767
rect 3617 12733 3651 12767
rect 6193 12733 6227 12767
rect 9045 12733 9079 12767
rect 10977 12733 11011 12767
rect 12633 12733 12667 12767
rect 14473 12733 14507 12767
rect 397 12665 431 12699
rect 765 12665 799 12699
rect 1409 12665 1443 12699
rect 5457 12665 5491 12699
rect 7021 12665 7055 12699
rect 15117 12665 15151 12699
rect 3525 12597 3559 12631
rect 6377 12597 6411 12631
rect 5825 12393 5859 12427
rect 14841 12393 14875 12427
rect 2973 12325 3007 12359
rect 3709 12325 3743 12359
rect 5641 12325 5675 12359
rect 6193 12325 6227 12359
rect 6653 12325 6687 12359
rect 581 12257 615 12291
rect 2789 12257 2823 12291
rect 5457 12257 5491 12291
rect 6101 12257 6135 12291
rect 6285 12257 6319 12291
rect 14933 12257 14967 12291
rect 15117 12257 15151 12291
rect 857 12189 891 12223
rect 3433 12189 3467 12223
rect 5181 12189 5215 12223
rect 6377 12189 6411 12223
rect 2329 12053 2363 12087
rect 3157 12053 3191 12087
rect 8125 12053 8159 12087
rect 15393 12053 15427 12087
rect 1225 11849 1259 11883
rect 3341 11849 3375 11883
rect 6193 11849 6227 11883
rect 1409 11781 1443 11815
rect 4353 11781 4387 11815
rect 673 11645 707 11679
rect 1041 11645 1075 11679
rect 1225 11645 1259 11679
rect 1685 11645 1719 11679
rect 3341 11645 3375 11679
rect 3525 11645 3559 11679
rect 3617 11645 3651 11679
rect 4169 11645 4203 11679
rect 4813 11645 4847 11679
rect 5917 11645 5951 11679
rect 6009 11645 6043 11679
rect 6745 11645 6779 11679
rect 8401 11645 8435 11679
rect 8769 11645 8803 11679
rect 1409 11577 1443 11611
rect 6193 11577 6227 11611
rect 8033 11577 8067 11611
rect 8217 11577 8251 11611
rect 489 11509 523 11543
rect 1593 11509 1627 11543
rect 4905 11509 4939 11543
rect 6837 11509 6871 11543
rect 8953 11509 8987 11543
rect 2329 11305 2363 11339
rect 5181 11305 5215 11339
rect 6469 11305 6503 11339
rect 8493 11305 8527 11339
rect 14841 11305 14875 11339
rect 3065 11237 3099 11271
rect 6101 11237 6135 11271
rect 6193 11237 6227 11271
rect 7021 11237 7055 11271
rect 581 11169 615 11203
rect 2697 11169 2731 11203
rect 2789 11169 2823 11203
rect 2973 11169 3007 11203
rect 3157 11169 3191 11203
rect 5917 11169 5951 11203
rect 6285 11169 6319 11203
rect 14933 11169 14967 11203
rect 15117 11169 15151 11203
rect 857 11101 891 11135
rect 3433 11101 3467 11135
rect 3709 11101 3743 11135
rect 6745 11101 6779 11135
rect 3341 11033 3375 11067
rect 15393 11033 15427 11067
rect 2605 10965 2639 10999
rect 1409 10761 1443 10795
rect 15117 10761 15151 10795
rect 11989 10693 12023 10727
rect 7941 10625 7975 10659
rect 673 10557 707 10591
rect 1593 10557 1627 10591
rect 1777 10557 1811 10591
rect 1869 10557 1903 10591
rect 6101 10557 6135 10591
rect 6469 10557 6503 10591
rect 9873 10557 9907 10591
rect 11805 10557 11839 10591
rect 12357 10557 12391 10591
rect 15025 10557 15059 10591
rect 6285 10489 6319 10523
rect 6377 10489 6411 10523
rect 8217 10489 8251 10523
rect 489 10421 523 10455
rect 6653 10421 6687 10455
rect 9689 10421 9723 10455
rect 10057 10421 10091 10455
rect 12449 10421 12483 10455
rect 6186 10217 6220 10251
rect 9321 10217 9355 10251
rect 3065 10149 3099 10183
rect 4905 10149 4939 10183
rect 6101 10149 6135 10183
rect 9137 10149 9171 10183
rect 2329 10081 2363 10115
rect 2513 10081 2547 10115
rect 4813 10081 4847 10115
rect 4997 10081 5031 10115
rect 5181 10081 5215 10115
rect 5733 10081 5767 10115
rect 5917 10081 5951 10115
rect 6009 10081 6043 10115
rect 6285 10081 6319 10115
rect 6469 10081 6503 10115
rect 8953 10081 8987 10115
rect 15117 10081 15151 10115
rect 397 10013 431 10047
rect 673 10013 707 10047
rect 2145 10013 2179 10047
rect 2789 10013 2823 10047
rect 6745 10013 6779 10047
rect 2697 9877 2731 9911
rect 4537 9877 4571 9911
rect 4629 9877 4663 9911
rect 5917 9877 5951 9911
rect 8217 9877 8251 9911
rect 15393 9877 15427 9911
rect 1133 9673 1167 9707
rect 1593 9605 1627 9639
rect 15025 9605 15059 9639
rect 4445 9537 4479 9571
rect 4721 9537 4755 9571
rect 6193 9537 6227 9571
rect 8217 9537 8251 9571
rect 10241 9537 10275 9571
rect 14289 9537 14323 9571
rect 14749 9537 14783 9571
rect 14933 9537 14967 9571
rect 673 9469 707 9503
rect 949 9469 983 9503
rect 1133 9469 1167 9503
rect 1869 9469 1903 9503
rect 2973 9469 3007 9503
rect 3341 9469 3375 9503
rect 10609 9469 10643 9503
rect 14657 9469 14691 9503
rect 1593 9401 1627 9435
rect 1777 9401 1811 9435
rect 3065 9401 3099 9435
rect 3157 9401 3191 9435
rect 8493 9401 8527 9435
rect 15393 9401 15427 9435
rect 489 9333 523 9367
rect 2789 9333 2823 9367
rect 9965 9333 9999 9367
rect 12035 9333 12069 9367
rect 2789 9129 2823 9163
rect 5457 9129 5491 9163
rect 6745 9129 6779 9163
rect 8769 9129 8803 9163
rect 9505 9129 9539 9163
rect 10701 9129 10735 9163
rect 3985 9061 4019 9095
rect 765 8993 799 9027
rect 2605 8993 2639 9027
rect 2881 8993 2915 9027
rect 3801 8993 3835 9027
rect 4169 8993 4203 9027
rect 5733 8993 5767 9027
rect 6929 8993 6963 9027
rect 8861 8993 8895 9027
rect 9597 8993 9631 9027
rect 10885 8993 10919 9027
rect 11437 8993 11471 9027
rect 11989 8993 12023 9027
rect 13921 8993 13955 9027
rect 14381 8993 14415 9027
rect 14565 8993 14599 9027
rect 14657 8993 14691 9027
rect 15117 8993 15151 9027
rect 1041 8925 1075 8959
rect 11529 8925 11563 8959
rect 11621 8925 11655 8959
rect 12357 8925 12391 8959
rect 11069 8857 11103 8891
rect 2513 8789 2547 8823
rect 2605 8789 2639 8823
rect 13783 8789 13817 8823
rect 14105 8789 14139 8823
rect 14197 8789 14231 8823
rect 15393 8789 15427 8823
rect 1317 8585 1351 8619
rect 5365 8585 5399 8619
rect 9781 8585 9815 8619
rect 13093 8585 13127 8619
rect 14565 8585 14599 8619
rect 3525 8517 3559 8551
rect 6009 8517 6043 8551
rect 14749 8517 14783 8551
rect 3893 8449 3927 8483
rect 5733 8449 5767 8483
rect 6561 8449 6595 8483
rect 8401 8449 8435 8483
rect 13553 8449 13587 8483
rect 765 8381 799 8415
rect 1133 8381 1167 8415
rect 1317 8381 1351 8415
rect 2973 8381 3007 8415
rect 3157 8381 3191 8415
rect 3249 8381 3283 8415
rect 3341 8381 3375 8415
rect 3617 8381 3651 8415
rect 5917 8381 5951 8415
rect 6377 8381 6411 8415
rect 7021 8381 7055 8415
rect 8217 8381 8251 8415
rect 8493 8381 8527 8415
rect 9597 8381 9631 8415
rect 9689 8381 9723 8415
rect 13277 8381 13311 8415
rect 13369 8381 13403 8415
rect 13645 8381 13679 8415
rect 14197 8381 14231 8415
rect 14933 8381 14967 8415
rect 15117 8381 15151 8415
rect 397 8313 431 8347
rect 2053 8313 2087 8347
rect 2237 8313 2271 8347
rect 2421 8313 2455 8347
rect 6469 8313 6503 8347
rect 9873 8313 9907 8347
rect 14381 8313 14415 8347
rect 6837 8245 6871 8279
rect 8033 8245 8067 8279
rect 3065 8041 3099 8075
rect 8585 8041 8619 8075
rect 9413 8041 9447 8075
rect 9581 8041 9615 8075
rect 10057 8041 10091 8075
rect 15301 8041 15335 8075
rect 1041 7973 1075 8007
rect 1225 7973 1259 8007
rect 2421 7973 2455 8007
rect 5733 7973 5767 8007
rect 7113 7973 7147 8007
rect 9781 7973 9815 8007
rect 673 7905 707 7939
rect 765 7905 799 7939
rect 949 7905 983 7939
rect 1317 7905 1351 7939
rect 1409 7905 1443 7939
rect 1777 7905 1811 7939
rect 2145 7905 2179 7939
rect 2329 7905 2363 7939
rect 2513 7905 2547 7939
rect 4537 7905 4571 7939
rect 4813 7905 4847 7939
rect 6285 7905 6319 7939
rect 6837 7905 6871 7939
rect 8677 7905 8711 7939
rect 8861 7905 8895 7939
rect 9873 7905 9907 7939
rect 10149 7905 10183 7939
rect 10793 7905 10827 7939
rect 10977 7905 11011 7939
rect 11897 7905 11931 7939
rect 14657 7905 14691 7939
rect 15393 7905 15427 7939
rect 12265 7837 12299 7871
rect 14749 7837 14783 7871
rect 1041 7769 1075 7803
rect 9873 7769 9907 7803
rect 13691 7769 13725 7803
rect 489 7701 523 7735
rect 765 7701 799 7735
rect 2697 7701 2731 7735
rect 4629 7701 4663 7735
rect 8769 7701 8803 7735
rect 9597 7701 9631 7735
rect 10885 7701 10919 7735
rect 14381 7701 14415 7735
rect 2145 7497 2179 7531
rect 3046 7497 3080 7531
rect 5181 7497 5215 7531
rect 13093 7497 13127 7531
rect 15301 7497 15335 7531
rect 5641 7429 5675 7463
rect 14013 7429 14047 7463
rect 673 7361 707 7395
rect 2789 7361 2823 7395
rect 6009 7361 6043 7395
rect 12081 7361 12115 7395
rect 13553 7361 13587 7395
rect 14197 7361 14231 7395
rect 15117 7361 15151 7395
rect 397 7293 431 7327
rect 4997 7293 5031 7327
rect 5457 7293 5491 7327
rect 5641 7293 5675 7327
rect 13277 7293 13311 7327
rect 13369 7293 13403 7327
rect 13645 7293 13679 7327
rect 13737 7293 13771 7327
rect 13921 7293 13955 7327
rect 14289 7293 14323 7327
rect 14933 7293 14967 7327
rect 15209 7293 15243 7327
rect 15393 7293 15427 7327
rect 6285 7225 6319 7259
rect 7941 7225 7975 7259
rect 11805 7225 11839 7259
rect 14749 7225 14783 7259
rect 4537 7157 4571 7191
rect 7757 7157 7791 7191
rect 9229 7157 9263 7191
rect 10333 7157 10367 7191
rect 13921 7157 13955 7191
rect 14657 7157 14691 7191
rect 6469 6953 6503 6987
rect 9781 6953 9815 6987
rect 9873 6953 9907 6987
rect 8585 6885 8619 6919
rect 673 6817 707 6851
rect 1685 6817 1719 6851
rect 4169 6817 4203 6851
rect 6653 6817 6687 6851
rect 7665 6817 7699 6851
rect 7849 6817 7883 6851
rect 8677 6817 8711 6851
rect 9045 6817 9079 6851
rect 9321 6817 9355 6851
rect 10977 6817 11011 6851
rect 11161 6817 11195 6851
rect 11345 6817 11379 6851
rect 15301 6817 15335 6851
rect 8033 6749 8067 6783
rect 8309 6749 8343 6783
rect 10057 6749 10091 6783
rect 489 6613 523 6647
rect 1501 6613 1535 6647
rect 4353 6613 4387 6647
rect 9413 6613 9447 6647
rect 15485 6613 15519 6647
rect 2237 6409 2271 6443
rect 4077 6409 4111 6443
rect 4518 6409 4552 6443
rect 6285 6409 6319 6443
rect 8769 6409 8803 6443
rect 12725 6409 12759 6443
rect 15209 6409 15243 6443
rect 6009 6341 6043 6375
rect 13645 6341 13679 6375
rect 14657 6341 14691 6375
rect 397 6273 431 6307
rect 2145 6273 2179 6307
rect 4261 6273 4295 6307
rect 8953 6273 8987 6307
rect 9045 6273 9079 6307
rect 9137 6273 9171 6307
rect 10977 6273 11011 6307
rect 13369 6273 13403 6307
rect 14013 6273 14047 6307
rect 2605 6205 2639 6239
rect 3433 6205 3467 6239
rect 3617 6205 3651 6239
rect 6101 6205 6135 6239
rect 6285 6205 6319 6239
rect 9229 6205 9263 6239
rect 9413 6205 9447 6239
rect 9597 6205 9631 6239
rect 9781 6205 9815 6239
rect 9965 6205 9999 6239
rect 13277 6205 13311 6239
rect 14105 6205 14139 6239
rect 15025 6205 15059 6239
rect 673 6137 707 6171
rect 2421 6137 2455 6171
rect 3709 6137 3743 6171
rect 3893 6137 3927 6171
rect 10517 6137 10551 6171
rect 11253 6137 11287 6171
rect 14381 6137 14415 6171
rect 3525 6069 3559 6103
rect 13737 6069 13771 6103
rect 14841 6069 14875 6103
rect 1133 5865 1167 5899
rect 1507 5865 1541 5899
rect 1593 5865 1627 5899
rect 3249 5865 3283 5899
rect 5917 5865 5951 5899
rect 14841 5865 14875 5899
rect 1409 5797 1443 5831
rect 8217 5797 8251 5831
rect 9965 5797 9999 5831
rect 765 5729 799 5763
rect 1041 5729 1075 5763
rect 1225 5729 1259 5763
rect 1685 5729 1719 5763
rect 4537 5729 4571 5763
rect 4629 5729 4663 5763
rect 4813 5729 4847 5763
rect 4997 5729 5031 5763
rect 5549 5729 5583 5763
rect 5703 5729 5737 5763
rect 7389 5729 7423 5763
rect 7665 5729 7699 5763
rect 7849 5729 7883 5763
rect 10057 5729 10091 5763
rect 10149 5729 10183 5763
rect 10333 5729 10367 5763
rect 10701 5729 10735 5763
rect 10885 5729 10919 5763
rect 10977 5729 11011 5763
rect 11069 5729 11103 5763
rect 11345 5729 11379 5763
rect 11529 5729 11563 5763
rect 14933 5729 14967 5763
rect 15117 5729 15151 5763
rect 7205 5593 7239 5627
rect 11253 5593 11287 5627
rect 489 5525 523 5559
rect 4813 5525 4847 5559
rect 5089 5525 5123 5559
rect 10333 5525 10367 5559
rect 11345 5525 11379 5559
rect 15393 5525 15427 5559
rect 3801 5321 3835 5355
rect 5181 5321 5215 5355
rect 7757 5253 7791 5287
rect 9873 5253 9907 5287
rect 10241 5253 10275 5287
rect 4813 5185 4847 5219
rect 10057 5185 10091 5219
rect 3341 5117 3375 5151
rect 3433 5117 3467 5151
rect 3525 5117 3559 5151
rect 3617 5117 3651 5151
rect 4537 5117 4571 5151
rect 4721 5117 4755 5151
rect 4997 5117 5031 5151
rect 5273 5117 5307 5151
rect 5641 5117 5675 5151
rect 5733 5117 5767 5151
rect 6101 5117 6135 5151
rect 6469 5117 6503 5151
rect 6837 5117 6871 5151
rect 7113 5117 7147 5151
rect 7321 5117 7355 5151
rect 7481 5117 7515 5151
rect 7573 5117 7607 5151
rect 8217 5117 8251 5151
rect 8309 5117 8343 5151
rect 8402 5117 8436 5151
rect 8585 5117 8619 5151
rect 8677 5117 8711 5151
rect 8774 5117 8808 5151
rect 9045 5117 9079 5151
rect 9229 5117 9263 5151
rect 9597 5117 9631 5151
rect 9781 5117 9815 5151
rect 10333 5117 10367 5151
rect 11161 5117 11195 5151
rect 12725 5117 12759 5151
rect 13093 5117 13127 5151
rect 3985 5049 4019 5083
rect 4077 5049 4111 5083
rect 5457 5049 5491 5083
rect 5825 5049 5859 5083
rect 13369 5049 13403 5083
rect 14933 5049 14967 5083
rect 15117 5049 15151 5083
rect 4169 4981 4203 5015
rect 6009 4981 6043 5015
rect 7021 4981 7055 5015
rect 7389 4981 7423 5015
rect 8125 4981 8159 5015
rect 8953 4981 8987 5015
rect 9045 4981 9079 5015
rect 10057 4981 10091 5015
rect 10977 4981 11011 5015
rect 12909 4981 12943 5015
rect 14841 4981 14875 5015
rect 15301 4981 15335 5015
rect 6193 4777 6227 4811
rect 7481 4777 7515 4811
rect 7665 4777 7699 4811
rect 13001 4777 13035 4811
rect 14013 4777 14047 4811
rect 14841 4777 14875 4811
rect 5181 4709 5215 4743
rect 9045 4709 9079 4743
rect 10241 4709 10275 4743
rect 397 4641 431 4675
rect 2789 4641 2823 4675
rect 3065 4641 3099 4675
rect 3249 4641 3283 4675
rect 3709 4641 3743 4675
rect 5457 4641 5491 4675
rect 5641 4641 5675 4675
rect 5825 4641 5859 4675
rect 6101 4641 6135 4675
rect 6285 4641 6319 4675
rect 6653 4641 6687 4675
rect 6929 4641 6963 4675
rect 7021 4641 7055 4675
rect 8309 4641 8343 4675
rect 8493 4641 8527 4675
rect 9229 4641 9263 4675
rect 9505 4641 9539 4675
rect 9965 4641 9999 4675
rect 13185 4641 13219 4675
rect 13829 4641 13863 4675
rect 14105 4641 14139 4675
rect 14657 4641 14691 4675
rect 15393 4641 15427 4675
rect 673 4573 707 4607
rect 3801 4573 3835 4607
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 5365 4573 5399 4607
rect 11069 4573 11103 4607
rect 11345 4573 11379 4607
rect 13369 4573 13403 4607
rect 13645 4573 13679 4607
rect 3065 4505 3099 4539
rect 5043 4505 5077 4539
rect 7205 4505 7239 4539
rect 8033 4505 8067 4539
rect 2145 4437 2179 4471
rect 3341 4437 3375 4471
rect 4537 4437 4571 4471
rect 4905 4437 4939 4471
rect 6469 4437 6503 4471
rect 6837 4437 6871 4471
rect 7673 4437 7707 4471
rect 8401 4437 8435 4471
rect 9413 4437 9447 4471
rect 12817 4437 12851 4471
rect 15301 4437 15335 4471
rect 1409 4233 1443 4267
rect 6837 4233 6871 4267
rect 11529 4233 11563 4267
rect 8217 4165 8251 4199
rect 10517 4165 10551 4199
rect 5917 4097 5951 4131
rect 6469 4097 6503 4131
rect 6929 4097 6963 4131
rect 13829 4097 13863 4131
rect 857 4029 891 4063
rect 1041 4029 1075 4063
rect 1133 4029 1167 4063
rect 1225 4029 1259 4063
rect 2421 4029 2455 4063
rect 3709 4029 3743 4063
rect 4261 4029 4295 4063
rect 4629 4029 4663 4063
rect 4721 4029 4755 4063
rect 4813 4029 4847 4063
rect 4997 4029 5031 4063
rect 5457 4029 5491 4063
rect 5641 4029 5675 4063
rect 6101 4029 6135 4063
rect 6193 4029 6227 4063
rect 6653 4029 6687 4063
rect 7021 4029 7055 4063
rect 7297 4029 7331 4063
rect 9413 4029 9447 4063
rect 9597 4029 9631 4063
rect 9689 4029 9723 4063
rect 10333 4029 10367 4063
rect 10977 4029 11011 4063
rect 11253 4029 11287 4063
rect 11345 4029 11379 4063
rect 13645 4029 13679 4063
rect 14473 4029 14507 4063
rect 15117 4029 15151 4063
rect 15393 4029 15427 4063
rect 5181 3961 5215 3995
rect 7481 3961 7515 3995
rect 8033 3961 8067 3995
rect 8953 3961 8987 3995
rect 10149 3961 10183 3995
rect 11161 3961 11195 3995
rect 2237 3893 2271 3927
rect 4445 3893 4479 3927
rect 5273 3893 5307 3927
rect 5549 3893 5583 3927
rect 7113 3893 7147 3927
rect 13461 3893 13495 3927
rect 14289 3893 14323 3927
rect 14933 3893 14967 3927
rect 15301 3893 15335 3927
rect 489 3689 523 3723
rect 949 3689 983 3723
rect 7665 3689 7699 3723
rect 10333 3689 10367 3723
rect 11253 3689 11287 3723
rect 15485 3689 15519 3723
rect 765 3621 799 3655
rect 2145 3621 2179 3655
rect 4721 3621 4755 3655
rect 7087 3621 7121 3655
rect 8125 3621 8159 3655
rect 10885 3621 10919 3655
rect 10977 3621 11011 3655
rect 11621 3621 11655 3655
rect 1133 3553 1167 3587
rect 1869 3553 1903 3587
rect 4537 3553 4571 3587
rect 7205 3553 7239 3587
rect 7297 3553 7331 3587
rect 7389 3553 7423 3587
rect 10701 3553 10735 3587
rect 11069 3553 11103 3587
rect 13185 3553 13219 3587
rect 15301 3553 15335 3587
rect 3617 3485 3651 3519
rect 4905 3485 4939 3519
rect 6929 3485 6963 3519
rect 8585 3485 8619 3519
rect 8861 3485 8895 3519
rect 11345 3485 11379 3519
rect 13461 3485 13495 3519
rect 13737 3485 13771 3519
rect 7757 3417 7791 3451
rect 13369 3417 13403 3451
rect 7573 3349 7607 3383
rect 13093 3349 13127 3383
rect 15209 3349 15243 3383
rect 581 3145 615 3179
rect 3525 3145 3559 3179
rect 4997 3145 5031 3179
rect 5181 3145 5215 3179
rect 9505 3145 9539 3179
rect 10241 3145 10275 3179
rect 13829 3145 13863 3179
rect 14933 3145 14967 3179
rect 15393 3145 15427 3179
rect 10609 3077 10643 3111
rect 6009 3009 6043 3043
rect 397 2941 431 2975
rect 3341 2941 3375 2975
rect 3893 2941 3927 2975
rect 4629 2941 4663 2975
rect 6285 2941 6319 2975
rect 8217 2941 8251 2975
rect 10793 2941 10827 2975
rect 11069 2941 11103 2975
rect 11437 2941 11471 2975
rect 14013 2941 14047 2975
rect 14289 2941 14323 2975
rect 14749 2941 14783 2975
rect 15117 2941 15151 2975
rect 4445 2873 4479 2907
rect 5006 2873 5040 2907
rect 10149 2873 10183 2907
rect 11253 2873 11287 2907
rect 11345 2873 11379 2907
rect 14565 2873 14599 2907
rect 11621 2805 11655 2839
rect 14197 2805 14231 2839
rect 3893 2601 3927 2635
rect 6653 2601 6687 2635
rect 10241 2601 10275 2635
rect 13185 2601 13219 2635
rect 2421 2533 2455 2567
rect 10885 2533 10919 2567
rect 11713 2533 11747 2567
rect 14565 2533 14599 2567
rect 15117 2533 15151 2567
rect 8401 2465 8435 2499
rect 8493 2465 8527 2499
rect 10701 2465 10735 2499
rect 10793 2465 10827 2499
rect 11069 2465 11103 2499
rect 11437 2465 11471 2499
rect 13553 2465 13587 2499
rect 14473 2465 14507 2499
rect 14749 2465 14783 2499
rect 2145 2397 2179 2431
rect 8125 2397 8159 2431
rect 8769 2397 8803 2431
rect 10517 2329 10551 2363
rect 13369 2261 13403 2295
rect 14289 2261 14323 2295
rect 14933 2261 14967 2295
rect 15393 2261 15427 2295
rect 13645 2057 13679 2091
rect 15209 2057 15243 2091
rect 6193 1989 6227 2023
rect 4445 1921 4479 1955
rect 4721 1921 4755 1955
rect 9597 1921 9631 1955
rect 13277 1921 13311 1955
rect 13461 1853 13495 1887
rect 13829 1853 13863 1887
rect 14013 1853 14047 1887
rect 14289 1853 14323 1887
rect 14381 1853 14415 1887
rect 15025 1853 15059 1887
rect 9873 1785 9907 1819
rect 11345 1717 11379 1751
rect 14197 1717 14231 1751
rect 14473 1717 14507 1751
rect 10149 1513 10183 1547
rect 10885 1513 10919 1547
rect 14841 1513 14875 1547
rect 11437 1445 11471 1479
rect 13369 1445 13403 1479
rect 15117 1445 15151 1479
rect 1409 1377 1443 1411
rect 3157 1377 3191 1411
rect 8769 1377 8803 1411
rect 9873 1377 9907 1411
rect 10057 1377 10091 1411
rect 10333 1377 10367 1411
rect 10701 1377 10735 1411
rect 10977 1377 11011 1411
rect 11253 1377 11287 1411
rect 9689 1309 9723 1343
rect 10517 1309 10551 1343
rect 13093 1309 13127 1343
rect 1317 1173 1351 1207
rect 3065 1173 3099 1207
rect 8677 1173 8711 1207
rect 11621 1173 11655 1207
rect 15393 1173 15427 1207
rect 581 969 615 1003
rect 15117 969 15151 1003
rect 397 765 431 799
rect 1501 765 1535 799
rect 3065 765 3099 799
rect 5457 765 5491 799
rect 7021 765 7055 799
rect 8769 765 8803 799
rect 10977 765 11011 799
rect 11069 765 11103 799
rect 12633 765 12667 799
rect 14473 765 14507 799
rect 14933 765 14967 799
rect 11161 697 11195 731
rect 1317 629 1351 663
rect 3249 629 3283 663
rect 5549 629 5583 663
rect 7113 629 7147 663
rect 8953 629 8987 663
rect 10793 629 10827 663
rect 12817 629 12851 663
rect 14657 629 14691 663
<< metal1 >>
rect 92 13082 15824 13104
rect 92 13030 1904 13082
rect 1956 13030 1968 13082
rect 2020 13030 2032 13082
rect 2084 13030 2096 13082
rect 2148 13030 2160 13082
rect 2212 13030 5837 13082
rect 5889 13030 5901 13082
rect 5953 13030 5965 13082
rect 6017 13030 6029 13082
rect 6081 13030 6093 13082
rect 6145 13030 9770 13082
rect 9822 13030 9834 13082
rect 9886 13030 9898 13082
rect 9950 13030 9962 13082
rect 10014 13030 10026 13082
rect 10078 13030 13703 13082
rect 13755 13030 13767 13082
rect 13819 13030 13831 13082
rect 13883 13030 13895 13082
rect 13947 13030 13959 13082
rect 14011 13030 15824 13082
rect 92 13008 15824 13030
rect 842 12928 848 12980
rect 900 12928 906 12980
rect 1118 12928 1124 12980
rect 1176 12928 1182 12980
rect 3145 12971 3203 12977
rect 3145 12937 3157 12971
rect 3191 12968 3203 12971
rect 3234 12968 3240 12980
rect 3191 12940 3240 12968
rect 3191 12937 3203 12940
rect 3145 12931 3203 12937
rect 3234 12928 3240 12940
rect 3292 12928 3298 12980
rect 5258 12928 5264 12980
rect 5316 12968 5322 12980
rect 5537 12971 5595 12977
rect 5537 12968 5549 12971
rect 5316 12940 5549 12968
rect 5316 12928 5322 12940
rect 5537 12937 5549 12940
rect 5583 12937 5595 12971
rect 5537 12931 5595 12937
rect 6638 12928 6644 12980
rect 6696 12968 6702 12980
rect 7101 12971 7159 12977
rect 7101 12968 7113 12971
rect 6696 12940 7113 12968
rect 6696 12928 6702 12940
rect 7101 12937 7113 12940
rect 7147 12937 7159 12971
rect 7101 12931 7159 12937
rect 8849 12971 8907 12977
rect 8849 12937 8861 12971
rect 8895 12968 8907 12971
rect 8938 12968 8944 12980
rect 8895 12940 8944 12968
rect 8895 12937 8907 12940
rect 8849 12931 8907 12937
rect 8938 12928 8944 12940
rect 8996 12928 9002 12980
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12968 10839 12971
rect 10870 12968 10876 12980
rect 10827 12940 10876 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 12802 12928 12808 12980
rect 12860 12928 12866 12980
rect 14642 12928 14648 12980
rect 14700 12928 14706 12980
rect 15381 12971 15439 12977
rect 15381 12937 15393 12971
rect 15427 12968 15439 12971
rect 15470 12968 15476 12980
rect 15427 12940 15476 12968
rect 15427 12937 15439 12940
rect 15381 12931 15439 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 860 12900 888 12928
rect 1673 12903 1731 12909
rect 1673 12900 1685 12903
rect 860 12872 1685 12900
rect 1673 12869 1685 12872
rect 1719 12869 1731 12903
rect 1673 12863 1731 12869
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12764 1915 12767
rect 2314 12764 2320 12776
rect 1903 12736 2320 12764
rect 1903 12733 1915 12736
rect 1857 12727 1915 12733
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 3234 12724 3240 12776
rect 3292 12764 3298 12776
rect 3329 12767 3387 12773
rect 3329 12764 3341 12767
rect 3292 12736 3341 12764
rect 3292 12724 3298 12736
rect 3329 12733 3341 12736
rect 3375 12733 3387 12767
rect 3329 12727 3387 12733
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12733 3479 12767
rect 3421 12727 3479 12733
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 382 12656 388 12708
rect 440 12656 446 12708
rect 753 12699 811 12705
rect 753 12665 765 12699
rect 799 12696 811 12699
rect 1302 12696 1308 12708
rect 799 12668 1308 12696
rect 799 12665 811 12668
rect 753 12659 811 12665
rect 1302 12656 1308 12668
rect 1360 12656 1366 12708
rect 1394 12656 1400 12708
rect 1452 12656 1458 12708
rect 3436 12696 3464 12727
rect 3344 12668 3464 12696
rect 3344 12640 3372 12668
rect 3326 12588 3332 12640
rect 3384 12588 3390 12640
rect 3510 12588 3516 12640
rect 3568 12588 3574 12640
rect 3620 12628 3648 12727
rect 5810 12724 5816 12776
rect 5868 12764 5874 12776
rect 6181 12767 6239 12773
rect 6181 12764 6193 12767
rect 5868 12736 6193 12764
rect 5868 12724 5874 12736
rect 6181 12733 6193 12736
rect 6227 12733 6239 12767
rect 6181 12727 6239 12733
rect 9030 12724 9036 12776
rect 9088 12724 9094 12776
rect 10962 12724 10968 12776
rect 11020 12724 11026 12776
rect 12342 12724 12348 12776
rect 12400 12764 12406 12776
rect 12621 12767 12679 12773
rect 12621 12764 12633 12767
rect 12400 12736 12633 12764
rect 12400 12724 12406 12736
rect 12621 12733 12633 12736
rect 12667 12733 12679 12767
rect 12621 12727 12679 12733
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14461 12767 14519 12773
rect 14461 12764 14473 12767
rect 14148 12736 14473 12764
rect 14148 12724 14154 12736
rect 14461 12733 14473 12736
rect 14507 12733 14519 12767
rect 14461 12727 14519 12733
rect 5442 12656 5448 12708
rect 5500 12656 5506 12708
rect 7009 12699 7067 12705
rect 7009 12696 7021 12699
rect 6886 12668 7021 12696
rect 6886 12640 6914 12668
rect 7009 12665 7021 12668
rect 7055 12665 7067 12699
rect 7009 12659 7067 12665
rect 15102 12656 15108 12708
rect 15160 12656 15166 12708
rect 5534 12628 5540 12640
rect 3620 12600 5540 12628
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 6365 12631 6423 12637
rect 6365 12597 6377 12631
rect 6411 12628 6423 12631
rect 6822 12628 6828 12640
rect 6411 12600 6828 12628
rect 6411 12597 6423 12600
rect 6365 12591 6423 12597
rect 6822 12588 6828 12600
rect 6880 12600 6914 12640
rect 6880 12588 6886 12600
rect 92 12538 15824 12560
rect 92 12486 2564 12538
rect 2616 12486 2628 12538
rect 2680 12486 2692 12538
rect 2744 12486 2756 12538
rect 2808 12486 2820 12538
rect 2872 12486 6497 12538
rect 6549 12486 6561 12538
rect 6613 12486 6625 12538
rect 6677 12486 6689 12538
rect 6741 12486 6753 12538
rect 6805 12486 10430 12538
rect 10482 12486 10494 12538
rect 10546 12486 10558 12538
rect 10610 12486 10622 12538
rect 10674 12486 10686 12538
rect 10738 12486 14363 12538
rect 14415 12486 14427 12538
rect 14479 12486 14491 12538
rect 14543 12486 14555 12538
rect 14607 12486 14619 12538
rect 14671 12486 15824 12538
rect 92 12464 15824 12486
rect 3050 12384 3056 12436
rect 3108 12424 3114 12436
rect 3108 12396 5212 12424
rect 3108 12384 3114 12396
rect 750 12356 756 12368
rect 584 12328 756 12356
rect 584 12297 612 12328
rect 750 12316 756 12328
rect 808 12316 814 12368
rect 1486 12316 1492 12368
rect 1544 12316 1550 12368
rect 2406 12316 2412 12368
rect 2464 12356 2470 12368
rect 2961 12359 3019 12365
rect 2961 12356 2973 12359
rect 2464 12328 2973 12356
rect 2464 12316 2470 12328
rect 2961 12325 2973 12328
rect 3007 12325 3019 12359
rect 2961 12319 3019 12325
rect 3694 12316 3700 12368
rect 3752 12316 3758 12368
rect 4154 12316 4160 12368
rect 4212 12316 4218 12368
rect 569 12291 627 12297
rect 569 12257 581 12291
rect 615 12257 627 12291
rect 2777 12291 2835 12297
rect 2777 12288 2789 12291
rect 569 12251 627 12257
rect 2332 12260 2789 12288
rect 842 12180 848 12232
rect 900 12180 906 12232
rect 2332 12096 2360 12260
rect 2777 12257 2789 12260
rect 2823 12257 2835 12291
rect 2777 12251 2835 12257
rect 5184 12288 5212 12396
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 5592 12396 5764 12424
rect 5592 12384 5598 12396
rect 5629 12359 5687 12365
rect 5629 12325 5641 12359
rect 5675 12325 5687 12359
rect 5629 12319 5687 12325
rect 5445 12291 5503 12297
rect 5445 12288 5457 12291
rect 5184 12260 5457 12288
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 5184 12229 5212 12260
rect 5445 12257 5457 12260
rect 5491 12257 5503 12291
rect 5445 12251 5503 12257
rect 5644 12232 5672 12319
rect 5736 12288 5764 12396
rect 5810 12384 5816 12436
rect 5868 12384 5874 12436
rect 14829 12427 14887 12433
rect 14829 12393 14841 12427
rect 14875 12424 14887 12427
rect 15102 12424 15108 12436
rect 14875 12396 15108 12424
rect 14875 12393 14887 12396
rect 14829 12387 14887 12393
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 6181 12359 6239 12365
rect 6181 12325 6193 12359
rect 6227 12356 6239 12359
rect 6641 12359 6699 12365
rect 6641 12356 6653 12359
rect 6227 12328 6653 12356
rect 6227 12325 6239 12328
rect 6181 12319 6239 12325
rect 6641 12325 6653 12328
rect 6687 12325 6699 12359
rect 6641 12319 6699 12325
rect 6089 12291 6147 12297
rect 6089 12288 6101 12291
rect 5736 12260 6101 12288
rect 6089 12257 6101 12260
rect 6135 12257 6147 12291
rect 6089 12251 6147 12257
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12257 6331 12291
rect 6273 12251 6331 12257
rect 5169 12223 5227 12229
rect 3476 12192 5120 12220
rect 3476 12180 3482 12192
rect 5092 12152 5120 12192
rect 5169 12189 5181 12223
rect 5215 12189 5227 12223
rect 5169 12183 5227 12189
rect 5626 12180 5632 12232
rect 5684 12180 5690 12232
rect 6178 12180 6184 12232
rect 6236 12220 6242 12232
rect 6288 12220 6316 12251
rect 7742 12248 7748 12300
rect 7800 12248 7806 12300
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 6236 12192 6316 12220
rect 6236 12180 6242 12192
rect 6362 12180 6368 12232
rect 6420 12220 6426 12232
rect 14936 12220 14964 12251
rect 15102 12248 15108 12300
rect 15160 12248 15166 12300
rect 15194 12220 15200 12232
rect 6420 12192 6500 12220
rect 14936 12192 15200 12220
rect 6420 12180 6426 12192
rect 6472 12152 6500 12192
rect 15194 12180 15200 12192
rect 15252 12180 15258 12232
rect 5092 12124 6500 12152
rect 2314 12044 2320 12096
rect 2372 12044 2378 12096
rect 3142 12044 3148 12096
rect 3200 12044 3206 12096
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8113 12087 8171 12093
rect 8113 12084 8125 12087
rect 8076 12056 8125 12084
rect 8076 12044 8082 12056
rect 8113 12053 8125 12056
rect 8159 12053 8171 12087
rect 8113 12047 8171 12053
rect 15378 12044 15384 12096
rect 15436 12044 15442 12096
rect 92 11994 15824 12016
rect 92 11942 1904 11994
rect 1956 11942 1968 11994
rect 2020 11942 2032 11994
rect 2084 11942 2096 11994
rect 2148 11942 2160 11994
rect 2212 11942 5837 11994
rect 5889 11942 5901 11994
rect 5953 11942 5965 11994
rect 6017 11942 6029 11994
rect 6081 11942 6093 11994
rect 6145 11942 9770 11994
rect 9822 11942 9834 11994
rect 9886 11942 9898 11994
rect 9950 11942 9962 11994
rect 10014 11942 10026 11994
rect 10078 11942 13703 11994
rect 13755 11942 13767 11994
rect 13819 11942 13831 11994
rect 13883 11942 13895 11994
rect 13947 11942 13959 11994
rect 14011 11942 15824 11994
rect 92 11920 15824 11942
rect 842 11840 848 11892
rect 900 11880 906 11892
rect 1213 11883 1271 11889
rect 1213 11880 1225 11883
rect 900 11852 1225 11880
rect 900 11840 906 11852
rect 1213 11849 1225 11852
rect 1259 11849 1271 11883
rect 1213 11843 1271 11849
rect 1302 11840 1308 11892
rect 1360 11880 1366 11892
rect 3050 11880 3056 11892
rect 1360 11852 3056 11880
rect 1360 11840 1366 11852
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 3142 11840 3148 11892
rect 3200 11840 3206 11892
rect 3326 11840 3332 11892
rect 3384 11840 3390 11892
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 4120 11852 5764 11880
rect 4120 11840 4126 11852
rect 1397 11815 1455 11821
rect 1397 11812 1409 11815
rect 1228 11784 1409 11812
rect 661 11679 719 11685
rect 661 11645 673 11679
rect 707 11645 719 11679
rect 661 11639 719 11645
rect 1029 11679 1087 11685
rect 1029 11645 1041 11679
rect 1075 11676 1087 11679
rect 1118 11676 1124 11688
rect 1075 11648 1124 11676
rect 1075 11645 1087 11648
rect 1029 11639 1087 11645
rect 676 11608 704 11639
rect 1118 11636 1124 11648
rect 1176 11636 1182 11688
rect 1228 11685 1256 11784
rect 1397 11781 1409 11784
rect 1443 11781 1455 11815
rect 1397 11775 1455 11781
rect 1320 11716 2774 11744
rect 1213 11679 1271 11685
rect 1213 11645 1225 11679
rect 1259 11645 1271 11679
rect 1213 11639 1271 11645
rect 1320 11608 1348 11716
rect 1578 11636 1584 11688
rect 1636 11676 1642 11688
rect 1673 11679 1731 11685
rect 1673 11676 1685 11679
rect 1636 11648 1685 11676
rect 1636 11636 1642 11648
rect 1673 11645 1685 11648
rect 1719 11645 1731 11679
rect 1673 11639 1731 11645
rect 676 11580 1348 11608
rect 1397 11611 1455 11617
rect 1397 11577 1409 11611
rect 1443 11608 1455 11611
rect 2314 11608 2320 11620
rect 1443 11580 2320 11608
rect 1443 11577 1455 11580
rect 1397 11571 1455 11577
rect 2314 11568 2320 11580
rect 2372 11568 2378 11620
rect 474 11500 480 11552
rect 532 11500 538 11552
rect 1581 11543 1639 11549
rect 1581 11509 1593 11543
rect 1627 11540 1639 11543
rect 1762 11540 1768 11552
rect 1627 11512 1768 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 1762 11500 1768 11512
rect 1820 11540 1826 11552
rect 2406 11540 2412 11552
rect 1820 11512 2412 11540
rect 1820 11500 1826 11512
rect 2406 11500 2412 11512
rect 2464 11500 2470 11552
rect 2746 11540 2774 11716
rect 3068 11676 3096 11840
rect 3160 11744 3188 11840
rect 4341 11815 4399 11821
rect 4341 11781 4353 11815
rect 4387 11812 4399 11815
rect 4387 11784 4844 11812
rect 4387 11781 4399 11784
rect 4341 11775 4399 11781
rect 3160 11716 4200 11744
rect 3329 11679 3387 11685
rect 3329 11678 3341 11679
rect 3252 11676 3341 11678
rect 3068 11650 3341 11676
rect 3068 11648 3280 11650
rect 3329 11645 3341 11650
rect 3375 11645 3387 11679
rect 3329 11639 3387 11645
rect 3513 11679 3571 11685
rect 3513 11645 3525 11679
rect 3559 11645 3571 11679
rect 3513 11639 3571 11645
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11676 3663 11679
rect 4062 11676 4068 11688
rect 3651 11648 4068 11676
rect 3651 11645 3663 11648
rect 3605 11639 3663 11645
rect 2958 11568 2964 11620
rect 3016 11608 3022 11620
rect 3528 11608 3556 11639
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4172 11685 4200 11716
rect 4816 11685 4844 11784
rect 5736 11688 5764 11852
rect 6178 11840 6184 11892
rect 6236 11840 6242 11892
rect 6012 11716 8248 11744
rect 6012 11688 6040 11716
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11676 4859 11679
rect 5442 11676 5448 11688
rect 4847 11648 5448 11676
rect 4847 11645 4859 11648
rect 4801 11639 4859 11645
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 5718 11636 5724 11688
rect 5776 11676 5782 11688
rect 5905 11679 5963 11685
rect 5905 11676 5917 11679
rect 5776 11648 5917 11676
rect 5776 11636 5782 11648
rect 5905 11645 5917 11648
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 5994 11636 6000 11688
rect 6052 11636 6058 11688
rect 6730 11636 6736 11688
rect 6788 11636 6794 11688
rect 6181 11611 6239 11617
rect 6181 11608 6193 11611
rect 3016 11580 3556 11608
rect 4816 11580 6193 11608
rect 3016 11568 3022 11580
rect 4816 11540 4844 11580
rect 6181 11577 6193 11580
rect 6227 11608 6239 11611
rect 8018 11608 8024 11620
rect 6227 11580 8024 11608
rect 6227 11577 6239 11580
rect 6181 11571 6239 11577
rect 8018 11568 8024 11580
rect 8076 11568 8082 11620
rect 8220 11617 8248 11716
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 8435 11648 8769 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 8757 11645 8769 11648
rect 8803 11645 8815 11679
rect 8757 11639 8815 11645
rect 8205 11611 8263 11617
rect 8205 11577 8217 11611
rect 8251 11608 8263 11611
rect 8478 11608 8484 11620
rect 8251 11580 8484 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 8478 11568 8484 11580
rect 8536 11568 8542 11620
rect 2746 11512 4844 11540
rect 4890 11500 4896 11552
rect 4948 11500 4954 11552
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6328 11512 6837 11540
rect 6328 11500 6334 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 8941 11543 8999 11549
rect 8941 11509 8953 11543
rect 8987 11540 8999 11543
rect 9030 11540 9036 11552
rect 8987 11512 9036 11540
rect 8987 11509 8999 11512
rect 8941 11503 8999 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 92 11450 15824 11472
rect 92 11398 2564 11450
rect 2616 11398 2628 11450
rect 2680 11398 2692 11450
rect 2744 11398 2756 11450
rect 2808 11398 2820 11450
rect 2872 11398 6497 11450
rect 6549 11398 6561 11450
rect 6613 11398 6625 11450
rect 6677 11398 6689 11450
rect 6741 11398 6753 11450
rect 6805 11398 10430 11450
rect 10482 11398 10494 11450
rect 10546 11398 10558 11450
rect 10610 11398 10622 11450
rect 10674 11398 10686 11450
rect 10738 11398 14363 11450
rect 14415 11398 14427 11450
rect 14479 11398 14491 11450
rect 14543 11398 14555 11450
rect 14607 11398 14619 11450
rect 14671 11398 15824 11450
rect 92 11376 15824 11398
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2363 11308 2452 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2424 11280 2452 11308
rect 2958 11296 2964 11348
rect 3016 11336 3022 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 3016 11308 5181 11336
rect 3016 11296 3022 11308
rect 5169 11305 5181 11308
rect 5215 11336 5227 11339
rect 5626 11336 5632 11348
rect 5215 11308 5632 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 5626 11296 5632 11308
rect 5684 11336 5690 11348
rect 6457 11339 6515 11345
rect 5684 11308 6224 11336
rect 5684 11296 5690 11308
rect 750 11268 756 11280
rect 584 11240 756 11268
rect 584 11209 612 11240
rect 750 11228 756 11240
rect 808 11228 814 11280
rect 1486 11228 1492 11280
rect 1544 11228 1550 11280
rect 2406 11228 2412 11280
rect 2464 11268 2470 11280
rect 3053 11271 3111 11277
rect 3053 11268 3065 11271
rect 2464 11240 3065 11268
rect 2464 11228 2470 11240
rect 3053 11237 3065 11240
rect 3099 11237 3111 11271
rect 3053 11231 3111 11237
rect 4154 11228 4160 11280
rect 4212 11228 4218 11280
rect 6196 11277 6224 11308
rect 6457 11305 6469 11339
rect 6503 11305 6515 11339
rect 6457 11299 6515 11305
rect 6089 11271 6147 11277
rect 6089 11268 6101 11271
rect 5644 11240 6101 11268
rect 5644 11212 5672 11240
rect 6089 11237 6101 11240
rect 6135 11237 6147 11271
rect 6089 11231 6147 11237
rect 6181 11271 6239 11277
rect 6181 11237 6193 11271
rect 6227 11237 6239 11271
rect 6472 11268 6500 11299
rect 8478 11296 8484 11348
rect 8536 11296 8542 11348
rect 14829 11339 14887 11345
rect 14829 11305 14841 11339
rect 14875 11336 14887 11339
rect 15102 11336 15108 11348
rect 14875 11308 15108 11336
rect 14875 11305 14887 11308
rect 14829 11299 14887 11305
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 7009 11271 7067 11277
rect 7009 11268 7021 11271
rect 6472 11240 7021 11268
rect 6181 11231 6239 11237
rect 7009 11237 7021 11240
rect 7055 11237 7067 11271
rect 7009 11231 7067 11237
rect 7742 11228 7748 11280
rect 7800 11228 7806 11280
rect 569 11203 627 11209
rect 569 11169 581 11203
rect 615 11169 627 11203
rect 569 11163 627 11169
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11169 2743 11203
rect 2685 11163 2743 11169
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 2866 11200 2872 11212
rect 2823 11172 2872 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 842 11092 848 11144
rect 900 11092 906 11144
rect 2700 11132 2728 11163
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 2961 11203 3019 11209
rect 2961 11169 2973 11203
rect 3007 11169 3019 11203
rect 3145 11203 3203 11209
rect 3145 11200 3157 11203
rect 2961 11163 3019 11169
rect 3068 11172 3157 11200
rect 2700 11104 2912 11132
rect 2590 10956 2596 11008
rect 2648 10956 2654 11008
rect 2884 10996 2912 11104
rect 2976 11064 3004 11163
rect 3068 11144 3096 11172
rect 3145 11169 3157 11172
rect 3191 11169 3203 11203
rect 3145 11163 3203 11169
rect 5626 11160 5632 11212
rect 5684 11160 5690 11212
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11200 5963 11203
rect 5994 11200 6000 11212
rect 5951 11172 6000 11200
rect 5951 11169 5963 11172
rect 5905 11163 5963 11169
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 6454 11200 6460 11212
rect 6319 11172 6460 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 14918 11160 14924 11212
rect 14976 11160 14982 11212
rect 15102 11160 15108 11212
rect 15160 11160 15166 11212
rect 3050 11092 3056 11144
rect 3108 11092 3114 11144
rect 3418 11092 3424 11144
rect 3476 11092 3482 11144
rect 3697 11135 3755 11141
rect 3697 11132 3709 11135
rect 3528 11104 3709 11132
rect 3329 11067 3387 11073
rect 2976 11036 3188 11064
rect 3160 11008 3188 11036
rect 3329 11033 3341 11067
rect 3375 11064 3387 11067
rect 3528 11064 3556 11104
rect 3697 11101 3709 11104
rect 3743 11101 3755 11135
rect 3697 11095 3755 11101
rect 6362 11092 6368 11144
rect 6420 11132 6426 11144
rect 6733 11135 6791 11141
rect 6733 11132 6745 11135
rect 6420 11104 6745 11132
rect 6420 11092 6426 11104
rect 6733 11101 6745 11104
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 3375 11036 3556 11064
rect 3375 11033 3387 11036
rect 3329 11027 3387 11033
rect 15378 11024 15384 11076
rect 15436 11024 15442 11076
rect 2958 10996 2964 11008
rect 2884 10968 2964 10996
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 3142 10956 3148 11008
rect 3200 10956 3206 11008
rect 92 10906 15824 10928
rect 92 10854 1904 10906
rect 1956 10854 1968 10906
rect 2020 10854 2032 10906
rect 2084 10854 2096 10906
rect 2148 10854 2160 10906
rect 2212 10854 5837 10906
rect 5889 10854 5901 10906
rect 5953 10854 5965 10906
rect 6017 10854 6029 10906
rect 6081 10854 6093 10906
rect 6145 10854 9770 10906
rect 9822 10854 9834 10906
rect 9886 10854 9898 10906
rect 9950 10854 9962 10906
rect 10014 10854 10026 10906
rect 10078 10854 13703 10906
rect 13755 10854 13767 10906
rect 13819 10854 13831 10906
rect 13883 10854 13895 10906
rect 13947 10854 13959 10906
rect 14011 10854 15824 10906
rect 92 10832 15824 10854
rect 842 10752 848 10804
rect 900 10792 906 10804
rect 1397 10795 1455 10801
rect 1397 10792 1409 10795
rect 900 10764 1409 10792
rect 900 10752 906 10764
rect 1397 10761 1409 10764
rect 1443 10761 1455 10795
rect 1397 10755 1455 10761
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 4120 10764 11836 10792
rect 4120 10752 4126 10764
rect 5810 10684 5816 10736
rect 5868 10724 5874 10736
rect 6454 10724 6460 10736
rect 5868 10696 6460 10724
rect 5868 10684 5874 10696
rect 6454 10684 6460 10696
rect 6512 10684 6518 10736
rect 5534 10656 5540 10668
rect 1596 10628 5540 10656
rect 661 10591 719 10597
rect 661 10557 673 10591
rect 707 10557 719 10591
rect 661 10551 719 10557
rect 676 10520 704 10551
rect 1118 10548 1124 10600
rect 1176 10588 1182 10600
rect 1596 10597 1624 10628
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 6362 10616 6368 10668
rect 6420 10656 6426 10668
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 6420 10628 7941 10656
rect 6420 10616 6426 10628
rect 7929 10625 7941 10628
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 1581 10591 1639 10597
rect 1581 10588 1593 10591
rect 1176 10560 1593 10588
rect 1176 10548 1182 10560
rect 1581 10557 1593 10560
rect 1627 10557 1639 10591
rect 1581 10551 1639 10557
rect 1762 10548 1768 10600
rect 1820 10548 1826 10600
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2590 10588 2596 10600
rect 1903 10560 2596 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 6086 10548 6092 10600
rect 6144 10548 6150 10600
rect 6178 10548 6184 10600
rect 6236 10588 6242 10600
rect 6236 10560 6408 10588
rect 6236 10548 6242 10560
rect 5994 10520 6000 10532
rect 676 10492 6000 10520
rect 5994 10480 6000 10492
rect 6052 10480 6058 10532
rect 6380 10529 6408 10560
rect 6454 10548 6460 10600
rect 6512 10588 6518 10600
rect 6822 10588 6828 10600
rect 6512 10560 6828 10588
rect 6512 10548 6518 10560
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 9858 10548 9864 10600
rect 9916 10548 9922 10600
rect 11808 10597 11836 10764
rect 15102 10752 15108 10804
rect 15160 10752 15166 10804
rect 11977 10727 12035 10733
rect 11977 10693 11989 10727
rect 12023 10724 12035 10727
rect 12023 10696 12388 10724
rect 12023 10693 12035 10696
rect 11977 10687 12035 10693
rect 12360 10600 12388 10696
rect 11793 10591 11851 10597
rect 11793 10557 11805 10591
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 12342 10548 12348 10600
rect 12400 10548 12406 10600
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15562 10588 15568 10600
rect 15059 10560 15568 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15562 10548 15568 10560
rect 15620 10548 15626 10600
rect 6273 10523 6331 10529
rect 6273 10489 6285 10523
rect 6319 10489 6331 10523
rect 6273 10483 6331 10489
rect 6365 10523 6423 10529
rect 6365 10489 6377 10523
rect 6411 10489 6423 10523
rect 8205 10523 8263 10529
rect 8205 10520 8217 10523
rect 6365 10483 6423 10489
rect 6656 10492 8217 10520
rect 474 10412 480 10464
rect 532 10412 538 10464
rect 5626 10412 5632 10464
rect 5684 10452 5690 10464
rect 6288 10452 6316 10483
rect 6656 10461 6684 10492
rect 8205 10489 8217 10492
rect 8251 10489 8263 10523
rect 9490 10520 9496 10532
rect 9430 10492 9496 10520
rect 8205 10483 8263 10489
rect 9490 10480 9496 10492
rect 9548 10480 9554 10532
rect 5684 10424 6316 10452
rect 6641 10455 6699 10461
rect 5684 10412 5690 10424
rect 6641 10421 6653 10455
rect 6687 10421 6699 10455
rect 6641 10415 6699 10421
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 9677 10455 9735 10461
rect 9677 10452 9689 10455
rect 9272 10424 9689 10452
rect 9272 10412 9278 10424
rect 9677 10421 9689 10424
rect 9723 10421 9735 10455
rect 9677 10415 9735 10421
rect 10045 10455 10103 10461
rect 10045 10421 10057 10455
rect 10091 10452 10103 10455
rect 11054 10452 11060 10464
rect 10091 10424 11060 10452
rect 10091 10421 10103 10424
rect 10045 10415 10103 10421
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 12434 10412 12440 10464
rect 12492 10412 12498 10464
rect 92 10362 15824 10384
rect 92 10310 2564 10362
rect 2616 10310 2628 10362
rect 2680 10310 2692 10362
rect 2744 10310 2756 10362
rect 2808 10310 2820 10362
rect 2872 10310 6497 10362
rect 6549 10310 6561 10362
rect 6613 10310 6625 10362
rect 6677 10310 6689 10362
rect 6741 10310 6753 10362
rect 6805 10310 10430 10362
rect 10482 10310 10494 10362
rect 10546 10310 10558 10362
rect 10610 10310 10622 10362
rect 10674 10310 10686 10362
rect 10738 10310 14363 10362
rect 14415 10310 14427 10362
rect 14479 10310 14491 10362
rect 14543 10310 14555 10362
rect 14607 10310 14619 10362
rect 14671 10310 15824 10362
rect 92 10288 15824 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 5810 10248 5816 10260
rect 1544 10220 4200 10248
rect 1544 10208 1550 10220
rect 1780 10098 1808 10220
rect 2774 10140 2780 10192
rect 2832 10180 2838 10192
rect 3053 10183 3111 10189
rect 3053 10180 3065 10183
rect 2832 10152 3065 10180
rect 2832 10140 2838 10152
rect 3053 10149 3065 10152
rect 3099 10149 3111 10183
rect 3053 10143 3111 10149
rect 4172 10124 4200 10220
rect 4816 10220 5816 10248
rect 2317 10115 2375 10121
rect 2317 10112 2329 10115
rect 2148 10084 2329 10112
rect 385 10047 443 10053
rect 385 10013 397 10047
rect 431 10013 443 10047
rect 385 10007 443 10013
rect 400 9908 428 10007
rect 658 10004 664 10056
rect 716 10004 722 10056
rect 1670 10004 1676 10056
rect 1728 10044 1734 10056
rect 2148 10053 2176 10084
rect 2317 10081 2329 10084
rect 2363 10081 2375 10115
rect 2317 10075 2375 10081
rect 2498 10072 2504 10124
rect 2556 10072 2562 10124
rect 4154 10072 4160 10124
rect 4212 10072 4218 10124
rect 4816 10121 4844 10220
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 5902 10208 5908 10260
rect 5960 10248 5966 10260
rect 6174 10251 6232 10257
rect 6174 10248 6186 10251
rect 5960 10220 6186 10248
rect 5960 10208 5966 10220
rect 6174 10217 6186 10220
rect 6220 10217 6232 10251
rect 9214 10248 9220 10260
rect 6174 10211 6232 10217
rect 6288 10220 9220 10248
rect 4893 10183 4951 10189
rect 4893 10149 4905 10183
rect 4939 10180 4951 10183
rect 6086 10180 6092 10192
rect 4939 10152 6092 10180
rect 4939 10149 4951 10152
rect 4893 10143 4951 10149
rect 6086 10140 6092 10152
rect 6144 10180 6150 10192
rect 6288 10180 6316 10220
rect 6144 10152 6316 10180
rect 6144 10140 6150 10152
rect 7742 10140 7748 10192
rect 7800 10140 7806 10192
rect 9140 10189 9168 10220
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 9309 10251 9367 10257
rect 9309 10217 9321 10251
rect 9355 10248 9367 10251
rect 9858 10248 9864 10260
rect 9355 10220 9864 10248
rect 9355 10217 9367 10220
rect 9309 10211 9367 10217
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 9125 10183 9183 10189
rect 9125 10149 9137 10183
rect 9171 10149 9183 10183
rect 9125 10143 9183 10149
rect 4801 10115 4859 10121
rect 4801 10081 4813 10115
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 4985 10115 5043 10121
rect 4985 10081 4997 10115
rect 5031 10081 5043 10115
rect 4985 10075 5043 10081
rect 2133 10047 2191 10053
rect 2133 10044 2145 10047
rect 1728 10016 2145 10044
rect 1728 10004 1734 10016
rect 2133 10013 2145 10016
rect 2179 10013 2191 10047
rect 2133 10007 2191 10013
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 3050 10044 3056 10056
rect 2823 10016 3056 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 2792 9976 2820 10007
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 3142 10004 3148 10056
rect 3200 10044 3206 10056
rect 5000 10044 5028 10075
rect 5166 10072 5172 10124
rect 5224 10072 5230 10124
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 5721 10115 5779 10121
rect 5721 10112 5733 10115
rect 5500 10084 5733 10112
rect 5500 10072 5506 10084
rect 5721 10081 5733 10084
rect 5767 10081 5779 10115
rect 5721 10075 5779 10081
rect 5902 10072 5908 10124
rect 5960 10072 5966 10124
rect 5997 10115 6055 10121
rect 5997 10081 6009 10115
rect 6043 10081 6055 10115
rect 5997 10075 6055 10081
rect 3200 10016 5580 10044
rect 3200 10004 3206 10016
rect 1688 9948 2820 9976
rect 750 9908 756 9920
rect 400 9880 756 9908
rect 750 9868 756 9880
rect 808 9908 814 9920
rect 1688 9908 1716 9948
rect 5552 9920 5580 10016
rect 5718 9936 5724 9988
rect 5776 9976 5782 9988
rect 6012 9976 6040 10075
rect 6178 10072 6184 10124
rect 6236 10112 6242 10124
rect 6273 10115 6331 10121
rect 6273 10112 6285 10115
rect 6236 10084 6285 10112
rect 6236 10072 6242 10084
rect 6273 10081 6285 10084
rect 6319 10081 6331 10115
rect 6273 10075 6331 10081
rect 6362 10072 6368 10124
rect 6420 10112 6426 10124
rect 6457 10115 6515 10121
rect 6457 10112 6469 10115
rect 6420 10084 6469 10112
rect 6420 10072 6426 10084
rect 6457 10081 6469 10084
rect 6503 10081 6515 10115
rect 8941 10115 8999 10121
rect 8941 10112 8953 10115
rect 6457 10075 6515 10081
rect 8220 10084 8953 10112
rect 6733 10047 6791 10053
rect 6733 10044 6745 10047
rect 5776 9948 6040 9976
rect 6104 10016 6745 10044
rect 5776 9936 5782 9948
rect 808 9880 1716 9908
rect 808 9868 814 9880
rect 2682 9868 2688 9920
rect 2740 9868 2746 9920
rect 4522 9868 4528 9920
rect 4580 9868 4586 9920
rect 4617 9911 4675 9917
rect 4617 9877 4629 9911
rect 4663 9908 4675 9911
rect 4706 9908 4712 9920
rect 4663 9880 4712 9908
rect 4663 9877 4675 9880
rect 4617 9871 4675 9877
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 5534 9868 5540 9920
rect 5592 9868 5598 9920
rect 5905 9911 5963 9917
rect 5905 9877 5917 9911
rect 5951 9908 5963 9911
rect 6104 9908 6132 10016
rect 6733 10013 6745 10016
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 6178 9936 6184 9988
rect 6236 9936 6242 9988
rect 5951 9880 6132 9908
rect 6196 9908 6224 9936
rect 8220 9917 8248 10084
rect 8941 10081 8953 10084
rect 8987 10081 8999 10115
rect 8941 10075 8999 10081
rect 15102 10072 15108 10124
rect 15160 10072 15166 10124
rect 8205 9911 8263 9917
rect 8205 9908 8217 9911
rect 6196 9880 8217 9908
rect 5951 9877 5963 9880
rect 5905 9871 5963 9877
rect 8205 9877 8217 9880
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 15378 9868 15384 9920
rect 15436 9868 15442 9920
rect 92 9818 15824 9840
rect 92 9766 1904 9818
rect 1956 9766 1968 9818
rect 2020 9766 2032 9818
rect 2084 9766 2096 9818
rect 2148 9766 2160 9818
rect 2212 9766 5837 9818
rect 5889 9766 5901 9818
rect 5953 9766 5965 9818
rect 6017 9766 6029 9818
rect 6081 9766 6093 9818
rect 6145 9766 9770 9818
rect 9822 9766 9834 9818
rect 9886 9766 9898 9818
rect 9950 9766 9962 9818
rect 10014 9766 10026 9818
rect 10078 9766 13703 9818
rect 13755 9766 13767 9818
rect 13819 9766 13831 9818
rect 13883 9766 13895 9818
rect 13947 9766 13959 9818
rect 14011 9766 15824 9818
rect 92 9744 15824 9766
rect 658 9664 664 9716
rect 716 9704 722 9716
rect 1121 9707 1179 9713
rect 1121 9704 1133 9707
rect 716 9676 1133 9704
rect 716 9664 722 9676
rect 1121 9673 1133 9676
rect 1167 9673 1179 9707
rect 1121 9667 1179 9673
rect 2682 9664 2688 9716
rect 2740 9664 2746 9716
rect 4062 9704 4068 9716
rect 2792 9676 4068 9704
rect 1581 9639 1639 9645
rect 1581 9605 1593 9639
rect 1627 9605 1639 9639
rect 2700 9636 2728 9664
rect 2792 9636 2820 9676
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 5166 9704 5172 9716
rect 4172 9676 5172 9704
rect 4172 9636 4200 9676
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 7742 9704 7748 9716
rect 6886 9676 7748 9704
rect 2700 9608 2820 9636
rect 2884 9608 4200 9636
rect 1581 9599 1639 9605
rect 661 9503 719 9509
rect 661 9469 673 9503
rect 707 9469 719 9503
rect 661 9463 719 9469
rect 937 9503 995 9509
rect 937 9469 949 9503
rect 983 9500 995 9503
rect 1026 9500 1032 9512
rect 983 9472 1032 9500
rect 983 9469 995 9472
rect 937 9463 995 9469
rect 676 9432 704 9463
rect 1026 9460 1032 9472
rect 1084 9460 1090 9512
rect 1121 9503 1179 9509
rect 1121 9469 1133 9503
rect 1167 9500 1179 9503
rect 1596 9500 1624 9599
rect 1762 9528 1768 9580
rect 1820 9528 1826 9580
rect 1167 9472 1624 9500
rect 1780 9500 1808 9528
rect 1857 9503 1915 9509
rect 1857 9500 1869 9503
rect 1780 9472 1869 9500
rect 1167 9469 1179 9472
rect 1121 9463 1179 9469
rect 1857 9469 1869 9472
rect 1903 9469 1915 9503
rect 1857 9463 1915 9469
rect 1581 9435 1639 9441
rect 1581 9432 1593 9435
rect 676 9404 1593 9432
rect 1581 9401 1593 9404
rect 1627 9432 1639 9435
rect 1670 9432 1676 9444
rect 1627 9404 1676 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 1670 9392 1676 9404
rect 1728 9392 1734 9444
rect 1765 9435 1823 9441
rect 1765 9401 1777 9435
rect 1811 9432 1823 9435
rect 2498 9432 2504 9444
rect 1811 9404 2504 9432
rect 1811 9401 1823 9404
rect 1765 9395 1823 9401
rect 2498 9392 2504 9404
rect 2556 9432 2562 9444
rect 2884 9432 2912 9608
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3418 9568 3424 9580
rect 3108 9540 3424 9568
rect 3108 9528 3114 9540
rect 3418 9528 3424 9540
rect 3476 9568 3482 9580
rect 4433 9571 4491 9577
rect 4433 9568 4445 9571
rect 3476 9540 4445 9568
rect 3476 9528 3482 9540
rect 4433 9537 4445 9540
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4706 9528 4712 9580
rect 4764 9528 4770 9580
rect 5166 9528 5172 9580
rect 5224 9568 5230 9580
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 5224 9540 6193 9568
rect 5224 9528 5230 9540
rect 6181 9537 6193 9540
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 3329 9503 3387 9509
rect 3016 9472 3280 9500
rect 3016 9460 3022 9472
rect 3053 9435 3111 9441
rect 3053 9432 3065 9435
rect 2556 9404 3065 9432
rect 2556 9392 2562 9404
rect 3053 9401 3065 9404
rect 3099 9401 3111 9435
rect 3053 9395 3111 9401
rect 3142 9392 3148 9444
rect 3200 9392 3206 9444
rect 474 9324 480 9376
rect 532 9324 538 9376
rect 2774 9324 2780 9376
rect 2832 9324 2838 9376
rect 2958 9324 2964 9376
rect 3016 9364 3022 9376
rect 3160 9364 3188 9392
rect 3016 9336 3188 9364
rect 3252 9364 3280 9472
rect 3329 9469 3341 9503
rect 3375 9469 3387 9503
rect 6886 9500 6914 9676
rect 7742 9664 7748 9676
rect 7800 9664 7806 9716
rect 15010 9596 15016 9648
rect 15068 9596 15074 9648
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9568 8263 9571
rect 10229 9571 10287 9577
rect 10229 9568 10241 9571
rect 8251 9540 10241 9568
rect 8251 9537 8263 9540
rect 8205 9531 8263 9537
rect 10229 9537 10241 9540
rect 10275 9568 10287 9571
rect 11698 9568 11704 9580
rect 10275 9540 11704 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 13504 9540 14289 9568
rect 13504 9528 13510 9540
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14277 9531 14335 9537
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9568 14795 9571
rect 14921 9571 14979 9577
rect 14921 9568 14933 9571
rect 14783 9540 14933 9568
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 14921 9537 14933 9540
rect 14967 9537 14979 9571
rect 14921 9531 14979 9537
rect 5842 9486 6914 9500
rect 3329 9463 3387 9469
rect 5828 9472 6914 9486
rect 10597 9503 10655 9509
rect 3344 9432 3372 9463
rect 3344 9404 4568 9432
rect 4540 9376 4568 9404
rect 3418 9364 3424 9376
rect 3252 9336 3424 9364
rect 3016 9324 3022 9336
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 4522 9324 4528 9376
rect 4580 9324 4586 9376
rect 5350 9324 5356 9376
rect 5408 9364 5414 9376
rect 5828 9364 5856 9472
rect 10597 9469 10609 9503
rect 10643 9500 10655 9503
rect 10686 9500 10692 9512
rect 10643 9472 10692 9500
rect 10643 9469 10655 9472
rect 10597 9463 10655 9469
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 14645 9503 14703 9509
rect 14645 9469 14657 9503
rect 14691 9500 14703 9503
rect 14691 9472 14780 9500
rect 14691 9469 14703 9472
rect 14645 9463 14703 9469
rect 8478 9392 8484 9444
rect 8536 9392 8542 9444
rect 9766 9432 9772 9444
rect 9706 9404 9772 9432
rect 9766 9392 9772 9404
rect 9824 9432 9830 9444
rect 13078 9432 13084 9444
rect 9824 9404 10272 9432
rect 9824 9392 9830 9404
rect 5408 9336 5856 9364
rect 9953 9367 10011 9373
rect 5408 9324 5414 9336
rect 9953 9333 9965 9367
rect 9999 9364 10011 9367
rect 10134 9364 10140 9376
rect 9999 9336 10140 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10244 9364 10272 9404
rect 10888 9404 10994 9432
rect 11716 9404 13084 9432
rect 10888 9376 10916 9404
rect 10870 9364 10876 9376
rect 10244 9336 10876 9364
rect 10870 9324 10876 9336
rect 10928 9364 10934 9376
rect 11716 9364 11744 9404
rect 13078 9392 13084 9404
rect 13136 9392 13142 9444
rect 14752 9376 14780 9472
rect 14826 9392 14832 9444
rect 14884 9432 14890 9444
rect 15381 9435 15439 9441
rect 15381 9432 15393 9435
rect 14884 9404 15393 9432
rect 14884 9392 14890 9404
rect 15381 9401 15393 9404
rect 15427 9401 15439 9435
rect 15381 9395 15439 9401
rect 10928 9336 11744 9364
rect 10928 9324 10934 9336
rect 11882 9324 11888 9376
rect 11940 9364 11946 9376
rect 12023 9367 12081 9373
rect 12023 9364 12035 9367
rect 11940 9336 12035 9364
rect 11940 9324 11946 9336
rect 12023 9333 12035 9336
rect 12069 9333 12081 9367
rect 12023 9327 12081 9333
rect 14734 9324 14740 9376
rect 14792 9324 14798 9376
rect 92 9274 15824 9296
rect 92 9222 2564 9274
rect 2616 9222 2628 9274
rect 2680 9222 2692 9274
rect 2744 9222 2756 9274
rect 2808 9222 2820 9274
rect 2872 9222 6497 9274
rect 6549 9222 6561 9274
rect 6613 9222 6625 9274
rect 6677 9222 6689 9274
rect 6741 9222 6753 9274
rect 6805 9222 10430 9274
rect 10482 9222 10494 9274
rect 10546 9222 10558 9274
rect 10610 9222 10622 9274
rect 10674 9222 10686 9274
rect 10738 9222 14363 9274
rect 14415 9222 14427 9274
rect 14479 9222 14491 9274
rect 14543 9222 14555 9274
rect 14607 9222 14619 9274
rect 14671 9222 15824 9274
rect 92 9200 15824 9222
rect 1762 9120 1768 9172
rect 1820 9160 1826 9172
rect 2682 9160 2688 9172
rect 1820 9132 2688 9160
rect 1820 9120 1826 9132
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 3234 9160 3240 9172
rect 2823 9132 3240 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 3234 9120 3240 9132
rect 3292 9160 3298 9172
rect 3292 9132 4016 9160
rect 3292 9120 3298 9132
rect 1486 9052 1492 9104
rect 1544 9052 1550 9104
rect 3988 9101 4016 9132
rect 5442 9120 5448 9172
rect 5500 9120 5506 9172
rect 6733 9163 6791 9169
rect 6733 9129 6745 9163
rect 6779 9160 6791 9163
rect 6822 9160 6828 9172
rect 6779 9132 6828 9160
rect 6779 9129 6791 9132
rect 6733 9123 6791 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 8757 9163 8815 9169
rect 8757 9160 8769 9163
rect 8536 9132 8769 9160
rect 8536 9120 8542 9132
rect 8757 9129 8769 9132
rect 8803 9129 8815 9163
rect 8757 9123 8815 9129
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 9766 9160 9772 9172
rect 9548 9132 9772 9160
rect 9548 9120 9554 9132
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 10689 9163 10747 9169
rect 10689 9129 10701 9163
rect 10735 9160 10747 9163
rect 10778 9160 10784 9172
rect 10735 9132 10784 9160
rect 10735 9129 10747 9132
rect 10689 9123 10747 9129
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 14826 9160 14832 9172
rect 10888 9132 13952 9160
rect 3973 9095 4031 9101
rect 2746 9064 3832 9092
rect 750 8984 756 9036
rect 808 8984 814 9036
rect 2593 9027 2651 9033
rect 2593 9024 2605 9027
rect 2516 8996 2605 9024
rect 1026 8916 1032 8968
rect 1084 8916 1090 8968
rect 750 8780 756 8832
rect 808 8820 814 8832
rect 2516 8829 2544 8996
rect 2593 8993 2605 8996
rect 2639 9024 2651 9027
rect 2746 9024 2774 9064
rect 3804 9033 3832 9064
rect 3973 9061 3985 9095
rect 4019 9092 4031 9095
rect 4522 9092 4528 9104
rect 4019 9064 4528 9092
rect 4019 9061 4031 9064
rect 3973 9055 4031 9061
rect 4522 9052 4528 9064
rect 4580 9052 4586 9104
rect 10888 9092 10916 9132
rect 11882 9092 11888 9104
rect 5644 9064 10916 9092
rect 11624 9064 11888 9092
rect 2639 8996 2774 9024
rect 2869 9027 2927 9033
rect 2639 8993 2651 8996
rect 2593 8987 2651 8993
rect 2869 8993 2881 9027
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 3789 9027 3847 9033
rect 3789 8993 3801 9027
rect 3835 8993 3847 9027
rect 3789 8987 3847 8993
rect 4157 9027 4215 9033
rect 4157 8993 4169 9027
rect 4203 9024 4215 9027
rect 5644 9024 5672 9064
rect 4203 8996 5672 9024
rect 5721 9027 5779 9033
rect 4203 8993 4215 8996
rect 4157 8987 4215 8993
rect 5721 8993 5733 9027
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 2884 8956 2912 8987
rect 2740 8928 2912 8956
rect 2740 8916 2774 8928
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 5736 8956 5764 8987
rect 6822 8984 6828 9036
rect 6880 9024 6886 9036
rect 6917 9027 6975 9033
rect 6917 9024 6929 9027
rect 6880 8996 6929 9024
rect 6880 8984 6886 8996
rect 6917 8993 6929 8996
rect 6963 8993 6975 9027
rect 6917 8987 6975 8993
rect 8846 8984 8852 9036
rect 8904 8984 8910 9036
rect 9582 8984 9588 9036
rect 9640 8984 9646 9036
rect 10873 9027 10931 9033
rect 10873 8993 10885 9027
rect 10919 9024 10931 9027
rect 10919 8996 11100 9024
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 5500 8928 5764 8956
rect 5500 8916 5506 8928
rect 2746 8888 2774 8916
rect 5718 8888 5724 8900
rect 2746 8860 5724 8888
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 11072 8897 11100 8996
rect 11422 8984 11428 9036
rect 11480 8984 11486 9036
rect 11624 8965 11652 9064
rect 11882 9052 11888 9064
rect 11940 9092 11946 9104
rect 11940 9064 12112 9092
rect 11940 9052 11946 9064
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 11977 9027 12035 9033
rect 11977 9024 11989 9027
rect 11756 8996 11989 9024
rect 11756 8984 11762 8996
rect 11977 8993 11989 8996
rect 12023 8993 12035 9027
rect 12084 9024 12112 9064
rect 13078 9052 13084 9104
rect 13136 9052 13142 9104
rect 13924 9033 13952 9132
rect 14384 9132 14832 9160
rect 14384 9033 14412 9132
rect 14826 9120 14832 9132
rect 14884 9120 14890 9172
rect 15010 9120 15016 9172
rect 15068 9120 15074 9172
rect 14734 9092 14740 9104
rect 14568 9064 14740 9092
rect 14568 9033 14596 9064
rect 14734 9052 14740 9064
rect 14792 9052 14798 9104
rect 13909 9027 13967 9033
rect 12084 8996 12480 9024
rect 11977 8987 12035 8993
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11057 8891 11115 8897
rect 11057 8857 11069 8891
rect 11103 8857 11115 8891
rect 11057 8851 11115 8857
rect 2501 8823 2559 8829
rect 2501 8820 2513 8823
rect 808 8792 2513 8820
rect 808 8780 814 8792
rect 2501 8789 2513 8792
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 2590 8780 2596 8832
rect 2648 8780 2654 8832
rect 2682 8780 2688 8832
rect 2740 8820 2746 8832
rect 4062 8820 4068 8832
rect 2740 8792 4068 8820
rect 2740 8780 2746 8792
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 11532 8820 11560 8919
rect 12342 8916 12348 8968
rect 12400 8916 12406 8968
rect 12452 8956 12480 8996
rect 13909 8993 13921 9027
rect 13955 8993 13967 9027
rect 13909 8987 13967 8993
rect 14369 9027 14427 9033
rect 14369 8993 14381 9027
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 14553 9027 14611 9033
rect 14553 8993 14565 9027
rect 14599 8993 14611 9027
rect 14553 8987 14611 8993
rect 14645 9027 14703 9033
rect 14645 8993 14657 9027
rect 14691 9024 14703 9027
rect 15028 9024 15056 9120
rect 14691 8996 15056 9024
rect 15105 9027 15163 9033
rect 14691 8993 14703 8996
rect 14645 8987 14703 8993
rect 15105 8993 15117 9027
rect 15151 8993 15163 9027
rect 15105 8987 15163 8993
rect 14568 8956 14596 8987
rect 12452 8928 14596 8956
rect 14734 8916 14740 8968
rect 14792 8956 14798 8968
rect 15120 8956 15148 8987
rect 14792 8928 15148 8956
rect 14792 8916 14798 8928
rect 13354 8820 13360 8832
rect 11532 8792 13360 8820
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 13538 8780 13544 8832
rect 13596 8820 13602 8832
rect 13771 8823 13829 8829
rect 13771 8820 13783 8823
rect 13596 8792 13783 8820
rect 13596 8780 13602 8792
rect 13771 8789 13783 8792
rect 13817 8789 13829 8823
rect 13771 8783 13829 8789
rect 14090 8780 14096 8832
rect 14148 8780 14154 8832
rect 14182 8780 14188 8832
rect 14240 8780 14246 8832
rect 15378 8780 15384 8832
rect 15436 8780 15442 8832
rect 92 8730 15824 8752
rect 92 8678 1904 8730
rect 1956 8678 1968 8730
rect 2020 8678 2032 8730
rect 2084 8678 2096 8730
rect 2148 8678 2160 8730
rect 2212 8678 5837 8730
rect 5889 8678 5901 8730
rect 5953 8678 5965 8730
rect 6017 8678 6029 8730
rect 6081 8678 6093 8730
rect 6145 8678 9770 8730
rect 9822 8678 9834 8730
rect 9886 8678 9898 8730
rect 9950 8678 9962 8730
rect 10014 8678 10026 8730
rect 10078 8678 13703 8730
rect 13755 8678 13767 8730
rect 13819 8678 13831 8730
rect 13883 8678 13895 8730
rect 13947 8678 13959 8730
rect 14011 8678 15824 8730
rect 92 8656 15824 8678
rect 1026 8576 1032 8628
rect 1084 8616 1090 8628
rect 1305 8619 1363 8625
rect 1305 8616 1317 8619
rect 1084 8588 1317 8616
rect 1084 8576 1090 8588
rect 1305 8585 1317 8588
rect 1351 8585 1363 8619
rect 1305 8579 1363 8585
rect 2590 8576 2596 8628
rect 2648 8576 2654 8628
rect 2958 8576 2964 8628
rect 3016 8576 3022 8628
rect 3234 8576 3240 8628
rect 3292 8576 3298 8628
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 5353 8619 5411 8625
rect 5353 8616 5365 8619
rect 4120 8588 5365 8616
rect 4120 8576 4126 8588
rect 5353 8585 5365 8588
rect 5399 8585 5411 8619
rect 5353 8579 5411 8585
rect 9769 8619 9827 8625
rect 9769 8585 9781 8619
rect 9815 8616 9827 8619
rect 11514 8616 11520 8628
rect 9815 8588 11520 8616
rect 9815 8585 9827 8588
rect 9769 8579 9827 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 12342 8576 12348 8628
rect 12400 8616 12406 8628
rect 13081 8619 13139 8625
rect 13081 8616 13093 8619
rect 12400 8588 13093 8616
rect 12400 8576 12406 8588
rect 13081 8585 13093 8588
rect 13127 8585 13139 8619
rect 13081 8579 13139 8585
rect 13446 8576 13452 8628
rect 13504 8576 13510 8628
rect 13538 8576 13544 8628
rect 13596 8576 13602 8628
rect 14553 8619 14611 8625
rect 14553 8585 14565 8619
rect 14599 8616 14611 8619
rect 15010 8616 15016 8628
rect 14599 8588 15016 8616
rect 14599 8585 14611 8588
rect 14553 8579 14611 8585
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 750 8372 756 8424
rect 808 8372 814 8424
rect 1118 8372 1124 8424
rect 1176 8372 1182 8424
rect 1305 8415 1363 8421
rect 1305 8381 1317 8415
rect 1351 8412 1363 8415
rect 2608 8412 2636 8576
rect 2976 8480 3004 8576
rect 2976 8452 3188 8480
rect 1351 8384 2636 8412
rect 1351 8381 1363 8384
rect 1305 8375 1363 8381
rect 2682 8372 2688 8424
rect 2740 8412 2746 8424
rect 3160 8421 3188 8452
rect 3252 8421 3280 8576
rect 3513 8551 3571 8557
rect 3513 8517 3525 8551
rect 3559 8517 3571 8551
rect 3513 8511 3571 8517
rect 5997 8551 6055 8557
rect 5997 8517 6009 8551
rect 6043 8517 6055 8551
rect 5997 8511 6055 8517
rect 6104 8520 9996 8548
rect 3528 8480 3556 8511
rect 3881 8483 3939 8489
rect 3881 8480 3893 8483
rect 3528 8452 3893 8480
rect 3881 8449 3893 8452
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 5718 8440 5724 8492
rect 5776 8440 5782 8492
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2740 8384 2973 8412
rect 2740 8372 2746 8384
rect 2961 8381 2973 8384
rect 3007 8381 3019 8415
rect 2961 8375 3019 8381
rect 3145 8415 3203 8421
rect 3145 8381 3157 8415
rect 3191 8381 3203 8415
rect 3145 8375 3203 8381
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 3418 8412 3424 8424
rect 3375 8384 3424 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 3602 8372 3608 8424
rect 3660 8372 3666 8424
rect 5350 8412 5356 8424
rect 5014 8384 5356 8412
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 5905 8415 5963 8421
rect 5905 8381 5917 8415
rect 5951 8412 5963 8415
rect 6012 8412 6040 8511
rect 5951 8384 6040 8412
rect 6104 8412 6132 8520
rect 6178 8440 6184 8492
rect 6236 8480 6242 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6236 8452 6561 8480
rect 6236 8440 6242 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8480 8447 8483
rect 9398 8480 9404 8492
rect 8435 8452 9404 8480
rect 8435 8449 8447 8452
rect 8389 8443 8447 8449
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 6104 8384 6377 8412
rect 5951 8381 5963 8384
rect 5905 8375 5963 8381
rect 382 8304 388 8356
rect 440 8304 446 8356
rect 2038 8304 2044 8356
rect 2096 8304 2102 8356
rect 2225 8347 2283 8353
rect 2225 8313 2237 8347
rect 2271 8344 2283 8347
rect 2314 8344 2320 8356
rect 2271 8316 2320 8344
rect 2271 8313 2283 8316
rect 2225 8307 2283 8313
rect 2314 8304 2320 8316
rect 2372 8304 2378 8356
rect 2409 8347 2467 8353
rect 2409 8313 2421 8347
rect 2455 8344 2467 8347
rect 2455 8316 3096 8344
rect 2455 8313 2467 8316
rect 2409 8307 2467 8313
rect 2056 8276 2084 8304
rect 2682 8276 2688 8288
rect 2056 8248 2688 8276
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 3068 8276 3096 8316
rect 3344 8316 4200 8344
rect 3344 8276 3372 8316
rect 3068 8248 3372 8276
rect 4172 8276 4200 8316
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 6104 8344 6132 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6564 8412 6592 8443
rect 9398 8440 9404 8452
rect 9456 8480 9462 8492
rect 9456 8452 9628 8480
rect 9456 8440 9462 8452
rect 6822 8412 6828 8424
rect 6564 8384 6828 8412
rect 6365 8375 6423 8381
rect 6822 8372 6828 8384
rect 6880 8412 6886 8424
rect 7009 8415 7067 8421
rect 7009 8412 7021 8415
rect 6880 8384 7021 8412
rect 6880 8372 6886 8384
rect 7009 8381 7021 8384
rect 7055 8381 7067 8415
rect 7009 8375 7067 8381
rect 7834 8372 7840 8424
rect 7892 8412 7898 8424
rect 8205 8415 8263 8421
rect 8205 8412 8217 8415
rect 7892 8384 8217 8412
rect 7892 8372 7898 8384
rect 8205 8381 8217 8384
rect 8251 8381 8263 8415
rect 8205 8375 8263 8381
rect 8478 8372 8484 8424
rect 8536 8372 8542 8424
rect 9600 8421 9628 8452
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 9674 8372 9680 8424
rect 9732 8372 9738 8424
rect 5500 8316 6132 8344
rect 6457 8347 6515 8353
rect 5500 8304 5506 8316
rect 6457 8313 6469 8347
rect 6503 8344 6515 8347
rect 9861 8347 9919 8353
rect 6503 8316 9812 8344
rect 6503 8313 6515 8316
rect 6457 8307 6515 8313
rect 4798 8276 4804 8288
rect 4172 8248 4804 8276
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 6822 8236 6828 8288
rect 6880 8236 6886 8288
rect 8018 8236 8024 8288
rect 8076 8236 8082 8288
rect 9784 8276 9812 8316
rect 9861 8313 9873 8347
rect 9907 8344 9919 8347
rect 9968 8344 9996 8520
rect 13464 8480 13492 8576
rect 13556 8548 13584 8576
rect 14737 8551 14795 8557
rect 13556 8520 13676 8548
rect 13280 8452 13492 8480
rect 13280 8421 13308 8452
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8381 13323 8415
rect 13265 8375 13323 8381
rect 13354 8372 13360 8424
rect 13412 8372 13418 8424
rect 13648 8421 13676 8520
rect 14737 8517 14749 8551
rect 14783 8548 14795 8551
rect 14826 8548 14832 8560
rect 14783 8520 14832 8548
rect 14783 8517 14795 8520
rect 14737 8511 14795 8517
rect 14826 8508 14832 8520
rect 14884 8508 14890 8560
rect 13633 8415 13691 8421
rect 13633 8381 13645 8415
rect 13679 8412 13691 8415
rect 14185 8415 14243 8421
rect 14185 8412 14197 8415
rect 13679 8384 14197 8412
rect 13679 8381 13691 8384
rect 13633 8375 13691 8381
rect 14185 8381 14197 8384
rect 14231 8412 14243 8415
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14231 8384 14933 8412
rect 14231 8381 14243 8384
rect 14185 8375 14243 8381
rect 14921 8381 14933 8384
rect 14967 8381 14979 8415
rect 14921 8375 14979 8381
rect 15105 8415 15163 8421
rect 15105 8381 15117 8415
rect 15151 8381 15163 8415
rect 15105 8375 15163 8381
rect 10962 8344 10968 8356
rect 9907 8316 10968 8344
rect 9907 8313 9919 8316
rect 9861 8307 9919 8313
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 14369 8347 14427 8353
rect 14369 8344 14381 8347
rect 11072 8316 14381 8344
rect 11072 8276 11100 8316
rect 14369 8313 14381 8316
rect 14415 8344 14427 8347
rect 15010 8344 15016 8356
rect 14415 8316 15016 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 15010 8304 15016 8316
rect 15068 8344 15074 8356
rect 15120 8344 15148 8375
rect 15068 8316 15148 8344
rect 15068 8304 15074 8316
rect 9784 8248 11100 8276
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 13538 8276 13544 8288
rect 13320 8248 13544 8276
rect 13320 8236 13326 8248
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 92 8186 15824 8208
rect 92 8134 2564 8186
rect 2616 8134 2628 8186
rect 2680 8134 2692 8186
rect 2744 8134 2756 8186
rect 2808 8134 2820 8186
rect 2872 8134 6497 8186
rect 6549 8134 6561 8186
rect 6613 8134 6625 8186
rect 6677 8134 6689 8186
rect 6741 8134 6753 8186
rect 6805 8134 10430 8186
rect 10482 8134 10494 8186
rect 10546 8134 10558 8186
rect 10610 8134 10622 8186
rect 10674 8134 10686 8186
rect 10738 8134 14363 8186
rect 14415 8134 14427 8186
rect 14479 8134 14491 8186
rect 14543 8134 14555 8186
rect 14607 8134 14619 8186
rect 14671 8134 15824 8186
rect 92 8112 15824 8134
rect 2314 8072 2320 8084
rect 1044 8044 2320 8072
rect 1044 8013 1072 8044
rect 2314 8032 2320 8044
rect 2372 8032 2378 8084
rect 3050 8032 3056 8084
rect 3108 8032 3114 8084
rect 6362 8032 6368 8084
rect 6420 8032 6426 8084
rect 8018 8072 8024 8084
rect 7116 8044 8024 8072
rect 1029 8007 1087 8013
rect 1029 8004 1041 8007
rect 676 7976 1041 8004
rect 676 7945 704 7976
rect 1029 7973 1041 7976
rect 1075 7973 1087 8007
rect 1029 7967 1087 7973
rect 1213 8007 1271 8013
rect 1213 7973 1225 8007
rect 1259 8004 1271 8007
rect 2038 8004 2044 8016
rect 1259 7976 2044 8004
rect 1259 7973 1271 7976
rect 1213 7967 1271 7973
rect 2038 7964 2044 7976
rect 2096 8004 2102 8016
rect 2409 8007 2467 8013
rect 2409 8004 2421 8007
rect 2096 7976 2421 8004
rect 2096 7964 2102 7976
rect 2409 7973 2421 7976
rect 2455 7973 2467 8007
rect 3418 8004 3424 8016
rect 2409 7967 2467 7973
rect 2746 7976 3424 8004
rect 661 7939 719 7945
rect 661 7905 673 7939
rect 707 7905 719 7939
rect 661 7899 719 7905
rect 753 7939 811 7945
rect 753 7905 765 7939
rect 799 7905 811 7939
rect 753 7899 811 7905
rect 937 7939 995 7945
rect 937 7905 949 7939
rect 983 7936 995 7939
rect 1305 7939 1363 7945
rect 983 7908 1164 7936
rect 983 7905 995 7908
rect 937 7899 995 7905
rect 768 7868 796 7899
rect 1136 7880 1164 7908
rect 1305 7905 1317 7939
rect 1351 7905 1363 7939
rect 1305 7899 1363 7905
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1486 7936 1492 7948
rect 1443 7908 1492 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 768 7840 1072 7868
rect 1044 7809 1072 7840
rect 1118 7828 1124 7880
rect 1176 7828 1182 7880
rect 1320 7868 1348 7899
rect 1486 7896 1492 7908
rect 1544 7896 1550 7948
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7905 1823 7939
rect 1765 7899 1823 7905
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2222 7936 2228 7948
rect 2179 7908 2228 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 1578 7868 1584 7880
rect 1320 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 1780 7812 1808 7899
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7905 2375 7939
rect 2317 7899 2375 7905
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7936 2559 7939
rect 2746 7936 2774 7976
rect 3418 7964 3424 7976
rect 3476 8004 3482 8016
rect 5721 8007 5779 8013
rect 5721 8004 5733 8007
rect 3476 7976 5733 8004
rect 3476 7964 3482 7976
rect 5721 7973 5733 7976
rect 5767 7973 5779 8007
rect 5721 7967 5779 7973
rect 2547 7908 2774 7936
rect 2547 7905 2559 7908
rect 2501 7899 2559 7905
rect 2332 7868 2360 7899
rect 2958 7896 2964 7948
rect 3016 7896 3022 7948
rect 4430 7896 4436 7948
rect 4488 7936 4494 7948
rect 4525 7939 4583 7945
rect 4525 7936 4537 7939
rect 4488 7908 4537 7936
rect 4488 7896 4494 7908
rect 4525 7905 4537 7908
rect 4571 7905 4583 7939
rect 4525 7899 4583 7905
rect 4798 7896 4804 7948
rect 4856 7896 4862 7948
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 5684 7908 6285 7936
rect 5684 7896 5690 7908
rect 6273 7905 6285 7908
rect 6319 7905 6331 7939
rect 6380 7936 6408 8032
rect 7116 8013 7144 8044
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 8478 8032 8484 8084
rect 8536 8072 8542 8084
rect 8573 8075 8631 8081
rect 8573 8072 8585 8075
rect 8536 8044 8585 8072
rect 8536 8032 8542 8044
rect 8573 8041 8585 8044
rect 8619 8041 8631 8075
rect 8573 8035 8631 8041
rect 9398 8032 9404 8084
rect 9456 8032 9462 8084
rect 9569 8075 9627 8081
rect 9569 8072 9581 8075
rect 9508 8044 9581 8072
rect 7101 8007 7159 8013
rect 7101 7973 7113 8007
rect 7147 7973 7159 8007
rect 7101 7967 7159 7973
rect 6825 7939 6883 7945
rect 6825 7936 6837 7939
rect 6380 7908 6837 7936
rect 6273 7899 6331 7905
rect 6825 7905 6837 7908
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 2976 7868 3004 7896
rect 2332 7840 3004 7868
rect 6288 7868 6316 7899
rect 8220 7868 8248 7922
rect 8662 7896 8668 7948
rect 8720 7896 8726 7948
rect 8849 7939 8907 7945
rect 8849 7905 8861 7939
rect 8895 7936 8907 7939
rect 9508 7936 9536 8044
rect 9569 8041 9581 8044
rect 9615 8072 9627 8075
rect 10045 8075 10103 8081
rect 9615 8044 9996 8072
rect 9615 8041 9627 8044
rect 9569 8035 9627 8041
rect 9769 8007 9827 8013
rect 9769 8004 9781 8007
rect 9692 7976 9781 8004
rect 9692 7948 9720 7976
rect 9769 7973 9781 7976
rect 9815 7973 9827 8007
rect 9968 8004 9996 8044
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 10134 8072 10140 8084
rect 10091 8044 10140 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 15010 8032 15016 8084
rect 15068 8072 15074 8084
rect 15289 8075 15347 8081
rect 15289 8072 15301 8075
rect 15068 8044 15301 8072
rect 15068 8032 15074 8044
rect 15289 8041 15301 8044
rect 15335 8041 15347 8075
rect 15289 8035 15347 8041
rect 9968 7976 10180 8004
rect 9769 7967 9827 7973
rect 8895 7908 9536 7936
rect 8895 7905 8907 7908
rect 8849 7899 8907 7905
rect 9674 7896 9680 7948
rect 9732 7934 9738 7948
rect 10152 7945 10180 7976
rect 13078 7964 13084 8016
rect 13136 7964 13142 8016
rect 9861 7939 9919 7945
rect 9861 7936 9873 7939
rect 9784 7934 9873 7936
rect 9732 7908 9873 7934
rect 9732 7906 9812 7908
rect 9732 7896 9738 7906
rect 9861 7905 9873 7908
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7936 10195 7939
rect 10318 7936 10324 7948
rect 10183 7908 10324 7936
rect 10183 7905 10195 7908
rect 10137 7899 10195 7905
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7936 11023 7939
rect 11011 7908 11192 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 6288 7840 6868 7868
rect 6840 7812 6868 7840
rect 6932 7840 8248 7868
rect 1029 7803 1087 7809
rect 1029 7769 1041 7803
rect 1075 7769 1087 7803
rect 1029 7763 1087 7769
rect 1762 7760 1768 7812
rect 1820 7800 1826 7812
rect 1820 7772 5028 7800
rect 1820 7760 1826 7772
rect 5000 7744 5028 7772
rect 6822 7760 6828 7812
rect 6880 7760 6886 7812
rect 474 7692 480 7744
rect 532 7692 538 7744
rect 750 7692 756 7744
rect 808 7692 814 7744
rect 2682 7692 2688 7744
rect 2740 7692 2746 7744
rect 3234 7692 3240 7744
rect 3292 7732 3298 7744
rect 4617 7735 4675 7741
rect 4617 7732 4629 7735
rect 3292 7704 4629 7732
rect 3292 7692 3298 7704
rect 4617 7701 4629 7704
rect 4663 7701 4675 7735
rect 4617 7695 4675 7701
rect 4982 7692 4988 7744
rect 5040 7692 5046 7744
rect 5074 7692 5080 7744
rect 5132 7732 5138 7744
rect 6932 7732 6960 7840
rect 8938 7828 8944 7880
rect 8996 7868 9002 7880
rect 10796 7868 10824 7899
rect 8996 7840 10824 7868
rect 8996 7828 9002 7840
rect 11164 7812 11192 7908
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 11885 7939 11943 7945
rect 11885 7936 11897 7939
rect 11756 7908 11897 7936
rect 11756 7896 11762 7908
rect 11885 7905 11897 7908
rect 11931 7905 11943 7939
rect 11885 7899 11943 7905
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 14645 7939 14703 7945
rect 14645 7936 14657 7939
rect 14240 7908 14657 7936
rect 14240 7896 14246 7908
rect 14645 7905 14657 7908
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 15378 7896 15384 7948
rect 15436 7896 15442 7948
rect 12250 7828 12256 7880
rect 12308 7828 12314 7880
rect 14734 7828 14740 7880
rect 14792 7828 14798 7880
rect 9858 7760 9864 7812
rect 9916 7760 9922 7812
rect 11146 7760 11152 7812
rect 11204 7760 11210 7812
rect 13679 7803 13737 7809
rect 13679 7800 13691 7803
rect 13464 7772 13691 7800
rect 13464 7744 13492 7772
rect 13679 7769 13691 7772
rect 13725 7769 13737 7803
rect 13679 7763 13737 7769
rect 5132 7704 6960 7732
rect 5132 7692 5138 7704
rect 7834 7692 7840 7744
rect 7892 7732 7898 7744
rect 8757 7735 8815 7741
rect 8757 7732 8769 7735
rect 7892 7704 8769 7732
rect 7892 7692 7898 7704
rect 8757 7701 8769 7704
rect 8803 7701 8815 7735
rect 8757 7695 8815 7701
rect 9585 7735 9643 7741
rect 9585 7701 9597 7735
rect 9631 7732 9643 7735
rect 10134 7732 10140 7744
rect 9631 7704 10140 7732
rect 9631 7701 9643 7704
rect 9585 7695 9643 7701
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 10873 7735 10931 7741
rect 10873 7701 10885 7735
rect 10919 7732 10931 7735
rect 13354 7732 13360 7744
rect 10919 7704 13360 7732
rect 10919 7701 10931 7704
rect 10873 7695 10931 7701
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 13446 7692 13452 7744
rect 13504 7692 13510 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 14369 7735 14427 7741
rect 14369 7732 14381 7735
rect 13596 7704 14381 7732
rect 13596 7692 13602 7704
rect 14369 7701 14381 7704
rect 14415 7701 14427 7735
rect 14369 7695 14427 7701
rect 92 7642 15824 7664
rect 92 7590 1904 7642
rect 1956 7590 1968 7642
rect 2020 7590 2032 7642
rect 2084 7590 2096 7642
rect 2148 7590 2160 7642
rect 2212 7590 5837 7642
rect 5889 7590 5901 7642
rect 5953 7590 5965 7642
rect 6017 7590 6029 7642
rect 6081 7590 6093 7642
rect 6145 7590 9770 7642
rect 9822 7590 9834 7642
rect 9886 7590 9898 7642
rect 9950 7590 9962 7642
rect 10014 7590 10026 7642
rect 10078 7590 13703 7642
rect 13755 7590 13767 7642
rect 13819 7590 13831 7642
rect 13883 7590 13895 7642
rect 13947 7590 13959 7642
rect 14011 7590 15824 7642
rect 92 7568 15824 7590
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 2314 7528 2320 7540
rect 2179 7500 2320 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 2314 7488 2320 7500
rect 2372 7488 2378 7540
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 3034 7531 3092 7537
rect 3034 7528 3046 7531
rect 2740 7500 3046 7528
rect 2740 7488 2746 7500
rect 3034 7497 3046 7500
rect 3080 7497 3092 7531
rect 3034 7491 3092 7497
rect 5169 7531 5227 7537
rect 5169 7497 5181 7531
rect 5215 7528 5227 7531
rect 5350 7528 5356 7540
rect 5215 7500 5356 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 5350 7488 5356 7500
rect 5408 7528 5414 7540
rect 5718 7528 5724 7540
rect 5408 7500 5724 7528
rect 5408 7488 5414 7500
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 13081 7531 13139 7537
rect 13081 7528 13093 7531
rect 12308 7500 13093 7528
rect 12308 7488 12314 7500
rect 13081 7497 13093 7500
rect 13127 7497 13139 7531
rect 13081 7491 13139 7497
rect 13538 7488 13544 7540
rect 13596 7488 13602 7540
rect 14182 7488 14188 7540
rect 14240 7488 14246 7540
rect 14734 7488 14740 7540
rect 14792 7528 14798 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 14792 7500 15301 7528
rect 14792 7488 14798 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 5629 7463 5687 7469
rect 5629 7460 5641 7463
rect 5592 7432 5641 7460
rect 5592 7420 5598 7432
rect 5629 7429 5641 7432
rect 5675 7429 5687 7463
rect 13556 7460 13584 7488
rect 5629 7423 5687 7429
rect 13280 7432 13584 7460
rect 661 7395 719 7401
rect 661 7361 673 7395
rect 707 7392 719 7395
rect 750 7392 756 7404
rect 707 7364 756 7392
rect 707 7361 719 7364
rect 661 7355 719 7361
rect 750 7352 756 7364
rect 808 7352 814 7404
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 3602 7392 3608 7404
rect 2823 7364 3608 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 3602 7352 3608 7364
rect 3660 7392 3666 7404
rect 4522 7392 4528 7404
rect 3660 7364 4528 7392
rect 3660 7352 3666 7364
rect 4522 7352 4528 7364
rect 4580 7392 4586 7404
rect 5997 7395 6055 7401
rect 5997 7392 6009 7395
rect 4580 7364 6009 7392
rect 4580 7352 4586 7364
rect 5997 7361 6009 7364
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 11698 7352 11704 7404
rect 11756 7392 11762 7404
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 11756 7364 12081 7392
rect 11756 7352 11762 7364
rect 12069 7361 12081 7364
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 382 7284 388 7336
rect 440 7284 446 7336
rect 1486 7148 1492 7200
rect 1544 7188 1550 7200
rect 1780 7188 1808 7310
rect 4982 7284 4988 7336
rect 5040 7284 5046 7336
rect 5074 7284 5080 7336
rect 5132 7284 5138 7336
rect 5442 7284 5448 7336
rect 5500 7284 5506 7336
rect 5626 7284 5632 7336
rect 5684 7284 5690 7336
rect 7742 7324 7748 7336
rect 7406 7296 7748 7324
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 13280 7333 13308 7432
rect 13906 7420 13912 7472
rect 13964 7460 13970 7472
rect 14001 7463 14059 7469
rect 14001 7460 14013 7463
rect 13964 7432 14013 7460
rect 13964 7420 13970 7432
rect 14001 7429 14013 7432
rect 14047 7429 14059 7463
rect 14200 7460 14228 7488
rect 14001 7423 14059 7429
rect 14108 7432 14228 7460
rect 13538 7352 13544 7404
rect 13596 7352 13602 7404
rect 13265 7327 13323 7333
rect 13265 7293 13277 7327
rect 13311 7293 13323 7327
rect 13265 7287 13323 7293
rect 13354 7284 13360 7336
rect 13412 7284 13418 7336
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 13633 7327 13691 7333
rect 13633 7324 13645 7327
rect 13504 7296 13645 7324
rect 13504 7284 13510 7296
rect 13633 7293 13645 7296
rect 13679 7324 13691 7327
rect 13725 7327 13783 7333
rect 13725 7324 13737 7327
rect 13679 7296 13737 7324
rect 13679 7293 13691 7296
rect 13633 7287 13691 7293
rect 13725 7293 13737 7296
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 13909 7327 13967 7333
rect 13909 7293 13921 7327
rect 13955 7324 13967 7327
rect 13998 7324 14004 7336
rect 13955 7296 14004 7324
rect 13955 7293 13967 7296
rect 13909 7287 13967 7293
rect 4338 7256 4344 7268
rect 4278 7228 4344 7256
rect 4338 7216 4344 7228
rect 4396 7256 4402 7268
rect 5092 7256 5120 7284
rect 4396 7228 5120 7256
rect 4396 7216 4402 7228
rect 6270 7216 6276 7268
rect 6328 7216 6334 7268
rect 7926 7216 7932 7268
rect 7984 7216 7990 7268
rect 10778 7216 10784 7268
rect 10836 7216 10842 7268
rect 11514 7216 11520 7268
rect 11572 7256 11578 7268
rect 11793 7259 11851 7265
rect 11793 7256 11805 7259
rect 11572 7228 11805 7256
rect 11572 7216 11578 7228
rect 11793 7225 11805 7228
rect 11839 7225 11851 7259
rect 13740 7256 13768 7287
rect 13998 7284 14004 7296
rect 14056 7284 14062 7336
rect 14108 7324 14136 7432
rect 14185 7395 14243 7401
rect 14185 7361 14197 7395
rect 14231 7392 14243 7395
rect 15105 7395 15163 7401
rect 15105 7392 15117 7395
rect 14231 7364 15117 7392
rect 14231 7361 14243 7364
rect 14185 7355 14243 7361
rect 15105 7361 15117 7364
rect 15151 7392 15163 7395
rect 15151 7364 15240 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 14108 7296 14289 7324
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 15010 7324 15016 7336
rect 14967 7296 15016 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 15212 7333 15240 7364
rect 15197 7327 15255 7333
rect 15197 7293 15209 7327
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 15381 7327 15439 7333
rect 15381 7293 15393 7327
rect 15427 7293 15439 7327
rect 15381 7287 15439 7293
rect 14737 7259 14795 7265
rect 14737 7256 14749 7259
rect 13740 7228 14749 7256
rect 11793 7219 11851 7225
rect 14737 7225 14749 7228
rect 14783 7225 14795 7259
rect 14737 7219 14795 7225
rect 1544 7160 1808 7188
rect 1544 7148 1550 7160
rect 2222 7148 2228 7200
rect 2280 7188 2286 7200
rect 2958 7188 2964 7200
rect 2280 7160 2964 7188
rect 2280 7148 2286 7160
rect 2958 7148 2964 7160
rect 3016 7188 3022 7200
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 3016 7160 4537 7188
rect 3016 7148 3022 7160
rect 4525 7157 4537 7160
rect 4571 7157 4583 7191
rect 4525 7151 4583 7157
rect 7742 7148 7748 7200
rect 7800 7148 7806 7200
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 8260 7160 9229 7188
rect 8260 7148 8266 7160
rect 9217 7157 9229 7160
rect 9263 7157 9275 7191
rect 9217 7151 9275 7157
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10321 7191 10379 7197
rect 10321 7188 10333 7191
rect 9916 7160 10333 7188
rect 9916 7148 9922 7160
rect 10321 7157 10333 7160
rect 10367 7157 10379 7191
rect 10321 7151 10379 7157
rect 13909 7191 13967 7197
rect 13909 7157 13921 7191
rect 13955 7188 13967 7191
rect 14645 7191 14703 7197
rect 14645 7188 14657 7191
rect 13955 7160 14657 7188
rect 13955 7157 13967 7160
rect 13909 7151 13967 7157
rect 14645 7157 14657 7160
rect 14691 7188 14703 7191
rect 15396 7188 15424 7287
rect 14691 7160 15424 7188
rect 14691 7157 14703 7160
rect 14645 7151 14703 7157
rect 92 7098 15824 7120
rect 92 7046 2564 7098
rect 2616 7046 2628 7098
rect 2680 7046 2692 7098
rect 2744 7046 2756 7098
rect 2808 7046 2820 7098
rect 2872 7046 6497 7098
rect 6549 7046 6561 7098
rect 6613 7046 6625 7098
rect 6677 7046 6689 7098
rect 6741 7046 6753 7098
rect 6805 7046 10430 7098
rect 10482 7046 10494 7098
rect 10546 7046 10558 7098
rect 10610 7046 10622 7098
rect 10674 7046 10686 7098
rect 10738 7046 14363 7098
rect 14415 7046 14427 7098
rect 14479 7046 14491 7098
rect 14543 7046 14555 7098
rect 14607 7046 14619 7098
rect 14671 7046 15824 7098
rect 92 7024 15824 7046
rect 1486 6944 1492 6996
rect 1544 6984 1550 6996
rect 4338 6984 4344 6996
rect 1544 6956 4344 6984
rect 1544 6944 1550 6956
rect 4338 6944 4344 6956
rect 4396 6944 4402 6996
rect 6270 6944 6276 6996
rect 6328 6984 6334 6996
rect 6457 6987 6515 6993
rect 6457 6984 6469 6987
rect 6328 6956 6469 6984
rect 6328 6944 6334 6956
rect 6457 6953 6469 6956
rect 6503 6953 6515 6987
rect 6457 6947 6515 6953
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 9769 6987 9827 6993
rect 9769 6984 9781 6987
rect 9272 6956 9781 6984
rect 9272 6944 9278 6956
rect 9769 6953 9781 6956
rect 9815 6953 9827 6987
rect 9769 6947 9827 6953
rect 9861 6987 9919 6993
rect 9861 6953 9873 6987
rect 9907 6984 9919 6987
rect 10318 6984 10324 6996
rect 9907 6956 10324 6984
rect 9907 6953 9919 6956
rect 9861 6947 9919 6953
rect 10318 6944 10324 6956
rect 10376 6944 10382 6996
rect 13998 6944 14004 6996
rect 14056 6984 14062 6996
rect 15010 6984 15016 6996
rect 14056 6956 15016 6984
rect 14056 6944 14062 6956
rect 15010 6944 15016 6956
rect 15068 6944 15074 6996
rect 8573 6919 8631 6925
rect 8573 6885 8585 6919
rect 8619 6916 8631 6919
rect 8938 6916 8944 6928
rect 8619 6888 8944 6916
rect 8619 6885 8631 6888
rect 8573 6879 8631 6885
rect 8938 6876 8944 6888
rect 8996 6876 9002 6928
rect 661 6851 719 6857
rect 661 6817 673 6851
rect 707 6848 719 6851
rect 1302 6848 1308 6860
rect 707 6820 1308 6848
rect 707 6817 719 6820
rect 661 6811 719 6817
rect 1302 6808 1308 6820
rect 1360 6808 1366 6860
rect 1670 6808 1676 6860
rect 1728 6808 1734 6860
rect 4154 6808 4160 6860
rect 4212 6808 4218 6860
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6848 6699 6851
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 6687 6820 7665 6848
rect 6687 6817 6699 6820
rect 6641 6811 6699 6817
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 7742 6808 7748 6860
rect 7800 6808 7806 6860
rect 7834 6808 7840 6860
rect 7892 6808 7898 6860
rect 8478 6808 8484 6860
rect 8536 6848 8542 6860
rect 8665 6851 8723 6857
rect 8665 6848 8677 6851
rect 8536 6820 8677 6848
rect 8536 6808 8542 6820
rect 8665 6817 8677 6820
rect 8711 6817 8723 6851
rect 8665 6811 8723 6817
rect 9033 6851 9091 6857
rect 9033 6817 9045 6851
rect 9079 6848 9091 6851
rect 9309 6851 9367 6857
rect 9079 6820 9168 6848
rect 9079 6817 9091 6820
rect 9033 6811 9091 6817
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 5442 6780 5448 6792
rect 4304 6752 5448 6780
rect 4304 6740 4310 6752
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 7760 6780 7788 6808
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7760 6752 8033 6780
rect 8021 6749 8033 6752
rect 8067 6780 8079 6783
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 8067 6752 8309 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 9140 6780 9168 6820
rect 9309 6817 9321 6851
rect 9355 6848 9367 6851
rect 9355 6820 10088 6848
rect 9355 6817 9367 6820
rect 9309 6811 9367 6817
rect 9858 6780 9864 6792
rect 9140 6752 9864 6780
rect 9140 6724 9168 6752
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10060 6789 10088 6820
rect 10962 6808 10968 6860
rect 11020 6808 11026 6860
rect 11146 6808 11152 6860
rect 11204 6808 11210 6860
rect 11333 6851 11391 6857
rect 11333 6817 11345 6851
rect 11379 6848 11391 6851
rect 11422 6848 11428 6860
rect 11379 6820 11428 6848
rect 11379 6817 11391 6820
rect 11333 6811 11391 6817
rect 11422 6808 11428 6820
rect 11480 6848 11486 6860
rect 13262 6848 13268 6860
rect 11480 6820 13268 6848
rect 11480 6808 11486 6820
rect 13262 6808 13268 6820
rect 13320 6848 13326 6860
rect 13538 6848 13544 6860
rect 13320 6820 13544 6848
rect 13320 6808 13326 6820
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 13906 6808 13912 6860
rect 13964 6848 13970 6860
rect 14090 6848 14096 6860
rect 13964 6820 14096 6848
rect 13964 6808 13970 6820
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 15286 6808 15292 6860
rect 15344 6808 15350 6860
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6780 10103 6783
rect 10134 6780 10140 6792
rect 10091 6752 10140 6780
rect 10091 6749 10103 6752
rect 10045 6743 10103 6749
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10980 6780 11008 6808
rect 10980 6752 11376 6780
rect 11348 6724 11376 6752
rect 3160 6684 8064 6712
rect 3160 6656 3188 6684
rect 8036 6656 8064 6684
rect 9122 6672 9128 6724
rect 9180 6672 9186 6724
rect 11330 6672 11336 6724
rect 11388 6672 11394 6724
rect 474 6604 480 6656
rect 532 6604 538 6656
rect 1394 6604 1400 6656
rect 1452 6644 1458 6656
rect 1489 6647 1547 6653
rect 1489 6644 1501 6647
rect 1452 6616 1501 6644
rect 1452 6604 1458 6616
rect 1489 6613 1501 6616
rect 1535 6613 1547 6647
rect 1489 6607 1547 6613
rect 3142 6604 3148 6656
rect 3200 6604 3206 6656
rect 4338 6604 4344 6656
rect 4396 6604 4402 6656
rect 8018 6604 8024 6656
rect 8076 6604 8082 6656
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 8904 6616 9413 6644
rect 8904 6604 8910 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9401 6607 9459 6613
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 14642 6644 14648 6656
rect 9548 6616 14648 6644
rect 9548 6604 9554 6616
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 15470 6604 15476 6656
rect 15528 6604 15534 6656
rect 92 6554 15824 6576
rect 92 6502 1904 6554
rect 1956 6502 1968 6554
rect 2020 6502 2032 6554
rect 2084 6502 2096 6554
rect 2148 6502 2160 6554
rect 2212 6502 5837 6554
rect 5889 6502 5901 6554
rect 5953 6502 5965 6554
rect 6017 6502 6029 6554
rect 6081 6502 6093 6554
rect 6145 6502 9770 6554
rect 9822 6502 9834 6554
rect 9886 6502 9898 6554
rect 9950 6502 9962 6554
rect 10014 6502 10026 6554
rect 10078 6502 13703 6554
rect 13755 6502 13767 6554
rect 13819 6502 13831 6554
rect 13883 6502 13895 6554
rect 13947 6502 13959 6554
rect 14011 6502 15824 6554
rect 92 6480 15824 6502
rect 1670 6400 1676 6452
rect 1728 6440 1734 6452
rect 2225 6443 2283 6449
rect 2225 6440 2237 6443
rect 1728 6412 2237 6440
rect 1728 6400 1734 6412
rect 2225 6409 2237 6412
rect 2271 6409 2283 6443
rect 2958 6440 2964 6452
rect 2225 6403 2283 6409
rect 2746 6412 2964 6440
rect 382 6264 388 6316
rect 440 6264 446 6316
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1360 6276 2145 6304
rect 1360 6264 1366 6276
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 1762 6196 1768 6248
rect 1820 6196 1826 6248
rect 658 6128 664 6180
rect 716 6128 722 6180
rect 2148 6100 2176 6267
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 2332 6208 2605 6236
rect 2332 6180 2360 6208
rect 2593 6205 2605 6208
rect 2639 6236 2651 6239
rect 2746 6236 2774 6412
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 4065 6443 4123 6449
rect 4065 6409 4077 6443
rect 4111 6440 4123 6443
rect 4154 6440 4160 6452
rect 4111 6412 4160 6440
rect 4111 6409 4123 6412
rect 4065 6403 4123 6409
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 4506 6443 4564 6449
rect 4506 6440 4518 6443
rect 4396 6412 4518 6440
rect 4396 6400 4402 6412
rect 4506 6409 4518 6412
rect 4552 6409 4564 6443
rect 4506 6403 4564 6409
rect 6178 6400 6184 6452
rect 6236 6440 6242 6452
rect 6273 6443 6331 6449
rect 6273 6440 6285 6443
rect 6236 6412 6285 6440
rect 6236 6400 6242 6412
rect 6273 6409 6285 6412
rect 6319 6409 6331 6443
rect 6273 6403 6331 6409
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 8720 6412 8769 6440
rect 8720 6400 8726 6412
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 9490 6440 9496 6452
rect 8757 6403 8815 6409
rect 8864 6412 9496 6440
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 5997 6375 6055 6381
rect 5997 6372 6009 6375
rect 5592 6344 6009 6372
rect 5592 6332 5598 6344
rect 5997 6341 6009 6344
rect 6043 6372 6055 6375
rect 8864 6372 8892 6412
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 10962 6400 10968 6452
rect 11020 6440 11026 6452
rect 12710 6440 12716 6452
rect 11020 6412 12716 6440
rect 11020 6400 11026 6412
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 15197 6443 15255 6449
rect 15197 6409 15209 6443
rect 15243 6440 15255 6443
rect 15286 6440 15292 6452
rect 15243 6412 15292 6440
rect 15243 6409 15255 6412
rect 15197 6403 15255 6409
rect 15286 6400 15292 6412
rect 15344 6400 15350 6452
rect 13633 6375 13691 6381
rect 6043 6344 8892 6372
rect 9048 6344 10180 6372
rect 6043 6341 6055 6344
rect 5997 6335 6055 6341
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6304 4307 6307
rect 4522 6304 4528 6316
rect 4295 6276 4528 6304
rect 4295 6273 4307 6276
rect 4249 6267 4307 6273
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 5718 6304 5724 6316
rect 5644 6276 5724 6304
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 2639 6208 3433 6236
rect 2639 6205 2651 6208
rect 2593 6199 2651 6205
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3421 6199 3479 6205
rect 3602 6196 3608 6248
rect 3660 6196 3666 6248
rect 5644 6222 5672 6276
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 9048 6313 9076 6344
rect 10152 6316 10180 6344
rect 13633 6341 13645 6375
rect 13679 6341 13691 6375
rect 13633 6335 13691 6341
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8536 6276 8953 6304
rect 8536 6264 8542 6276
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 9122 6264 9128 6316
rect 9180 6264 9186 6316
rect 10134 6264 10140 6316
rect 10192 6264 10198 6316
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11238 6304 11244 6316
rect 11011 6276 11244 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 11238 6264 11244 6276
rect 11296 6304 11302 6316
rect 11698 6304 11704 6316
rect 11296 6276 11704 6304
rect 11296 6264 11302 6276
rect 11698 6264 11704 6276
rect 11756 6304 11762 6316
rect 11974 6304 11980 6316
rect 11756 6276 11980 6304
rect 11756 6264 11762 6276
rect 11974 6264 11980 6276
rect 12032 6264 12038 6316
rect 13357 6307 13415 6313
rect 13357 6273 13369 6307
rect 13403 6304 13415 6307
rect 13538 6304 13544 6316
rect 13403 6276 13544 6304
rect 13403 6273 13415 6276
rect 13357 6267 13415 6273
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 13648 6304 13676 6335
rect 14642 6332 14648 6384
rect 14700 6332 14706 6384
rect 14001 6307 14059 6313
rect 14001 6304 14013 6307
rect 13648 6276 14013 6304
rect 14001 6273 14013 6276
rect 14047 6273 14059 6307
rect 14001 6267 14059 6273
rect 6086 6196 6092 6248
rect 6144 6196 6150 6248
rect 6273 6239 6331 6245
rect 6273 6236 6285 6239
rect 6196 6208 6285 6236
rect 6196 6180 6224 6208
rect 6273 6205 6285 6208
rect 6319 6236 6331 6239
rect 6822 6236 6828 6248
rect 6319 6208 6828 6236
rect 6319 6205 6331 6208
rect 6273 6199 6331 6205
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 9214 6196 9220 6248
rect 9272 6196 9278 6248
rect 9398 6196 9404 6248
rect 9456 6196 9462 6248
rect 9585 6239 9643 6245
rect 9585 6205 9597 6239
rect 9631 6205 9643 6239
rect 9585 6199 9643 6205
rect 9769 6239 9827 6245
rect 9769 6205 9781 6239
rect 9815 6236 9827 6239
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9815 6208 9965 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 2314 6128 2320 6180
rect 2372 6128 2378 6180
rect 2409 6171 2467 6177
rect 2409 6137 2421 6171
rect 2455 6137 2467 6171
rect 2409 6131 2467 6137
rect 2424 6100 2452 6131
rect 3694 6128 3700 6180
rect 3752 6128 3758 6180
rect 3881 6171 3939 6177
rect 3881 6137 3893 6171
rect 3927 6168 3939 6171
rect 4154 6168 4160 6180
rect 3927 6140 4160 6168
rect 3927 6137 3939 6140
rect 3881 6131 3939 6137
rect 4154 6128 4160 6140
rect 4212 6128 4218 6180
rect 6178 6128 6184 6180
rect 6236 6128 6242 6180
rect 8938 6128 8944 6180
rect 8996 6168 9002 6180
rect 9600 6168 9628 6199
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 13265 6239 13323 6245
rect 13265 6236 13277 6239
rect 12768 6208 13277 6236
rect 12768 6196 12774 6208
rect 13265 6205 13277 6208
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 14090 6196 14096 6248
rect 14148 6196 14154 6248
rect 15013 6239 15071 6245
rect 15013 6236 15025 6239
rect 14844 6208 15025 6236
rect 8996 6140 9628 6168
rect 10505 6171 10563 6177
rect 8996 6128 9002 6140
rect 10505 6137 10517 6171
rect 10551 6168 10563 6171
rect 10778 6168 10784 6180
rect 10551 6140 10784 6168
rect 10551 6137 10563 6140
rect 10505 6131 10563 6137
rect 2148 6072 2452 6100
rect 3513 6103 3571 6109
rect 3513 6069 3525 6103
rect 3559 6100 3571 6103
rect 5166 6100 5172 6112
rect 3559 6072 5172 6100
rect 3559 6069 3571 6072
rect 3513 6063 3571 6069
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 10520 6100 10548 6131
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 11241 6171 11299 6177
rect 11241 6137 11253 6171
rect 11287 6137 11299 6171
rect 12526 6168 12532 6180
rect 12466 6140 12532 6168
rect 11241 6131 11299 6137
rect 7340 6072 10548 6100
rect 11256 6100 11284 6131
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 14369 6171 14427 6177
rect 14369 6168 14381 6171
rect 12636 6140 14381 6168
rect 11422 6100 11428 6112
rect 11256 6072 11428 6100
rect 7340 6060 7346 6072
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 11974 6060 11980 6112
rect 12032 6100 12038 6112
rect 12636 6100 12664 6140
rect 14369 6137 14381 6140
rect 14415 6137 14427 6171
rect 14369 6131 14427 6137
rect 12032 6072 12664 6100
rect 12032 6060 12038 6072
rect 13722 6060 13728 6112
rect 13780 6060 13786 6112
rect 14844 6109 14872 6208
rect 15013 6205 15025 6208
rect 15059 6205 15071 6239
rect 15013 6199 15071 6205
rect 14829 6103 14887 6109
rect 14829 6069 14841 6103
rect 14875 6069 14887 6103
rect 14829 6063 14887 6069
rect 92 6010 15824 6032
rect 92 5958 2564 6010
rect 2616 5958 2628 6010
rect 2680 5958 2692 6010
rect 2744 5958 2756 6010
rect 2808 5958 2820 6010
rect 2872 5958 6497 6010
rect 6549 5958 6561 6010
rect 6613 5958 6625 6010
rect 6677 5958 6689 6010
rect 6741 5958 6753 6010
rect 6805 5958 10430 6010
rect 10482 5958 10494 6010
rect 10546 5958 10558 6010
rect 10610 5958 10622 6010
rect 10674 5958 10686 6010
rect 10738 5958 14363 6010
rect 14415 5958 14427 6010
rect 14479 5958 14491 6010
rect 14543 5958 14555 6010
rect 14607 5958 14619 6010
rect 14671 5958 15824 6010
rect 92 5936 15824 5958
rect 658 5856 664 5908
rect 716 5896 722 5908
rect 1121 5899 1179 5905
rect 1121 5896 1133 5899
rect 716 5868 1133 5896
rect 716 5856 722 5868
rect 1121 5865 1133 5868
rect 1167 5865 1179 5899
rect 1495 5899 1553 5905
rect 1495 5896 1507 5899
rect 1121 5859 1179 5865
rect 1228 5868 1507 5896
rect 753 5763 811 5769
rect 753 5729 765 5763
rect 799 5729 811 5763
rect 753 5723 811 5729
rect 768 5692 796 5723
rect 1026 5720 1032 5772
rect 1084 5720 1090 5772
rect 1228 5769 1256 5868
rect 1495 5865 1507 5868
rect 1541 5865 1553 5899
rect 1495 5859 1553 5865
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 2314 5896 2320 5908
rect 1627 5868 2320 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 4522 5896 4528 5908
rect 3283 5868 4528 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 1302 5788 1308 5840
rect 1360 5828 1366 5840
rect 1397 5831 1455 5837
rect 1397 5828 1409 5831
rect 1360 5800 1409 5828
rect 1360 5788 1366 5800
rect 1397 5797 1409 5800
rect 1443 5797 1455 5831
rect 1397 5791 1455 5797
rect 1213 5763 1271 5769
rect 1213 5729 1225 5763
rect 1259 5729 1271 5763
rect 1213 5723 1271 5729
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 1673 5763 1731 5769
rect 1673 5760 1685 5763
rect 1636 5732 1685 5760
rect 1636 5720 1642 5732
rect 1673 5729 1685 5732
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 3142 5692 3148 5704
rect 768 5664 3148 5692
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 1670 5624 1676 5636
rect 400 5596 1676 5624
rect 400 5568 428 5596
rect 1670 5584 1676 5596
rect 1728 5624 1734 5636
rect 3252 5624 3280 5859
rect 4522 5856 4528 5868
rect 4580 5856 4586 5908
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 5905 5899 5963 5905
rect 5905 5896 5917 5899
rect 5776 5868 5917 5896
rect 5776 5856 5782 5868
rect 5905 5865 5917 5868
rect 5951 5896 5963 5899
rect 6086 5896 6092 5908
rect 5951 5868 6092 5896
rect 5951 5865 5963 5868
rect 5905 5859 5963 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 9398 5896 9404 5908
rect 8720 5868 9404 5896
rect 8720 5856 8726 5868
rect 9398 5856 9404 5868
rect 9456 5896 9462 5908
rect 11146 5896 11152 5908
rect 9456 5868 11152 5896
rect 9456 5856 9462 5868
rect 11146 5856 11152 5868
rect 11204 5896 11210 5908
rect 11204 5868 11560 5896
rect 11204 5856 11210 5868
rect 4430 5788 4436 5840
rect 4488 5828 4494 5840
rect 8202 5828 8208 5840
rect 4488 5800 8208 5828
rect 4488 5788 4494 5800
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 9953 5831 10011 5837
rect 9953 5797 9965 5831
rect 9999 5828 10011 5831
rect 11238 5828 11244 5840
rect 9999 5800 11244 5828
rect 9999 5797 10011 5800
rect 9953 5791 10011 5797
rect 11238 5788 11244 5800
rect 11296 5788 11302 5840
rect 4154 5720 4160 5772
rect 4212 5720 4218 5772
rect 4448 5760 4476 5788
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 4448 5732 4537 5760
rect 4525 5729 4537 5732
rect 4571 5729 4583 5763
rect 4525 5723 4583 5729
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5760 4675 5763
rect 4706 5760 4712 5772
rect 4663 5732 4712 5760
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 4801 5763 4859 5769
rect 4801 5729 4813 5763
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 4985 5763 5043 5769
rect 4985 5729 4997 5763
rect 5031 5729 5043 5763
rect 4985 5723 5043 5729
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 5691 5763 5749 5769
rect 5691 5729 5703 5763
rect 5737 5760 5749 5763
rect 6178 5760 6184 5772
rect 5737 5732 6184 5760
rect 5737 5729 5749 5732
rect 5691 5723 5749 5729
rect 4172 5692 4200 5720
rect 4816 5692 4844 5723
rect 4172 5664 4844 5692
rect 5000 5692 5028 5723
rect 5074 5692 5080 5704
rect 5000 5664 5080 5692
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 5552 5692 5580 5723
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 7190 5760 7196 5772
rect 6288 5732 7196 5760
rect 6288 5692 6316 5732
rect 7190 5720 7196 5732
rect 7248 5760 7254 5772
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 7248 5732 7389 5760
rect 7248 5720 7254 5732
rect 7377 5729 7389 5732
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 7650 5720 7656 5772
rect 7708 5720 7714 5772
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 8110 5760 8116 5772
rect 7883 5732 8116 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 9732 5732 10057 5760
rect 9732 5720 9738 5732
rect 10045 5729 10057 5732
rect 10091 5729 10103 5763
rect 10045 5723 10103 5729
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 10689 5763 10747 5769
rect 10367 5732 10640 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 5552 5664 6316 5692
rect 1728 5596 3280 5624
rect 1728 5584 1734 5596
rect 3878 5584 3884 5636
rect 3936 5624 3942 5636
rect 5552 5624 5580 5664
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 10152 5692 10180 5723
rect 8904 5664 10180 5692
rect 8904 5652 8910 5664
rect 3936 5596 5580 5624
rect 7193 5627 7251 5633
rect 3936 5584 3942 5596
rect 7193 5593 7205 5627
rect 7239 5593 7251 5627
rect 10612 5624 10640 5732
rect 10689 5729 10701 5763
rect 10735 5760 10747 5763
rect 10778 5760 10784 5772
rect 10735 5732 10784 5760
rect 10735 5729 10747 5732
rect 10689 5723 10747 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 10870 5720 10876 5772
rect 10928 5720 10934 5772
rect 10962 5720 10968 5772
rect 11020 5720 11026 5772
rect 11057 5763 11115 5769
rect 11057 5729 11069 5763
rect 11103 5760 11115 5763
rect 11103 5732 11192 5760
rect 11103 5729 11115 5732
rect 11057 5723 11115 5729
rect 11164 5624 11192 5732
rect 11330 5720 11336 5772
rect 11388 5720 11394 5772
rect 11532 5769 11560 5868
rect 14826 5856 14832 5908
rect 14884 5856 14890 5908
rect 13078 5788 13084 5840
rect 13136 5828 13142 5840
rect 14844 5828 14872 5856
rect 13136 5800 14872 5828
rect 13136 5788 13142 5800
rect 11517 5763 11575 5769
rect 11517 5729 11529 5763
rect 11563 5729 11575 5763
rect 14921 5763 14979 5769
rect 14921 5760 14933 5763
rect 11517 5723 11575 5729
rect 14844 5732 14933 5760
rect 14844 5704 14872 5732
rect 14921 5729 14933 5732
rect 14967 5760 14979 5763
rect 15105 5763 15163 5769
rect 15105 5760 15117 5763
rect 14967 5732 15117 5760
rect 14967 5729 14979 5732
rect 14921 5723 14979 5729
rect 15105 5729 15117 5732
rect 15151 5729 15163 5763
rect 15105 5723 15163 5729
rect 14826 5652 14832 5704
rect 14884 5652 14890 5704
rect 10612 5596 11192 5624
rect 7193 5587 7251 5593
rect 382 5516 388 5568
rect 440 5516 446 5568
rect 474 5516 480 5568
rect 532 5516 538 5568
rect 3510 5516 3516 5568
rect 3568 5556 3574 5568
rect 4706 5556 4712 5568
rect 3568 5528 4712 5556
rect 3568 5516 3574 5528
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 4798 5516 4804 5568
rect 4856 5516 4862 5568
rect 5077 5559 5135 5565
rect 5077 5525 5089 5559
rect 5123 5556 5135 5559
rect 5442 5556 5448 5568
rect 5123 5528 5448 5556
rect 5123 5525 5135 5528
rect 5077 5519 5135 5525
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 7208 5556 7236 5587
rect 9214 5556 9220 5568
rect 5684 5528 9220 5556
rect 5684 5516 5690 5528
rect 9214 5516 9220 5528
rect 9272 5556 9278 5568
rect 9582 5556 9588 5568
rect 9272 5528 9588 5556
rect 9272 5516 9278 5528
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 10318 5516 10324 5568
rect 10376 5516 10382 5568
rect 11164 5556 11192 5596
rect 11241 5627 11299 5633
rect 11241 5593 11253 5627
rect 11287 5624 11299 5627
rect 11422 5624 11428 5636
rect 11287 5596 11428 5624
rect 11287 5593 11299 5596
rect 11241 5587 11299 5593
rect 11422 5584 11428 5596
rect 11480 5584 11486 5636
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 11164 5528 11345 5556
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 11333 5519 11391 5525
rect 15378 5516 15384 5568
rect 15436 5516 15442 5568
rect 92 5466 15824 5488
rect 92 5414 1904 5466
rect 1956 5414 1968 5466
rect 2020 5414 2032 5466
rect 2084 5414 2096 5466
rect 2148 5414 2160 5466
rect 2212 5414 5837 5466
rect 5889 5414 5901 5466
rect 5953 5414 5965 5466
rect 6017 5414 6029 5466
rect 6081 5414 6093 5466
rect 6145 5414 9770 5466
rect 9822 5414 9834 5466
rect 9886 5414 9898 5466
rect 9950 5414 9962 5466
rect 10014 5414 10026 5466
rect 10078 5414 13703 5466
rect 13755 5414 13767 5466
rect 13819 5414 13831 5466
rect 13883 5414 13895 5466
rect 13947 5414 13959 5466
rect 14011 5414 15824 5466
rect 92 5392 15824 5414
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 3789 5355 3847 5361
rect 3789 5352 3801 5355
rect 3752 5324 3801 5352
rect 3752 5312 3758 5324
rect 3789 5321 3801 5324
rect 3835 5321 3847 5355
rect 4062 5352 4068 5364
rect 3789 5315 3847 5321
rect 3896 5324 4068 5352
rect 3896 5284 3924 5324
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 5166 5312 5172 5364
rect 5224 5312 5230 5364
rect 5350 5312 5356 5364
rect 5408 5352 5414 5364
rect 7282 5352 7288 5364
rect 5408 5324 7288 5352
rect 5408 5312 5414 5324
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 10962 5352 10968 5364
rect 9232 5324 10968 5352
rect 3344 5256 3924 5284
rect 3344 5157 3372 5256
rect 4706 5244 4712 5296
rect 4764 5284 4770 5296
rect 5368 5284 5396 5312
rect 4764 5256 5396 5284
rect 7745 5287 7803 5293
rect 4764 5244 4770 5256
rect 7745 5253 7757 5287
rect 7791 5284 7803 5287
rect 8294 5284 8300 5296
rect 7791 5256 8300 5284
rect 7791 5253 7803 5256
rect 7745 5247 7803 5253
rect 3970 5216 3976 5228
rect 3436 5188 3976 5216
rect 3436 5157 3464 5188
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 4801 5219 4859 5225
rect 4801 5216 4813 5219
rect 4212 5188 4813 5216
rect 4212 5176 4218 5188
rect 4801 5185 4813 5188
rect 4847 5185 4859 5219
rect 7760 5216 7788 5247
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 8754 5244 8760 5296
rect 8812 5284 8818 5296
rect 8812 5256 9168 5284
rect 8812 5244 8818 5256
rect 4801 5179 4859 5185
rect 7484 5188 7788 5216
rect 8220 5188 8984 5216
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 3421 5151 3479 5157
rect 3421 5117 3433 5151
rect 3467 5117 3479 5151
rect 3421 5111 3479 5117
rect 3436 5080 3464 5111
rect 3510 5108 3516 5160
rect 3568 5108 3574 5160
rect 3605 5151 3663 5157
rect 3605 5117 3617 5151
rect 3651 5148 3663 5151
rect 3786 5148 3792 5160
rect 3651 5120 3792 5148
rect 3651 5117 3663 5120
rect 3605 5111 3663 5117
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 3878 5108 3884 5160
rect 3936 5108 3942 5160
rect 4522 5108 4528 5160
rect 4580 5108 4586 5160
rect 4706 5108 4712 5160
rect 4764 5148 4770 5160
rect 4985 5151 5043 5157
rect 4985 5148 4997 5151
rect 4764 5120 4997 5148
rect 4764 5108 4770 5120
rect 4985 5117 4997 5120
rect 5031 5117 5043 5151
rect 4985 5111 5043 5117
rect 5166 5108 5172 5160
rect 5224 5148 5230 5160
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 5224 5120 5273 5148
rect 5224 5108 5230 5120
rect 5261 5117 5273 5120
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 5626 5108 5632 5160
rect 5684 5108 5690 5160
rect 5718 5108 5724 5160
rect 5776 5108 5782 5160
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 6089 5151 6147 5157
rect 6089 5148 6101 5151
rect 5960 5120 6101 5148
rect 5960 5108 5966 5120
rect 6089 5117 6101 5120
rect 6135 5148 6147 5151
rect 6178 5148 6184 5160
rect 6135 5120 6184 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 6178 5108 6184 5120
rect 6236 5108 6242 5160
rect 6457 5151 6515 5157
rect 6457 5117 6469 5151
rect 6503 5117 6515 5151
rect 6457 5111 6515 5117
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 7006 5148 7012 5160
rect 6871 5120 7012 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 2976 5052 3464 5080
rect 3896 5080 3924 5108
rect 3973 5083 4031 5089
rect 3973 5080 3985 5083
rect 3896 5052 3985 5080
rect 2976 5024 3004 5052
rect 3973 5049 3985 5052
rect 4019 5049 4031 5083
rect 3973 5043 4031 5049
rect 4065 5083 4123 5089
rect 4065 5049 4077 5083
rect 4111 5080 4123 5083
rect 4246 5080 4252 5092
rect 4111 5052 4252 5080
rect 4111 5049 4123 5052
rect 4065 5043 4123 5049
rect 4246 5040 4252 5052
rect 4304 5080 4310 5092
rect 5445 5083 5503 5089
rect 5445 5080 5457 5083
rect 4304 5052 5457 5080
rect 4304 5040 4310 5052
rect 5445 5049 5457 5052
rect 5491 5049 5503 5083
rect 5445 5043 5503 5049
rect 5534 5040 5540 5092
rect 5592 5080 5598 5092
rect 5813 5083 5871 5089
rect 5813 5080 5825 5083
rect 5592 5052 5825 5080
rect 5592 5040 5598 5052
rect 5813 5049 5825 5052
rect 5859 5049 5871 5083
rect 6270 5080 6276 5092
rect 5813 5043 5871 5049
rect 5920 5052 6276 5080
rect 2958 4972 2964 5024
rect 3016 4972 3022 5024
rect 3694 4972 3700 5024
rect 3752 5012 3758 5024
rect 4157 5015 4215 5021
rect 4157 5012 4169 5015
rect 3752 4984 4169 5012
rect 3752 4972 3758 4984
rect 4157 4981 4169 4984
rect 4203 5012 4215 5015
rect 5626 5012 5632 5024
rect 4203 4984 5632 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 5626 4972 5632 4984
rect 5684 5012 5690 5024
rect 5920 5012 5948 5052
rect 6270 5040 6276 5052
rect 6328 5080 6334 5092
rect 6472 5080 6500 5111
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5148 7159 5151
rect 7190 5148 7196 5160
rect 7147 5120 7196 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 7282 5108 7288 5160
rect 7340 5157 7346 5160
rect 7484 5157 7512 5188
rect 7340 5151 7367 5157
rect 7355 5117 7367 5151
rect 7340 5111 7367 5117
rect 7469 5151 7527 5157
rect 7469 5117 7481 5151
rect 7515 5117 7527 5151
rect 7469 5111 7527 5117
rect 7561 5151 7619 5157
rect 7561 5117 7573 5151
rect 7607 5117 7619 5151
rect 7561 5111 7619 5117
rect 7340 5108 7346 5111
rect 7576 5080 7604 5111
rect 7650 5108 7656 5160
rect 7708 5148 7714 5160
rect 8220 5157 8248 5188
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 7708 5120 8217 5148
rect 7708 5108 7714 5120
rect 8205 5117 8217 5120
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 8294 5108 8300 5160
rect 8352 5108 8358 5160
rect 8390 5151 8448 5157
rect 8390 5117 8402 5151
rect 8436 5117 8448 5151
rect 8390 5111 8448 5117
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 8405 5080 8433 5111
rect 6328 5052 6500 5080
rect 7024 5052 7604 5080
rect 8312 5052 8433 5080
rect 8588 5080 8616 5111
rect 8662 5108 8668 5160
rect 8720 5108 8726 5160
rect 8754 5108 8760 5160
rect 8812 5157 8818 5160
rect 8812 5148 8820 5157
rect 8956 5150 8984 5188
rect 9033 5151 9091 5157
rect 9033 5150 9045 5151
rect 8812 5120 8857 5148
rect 8956 5122 9045 5150
rect 8812 5111 8820 5120
rect 9033 5117 9045 5122
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 8812 5108 8818 5111
rect 9140 5080 9168 5256
rect 9232 5157 9260 5324
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 12584 5324 14412 5352
rect 12584 5312 12590 5324
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 9861 5287 9919 5293
rect 9861 5284 9873 5287
rect 9732 5256 9873 5284
rect 9732 5244 9738 5256
rect 9861 5253 9873 5256
rect 9907 5284 9919 5287
rect 10229 5287 10287 5293
rect 9907 5256 10180 5284
rect 9907 5253 9919 5256
rect 9861 5247 9919 5253
rect 9646 5188 9904 5216
rect 9646 5160 9674 5188
rect 9217 5151 9275 5157
rect 9217 5117 9229 5151
rect 9263 5117 9275 5151
rect 9217 5111 9275 5117
rect 9582 5108 9588 5160
rect 9640 5120 9674 5160
rect 9769 5151 9827 5157
rect 9640 5108 9646 5120
rect 9769 5117 9781 5151
rect 9815 5117 9827 5151
rect 9876 5148 9904 5188
rect 9950 5176 9956 5228
rect 10008 5216 10014 5228
rect 10045 5219 10103 5225
rect 10045 5216 10057 5219
rect 10008 5188 10057 5216
rect 10008 5176 10014 5188
rect 10045 5185 10057 5188
rect 10091 5185 10103 5219
rect 10152 5216 10180 5256
rect 10229 5253 10241 5287
rect 10275 5284 10287 5287
rect 13078 5284 13084 5296
rect 10275 5256 13084 5284
rect 10275 5253 10287 5256
rect 10229 5247 10287 5253
rect 13078 5244 13084 5256
rect 13136 5244 13142 5296
rect 10778 5216 10784 5228
rect 10152 5188 10784 5216
rect 10045 5179 10103 5185
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 13906 5216 13912 5228
rect 11164 5188 13912 5216
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 9876 5120 10333 5148
rect 9769 5111 9827 5117
rect 10321 5117 10333 5120
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 9784 5080 9812 5111
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 11164 5157 11192 5188
rect 13906 5176 13912 5188
rect 13964 5176 13970 5228
rect 11149 5151 11207 5157
rect 11149 5148 11161 5151
rect 11112 5120 11161 5148
rect 11112 5108 11118 5120
rect 11149 5117 11161 5120
rect 11195 5117 11207 5151
rect 11149 5111 11207 5117
rect 12710 5108 12716 5160
rect 12768 5108 12774 5160
rect 13078 5108 13084 5160
rect 13136 5108 13142 5160
rect 14384 5148 14412 5324
rect 14384 5120 14490 5148
rect 13357 5083 13415 5089
rect 13357 5080 13369 5083
rect 8588 5052 9076 5080
rect 9140 5052 9812 5080
rect 12912 5052 13369 5080
rect 6328 5040 6334 5052
rect 7024 5024 7052 5052
rect 8312 5024 8340 5052
rect 5684 4984 5948 5012
rect 5684 4972 5690 4984
rect 5994 4972 6000 5024
rect 6052 4972 6058 5024
rect 7006 4972 7012 5024
rect 7064 4972 7070 5024
rect 7374 4972 7380 5024
rect 7432 4972 7438 5024
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 8113 5015 8171 5021
rect 8113 5012 8125 5015
rect 7892 4984 8125 5012
rect 7892 4972 7898 4984
rect 8113 4981 8125 4984
rect 8159 4981 8171 5015
rect 8113 4975 8171 4981
rect 8294 4972 8300 5024
rect 8352 4972 8358 5024
rect 8938 4972 8944 5024
rect 8996 4972 9002 5024
rect 9048 5021 9076 5052
rect 9033 5015 9091 5021
rect 9033 4981 9045 5015
rect 9079 4981 9091 5015
rect 9033 4975 9091 4981
rect 10045 5015 10103 5021
rect 10045 4981 10057 5015
rect 10091 5012 10103 5015
rect 10134 5012 10140 5024
rect 10091 4984 10140 5012
rect 10091 4981 10103 4984
rect 10045 4975 10103 4981
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 10962 4972 10968 5024
rect 11020 4972 11026 5024
rect 12912 5021 12940 5052
rect 13357 5049 13369 5052
rect 13403 5049 13415 5083
rect 14921 5083 14979 5089
rect 14921 5080 14933 5083
rect 13357 5043 13415 5049
rect 14660 5052 14933 5080
rect 12897 5015 12955 5021
rect 12897 4981 12909 5015
rect 12943 4981 12955 5015
rect 12897 4975 12955 4981
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14660 5012 14688 5052
rect 14921 5049 14933 5052
rect 14967 5049 14979 5083
rect 14921 5043 14979 5049
rect 15105 5083 15163 5089
rect 15105 5049 15117 5083
rect 15151 5049 15163 5083
rect 15105 5043 15163 5049
rect 14056 4984 14688 5012
rect 14056 4972 14062 4984
rect 14734 4972 14740 5024
rect 14792 5012 14798 5024
rect 14829 5015 14887 5021
rect 14829 5012 14841 5015
rect 14792 4984 14841 5012
rect 14792 4972 14798 4984
rect 14829 4981 14841 4984
rect 14875 5012 14887 5015
rect 15120 5012 15148 5043
rect 14875 4984 15148 5012
rect 14875 4981 14887 4984
rect 14829 4975 14887 4981
rect 15194 4972 15200 5024
rect 15252 5012 15258 5024
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 15252 4984 15301 5012
rect 15252 4972 15258 4984
rect 15289 4981 15301 4984
rect 15335 4981 15347 5015
rect 15289 4975 15347 4981
rect 92 4922 15824 4944
rect 92 4870 2564 4922
rect 2616 4870 2628 4922
rect 2680 4870 2692 4922
rect 2744 4870 2756 4922
rect 2808 4870 2820 4922
rect 2872 4870 6497 4922
rect 6549 4870 6561 4922
rect 6613 4870 6625 4922
rect 6677 4870 6689 4922
rect 6741 4870 6753 4922
rect 6805 4870 10430 4922
rect 10482 4870 10494 4922
rect 10546 4870 10558 4922
rect 10610 4870 10622 4922
rect 10674 4870 10686 4922
rect 10738 4870 14363 4922
rect 14415 4870 14427 4922
rect 14479 4870 14491 4922
rect 14543 4870 14555 4922
rect 14607 4870 14619 4922
rect 14671 4870 15824 4922
rect 92 4848 15824 4870
rect 6181 4811 6239 4817
rect 6181 4808 6193 4811
rect 3068 4780 6193 4808
rect 382 4632 388 4684
rect 440 4632 446 4684
rect 1762 4632 1768 4684
rect 1820 4672 1826 4684
rect 2314 4672 2320 4684
rect 1820 4644 2320 4672
rect 1820 4632 1826 4644
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 2777 4675 2835 4681
rect 2777 4641 2789 4675
rect 2823 4672 2835 4675
rect 2958 4672 2964 4684
rect 2823 4644 2964 4672
rect 2823 4641 2835 4644
rect 2777 4635 2835 4641
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 3068 4681 3096 4780
rect 6181 4777 6193 4780
rect 6227 4777 6239 4811
rect 6181 4771 6239 4777
rect 7006 4768 7012 4820
rect 7064 4768 7070 4820
rect 7374 4768 7380 4820
rect 7432 4768 7438 4820
rect 7466 4768 7472 4820
rect 7524 4768 7530 4820
rect 7653 4811 7711 4817
rect 7653 4777 7665 4811
rect 7699 4808 7711 4811
rect 8846 4808 8852 4820
rect 7699 4780 8852 4808
rect 7699 4777 7711 4780
rect 7653 4771 7711 4777
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 11054 4768 11060 4820
rect 11112 4768 11118 4820
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 12989 4811 13047 4817
rect 12989 4808 13001 4811
rect 12768 4780 13001 4808
rect 12768 4768 12774 4780
rect 12989 4777 13001 4780
rect 13035 4777 13047 4811
rect 13998 4808 14004 4820
rect 12989 4771 13047 4777
rect 13096 4780 14004 4808
rect 4798 4700 4804 4752
rect 4856 4700 4862 4752
rect 5169 4743 5227 4749
rect 5169 4709 5181 4743
rect 5215 4740 5227 4743
rect 5350 4740 5356 4752
rect 5215 4712 5356 4740
rect 5215 4709 5227 4712
rect 5169 4703 5227 4709
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 7024 4740 7052 4768
rect 6288 4712 7052 4740
rect 3053 4675 3111 4681
rect 3053 4641 3065 4675
rect 3099 4641 3111 4675
rect 3053 4635 3111 4641
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 3510 4672 3516 4684
rect 3283 4644 3516 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 3510 4632 3516 4644
rect 3568 4632 3574 4684
rect 3694 4632 3700 4684
rect 3752 4632 3758 4684
rect 4816 4672 4844 4700
rect 3988 4644 4844 4672
rect 658 4564 664 4616
rect 716 4564 722 4616
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 3988 4613 4016 4644
rect 5442 4632 5448 4684
rect 5500 4632 5506 4684
rect 5626 4632 5632 4684
rect 5684 4632 5690 4684
rect 5810 4632 5816 4684
rect 5868 4632 5874 4684
rect 5994 4632 6000 4684
rect 6052 4672 6058 4684
rect 6089 4675 6147 4681
rect 6089 4672 6101 4675
rect 6052 4644 6101 4672
rect 6052 4632 6058 4644
rect 6089 4641 6101 4644
rect 6135 4672 6147 4675
rect 6178 4672 6184 4684
rect 6135 4644 6184 4672
rect 6135 4641 6147 4644
rect 6089 4635 6147 4641
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6288 4681 6316 4712
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4641 6331 4675
rect 6273 4635 6331 4641
rect 6641 4675 6699 4681
rect 6641 4641 6653 4675
rect 6687 4672 6699 4675
rect 6822 4672 6828 4684
rect 6687 4644 6828 4672
rect 6687 4641 6699 4644
rect 6641 4635 6699 4641
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4641 6975 4675
rect 6917 4635 6975 4641
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 4764 4576 4813 4604
rect 4764 4564 4770 4576
rect 4801 4573 4813 4576
rect 4847 4604 4859 4607
rect 5258 4604 5264 4616
rect 4847 4576 5264 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 5258 4564 5264 4576
rect 5316 4604 5322 4616
rect 5353 4607 5411 4613
rect 5353 4604 5365 4607
rect 5316 4576 5365 4604
rect 5316 4564 5322 4576
rect 5353 4573 5365 4576
rect 5399 4573 5411 4607
rect 6932 4604 6960 4635
rect 7006 4632 7012 4684
rect 7064 4632 7070 4684
rect 7392 4672 7420 4768
rect 8938 4700 8944 4752
rect 8996 4740 9002 4752
rect 9033 4743 9091 4749
rect 9033 4740 9045 4743
rect 8996 4712 9045 4740
rect 8996 4700 9002 4712
rect 9033 4709 9045 4712
rect 9079 4740 9091 4743
rect 9079 4712 9536 4740
rect 9079 4709 9091 4712
rect 9033 4703 9091 4709
rect 8297 4675 8355 4681
rect 8297 4672 8309 4675
rect 7392 4644 8309 4672
rect 8297 4641 8309 4644
rect 8343 4641 8355 4675
rect 8297 4635 8355 4641
rect 8478 4632 8484 4684
rect 8536 4632 8542 4684
rect 9508 4681 9536 4712
rect 10226 4700 10232 4752
rect 10284 4740 10290 4752
rect 11072 4740 11100 4768
rect 13096 4740 13124 4780
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14826 4768 14832 4820
rect 14884 4768 14890 4820
rect 14734 4740 14740 4752
rect 10284 4712 11100 4740
rect 12820 4712 13124 4740
rect 13832 4712 14740 4740
rect 10284 4700 10290 4712
rect 9217 4675 9275 4681
rect 9217 4641 9229 4675
rect 9263 4641 9275 4675
rect 9217 4635 9275 4641
rect 9493 4675 9551 4681
rect 9493 4641 9505 4675
rect 9539 4641 9551 4675
rect 9493 4635 9551 4641
rect 7098 4604 7104 4616
rect 6932 4576 7104 4604
rect 5353 4567 5411 4573
rect 7098 4564 7104 4576
rect 7156 4564 7162 4616
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 9232 4604 9260 4635
rect 9582 4632 9588 4684
rect 9640 4672 9646 4684
rect 9953 4675 10011 4681
rect 9953 4672 9965 4675
rect 9640 4644 9965 4672
rect 9640 4632 9646 4644
rect 9953 4641 9965 4644
rect 9999 4641 10011 4675
rect 9953 4635 10011 4641
rect 12434 4632 12440 4684
rect 12492 4632 12498 4684
rect 7616 4576 9260 4604
rect 11057 4607 11115 4613
rect 7616 4564 7622 4576
rect 11057 4573 11069 4607
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4604 11391 4607
rect 11422 4604 11428 4616
rect 11379 4576 11428 4604
rect 11379 4573 11391 4576
rect 11333 4567 11391 4573
rect 2406 4496 2412 4548
rect 2464 4536 2470 4548
rect 3053 4539 3111 4545
rect 3053 4536 3065 4539
rect 2464 4508 3065 4536
rect 2464 4496 2470 4508
rect 3053 4505 3065 4508
rect 3099 4505 3111 4539
rect 3804 4536 3832 4564
rect 5031 4539 5089 4545
rect 5031 4536 5043 4539
rect 3804 4508 5043 4536
rect 3053 4499 3111 4505
rect 5031 4505 5043 4508
rect 5077 4505 5089 4539
rect 5031 4499 5089 4505
rect 1118 4428 1124 4480
rect 1176 4468 1182 4480
rect 2133 4471 2191 4477
rect 2133 4468 2145 4471
rect 1176 4440 2145 4468
rect 1176 4428 1182 4440
rect 2133 4437 2145 4440
rect 2179 4437 2191 4471
rect 2133 4431 2191 4437
rect 3326 4428 3332 4480
rect 3384 4428 3390 4480
rect 4522 4428 4528 4480
rect 4580 4428 4586 4480
rect 4614 4428 4620 4480
rect 4672 4468 4678 4480
rect 4893 4471 4951 4477
rect 4893 4468 4905 4471
rect 4672 4440 4905 4468
rect 4672 4428 4678 4440
rect 4893 4437 4905 4440
rect 4939 4437 4951 4471
rect 5046 4468 5074 4499
rect 5166 4496 5172 4548
rect 5224 4536 5230 4548
rect 7193 4539 7251 4545
rect 7193 4536 7205 4539
rect 5224 4508 7205 4536
rect 5224 4496 5230 4508
rect 7193 4505 7205 4508
rect 7239 4536 7251 4539
rect 8021 4539 8079 4545
rect 7239 4508 7788 4536
rect 7239 4505 7251 4508
rect 7193 4499 7251 4505
rect 5718 4468 5724 4480
rect 5046 4440 5724 4468
rect 4893 4431 4951 4437
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 6457 4471 6515 4477
rect 6457 4437 6469 4471
rect 6503 4468 6515 4471
rect 6546 4468 6552 4480
rect 6503 4440 6552 4468
rect 6503 4437 6515 4440
rect 6457 4431 6515 4437
rect 6546 4428 6552 4440
rect 6604 4428 6610 4480
rect 6638 4428 6644 4480
rect 6696 4468 6702 4480
rect 6825 4471 6883 4477
rect 6825 4468 6837 4471
rect 6696 4440 6837 4468
rect 6696 4428 6702 4440
rect 6825 4437 6837 4440
rect 6871 4468 6883 4471
rect 7558 4468 7564 4480
rect 6871 4440 7564 4468
rect 6871 4437 6883 4440
rect 6825 4431 6883 4437
rect 7558 4428 7564 4440
rect 7616 4428 7622 4480
rect 7661 4471 7719 4477
rect 7661 4437 7673 4471
rect 7707 4468 7719 4471
rect 7760 4468 7788 4508
rect 8021 4505 8033 4539
rect 8067 4536 8079 4539
rect 8110 4536 8116 4548
rect 8067 4508 8116 4536
rect 8067 4505 8079 4508
rect 8021 4499 8079 4505
rect 8110 4496 8116 4508
rect 8168 4496 8174 4548
rect 8478 4496 8484 4548
rect 8536 4536 8542 4548
rect 9950 4536 9956 4548
rect 8536 4508 9956 4536
rect 8536 4496 8542 4508
rect 9950 4496 9956 4508
rect 10008 4496 10014 4548
rect 8294 4468 8300 4480
rect 7707 4440 8300 4468
rect 7707 4437 7719 4440
rect 7661 4431 7719 4437
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 8386 4428 8392 4480
rect 8444 4428 8450 4480
rect 9401 4471 9459 4477
rect 9401 4437 9413 4471
rect 9447 4468 9459 4471
rect 9674 4468 9680 4480
rect 9447 4440 9680 4468
rect 9447 4437 9459 4440
rect 9401 4431 9459 4437
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 11072 4468 11100 4567
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 12820 4480 12848 4712
rect 13173 4675 13231 4681
rect 13173 4641 13185 4675
rect 13219 4672 13231 4675
rect 13262 4672 13268 4684
rect 13219 4644 13268 4672
rect 13219 4641 13231 4644
rect 13173 4635 13231 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 13832 4681 13860 4712
rect 14734 4700 14740 4712
rect 14792 4700 14798 4752
rect 13817 4675 13875 4681
rect 13817 4641 13829 4675
rect 13863 4641 13875 4675
rect 13817 4635 13875 4641
rect 13906 4632 13912 4684
rect 13964 4672 13970 4684
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 13964 4644 14105 4672
rect 13964 4632 13970 4644
rect 14093 4641 14105 4644
rect 14139 4672 14151 4675
rect 14458 4672 14464 4684
rect 14139 4644 14464 4672
rect 14139 4641 14151 4644
rect 14093 4635 14151 4641
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 14642 4632 14648 4684
rect 14700 4632 14706 4684
rect 15378 4632 15384 4684
rect 15436 4632 15442 4684
rect 13357 4607 13415 4613
rect 13357 4573 13369 4607
rect 13403 4604 13415 4607
rect 13633 4607 13691 4613
rect 13633 4604 13645 4607
rect 13403 4576 13645 4604
rect 13403 4573 13415 4576
rect 13357 4567 13415 4573
rect 13633 4573 13645 4576
rect 13679 4573 13691 4607
rect 13633 4567 13691 4573
rect 11330 4468 11336 4480
rect 11072 4440 11336 4468
rect 11330 4428 11336 4440
rect 11388 4428 11394 4480
rect 12802 4428 12808 4480
rect 12860 4428 12866 4480
rect 15286 4428 15292 4480
rect 15344 4428 15350 4480
rect 92 4378 15824 4400
rect 92 4326 1904 4378
rect 1956 4326 1968 4378
rect 2020 4326 2032 4378
rect 2084 4326 2096 4378
rect 2148 4326 2160 4378
rect 2212 4326 5837 4378
rect 5889 4326 5901 4378
rect 5953 4326 5965 4378
rect 6017 4326 6029 4378
rect 6081 4326 6093 4378
rect 6145 4326 9770 4378
rect 9822 4326 9834 4378
rect 9886 4326 9898 4378
rect 9950 4326 9962 4378
rect 10014 4326 10026 4378
rect 10078 4326 13703 4378
rect 13755 4326 13767 4378
rect 13819 4326 13831 4378
rect 13883 4326 13895 4378
rect 13947 4326 13959 4378
rect 14011 4326 15824 4378
rect 92 4304 15824 4326
rect 658 4224 664 4276
rect 716 4264 722 4276
rect 1397 4267 1455 4273
rect 1397 4264 1409 4267
rect 716 4236 1409 4264
rect 716 4224 722 4236
rect 1397 4233 1409 4236
rect 1443 4233 1455 4267
rect 6825 4267 6883 4273
rect 1397 4227 1455 4233
rect 2746 4236 6776 4264
rect 2746 4196 2774 4236
rect 5166 4196 5172 4208
rect 1136 4168 2774 4196
rect 4724 4168 5172 4196
rect 1136 4072 1164 4168
rect 4522 4128 4528 4140
rect 1228 4100 4528 4128
rect 845 4063 903 4069
rect 845 4029 857 4063
rect 891 4060 903 4063
rect 891 4032 980 4060
rect 891 4029 903 4032
rect 845 4023 903 4029
rect 952 3936 980 4032
rect 1026 4020 1032 4072
rect 1084 4020 1090 4072
rect 1118 4020 1124 4072
rect 1176 4020 1182 4072
rect 1228 4069 1256 4100
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 1213 4063 1271 4069
rect 1213 4029 1225 4063
rect 1259 4029 1271 4063
rect 1213 4023 1271 4029
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4060 2467 4063
rect 3326 4060 3332 4072
rect 2455 4032 3332 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 3694 4020 3700 4072
rect 3752 4020 3758 4072
rect 4724 4069 4752 4168
rect 5166 4156 5172 4168
rect 5224 4156 5230 4208
rect 6546 4196 6552 4208
rect 5552 4168 6552 4196
rect 5552 4128 5580 4168
rect 6546 4156 6552 4168
rect 6604 4156 6610 4208
rect 6748 4196 6776 4236
rect 6825 4233 6837 4267
rect 6871 4264 6883 4267
rect 7466 4264 7472 4276
rect 6871 4236 7472 4264
rect 6871 4233 6883 4236
rect 6825 4227 6883 4233
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 8846 4224 8852 4276
rect 8904 4264 8910 4276
rect 8904 4236 11284 4264
rect 8904 4224 8910 4236
rect 7098 4196 7104 4208
rect 6748 4168 7104 4196
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 8018 4156 8024 4208
rect 8076 4196 8082 4208
rect 8205 4199 8263 4205
rect 8205 4196 8217 4199
rect 8076 4168 8217 4196
rect 8076 4156 8082 4168
rect 8205 4165 8217 4168
rect 8251 4196 8263 4199
rect 8478 4196 8484 4208
rect 8251 4168 8484 4196
rect 8251 4165 8263 4168
rect 8205 4159 8263 4165
rect 8478 4156 8484 4168
rect 8536 4156 8542 4208
rect 10134 4156 10140 4208
rect 10192 4156 10198 4208
rect 10502 4156 10508 4208
rect 10560 4156 10566 4208
rect 11256 4196 11284 4236
rect 11422 4224 11428 4276
rect 11480 4264 11486 4276
rect 11517 4267 11575 4273
rect 11517 4264 11529 4267
rect 11480 4236 11529 4264
rect 11480 4224 11486 4236
rect 11517 4233 11529 4236
rect 11563 4233 11575 4267
rect 11517 4227 11575 4233
rect 12802 4196 12808 4208
rect 11256 4168 12808 4196
rect 5000 4100 5580 4128
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4617 4063 4675 4069
rect 4617 4029 4629 4063
rect 4663 4029 4675 4063
rect 4617 4023 4675 4029
rect 4709 4063 4767 4069
rect 4709 4029 4721 4063
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 4264 3936 4292 4023
rect 934 3884 940 3936
rect 992 3884 998 3936
rect 2222 3884 2228 3936
rect 2280 3884 2286 3936
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 3142 3924 3148 3936
rect 2372 3896 3148 3924
rect 2372 3884 2378 3896
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 4246 3884 4252 3936
rect 4304 3884 4310 3936
rect 4430 3884 4436 3936
rect 4488 3884 4494 3936
rect 4632 3924 4660 4023
rect 4798 4020 4804 4072
rect 4856 4020 4862 4072
rect 5000 4069 5028 4100
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5776 4100 5917 4128
rect 5776 4088 5782 4100
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 5905 4091 5963 4097
rect 6104 4100 6469 4128
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4029 5043 4063
rect 5445 4063 5503 4069
rect 5445 4060 5457 4063
rect 4985 4023 5043 4029
rect 5092 4032 5457 4060
rect 4798 3924 4804 3936
rect 4632 3896 4804 3924
rect 4798 3884 4804 3896
rect 4856 3924 4862 3936
rect 5092 3924 5120 4032
rect 5445 4029 5457 4032
rect 5491 4060 5503 4063
rect 5534 4060 5540 4072
rect 5491 4032 5540 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 6104 4069 6132 4100
rect 6457 4097 6469 4100
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6880 4100 6929 4128
rect 6880 4088 6886 4100
rect 6917 4097 6929 4100
rect 6963 4128 6975 4131
rect 8386 4128 8392 4140
rect 6963 4100 7052 4128
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4029 5687 4063
rect 5629 4023 5687 4029
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4029 6147 4063
rect 6089 4023 6147 4029
rect 5166 3952 5172 4004
rect 5224 3952 5230 4004
rect 5644 3992 5672 4023
rect 6178 4020 6184 4072
rect 6236 4020 6242 4072
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 6638 4060 6644 4072
rect 6328 4032 6644 4060
rect 6328 4020 6334 4032
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 6730 4020 6736 4072
rect 6788 4020 6794 4072
rect 7024 4069 7052 4100
rect 7208 4100 8392 4128
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4029 7067 4063
rect 7009 4023 7067 4029
rect 5460 3964 5672 3992
rect 5460 3936 5488 3964
rect 4856 3896 5120 3924
rect 4856 3884 4862 3896
rect 5258 3884 5264 3936
rect 5316 3884 5322 3936
rect 5442 3884 5448 3936
rect 5500 3884 5506 3936
rect 5534 3884 5540 3936
rect 5592 3884 5598 3936
rect 6748 3924 6776 4020
rect 6822 3952 6828 4004
rect 6880 3992 6886 4004
rect 7208 3992 7236 4100
rect 8386 4088 8392 4100
rect 8444 4128 8450 4140
rect 9306 4128 9312 4140
rect 8444 4100 9312 4128
rect 8444 4088 8450 4100
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 10152 4128 10180 4156
rect 9600 4100 10180 4128
rect 7282 4020 7288 4072
rect 7340 4060 7346 4072
rect 8662 4060 8668 4072
rect 7340 4032 8668 4060
rect 7340 4020 7346 4032
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9600 4069 9628 4100
rect 9401 4063 9459 4069
rect 9401 4029 9413 4063
rect 9447 4029 9459 4063
rect 9401 4023 9459 4029
rect 9585 4063 9643 4069
rect 9585 4029 9597 4063
rect 9631 4029 9643 4063
rect 9585 4023 9643 4029
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4060 9735 4063
rect 10318 4060 10324 4072
rect 9723 4032 10324 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 6880 3964 7236 3992
rect 7469 3995 7527 4001
rect 6880 3952 6886 3964
rect 7469 3961 7481 3995
rect 7515 3992 7527 3995
rect 8021 3995 8079 4001
rect 8021 3992 8033 3995
rect 7515 3964 8033 3992
rect 7515 3961 7527 3964
rect 7469 3955 7527 3961
rect 8021 3961 8033 3964
rect 8067 3961 8079 3995
rect 8021 3955 8079 3961
rect 8938 3952 8944 4004
rect 8996 3952 9002 4004
rect 9416 3992 9444 4023
rect 10318 4020 10324 4032
rect 10376 4020 10382 4072
rect 10870 4060 10876 4072
rect 10428 4032 10876 4060
rect 9416 3964 9674 3992
rect 7101 3927 7159 3933
rect 7101 3924 7113 3927
rect 6748 3896 7113 3924
rect 7101 3893 7113 3896
rect 7147 3924 7159 3927
rect 7374 3924 7380 3936
rect 7147 3896 7380 3924
rect 7147 3893 7159 3896
rect 7101 3887 7159 3893
rect 7374 3884 7380 3896
rect 7432 3924 7438 3936
rect 7834 3924 7840 3936
rect 7432 3896 7840 3924
rect 7432 3884 7438 3896
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 9646 3924 9674 3964
rect 10134 3952 10140 4004
rect 10192 3992 10198 4004
rect 10428 3992 10456 4032
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11054 4060 11060 4072
rect 11011 4032 11060 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 11256 4069 11284 4168
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13280 4100 13829 4128
rect 13280 4072 13308 4100
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 15562 4088 15568 4140
rect 15620 4088 15626 4140
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4029 11299 4063
rect 11241 4023 11299 4029
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4029 11391 4063
rect 11333 4023 11391 4029
rect 10192 3964 10456 3992
rect 10192 3952 10198 3964
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 11149 3995 11207 4001
rect 11149 3992 11161 3995
rect 10836 3964 11161 3992
rect 10836 3952 10842 3964
rect 11149 3961 11161 3964
rect 11195 3961 11207 3995
rect 11149 3955 11207 3961
rect 10226 3924 10232 3936
rect 9646 3896 10232 3924
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 11348 3924 11376 4023
rect 13262 4020 13268 4072
rect 13320 4020 13326 4072
rect 13538 4020 13544 4072
rect 13596 4060 13602 4072
rect 13633 4063 13691 4069
rect 13633 4060 13645 4063
rect 13596 4032 13645 4060
rect 13596 4020 13602 4032
rect 13633 4029 13645 4032
rect 13679 4029 13691 4063
rect 13633 4023 13691 4029
rect 14458 4020 14464 4072
rect 14516 4060 14522 4072
rect 15105 4063 15163 4069
rect 14516 4032 14780 4060
rect 14516 4020 14522 4032
rect 14752 4004 14780 4032
rect 15105 4029 15117 4063
rect 15151 4060 15163 4063
rect 15194 4060 15200 4072
rect 15151 4032 15200 4060
rect 15151 4029 15163 4032
rect 15105 4023 15163 4029
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 15378 4020 15384 4072
rect 15436 4020 15442 4072
rect 14734 3952 14740 4004
rect 14792 3952 14798 4004
rect 15010 3992 15016 4004
rect 14936 3964 15016 3992
rect 10928 3896 11376 3924
rect 10928 3884 10934 3896
rect 13354 3884 13360 3936
rect 13412 3924 13418 3936
rect 13449 3927 13507 3933
rect 13449 3924 13461 3927
rect 13412 3896 13461 3924
rect 13412 3884 13418 3896
rect 13449 3893 13461 3896
rect 13495 3893 13507 3927
rect 13449 3887 13507 3893
rect 14274 3884 14280 3936
rect 14332 3884 14338 3936
rect 14936 3933 14964 3964
rect 15010 3952 15016 3964
rect 15068 3992 15074 4004
rect 15580 3992 15608 4088
rect 15068 3964 15608 3992
rect 15068 3952 15074 3964
rect 14921 3927 14979 3933
rect 14921 3893 14933 3927
rect 14967 3893 14979 3927
rect 14921 3887 14979 3893
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 15160 3896 15301 3924
rect 15160 3884 15166 3896
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 15289 3887 15347 3893
rect 92 3834 15824 3856
rect 92 3782 2564 3834
rect 2616 3782 2628 3834
rect 2680 3782 2692 3834
rect 2744 3782 2756 3834
rect 2808 3782 2820 3834
rect 2872 3782 6497 3834
rect 6549 3782 6561 3834
rect 6613 3782 6625 3834
rect 6677 3782 6689 3834
rect 6741 3782 6753 3834
rect 6805 3782 10430 3834
rect 10482 3782 10494 3834
rect 10546 3782 10558 3834
rect 10610 3782 10622 3834
rect 10674 3782 10686 3834
rect 10738 3782 14363 3834
rect 14415 3782 14427 3834
rect 14479 3782 14491 3834
rect 14543 3782 14555 3834
rect 14607 3782 14619 3834
rect 14671 3782 15824 3834
rect 92 3760 15824 3782
rect 474 3680 480 3732
rect 532 3680 538 3732
rect 934 3680 940 3732
rect 992 3680 998 3732
rect 5534 3720 5540 3732
rect 1780 3692 5540 3720
rect 753 3655 811 3661
rect 753 3621 765 3655
rect 799 3652 811 3655
rect 1780 3652 1808 3692
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 6914 3680 6920 3732
rect 6972 3720 6978 3732
rect 7558 3720 7564 3732
rect 6972 3692 7564 3720
rect 6972 3680 6978 3692
rect 7558 3680 7564 3692
rect 7616 3720 7622 3732
rect 7653 3723 7711 3729
rect 7653 3720 7665 3723
rect 7616 3692 7665 3720
rect 7616 3680 7622 3692
rect 7653 3689 7665 3692
rect 7699 3689 7711 3723
rect 10134 3720 10140 3732
rect 7653 3683 7711 3689
rect 8220 3692 10140 3720
rect 799 3624 1808 3652
rect 2133 3655 2191 3661
rect 799 3621 811 3624
rect 753 3615 811 3621
rect 2133 3621 2145 3655
rect 2179 3652 2191 3655
rect 2222 3652 2228 3664
rect 2179 3624 2228 3652
rect 2179 3621 2191 3624
rect 2133 3615 2191 3621
rect 2222 3612 2228 3624
rect 2280 3612 2286 3664
rect 3142 3612 3148 3664
rect 3200 3612 3206 3664
rect 4709 3655 4767 3661
rect 4709 3621 4721 3655
rect 4755 3652 4767 3655
rect 5258 3652 5264 3664
rect 4755 3624 5264 3652
rect 4755 3621 4767 3624
rect 4709 3615 4767 3621
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 6822 3612 6828 3664
rect 6880 3652 6886 3664
rect 7075 3655 7133 3661
rect 7075 3652 7087 3655
rect 6880 3624 7087 3652
rect 6880 3612 6886 3624
rect 7075 3621 7087 3624
rect 7121 3621 7133 3655
rect 7075 3615 7133 3621
rect 7466 3612 7472 3664
rect 7524 3652 7530 3664
rect 8113 3655 8171 3661
rect 8113 3652 8125 3655
rect 7524 3624 8125 3652
rect 7524 3612 7530 3624
rect 8113 3621 8125 3624
rect 8159 3621 8171 3655
rect 8113 3615 8171 3621
rect 1118 3544 1124 3596
rect 1176 3544 1182 3596
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 1857 3587 1915 3593
rect 1857 3584 1869 3587
rect 1728 3556 1869 3584
rect 1728 3544 1734 3556
rect 1857 3553 1869 3556
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 4571 3556 4752 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 4246 3516 4252 3528
rect 3651 3488 4252 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 4246 3476 4252 3488
rect 4304 3516 4310 3528
rect 4724 3516 4752 3556
rect 4798 3544 4804 3596
rect 4856 3544 4862 3596
rect 7190 3544 7196 3596
rect 7248 3544 7254 3596
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3553 7343 3587
rect 7285 3547 7343 3553
rect 7377 3587 7435 3593
rect 7377 3553 7389 3587
rect 7423 3584 7435 3587
rect 7558 3584 7564 3596
rect 7423 3556 7564 3584
rect 7423 3553 7435 3556
rect 7377 3547 7435 3553
rect 4304 3488 4752 3516
rect 4816 3516 4844 3544
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4816 3488 4905 3516
rect 4304 3476 4310 3488
rect 4724 3392 4752 3488
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 6822 3476 6828 3528
rect 6880 3516 6886 3528
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 6880 3488 6929 3516
rect 6880 3476 6886 3488
rect 6917 3485 6929 3488
rect 6963 3516 6975 3519
rect 6963 3488 7236 3516
rect 6963 3485 6975 3488
rect 6917 3479 6975 3485
rect 4706 3340 4712 3392
rect 4764 3340 4770 3392
rect 7208 3380 7236 3488
rect 7300 3448 7328 3547
rect 7558 3544 7564 3556
rect 7616 3544 7622 3596
rect 8220 3516 8248 3692
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10318 3680 10324 3732
rect 10376 3680 10382 3732
rect 11054 3680 11060 3732
rect 11112 3680 11118 3732
rect 11241 3723 11299 3729
rect 11241 3689 11253 3723
rect 11287 3689 11299 3723
rect 11241 3683 11299 3689
rect 10226 3652 10232 3664
rect 10074 3624 10232 3652
rect 10226 3612 10232 3624
rect 10284 3612 10290 3664
rect 10778 3612 10784 3664
rect 10836 3652 10842 3664
rect 10873 3655 10931 3661
rect 10873 3652 10885 3655
rect 10836 3624 10885 3652
rect 10836 3612 10842 3624
rect 10873 3621 10885 3624
rect 10919 3621 10931 3655
rect 10873 3615 10931 3621
rect 10965 3655 11023 3661
rect 10965 3621 10977 3655
rect 11011 3652 11023 3655
rect 11072 3652 11100 3680
rect 11256 3652 11284 3683
rect 12526 3680 12532 3732
rect 12584 3720 12590 3732
rect 12584 3692 13216 3720
rect 12584 3680 12590 3692
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 11011 3624 11192 3652
rect 11256 3624 11621 3652
rect 11011 3621 11023 3624
rect 10965 3615 11023 3621
rect 10686 3544 10692 3596
rect 10744 3544 10750 3596
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3553 11115 3587
rect 11164 3584 11192 3624
rect 11609 3621 11621 3624
rect 11655 3621 11667 3655
rect 11609 3615 11667 3621
rect 12728 3596 12756 3692
rect 13188 3652 13216 3692
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 15436 3692 15485 3720
rect 15436 3680 15442 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 15473 3683 15531 3689
rect 13188 3624 14214 3652
rect 11164 3556 11284 3584
rect 11057 3547 11115 3553
rect 7484 3488 8248 3516
rect 7374 3448 7380 3460
rect 7300 3420 7380 3448
rect 7374 3408 7380 3420
rect 7432 3408 7438 3460
rect 7484 3380 7512 3488
rect 8570 3476 8576 3528
rect 8628 3476 8634 3528
rect 8846 3476 8852 3528
rect 8904 3476 8910 3528
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 10318 3516 10324 3528
rect 9364 3488 10324 3516
rect 9364 3476 9370 3488
rect 10318 3476 10324 3488
rect 10376 3516 10382 3528
rect 10870 3516 10876 3528
rect 10376 3488 10876 3516
rect 10376 3476 10382 3488
rect 10870 3476 10876 3488
rect 10928 3516 10934 3528
rect 11072 3516 11100 3547
rect 10928 3488 11100 3516
rect 10928 3476 10934 3488
rect 7742 3408 7748 3460
rect 7800 3448 7806 3460
rect 8110 3448 8116 3460
rect 7800 3420 8116 3448
rect 7800 3408 7806 3420
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 7208 3352 7512 3380
rect 7558 3340 7564 3392
rect 7616 3340 7622 3392
rect 11256 3380 11284 3556
rect 12710 3544 12716 3596
rect 12768 3544 12774 3596
rect 13078 3544 13084 3596
rect 13136 3544 13142 3596
rect 13173 3587 13231 3593
rect 13173 3553 13185 3587
rect 13219 3584 13231 3587
rect 13354 3584 13360 3596
rect 13219 3556 13360 3584
rect 13219 3553 13231 3556
rect 13173 3547 13231 3553
rect 13354 3544 13360 3556
rect 13412 3544 13418 3596
rect 15286 3544 15292 3596
rect 15344 3544 15350 3596
rect 11330 3476 11336 3528
rect 11388 3516 11394 3528
rect 13096 3516 13124 3544
rect 13449 3519 13507 3525
rect 13449 3516 13461 3519
rect 11388 3488 13461 3516
rect 11388 3476 11394 3488
rect 13449 3485 13461 3488
rect 13495 3485 13507 3519
rect 13725 3519 13783 3525
rect 13725 3516 13737 3519
rect 13449 3479 13507 3485
rect 13556 3488 13737 3516
rect 13357 3451 13415 3457
rect 13357 3417 13369 3451
rect 13403 3448 13415 3451
rect 13556 3448 13584 3488
rect 13725 3485 13737 3488
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 13403 3420 13584 3448
rect 13403 3417 13415 3420
rect 13357 3411 13415 3417
rect 13081 3383 13139 3389
rect 13081 3380 13093 3383
rect 11256 3352 13093 3380
rect 13081 3349 13093 3352
rect 13127 3380 13139 3383
rect 13446 3380 13452 3392
rect 13127 3352 13452 3380
rect 13127 3349 13139 3352
rect 13081 3343 13139 3349
rect 13446 3340 13452 3352
rect 13504 3340 13510 3392
rect 14826 3340 14832 3392
rect 14884 3380 14890 3392
rect 15197 3383 15255 3389
rect 15197 3380 15209 3383
rect 14884 3352 15209 3380
rect 14884 3340 14890 3352
rect 15197 3349 15209 3352
rect 15243 3349 15255 3383
rect 15197 3343 15255 3349
rect 92 3290 15824 3312
rect 92 3238 1904 3290
rect 1956 3238 1968 3290
rect 2020 3238 2032 3290
rect 2084 3238 2096 3290
rect 2148 3238 2160 3290
rect 2212 3238 5837 3290
rect 5889 3238 5901 3290
rect 5953 3238 5965 3290
rect 6017 3238 6029 3290
rect 6081 3238 6093 3290
rect 6145 3238 9770 3290
rect 9822 3238 9834 3290
rect 9886 3238 9898 3290
rect 9950 3238 9962 3290
rect 10014 3238 10026 3290
rect 10078 3238 13703 3290
rect 13755 3238 13767 3290
rect 13819 3238 13831 3290
rect 13883 3238 13895 3290
rect 13947 3238 13959 3290
rect 14011 3238 15824 3290
rect 92 3216 15824 3238
rect 569 3179 627 3185
rect 569 3145 581 3179
rect 615 3176 627 3179
rect 615 3148 2774 3176
rect 615 3145 627 3148
rect 569 3139 627 3145
rect 2746 3108 2774 3148
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 3510 3176 3516 3188
rect 3200 3148 3516 3176
rect 3200 3136 3206 3148
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 4985 3179 5043 3185
rect 4985 3145 4997 3179
rect 5031 3176 5043 3179
rect 5074 3176 5080 3188
rect 5031 3148 5080 3176
rect 5031 3145 5043 3148
rect 4985 3139 5043 3145
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5169 3179 5227 3185
rect 5169 3145 5181 3179
rect 5215 3176 5227 3179
rect 7282 3176 7288 3188
rect 5215 3148 7288 3176
rect 5215 3145 5227 3148
rect 5169 3139 5227 3145
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 9493 3179 9551 3185
rect 9493 3176 9505 3179
rect 8628 3148 9505 3176
rect 8628 3136 8634 3148
rect 9493 3145 9505 3148
rect 9539 3176 9551 3179
rect 9582 3176 9588 3188
rect 9539 3148 9588 3176
rect 9539 3145 9551 3148
rect 9493 3139 9551 3145
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 10226 3136 10232 3188
rect 10284 3136 10290 3188
rect 10870 3136 10876 3188
rect 10928 3136 10934 3188
rect 13446 3136 13452 3188
rect 13504 3136 13510 3188
rect 13538 3136 13544 3188
rect 13596 3176 13602 3188
rect 13817 3179 13875 3185
rect 13817 3176 13829 3179
rect 13596 3148 13829 3176
rect 13596 3136 13602 3148
rect 13817 3145 13829 3148
rect 13863 3145 13875 3179
rect 13817 3139 13875 3145
rect 14826 3136 14832 3188
rect 14884 3136 14890 3188
rect 14921 3179 14979 3185
rect 14921 3145 14933 3179
rect 14967 3176 14979 3179
rect 15286 3176 15292 3188
rect 14967 3148 15292 3176
rect 14967 3145 14979 3148
rect 14921 3139 14979 3145
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 15381 3179 15439 3185
rect 15381 3145 15393 3179
rect 15427 3176 15439 3179
rect 15470 3176 15476 3188
rect 15427 3148 15476 3176
rect 15427 3145 15439 3148
rect 15381 3139 15439 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 4062 3108 4068 3120
rect 2746 3080 4068 3108
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 4172 3080 7403 3108
rect 4172 3040 4200 3080
rect 3344 3012 4200 3040
rect 5997 3043 6055 3049
rect 3344 2984 3372 3012
rect 5997 3009 6009 3043
rect 6043 3040 6055 3043
rect 7282 3040 7288 3052
rect 6043 3012 7288 3040
rect 6043 3009 6055 3012
rect 5997 3003 6055 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 382 2932 388 2984
rect 440 2932 446 2984
rect 3326 2932 3332 2984
rect 3384 2932 3390 2984
rect 3878 2932 3884 2984
rect 3936 2972 3942 2984
rect 4617 2975 4675 2981
rect 4617 2972 4629 2975
rect 3936 2944 4629 2972
rect 3936 2932 3942 2944
rect 4617 2941 4629 2944
rect 4663 2972 4675 2975
rect 5166 2972 5172 2984
rect 4663 2944 5172 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 5258 2932 5264 2984
rect 5316 2972 5322 2984
rect 6178 2972 6184 2984
rect 5316 2944 6184 2972
rect 5316 2932 5322 2944
rect 6178 2932 6184 2944
rect 6236 2972 6242 2984
rect 6273 2975 6331 2981
rect 6273 2972 6285 2975
rect 6236 2944 6285 2972
rect 6236 2932 6242 2944
rect 6273 2941 6285 2944
rect 6319 2972 6331 2975
rect 7006 2972 7012 2984
rect 6319 2944 7012 2972
rect 6319 2941 6331 2944
rect 6273 2935 6331 2941
rect 7006 2932 7012 2944
rect 7064 2932 7070 2984
rect 4433 2907 4491 2913
rect 4433 2873 4445 2907
rect 4479 2873 4491 2907
rect 4433 2867 4491 2873
rect 4448 2836 4476 2867
rect 4706 2864 4712 2916
rect 4764 2904 4770 2916
rect 4994 2907 5052 2913
rect 4994 2904 5006 2907
rect 4764 2876 5006 2904
rect 4764 2864 4770 2876
rect 4994 2873 5006 2876
rect 5040 2873 5052 2907
rect 7375 2904 7403 3080
rect 8846 3068 8852 3120
rect 8904 3108 8910 3120
rect 10597 3111 10655 3117
rect 10597 3108 10609 3111
rect 8904 3080 10609 3108
rect 8904 3068 8910 3080
rect 10597 3077 10609 3080
rect 10643 3077 10655 3111
rect 10888 3108 10916 3136
rect 10888 3080 11468 3108
rect 10597 3071 10655 3077
rect 8938 3000 8944 3052
rect 8996 3000 9002 3052
rect 10686 3000 10692 3052
rect 10744 3040 10750 3052
rect 10744 3012 11376 3040
rect 10744 3000 10750 3012
rect 8202 2932 8208 2984
rect 8260 2932 8266 2984
rect 8956 2972 8984 3000
rect 10781 2975 10839 2981
rect 10781 2972 10793 2975
rect 8956 2944 10793 2972
rect 10781 2941 10793 2944
rect 10827 2941 10839 2975
rect 10781 2935 10839 2941
rect 11057 2975 11115 2981
rect 11057 2941 11069 2975
rect 11103 2972 11115 2975
rect 11146 2972 11152 2984
rect 11103 2944 11152 2972
rect 11103 2941 11115 2944
rect 11057 2935 11115 2941
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 9490 2904 9496 2916
rect 7375 2876 9496 2904
rect 4994 2867 5052 2873
rect 9490 2864 9496 2876
rect 9548 2904 9554 2916
rect 10137 2907 10195 2913
rect 10137 2904 10149 2907
rect 9548 2876 10149 2904
rect 9548 2864 9554 2876
rect 10137 2873 10149 2876
rect 10183 2873 10195 2907
rect 10137 2867 10195 2873
rect 10870 2864 10876 2916
rect 10928 2904 10934 2916
rect 11348 2913 11376 3012
rect 11440 2981 11468 3080
rect 11425 2975 11483 2981
rect 11425 2941 11437 2975
rect 11471 2941 11483 2975
rect 11425 2935 11483 2941
rect 11241 2907 11299 2913
rect 11241 2904 11253 2907
rect 10928 2876 11253 2904
rect 10928 2864 10934 2876
rect 11241 2873 11253 2876
rect 11287 2873 11299 2907
rect 11241 2867 11299 2873
rect 11333 2907 11391 2913
rect 11333 2873 11345 2907
rect 11379 2904 11391 2907
rect 13170 2904 13176 2916
rect 11379 2876 13176 2904
rect 11379 2873 11391 2876
rect 11333 2867 11391 2873
rect 13170 2864 13176 2876
rect 13228 2864 13234 2916
rect 5626 2836 5632 2848
rect 4448 2808 5632 2836
rect 5626 2796 5632 2808
rect 5684 2836 5690 2848
rect 7742 2836 7748 2848
rect 5684 2808 7748 2836
rect 5684 2796 5690 2808
rect 7742 2796 7748 2808
rect 7800 2796 7806 2848
rect 9582 2796 9588 2848
rect 9640 2836 9646 2848
rect 11422 2836 11428 2848
rect 9640 2808 11428 2836
rect 9640 2796 9646 2808
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 11606 2796 11612 2848
rect 11664 2796 11670 2848
rect 13464 2836 13492 3136
rect 14844 3040 14872 3136
rect 14016 3012 14872 3040
rect 14016 2981 14044 3012
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2941 14059 2975
rect 14001 2935 14059 2941
rect 14277 2975 14335 2981
rect 14277 2941 14289 2975
rect 14323 2972 14335 2975
rect 14366 2972 14372 2984
rect 14323 2944 14372 2972
rect 14323 2941 14335 2944
rect 14277 2935 14335 2941
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2972 14795 2975
rect 14844 2972 14872 3012
rect 14783 2944 14872 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 15010 2932 15016 2984
rect 15068 2972 15074 2984
rect 15105 2975 15163 2981
rect 15105 2972 15117 2975
rect 15068 2944 15117 2972
rect 15068 2932 15074 2944
rect 15105 2941 15117 2944
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 14553 2907 14611 2913
rect 14553 2873 14565 2907
rect 14599 2873 14611 2907
rect 14553 2867 14611 2873
rect 14185 2839 14243 2845
rect 14185 2836 14197 2839
rect 13464 2808 14197 2836
rect 14185 2805 14197 2808
rect 14231 2836 14243 2839
rect 14568 2836 14596 2867
rect 14231 2808 14596 2836
rect 14231 2805 14243 2808
rect 14185 2799 14243 2805
rect 92 2746 15824 2768
rect 92 2694 2564 2746
rect 2616 2694 2628 2746
rect 2680 2694 2692 2746
rect 2744 2694 2756 2746
rect 2808 2694 2820 2746
rect 2872 2694 6497 2746
rect 6549 2694 6561 2746
rect 6613 2694 6625 2746
rect 6677 2694 6689 2746
rect 6741 2694 6753 2746
rect 6805 2694 10430 2746
rect 10482 2694 10494 2746
rect 10546 2694 10558 2746
rect 10610 2694 10622 2746
rect 10674 2694 10686 2746
rect 10738 2694 14363 2746
rect 14415 2694 14427 2746
rect 14479 2694 14491 2746
rect 14543 2694 14555 2746
rect 14607 2694 14619 2746
rect 14671 2694 15824 2746
rect 92 2672 15824 2694
rect 3878 2592 3884 2644
rect 3936 2592 3942 2644
rect 6641 2635 6699 2641
rect 6641 2601 6653 2635
rect 6687 2632 6699 2635
rect 6822 2632 6828 2644
rect 6687 2604 6828 2632
rect 6687 2601 6699 2604
rect 6641 2595 6699 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 9582 2632 9588 2644
rect 8496 2604 9588 2632
rect 2406 2524 2412 2576
rect 2464 2524 2470 2576
rect 3510 2456 3516 2508
rect 3568 2496 3574 2508
rect 7006 2496 7012 2508
rect 3568 2468 7012 2496
rect 3568 2456 3574 2468
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 8496 2505 8524 2604
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10275 2604 11008 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10870 2524 10876 2576
rect 10928 2524 10934 2576
rect 10980 2564 11008 2604
rect 13170 2592 13176 2644
rect 13228 2592 13234 2644
rect 11146 2564 11152 2576
rect 10980 2536 11152 2564
rect 8389 2499 8447 2505
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 8435 2468 8493 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 8481 2465 8493 2468
rect 8527 2465 8539 2499
rect 10226 2496 10232 2508
rect 9890 2468 10232 2496
rect 8481 2459 8539 2465
rect 10226 2456 10232 2468
rect 10284 2456 10290 2508
rect 10318 2456 10324 2508
rect 10376 2496 10382 2508
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 10376 2468 10701 2496
rect 10376 2456 10382 2468
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 10689 2459 10747 2465
rect 10781 2499 10839 2505
rect 10781 2465 10793 2499
rect 10827 2496 10839 2499
rect 10980 2496 11008 2536
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 11698 2524 11704 2576
rect 11756 2524 11762 2576
rect 13188 2564 13216 2592
rect 14553 2567 14611 2573
rect 14553 2564 14565 2567
rect 13188 2536 14565 2564
rect 14553 2533 14565 2536
rect 14599 2533 14611 2567
rect 14553 2527 14611 2533
rect 14918 2524 14924 2576
rect 14976 2564 14982 2576
rect 15105 2567 15163 2573
rect 15105 2564 15117 2567
rect 14976 2536 15117 2564
rect 14976 2524 14982 2536
rect 15105 2533 15117 2536
rect 15151 2564 15163 2567
rect 15194 2564 15200 2576
rect 15151 2536 15200 2564
rect 15151 2533 15163 2536
rect 15105 2527 15163 2533
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 10827 2468 11008 2496
rect 11057 2499 11115 2505
rect 10827 2465 10839 2468
rect 10781 2459 10839 2465
rect 11057 2465 11069 2499
rect 11103 2496 11115 2499
rect 11238 2496 11244 2508
rect 11103 2468 11244 2496
rect 11103 2465 11115 2468
rect 11057 2459 11115 2465
rect 11238 2456 11244 2468
rect 11296 2456 11302 2508
rect 11422 2456 11428 2508
rect 11480 2456 11486 2508
rect 12710 2456 12716 2508
rect 12768 2496 12774 2508
rect 13446 2496 13452 2508
rect 12768 2468 13452 2496
rect 12768 2456 12774 2468
rect 13446 2456 13452 2468
rect 13504 2456 13510 2508
rect 13538 2456 13544 2508
rect 13596 2456 13602 2508
rect 14461 2499 14519 2505
rect 14461 2465 14473 2499
rect 14507 2496 14519 2499
rect 14642 2496 14648 2508
rect 14507 2468 14648 2496
rect 14507 2465 14519 2468
rect 14461 2459 14519 2465
rect 14642 2456 14648 2468
rect 14700 2456 14706 2508
rect 14737 2499 14795 2505
rect 14737 2465 14749 2499
rect 14783 2496 14795 2499
rect 14783 2468 14872 2496
rect 14783 2465 14795 2468
rect 14737 2459 14795 2465
rect 1762 2388 1768 2440
rect 1820 2428 1826 2440
rect 2133 2431 2191 2437
rect 2133 2428 2145 2431
rect 1820 2400 2145 2428
rect 1820 2388 1826 2400
rect 2133 2397 2145 2400
rect 2179 2428 2191 2431
rect 2179 2400 2268 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2240 2292 2268 2400
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7616 2400 8125 2428
rect 7616 2388 7622 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 8803 2400 10548 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 10520 2369 10548 2400
rect 10505 2363 10563 2369
rect 3528 2332 4476 2360
rect 3528 2292 3556 2332
rect 4448 2304 4476 2332
rect 10505 2329 10517 2363
rect 10551 2329 10563 2363
rect 10505 2323 10563 2329
rect 14844 2304 14872 2468
rect 2240 2264 3556 2292
rect 4430 2252 4436 2304
rect 4488 2252 4494 2304
rect 13354 2252 13360 2304
rect 13412 2252 13418 2304
rect 14274 2252 14280 2304
rect 14332 2252 14338 2304
rect 14826 2252 14832 2304
rect 14884 2252 14890 2304
rect 14918 2252 14924 2304
rect 14976 2252 14982 2304
rect 15378 2252 15384 2304
rect 15436 2252 15442 2304
rect 92 2202 15824 2224
rect 92 2150 1904 2202
rect 1956 2150 1968 2202
rect 2020 2150 2032 2202
rect 2084 2150 2096 2202
rect 2148 2150 2160 2202
rect 2212 2150 5837 2202
rect 5889 2150 5901 2202
rect 5953 2150 5965 2202
rect 6017 2150 6029 2202
rect 6081 2150 6093 2202
rect 6145 2150 9770 2202
rect 9822 2150 9834 2202
rect 9886 2150 9898 2202
rect 9950 2150 9962 2202
rect 10014 2150 10026 2202
rect 10078 2150 13703 2202
rect 13755 2150 13767 2202
rect 13819 2150 13831 2202
rect 13883 2150 13895 2202
rect 13947 2150 13959 2202
rect 14011 2150 15824 2202
rect 92 2128 15824 2150
rect 4062 2048 4068 2100
rect 4120 2088 4126 2100
rect 7926 2088 7932 2100
rect 4120 2060 7932 2088
rect 4120 2048 4126 2060
rect 7926 2048 7932 2060
rect 7984 2048 7990 2100
rect 13538 2048 13544 2100
rect 13596 2088 13602 2100
rect 13633 2091 13691 2097
rect 13633 2088 13645 2091
rect 13596 2060 13645 2088
rect 13596 2048 13602 2060
rect 13633 2057 13645 2060
rect 13679 2057 13691 2091
rect 13633 2051 13691 2057
rect 14274 2048 14280 2100
rect 14332 2048 14338 2100
rect 14918 2048 14924 2100
rect 14976 2048 14982 2100
rect 15194 2048 15200 2100
rect 15252 2048 15258 2100
rect 6178 1980 6184 2032
rect 6236 1980 6242 2032
rect 7006 1980 7012 2032
rect 7064 1980 7070 2032
rect 4430 1912 4436 1964
rect 4488 1912 4494 1964
rect 4706 1912 4712 1964
rect 4764 1912 4770 1964
rect 7024 1884 7052 1980
rect 9582 1912 9588 1964
rect 9640 1912 9646 1964
rect 13262 1952 13268 1964
rect 12452 1924 13268 1952
rect 12452 1896 12480 1924
rect 13262 1912 13268 1924
rect 13320 1912 13326 1964
rect 5842 1856 7052 1884
rect 12434 1844 12440 1896
rect 12492 1844 12498 1896
rect 12710 1844 12716 1896
rect 12768 1844 12774 1896
rect 13170 1844 13176 1896
rect 13228 1844 13234 1896
rect 14292 1893 14320 2048
rect 13449 1887 13507 1893
rect 13449 1853 13461 1887
rect 13495 1884 13507 1887
rect 13817 1887 13875 1893
rect 13817 1884 13829 1887
rect 13495 1856 13829 1884
rect 13495 1853 13507 1856
rect 13449 1847 13507 1853
rect 13817 1853 13829 1856
rect 13863 1853 13875 1887
rect 13817 1847 13875 1853
rect 14001 1887 14059 1893
rect 14001 1853 14013 1887
rect 14047 1853 14059 1887
rect 14001 1847 14059 1853
rect 14277 1887 14335 1893
rect 14277 1853 14289 1887
rect 14323 1853 14335 1887
rect 14277 1847 14335 1853
rect 9858 1776 9864 1828
rect 9916 1776 9922 1828
rect 12728 1816 12756 1844
rect 11086 1788 12756 1816
rect 10226 1708 10232 1760
rect 10284 1748 10290 1760
rect 11164 1748 11192 1788
rect 10284 1720 11192 1748
rect 10284 1708 10290 1720
rect 11330 1708 11336 1760
rect 11388 1708 11394 1760
rect 13188 1748 13216 1844
rect 14016 1816 14044 1847
rect 14366 1844 14372 1896
rect 14424 1844 14430 1896
rect 14826 1844 14832 1896
rect 14884 1844 14890 1896
rect 14936 1884 14964 2048
rect 15013 1887 15071 1893
rect 15013 1884 15025 1887
rect 14936 1856 15025 1884
rect 15013 1853 15025 1856
rect 15059 1853 15071 1887
rect 15013 1847 15071 1853
rect 14844 1816 14872 1844
rect 14016 1788 14872 1816
rect 14185 1751 14243 1757
rect 14185 1748 14197 1751
rect 13188 1720 14197 1748
rect 14185 1717 14197 1720
rect 14231 1717 14243 1751
rect 14185 1711 14243 1717
rect 14274 1708 14280 1760
rect 14332 1748 14338 1760
rect 14461 1751 14519 1757
rect 14461 1748 14473 1751
rect 14332 1720 14473 1748
rect 14332 1708 14338 1720
rect 14461 1717 14473 1720
rect 14507 1717 14519 1751
rect 14461 1711 14519 1717
rect 92 1658 15824 1680
rect 92 1606 2564 1658
rect 2616 1606 2628 1658
rect 2680 1606 2692 1658
rect 2744 1606 2756 1658
rect 2808 1606 2820 1658
rect 2872 1606 6497 1658
rect 6549 1606 6561 1658
rect 6613 1606 6625 1658
rect 6677 1606 6689 1658
rect 6741 1606 6753 1658
rect 6805 1606 10430 1658
rect 10482 1606 10494 1658
rect 10546 1606 10558 1658
rect 10610 1606 10622 1658
rect 10674 1606 10686 1658
rect 10738 1606 14363 1658
rect 14415 1606 14427 1658
rect 14479 1606 14491 1658
rect 14543 1606 14555 1658
rect 14607 1606 14619 1658
rect 14671 1606 15824 1658
rect 92 1584 15824 1606
rect 9858 1504 9864 1556
rect 9916 1544 9922 1556
rect 10137 1547 10195 1553
rect 10137 1544 10149 1547
rect 9916 1516 10149 1544
rect 9916 1504 9922 1516
rect 10137 1513 10149 1516
rect 10183 1513 10195 1547
rect 10137 1507 10195 1513
rect 10873 1547 10931 1553
rect 10873 1513 10885 1547
rect 10919 1544 10931 1547
rect 11146 1544 11152 1556
rect 10919 1516 11152 1544
rect 10919 1513 10931 1516
rect 10873 1507 10931 1513
rect 11146 1504 11152 1516
rect 11204 1504 11210 1556
rect 11330 1504 11336 1556
rect 11388 1504 11394 1556
rect 14826 1504 14832 1556
rect 14884 1504 14890 1556
rect 11348 1476 11376 1504
rect 11425 1479 11483 1485
rect 11425 1476 11437 1479
rect 10704 1448 11437 1476
rect 1394 1368 1400 1420
rect 1452 1368 1458 1420
rect 3142 1368 3148 1420
rect 3200 1368 3206 1420
rect 8757 1411 8815 1417
rect 8757 1377 8769 1411
rect 8803 1408 8815 1411
rect 9030 1408 9036 1420
rect 8803 1380 9036 1408
rect 8803 1377 8815 1380
rect 8757 1371 8815 1377
rect 9030 1368 9036 1380
rect 9088 1368 9094 1420
rect 10704 1417 10732 1448
rect 11425 1445 11437 1448
rect 11471 1445 11483 1479
rect 11425 1439 11483 1445
rect 13354 1436 13360 1488
rect 13412 1436 13418 1488
rect 13446 1436 13452 1488
rect 13504 1476 13510 1488
rect 13504 1448 13846 1476
rect 13504 1436 13510 1448
rect 15102 1436 15108 1488
rect 15160 1436 15166 1488
rect 9861 1411 9919 1417
rect 9861 1377 9873 1411
rect 9907 1377 9919 1411
rect 9861 1371 9919 1377
rect 10045 1411 10103 1417
rect 10045 1377 10057 1411
rect 10091 1408 10103 1411
rect 10321 1411 10379 1417
rect 10321 1408 10333 1411
rect 10091 1380 10333 1408
rect 10091 1377 10103 1380
rect 10045 1371 10103 1377
rect 10321 1377 10333 1380
rect 10367 1377 10379 1411
rect 10321 1371 10379 1377
rect 10689 1411 10747 1417
rect 10689 1377 10701 1411
rect 10735 1377 10747 1411
rect 10689 1371 10747 1377
rect 9674 1300 9680 1352
rect 9732 1300 9738 1352
rect 9876 1340 9904 1371
rect 10962 1368 10968 1420
rect 11020 1368 11026 1420
rect 11146 1368 11152 1420
rect 11204 1408 11210 1420
rect 11241 1411 11299 1417
rect 11241 1408 11253 1411
rect 11204 1380 11253 1408
rect 11204 1368 11210 1380
rect 11241 1377 11253 1380
rect 11287 1377 11299 1411
rect 12434 1408 12440 1420
rect 11241 1371 11299 1377
rect 12406 1368 12440 1408
rect 12492 1368 12498 1420
rect 10505 1343 10563 1349
rect 10505 1340 10517 1343
rect 9876 1312 10517 1340
rect 10505 1309 10517 1312
rect 10551 1309 10563 1343
rect 12406 1340 12434 1368
rect 10505 1303 10563 1309
rect 10612 1312 12434 1340
rect 9692 1272 9720 1300
rect 10612 1272 10640 1312
rect 13078 1300 13084 1352
rect 13136 1300 13142 1352
rect 9692 1244 10640 1272
rect 1302 1164 1308 1216
rect 1360 1164 1366 1216
rect 3050 1164 3056 1216
rect 3108 1164 3114 1216
rect 8662 1164 8668 1216
rect 8720 1164 8726 1216
rect 11606 1164 11612 1216
rect 11664 1164 11670 1216
rect 15378 1164 15384 1216
rect 15436 1164 15442 1216
rect 92 1114 15824 1136
rect 92 1062 1904 1114
rect 1956 1062 1968 1114
rect 2020 1062 2032 1114
rect 2084 1062 2096 1114
rect 2148 1062 2160 1114
rect 2212 1062 5837 1114
rect 5889 1062 5901 1114
rect 5953 1062 5965 1114
rect 6017 1062 6029 1114
rect 6081 1062 6093 1114
rect 6145 1062 9770 1114
rect 9822 1062 9834 1114
rect 9886 1062 9898 1114
rect 9950 1062 9962 1114
rect 10014 1062 10026 1114
rect 10078 1062 13703 1114
rect 13755 1062 13767 1114
rect 13819 1062 13831 1114
rect 13883 1062 13895 1114
rect 13947 1062 13959 1114
rect 14011 1062 15824 1114
rect 92 1040 15824 1062
rect 569 1003 627 1009
rect 569 969 581 1003
rect 615 1000 627 1003
rect 3326 1000 3332 1012
rect 615 972 3332 1000
rect 615 969 627 972
rect 569 963 627 969
rect 3326 960 3332 972
rect 3384 960 3390 1012
rect 11606 960 11612 1012
rect 11664 1000 11670 1012
rect 11664 972 12434 1000
rect 11664 960 11670 972
rect 12406 864 12434 972
rect 15102 960 15108 1012
rect 15160 960 15166 1012
rect 12406 836 14964 864
rect 382 756 388 808
rect 440 756 446 808
rect 1302 756 1308 808
rect 1360 796 1366 808
rect 1489 799 1547 805
rect 1489 796 1501 799
rect 1360 768 1501 796
rect 1360 756 1366 768
rect 1489 765 1501 768
rect 1535 765 1547 799
rect 1489 759 1547 765
rect 3050 756 3056 808
rect 3108 756 3114 808
rect 4982 756 4988 808
rect 5040 796 5046 808
rect 5445 799 5503 805
rect 5445 796 5457 799
rect 5040 768 5457 796
rect 5040 756 5046 768
rect 5445 765 5457 768
rect 5491 765 5503 799
rect 5445 759 5503 765
rect 6362 756 6368 808
rect 6420 796 6426 808
rect 7009 799 7067 805
rect 7009 796 7021 799
rect 6420 768 7021 796
rect 6420 756 6426 768
rect 7009 765 7021 768
rect 7055 765 7067 799
rect 7009 759 7067 765
rect 8662 756 8668 808
rect 8720 796 8726 808
rect 8757 799 8815 805
rect 8757 796 8769 799
rect 8720 768 8769 796
rect 8720 756 8726 768
rect 8757 765 8769 768
rect 8803 765 8815 799
rect 8757 759 8815 765
rect 10965 799 11023 805
rect 10965 765 10977 799
rect 11011 765 11023 799
rect 10965 759 11023 765
rect 10980 728 11008 759
rect 11054 756 11060 808
rect 11112 756 11118 808
rect 12618 756 12624 808
rect 12676 756 12682 808
rect 14274 756 14280 808
rect 14332 796 14338 808
rect 14936 805 14964 836
rect 14461 799 14519 805
rect 14461 796 14473 799
rect 14332 768 14473 796
rect 14332 756 14338 768
rect 14461 765 14473 768
rect 14507 765 14519 799
rect 14461 759 14519 765
rect 14921 799 14979 805
rect 14921 765 14933 799
rect 14967 765 14979 799
rect 14921 759 14979 765
rect 11149 731 11207 737
rect 11149 728 11161 731
rect 10980 700 11161 728
rect 11149 697 11161 700
rect 11195 697 11207 731
rect 11149 691 11207 697
rect 1302 620 1308 672
rect 1360 620 1366 672
rect 3234 620 3240 672
rect 3292 620 3298 672
rect 5258 620 5264 672
rect 5316 660 5322 672
rect 5537 663 5595 669
rect 5537 660 5549 663
rect 5316 632 5549 660
rect 5316 620 5322 632
rect 5537 629 5549 632
rect 5583 629 5595 663
rect 5537 623 5595 629
rect 7098 620 7104 672
rect 7156 620 7162 672
rect 8938 620 8944 672
rect 8996 620 9002 672
rect 10778 620 10784 672
rect 10836 620 10842 672
rect 12802 620 12808 672
rect 12860 620 12866 672
rect 14645 663 14703 669
rect 14645 629 14657 663
rect 14691 660 14703 663
rect 14734 660 14740 672
rect 14691 632 14740 660
rect 14691 629 14703 632
rect 14645 623 14703 629
rect 14734 620 14740 632
rect 14792 620 14798 672
rect 92 570 15824 592
rect 92 518 2564 570
rect 2616 518 2628 570
rect 2680 518 2692 570
rect 2744 518 2756 570
rect 2808 518 2820 570
rect 2872 518 6497 570
rect 6549 518 6561 570
rect 6613 518 6625 570
rect 6677 518 6689 570
rect 6741 518 6753 570
rect 6805 518 10430 570
rect 10482 518 10494 570
rect 10546 518 10558 570
rect 10610 518 10622 570
rect 10674 518 10686 570
rect 10738 518 14363 570
rect 14415 518 14427 570
rect 14479 518 14491 570
rect 14543 518 14555 570
rect 14607 518 14619 570
rect 14671 518 15824 570
rect 92 496 15824 518
<< via1 >>
rect 1904 13030 1956 13082
rect 1968 13030 2020 13082
rect 2032 13030 2084 13082
rect 2096 13030 2148 13082
rect 2160 13030 2212 13082
rect 5837 13030 5889 13082
rect 5901 13030 5953 13082
rect 5965 13030 6017 13082
rect 6029 13030 6081 13082
rect 6093 13030 6145 13082
rect 9770 13030 9822 13082
rect 9834 13030 9886 13082
rect 9898 13030 9950 13082
rect 9962 13030 10014 13082
rect 10026 13030 10078 13082
rect 13703 13030 13755 13082
rect 13767 13030 13819 13082
rect 13831 13030 13883 13082
rect 13895 13030 13947 13082
rect 13959 13030 14011 13082
rect 848 12928 900 12980
rect 1124 12971 1176 12980
rect 1124 12937 1133 12971
rect 1133 12937 1167 12971
rect 1167 12937 1176 12971
rect 1124 12928 1176 12937
rect 3240 12928 3292 12980
rect 5264 12928 5316 12980
rect 6644 12928 6696 12980
rect 8944 12928 8996 12980
rect 10876 12928 10928 12980
rect 12808 12971 12860 12980
rect 12808 12937 12817 12971
rect 12817 12937 12851 12971
rect 12851 12937 12860 12971
rect 12808 12928 12860 12937
rect 14648 12971 14700 12980
rect 14648 12937 14657 12971
rect 14657 12937 14691 12971
rect 14691 12937 14700 12971
rect 14648 12928 14700 12937
rect 15476 12928 15528 12980
rect 2320 12724 2372 12776
rect 3240 12724 3292 12776
rect 388 12699 440 12708
rect 388 12665 397 12699
rect 397 12665 431 12699
rect 431 12665 440 12699
rect 388 12656 440 12665
rect 1308 12656 1360 12708
rect 1400 12699 1452 12708
rect 1400 12665 1409 12699
rect 1409 12665 1443 12699
rect 1443 12665 1452 12699
rect 1400 12656 1452 12665
rect 3332 12588 3384 12640
rect 3516 12631 3568 12640
rect 3516 12597 3525 12631
rect 3525 12597 3559 12631
rect 3559 12597 3568 12631
rect 3516 12588 3568 12597
rect 5816 12724 5868 12776
rect 9036 12767 9088 12776
rect 9036 12733 9045 12767
rect 9045 12733 9079 12767
rect 9079 12733 9088 12767
rect 9036 12724 9088 12733
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 12348 12724 12400 12776
rect 14096 12724 14148 12776
rect 5448 12699 5500 12708
rect 5448 12665 5457 12699
rect 5457 12665 5491 12699
rect 5491 12665 5500 12699
rect 5448 12656 5500 12665
rect 15108 12699 15160 12708
rect 15108 12665 15117 12699
rect 15117 12665 15151 12699
rect 15151 12665 15160 12699
rect 15108 12656 15160 12665
rect 5540 12588 5592 12640
rect 6828 12588 6880 12640
rect 2564 12486 2616 12538
rect 2628 12486 2680 12538
rect 2692 12486 2744 12538
rect 2756 12486 2808 12538
rect 2820 12486 2872 12538
rect 6497 12486 6549 12538
rect 6561 12486 6613 12538
rect 6625 12486 6677 12538
rect 6689 12486 6741 12538
rect 6753 12486 6805 12538
rect 10430 12486 10482 12538
rect 10494 12486 10546 12538
rect 10558 12486 10610 12538
rect 10622 12486 10674 12538
rect 10686 12486 10738 12538
rect 14363 12486 14415 12538
rect 14427 12486 14479 12538
rect 14491 12486 14543 12538
rect 14555 12486 14607 12538
rect 14619 12486 14671 12538
rect 3056 12384 3108 12436
rect 756 12316 808 12368
rect 1492 12316 1544 12368
rect 2412 12316 2464 12368
rect 3700 12359 3752 12368
rect 3700 12325 3709 12359
rect 3709 12325 3743 12359
rect 3743 12325 3752 12359
rect 3700 12316 3752 12325
rect 4160 12316 4212 12368
rect 848 12223 900 12232
rect 848 12189 857 12223
rect 857 12189 891 12223
rect 891 12189 900 12223
rect 848 12180 900 12189
rect 5540 12384 5592 12436
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 5816 12427 5868 12436
rect 5816 12393 5825 12427
rect 5825 12393 5859 12427
rect 5859 12393 5868 12427
rect 5816 12384 5868 12393
rect 15108 12384 15160 12436
rect 3424 12180 3476 12189
rect 5632 12180 5684 12232
rect 6184 12180 6236 12232
rect 7748 12248 7800 12300
rect 6368 12223 6420 12232
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 15108 12291 15160 12300
rect 15108 12257 15117 12291
rect 15117 12257 15151 12291
rect 15151 12257 15160 12291
rect 15108 12248 15160 12257
rect 6368 12180 6420 12189
rect 15200 12180 15252 12232
rect 2320 12087 2372 12096
rect 2320 12053 2329 12087
rect 2329 12053 2363 12087
rect 2363 12053 2372 12087
rect 2320 12044 2372 12053
rect 3148 12087 3200 12096
rect 3148 12053 3157 12087
rect 3157 12053 3191 12087
rect 3191 12053 3200 12087
rect 3148 12044 3200 12053
rect 8024 12044 8076 12096
rect 15384 12087 15436 12096
rect 15384 12053 15393 12087
rect 15393 12053 15427 12087
rect 15427 12053 15436 12087
rect 15384 12044 15436 12053
rect 1904 11942 1956 11994
rect 1968 11942 2020 11994
rect 2032 11942 2084 11994
rect 2096 11942 2148 11994
rect 2160 11942 2212 11994
rect 5837 11942 5889 11994
rect 5901 11942 5953 11994
rect 5965 11942 6017 11994
rect 6029 11942 6081 11994
rect 6093 11942 6145 11994
rect 9770 11942 9822 11994
rect 9834 11942 9886 11994
rect 9898 11942 9950 11994
rect 9962 11942 10014 11994
rect 10026 11942 10078 11994
rect 13703 11942 13755 11994
rect 13767 11942 13819 11994
rect 13831 11942 13883 11994
rect 13895 11942 13947 11994
rect 13959 11942 14011 11994
rect 848 11840 900 11892
rect 1308 11840 1360 11892
rect 3056 11840 3108 11892
rect 3148 11840 3200 11892
rect 3332 11883 3384 11892
rect 3332 11849 3341 11883
rect 3341 11849 3375 11883
rect 3375 11849 3384 11883
rect 3332 11840 3384 11849
rect 4068 11840 4120 11892
rect 1124 11636 1176 11688
rect 1584 11636 1636 11688
rect 2320 11568 2372 11620
rect 480 11543 532 11552
rect 480 11509 489 11543
rect 489 11509 523 11543
rect 523 11509 532 11543
rect 480 11500 532 11509
rect 1768 11500 1820 11552
rect 2412 11500 2464 11552
rect 2964 11568 3016 11620
rect 4068 11636 4120 11688
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 5448 11636 5500 11688
rect 5724 11636 5776 11688
rect 6000 11679 6052 11688
rect 6000 11645 6009 11679
rect 6009 11645 6043 11679
rect 6043 11645 6052 11679
rect 6000 11636 6052 11645
rect 6736 11679 6788 11688
rect 6736 11645 6745 11679
rect 6745 11645 6779 11679
rect 6779 11645 6788 11679
rect 6736 11636 6788 11645
rect 8024 11611 8076 11620
rect 8024 11577 8033 11611
rect 8033 11577 8067 11611
rect 8067 11577 8076 11611
rect 8024 11568 8076 11577
rect 8484 11568 8536 11620
rect 4896 11543 4948 11552
rect 4896 11509 4905 11543
rect 4905 11509 4939 11543
rect 4939 11509 4948 11543
rect 4896 11500 4948 11509
rect 6276 11500 6328 11552
rect 9036 11500 9088 11552
rect 2564 11398 2616 11450
rect 2628 11398 2680 11450
rect 2692 11398 2744 11450
rect 2756 11398 2808 11450
rect 2820 11398 2872 11450
rect 6497 11398 6549 11450
rect 6561 11398 6613 11450
rect 6625 11398 6677 11450
rect 6689 11398 6741 11450
rect 6753 11398 6805 11450
rect 10430 11398 10482 11450
rect 10494 11398 10546 11450
rect 10558 11398 10610 11450
rect 10622 11398 10674 11450
rect 10686 11398 10738 11450
rect 14363 11398 14415 11450
rect 14427 11398 14479 11450
rect 14491 11398 14543 11450
rect 14555 11398 14607 11450
rect 14619 11398 14671 11450
rect 2964 11296 3016 11348
rect 5632 11296 5684 11348
rect 756 11228 808 11280
rect 1492 11228 1544 11280
rect 2412 11228 2464 11280
rect 4160 11228 4212 11280
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 15108 11296 15160 11348
rect 7748 11228 7800 11280
rect 848 11135 900 11144
rect 848 11101 857 11135
rect 857 11101 891 11135
rect 891 11101 900 11135
rect 848 11092 900 11101
rect 2872 11160 2924 11212
rect 2596 10999 2648 11008
rect 2596 10965 2605 10999
rect 2605 10965 2639 10999
rect 2639 10965 2648 10999
rect 2596 10956 2648 10965
rect 5632 11160 5684 11212
rect 6000 11160 6052 11212
rect 6460 11160 6512 11212
rect 14924 11203 14976 11212
rect 14924 11169 14933 11203
rect 14933 11169 14967 11203
rect 14967 11169 14976 11203
rect 14924 11160 14976 11169
rect 15108 11203 15160 11212
rect 15108 11169 15117 11203
rect 15117 11169 15151 11203
rect 15151 11169 15160 11203
rect 15108 11160 15160 11169
rect 3056 11092 3108 11144
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 6368 11092 6420 11144
rect 15384 11067 15436 11076
rect 15384 11033 15393 11067
rect 15393 11033 15427 11067
rect 15427 11033 15436 11067
rect 15384 11024 15436 11033
rect 2964 10956 3016 11008
rect 3148 10956 3200 11008
rect 1904 10854 1956 10906
rect 1968 10854 2020 10906
rect 2032 10854 2084 10906
rect 2096 10854 2148 10906
rect 2160 10854 2212 10906
rect 5837 10854 5889 10906
rect 5901 10854 5953 10906
rect 5965 10854 6017 10906
rect 6029 10854 6081 10906
rect 6093 10854 6145 10906
rect 9770 10854 9822 10906
rect 9834 10854 9886 10906
rect 9898 10854 9950 10906
rect 9962 10854 10014 10906
rect 10026 10854 10078 10906
rect 13703 10854 13755 10906
rect 13767 10854 13819 10906
rect 13831 10854 13883 10906
rect 13895 10854 13947 10906
rect 13959 10854 14011 10906
rect 848 10752 900 10804
rect 4068 10752 4120 10804
rect 5816 10684 5868 10736
rect 6460 10684 6512 10736
rect 1124 10548 1176 10600
rect 5540 10616 5592 10668
rect 6368 10616 6420 10668
rect 1768 10591 1820 10600
rect 1768 10557 1777 10591
rect 1777 10557 1811 10591
rect 1811 10557 1820 10591
rect 1768 10548 1820 10557
rect 2596 10548 2648 10600
rect 6092 10591 6144 10600
rect 6092 10557 6101 10591
rect 6101 10557 6135 10591
rect 6135 10557 6144 10591
rect 6092 10548 6144 10557
rect 6184 10548 6236 10600
rect 6000 10480 6052 10532
rect 6460 10591 6512 10600
rect 6460 10557 6469 10591
rect 6469 10557 6503 10591
rect 6503 10557 6512 10591
rect 6460 10548 6512 10557
rect 6828 10548 6880 10600
rect 9864 10591 9916 10600
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 15108 10795 15160 10804
rect 15108 10761 15117 10795
rect 15117 10761 15151 10795
rect 15151 10761 15160 10795
rect 15108 10752 15160 10761
rect 12348 10591 12400 10600
rect 12348 10557 12357 10591
rect 12357 10557 12391 10591
rect 12391 10557 12400 10591
rect 12348 10548 12400 10557
rect 15568 10548 15620 10600
rect 480 10455 532 10464
rect 480 10421 489 10455
rect 489 10421 523 10455
rect 523 10421 532 10455
rect 480 10412 532 10421
rect 5632 10412 5684 10464
rect 9496 10480 9548 10532
rect 9220 10412 9272 10464
rect 11060 10412 11112 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 2564 10310 2616 10362
rect 2628 10310 2680 10362
rect 2692 10310 2744 10362
rect 2756 10310 2808 10362
rect 2820 10310 2872 10362
rect 6497 10310 6549 10362
rect 6561 10310 6613 10362
rect 6625 10310 6677 10362
rect 6689 10310 6741 10362
rect 6753 10310 6805 10362
rect 10430 10310 10482 10362
rect 10494 10310 10546 10362
rect 10558 10310 10610 10362
rect 10622 10310 10674 10362
rect 10686 10310 10738 10362
rect 14363 10310 14415 10362
rect 14427 10310 14479 10362
rect 14491 10310 14543 10362
rect 14555 10310 14607 10362
rect 14619 10310 14671 10362
rect 1492 10208 1544 10260
rect 2780 10140 2832 10192
rect 664 10047 716 10056
rect 664 10013 673 10047
rect 673 10013 707 10047
rect 707 10013 716 10047
rect 664 10004 716 10013
rect 1676 10004 1728 10056
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 4160 10072 4212 10124
rect 5816 10208 5868 10260
rect 5908 10208 5960 10260
rect 6092 10183 6144 10192
rect 6092 10149 6101 10183
rect 6101 10149 6135 10183
rect 6135 10149 6144 10183
rect 6092 10140 6144 10149
rect 7748 10140 7800 10192
rect 9220 10208 9272 10260
rect 9864 10208 9916 10260
rect 3056 10004 3108 10056
rect 3148 10004 3200 10056
rect 5172 10115 5224 10124
rect 5172 10081 5181 10115
rect 5181 10081 5215 10115
rect 5215 10081 5224 10115
rect 5172 10072 5224 10081
rect 5448 10072 5500 10124
rect 5908 10115 5960 10124
rect 5908 10081 5917 10115
rect 5917 10081 5951 10115
rect 5951 10081 5960 10115
rect 5908 10072 5960 10081
rect 756 9868 808 9920
rect 5724 9936 5776 9988
rect 6184 10072 6236 10124
rect 6368 10072 6420 10124
rect 2688 9911 2740 9920
rect 2688 9877 2697 9911
rect 2697 9877 2731 9911
rect 2731 9877 2740 9911
rect 2688 9868 2740 9877
rect 4528 9911 4580 9920
rect 4528 9877 4537 9911
rect 4537 9877 4571 9911
rect 4571 9877 4580 9911
rect 4528 9868 4580 9877
rect 4712 9868 4764 9920
rect 5540 9868 5592 9920
rect 6184 9936 6236 9988
rect 15108 10115 15160 10124
rect 15108 10081 15117 10115
rect 15117 10081 15151 10115
rect 15151 10081 15160 10115
rect 15108 10072 15160 10081
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15384 9868 15436 9877
rect 1904 9766 1956 9818
rect 1968 9766 2020 9818
rect 2032 9766 2084 9818
rect 2096 9766 2148 9818
rect 2160 9766 2212 9818
rect 5837 9766 5889 9818
rect 5901 9766 5953 9818
rect 5965 9766 6017 9818
rect 6029 9766 6081 9818
rect 6093 9766 6145 9818
rect 9770 9766 9822 9818
rect 9834 9766 9886 9818
rect 9898 9766 9950 9818
rect 9962 9766 10014 9818
rect 10026 9766 10078 9818
rect 13703 9766 13755 9818
rect 13767 9766 13819 9818
rect 13831 9766 13883 9818
rect 13895 9766 13947 9818
rect 13959 9766 14011 9818
rect 664 9664 716 9716
rect 2688 9664 2740 9716
rect 4068 9664 4120 9716
rect 5172 9664 5224 9716
rect 1032 9460 1084 9512
rect 1768 9528 1820 9580
rect 1676 9392 1728 9444
rect 2504 9392 2556 9444
rect 3056 9528 3108 9580
rect 3424 9528 3476 9580
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 5172 9528 5224 9580
rect 2964 9503 3016 9512
rect 2964 9469 2973 9503
rect 2973 9469 3007 9503
rect 3007 9469 3016 9503
rect 2964 9460 3016 9469
rect 3148 9435 3200 9444
rect 3148 9401 3157 9435
rect 3157 9401 3191 9435
rect 3191 9401 3200 9435
rect 3148 9392 3200 9401
rect 480 9367 532 9376
rect 480 9333 489 9367
rect 489 9333 523 9367
rect 523 9333 532 9367
rect 480 9324 532 9333
rect 2780 9367 2832 9376
rect 2780 9333 2789 9367
rect 2789 9333 2823 9367
rect 2823 9333 2832 9367
rect 2780 9324 2832 9333
rect 2964 9324 3016 9376
rect 7748 9664 7800 9716
rect 15016 9639 15068 9648
rect 15016 9605 15025 9639
rect 15025 9605 15059 9639
rect 15059 9605 15068 9639
rect 15016 9596 15068 9605
rect 11704 9528 11756 9580
rect 13452 9528 13504 9580
rect 3424 9324 3476 9376
rect 4528 9324 4580 9376
rect 5356 9324 5408 9376
rect 10692 9460 10744 9512
rect 8484 9435 8536 9444
rect 8484 9401 8493 9435
rect 8493 9401 8527 9435
rect 8527 9401 8536 9435
rect 8484 9392 8536 9401
rect 9772 9392 9824 9444
rect 10140 9324 10192 9376
rect 10876 9324 10928 9376
rect 13084 9392 13136 9444
rect 14832 9392 14884 9444
rect 11888 9324 11940 9376
rect 14740 9324 14792 9376
rect 2564 9222 2616 9274
rect 2628 9222 2680 9274
rect 2692 9222 2744 9274
rect 2756 9222 2808 9274
rect 2820 9222 2872 9274
rect 6497 9222 6549 9274
rect 6561 9222 6613 9274
rect 6625 9222 6677 9274
rect 6689 9222 6741 9274
rect 6753 9222 6805 9274
rect 10430 9222 10482 9274
rect 10494 9222 10546 9274
rect 10558 9222 10610 9274
rect 10622 9222 10674 9274
rect 10686 9222 10738 9274
rect 14363 9222 14415 9274
rect 14427 9222 14479 9274
rect 14491 9222 14543 9274
rect 14555 9222 14607 9274
rect 14619 9222 14671 9274
rect 1768 9120 1820 9172
rect 2688 9120 2740 9172
rect 3240 9120 3292 9172
rect 1492 9052 1544 9104
rect 5448 9163 5500 9172
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 6828 9120 6880 9172
rect 8484 9120 8536 9172
rect 9496 9163 9548 9172
rect 9496 9129 9505 9163
rect 9505 9129 9539 9163
rect 9539 9129 9548 9163
rect 9496 9120 9548 9129
rect 9772 9120 9824 9172
rect 10784 9120 10836 9172
rect 756 9027 808 9036
rect 756 8993 765 9027
rect 765 8993 799 9027
rect 799 8993 808 9027
rect 756 8984 808 8993
rect 1032 8959 1084 8968
rect 1032 8925 1041 8959
rect 1041 8925 1075 8959
rect 1075 8925 1084 8959
rect 1032 8916 1084 8925
rect 756 8780 808 8832
rect 4528 9052 4580 9104
rect 2688 8916 2740 8968
rect 5448 8916 5500 8968
rect 6828 8984 6880 9036
rect 8852 9027 8904 9036
rect 8852 8993 8861 9027
rect 8861 8993 8895 9027
rect 8895 8993 8904 9027
rect 8852 8984 8904 8993
rect 9588 9027 9640 9036
rect 9588 8993 9597 9027
rect 9597 8993 9631 9027
rect 9631 8993 9640 9027
rect 9588 8984 9640 8993
rect 5724 8848 5776 8900
rect 11428 9027 11480 9036
rect 11428 8993 11437 9027
rect 11437 8993 11471 9027
rect 11471 8993 11480 9027
rect 11428 8984 11480 8993
rect 11888 9052 11940 9104
rect 11704 8984 11756 9036
rect 13084 9052 13136 9104
rect 14832 9120 14884 9172
rect 15016 9120 15068 9172
rect 14740 9052 14792 9104
rect 2596 8823 2648 8832
rect 2596 8789 2605 8823
rect 2605 8789 2639 8823
rect 2639 8789 2648 8823
rect 2596 8780 2648 8789
rect 2688 8780 2740 8832
rect 4068 8780 4120 8832
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 14740 8916 14792 8968
rect 13360 8780 13412 8832
rect 13544 8780 13596 8832
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 14188 8823 14240 8832
rect 14188 8789 14197 8823
rect 14197 8789 14231 8823
rect 14231 8789 14240 8823
rect 14188 8780 14240 8789
rect 15384 8823 15436 8832
rect 15384 8789 15393 8823
rect 15393 8789 15427 8823
rect 15427 8789 15436 8823
rect 15384 8780 15436 8789
rect 1904 8678 1956 8730
rect 1968 8678 2020 8730
rect 2032 8678 2084 8730
rect 2096 8678 2148 8730
rect 2160 8678 2212 8730
rect 5837 8678 5889 8730
rect 5901 8678 5953 8730
rect 5965 8678 6017 8730
rect 6029 8678 6081 8730
rect 6093 8678 6145 8730
rect 9770 8678 9822 8730
rect 9834 8678 9886 8730
rect 9898 8678 9950 8730
rect 9962 8678 10014 8730
rect 10026 8678 10078 8730
rect 13703 8678 13755 8730
rect 13767 8678 13819 8730
rect 13831 8678 13883 8730
rect 13895 8678 13947 8730
rect 13959 8678 14011 8730
rect 1032 8576 1084 8628
rect 2596 8576 2648 8628
rect 2964 8576 3016 8628
rect 3240 8576 3292 8628
rect 4068 8576 4120 8628
rect 11520 8576 11572 8628
rect 12348 8576 12400 8628
rect 13452 8576 13504 8628
rect 13544 8576 13596 8628
rect 15016 8576 15068 8628
rect 756 8415 808 8424
rect 756 8381 765 8415
rect 765 8381 799 8415
rect 799 8381 808 8415
rect 756 8372 808 8381
rect 1124 8415 1176 8424
rect 1124 8381 1133 8415
rect 1133 8381 1167 8415
rect 1167 8381 1176 8415
rect 1124 8372 1176 8381
rect 2688 8372 2740 8424
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 5724 8440 5776 8449
rect 3424 8372 3476 8424
rect 3608 8415 3660 8424
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 5356 8372 5408 8424
rect 6184 8440 6236 8492
rect 388 8347 440 8356
rect 388 8313 397 8347
rect 397 8313 431 8347
rect 431 8313 440 8347
rect 388 8304 440 8313
rect 2044 8347 2096 8356
rect 2044 8313 2053 8347
rect 2053 8313 2087 8347
rect 2087 8313 2096 8347
rect 2044 8304 2096 8313
rect 2320 8304 2372 8356
rect 2688 8236 2740 8288
rect 5448 8304 5500 8356
rect 9404 8440 9456 8492
rect 6828 8372 6880 8424
rect 7840 8372 7892 8424
rect 8484 8415 8536 8424
rect 8484 8381 8493 8415
rect 8493 8381 8527 8415
rect 8527 8381 8536 8415
rect 8484 8372 8536 8381
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 4804 8236 4856 8288
rect 6828 8279 6880 8288
rect 6828 8245 6837 8279
rect 6837 8245 6871 8279
rect 6871 8245 6880 8279
rect 6828 8236 6880 8245
rect 8024 8279 8076 8288
rect 8024 8245 8033 8279
rect 8033 8245 8067 8279
rect 8067 8245 8076 8279
rect 8024 8236 8076 8245
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 13360 8415 13412 8424
rect 13360 8381 13369 8415
rect 13369 8381 13403 8415
rect 13403 8381 13412 8415
rect 13360 8372 13412 8381
rect 14832 8508 14884 8560
rect 10968 8304 11020 8356
rect 15016 8304 15068 8356
rect 13268 8236 13320 8288
rect 13544 8236 13596 8288
rect 2564 8134 2616 8186
rect 2628 8134 2680 8186
rect 2692 8134 2744 8186
rect 2756 8134 2808 8186
rect 2820 8134 2872 8186
rect 6497 8134 6549 8186
rect 6561 8134 6613 8186
rect 6625 8134 6677 8186
rect 6689 8134 6741 8186
rect 6753 8134 6805 8186
rect 10430 8134 10482 8186
rect 10494 8134 10546 8186
rect 10558 8134 10610 8186
rect 10622 8134 10674 8186
rect 10686 8134 10738 8186
rect 14363 8134 14415 8186
rect 14427 8134 14479 8186
rect 14491 8134 14543 8186
rect 14555 8134 14607 8186
rect 14619 8134 14671 8186
rect 2320 8032 2372 8084
rect 3056 8075 3108 8084
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 6368 8032 6420 8084
rect 2044 7964 2096 8016
rect 1124 7828 1176 7880
rect 1492 7896 1544 7948
rect 1584 7828 1636 7880
rect 2228 7896 2280 7948
rect 3424 7964 3476 8016
rect 2964 7896 3016 7948
rect 4436 7896 4488 7948
rect 4804 7939 4856 7948
rect 4804 7905 4813 7939
rect 4813 7905 4847 7939
rect 4847 7905 4856 7939
rect 4804 7896 4856 7905
rect 5632 7896 5684 7948
rect 8024 8032 8076 8084
rect 8484 8032 8536 8084
rect 9404 8075 9456 8084
rect 9404 8041 9413 8075
rect 9413 8041 9447 8075
rect 9447 8041 9456 8075
rect 9404 8032 9456 8041
rect 8668 7939 8720 7948
rect 8668 7905 8677 7939
rect 8677 7905 8711 7939
rect 8711 7905 8720 7939
rect 8668 7896 8720 7905
rect 10140 8032 10192 8084
rect 15016 8032 15068 8084
rect 9680 7896 9732 7948
rect 13084 7964 13136 8016
rect 10324 7896 10376 7948
rect 1768 7760 1820 7812
rect 6828 7760 6880 7812
rect 480 7735 532 7744
rect 480 7701 489 7735
rect 489 7701 523 7735
rect 523 7701 532 7735
rect 480 7692 532 7701
rect 756 7735 808 7744
rect 756 7701 765 7735
rect 765 7701 799 7735
rect 799 7701 808 7735
rect 756 7692 808 7701
rect 2688 7735 2740 7744
rect 2688 7701 2697 7735
rect 2697 7701 2731 7735
rect 2731 7701 2740 7735
rect 2688 7692 2740 7701
rect 3240 7692 3292 7744
rect 4988 7692 5040 7744
rect 5080 7692 5132 7744
rect 8944 7828 8996 7880
rect 11704 7896 11756 7948
rect 14188 7896 14240 7948
rect 15384 7939 15436 7948
rect 15384 7905 15393 7939
rect 15393 7905 15427 7939
rect 15427 7905 15436 7939
rect 15384 7896 15436 7905
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 14740 7871 14792 7880
rect 14740 7837 14749 7871
rect 14749 7837 14783 7871
rect 14783 7837 14792 7871
rect 14740 7828 14792 7837
rect 9864 7803 9916 7812
rect 9864 7769 9873 7803
rect 9873 7769 9907 7803
rect 9907 7769 9916 7803
rect 9864 7760 9916 7769
rect 11152 7760 11204 7812
rect 7840 7692 7892 7744
rect 10140 7692 10192 7744
rect 13360 7692 13412 7744
rect 13452 7692 13504 7744
rect 13544 7692 13596 7744
rect 1904 7590 1956 7642
rect 1968 7590 2020 7642
rect 2032 7590 2084 7642
rect 2096 7590 2148 7642
rect 2160 7590 2212 7642
rect 5837 7590 5889 7642
rect 5901 7590 5953 7642
rect 5965 7590 6017 7642
rect 6029 7590 6081 7642
rect 6093 7590 6145 7642
rect 9770 7590 9822 7642
rect 9834 7590 9886 7642
rect 9898 7590 9950 7642
rect 9962 7590 10014 7642
rect 10026 7590 10078 7642
rect 13703 7590 13755 7642
rect 13767 7590 13819 7642
rect 13831 7590 13883 7642
rect 13895 7590 13947 7642
rect 13959 7590 14011 7642
rect 2320 7488 2372 7540
rect 2688 7488 2740 7540
rect 5356 7488 5408 7540
rect 5724 7488 5776 7540
rect 12256 7488 12308 7540
rect 13544 7488 13596 7540
rect 14188 7488 14240 7540
rect 14740 7488 14792 7540
rect 5540 7420 5592 7472
rect 756 7352 808 7404
rect 3608 7352 3660 7404
rect 4528 7352 4580 7404
rect 11704 7352 11756 7404
rect 388 7327 440 7336
rect 388 7293 397 7327
rect 397 7293 431 7327
rect 431 7293 440 7327
rect 388 7284 440 7293
rect 1492 7148 1544 7200
rect 4988 7327 5040 7336
rect 4988 7293 4997 7327
rect 4997 7293 5031 7327
rect 5031 7293 5040 7327
rect 4988 7284 5040 7293
rect 5080 7284 5132 7336
rect 5448 7327 5500 7336
rect 5448 7293 5457 7327
rect 5457 7293 5491 7327
rect 5491 7293 5500 7327
rect 5448 7284 5500 7293
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 7748 7284 7800 7336
rect 13912 7420 13964 7472
rect 13544 7395 13596 7404
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 13360 7327 13412 7336
rect 13360 7293 13369 7327
rect 13369 7293 13403 7327
rect 13403 7293 13412 7327
rect 13360 7284 13412 7293
rect 13452 7284 13504 7336
rect 4344 7216 4396 7268
rect 6276 7259 6328 7268
rect 6276 7225 6285 7259
rect 6285 7225 6319 7259
rect 6319 7225 6328 7259
rect 6276 7216 6328 7225
rect 7932 7259 7984 7268
rect 7932 7225 7941 7259
rect 7941 7225 7975 7259
rect 7975 7225 7984 7259
rect 7932 7216 7984 7225
rect 10784 7216 10836 7268
rect 11520 7216 11572 7268
rect 14004 7284 14056 7336
rect 15016 7284 15068 7336
rect 2228 7148 2280 7200
rect 2964 7148 3016 7200
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 8208 7148 8260 7200
rect 9864 7148 9916 7200
rect 2564 7046 2616 7098
rect 2628 7046 2680 7098
rect 2692 7046 2744 7098
rect 2756 7046 2808 7098
rect 2820 7046 2872 7098
rect 6497 7046 6549 7098
rect 6561 7046 6613 7098
rect 6625 7046 6677 7098
rect 6689 7046 6741 7098
rect 6753 7046 6805 7098
rect 10430 7046 10482 7098
rect 10494 7046 10546 7098
rect 10558 7046 10610 7098
rect 10622 7046 10674 7098
rect 10686 7046 10738 7098
rect 14363 7046 14415 7098
rect 14427 7046 14479 7098
rect 14491 7046 14543 7098
rect 14555 7046 14607 7098
rect 14619 7046 14671 7098
rect 1492 6944 1544 6996
rect 4344 6944 4396 6996
rect 6276 6944 6328 6996
rect 9220 6944 9272 6996
rect 10324 6944 10376 6996
rect 14004 6944 14056 6996
rect 15016 6944 15068 6996
rect 8944 6876 8996 6928
rect 1308 6808 1360 6860
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 4160 6851 4212 6860
rect 4160 6817 4169 6851
rect 4169 6817 4203 6851
rect 4203 6817 4212 6851
rect 4160 6808 4212 6817
rect 7748 6808 7800 6860
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 8484 6808 8536 6860
rect 4252 6740 4304 6792
rect 5448 6740 5500 6792
rect 9864 6740 9916 6792
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 11152 6851 11204 6860
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 11152 6808 11204 6817
rect 11428 6808 11480 6860
rect 13268 6808 13320 6860
rect 13544 6808 13596 6860
rect 13912 6808 13964 6860
rect 14096 6808 14148 6860
rect 15292 6851 15344 6860
rect 15292 6817 15301 6851
rect 15301 6817 15335 6851
rect 15335 6817 15344 6851
rect 15292 6808 15344 6817
rect 10140 6740 10192 6792
rect 9128 6672 9180 6724
rect 11336 6672 11388 6724
rect 480 6647 532 6656
rect 480 6613 489 6647
rect 489 6613 523 6647
rect 523 6613 532 6647
rect 480 6604 532 6613
rect 1400 6604 1452 6656
rect 3148 6604 3200 6656
rect 4344 6647 4396 6656
rect 4344 6613 4353 6647
rect 4353 6613 4387 6647
rect 4387 6613 4396 6647
rect 4344 6604 4396 6613
rect 8024 6604 8076 6656
rect 8852 6604 8904 6656
rect 9496 6604 9548 6656
rect 14648 6604 14700 6656
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 1904 6502 1956 6554
rect 1968 6502 2020 6554
rect 2032 6502 2084 6554
rect 2096 6502 2148 6554
rect 2160 6502 2212 6554
rect 5837 6502 5889 6554
rect 5901 6502 5953 6554
rect 5965 6502 6017 6554
rect 6029 6502 6081 6554
rect 6093 6502 6145 6554
rect 9770 6502 9822 6554
rect 9834 6502 9886 6554
rect 9898 6502 9950 6554
rect 9962 6502 10014 6554
rect 10026 6502 10078 6554
rect 13703 6502 13755 6554
rect 13767 6502 13819 6554
rect 13831 6502 13883 6554
rect 13895 6502 13947 6554
rect 13959 6502 14011 6554
rect 1676 6400 1728 6452
rect 388 6307 440 6316
rect 388 6273 397 6307
rect 397 6273 431 6307
rect 431 6273 440 6307
rect 388 6264 440 6273
rect 1308 6264 1360 6316
rect 1768 6196 1820 6248
rect 664 6171 716 6180
rect 664 6137 673 6171
rect 673 6137 707 6171
rect 707 6137 716 6171
rect 664 6128 716 6137
rect 2964 6400 3016 6452
rect 4160 6400 4212 6452
rect 4344 6400 4396 6452
rect 6184 6400 6236 6452
rect 8668 6400 8720 6452
rect 5540 6332 5592 6384
rect 9496 6400 9548 6452
rect 10968 6400 11020 6452
rect 12716 6443 12768 6452
rect 12716 6409 12725 6443
rect 12725 6409 12759 6443
rect 12759 6409 12768 6443
rect 12716 6400 12768 6409
rect 15292 6400 15344 6452
rect 4528 6264 4580 6316
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 5724 6264 5776 6316
rect 8484 6264 8536 6316
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 10140 6264 10192 6316
rect 11244 6264 11296 6316
rect 11704 6264 11756 6316
rect 11980 6264 12032 6316
rect 13544 6264 13596 6316
rect 14648 6375 14700 6384
rect 14648 6341 14657 6375
rect 14657 6341 14691 6375
rect 14691 6341 14700 6375
rect 14648 6332 14700 6341
rect 6092 6239 6144 6248
rect 6092 6205 6101 6239
rect 6101 6205 6135 6239
rect 6135 6205 6144 6239
rect 6092 6196 6144 6205
rect 6828 6196 6880 6248
rect 9220 6239 9272 6248
rect 9220 6205 9229 6239
rect 9229 6205 9263 6239
rect 9263 6205 9272 6239
rect 9220 6196 9272 6205
rect 9404 6239 9456 6248
rect 9404 6205 9413 6239
rect 9413 6205 9447 6239
rect 9447 6205 9456 6239
rect 9404 6196 9456 6205
rect 2320 6128 2372 6180
rect 3700 6171 3752 6180
rect 3700 6137 3709 6171
rect 3709 6137 3743 6171
rect 3743 6137 3752 6171
rect 3700 6128 3752 6137
rect 4160 6128 4212 6180
rect 6184 6128 6236 6180
rect 8944 6128 8996 6180
rect 12716 6196 12768 6248
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 5172 6060 5224 6112
rect 7288 6060 7340 6112
rect 10784 6128 10836 6180
rect 12532 6128 12584 6180
rect 11428 6060 11480 6112
rect 11980 6060 12032 6112
rect 13728 6103 13780 6112
rect 13728 6069 13737 6103
rect 13737 6069 13771 6103
rect 13771 6069 13780 6103
rect 13728 6060 13780 6069
rect 2564 5958 2616 6010
rect 2628 5958 2680 6010
rect 2692 5958 2744 6010
rect 2756 5958 2808 6010
rect 2820 5958 2872 6010
rect 6497 5958 6549 6010
rect 6561 5958 6613 6010
rect 6625 5958 6677 6010
rect 6689 5958 6741 6010
rect 6753 5958 6805 6010
rect 10430 5958 10482 6010
rect 10494 5958 10546 6010
rect 10558 5958 10610 6010
rect 10622 5958 10674 6010
rect 10686 5958 10738 6010
rect 14363 5958 14415 6010
rect 14427 5958 14479 6010
rect 14491 5958 14543 6010
rect 14555 5958 14607 6010
rect 14619 5958 14671 6010
rect 664 5856 716 5908
rect 1032 5763 1084 5772
rect 1032 5729 1041 5763
rect 1041 5729 1075 5763
rect 1075 5729 1084 5763
rect 1032 5720 1084 5729
rect 2320 5856 2372 5908
rect 1308 5788 1360 5840
rect 1584 5720 1636 5772
rect 3148 5652 3200 5704
rect 1676 5584 1728 5636
rect 4528 5856 4580 5908
rect 5724 5856 5776 5908
rect 6092 5856 6144 5908
rect 8668 5856 8720 5908
rect 9404 5856 9456 5908
rect 11152 5856 11204 5908
rect 4436 5788 4488 5840
rect 8208 5831 8260 5840
rect 8208 5797 8217 5831
rect 8217 5797 8251 5831
rect 8251 5797 8260 5831
rect 8208 5788 8260 5797
rect 11244 5788 11296 5840
rect 4160 5720 4212 5772
rect 4712 5720 4764 5772
rect 5080 5652 5132 5704
rect 6184 5720 6236 5772
rect 7196 5720 7248 5772
rect 7656 5763 7708 5772
rect 7656 5729 7665 5763
rect 7665 5729 7699 5763
rect 7699 5729 7708 5763
rect 7656 5720 7708 5729
rect 8116 5720 8168 5772
rect 9680 5720 9732 5772
rect 3884 5584 3936 5636
rect 8852 5652 8904 5704
rect 10784 5720 10836 5772
rect 10876 5763 10928 5772
rect 10876 5729 10885 5763
rect 10885 5729 10919 5763
rect 10919 5729 10928 5763
rect 10876 5720 10928 5729
rect 10968 5763 11020 5772
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 11336 5763 11388 5772
rect 11336 5729 11345 5763
rect 11345 5729 11379 5763
rect 11379 5729 11388 5763
rect 11336 5720 11388 5729
rect 14832 5899 14884 5908
rect 14832 5865 14841 5899
rect 14841 5865 14875 5899
rect 14875 5865 14884 5899
rect 14832 5856 14884 5865
rect 13084 5788 13136 5840
rect 14832 5652 14884 5704
rect 388 5516 440 5568
rect 480 5559 532 5568
rect 480 5525 489 5559
rect 489 5525 523 5559
rect 523 5525 532 5559
rect 480 5516 532 5525
rect 3516 5516 3568 5568
rect 4712 5516 4764 5568
rect 4804 5559 4856 5568
rect 4804 5525 4813 5559
rect 4813 5525 4847 5559
rect 4847 5525 4856 5559
rect 4804 5516 4856 5525
rect 5448 5516 5500 5568
rect 5632 5516 5684 5568
rect 9220 5516 9272 5568
rect 9588 5516 9640 5568
rect 10324 5559 10376 5568
rect 10324 5525 10333 5559
rect 10333 5525 10367 5559
rect 10367 5525 10376 5559
rect 10324 5516 10376 5525
rect 11428 5584 11480 5636
rect 15384 5559 15436 5568
rect 15384 5525 15393 5559
rect 15393 5525 15427 5559
rect 15427 5525 15436 5559
rect 15384 5516 15436 5525
rect 1904 5414 1956 5466
rect 1968 5414 2020 5466
rect 2032 5414 2084 5466
rect 2096 5414 2148 5466
rect 2160 5414 2212 5466
rect 5837 5414 5889 5466
rect 5901 5414 5953 5466
rect 5965 5414 6017 5466
rect 6029 5414 6081 5466
rect 6093 5414 6145 5466
rect 9770 5414 9822 5466
rect 9834 5414 9886 5466
rect 9898 5414 9950 5466
rect 9962 5414 10014 5466
rect 10026 5414 10078 5466
rect 13703 5414 13755 5466
rect 13767 5414 13819 5466
rect 13831 5414 13883 5466
rect 13895 5414 13947 5466
rect 13959 5414 14011 5466
rect 3700 5312 3752 5364
rect 4068 5312 4120 5364
rect 5172 5355 5224 5364
rect 5172 5321 5181 5355
rect 5181 5321 5215 5355
rect 5215 5321 5224 5355
rect 5172 5312 5224 5321
rect 5356 5312 5408 5364
rect 7288 5312 7340 5364
rect 4712 5244 4764 5296
rect 3976 5176 4028 5228
rect 4160 5176 4212 5228
rect 8300 5244 8352 5296
rect 8760 5244 8812 5296
rect 3516 5151 3568 5160
rect 3516 5117 3525 5151
rect 3525 5117 3559 5151
rect 3559 5117 3568 5151
rect 3516 5108 3568 5117
rect 3792 5108 3844 5160
rect 3884 5108 3936 5160
rect 4528 5151 4580 5160
rect 4528 5117 4537 5151
rect 4537 5117 4571 5151
rect 4571 5117 4580 5151
rect 4528 5108 4580 5117
rect 4712 5151 4764 5160
rect 4712 5117 4721 5151
rect 4721 5117 4755 5151
rect 4755 5117 4764 5151
rect 4712 5108 4764 5117
rect 5172 5108 5224 5160
rect 5632 5151 5684 5160
rect 5632 5117 5641 5151
rect 5641 5117 5675 5151
rect 5675 5117 5684 5151
rect 5632 5108 5684 5117
rect 5724 5151 5776 5160
rect 5724 5117 5733 5151
rect 5733 5117 5767 5151
rect 5767 5117 5776 5151
rect 5724 5108 5776 5117
rect 5908 5108 5960 5160
rect 6184 5108 6236 5160
rect 4252 5040 4304 5092
rect 5540 5040 5592 5092
rect 2964 4972 3016 5024
rect 3700 4972 3752 5024
rect 5632 4972 5684 5024
rect 6276 5040 6328 5092
rect 7012 5108 7064 5160
rect 7196 5108 7248 5160
rect 7288 5151 7340 5160
rect 7288 5117 7321 5151
rect 7321 5117 7340 5151
rect 7288 5108 7340 5117
rect 7656 5108 7708 5160
rect 8300 5151 8352 5160
rect 8300 5117 8309 5151
rect 8309 5117 8343 5151
rect 8343 5117 8352 5151
rect 8300 5108 8352 5117
rect 8668 5151 8720 5160
rect 8668 5117 8677 5151
rect 8677 5117 8711 5151
rect 8711 5117 8720 5151
rect 8668 5108 8720 5117
rect 8760 5151 8812 5160
rect 8760 5117 8774 5151
rect 8774 5117 8808 5151
rect 8808 5117 8812 5151
rect 8760 5108 8812 5117
rect 10968 5312 11020 5364
rect 12532 5312 12584 5364
rect 9680 5244 9732 5296
rect 9588 5151 9640 5160
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 9956 5176 10008 5228
rect 13084 5244 13136 5296
rect 10784 5176 10836 5228
rect 11060 5108 11112 5160
rect 13912 5176 13964 5228
rect 12716 5151 12768 5160
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 12716 5108 12768 5117
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 6000 5015 6052 5024
rect 6000 4981 6009 5015
rect 6009 4981 6043 5015
rect 6043 4981 6052 5015
rect 6000 4972 6052 4981
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 7840 4972 7892 5024
rect 8300 4972 8352 5024
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 8944 4972 8996 4981
rect 10140 4972 10192 5024
rect 10968 5015 11020 5024
rect 10968 4981 10977 5015
rect 10977 4981 11011 5015
rect 11011 4981 11020 5015
rect 10968 4972 11020 4981
rect 14004 4972 14056 5024
rect 14740 4972 14792 5024
rect 15200 4972 15252 5024
rect 2564 4870 2616 4922
rect 2628 4870 2680 4922
rect 2692 4870 2744 4922
rect 2756 4870 2808 4922
rect 2820 4870 2872 4922
rect 6497 4870 6549 4922
rect 6561 4870 6613 4922
rect 6625 4870 6677 4922
rect 6689 4870 6741 4922
rect 6753 4870 6805 4922
rect 10430 4870 10482 4922
rect 10494 4870 10546 4922
rect 10558 4870 10610 4922
rect 10622 4870 10674 4922
rect 10686 4870 10738 4922
rect 14363 4870 14415 4922
rect 14427 4870 14479 4922
rect 14491 4870 14543 4922
rect 14555 4870 14607 4922
rect 14619 4870 14671 4922
rect 388 4675 440 4684
rect 388 4641 397 4675
rect 397 4641 431 4675
rect 431 4641 440 4675
rect 388 4632 440 4641
rect 1768 4632 1820 4684
rect 2320 4632 2372 4684
rect 2964 4632 3016 4684
rect 7012 4768 7064 4820
rect 7380 4768 7432 4820
rect 7472 4811 7524 4820
rect 7472 4777 7481 4811
rect 7481 4777 7515 4811
rect 7515 4777 7524 4811
rect 7472 4768 7524 4777
rect 8852 4768 8904 4820
rect 11060 4768 11112 4820
rect 12716 4768 12768 4820
rect 14004 4811 14056 4820
rect 4804 4700 4856 4752
rect 5356 4700 5408 4752
rect 3516 4632 3568 4684
rect 3700 4675 3752 4684
rect 3700 4641 3709 4675
rect 3709 4641 3743 4675
rect 3743 4641 3752 4675
rect 3700 4632 3752 4641
rect 664 4607 716 4616
rect 664 4573 673 4607
rect 673 4573 707 4607
rect 707 4573 716 4607
rect 664 4564 716 4573
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 5448 4632 5500 4641
rect 5632 4675 5684 4684
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5632 4632 5684 4641
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 6000 4632 6052 4684
rect 6184 4632 6236 4684
rect 6828 4632 6880 4684
rect 4712 4564 4764 4616
rect 5264 4564 5316 4616
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 8944 4700 8996 4752
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 10232 4743 10284 4752
rect 10232 4709 10241 4743
rect 10241 4709 10275 4743
rect 10275 4709 10284 4743
rect 14004 4777 14013 4811
rect 14013 4777 14047 4811
rect 14047 4777 14056 4811
rect 14004 4768 14056 4777
rect 14832 4811 14884 4820
rect 14832 4777 14841 4811
rect 14841 4777 14875 4811
rect 14875 4777 14884 4811
rect 14832 4768 14884 4777
rect 10232 4700 10284 4709
rect 7104 4564 7156 4616
rect 7564 4564 7616 4616
rect 9588 4632 9640 4684
rect 12440 4632 12492 4684
rect 2412 4496 2464 4548
rect 1124 4428 1176 4480
rect 3332 4471 3384 4480
rect 3332 4437 3341 4471
rect 3341 4437 3375 4471
rect 3375 4437 3384 4471
rect 3332 4428 3384 4437
rect 4528 4471 4580 4480
rect 4528 4437 4537 4471
rect 4537 4437 4571 4471
rect 4571 4437 4580 4471
rect 4528 4428 4580 4437
rect 4620 4428 4672 4480
rect 5172 4496 5224 4548
rect 5724 4428 5776 4480
rect 6552 4428 6604 4480
rect 6644 4428 6696 4480
rect 7564 4428 7616 4480
rect 8116 4496 8168 4548
rect 8484 4496 8536 4548
rect 9956 4496 10008 4548
rect 8300 4428 8352 4480
rect 8392 4471 8444 4480
rect 8392 4437 8401 4471
rect 8401 4437 8435 4471
rect 8435 4437 8444 4471
rect 8392 4428 8444 4437
rect 9680 4428 9732 4480
rect 11428 4564 11480 4616
rect 13268 4632 13320 4684
rect 14740 4700 14792 4752
rect 13912 4632 13964 4684
rect 14464 4632 14516 4684
rect 14648 4675 14700 4684
rect 14648 4641 14657 4675
rect 14657 4641 14691 4675
rect 14691 4641 14700 4675
rect 14648 4632 14700 4641
rect 15384 4675 15436 4684
rect 15384 4641 15393 4675
rect 15393 4641 15427 4675
rect 15427 4641 15436 4675
rect 15384 4632 15436 4641
rect 11336 4428 11388 4480
rect 12808 4471 12860 4480
rect 12808 4437 12817 4471
rect 12817 4437 12851 4471
rect 12851 4437 12860 4471
rect 12808 4428 12860 4437
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 1904 4326 1956 4378
rect 1968 4326 2020 4378
rect 2032 4326 2084 4378
rect 2096 4326 2148 4378
rect 2160 4326 2212 4378
rect 5837 4326 5889 4378
rect 5901 4326 5953 4378
rect 5965 4326 6017 4378
rect 6029 4326 6081 4378
rect 6093 4326 6145 4378
rect 9770 4326 9822 4378
rect 9834 4326 9886 4378
rect 9898 4326 9950 4378
rect 9962 4326 10014 4378
rect 10026 4326 10078 4378
rect 13703 4326 13755 4378
rect 13767 4326 13819 4378
rect 13831 4326 13883 4378
rect 13895 4326 13947 4378
rect 13959 4326 14011 4378
rect 664 4224 716 4276
rect 1032 4063 1084 4072
rect 1032 4029 1041 4063
rect 1041 4029 1075 4063
rect 1075 4029 1084 4063
rect 1032 4020 1084 4029
rect 1124 4063 1176 4072
rect 1124 4029 1133 4063
rect 1133 4029 1167 4063
rect 1167 4029 1176 4063
rect 1124 4020 1176 4029
rect 4528 4088 4580 4140
rect 3332 4020 3384 4072
rect 3700 4063 3752 4072
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 5172 4156 5224 4208
rect 6552 4156 6604 4208
rect 7472 4224 7524 4276
rect 8852 4224 8904 4276
rect 7104 4156 7156 4208
rect 8024 4156 8076 4208
rect 8484 4156 8536 4208
rect 10140 4156 10192 4208
rect 10508 4199 10560 4208
rect 10508 4165 10517 4199
rect 10517 4165 10551 4199
rect 10551 4165 10560 4199
rect 10508 4156 10560 4165
rect 11428 4224 11480 4276
rect 940 3884 992 3936
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 2228 3884 2280 3893
rect 2320 3884 2372 3936
rect 3148 3884 3200 3936
rect 4252 3884 4304 3936
rect 4436 3927 4488 3936
rect 4436 3893 4445 3927
rect 4445 3893 4479 3927
rect 4479 3893 4488 3927
rect 4436 3884 4488 3893
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 5724 4088 5776 4140
rect 4804 3884 4856 3936
rect 5540 4020 5592 4072
rect 6828 4088 6880 4140
rect 5172 3995 5224 4004
rect 5172 3961 5181 3995
rect 5181 3961 5215 3995
rect 5215 3961 5224 3995
rect 5172 3952 5224 3961
rect 6184 4063 6236 4072
rect 6184 4029 6193 4063
rect 6193 4029 6227 4063
rect 6227 4029 6236 4063
rect 6184 4020 6236 4029
rect 6276 4020 6328 4072
rect 6644 4063 6696 4072
rect 6644 4029 6653 4063
rect 6653 4029 6687 4063
rect 6687 4029 6696 4063
rect 6644 4020 6696 4029
rect 6736 4020 6788 4072
rect 5264 3927 5316 3936
rect 5264 3893 5273 3927
rect 5273 3893 5307 3927
rect 5307 3893 5316 3927
rect 5264 3884 5316 3893
rect 5448 3884 5500 3936
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 6828 3952 6880 4004
rect 8392 4088 8444 4140
rect 9312 4088 9364 4140
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 8668 4020 8720 4072
rect 10324 4063 10376 4072
rect 8944 3995 8996 4004
rect 8944 3961 8953 3995
rect 8953 3961 8987 3995
rect 8987 3961 8996 3995
rect 8944 3952 8996 3961
rect 10324 4029 10333 4063
rect 10333 4029 10367 4063
rect 10367 4029 10376 4063
rect 10324 4020 10376 4029
rect 7380 3884 7432 3936
rect 7840 3884 7892 3936
rect 10140 3995 10192 4004
rect 10140 3961 10149 3995
rect 10149 3961 10183 3995
rect 10183 3961 10192 3995
rect 10876 4020 10928 4072
rect 11060 4020 11112 4072
rect 12808 4156 12860 4208
rect 15568 4088 15620 4140
rect 10140 3952 10192 3961
rect 10784 3952 10836 4004
rect 10232 3884 10284 3936
rect 10876 3884 10928 3936
rect 13268 4020 13320 4072
rect 13544 4020 13596 4072
rect 14464 4063 14516 4072
rect 14464 4029 14473 4063
rect 14473 4029 14507 4063
rect 14507 4029 14516 4063
rect 14464 4020 14516 4029
rect 15200 4020 15252 4072
rect 15384 4063 15436 4072
rect 15384 4029 15393 4063
rect 15393 4029 15427 4063
rect 15427 4029 15436 4063
rect 15384 4020 15436 4029
rect 14740 3952 14792 4004
rect 13360 3884 13412 3936
rect 14280 3927 14332 3936
rect 14280 3893 14289 3927
rect 14289 3893 14323 3927
rect 14323 3893 14332 3927
rect 14280 3884 14332 3893
rect 15016 3952 15068 4004
rect 15108 3884 15160 3936
rect 2564 3782 2616 3834
rect 2628 3782 2680 3834
rect 2692 3782 2744 3834
rect 2756 3782 2808 3834
rect 2820 3782 2872 3834
rect 6497 3782 6549 3834
rect 6561 3782 6613 3834
rect 6625 3782 6677 3834
rect 6689 3782 6741 3834
rect 6753 3782 6805 3834
rect 10430 3782 10482 3834
rect 10494 3782 10546 3834
rect 10558 3782 10610 3834
rect 10622 3782 10674 3834
rect 10686 3782 10738 3834
rect 14363 3782 14415 3834
rect 14427 3782 14479 3834
rect 14491 3782 14543 3834
rect 14555 3782 14607 3834
rect 14619 3782 14671 3834
rect 480 3723 532 3732
rect 480 3689 489 3723
rect 489 3689 523 3723
rect 523 3689 532 3723
rect 480 3680 532 3689
rect 940 3723 992 3732
rect 940 3689 949 3723
rect 949 3689 983 3723
rect 983 3689 992 3723
rect 940 3680 992 3689
rect 5540 3680 5592 3732
rect 6920 3680 6972 3732
rect 7564 3680 7616 3732
rect 2228 3612 2280 3664
rect 3148 3612 3200 3664
rect 5264 3612 5316 3664
rect 6828 3612 6880 3664
rect 7472 3612 7524 3664
rect 1124 3587 1176 3596
rect 1124 3553 1133 3587
rect 1133 3553 1167 3587
rect 1167 3553 1176 3587
rect 1124 3544 1176 3553
rect 1676 3544 1728 3596
rect 4252 3476 4304 3528
rect 4804 3544 4856 3596
rect 7196 3587 7248 3596
rect 7196 3553 7205 3587
rect 7205 3553 7239 3587
rect 7239 3553 7248 3587
rect 7196 3544 7248 3553
rect 6828 3476 6880 3528
rect 4712 3340 4764 3392
rect 7564 3544 7616 3596
rect 10140 3680 10192 3732
rect 10324 3723 10376 3732
rect 10324 3689 10333 3723
rect 10333 3689 10367 3723
rect 10367 3689 10376 3723
rect 10324 3680 10376 3689
rect 11060 3680 11112 3732
rect 10232 3612 10284 3664
rect 10784 3612 10836 3664
rect 12532 3680 12584 3732
rect 10692 3587 10744 3596
rect 10692 3553 10701 3587
rect 10701 3553 10735 3587
rect 10735 3553 10744 3587
rect 10692 3544 10744 3553
rect 15384 3680 15436 3732
rect 7380 3408 7432 3460
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 8852 3519 8904 3528
rect 8852 3485 8861 3519
rect 8861 3485 8895 3519
rect 8895 3485 8904 3519
rect 8852 3476 8904 3485
rect 9312 3476 9364 3528
rect 10324 3476 10376 3528
rect 10876 3476 10928 3528
rect 7748 3451 7800 3460
rect 7748 3417 7757 3451
rect 7757 3417 7791 3451
rect 7791 3417 7800 3451
rect 7748 3408 7800 3417
rect 8116 3408 8168 3460
rect 7564 3383 7616 3392
rect 7564 3349 7573 3383
rect 7573 3349 7607 3383
rect 7607 3349 7616 3383
rect 7564 3340 7616 3349
rect 12716 3544 12768 3596
rect 13084 3544 13136 3596
rect 13360 3544 13412 3596
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 11336 3519 11388 3528
rect 11336 3485 11345 3519
rect 11345 3485 11379 3519
rect 11379 3485 11388 3519
rect 11336 3476 11388 3485
rect 13452 3340 13504 3392
rect 14832 3340 14884 3392
rect 1904 3238 1956 3290
rect 1968 3238 2020 3290
rect 2032 3238 2084 3290
rect 2096 3238 2148 3290
rect 2160 3238 2212 3290
rect 5837 3238 5889 3290
rect 5901 3238 5953 3290
rect 5965 3238 6017 3290
rect 6029 3238 6081 3290
rect 6093 3238 6145 3290
rect 9770 3238 9822 3290
rect 9834 3238 9886 3290
rect 9898 3238 9950 3290
rect 9962 3238 10014 3290
rect 10026 3238 10078 3290
rect 13703 3238 13755 3290
rect 13767 3238 13819 3290
rect 13831 3238 13883 3290
rect 13895 3238 13947 3290
rect 13959 3238 14011 3290
rect 3148 3136 3200 3188
rect 3516 3179 3568 3188
rect 3516 3145 3525 3179
rect 3525 3145 3559 3179
rect 3559 3145 3568 3179
rect 3516 3136 3568 3145
rect 5080 3136 5132 3188
rect 7288 3136 7340 3188
rect 8576 3136 8628 3188
rect 9588 3136 9640 3188
rect 10232 3179 10284 3188
rect 10232 3145 10241 3179
rect 10241 3145 10275 3179
rect 10275 3145 10284 3179
rect 10232 3136 10284 3145
rect 10876 3136 10928 3188
rect 13452 3136 13504 3188
rect 13544 3136 13596 3188
rect 14832 3136 14884 3188
rect 15292 3136 15344 3188
rect 15476 3136 15528 3188
rect 4068 3068 4120 3120
rect 7288 3000 7340 3052
rect 388 2975 440 2984
rect 388 2941 397 2975
rect 397 2941 431 2975
rect 431 2941 440 2975
rect 388 2932 440 2941
rect 3332 2975 3384 2984
rect 3332 2941 3341 2975
rect 3341 2941 3375 2975
rect 3375 2941 3384 2975
rect 3332 2932 3384 2941
rect 3884 2975 3936 2984
rect 3884 2941 3893 2975
rect 3893 2941 3927 2975
rect 3927 2941 3936 2975
rect 3884 2932 3936 2941
rect 5172 2932 5224 2984
rect 5264 2932 5316 2984
rect 6184 2932 6236 2984
rect 7012 2932 7064 2984
rect 4712 2864 4764 2916
rect 8852 3068 8904 3120
rect 8944 3000 8996 3052
rect 10692 3000 10744 3052
rect 8208 2975 8260 2984
rect 8208 2941 8217 2975
rect 8217 2941 8251 2975
rect 8251 2941 8260 2975
rect 8208 2932 8260 2941
rect 11152 2932 11204 2984
rect 9496 2864 9548 2916
rect 10876 2864 10928 2916
rect 13176 2864 13228 2916
rect 5632 2796 5684 2848
rect 7748 2796 7800 2848
rect 9588 2796 9640 2848
rect 11428 2796 11480 2848
rect 11612 2839 11664 2848
rect 11612 2805 11621 2839
rect 11621 2805 11655 2839
rect 11655 2805 11664 2839
rect 11612 2796 11664 2805
rect 14372 2932 14424 2984
rect 15016 2932 15068 2984
rect 2564 2694 2616 2746
rect 2628 2694 2680 2746
rect 2692 2694 2744 2746
rect 2756 2694 2808 2746
rect 2820 2694 2872 2746
rect 6497 2694 6549 2746
rect 6561 2694 6613 2746
rect 6625 2694 6677 2746
rect 6689 2694 6741 2746
rect 6753 2694 6805 2746
rect 10430 2694 10482 2746
rect 10494 2694 10546 2746
rect 10558 2694 10610 2746
rect 10622 2694 10674 2746
rect 10686 2694 10738 2746
rect 14363 2694 14415 2746
rect 14427 2694 14479 2746
rect 14491 2694 14543 2746
rect 14555 2694 14607 2746
rect 14619 2694 14671 2746
rect 3884 2635 3936 2644
rect 3884 2601 3893 2635
rect 3893 2601 3927 2635
rect 3927 2601 3936 2635
rect 3884 2592 3936 2601
rect 6828 2592 6880 2644
rect 2412 2567 2464 2576
rect 2412 2533 2421 2567
rect 2421 2533 2455 2567
rect 2455 2533 2464 2567
rect 2412 2524 2464 2533
rect 3516 2456 3568 2508
rect 7012 2456 7064 2508
rect 9588 2592 9640 2644
rect 10876 2567 10928 2576
rect 10876 2533 10885 2567
rect 10885 2533 10919 2567
rect 10919 2533 10928 2567
rect 10876 2524 10928 2533
rect 13176 2635 13228 2644
rect 13176 2601 13185 2635
rect 13185 2601 13219 2635
rect 13219 2601 13228 2635
rect 13176 2592 13228 2601
rect 10232 2456 10284 2508
rect 10324 2456 10376 2508
rect 11152 2524 11204 2576
rect 11704 2567 11756 2576
rect 11704 2533 11713 2567
rect 11713 2533 11747 2567
rect 11747 2533 11756 2567
rect 11704 2524 11756 2533
rect 14924 2524 14976 2576
rect 15200 2524 15252 2576
rect 11244 2456 11296 2508
rect 11428 2499 11480 2508
rect 11428 2465 11437 2499
rect 11437 2465 11471 2499
rect 11471 2465 11480 2499
rect 11428 2456 11480 2465
rect 12716 2456 12768 2508
rect 13452 2456 13504 2508
rect 13544 2499 13596 2508
rect 13544 2465 13553 2499
rect 13553 2465 13587 2499
rect 13587 2465 13596 2499
rect 13544 2456 13596 2465
rect 14648 2456 14700 2508
rect 1768 2388 1820 2440
rect 7564 2388 7616 2440
rect 4436 2252 4488 2304
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 14832 2252 14884 2304
rect 14924 2295 14976 2304
rect 14924 2261 14933 2295
rect 14933 2261 14967 2295
rect 14967 2261 14976 2295
rect 14924 2252 14976 2261
rect 15384 2295 15436 2304
rect 15384 2261 15393 2295
rect 15393 2261 15427 2295
rect 15427 2261 15436 2295
rect 15384 2252 15436 2261
rect 1904 2150 1956 2202
rect 1968 2150 2020 2202
rect 2032 2150 2084 2202
rect 2096 2150 2148 2202
rect 2160 2150 2212 2202
rect 5837 2150 5889 2202
rect 5901 2150 5953 2202
rect 5965 2150 6017 2202
rect 6029 2150 6081 2202
rect 6093 2150 6145 2202
rect 9770 2150 9822 2202
rect 9834 2150 9886 2202
rect 9898 2150 9950 2202
rect 9962 2150 10014 2202
rect 10026 2150 10078 2202
rect 13703 2150 13755 2202
rect 13767 2150 13819 2202
rect 13831 2150 13883 2202
rect 13895 2150 13947 2202
rect 13959 2150 14011 2202
rect 4068 2048 4120 2100
rect 7932 2048 7984 2100
rect 13544 2048 13596 2100
rect 14280 2048 14332 2100
rect 14924 2048 14976 2100
rect 15200 2091 15252 2100
rect 15200 2057 15209 2091
rect 15209 2057 15243 2091
rect 15243 2057 15252 2091
rect 15200 2048 15252 2057
rect 6184 2023 6236 2032
rect 6184 1989 6193 2023
rect 6193 1989 6227 2023
rect 6227 1989 6236 2023
rect 6184 1980 6236 1989
rect 7012 1980 7064 2032
rect 4436 1955 4488 1964
rect 4436 1921 4445 1955
rect 4445 1921 4479 1955
rect 4479 1921 4488 1955
rect 4436 1912 4488 1921
rect 4712 1955 4764 1964
rect 4712 1921 4721 1955
rect 4721 1921 4755 1955
rect 4755 1921 4764 1955
rect 4712 1912 4764 1921
rect 9588 1955 9640 1964
rect 9588 1921 9597 1955
rect 9597 1921 9631 1955
rect 9631 1921 9640 1955
rect 9588 1912 9640 1921
rect 13268 1955 13320 1964
rect 13268 1921 13277 1955
rect 13277 1921 13311 1955
rect 13311 1921 13320 1955
rect 13268 1912 13320 1921
rect 12440 1844 12492 1896
rect 12716 1844 12768 1896
rect 13176 1844 13228 1896
rect 9864 1819 9916 1828
rect 9864 1785 9873 1819
rect 9873 1785 9907 1819
rect 9907 1785 9916 1819
rect 9864 1776 9916 1785
rect 10232 1708 10284 1760
rect 11336 1751 11388 1760
rect 11336 1717 11345 1751
rect 11345 1717 11379 1751
rect 11379 1717 11388 1751
rect 11336 1708 11388 1717
rect 14372 1887 14424 1896
rect 14372 1853 14381 1887
rect 14381 1853 14415 1887
rect 14415 1853 14424 1887
rect 14372 1844 14424 1853
rect 14832 1844 14884 1896
rect 14280 1708 14332 1760
rect 2564 1606 2616 1658
rect 2628 1606 2680 1658
rect 2692 1606 2744 1658
rect 2756 1606 2808 1658
rect 2820 1606 2872 1658
rect 6497 1606 6549 1658
rect 6561 1606 6613 1658
rect 6625 1606 6677 1658
rect 6689 1606 6741 1658
rect 6753 1606 6805 1658
rect 10430 1606 10482 1658
rect 10494 1606 10546 1658
rect 10558 1606 10610 1658
rect 10622 1606 10674 1658
rect 10686 1606 10738 1658
rect 14363 1606 14415 1658
rect 14427 1606 14479 1658
rect 14491 1606 14543 1658
rect 14555 1606 14607 1658
rect 14619 1606 14671 1658
rect 9864 1504 9916 1556
rect 11152 1504 11204 1556
rect 11336 1504 11388 1556
rect 14832 1547 14884 1556
rect 14832 1513 14841 1547
rect 14841 1513 14875 1547
rect 14875 1513 14884 1547
rect 14832 1504 14884 1513
rect 1400 1411 1452 1420
rect 1400 1377 1409 1411
rect 1409 1377 1443 1411
rect 1443 1377 1452 1411
rect 1400 1368 1452 1377
rect 3148 1411 3200 1420
rect 3148 1377 3157 1411
rect 3157 1377 3191 1411
rect 3191 1377 3200 1411
rect 3148 1368 3200 1377
rect 9036 1368 9088 1420
rect 13360 1479 13412 1488
rect 13360 1445 13369 1479
rect 13369 1445 13403 1479
rect 13403 1445 13412 1479
rect 13360 1436 13412 1445
rect 13452 1436 13504 1488
rect 15108 1479 15160 1488
rect 15108 1445 15117 1479
rect 15117 1445 15151 1479
rect 15151 1445 15160 1479
rect 15108 1436 15160 1445
rect 9680 1343 9732 1352
rect 9680 1309 9689 1343
rect 9689 1309 9723 1343
rect 9723 1309 9732 1343
rect 9680 1300 9732 1309
rect 10968 1411 11020 1420
rect 10968 1377 10977 1411
rect 10977 1377 11011 1411
rect 11011 1377 11020 1411
rect 10968 1368 11020 1377
rect 11152 1368 11204 1420
rect 12440 1368 12492 1420
rect 13084 1343 13136 1352
rect 13084 1309 13093 1343
rect 13093 1309 13127 1343
rect 13127 1309 13136 1343
rect 13084 1300 13136 1309
rect 1308 1207 1360 1216
rect 1308 1173 1317 1207
rect 1317 1173 1351 1207
rect 1351 1173 1360 1207
rect 1308 1164 1360 1173
rect 3056 1207 3108 1216
rect 3056 1173 3065 1207
rect 3065 1173 3099 1207
rect 3099 1173 3108 1207
rect 3056 1164 3108 1173
rect 8668 1207 8720 1216
rect 8668 1173 8677 1207
rect 8677 1173 8711 1207
rect 8711 1173 8720 1207
rect 8668 1164 8720 1173
rect 11612 1207 11664 1216
rect 11612 1173 11621 1207
rect 11621 1173 11655 1207
rect 11655 1173 11664 1207
rect 11612 1164 11664 1173
rect 15384 1207 15436 1216
rect 15384 1173 15393 1207
rect 15393 1173 15427 1207
rect 15427 1173 15436 1207
rect 15384 1164 15436 1173
rect 1904 1062 1956 1114
rect 1968 1062 2020 1114
rect 2032 1062 2084 1114
rect 2096 1062 2148 1114
rect 2160 1062 2212 1114
rect 5837 1062 5889 1114
rect 5901 1062 5953 1114
rect 5965 1062 6017 1114
rect 6029 1062 6081 1114
rect 6093 1062 6145 1114
rect 9770 1062 9822 1114
rect 9834 1062 9886 1114
rect 9898 1062 9950 1114
rect 9962 1062 10014 1114
rect 10026 1062 10078 1114
rect 13703 1062 13755 1114
rect 13767 1062 13819 1114
rect 13831 1062 13883 1114
rect 13895 1062 13947 1114
rect 13959 1062 14011 1114
rect 3332 960 3384 1012
rect 11612 960 11664 1012
rect 15108 1003 15160 1012
rect 15108 969 15117 1003
rect 15117 969 15151 1003
rect 15151 969 15160 1003
rect 15108 960 15160 969
rect 388 799 440 808
rect 388 765 397 799
rect 397 765 431 799
rect 431 765 440 799
rect 388 756 440 765
rect 1308 756 1360 808
rect 3056 799 3108 808
rect 3056 765 3065 799
rect 3065 765 3099 799
rect 3099 765 3108 799
rect 3056 756 3108 765
rect 4988 756 5040 808
rect 6368 756 6420 808
rect 8668 756 8720 808
rect 11060 799 11112 808
rect 11060 765 11069 799
rect 11069 765 11103 799
rect 11103 765 11112 799
rect 11060 756 11112 765
rect 12624 799 12676 808
rect 12624 765 12633 799
rect 12633 765 12667 799
rect 12667 765 12676 799
rect 12624 756 12676 765
rect 14280 756 14332 808
rect 1308 663 1360 672
rect 1308 629 1317 663
rect 1317 629 1351 663
rect 1351 629 1360 663
rect 1308 620 1360 629
rect 3240 663 3292 672
rect 3240 629 3249 663
rect 3249 629 3283 663
rect 3283 629 3292 663
rect 3240 620 3292 629
rect 5264 620 5316 672
rect 7104 663 7156 672
rect 7104 629 7113 663
rect 7113 629 7147 663
rect 7147 629 7156 663
rect 7104 620 7156 629
rect 8944 663 8996 672
rect 8944 629 8953 663
rect 8953 629 8987 663
rect 8987 629 8996 663
rect 8944 620 8996 629
rect 10784 663 10836 672
rect 10784 629 10793 663
rect 10793 629 10827 663
rect 10827 629 10836 663
rect 10784 620 10836 629
rect 12808 663 12860 672
rect 12808 629 12817 663
rect 12817 629 12851 663
rect 12851 629 12860 663
rect 12808 620 12860 629
rect 14740 620 14792 672
rect 2564 518 2616 570
rect 2628 518 2680 570
rect 2692 518 2744 570
rect 2756 518 2808 570
rect 2820 518 2872 570
rect 6497 518 6549 570
rect 6561 518 6613 570
rect 6625 518 6677 570
rect 6689 518 6741 570
rect 6753 518 6805 570
rect 10430 518 10482 570
rect 10494 518 10546 570
rect 10558 518 10610 570
rect 10622 518 10674 570
rect 10686 518 10738 570
rect 14363 518 14415 570
rect 14427 518 14479 570
rect 14491 518 14543 570
rect 14555 518 14607 570
rect 14619 518 14671 570
<< metal2 >>
rect 12806 13968 12862 13977
rect 12806 13903 12862 13912
rect 3238 13832 3294 13841
rect 3238 13767 3294 13776
rect 5262 13832 5318 13841
rect 5262 13767 5318 13776
rect 6642 13832 6698 13841
rect 6642 13767 6698 13776
rect 8942 13832 8998 13841
rect 8942 13767 8998 13776
rect 10874 13832 10930 13841
rect 10874 13767 10930 13776
rect 1122 13288 1178 13297
rect 1122 13223 1178 13232
rect 846 13152 902 13161
rect 846 13087 902 13096
rect 860 12986 888 13087
rect 1136 12986 1164 13223
rect 1904 13084 2212 13093
rect 1904 13082 1910 13084
rect 1966 13082 1990 13084
rect 2046 13082 2070 13084
rect 2126 13082 2150 13084
rect 2206 13082 2212 13084
rect 1966 13030 1968 13082
rect 2148 13030 2150 13082
rect 1904 13028 1910 13030
rect 1966 13028 1990 13030
rect 2046 13028 2070 13030
rect 2126 13028 2150 13030
rect 2206 13028 2212 13030
rect 1904 13019 2212 13028
rect 3252 12986 3280 13767
rect 5276 12986 5304 13767
rect 5837 13084 6145 13093
rect 5837 13082 5843 13084
rect 5899 13082 5923 13084
rect 5979 13082 6003 13084
rect 6059 13082 6083 13084
rect 6139 13082 6145 13084
rect 5899 13030 5901 13082
rect 6081 13030 6083 13082
rect 5837 13028 5843 13030
rect 5899 13028 5923 13030
rect 5979 13028 6003 13030
rect 6059 13028 6083 13030
rect 6139 13028 6145 13030
rect 5837 13019 6145 13028
rect 6656 12986 6684 13767
rect 8956 12986 8984 13767
rect 9770 13084 10078 13093
rect 9770 13082 9776 13084
rect 9832 13082 9856 13084
rect 9912 13082 9936 13084
rect 9992 13082 10016 13084
rect 10072 13082 10078 13084
rect 9832 13030 9834 13082
rect 10014 13030 10016 13082
rect 9770 13028 9776 13030
rect 9832 13028 9856 13030
rect 9912 13028 9936 13030
rect 9992 13028 10016 13030
rect 10072 13028 10078 13030
rect 9770 13019 10078 13028
rect 10888 12986 10916 13767
rect 12820 12986 12848 13903
rect 14646 13832 14702 13841
rect 14646 13767 14702 13776
rect 13703 13084 14011 13093
rect 13703 13082 13709 13084
rect 13765 13082 13789 13084
rect 13845 13082 13869 13084
rect 13925 13082 13949 13084
rect 14005 13082 14011 13084
rect 13765 13030 13767 13082
rect 13947 13030 13949 13082
rect 13703 13028 13709 13030
rect 13765 13028 13789 13030
rect 13845 13028 13869 13030
rect 13925 13028 13949 13030
rect 14005 13028 14011 13030
rect 13703 13019 14011 13028
rect 14660 12986 14688 13767
rect 15474 13016 15530 13025
rect 848 12980 900 12986
rect 848 12922 900 12928
rect 1124 12980 1176 12986
rect 1124 12922 1176 12928
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 14648 12980 14700 12986
rect 15474 12951 15476 12960
rect 14648 12922 14700 12928
rect 15528 12951 15530 12960
rect 15476 12922 15528 12928
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 388 12708 440 12714
rect 388 12650 440 12656
rect 1308 12708 1360 12714
rect 1308 12650 1360 12656
rect 1400 12708 1452 12714
rect 1400 12650 1452 12656
rect 400 12209 428 12650
rect 756 12368 808 12374
rect 756 12310 808 12316
rect 386 12200 442 12209
rect 386 12135 442 12144
rect 480 11552 532 11558
rect 480 11494 532 11500
rect 492 11257 520 11494
rect 768 11286 796 12310
rect 848 12232 900 12238
rect 848 12174 900 12180
rect 860 11898 888 12174
rect 1320 11898 1348 12650
rect 848 11892 900 11898
rect 848 11834 900 11840
rect 1308 11892 1360 11898
rect 1308 11834 1360 11840
rect 1124 11688 1176 11694
rect 1124 11630 1176 11636
rect 756 11280 808 11286
rect 478 11248 534 11257
rect 756 11222 808 11228
rect 478 11183 534 11192
rect 480 10464 532 10470
rect 480 10406 532 10412
rect 492 10305 520 10406
rect 478 10296 534 10305
rect 478 10231 534 10240
rect 664 10056 716 10062
rect 664 9998 716 10004
rect 676 9722 704 9998
rect 768 9926 796 11222
rect 848 11144 900 11150
rect 848 11086 900 11092
rect 860 10810 888 11086
rect 848 10804 900 10810
rect 848 10746 900 10752
rect 1136 10606 1164 11630
rect 1124 10600 1176 10606
rect 1124 10542 1176 10548
rect 756 9920 808 9926
rect 756 9862 808 9868
rect 664 9716 716 9722
rect 664 9658 716 9664
rect 480 9376 532 9382
rect 478 9344 480 9353
rect 532 9344 534 9353
rect 478 9279 534 9288
rect 768 9042 796 9862
rect 1032 9512 1084 9518
rect 1136 9500 1164 10542
rect 1084 9472 1164 9500
rect 1032 9454 1084 9460
rect 756 9036 808 9042
rect 756 8978 808 8984
rect 1032 8968 1084 8974
rect 1032 8910 1084 8916
rect 756 8832 808 8838
rect 756 8774 808 8780
rect 768 8430 796 8774
rect 1044 8634 1072 8910
rect 1032 8628 1084 8634
rect 1032 8570 1084 8576
rect 1136 8430 1164 9472
rect 756 8424 808 8430
rect 386 8392 442 8401
rect 756 8366 808 8372
rect 1124 8424 1176 8430
rect 1124 8366 1176 8372
rect 386 8327 388 8336
rect 440 8327 442 8336
rect 388 8298 440 8304
rect 1136 7886 1164 8366
rect 1124 7880 1176 7886
rect 1044 7840 1124 7868
rect 480 7744 532 7750
rect 480 7686 532 7692
rect 756 7744 808 7750
rect 756 7686 808 7692
rect 492 7449 520 7686
rect 478 7440 534 7449
rect 768 7410 796 7686
rect 478 7375 534 7384
rect 756 7404 808 7410
rect 756 7346 808 7352
rect 388 7336 440 7342
rect 388 7278 440 7284
rect 400 6322 428 7278
rect 480 6656 532 6662
rect 480 6598 532 6604
rect 492 6497 520 6598
rect 478 6488 534 6497
rect 478 6423 534 6432
rect 388 6316 440 6322
rect 388 6258 440 6264
rect 400 5574 428 6258
rect 664 6180 716 6186
rect 664 6122 716 6128
rect 676 5914 704 6122
rect 664 5908 716 5914
rect 664 5850 716 5856
rect 1044 5778 1072 7840
rect 1124 7822 1176 7828
rect 1308 6860 1360 6866
rect 1308 6802 1360 6808
rect 1320 6322 1348 6802
rect 1412 6662 1440 12650
rect 1492 12368 1544 12374
rect 1492 12310 1544 12316
rect 1504 11286 1532 12310
rect 2332 12102 2360 12718
rect 2564 12540 2872 12549
rect 2564 12538 2570 12540
rect 2626 12538 2650 12540
rect 2706 12538 2730 12540
rect 2786 12538 2810 12540
rect 2866 12538 2872 12540
rect 2626 12486 2628 12538
rect 2808 12486 2810 12538
rect 2564 12484 2570 12486
rect 2626 12484 2650 12486
rect 2706 12484 2730 12486
rect 2786 12484 2810 12486
rect 2866 12484 2872 12486
rect 2564 12475 2872 12484
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 2412 12368 2464 12374
rect 2412 12310 2464 12316
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 1904 11996 2212 12005
rect 1904 11994 1910 11996
rect 1966 11994 1990 11996
rect 2046 11994 2070 11996
rect 2126 11994 2150 11996
rect 2206 11994 2212 11996
rect 1966 11942 1968 11994
rect 2148 11942 2150 11994
rect 1904 11940 1910 11942
rect 1966 11940 1990 11942
rect 2046 11940 2070 11942
rect 2126 11940 2150 11942
rect 2206 11940 2212 11942
rect 1904 11931 2212 11940
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1492 11280 1544 11286
rect 1492 11222 1544 11228
rect 1504 10266 1532 11222
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1504 9110 1532 10202
rect 1596 9330 1624 11630
rect 2332 11626 2360 12038
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2424 11558 2452 12310
rect 3068 11898 3096 12378
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3160 11898 3188 12038
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 1780 10606 1808 11494
rect 2424 11286 2452 11494
rect 2564 11452 2872 11461
rect 2564 11450 2570 11452
rect 2626 11450 2650 11452
rect 2706 11450 2730 11452
rect 2786 11450 2810 11452
rect 2866 11450 2872 11452
rect 2626 11398 2628 11450
rect 2808 11398 2810 11450
rect 2564 11396 2570 11398
rect 2626 11396 2650 11398
rect 2706 11396 2730 11398
rect 2786 11396 2810 11398
rect 2866 11396 2872 11398
rect 2564 11387 2872 11396
rect 2976 11354 3004 11562
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2412 11280 2464 11286
rect 2976 11234 3004 11290
rect 2412 11222 2464 11228
rect 2884 11218 3004 11234
rect 2872 11212 3004 11218
rect 2924 11206 3004 11212
rect 2872 11154 2924 11160
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2964 11008 3016 11014
rect 3068 10996 3096 11086
rect 3016 10968 3096 10996
rect 3148 11008 3200 11014
rect 2964 10950 3016 10956
rect 3148 10950 3200 10956
rect 1904 10908 2212 10917
rect 1904 10906 1910 10908
rect 1966 10906 1990 10908
rect 2046 10906 2070 10908
rect 2126 10906 2150 10908
rect 2206 10906 2212 10908
rect 1966 10854 1968 10906
rect 2148 10854 2150 10906
rect 1904 10852 1910 10854
rect 1966 10852 1990 10854
rect 2046 10852 2070 10854
rect 2126 10852 2150 10854
rect 2206 10852 2212 10854
rect 1904 10843 2212 10852
rect 2608 10606 2636 10950
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2564 10364 2872 10373
rect 2564 10362 2570 10364
rect 2626 10362 2650 10364
rect 2706 10362 2730 10364
rect 2786 10362 2810 10364
rect 2866 10362 2872 10364
rect 2626 10310 2628 10362
rect 2808 10310 2810 10362
rect 2564 10308 2570 10310
rect 2626 10308 2650 10310
rect 2706 10308 2730 10310
rect 2786 10308 2810 10310
rect 2866 10308 2872 10310
rect 2564 10299 2872 10308
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1688 9450 1716 9998
rect 1904 9820 2212 9829
rect 1904 9818 1910 9820
rect 1966 9818 1990 9820
rect 2046 9818 2070 9820
rect 2126 9818 2150 9820
rect 2206 9818 2212 9820
rect 1966 9766 1968 9818
rect 2148 9766 2150 9818
rect 1904 9764 1910 9766
rect 1966 9764 1990 9766
rect 2046 9764 2070 9766
rect 2126 9764 2150 9766
rect 2206 9764 2212 9766
rect 1904 9755 2212 9764
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 1780 9330 1808 9522
rect 2516 9450 2544 10066
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2700 9722 2728 9862
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2792 9382 2820 10134
rect 2976 9518 3004 10950
rect 3160 10062 3188 10950
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3068 9586 3096 9998
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 1596 9302 1808 9330
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 1492 9104 1544 9110
rect 1492 9046 1544 9052
rect 1504 7954 1532 9046
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1504 7206 1532 7890
rect 1596 7886 1624 9302
rect 1780 9178 1808 9302
rect 2564 9276 2872 9285
rect 2564 9274 2570 9276
rect 2626 9274 2650 9276
rect 2706 9274 2730 9276
rect 2786 9274 2810 9276
rect 2866 9274 2872 9276
rect 2626 9222 2628 9274
rect 2808 9222 2810 9274
rect 2564 9220 2570 9222
rect 2626 9220 2650 9222
rect 2706 9220 2730 9222
rect 2786 9220 2810 9222
rect 2866 9220 2872 9222
rect 2564 9211 2872 9220
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2700 8974 2728 9114
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 1904 8732 2212 8741
rect 1904 8730 1910 8732
rect 1966 8730 1990 8732
rect 2046 8730 2070 8732
rect 2126 8730 2150 8732
rect 2206 8730 2212 8732
rect 1966 8678 1968 8730
rect 2148 8678 2150 8730
rect 1904 8676 1910 8678
rect 1966 8676 1990 8678
rect 2046 8676 2070 8678
rect 2126 8676 2150 8678
rect 2206 8676 2212 8678
rect 1904 8667 2212 8676
rect 2608 8634 2636 8774
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2700 8430 2728 8774
rect 2976 8634 3004 9318
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2056 8022 2084 8298
rect 2332 8090 2360 8298
rect 2700 8294 2728 8366
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2564 8188 2872 8197
rect 2564 8186 2570 8188
rect 2626 8186 2650 8188
rect 2706 8186 2730 8188
rect 2786 8186 2810 8188
rect 2866 8186 2872 8188
rect 2626 8134 2628 8186
rect 2808 8134 2810 8186
rect 2564 8132 2570 8134
rect 2626 8132 2650 8134
rect 2706 8132 2730 8134
rect 2786 8132 2810 8134
rect 2866 8132 2872 8134
rect 2564 8123 2872 8132
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2044 8016 2096 8022
rect 2044 7958 2096 7964
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 7002 1532 7142
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 5846 1348 6258
rect 1308 5840 1360 5846
rect 1308 5782 1360 5788
rect 1032 5772 1084 5778
rect 1032 5714 1084 5720
rect 388 5568 440 5574
rect 480 5568 532 5574
rect 388 5510 440 5516
rect 478 5536 480 5545
rect 532 5536 534 5545
rect 400 4690 428 5510
rect 478 5471 534 5480
rect 388 4684 440 4690
rect 388 4626 440 4632
rect 664 4616 716 4622
rect 664 4558 716 4564
rect 676 4282 704 4558
rect 664 4276 716 4282
rect 664 4218 716 4224
rect 478 4176 534 4185
rect 478 4111 534 4120
rect 492 3738 520 4111
rect 1044 4078 1072 5714
rect 1124 4480 1176 4486
rect 1124 4422 1176 4428
rect 1136 4078 1164 4422
rect 1032 4072 1084 4078
rect 1032 4014 1084 4020
rect 1124 4072 1176 4078
rect 1124 4014 1176 4020
rect 940 3936 992 3942
rect 940 3878 992 3884
rect 952 3738 980 3878
rect 480 3732 532 3738
rect 480 3674 532 3680
rect 940 3732 992 3738
rect 940 3674 992 3680
rect 1122 3632 1178 3641
rect 1122 3567 1124 3576
rect 1176 3567 1178 3576
rect 1124 3538 1176 3544
rect 388 2984 440 2990
rect 388 2926 440 2932
rect 400 2689 428 2926
rect 386 2680 442 2689
rect 386 2615 442 2624
rect 1412 1426 1440 6598
rect 1596 5778 1624 7822
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1688 6458 1716 6802
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1780 6254 1808 7754
rect 1904 7644 2212 7653
rect 1904 7642 1910 7644
rect 1966 7642 1990 7644
rect 2046 7642 2070 7644
rect 2126 7642 2150 7644
rect 2206 7642 2212 7644
rect 1966 7590 1968 7642
rect 2148 7590 2150 7642
rect 1904 7588 1910 7590
rect 1966 7588 1990 7590
rect 2046 7588 2070 7590
rect 2126 7588 2150 7590
rect 2206 7588 2212 7590
rect 1904 7579 2212 7588
rect 2240 7206 2268 7890
rect 2332 7546 2360 8026
rect 2976 7954 3004 8570
rect 3068 8090 3096 9522
rect 3160 9450 3188 9998
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3252 9330 3280 12718
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3344 11898 3372 12582
rect 3528 12434 3556 12582
rect 3528 12406 3740 12434
rect 3712 12374 3740 12406
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3436 11150 3464 12174
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4080 11694 4108 11834
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4172 11286 4200 12310
rect 5460 11694 5488 12650
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 12442 5580 12582
rect 5828 12442 5856 12718
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6497 12540 6805 12549
rect 6497 12538 6503 12540
rect 6559 12538 6583 12540
rect 6639 12538 6663 12540
rect 6719 12538 6743 12540
rect 6799 12538 6805 12540
rect 6559 12486 6561 12538
rect 6741 12486 6743 12538
rect 6497 12484 6503 12486
rect 6559 12484 6583 12486
rect 6639 12484 6663 12486
rect 6719 12484 6743 12486
rect 6799 12484 6805 12486
rect 6497 12475 6805 12484
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5816 12436 5868 12442
rect 6840 12434 6868 12582
rect 5816 12378 5868 12384
rect 6748 12406 6868 12434
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3436 9586 3464 11086
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4080 9722 4108 10746
rect 4172 10130 4200 11222
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 4540 9382 4568 9862
rect 4724 9586 4752 9862
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 3160 9302 3280 9330
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2688 7744 2740 7750
rect 3160 7732 3188 9302
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3252 8634 3280 9114
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3436 8430 3464 9318
rect 4540 9110 4568 9318
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4080 8634 4108 8774
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3436 8022 3464 8366
rect 3424 8016 3476 8022
rect 3424 7958 3476 7964
rect 3240 7744 3292 7750
rect 3160 7704 3240 7732
rect 2688 7686 2740 7692
rect 3240 7686 3292 7692
rect 2700 7546 2728 7686
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2564 7100 2872 7109
rect 2564 7098 2570 7100
rect 2626 7098 2650 7100
rect 2706 7098 2730 7100
rect 2786 7098 2810 7100
rect 2866 7098 2872 7100
rect 2626 7046 2628 7098
rect 2808 7046 2810 7098
rect 2564 7044 2570 7046
rect 2626 7044 2650 7046
rect 2706 7044 2730 7046
rect 2786 7044 2810 7046
rect 2866 7044 2872 7046
rect 2564 7035 2872 7044
rect 1904 6556 2212 6565
rect 1904 6554 1910 6556
rect 1966 6554 1990 6556
rect 2046 6554 2070 6556
rect 2126 6554 2150 6556
rect 2206 6554 2212 6556
rect 1966 6502 1968 6554
rect 2148 6502 2150 6554
rect 1904 6500 1910 6502
rect 1966 6500 1990 6502
rect 2046 6500 2070 6502
rect 2126 6500 2150 6502
rect 2206 6500 2212 6502
rect 1904 6491 2212 6500
rect 2976 6458 3004 7142
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 1688 3602 1716 5578
rect 1780 4690 1808 6190
rect 2320 6180 2372 6186
rect 2320 6122 2372 6128
rect 2332 5914 2360 6122
rect 2564 6012 2872 6021
rect 2564 6010 2570 6012
rect 2626 6010 2650 6012
rect 2706 6010 2730 6012
rect 2786 6010 2810 6012
rect 2866 6010 2872 6012
rect 2626 5958 2628 6010
rect 2808 5958 2810 6010
rect 2564 5956 2570 5958
rect 2626 5956 2650 5958
rect 2706 5956 2730 5958
rect 2786 5956 2810 5958
rect 2866 5956 2872 5958
rect 2564 5947 2872 5956
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 3160 5710 3188 6598
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 1904 5468 2212 5477
rect 1904 5466 1910 5468
rect 1966 5466 1990 5468
rect 2046 5466 2070 5468
rect 2126 5466 2150 5468
rect 2206 5466 2212 5468
rect 1966 5414 1968 5466
rect 2148 5414 2150 5466
rect 1904 5412 1910 5414
rect 1966 5412 1990 5414
rect 2046 5412 2070 5414
rect 2126 5412 2150 5414
rect 2206 5412 2212 5414
rect 1904 5403 2212 5412
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2564 4924 2872 4933
rect 2564 4922 2570 4924
rect 2626 4922 2650 4924
rect 2706 4922 2730 4924
rect 2786 4922 2810 4924
rect 2866 4922 2872 4924
rect 2626 4870 2628 4922
rect 2808 4870 2810 4922
rect 2564 4868 2570 4870
rect 2626 4868 2650 4870
rect 2706 4868 2730 4870
rect 2786 4868 2810 4870
rect 2866 4868 2872 4870
rect 2564 4859 2872 4868
rect 2976 4690 3004 4966
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 1904 4380 2212 4389
rect 1904 4378 1910 4380
rect 1966 4378 1990 4380
rect 2046 4378 2070 4380
rect 2126 4378 2150 4380
rect 2206 4378 2212 4380
rect 1966 4326 1968 4378
rect 2148 4326 2150 4378
rect 1904 4324 1910 4326
rect 1966 4324 1990 4326
rect 2046 4324 2070 4326
rect 2126 4324 2150 4326
rect 2206 4324 2212 4326
rect 1904 4315 2212 4324
rect 2332 3942 2360 4626
rect 2412 4548 2464 4554
rect 2412 4490 2464 4496
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2240 3670 2268 3878
rect 2228 3664 2280 3670
rect 2228 3606 2280 3612
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1688 2774 1716 3538
rect 1904 3292 2212 3301
rect 1904 3290 1910 3292
rect 1966 3290 1990 3292
rect 2046 3290 2070 3292
rect 2126 3290 2150 3292
rect 2206 3290 2212 3292
rect 1966 3238 1968 3290
rect 2148 3238 2150 3290
rect 1904 3236 1910 3238
rect 1966 3236 1990 3238
rect 2046 3236 2070 3238
rect 2126 3236 2150 3238
rect 2206 3236 2212 3238
rect 1904 3227 2212 3236
rect 1688 2746 1808 2774
rect 1780 2446 1808 2746
rect 2424 2582 2452 4490
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 2564 3836 2872 3845
rect 2564 3834 2570 3836
rect 2626 3834 2650 3836
rect 2706 3834 2730 3836
rect 2786 3834 2810 3836
rect 2866 3834 2872 3836
rect 2626 3782 2628 3834
rect 2808 3782 2810 3834
rect 2564 3780 2570 3782
rect 2626 3780 2650 3782
rect 2706 3780 2730 3782
rect 2786 3780 2810 3782
rect 2866 3780 2872 3782
rect 2564 3771 2872 3780
rect 3160 3670 3188 3878
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3160 3194 3188 3606
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3252 3074 3280 7686
rect 3620 7410 3648 8366
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4816 7954 4844 8230
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 4344 7268 4396 7274
rect 4344 7210 4396 7216
rect 4356 7002 4384 7210
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4172 6458 4200 6802
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3608 6248 3660 6254
rect 3606 6216 3608 6225
rect 3660 6216 3662 6225
rect 3606 6151 3662 6160
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 4160 6180 4212 6186
rect 4264 6168 4292 6734
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4356 6458 4384 6598
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4212 6140 4384 6168
rect 4160 6122 4212 6128
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3528 5166 3556 5510
rect 3712 5370 3740 6122
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3896 5166 3924 5578
rect 4066 5536 4122 5545
rect 4066 5471 4122 5480
rect 4080 5370 4108 5471
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4172 5250 4200 5714
rect 4356 5658 4384 6140
rect 4448 5846 4476 7890
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4540 6322 4568 7346
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4540 5914 4568 6258
rect 4618 6216 4674 6225
rect 4618 6151 4674 6160
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4356 5630 4568 5658
rect 3988 5234 4200 5250
rect 3976 5228 4212 5234
rect 4028 5222 4160 5228
rect 3976 5170 4028 5176
rect 4160 5170 4212 5176
rect 4540 5166 4568 5630
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 3528 4690 3556 5102
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3712 4690 3740 4966
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4078 3372 4422
rect 3712 4078 3740 4626
rect 3804 4622 3832 5102
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4264 4978 4292 5034
rect 4080 4950 4292 4978
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3160 3046 3280 3074
rect 2564 2748 2872 2757
rect 2564 2746 2570 2748
rect 2626 2746 2650 2748
rect 2706 2746 2730 2748
rect 2786 2746 2810 2748
rect 2866 2746 2872 2748
rect 2626 2694 2628 2746
rect 2808 2694 2810 2746
rect 2564 2692 2570 2694
rect 2626 2692 2650 2694
rect 2706 2692 2730 2694
rect 2786 2692 2810 2694
rect 2866 2692 2872 2694
rect 2564 2683 2872 2692
rect 2412 2576 2464 2582
rect 2412 2518 2464 2524
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 1904 2204 2212 2213
rect 1904 2202 1910 2204
rect 1966 2202 1990 2204
rect 2046 2202 2070 2204
rect 2126 2202 2150 2204
rect 2206 2202 2212 2204
rect 1966 2150 1968 2202
rect 2148 2150 2150 2202
rect 1904 2148 1910 2150
rect 1966 2148 1990 2150
rect 2046 2148 2070 2150
rect 2126 2148 2150 2150
rect 2206 2148 2212 2150
rect 1904 2139 2212 2148
rect 2564 1660 2872 1669
rect 2564 1658 2570 1660
rect 2626 1658 2650 1660
rect 2706 1658 2730 1660
rect 2786 1658 2810 1660
rect 2866 1658 2872 1660
rect 2626 1606 2628 1658
rect 2808 1606 2810 1658
rect 2564 1604 2570 1606
rect 2626 1604 2650 1606
rect 2706 1604 2730 1606
rect 2786 1604 2810 1606
rect 2866 1604 2872 1606
rect 2564 1595 2872 1604
rect 3160 1426 3188 3046
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 1400 1420 1452 1426
rect 1400 1362 1452 1368
rect 3148 1420 3200 1426
rect 3148 1362 3200 1368
rect 1308 1216 1360 1222
rect 1308 1158 1360 1164
rect 3056 1216 3108 1222
rect 3056 1158 3108 1164
rect 1320 814 1348 1158
rect 1904 1116 2212 1125
rect 1904 1114 1910 1116
rect 1966 1114 1990 1116
rect 2046 1114 2070 1116
rect 2126 1114 2150 1116
rect 2206 1114 2212 1116
rect 1966 1062 1968 1114
rect 2148 1062 2150 1114
rect 1904 1060 1910 1062
rect 1966 1060 1990 1062
rect 2046 1060 2070 1062
rect 2126 1060 2150 1062
rect 2206 1060 2212 1062
rect 1904 1051 2212 1060
rect 3068 814 3096 1158
rect 3344 1018 3372 2926
rect 3528 2514 3556 3130
rect 4080 3126 4108 4950
rect 4632 4486 4660 6151
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4724 5574 4752 5714
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4724 5302 4752 5510
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4724 4622 4752 5102
rect 4816 4758 4844 5510
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4540 4146 4568 4422
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4816 4078 4844 4694
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4264 3534 4292 3878
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3896 2650 3924 2926
rect 4448 2774 4476 3878
rect 4816 3602 4844 3878
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4724 2922 4752 3334
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4908 2774 4936 11494
rect 5552 10674 5580 12378
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 5644 11354 5672 12174
rect 5837 11996 6145 12005
rect 5837 11994 5843 11996
rect 5899 11994 5923 11996
rect 5979 11994 6003 11996
rect 6059 11994 6083 11996
rect 6139 11994 6145 11996
rect 5899 11942 5901 11994
rect 6081 11942 6083 11994
rect 5837 11940 5843 11942
rect 5899 11940 5923 11942
rect 5979 11940 6003 11942
rect 6059 11940 6083 11942
rect 6139 11940 6145 11942
rect 5837 11931 6145 11940
rect 6196 11898 6224 12174
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5448 10124 5500 10130
rect 5552 10112 5580 10610
rect 5644 10470 5672 11154
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5500 10084 5580 10112
rect 5448 10066 5500 10072
rect 5184 9722 5212 10066
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5184 9586 5212 9658
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5368 8430 5396 9318
rect 5460 9178 5488 10066
rect 5540 9920 5592 9926
rect 5644 9908 5672 10406
rect 5736 9994 5764 11630
rect 6012 11218 6040 11630
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6012 10996 6040 11154
rect 6012 10968 6224 10996
rect 5837 10908 6145 10917
rect 5837 10906 5843 10908
rect 5899 10906 5923 10908
rect 5979 10906 6003 10908
rect 6059 10906 6083 10908
rect 6139 10906 6145 10908
rect 5899 10854 5901 10906
rect 6081 10854 6083 10906
rect 5837 10852 5843 10854
rect 5899 10852 5923 10854
rect 5979 10852 6003 10854
rect 6059 10852 6083 10854
rect 6139 10852 6145 10854
rect 5837 10843 6145 10852
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5828 10266 5856 10678
rect 6196 10606 6224 10968
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5920 10130 5948 10202
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 6012 10010 6040 10474
rect 6104 10198 6132 10542
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6196 10010 6224 10066
rect 6012 9994 6224 10010
rect 5724 9988 5776 9994
rect 6012 9988 6236 9994
rect 6012 9982 6184 9988
rect 5724 9930 5776 9936
rect 6184 9930 6236 9936
rect 5592 9880 5672 9908
rect 5540 9862 5592 9868
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5000 7342 5028 7686
rect 5092 7342 5120 7686
rect 5368 7546 5396 8366
rect 5460 8362 5488 8910
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5460 7342 5488 8298
rect 5552 7478 5580 9862
rect 5736 8906 5764 9930
rect 5837 9820 6145 9829
rect 5837 9818 5843 9820
rect 5899 9818 5923 9820
rect 5979 9818 6003 9820
rect 6059 9818 6083 9820
rect 6139 9818 6145 9820
rect 5899 9766 5901 9818
rect 6081 9766 6083 9818
rect 5837 9764 5843 9766
rect 5899 9764 5923 9766
rect 5979 9764 6003 9766
rect 6059 9764 6083 9766
rect 6139 9764 6145 9766
rect 5837 9755 6145 9764
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5736 8498 5764 8842
rect 5837 8732 6145 8741
rect 5837 8730 5843 8732
rect 5899 8730 5923 8732
rect 5979 8730 6003 8732
rect 6059 8730 6083 8732
rect 6139 8730 6145 8732
rect 5899 8678 5901 8730
rect 6081 8678 6083 8730
rect 5837 8676 5843 8678
rect 5899 8676 5923 8678
rect 5979 8676 6003 8678
rect 6059 8676 6083 8678
rect 6139 8676 6145 8678
rect 5837 8667 6145 8676
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5644 7342 5672 7890
rect 5837 7644 6145 7653
rect 5837 7642 5843 7644
rect 5899 7642 5923 7644
rect 5979 7642 6003 7644
rect 6059 7642 6083 7644
rect 6139 7642 6145 7644
rect 5899 7590 5901 7642
rect 6081 7590 6083 7642
rect 5837 7588 5843 7590
rect 5899 7588 5923 7590
rect 5979 7588 6003 7590
rect 6059 7588 6083 7590
rect 6139 7588 6145 7590
rect 5837 7579 6145 7588
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5460 6798 5488 7278
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5092 5148 5120 5646
rect 5184 5370 5212 6054
rect 5448 5568 5500 5574
rect 5552 5545 5580 6326
rect 5736 6322 5764 7482
rect 5837 6556 6145 6565
rect 5837 6554 5843 6556
rect 5899 6554 5923 6556
rect 5979 6554 6003 6556
rect 6059 6554 6083 6556
rect 6139 6554 6145 6556
rect 5899 6502 5901 6554
rect 6081 6502 6083 6554
rect 5837 6500 5843 6502
rect 5899 6500 5923 6502
rect 5979 6500 6003 6502
rect 6059 6500 6083 6502
rect 6139 6500 6145 6502
rect 5837 6491 6145 6500
rect 6196 6458 6224 8434
rect 6288 7426 6316 11494
rect 6380 11150 6408 12174
rect 6748 11694 6776 12406
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6497 11452 6805 11461
rect 6497 11450 6503 11452
rect 6559 11450 6583 11452
rect 6639 11450 6663 11452
rect 6719 11450 6743 11452
rect 6799 11450 6805 11452
rect 6559 11398 6561 11450
rect 6741 11398 6743 11450
rect 6497 11396 6503 11398
rect 6559 11396 6583 11398
rect 6639 11396 6663 11398
rect 6719 11396 6743 11398
rect 6799 11396 6805 11398
rect 6497 11387 6805 11396
rect 7760 11286 7788 12242
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11626 8064 12038
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8496 11354 8524 11562
rect 9048 11558 9076 12718
rect 10430 12540 10738 12549
rect 10430 12538 10436 12540
rect 10492 12538 10516 12540
rect 10572 12538 10596 12540
rect 10652 12538 10676 12540
rect 10732 12538 10738 12540
rect 10492 12486 10494 12538
rect 10674 12486 10676 12538
rect 10430 12484 10436 12486
rect 10492 12484 10516 12486
rect 10572 12484 10596 12486
rect 10652 12484 10676 12486
rect 10732 12484 10738 12486
rect 10430 12475 10738 12484
rect 9770 11996 10078 12005
rect 9770 11994 9776 11996
rect 9832 11994 9856 11996
rect 9912 11994 9936 11996
rect 9992 11994 10016 11996
rect 10072 11994 10078 11996
rect 9832 11942 9834 11994
rect 10014 11942 10016 11994
rect 9770 11940 9776 11942
rect 9832 11940 9856 11942
rect 9912 11940 9936 11942
rect 9992 11940 10016 11942
rect 10072 11940 10078 11942
rect 9770 11931 10078 11940
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6380 10674 6408 11086
rect 6472 10742 6500 11154
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6380 10130 6408 10610
rect 6472 10606 6500 10678
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6497 10364 6805 10373
rect 6497 10362 6503 10364
rect 6559 10362 6583 10364
rect 6639 10362 6663 10364
rect 6719 10362 6743 10364
rect 6799 10362 6805 10364
rect 6559 10310 6561 10362
rect 6741 10310 6743 10362
rect 6497 10308 6503 10310
rect 6559 10308 6583 10310
rect 6639 10308 6663 10310
rect 6719 10308 6743 10310
rect 6799 10308 6805 10310
rect 6497 10299 6805 10308
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6380 8090 6408 10066
rect 6497 9276 6805 9285
rect 6497 9274 6503 9276
rect 6559 9274 6583 9276
rect 6639 9274 6663 9276
rect 6719 9274 6743 9276
rect 6799 9274 6805 9276
rect 6559 9222 6561 9274
rect 6741 9222 6743 9274
rect 6497 9220 6503 9222
rect 6559 9220 6583 9222
rect 6639 9220 6663 9222
rect 6719 9220 6743 9222
rect 6799 9220 6805 9222
rect 6497 9211 6805 9220
rect 6840 9178 6868 10542
rect 7760 10198 7788 11222
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7760 9722 7788 10134
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8430 6868 8978
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6497 8188 6805 8197
rect 6497 8186 6503 8188
rect 6559 8186 6583 8188
rect 6639 8186 6663 8188
rect 6719 8186 6743 8188
rect 6799 8186 6805 8188
rect 6559 8134 6561 8186
rect 6741 8134 6743 8186
rect 6497 8132 6503 8134
rect 6559 8132 6583 8134
rect 6639 8132 6663 8134
rect 6719 8132 6743 8134
rect 6799 8132 6805 8134
rect 6497 8123 6805 8132
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6840 7818 6868 8230
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6288 7398 6408 7426
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6288 7002 6316 7210
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6182 6216 6238 6225
rect 6104 5914 6132 6190
rect 6182 6151 6184 6160
rect 6236 6151 6238 6160
rect 6184 6122 6236 6128
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 5632 5568 5684 5574
rect 5448 5510 5500 5516
rect 5538 5536 5594 5545
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5172 5160 5224 5166
rect 5092 5120 5172 5148
rect 5172 5102 5224 5108
rect 5184 4554 5212 5102
rect 5368 4758 5396 5306
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5460 4690 5488 5510
rect 5632 5510 5684 5516
rect 5538 5471 5594 5480
rect 5644 5166 5672 5510
rect 5736 5166 5764 5850
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 5837 5468 6145 5477
rect 5837 5466 5843 5468
rect 5899 5466 5923 5468
rect 5979 5466 6003 5468
rect 6059 5466 6083 5468
rect 6139 5466 6145 5468
rect 5899 5414 5901 5466
rect 6081 5414 6083 5466
rect 5837 5412 5843 5414
rect 5899 5412 5923 5414
rect 5979 5412 6003 5414
rect 6059 5412 6083 5414
rect 6139 5412 6145 5414
rect 5837 5403 6145 5412
rect 6196 5166 6224 5714
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5184 4214 5212 4490
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5092 2836 5120 3130
rect 5184 2990 5212 3946
rect 5276 3942 5304 4558
rect 5460 3942 5488 4626
rect 5552 4078 5580 5034
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4690 5672 4966
rect 5814 4720 5870 4729
rect 5632 4684 5684 4690
rect 5814 4655 5816 4664
rect 5632 4626 5684 4632
rect 5868 4655 5870 4664
rect 5816 4626 5868 4632
rect 5920 4570 5948 5102
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4690 6040 4966
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 5644 4542 5948 4570
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5276 3670 5304 3878
rect 5552 3738 5580 3878
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5276 2836 5304 2926
rect 5644 2854 5672 4542
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5736 4146 5764 4422
rect 5837 4380 6145 4389
rect 5837 4378 5843 4380
rect 5899 4378 5923 4380
rect 5979 4378 6003 4380
rect 6059 4378 6083 4380
rect 6139 4378 6145 4380
rect 5899 4326 5901 4378
rect 6081 4326 6083 4378
rect 5837 4324 5843 4326
rect 5899 4324 5923 4326
rect 5979 4324 6003 4326
rect 6059 4324 6083 4326
rect 6139 4324 6145 4326
rect 5837 4315 6145 4324
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 6196 4078 6224 4626
rect 6288 4078 6316 5034
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 5837 3292 6145 3301
rect 5837 3290 5843 3292
rect 5899 3290 5923 3292
rect 5979 3290 6003 3292
rect 6059 3290 6083 3292
rect 6139 3290 6145 3292
rect 5899 3238 5901 3290
rect 6081 3238 6083 3290
rect 5837 3236 5843 3238
rect 5899 3236 5923 3238
rect 5979 3236 6003 3238
rect 6059 3236 6083 3238
rect 6139 3236 6145 3238
rect 5837 3227 6145 3236
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 5092 2808 5304 2836
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 4448 2746 4752 2774
rect 4908 2746 5028 2774
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4080 1873 4108 2042
rect 4448 1970 4476 2246
rect 4724 1970 4752 2746
rect 4436 1964 4488 1970
rect 4436 1906 4488 1912
rect 4712 1964 4764 1970
rect 4712 1906 4764 1912
rect 4066 1864 4122 1873
rect 4066 1799 4122 1808
rect 3332 1012 3384 1018
rect 3332 954 3384 960
rect 5000 814 5028 2746
rect 5837 2204 6145 2213
rect 5837 2202 5843 2204
rect 5899 2202 5923 2204
rect 5979 2202 6003 2204
rect 6059 2202 6083 2204
rect 6139 2202 6145 2204
rect 5899 2150 5901 2202
rect 6081 2150 6083 2202
rect 5837 2148 5843 2150
rect 5899 2148 5923 2150
rect 5979 2148 6003 2150
rect 6059 2148 6083 2150
rect 6139 2148 6145 2150
rect 5837 2139 6145 2148
rect 6196 2038 6224 2926
rect 6184 2032 6236 2038
rect 6184 1974 6236 1980
rect 5837 1116 6145 1125
rect 5837 1114 5843 1116
rect 5899 1114 5923 1116
rect 5979 1114 6003 1116
rect 6059 1114 6083 1116
rect 6139 1114 6145 1116
rect 5899 1062 5901 1114
rect 6081 1062 6083 1114
rect 5837 1060 5843 1062
rect 5899 1060 5923 1062
rect 5979 1060 6003 1062
rect 6059 1060 6083 1062
rect 6139 1060 6145 1062
rect 5837 1051 6145 1060
rect 6380 814 6408 7398
rect 7760 7342 7788 9658
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8496 9178 8524 9386
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 7852 7750 7880 8366
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8036 8090 8064 8230
rect 8496 8090 8524 8366
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 6497 7100 6805 7109
rect 6497 7098 6503 7100
rect 6559 7098 6583 7100
rect 6639 7098 6663 7100
rect 6719 7098 6743 7100
rect 6799 7098 6805 7100
rect 6559 7046 6561 7098
rect 6741 7046 6743 7098
rect 6497 7044 6503 7046
rect 6559 7044 6583 7046
rect 6639 7044 6663 7046
rect 6719 7044 6743 7046
rect 6799 7044 6805 7046
rect 6497 7035 6805 7044
rect 7760 6866 7788 7142
rect 7852 6866 7880 7686
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6497 6012 6805 6021
rect 6497 6010 6503 6012
rect 6559 6010 6583 6012
rect 6639 6010 6663 6012
rect 6719 6010 6743 6012
rect 6799 6010 6805 6012
rect 6559 5958 6561 6010
rect 6741 5958 6743 6010
rect 6497 5956 6503 5958
rect 6559 5956 6583 5958
rect 6639 5956 6663 5958
rect 6719 5956 6743 5958
rect 6799 5956 6805 5958
rect 6497 5947 6805 5956
rect 6497 4924 6805 4933
rect 6497 4922 6503 4924
rect 6559 4922 6583 4924
rect 6639 4922 6663 4924
rect 6719 4922 6743 4924
rect 6799 4922 6805 4924
rect 6559 4870 6561 4922
rect 6741 4870 6743 4922
rect 6497 4868 6503 4870
rect 6559 4868 6583 4870
rect 6639 4868 6663 4870
rect 6719 4868 6743 4870
rect 6799 4868 6805 4870
rect 6497 4859 6805 4868
rect 6840 4808 6868 6190
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7208 5166 7236 5714
rect 7300 5370 7328 6054
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7300 5166 7328 5306
rect 7668 5166 7696 5714
rect 7012 5160 7064 5166
rect 7196 5160 7248 5166
rect 7064 5120 7144 5148
rect 7012 5102 7064 5108
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7024 4826 7052 4966
rect 6748 4780 6868 4808
rect 7012 4820 7064 4826
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6564 4214 6592 4422
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6656 4078 6684 4422
rect 6748 4078 6776 4780
rect 7012 4762 7064 4768
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6840 4146 6868 4626
rect 6828 4140 6880 4146
rect 6880 4100 6960 4128
rect 6828 4082 6880 4088
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6497 3836 6805 3845
rect 6497 3834 6503 3836
rect 6559 3834 6583 3836
rect 6639 3834 6663 3836
rect 6719 3834 6743 3836
rect 6799 3834 6805 3836
rect 6559 3782 6561 3834
rect 6741 3782 6743 3834
rect 6497 3780 6503 3782
rect 6559 3780 6583 3782
rect 6639 3780 6663 3782
rect 6719 3780 6743 3782
rect 6799 3780 6805 3782
rect 6497 3771 6805 3780
rect 6840 3670 6868 3946
rect 6932 3738 6960 4100
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6497 2748 6805 2757
rect 6497 2746 6503 2748
rect 6559 2746 6583 2748
rect 6639 2746 6663 2748
rect 6719 2746 6743 2748
rect 6799 2746 6805 2748
rect 6559 2694 6561 2746
rect 6741 2694 6743 2746
rect 6497 2692 6503 2694
rect 6559 2692 6583 2694
rect 6639 2692 6663 2694
rect 6719 2692 6743 2694
rect 6799 2692 6805 2694
rect 6497 2683 6805 2692
rect 6840 2650 6868 3470
rect 7024 2990 7052 4626
rect 7116 4622 7144 5120
rect 7196 5102 7248 5108
rect 7288 5160 7340 5166
rect 7656 5160 7708 5166
rect 7288 5102 7340 5108
rect 7576 5120 7656 5148
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7116 4214 7144 4558
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 7208 4162 7236 5102
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4826 7420 4966
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7484 4282 7512 4762
rect 7576 4622 7604 5120
rect 7656 5102 7708 5108
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7576 4486 7604 4558
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7116 3584 7144 4150
rect 7208 4134 7512 4162
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7196 3596 7248 3602
rect 7116 3556 7196 3584
rect 7196 3538 7248 3544
rect 7300 3194 7328 4014
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3466 7420 3878
rect 7484 3670 7512 4134
rect 7852 3942 7880 4966
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7288 3052 7340 3058
rect 7484 3040 7512 3606
rect 7576 3602 7604 3674
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7340 3012 7512 3040
rect 7288 2994 7340 3000
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7024 2038 7052 2450
rect 7576 2446 7604 3334
rect 7760 2854 7788 3402
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7944 2106 7972 7210
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 4214 8064 6598
rect 8220 5846 8248 7142
rect 8496 6866 8524 8026
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8496 6322 8524 6802
rect 8680 6458 8708 7890
rect 8864 6662 8892 8978
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8956 6934 8984 7822
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8956 6186 8984 6870
rect 8944 6180 8996 6186
rect 8772 6140 8944 6168
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8128 4554 8156 5714
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 8128 3466 8156 4490
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 8220 2990 8248 5782
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8312 5166 8340 5238
rect 8680 5166 8708 5850
rect 8772 5302 8800 6140
rect 8944 6122 8996 6128
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 8772 5166 8800 5238
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4486 8340 4966
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8496 4554 8524 4626
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8404 4146 8432 4422
rect 8496 4214 8524 4490
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8680 4078 8708 5102
rect 8864 4826 8892 5646
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8864 4282 8892 4762
rect 8956 4758 8984 4966
rect 8944 4752 8996 4758
rect 8944 4694 8996 4700
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8588 3194 8616 3470
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8864 3126 8892 3470
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 8956 3058 8984 3946
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 7012 2032 7064 2038
rect 7012 1974 7064 1980
rect 6497 1660 6805 1669
rect 6497 1658 6503 1660
rect 6559 1658 6583 1660
rect 6639 1658 6663 1660
rect 6719 1658 6743 1660
rect 6799 1658 6805 1660
rect 6559 1606 6561 1658
rect 6741 1606 6743 1658
rect 6497 1604 6503 1606
rect 6559 1604 6583 1606
rect 6639 1604 6663 1606
rect 6719 1604 6743 1606
rect 6799 1604 6805 1606
rect 6497 1595 6805 1604
rect 9048 1426 9076 11494
rect 10430 11452 10738 11461
rect 10430 11450 10436 11452
rect 10492 11450 10516 11452
rect 10572 11450 10596 11452
rect 10652 11450 10676 11452
rect 10732 11450 10738 11452
rect 10492 11398 10494 11450
rect 10674 11398 10676 11450
rect 10430 11396 10436 11398
rect 10492 11396 10516 11398
rect 10572 11396 10596 11398
rect 10652 11396 10676 11398
rect 10732 11396 10738 11398
rect 10430 11387 10738 11396
rect 9770 10908 10078 10917
rect 9770 10906 9776 10908
rect 9832 10906 9856 10908
rect 9912 10906 9936 10908
rect 9992 10906 10016 10908
rect 10072 10906 10078 10908
rect 9832 10854 9834 10906
rect 10014 10854 10016 10906
rect 9770 10852 9776 10854
rect 9832 10852 9856 10854
rect 9912 10852 9936 10854
rect 9992 10852 10016 10854
rect 10072 10852 10078 10854
rect 9770 10843 10078 10852
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9232 10266 9260 10406
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9508 9178 9536 10474
rect 9876 10266 9904 10542
rect 10980 10452 11008 12718
rect 12360 10606 12388 12718
rect 13703 11996 14011 12005
rect 13703 11994 13709 11996
rect 13765 11994 13789 11996
rect 13845 11994 13869 11996
rect 13925 11994 13949 11996
rect 14005 11994 14011 11996
rect 13765 11942 13767 11994
rect 13947 11942 13949 11994
rect 13703 11940 13709 11942
rect 13765 11940 13789 11942
rect 13845 11940 13869 11942
rect 13925 11940 13949 11942
rect 14005 11940 14011 11942
rect 13703 11931 14011 11940
rect 13703 10908 14011 10917
rect 13703 10906 13709 10908
rect 13765 10906 13789 10908
rect 13845 10906 13869 10908
rect 13925 10906 13949 10908
rect 14005 10906 14011 10908
rect 13765 10854 13767 10906
rect 13947 10854 13949 10906
rect 13703 10852 13709 10854
rect 13765 10852 13789 10854
rect 13845 10852 13869 10854
rect 13925 10852 13949 10854
rect 14005 10852 14011 10854
rect 13703 10843 14011 10852
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 11060 10464 11112 10470
rect 10980 10424 11060 10452
rect 11060 10406 11112 10412
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 10430 10364 10738 10373
rect 10430 10362 10436 10364
rect 10492 10362 10516 10364
rect 10572 10362 10596 10364
rect 10652 10362 10676 10364
rect 10732 10362 10738 10364
rect 10492 10310 10494 10362
rect 10674 10310 10676 10362
rect 10430 10308 10436 10310
rect 10492 10308 10516 10310
rect 10572 10308 10596 10310
rect 10652 10308 10676 10310
rect 10732 10308 10738 10310
rect 10430 10299 10738 10308
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9770 9820 10078 9829
rect 9770 9818 9776 9820
rect 9832 9818 9856 9820
rect 9912 9818 9936 9820
rect 9992 9818 10016 9820
rect 10072 9818 10078 9820
rect 9832 9766 9834 9818
rect 10014 9766 10016 9818
rect 9770 9764 9776 9766
rect 9832 9764 9856 9766
rect 9912 9764 9936 9766
rect 9992 9764 10016 9766
rect 10072 9764 10078 9766
rect 9770 9755 10078 9764
rect 10692 9512 10744 9518
rect 10744 9460 10824 9466
rect 10692 9454 10824 9460
rect 9772 9444 9824 9450
rect 10704 9438 10824 9454
rect 9772 9386 9824 9392
rect 9784 9178 9812 9386
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9416 8090 9444 8434
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9140 6322 9168 6666
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9232 6254 9260 6938
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6458 9536 6598
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9232 5574 9260 6190
rect 9416 5914 9444 6190
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9600 5760 9628 8978
rect 9770 8732 10078 8741
rect 9770 8730 9776 8732
rect 9832 8730 9856 8732
rect 9912 8730 9936 8732
rect 9992 8730 10016 8732
rect 10072 8730 10078 8732
rect 9832 8678 9834 8730
rect 10014 8678 10016 8730
rect 9770 8676 9776 8678
rect 9832 8676 9856 8678
rect 9912 8676 9936 8678
rect 9992 8676 10016 8678
rect 10072 8676 10078 8678
rect 9770 8667 10078 8676
rect 9680 8424 9732 8430
rect 9732 8384 9904 8412
rect 9680 8366 9732 8372
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 7188 9720 7890
rect 9876 7818 9904 8384
rect 10152 8090 10180 9318
rect 10430 9276 10738 9285
rect 10430 9274 10436 9276
rect 10492 9274 10516 9276
rect 10572 9274 10596 9276
rect 10652 9274 10676 9276
rect 10732 9274 10738 9276
rect 10492 9222 10494 9274
rect 10674 9222 10676 9274
rect 10430 9220 10436 9222
rect 10492 9220 10516 9222
rect 10572 9220 10596 9222
rect 10652 9220 10676 9222
rect 10732 9220 10738 9222
rect 10430 9211 10738 9220
rect 10796 9178 10824 9438
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10430 8188 10738 8197
rect 10430 8186 10436 8188
rect 10492 8186 10516 8188
rect 10572 8186 10596 8188
rect 10652 8186 10676 8188
rect 10732 8186 10738 8188
rect 10492 8134 10494 8186
rect 10674 8134 10676 8186
rect 10430 8132 10436 8134
rect 10492 8132 10516 8134
rect 10572 8132 10596 8134
rect 10652 8132 10676 8134
rect 10732 8132 10738 8134
rect 10430 8123 10738 8132
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 10152 7750 10180 8026
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 9770 7644 10078 7653
rect 9770 7642 9776 7644
rect 9832 7642 9856 7644
rect 9912 7642 9936 7644
rect 9992 7642 10016 7644
rect 10072 7642 10078 7644
rect 9832 7590 9834 7642
rect 10014 7590 10016 7642
rect 9770 7588 9776 7590
rect 9832 7588 9856 7590
rect 9912 7588 9936 7590
rect 9992 7588 10016 7590
rect 10072 7588 10078 7590
rect 9770 7579 10078 7588
rect 9864 7200 9916 7206
rect 9692 7160 9864 7188
rect 9864 7142 9916 7148
rect 9876 6798 9904 7142
rect 10152 6798 10180 7686
rect 10336 7002 10364 7890
rect 10888 7426 10916 9318
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10796 7398 10916 7426
rect 10796 7274 10824 7398
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 10430 7100 10738 7109
rect 10430 7098 10436 7100
rect 10492 7098 10516 7100
rect 10572 7098 10596 7100
rect 10652 7098 10676 7100
rect 10732 7098 10738 7100
rect 10492 7046 10494 7098
rect 10674 7046 10676 7098
rect 10430 7044 10436 7046
rect 10492 7044 10516 7046
rect 10572 7044 10596 7046
rect 10652 7044 10676 7046
rect 10732 7044 10738 7046
rect 10430 7035 10738 7044
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 9770 6556 10078 6565
rect 9770 6554 9776 6556
rect 9832 6554 9856 6556
rect 9912 6554 9936 6556
rect 9992 6554 10016 6556
rect 10072 6554 10078 6556
rect 9832 6502 9834 6554
rect 10014 6502 10016 6554
rect 9770 6500 9776 6502
rect 9832 6500 9856 6502
rect 9912 6500 9936 6502
rect 9992 6500 10016 6502
rect 10072 6500 10078 6502
rect 9770 6491 10078 6500
rect 10152 6322 10180 6734
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 9508 5732 9628 5760
rect 9680 5772 9732 5778
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9324 3534 9352 4082
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9508 2922 9536 5732
rect 9680 5714 9732 5720
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 5166 9628 5510
rect 9692 5302 9720 5714
rect 10336 5574 10364 6938
rect 10980 6866 11008 8298
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10430 6012 10738 6021
rect 10430 6010 10436 6012
rect 10492 6010 10516 6012
rect 10572 6010 10596 6012
rect 10652 6010 10676 6012
rect 10732 6010 10738 6012
rect 10492 5958 10494 6010
rect 10674 5958 10676 6010
rect 10430 5956 10436 5958
rect 10492 5956 10516 5958
rect 10572 5956 10596 5958
rect 10652 5956 10676 5958
rect 10732 5956 10738 5958
rect 10430 5947 10738 5956
rect 10796 5778 10824 6122
rect 10874 5944 10930 5953
rect 10874 5879 10930 5888
rect 10888 5778 10916 5879
rect 10980 5778 11008 6394
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 9770 5468 10078 5477
rect 9770 5466 9776 5468
rect 9832 5466 9856 5468
rect 9912 5466 9936 5468
rect 9992 5466 10016 5468
rect 10072 5466 10078 5468
rect 9832 5414 9834 5466
rect 10014 5414 10016 5466
rect 9770 5412 9776 5414
rect 9832 5412 9856 5414
rect 9912 5412 9936 5414
rect 9992 5412 10016 5414
rect 10072 5412 10078 5414
rect 9770 5403 10078 5412
rect 10980 5370 11008 5714
rect 11072 5658 11100 10406
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11716 9042 11744 9522
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9110 11928 9318
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11164 6866 11192 7754
rect 11440 6866 11468 8978
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11532 7274 11560 8570
rect 11716 7954 11744 8978
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 8634 12388 8910
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11716 7410 11744 7890
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7546 12296 7822
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11164 5914 11192 6802
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11256 5846 11284 6258
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11348 5778 11376 6666
rect 11716 6322 11744 7346
rect 12452 6610 12480 10406
rect 13703 9820 14011 9829
rect 13703 9818 13709 9820
rect 13765 9818 13789 9820
rect 13845 9818 13869 9820
rect 13925 9818 13949 9820
rect 14005 9818 14011 9820
rect 13765 9766 13767 9818
rect 13947 9766 13949 9818
rect 13703 9764 13709 9766
rect 13765 9764 13789 9766
rect 13845 9764 13869 9766
rect 13925 9764 13949 9766
rect 14005 9764 14011 9766
rect 13703 9755 14011 9764
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 13096 9110 13124 9386
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 13096 8022 13124 9046
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 8430 13400 8774
rect 13464 8634 13492 9522
rect 14108 8838 14136 12718
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 14363 12540 14671 12549
rect 14363 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14585 12538 14609 12540
rect 14665 12538 14671 12540
rect 14425 12486 14427 12538
rect 14607 12486 14609 12538
rect 14363 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14585 12484 14609 12486
rect 14665 12484 14671 12486
rect 14363 12475 14671 12484
rect 15120 12442 15148 12650
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 14363 11452 14671 11461
rect 14363 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14585 11450 14609 11452
rect 14665 11450 14671 11452
rect 14425 11398 14427 11450
rect 14607 11398 14609 11450
rect 14363 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14585 11396 14609 11398
rect 14665 11396 14671 11398
rect 14363 11387 14671 11396
rect 15120 11354 15148 12242
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 14363 10364 14671 10373
rect 14363 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14585 10362 14609 10364
rect 14665 10362 14671 10364
rect 14425 10310 14427 10362
rect 14607 10310 14609 10362
rect 14363 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14585 10308 14609 10310
rect 14665 10308 14671 10310
rect 14363 10299 14671 10308
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14363 9276 14671 9285
rect 14363 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14585 9274 14609 9276
rect 14665 9274 14671 9276
rect 14425 9222 14427 9274
rect 14607 9222 14609 9274
rect 14363 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14585 9220 14609 9222
rect 14665 9220 14671 9222
rect 14363 9211 14671 9220
rect 14752 9110 14780 9318
rect 14844 9178 14872 9386
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14740 9104 14792 9110
rect 14740 9046 14792 9052
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 13556 8634 13584 8774
rect 13703 8732 14011 8741
rect 13703 8730 13709 8732
rect 13765 8730 13789 8732
rect 13845 8730 13869 8732
rect 13925 8730 13949 8732
rect 14005 8730 14011 8732
rect 13765 8678 13767 8730
rect 13947 8678 13949 8730
rect 13703 8676 13709 8678
rect 13765 8676 13789 8678
rect 13845 8676 13869 8678
rect 13925 8676 13949 8678
rect 14005 8676 14011 8678
rect 13703 8667 14011 8676
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 13280 6866 13308 8230
rect 13372 7750 13400 8366
rect 13556 8294 13584 8434
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13372 7342 13400 7686
rect 13464 7342 13492 7686
rect 13556 7546 13584 7686
rect 13703 7644 14011 7653
rect 13703 7642 13709 7644
rect 13765 7642 13789 7644
rect 13845 7642 13869 7644
rect 13925 7642 13949 7644
rect 14005 7642 14011 7644
rect 13765 7590 13767 7642
rect 13947 7590 13949 7642
rect 13703 7588 13709 7590
rect 13765 7588 13789 7590
rect 13845 7588 13869 7590
rect 13925 7588 13949 7590
rect 14005 7588 14011 7590
rect 13703 7579 14011 7588
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13556 6866 13584 7346
rect 13924 6866 13952 7414
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14016 7002 14044 7278
rect 14004 6996 14056 7002
rect 14108 6984 14136 8774
rect 14200 7954 14228 8774
rect 14363 8188 14671 8197
rect 14363 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14585 8186 14609 8188
rect 14665 8186 14671 8188
rect 14425 8134 14427 8186
rect 14607 8134 14609 8186
rect 14363 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14585 8132 14609 8134
rect 14665 8132 14671 8134
rect 14363 8123 14671 8132
rect 14752 7970 14780 8910
rect 14844 8566 14872 9114
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14188 7948 14240 7954
rect 14752 7942 14872 7970
rect 14188 7890 14240 7896
rect 14200 7546 14228 7890
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14752 7546 14780 7822
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14363 7100 14671 7109
rect 14363 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14585 7098 14609 7100
rect 14665 7098 14671 7100
rect 14425 7046 14427 7098
rect 14607 7046 14609 7098
rect 14363 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14585 7044 14609 7046
rect 14665 7044 14671 7046
rect 14363 7035 14671 7044
rect 14108 6956 14228 6984
rect 14004 6938 14056 6944
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 14016 6746 14044 6938
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 13556 6718 14044 6746
rect 12452 6582 12664 6610
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11992 6118 12020 6258
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11072 5630 11192 5658
rect 11440 5642 11468 6054
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9586 4720 9642 4729
rect 9586 4655 9588 4664
rect 9640 4655 9642 4664
rect 9588 4626 9640 4632
rect 9968 4554 9996 5170
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9600 2854 9628 3130
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9600 2650 9628 2790
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9600 1970 9628 2586
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 9036 1420 9088 1426
rect 9036 1362 9088 1368
rect 9692 1358 9720 4422
rect 9770 4380 10078 4389
rect 9770 4378 9776 4380
rect 9832 4378 9856 4380
rect 9912 4378 9936 4380
rect 9992 4378 10016 4380
rect 10072 4378 10078 4380
rect 9832 4326 9834 4378
rect 10014 4326 10016 4378
rect 9770 4324 9776 4326
rect 9832 4324 9856 4326
rect 9912 4324 9936 4326
rect 9992 4324 10016 4326
rect 10072 4324 10078 4326
rect 9770 4315 10078 4324
rect 10152 4214 10180 4966
rect 10430 4924 10738 4933
rect 10430 4922 10436 4924
rect 10492 4922 10516 4924
rect 10572 4922 10596 4924
rect 10652 4922 10676 4924
rect 10732 4922 10738 4924
rect 10492 4870 10494 4922
rect 10674 4870 10676 4922
rect 10430 4868 10436 4870
rect 10492 4868 10516 4870
rect 10572 4868 10596 4870
rect 10652 4868 10676 4870
rect 10732 4868 10738 4870
rect 10430 4859 10738 4868
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10152 3738 10180 3946
rect 10244 3942 10272 4694
rect 10506 4584 10562 4593
rect 10506 4519 10562 4528
rect 10520 4214 10548 4519
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10336 3738 10364 4014
rect 10796 4010 10824 5170
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10876 4072 10928 4078
rect 10874 4040 10876 4049
rect 10928 4040 10930 4049
rect 10784 4004 10836 4010
rect 10874 3975 10930 3984
rect 10784 3946 10836 3952
rect 10430 3836 10738 3845
rect 10430 3834 10436 3836
rect 10492 3834 10516 3836
rect 10572 3834 10596 3836
rect 10652 3834 10676 3836
rect 10732 3834 10738 3836
rect 10492 3782 10494 3834
rect 10674 3782 10676 3834
rect 10430 3780 10436 3782
rect 10492 3780 10516 3782
rect 10572 3780 10596 3782
rect 10652 3780 10676 3782
rect 10732 3780 10738 3782
rect 10430 3771 10738 3780
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10796 3670 10824 3946
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 9770 3292 10078 3301
rect 9770 3290 9776 3292
rect 9832 3290 9856 3292
rect 9912 3290 9936 3292
rect 9992 3290 10016 3292
rect 10072 3290 10078 3292
rect 9832 3238 9834 3290
rect 10014 3238 10016 3290
rect 9770 3236 9776 3238
rect 9832 3236 9856 3238
rect 9912 3236 9936 3238
rect 9992 3236 10016 3238
rect 10072 3236 10078 3238
rect 9770 3227 10078 3236
rect 10244 3194 10272 3606
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10244 2514 10272 3130
rect 10336 2514 10364 3470
rect 10704 3058 10732 3538
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10796 2774 10824 3606
rect 10888 3534 10916 3878
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 3194 10916 3470
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 10888 2774 10916 2858
rect 10430 2748 10738 2757
rect 10430 2746 10436 2748
rect 10492 2746 10516 2748
rect 10572 2746 10596 2748
rect 10652 2746 10676 2748
rect 10732 2746 10738 2748
rect 10796 2746 10916 2774
rect 10492 2694 10494 2746
rect 10674 2694 10676 2746
rect 10430 2692 10436 2694
rect 10492 2692 10516 2694
rect 10572 2692 10596 2694
rect 10652 2692 10676 2694
rect 10732 2692 10738 2694
rect 10430 2683 10738 2692
rect 10888 2582 10916 2746
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 9770 2204 10078 2213
rect 9770 2202 9776 2204
rect 9832 2202 9856 2204
rect 9912 2202 9936 2204
rect 9992 2202 10016 2204
rect 10072 2202 10078 2204
rect 9832 2150 9834 2202
rect 10014 2150 10016 2202
rect 9770 2148 9776 2150
rect 9832 2148 9856 2150
rect 9912 2148 9936 2150
rect 9992 2148 10016 2150
rect 10072 2148 10078 2150
rect 9770 2139 10078 2148
rect 9864 1828 9916 1834
rect 9864 1770 9916 1776
rect 9876 1562 9904 1770
rect 10244 1766 10272 2450
rect 10232 1760 10284 1766
rect 10232 1702 10284 1708
rect 10430 1660 10738 1669
rect 10430 1658 10436 1660
rect 10492 1658 10516 1660
rect 10572 1658 10596 1660
rect 10652 1658 10676 1660
rect 10732 1658 10738 1660
rect 10492 1606 10494 1658
rect 10674 1606 10676 1658
rect 10430 1604 10436 1606
rect 10492 1604 10516 1606
rect 10572 1604 10596 1606
rect 10652 1604 10676 1606
rect 10732 1604 10738 1606
rect 10430 1595 10738 1604
rect 9864 1556 9916 1562
rect 9864 1498 9916 1504
rect 10980 1426 11008 4966
rect 11072 4826 11100 5102
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11072 3738 11100 4014
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11164 3618 11192 5630
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 12544 5370 12572 6122
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12544 4706 12572 5306
rect 12452 4690 12572 4706
rect 12440 4684 12572 4690
rect 12492 4678 12572 4684
rect 12440 4626 12492 4632
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11242 4040 11298 4049
rect 11242 3975 11298 3984
rect 11072 3590 11192 3618
rect 10968 1420 11020 1426
rect 10968 1362 11020 1368
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 8668 1216 8720 1222
rect 8668 1158 8720 1164
rect 8680 814 8708 1158
rect 9770 1116 10078 1125
rect 9770 1114 9776 1116
rect 9832 1114 9856 1116
rect 9912 1114 9936 1116
rect 9992 1114 10016 1116
rect 10072 1114 10078 1116
rect 9832 1062 9834 1114
rect 10014 1062 10016 1114
rect 9770 1060 9776 1062
rect 9832 1060 9856 1062
rect 9912 1060 9936 1062
rect 9992 1060 10016 1062
rect 10072 1060 10078 1062
rect 9770 1051 10078 1060
rect 11072 814 11100 3590
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11164 2582 11192 2926
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11164 1562 11192 2518
rect 11256 2514 11284 3975
rect 11348 3534 11376 4422
rect 11440 4282 11468 4558
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 12544 3738 12572 4678
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11348 3346 11376 3470
rect 11348 3318 11468 3346
rect 11440 2854 11468 3318
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11440 2514 11468 2790
rect 11624 2564 11652 2790
rect 11704 2576 11756 2582
rect 11624 2536 11704 2564
rect 11704 2518 11756 2524
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 12440 1896 12492 1902
rect 12440 1838 12492 1844
rect 11336 1760 11388 1766
rect 11336 1702 11388 1708
rect 11348 1562 11376 1702
rect 11152 1556 11204 1562
rect 11152 1498 11204 1504
rect 11336 1556 11388 1562
rect 11336 1498 11388 1504
rect 11164 1426 11192 1498
rect 12452 1426 12480 1838
rect 11152 1420 11204 1426
rect 11152 1362 11204 1368
rect 12440 1420 12492 1426
rect 12440 1362 12492 1368
rect 11612 1216 11664 1222
rect 11612 1158 11664 1164
rect 11624 1018 11652 1158
rect 11612 1012 11664 1018
rect 11612 954 11664 960
rect 12636 814 12664 6582
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12728 6254 12756 6394
rect 13556 6322 13584 6718
rect 13703 6556 14011 6565
rect 13703 6554 13709 6556
rect 13765 6554 13789 6556
rect 13845 6554 13869 6556
rect 13925 6554 13949 6556
rect 14005 6554 14011 6556
rect 13765 6502 13767 6554
rect 13947 6502 13949 6554
rect 13703 6500 13709 6502
rect 13765 6500 13789 6502
rect 13845 6500 13869 6502
rect 13925 6500 13949 6502
rect 14005 6500 14011 6502
rect 13703 6491 14011 6500
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 14108 6254 14136 6802
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5953 13768 6054
rect 13726 5944 13782 5953
rect 13726 5879 13782 5888
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 13096 5302 13124 5782
rect 13703 5468 14011 5477
rect 13703 5466 13709 5468
rect 13765 5466 13789 5468
rect 13845 5466 13869 5468
rect 13925 5466 13949 5468
rect 14005 5466 14011 5468
rect 13765 5414 13767 5466
rect 13947 5414 13949 5466
rect 13703 5412 13709 5414
rect 13765 5412 13789 5414
rect 13845 5412 13869 5414
rect 13925 5412 13949 5414
rect 14005 5412 14011 5414
rect 13703 5403 14011 5412
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12728 4826 12756 5102
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12820 4214 12848 4422
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 13096 3602 13124 5102
rect 13924 4690 13952 5170
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14016 4826 14044 4966
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 13280 4078 13308 4626
rect 13703 4380 14011 4389
rect 13703 4378 13709 4380
rect 13765 4378 13789 4380
rect 13845 4378 13869 4380
rect 13925 4378 13949 4380
rect 14005 4378 14011 4380
rect 13765 4326 13767 4378
rect 13947 4326 13949 4378
rect 13703 4324 13709 4326
rect 13765 4324 13789 4326
rect 13845 4324 13869 4326
rect 13925 4324 13949 4326
rect 14005 4324 14011 4326
rect 13703 4315 14011 4324
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 12728 2514 12756 3538
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 12728 1902 12756 2450
rect 12716 1896 12768 1902
rect 12716 1838 12768 1844
rect 13096 1358 13124 3538
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 13188 2650 13216 2858
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13188 1902 13216 2586
rect 13280 1970 13308 4014
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13372 3602 13400 3878
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13464 3194 13492 3334
rect 13556 3194 13584 4014
rect 14200 3516 14228 6956
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14660 6390 14688 6598
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14363 6012 14671 6021
rect 14363 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14585 6010 14609 6012
rect 14665 6010 14671 6012
rect 14425 5958 14427 6010
rect 14607 5958 14609 6010
rect 14363 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14585 5956 14609 5958
rect 14665 5956 14671 5958
rect 14363 5947 14671 5956
rect 14844 5914 14872 7942
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14363 4924 14671 4933
rect 14363 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14585 4922 14609 4924
rect 14665 4922 14671 4924
rect 14425 4870 14427 4922
rect 14607 4870 14609 4922
rect 14363 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14585 4868 14609 4870
rect 14665 4868 14671 4870
rect 14363 4859 14671 4868
rect 14752 4758 14780 4966
rect 14844 4826 14872 5646
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14476 4078 14504 4626
rect 14660 4593 14688 4626
rect 14646 4584 14702 4593
rect 14646 4519 14702 4528
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14292 3618 14320 3878
rect 14363 3836 14671 3845
rect 14363 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14585 3834 14609 3836
rect 14665 3834 14671 3836
rect 14425 3782 14427 3834
rect 14607 3782 14609 3834
rect 14363 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14585 3780 14609 3782
rect 14665 3780 14671 3782
rect 14363 3771 14671 3780
rect 14292 3590 14412 3618
rect 14200 3488 14320 3516
rect 13703 3292 14011 3301
rect 13703 3290 13709 3292
rect 13765 3290 13789 3292
rect 13845 3290 13869 3292
rect 13925 3290 13949 3292
rect 14005 3290 14011 3292
rect 13765 3238 13767 3290
rect 13947 3238 13949 3290
rect 13703 3236 13709 3238
rect 13765 3236 13789 3238
rect 13845 3236 13869 3238
rect 13925 3236 13949 3238
rect 14005 3236 14011 3238
rect 13703 3227 14011 3236
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 14292 2632 14320 3488
rect 14384 2990 14412 3590
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14363 2748 14671 2757
rect 14363 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14585 2746 14609 2748
rect 14665 2746 14671 2748
rect 14425 2694 14427 2746
rect 14607 2694 14609 2746
rect 14363 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14585 2692 14609 2694
rect 14665 2692 14671 2694
rect 14363 2683 14671 2692
rect 14292 2604 14412 2632
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13268 1964 13320 1970
rect 13268 1906 13320 1912
rect 13176 1896 13228 1902
rect 13176 1838 13228 1844
rect 13372 1494 13400 2246
rect 13464 1494 13492 2450
rect 13556 2106 13584 2450
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 13703 2204 14011 2213
rect 13703 2202 13709 2204
rect 13765 2202 13789 2204
rect 13845 2202 13869 2204
rect 13925 2202 13949 2204
rect 14005 2202 14011 2204
rect 13765 2150 13767 2202
rect 13947 2150 13949 2202
rect 13703 2148 13709 2150
rect 13765 2148 13789 2150
rect 13845 2148 13869 2150
rect 13925 2148 13949 2150
rect 14005 2148 14011 2150
rect 13703 2139 14011 2148
rect 14292 2106 14320 2246
rect 13544 2100 13596 2106
rect 13544 2042 13596 2048
rect 14280 2100 14332 2106
rect 14280 2042 14332 2048
rect 14384 1902 14412 2604
rect 14648 2508 14700 2514
rect 14752 2496 14780 3946
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 14844 3194 14872 3334
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 14936 2582 14964 11154
rect 15120 10810 15148 11154
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 15028 9178 15056 9590
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15028 8634 15056 9114
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 15028 8090 15056 8298
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 15028 7342 15056 8026
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15028 7002 15056 7278
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 15028 2990 15056 3946
rect 15120 3942 15148 10066
rect 15212 5114 15240 12174
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 11937 15424 12038
rect 15382 11928 15438 11937
rect 15382 11863 15438 11872
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15396 10985 15424 11018
rect 15382 10976 15438 10985
rect 15382 10911 15438 10920
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 9761 15424 9862
rect 15382 9752 15438 9761
rect 15382 9687 15438 9696
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15396 8673 15424 8774
rect 15382 8664 15438 8673
rect 15382 8599 15438 8608
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 15396 7585 15424 7890
rect 15382 7576 15438 7585
rect 15382 7511 15438 7520
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15304 6458 15332 6802
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15488 6497 15516 6598
rect 15474 6488 15530 6497
rect 15292 6452 15344 6458
rect 15474 6423 15530 6432
rect 15292 6394 15344 6400
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15396 5409 15424 5510
rect 15382 5400 15438 5409
rect 15382 5335 15438 5344
rect 15212 5086 15516 5114
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15212 4078 15240 4966
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15304 4321 15332 4422
rect 15290 4312 15346 4321
rect 15290 4247 15346 4256
rect 15396 4078 15424 4626
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15396 3738 15424 4014
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15304 3194 15332 3538
rect 15488 3346 15516 5086
rect 15580 4146 15608 10542
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15396 3318 15516 3346
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 15396 2774 15424 3318
rect 15474 3224 15530 3233
rect 15474 3159 15476 3168
rect 15528 3159 15530 3168
rect 15476 3130 15528 3136
rect 15120 2746 15424 2774
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 14700 2468 14780 2496
rect 14648 2450 14700 2456
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 14844 1902 14872 2246
rect 14936 2106 14964 2246
rect 14924 2100 14976 2106
rect 14924 2042 14976 2048
rect 14372 1896 14424 1902
rect 14372 1838 14424 1844
rect 14832 1896 14884 1902
rect 14832 1838 14884 1844
rect 14280 1760 14332 1766
rect 14280 1702 14332 1708
rect 13360 1488 13412 1494
rect 13360 1430 13412 1436
rect 13452 1488 13504 1494
rect 13452 1430 13504 1436
rect 13084 1352 13136 1358
rect 13084 1294 13136 1300
rect 13703 1116 14011 1125
rect 13703 1114 13709 1116
rect 13765 1114 13789 1116
rect 13845 1114 13869 1116
rect 13925 1114 13949 1116
rect 14005 1114 14011 1116
rect 13765 1062 13767 1114
rect 13947 1062 13949 1114
rect 13703 1060 13709 1062
rect 13765 1060 13789 1062
rect 13845 1060 13869 1062
rect 13925 1060 13949 1062
rect 14005 1060 14011 1062
rect 13703 1051 14011 1060
rect 14292 814 14320 1702
rect 14363 1660 14671 1669
rect 14363 1658 14369 1660
rect 14425 1658 14449 1660
rect 14505 1658 14529 1660
rect 14585 1658 14609 1660
rect 14665 1658 14671 1660
rect 14425 1606 14427 1658
rect 14607 1606 14609 1658
rect 14363 1604 14369 1606
rect 14425 1604 14449 1606
rect 14505 1604 14529 1606
rect 14585 1604 14609 1606
rect 14665 1604 14671 1606
rect 14363 1595 14671 1604
rect 14844 1562 14872 1838
rect 14832 1556 14884 1562
rect 14832 1498 14884 1504
rect 15120 1494 15148 2746
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 15212 2106 15240 2518
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 15396 2145 15424 2246
rect 15382 2136 15438 2145
rect 15200 2100 15252 2106
rect 15382 2071 15438 2080
rect 15200 2042 15252 2048
rect 15108 1488 15160 1494
rect 15108 1430 15160 1436
rect 15120 1018 15148 1430
rect 15384 1216 15436 1222
rect 15384 1158 15436 1164
rect 15396 1057 15424 1158
rect 15382 1048 15438 1057
rect 15108 1012 15160 1018
rect 15382 983 15438 992
rect 15108 954 15160 960
rect 388 808 440 814
rect 386 776 388 785
rect 1308 808 1360 814
rect 440 776 442 785
rect 1308 750 1360 756
rect 3056 808 3108 814
rect 3056 750 3108 756
rect 4988 808 5040 814
rect 4988 750 5040 756
rect 6368 808 6420 814
rect 6368 750 6420 756
rect 8668 808 8720 814
rect 8668 750 8720 756
rect 11060 808 11112 814
rect 11060 750 11112 756
rect 12624 808 12676 814
rect 12624 750 12676 756
rect 14280 808 14332 814
rect 14280 750 14332 756
rect 386 711 442 720
rect 1308 672 1360 678
rect 1308 614 1360 620
rect 3240 672 3292 678
rect 3240 614 3292 620
rect 5264 672 5316 678
rect 5264 614 5316 620
rect 7104 672 7156 678
rect 7104 614 7156 620
rect 8944 672 8996 678
rect 8944 614 8996 620
rect 10784 672 10836 678
rect 10784 614 10836 620
rect 12808 672 12860 678
rect 12808 614 12860 620
rect 14740 672 14792 678
rect 14740 614 14792 620
rect 1320 105 1348 614
rect 2564 572 2872 581
rect 2564 570 2570 572
rect 2626 570 2650 572
rect 2706 570 2730 572
rect 2786 570 2810 572
rect 2866 570 2872 572
rect 2626 518 2628 570
rect 2808 518 2810 570
rect 2564 516 2570 518
rect 2626 516 2650 518
rect 2706 516 2730 518
rect 2786 516 2810 518
rect 2866 516 2872 518
rect 2564 507 2872 516
rect 3252 105 3280 614
rect 5276 105 5304 614
rect 6497 572 6805 581
rect 6497 570 6503 572
rect 6559 570 6583 572
rect 6639 570 6663 572
rect 6719 570 6743 572
rect 6799 570 6805 572
rect 6559 518 6561 570
rect 6741 518 6743 570
rect 6497 516 6503 518
rect 6559 516 6583 518
rect 6639 516 6663 518
rect 6719 516 6743 518
rect 6799 516 6805 518
rect 6497 507 6805 516
rect 7116 105 7144 614
rect 8956 105 8984 614
rect 10430 572 10738 581
rect 10430 570 10436 572
rect 10492 570 10516 572
rect 10572 570 10596 572
rect 10652 570 10676 572
rect 10732 570 10738 572
rect 10492 518 10494 570
rect 10674 518 10676 570
rect 10430 516 10436 518
rect 10492 516 10516 518
rect 10572 516 10596 518
rect 10652 516 10676 518
rect 10732 516 10738 518
rect 10430 507 10738 516
rect 10796 377 10824 614
rect 10782 368 10838 377
rect 10782 303 10838 312
rect 12820 105 12848 614
rect 14363 572 14671 581
rect 14363 570 14369 572
rect 14425 570 14449 572
rect 14505 570 14529 572
rect 14585 570 14609 572
rect 14665 570 14671 572
rect 14425 518 14427 570
rect 14607 518 14609 570
rect 14363 516 14369 518
rect 14425 516 14449 518
rect 14505 516 14529 518
rect 14585 516 14609 518
rect 14665 516 14671 518
rect 14363 507 14671 516
rect 14752 105 14780 614
rect 1306 96 1362 105
rect 1306 31 1362 40
rect 3238 96 3294 105
rect 3238 31 3294 40
rect 5262 96 5318 105
rect 5262 31 5318 40
rect 7102 96 7158 105
rect 7102 31 7158 40
rect 8942 96 8998 105
rect 8942 31 8998 40
rect 12806 96 12862 105
rect 12806 31 12862 40
rect 14738 96 14794 105
rect 14738 31 14794 40
<< via2 >>
rect 12806 13912 12862 13968
rect 3238 13776 3294 13832
rect 5262 13776 5318 13832
rect 6642 13776 6698 13832
rect 8942 13776 8998 13832
rect 10874 13776 10930 13832
rect 1122 13232 1178 13288
rect 846 13096 902 13152
rect 1910 13082 1966 13084
rect 1990 13082 2046 13084
rect 2070 13082 2126 13084
rect 2150 13082 2206 13084
rect 1910 13030 1956 13082
rect 1956 13030 1966 13082
rect 1990 13030 2020 13082
rect 2020 13030 2032 13082
rect 2032 13030 2046 13082
rect 2070 13030 2084 13082
rect 2084 13030 2096 13082
rect 2096 13030 2126 13082
rect 2150 13030 2160 13082
rect 2160 13030 2206 13082
rect 1910 13028 1966 13030
rect 1990 13028 2046 13030
rect 2070 13028 2126 13030
rect 2150 13028 2206 13030
rect 5843 13082 5899 13084
rect 5923 13082 5979 13084
rect 6003 13082 6059 13084
rect 6083 13082 6139 13084
rect 5843 13030 5889 13082
rect 5889 13030 5899 13082
rect 5923 13030 5953 13082
rect 5953 13030 5965 13082
rect 5965 13030 5979 13082
rect 6003 13030 6017 13082
rect 6017 13030 6029 13082
rect 6029 13030 6059 13082
rect 6083 13030 6093 13082
rect 6093 13030 6139 13082
rect 5843 13028 5899 13030
rect 5923 13028 5979 13030
rect 6003 13028 6059 13030
rect 6083 13028 6139 13030
rect 9776 13082 9832 13084
rect 9856 13082 9912 13084
rect 9936 13082 9992 13084
rect 10016 13082 10072 13084
rect 9776 13030 9822 13082
rect 9822 13030 9832 13082
rect 9856 13030 9886 13082
rect 9886 13030 9898 13082
rect 9898 13030 9912 13082
rect 9936 13030 9950 13082
rect 9950 13030 9962 13082
rect 9962 13030 9992 13082
rect 10016 13030 10026 13082
rect 10026 13030 10072 13082
rect 9776 13028 9832 13030
rect 9856 13028 9912 13030
rect 9936 13028 9992 13030
rect 10016 13028 10072 13030
rect 14646 13776 14702 13832
rect 13709 13082 13765 13084
rect 13789 13082 13845 13084
rect 13869 13082 13925 13084
rect 13949 13082 14005 13084
rect 13709 13030 13755 13082
rect 13755 13030 13765 13082
rect 13789 13030 13819 13082
rect 13819 13030 13831 13082
rect 13831 13030 13845 13082
rect 13869 13030 13883 13082
rect 13883 13030 13895 13082
rect 13895 13030 13925 13082
rect 13949 13030 13959 13082
rect 13959 13030 14005 13082
rect 13709 13028 13765 13030
rect 13789 13028 13845 13030
rect 13869 13028 13925 13030
rect 13949 13028 14005 13030
rect 15474 12980 15530 13016
rect 15474 12960 15476 12980
rect 15476 12960 15528 12980
rect 15528 12960 15530 12980
rect 386 12144 442 12200
rect 478 11192 534 11248
rect 478 10240 534 10296
rect 478 9324 480 9344
rect 480 9324 532 9344
rect 532 9324 534 9344
rect 478 9288 534 9324
rect 386 8356 442 8392
rect 386 8336 388 8356
rect 388 8336 440 8356
rect 440 8336 442 8356
rect 478 7384 534 7440
rect 478 6432 534 6488
rect 2570 12538 2626 12540
rect 2650 12538 2706 12540
rect 2730 12538 2786 12540
rect 2810 12538 2866 12540
rect 2570 12486 2616 12538
rect 2616 12486 2626 12538
rect 2650 12486 2680 12538
rect 2680 12486 2692 12538
rect 2692 12486 2706 12538
rect 2730 12486 2744 12538
rect 2744 12486 2756 12538
rect 2756 12486 2786 12538
rect 2810 12486 2820 12538
rect 2820 12486 2866 12538
rect 2570 12484 2626 12486
rect 2650 12484 2706 12486
rect 2730 12484 2786 12486
rect 2810 12484 2866 12486
rect 1910 11994 1966 11996
rect 1990 11994 2046 11996
rect 2070 11994 2126 11996
rect 2150 11994 2206 11996
rect 1910 11942 1956 11994
rect 1956 11942 1966 11994
rect 1990 11942 2020 11994
rect 2020 11942 2032 11994
rect 2032 11942 2046 11994
rect 2070 11942 2084 11994
rect 2084 11942 2096 11994
rect 2096 11942 2126 11994
rect 2150 11942 2160 11994
rect 2160 11942 2206 11994
rect 1910 11940 1966 11942
rect 1990 11940 2046 11942
rect 2070 11940 2126 11942
rect 2150 11940 2206 11942
rect 2570 11450 2626 11452
rect 2650 11450 2706 11452
rect 2730 11450 2786 11452
rect 2810 11450 2866 11452
rect 2570 11398 2616 11450
rect 2616 11398 2626 11450
rect 2650 11398 2680 11450
rect 2680 11398 2692 11450
rect 2692 11398 2706 11450
rect 2730 11398 2744 11450
rect 2744 11398 2756 11450
rect 2756 11398 2786 11450
rect 2810 11398 2820 11450
rect 2820 11398 2866 11450
rect 2570 11396 2626 11398
rect 2650 11396 2706 11398
rect 2730 11396 2786 11398
rect 2810 11396 2866 11398
rect 1910 10906 1966 10908
rect 1990 10906 2046 10908
rect 2070 10906 2126 10908
rect 2150 10906 2206 10908
rect 1910 10854 1956 10906
rect 1956 10854 1966 10906
rect 1990 10854 2020 10906
rect 2020 10854 2032 10906
rect 2032 10854 2046 10906
rect 2070 10854 2084 10906
rect 2084 10854 2096 10906
rect 2096 10854 2126 10906
rect 2150 10854 2160 10906
rect 2160 10854 2206 10906
rect 1910 10852 1966 10854
rect 1990 10852 2046 10854
rect 2070 10852 2126 10854
rect 2150 10852 2206 10854
rect 2570 10362 2626 10364
rect 2650 10362 2706 10364
rect 2730 10362 2786 10364
rect 2810 10362 2866 10364
rect 2570 10310 2616 10362
rect 2616 10310 2626 10362
rect 2650 10310 2680 10362
rect 2680 10310 2692 10362
rect 2692 10310 2706 10362
rect 2730 10310 2744 10362
rect 2744 10310 2756 10362
rect 2756 10310 2786 10362
rect 2810 10310 2820 10362
rect 2820 10310 2866 10362
rect 2570 10308 2626 10310
rect 2650 10308 2706 10310
rect 2730 10308 2786 10310
rect 2810 10308 2866 10310
rect 1910 9818 1966 9820
rect 1990 9818 2046 9820
rect 2070 9818 2126 9820
rect 2150 9818 2206 9820
rect 1910 9766 1956 9818
rect 1956 9766 1966 9818
rect 1990 9766 2020 9818
rect 2020 9766 2032 9818
rect 2032 9766 2046 9818
rect 2070 9766 2084 9818
rect 2084 9766 2096 9818
rect 2096 9766 2126 9818
rect 2150 9766 2160 9818
rect 2160 9766 2206 9818
rect 1910 9764 1966 9766
rect 1990 9764 2046 9766
rect 2070 9764 2126 9766
rect 2150 9764 2206 9766
rect 2570 9274 2626 9276
rect 2650 9274 2706 9276
rect 2730 9274 2786 9276
rect 2810 9274 2866 9276
rect 2570 9222 2616 9274
rect 2616 9222 2626 9274
rect 2650 9222 2680 9274
rect 2680 9222 2692 9274
rect 2692 9222 2706 9274
rect 2730 9222 2744 9274
rect 2744 9222 2756 9274
rect 2756 9222 2786 9274
rect 2810 9222 2820 9274
rect 2820 9222 2866 9274
rect 2570 9220 2626 9222
rect 2650 9220 2706 9222
rect 2730 9220 2786 9222
rect 2810 9220 2866 9222
rect 1910 8730 1966 8732
rect 1990 8730 2046 8732
rect 2070 8730 2126 8732
rect 2150 8730 2206 8732
rect 1910 8678 1956 8730
rect 1956 8678 1966 8730
rect 1990 8678 2020 8730
rect 2020 8678 2032 8730
rect 2032 8678 2046 8730
rect 2070 8678 2084 8730
rect 2084 8678 2096 8730
rect 2096 8678 2126 8730
rect 2150 8678 2160 8730
rect 2160 8678 2206 8730
rect 1910 8676 1966 8678
rect 1990 8676 2046 8678
rect 2070 8676 2126 8678
rect 2150 8676 2206 8678
rect 2570 8186 2626 8188
rect 2650 8186 2706 8188
rect 2730 8186 2786 8188
rect 2810 8186 2866 8188
rect 2570 8134 2616 8186
rect 2616 8134 2626 8186
rect 2650 8134 2680 8186
rect 2680 8134 2692 8186
rect 2692 8134 2706 8186
rect 2730 8134 2744 8186
rect 2744 8134 2756 8186
rect 2756 8134 2786 8186
rect 2810 8134 2820 8186
rect 2820 8134 2866 8186
rect 2570 8132 2626 8134
rect 2650 8132 2706 8134
rect 2730 8132 2786 8134
rect 2810 8132 2866 8134
rect 478 5516 480 5536
rect 480 5516 532 5536
rect 532 5516 534 5536
rect 478 5480 534 5516
rect 478 4120 534 4176
rect 1122 3596 1178 3632
rect 1122 3576 1124 3596
rect 1124 3576 1176 3596
rect 1176 3576 1178 3596
rect 386 2624 442 2680
rect 1910 7642 1966 7644
rect 1990 7642 2046 7644
rect 2070 7642 2126 7644
rect 2150 7642 2206 7644
rect 1910 7590 1956 7642
rect 1956 7590 1966 7642
rect 1990 7590 2020 7642
rect 2020 7590 2032 7642
rect 2032 7590 2046 7642
rect 2070 7590 2084 7642
rect 2084 7590 2096 7642
rect 2096 7590 2126 7642
rect 2150 7590 2160 7642
rect 2160 7590 2206 7642
rect 1910 7588 1966 7590
rect 1990 7588 2046 7590
rect 2070 7588 2126 7590
rect 2150 7588 2206 7590
rect 6503 12538 6559 12540
rect 6583 12538 6639 12540
rect 6663 12538 6719 12540
rect 6743 12538 6799 12540
rect 6503 12486 6549 12538
rect 6549 12486 6559 12538
rect 6583 12486 6613 12538
rect 6613 12486 6625 12538
rect 6625 12486 6639 12538
rect 6663 12486 6677 12538
rect 6677 12486 6689 12538
rect 6689 12486 6719 12538
rect 6743 12486 6753 12538
rect 6753 12486 6799 12538
rect 6503 12484 6559 12486
rect 6583 12484 6639 12486
rect 6663 12484 6719 12486
rect 6743 12484 6799 12486
rect 2570 7098 2626 7100
rect 2650 7098 2706 7100
rect 2730 7098 2786 7100
rect 2810 7098 2866 7100
rect 2570 7046 2616 7098
rect 2616 7046 2626 7098
rect 2650 7046 2680 7098
rect 2680 7046 2692 7098
rect 2692 7046 2706 7098
rect 2730 7046 2744 7098
rect 2744 7046 2756 7098
rect 2756 7046 2786 7098
rect 2810 7046 2820 7098
rect 2820 7046 2866 7098
rect 2570 7044 2626 7046
rect 2650 7044 2706 7046
rect 2730 7044 2786 7046
rect 2810 7044 2866 7046
rect 1910 6554 1966 6556
rect 1990 6554 2046 6556
rect 2070 6554 2126 6556
rect 2150 6554 2206 6556
rect 1910 6502 1956 6554
rect 1956 6502 1966 6554
rect 1990 6502 2020 6554
rect 2020 6502 2032 6554
rect 2032 6502 2046 6554
rect 2070 6502 2084 6554
rect 2084 6502 2096 6554
rect 2096 6502 2126 6554
rect 2150 6502 2160 6554
rect 2160 6502 2206 6554
rect 1910 6500 1966 6502
rect 1990 6500 2046 6502
rect 2070 6500 2126 6502
rect 2150 6500 2206 6502
rect 2570 6010 2626 6012
rect 2650 6010 2706 6012
rect 2730 6010 2786 6012
rect 2810 6010 2866 6012
rect 2570 5958 2616 6010
rect 2616 5958 2626 6010
rect 2650 5958 2680 6010
rect 2680 5958 2692 6010
rect 2692 5958 2706 6010
rect 2730 5958 2744 6010
rect 2744 5958 2756 6010
rect 2756 5958 2786 6010
rect 2810 5958 2820 6010
rect 2820 5958 2866 6010
rect 2570 5956 2626 5958
rect 2650 5956 2706 5958
rect 2730 5956 2786 5958
rect 2810 5956 2866 5958
rect 1910 5466 1966 5468
rect 1990 5466 2046 5468
rect 2070 5466 2126 5468
rect 2150 5466 2206 5468
rect 1910 5414 1956 5466
rect 1956 5414 1966 5466
rect 1990 5414 2020 5466
rect 2020 5414 2032 5466
rect 2032 5414 2046 5466
rect 2070 5414 2084 5466
rect 2084 5414 2096 5466
rect 2096 5414 2126 5466
rect 2150 5414 2160 5466
rect 2160 5414 2206 5466
rect 1910 5412 1966 5414
rect 1990 5412 2046 5414
rect 2070 5412 2126 5414
rect 2150 5412 2206 5414
rect 2570 4922 2626 4924
rect 2650 4922 2706 4924
rect 2730 4922 2786 4924
rect 2810 4922 2866 4924
rect 2570 4870 2616 4922
rect 2616 4870 2626 4922
rect 2650 4870 2680 4922
rect 2680 4870 2692 4922
rect 2692 4870 2706 4922
rect 2730 4870 2744 4922
rect 2744 4870 2756 4922
rect 2756 4870 2786 4922
rect 2810 4870 2820 4922
rect 2820 4870 2866 4922
rect 2570 4868 2626 4870
rect 2650 4868 2706 4870
rect 2730 4868 2786 4870
rect 2810 4868 2866 4870
rect 1910 4378 1966 4380
rect 1990 4378 2046 4380
rect 2070 4378 2126 4380
rect 2150 4378 2206 4380
rect 1910 4326 1956 4378
rect 1956 4326 1966 4378
rect 1990 4326 2020 4378
rect 2020 4326 2032 4378
rect 2032 4326 2046 4378
rect 2070 4326 2084 4378
rect 2084 4326 2096 4378
rect 2096 4326 2126 4378
rect 2150 4326 2160 4378
rect 2160 4326 2206 4378
rect 1910 4324 1966 4326
rect 1990 4324 2046 4326
rect 2070 4324 2126 4326
rect 2150 4324 2206 4326
rect 1910 3290 1966 3292
rect 1990 3290 2046 3292
rect 2070 3290 2126 3292
rect 2150 3290 2206 3292
rect 1910 3238 1956 3290
rect 1956 3238 1966 3290
rect 1990 3238 2020 3290
rect 2020 3238 2032 3290
rect 2032 3238 2046 3290
rect 2070 3238 2084 3290
rect 2084 3238 2096 3290
rect 2096 3238 2126 3290
rect 2150 3238 2160 3290
rect 2160 3238 2206 3290
rect 1910 3236 1966 3238
rect 1990 3236 2046 3238
rect 2070 3236 2126 3238
rect 2150 3236 2206 3238
rect 2570 3834 2626 3836
rect 2650 3834 2706 3836
rect 2730 3834 2786 3836
rect 2810 3834 2866 3836
rect 2570 3782 2616 3834
rect 2616 3782 2626 3834
rect 2650 3782 2680 3834
rect 2680 3782 2692 3834
rect 2692 3782 2706 3834
rect 2730 3782 2744 3834
rect 2744 3782 2756 3834
rect 2756 3782 2786 3834
rect 2810 3782 2820 3834
rect 2820 3782 2866 3834
rect 2570 3780 2626 3782
rect 2650 3780 2706 3782
rect 2730 3780 2786 3782
rect 2810 3780 2866 3782
rect 3606 6196 3608 6216
rect 3608 6196 3660 6216
rect 3660 6196 3662 6216
rect 3606 6160 3662 6196
rect 4066 5480 4122 5536
rect 4618 6160 4674 6216
rect 2570 2746 2626 2748
rect 2650 2746 2706 2748
rect 2730 2746 2786 2748
rect 2810 2746 2866 2748
rect 2570 2694 2616 2746
rect 2616 2694 2626 2746
rect 2650 2694 2680 2746
rect 2680 2694 2692 2746
rect 2692 2694 2706 2746
rect 2730 2694 2744 2746
rect 2744 2694 2756 2746
rect 2756 2694 2786 2746
rect 2810 2694 2820 2746
rect 2820 2694 2866 2746
rect 2570 2692 2626 2694
rect 2650 2692 2706 2694
rect 2730 2692 2786 2694
rect 2810 2692 2866 2694
rect 1910 2202 1966 2204
rect 1990 2202 2046 2204
rect 2070 2202 2126 2204
rect 2150 2202 2206 2204
rect 1910 2150 1956 2202
rect 1956 2150 1966 2202
rect 1990 2150 2020 2202
rect 2020 2150 2032 2202
rect 2032 2150 2046 2202
rect 2070 2150 2084 2202
rect 2084 2150 2096 2202
rect 2096 2150 2126 2202
rect 2150 2150 2160 2202
rect 2160 2150 2206 2202
rect 1910 2148 1966 2150
rect 1990 2148 2046 2150
rect 2070 2148 2126 2150
rect 2150 2148 2206 2150
rect 2570 1658 2626 1660
rect 2650 1658 2706 1660
rect 2730 1658 2786 1660
rect 2810 1658 2866 1660
rect 2570 1606 2616 1658
rect 2616 1606 2626 1658
rect 2650 1606 2680 1658
rect 2680 1606 2692 1658
rect 2692 1606 2706 1658
rect 2730 1606 2744 1658
rect 2744 1606 2756 1658
rect 2756 1606 2786 1658
rect 2810 1606 2820 1658
rect 2820 1606 2866 1658
rect 2570 1604 2626 1606
rect 2650 1604 2706 1606
rect 2730 1604 2786 1606
rect 2810 1604 2866 1606
rect 1910 1114 1966 1116
rect 1990 1114 2046 1116
rect 2070 1114 2126 1116
rect 2150 1114 2206 1116
rect 1910 1062 1956 1114
rect 1956 1062 1966 1114
rect 1990 1062 2020 1114
rect 2020 1062 2032 1114
rect 2032 1062 2046 1114
rect 2070 1062 2084 1114
rect 2084 1062 2096 1114
rect 2096 1062 2126 1114
rect 2150 1062 2160 1114
rect 2160 1062 2206 1114
rect 1910 1060 1966 1062
rect 1990 1060 2046 1062
rect 2070 1060 2126 1062
rect 2150 1060 2206 1062
rect 5843 11994 5899 11996
rect 5923 11994 5979 11996
rect 6003 11994 6059 11996
rect 6083 11994 6139 11996
rect 5843 11942 5889 11994
rect 5889 11942 5899 11994
rect 5923 11942 5953 11994
rect 5953 11942 5965 11994
rect 5965 11942 5979 11994
rect 6003 11942 6017 11994
rect 6017 11942 6029 11994
rect 6029 11942 6059 11994
rect 6083 11942 6093 11994
rect 6093 11942 6139 11994
rect 5843 11940 5899 11942
rect 5923 11940 5979 11942
rect 6003 11940 6059 11942
rect 6083 11940 6139 11942
rect 5843 10906 5899 10908
rect 5923 10906 5979 10908
rect 6003 10906 6059 10908
rect 6083 10906 6139 10908
rect 5843 10854 5889 10906
rect 5889 10854 5899 10906
rect 5923 10854 5953 10906
rect 5953 10854 5965 10906
rect 5965 10854 5979 10906
rect 6003 10854 6017 10906
rect 6017 10854 6029 10906
rect 6029 10854 6059 10906
rect 6083 10854 6093 10906
rect 6093 10854 6139 10906
rect 5843 10852 5899 10854
rect 5923 10852 5979 10854
rect 6003 10852 6059 10854
rect 6083 10852 6139 10854
rect 5843 9818 5899 9820
rect 5923 9818 5979 9820
rect 6003 9818 6059 9820
rect 6083 9818 6139 9820
rect 5843 9766 5889 9818
rect 5889 9766 5899 9818
rect 5923 9766 5953 9818
rect 5953 9766 5965 9818
rect 5965 9766 5979 9818
rect 6003 9766 6017 9818
rect 6017 9766 6029 9818
rect 6029 9766 6059 9818
rect 6083 9766 6093 9818
rect 6093 9766 6139 9818
rect 5843 9764 5899 9766
rect 5923 9764 5979 9766
rect 6003 9764 6059 9766
rect 6083 9764 6139 9766
rect 5843 8730 5899 8732
rect 5923 8730 5979 8732
rect 6003 8730 6059 8732
rect 6083 8730 6139 8732
rect 5843 8678 5889 8730
rect 5889 8678 5899 8730
rect 5923 8678 5953 8730
rect 5953 8678 5965 8730
rect 5965 8678 5979 8730
rect 6003 8678 6017 8730
rect 6017 8678 6029 8730
rect 6029 8678 6059 8730
rect 6083 8678 6093 8730
rect 6093 8678 6139 8730
rect 5843 8676 5899 8678
rect 5923 8676 5979 8678
rect 6003 8676 6059 8678
rect 6083 8676 6139 8678
rect 5843 7642 5899 7644
rect 5923 7642 5979 7644
rect 6003 7642 6059 7644
rect 6083 7642 6139 7644
rect 5843 7590 5889 7642
rect 5889 7590 5899 7642
rect 5923 7590 5953 7642
rect 5953 7590 5965 7642
rect 5965 7590 5979 7642
rect 6003 7590 6017 7642
rect 6017 7590 6029 7642
rect 6029 7590 6059 7642
rect 6083 7590 6093 7642
rect 6093 7590 6139 7642
rect 5843 7588 5899 7590
rect 5923 7588 5979 7590
rect 6003 7588 6059 7590
rect 6083 7588 6139 7590
rect 5843 6554 5899 6556
rect 5923 6554 5979 6556
rect 6003 6554 6059 6556
rect 6083 6554 6139 6556
rect 5843 6502 5889 6554
rect 5889 6502 5899 6554
rect 5923 6502 5953 6554
rect 5953 6502 5965 6554
rect 5965 6502 5979 6554
rect 6003 6502 6017 6554
rect 6017 6502 6029 6554
rect 6029 6502 6059 6554
rect 6083 6502 6093 6554
rect 6093 6502 6139 6554
rect 5843 6500 5899 6502
rect 5923 6500 5979 6502
rect 6003 6500 6059 6502
rect 6083 6500 6139 6502
rect 6503 11450 6559 11452
rect 6583 11450 6639 11452
rect 6663 11450 6719 11452
rect 6743 11450 6799 11452
rect 6503 11398 6549 11450
rect 6549 11398 6559 11450
rect 6583 11398 6613 11450
rect 6613 11398 6625 11450
rect 6625 11398 6639 11450
rect 6663 11398 6677 11450
rect 6677 11398 6689 11450
rect 6689 11398 6719 11450
rect 6743 11398 6753 11450
rect 6753 11398 6799 11450
rect 6503 11396 6559 11398
rect 6583 11396 6639 11398
rect 6663 11396 6719 11398
rect 6743 11396 6799 11398
rect 10436 12538 10492 12540
rect 10516 12538 10572 12540
rect 10596 12538 10652 12540
rect 10676 12538 10732 12540
rect 10436 12486 10482 12538
rect 10482 12486 10492 12538
rect 10516 12486 10546 12538
rect 10546 12486 10558 12538
rect 10558 12486 10572 12538
rect 10596 12486 10610 12538
rect 10610 12486 10622 12538
rect 10622 12486 10652 12538
rect 10676 12486 10686 12538
rect 10686 12486 10732 12538
rect 10436 12484 10492 12486
rect 10516 12484 10572 12486
rect 10596 12484 10652 12486
rect 10676 12484 10732 12486
rect 9776 11994 9832 11996
rect 9856 11994 9912 11996
rect 9936 11994 9992 11996
rect 10016 11994 10072 11996
rect 9776 11942 9822 11994
rect 9822 11942 9832 11994
rect 9856 11942 9886 11994
rect 9886 11942 9898 11994
rect 9898 11942 9912 11994
rect 9936 11942 9950 11994
rect 9950 11942 9962 11994
rect 9962 11942 9992 11994
rect 10016 11942 10026 11994
rect 10026 11942 10072 11994
rect 9776 11940 9832 11942
rect 9856 11940 9912 11942
rect 9936 11940 9992 11942
rect 10016 11940 10072 11942
rect 6503 10362 6559 10364
rect 6583 10362 6639 10364
rect 6663 10362 6719 10364
rect 6743 10362 6799 10364
rect 6503 10310 6549 10362
rect 6549 10310 6559 10362
rect 6583 10310 6613 10362
rect 6613 10310 6625 10362
rect 6625 10310 6639 10362
rect 6663 10310 6677 10362
rect 6677 10310 6689 10362
rect 6689 10310 6719 10362
rect 6743 10310 6753 10362
rect 6753 10310 6799 10362
rect 6503 10308 6559 10310
rect 6583 10308 6639 10310
rect 6663 10308 6719 10310
rect 6743 10308 6799 10310
rect 6503 9274 6559 9276
rect 6583 9274 6639 9276
rect 6663 9274 6719 9276
rect 6743 9274 6799 9276
rect 6503 9222 6549 9274
rect 6549 9222 6559 9274
rect 6583 9222 6613 9274
rect 6613 9222 6625 9274
rect 6625 9222 6639 9274
rect 6663 9222 6677 9274
rect 6677 9222 6689 9274
rect 6689 9222 6719 9274
rect 6743 9222 6753 9274
rect 6753 9222 6799 9274
rect 6503 9220 6559 9222
rect 6583 9220 6639 9222
rect 6663 9220 6719 9222
rect 6743 9220 6799 9222
rect 6503 8186 6559 8188
rect 6583 8186 6639 8188
rect 6663 8186 6719 8188
rect 6743 8186 6799 8188
rect 6503 8134 6549 8186
rect 6549 8134 6559 8186
rect 6583 8134 6613 8186
rect 6613 8134 6625 8186
rect 6625 8134 6639 8186
rect 6663 8134 6677 8186
rect 6677 8134 6689 8186
rect 6689 8134 6719 8186
rect 6743 8134 6753 8186
rect 6753 8134 6799 8186
rect 6503 8132 6559 8134
rect 6583 8132 6639 8134
rect 6663 8132 6719 8134
rect 6743 8132 6799 8134
rect 6182 6180 6238 6216
rect 6182 6160 6184 6180
rect 6184 6160 6236 6180
rect 6236 6160 6238 6180
rect 5538 5480 5594 5536
rect 5843 5466 5899 5468
rect 5923 5466 5979 5468
rect 6003 5466 6059 5468
rect 6083 5466 6139 5468
rect 5843 5414 5889 5466
rect 5889 5414 5899 5466
rect 5923 5414 5953 5466
rect 5953 5414 5965 5466
rect 5965 5414 5979 5466
rect 6003 5414 6017 5466
rect 6017 5414 6029 5466
rect 6029 5414 6059 5466
rect 6083 5414 6093 5466
rect 6093 5414 6139 5466
rect 5843 5412 5899 5414
rect 5923 5412 5979 5414
rect 6003 5412 6059 5414
rect 6083 5412 6139 5414
rect 5814 4684 5870 4720
rect 5814 4664 5816 4684
rect 5816 4664 5868 4684
rect 5868 4664 5870 4684
rect 5843 4378 5899 4380
rect 5923 4378 5979 4380
rect 6003 4378 6059 4380
rect 6083 4378 6139 4380
rect 5843 4326 5889 4378
rect 5889 4326 5899 4378
rect 5923 4326 5953 4378
rect 5953 4326 5965 4378
rect 5965 4326 5979 4378
rect 6003 4326 6017 4378
rect 6017 4326 6029 4378
rect 6029 4326 6059 4378
rect 6083 4326 6093 4378
rect 6093 4326 6139 4378
rect 5843 4324 5899 4326
rect 5923 4324 5979 4326
rect 6003 4324 6059 4326
rect 6083 4324 6139 4326
rect 5843 3290 5899 3292
rect 5923 3290 5979 3292
rect 6003 3290 6059 3292
rect 6083 3290 6139 3292
rect 5843 3238 5889 3290
rect 5889 3238 5899 3290
rect 5923 3238 5953 3290
rect 5953 3238 5965 3290
rect 5965 3238 5979 3290
rect 6003 3238 6017 3290
rect 6017 3238 6029 3290
rect 6029 3238 6059 3290
rect 6083 3238 6093 3290
rect 6093 3238 6139 3290
rect 5843 3236 5899 3238
rect 5923 3236 5979 3238
rect 6003 3236 6059 3238
rect 6083 3236 6139 3238
rect 4066 1808 4122 1864
rect 5843 2202 5899 2204
rect 5923 2202 5979 2204
rect 6003 2202 6059 2204
rect 6083 2202 6139 2204
rect 5843 2150 5889 2202
rect 5889 2150 5899 2202
rect 5923 2150 5953 2202
rect 5953 2150 5965 2202
rect 5965 2150 5979 2202
rect 6003 2150 6017 2202
rect 6017 2150 6029 2202
rect 6029 2150 6059 2202
rect 6083 2150 6093 2202
rect 6093 2150 6139 2202
rect 5843 2148 5899 2150
rect 5923 2148 5979 2150
rect 6003 2148 6059 2150
rect 6083 2148 6139 2150
rect 5843 1114 5899 1116
rect 5923 1114 5979 1116
rect 6003 1114 6059 1116
rect 6083 1114 6139 1116
rect 5843 1062 5889 1114
rect 5889 1062 5899 1114
rect 5923 1062 5953 1114
rect 5953 1062 5965 1114
rect 5965 1062 5979 1114
rect 6003 1062 6017 1114
rect 6017 1062 6029 1114
rect 6029 1062 6059 1114
rect 6083 1062 6093 1114
rect 6093 1062 6139 1114
rect 5843 1060 5899 1062
rect 5923 1060 5979 1062
rect 6003 1060 6059 1062
rect 6083 1060 6139 1062
rect 6503 7098 6559 7100
rect 6583 7098 6639 7100
rect 6663 7098 6719 7100
rect 6743 7098 6799 7100
rect 6503 7046 6549 7098
rect 6549 7046 6559 7098
rect 6583 7046 6613 7098
rect 6613 7046 6625 7098
rect 6625 7046 6639 7098
rect 6663 7046 6677 7098
rect 6677 7046 6689 7098
rect 6689 7046 6719 7098
rect 6743 7046 6753 7098
rect 6753 7046 6799 7098
rect 6503 7044 6559 7046
rect 6583 7044 6639 7046
rect 6663 7044 6719 7046
rect 6743 7044 6799 7046
rect 6503 6010 6559 6012
rect 6583 6010 6639 6012
rect 6663 6010 6719 6012
rect 6743 6010 6799 6012
rect 6503 5958 6549 6010
rect 6549 5958 6559 6010
rect 6583 5958 6613 6010
rect 6613 5958 6625 6010
rect 6625 5958 6639 6010
rect 6663 5958 6677 6010
rect 6677 5958 6689 6010
rect 6689 5958 6719 6010
rect 6743 5958 6753 6010
rect 6753 5958 6799 6010
rect 6503 5956 6559 5958
rect 6583 5956 6639 5958
rect 6663 5956 6719 5958
rect 6743 5956 6799 5958
rect 6503 4922 6559 4924
rect 6583 4922 6639 4924
rect 6663 4922 6719 4924
rect 6743 4922 6799 4924
rect 6503 4870 6549 4922
rect 6549 4870 6559 4922
rect 6583 4870 6613 4922
rect 6613 4870 6625 4922
rect 6625 4870 6639 4922
rect 6663 4870 6677 4922
rect 6677 4870 6689 4922
rect 6689 4870 6719 4922
rect 6743 4870 6753 4922
rect 6753 4870 6799 4922
rect 6503 4868 6559 4870
rect 6583 4868 6639 4870
rect 6663 4868 6719 4870
rect 6743 4868 6799 4870
rect 6503 3834 6559 3836
rect 6583 3834 6639 3836
rect 6663 3834 6719 3836
rect 6743 3834 6799 3836
rect 6503 3782 6549 3834
rect 6549 3782 6559 3834
rect 6583 3782 6613 3834
rect 6613 3782 6625 3834
rect 6625 3782 6639 3834
rect 6663 3782 6677 3834
rect 6677 3782 6689 3834
rect 6689 3782 6719 3834
rect 6743 3782 6753 3834
rect 6753 3782 6799 3834
rect 6503 3780 6559 3782
rect 6583 3780 6639 3782
rect 6663 3780 6719 3782
rect 6743 3780 6799 3782
rect 6503 2746 6559 2748
rect 6583 2746 6639 2748
rect 6663 2746 6719 2748
rect 6743 2746 6799 2748
rect 6503 2694 6549 2746
rect 6549 2694 6559 2746
rect 6583 2694 6613 2746
rect 6613 2694 6625 2746
rect 6625 2694 6639 2746
rect 6663 2694 6677 2746
rect 6677 2694 6689 2746
rect 6689 2694 6719 2746
rect 6743 2694 6753 2746
rect 6753 2694 6799 2746
rect 6503 2692 6559 2694
rect 6583 2692 6639 2694
rect 6663 2692 6719 2694
rect 6743 2692 6799 2694
rect 6503 1658 6559 1660
rect 6583 1658 6639 1660
rect 6663 1658 6719 1660
rect 6743 1658 6799 1660
rect 6503 1606 6549 1658
rect 6549 1606 6559 1658
rect 6583 1606 6613 1658
rect 6613 1606 6625 1658
rect 6625 1606 6639 1658
rect 6663 1606 6677 1658
rect 6677 1606 6689 1658
rect 6689 1606 6719 1658
rect 6743 1606 6753 1658
rect 6753 1606 6799 1658
rect 6503 1604 6559 1606
rect 6583 1604 6639 1606
rect 6663 1604 6719 1606
rect 6743 1604 6799 1606
rect 10436 11450 10492 11452
rect 10516 11450 10572 11452
rect 10596 11450 10652 11452
rect 10676 11450 10732 11452
rect 10436 11398 10482 11450
rect 10482 11398 10492 11450
rect 10516 11398 10546 11450
rect 10546 11398 10558 11450
rect 10558 11398 10572 11450
rect 10596 11398 10610 11450
rect 10610 11398 10622 11450
rect 10622 11398 10652 11450
rect 10676 11398 10686 11450
rect 10686 11398 10732 11450
rect 10436 11396 10492 11398
rect 10516 11396 10572 11398
rect 10596 11396 10652 11398
rect 10676 11396 10732 11398
rect 9776 10906 9832 10908
rect 9856 10906 9912 10908
rect 9936 10906 9992 10908
rect 10016 10906 10072 10908
rect 9776 10854 9822 10906
rect 9822 10854 9832 10906
rect 9856 10854 9886 10906
rect 9886 10854 9898 10906
rect 9898 10854 9912 10906
rect 9936 10854 9950 10906
rect 9950 10854 9962 10906
rect 9962 10854 9992 10906
rect 10016 10854 10026 10906
rect 10026 10854 10072 10906
rect 9776 10852 9832 10854
rect 9856 10852 9912 10854
rect 9936 10852 9992 10854
rect 10016 10852 10072 10854
rect 13709 11994 13765 11996
rect 13789 11994 13845 11996
rect 13869 11994 13925 11996
rect 13949 11994 14005 11996
rect 13709 11942 13755 11994
rect 13755 11942 13765 11994
rect 13789 11942 13819 11994
rect 13819 11942 13831 11994
rect 13831 11942 13845 11994
rect 13869 11942 13883 11994
rect 13883 11942 13895 11994
rect 13895 11942 13925 11994
rect 13949 11942 13959 11994
rect 13959 11942 14005 11994
rect 13709 11940 13765 11942
rect 13789 11940 13845 11942
rect 13869 11940 13925 11942
rect 13949 11940 14005 11942
rect 13709 10906 13765 10908
rect 13789 10906 13845 10908
rect 13869 10906 13925 10908
rect 13949 10906 14005 10908
rect 13709 10854 13755 10906
rect 13755 10854 13765 10906
rect 13789 10854 13819 10906
rect 13819 10854 13831 10906
rect 13831 10854 13845 10906
rect 13869 10854 13883 10906
rect 13883 10854 13895 10906
rect 13895 10854 13925 10906
rect 13949 10854 13959 10906
rect 13959 10854 14005 10906
rect 13709 10852 13765 10854
rect 13789 10852 13845 10854
rect 13869 10852 13925 10854
rect 13949 10852 14005 10854
rect 10436 10362 10492 10364
rect 10516 10362 10572 10364
rect 10596 10362 10652 10364
rect 10676 10362 10732 10364
rect 10436 10310 10482 10362
rect 10482 10310 10492 10362
rect 10516 10310 10546 10362
rect 10546 10310 10558 10362
rect 10558 10310 10572 10362
rect 10596 10310 10610 10362
rect 10610 10310 10622 10362
rect 10622 10310 10652 10362
rect 10676 10310 10686 10362
rect 10686 10310 10732 10362
rect 10436 10308 10492 10310
rect 10516 10308 10572 10310
rect 10596 10308 10652 10310
rect 10676 10308 10732 10310
rect 9776 9818 9832 9820
rect 9856 9818 9912 9820
rect 9936 9818 9992 9820
rect 10016 9818 10072 9820
rect 9776 9766 9822 9818
rect 9822 9766 9832 9818
rect 9856 9766 9886 9818
rect 9886 9766 9898 9818
rect 9898 9766 9912 9818
rect 9936 9766 9950 9818
rect 9950 9766 9962 9818
rect 9962 9766 9992 9818
rect 10016 9766 10026 9818
rect 10026 9766 10072 9818
rect 9776 9764 9832 9766
rect 9856 9764 9912 9766
rect 9936 9764 9992 9766
rect 10016 9764 10072 9766
rect 9776 8730 9832 8732
rect 9856 8730 9912 8732
rect 9936 8730 9992 8732
rect 10016 8730 10072 8732
rect 9776 8678 9822 8730
rect 9822 8678 9832 8730
rect 9856 8678 9886 8730
rect 9886 8678 9898 8730
rect 9898 8678 9912 8730
rect 9936 8678 9950 8730
rect 9950 8678 9962 8730
rect 9962 8678 9992 8730
rect 10016 8678 10026 8730
rect 10026 8678 10072 8730
rect 9776 8676 9832 8678
rect 9856 8676 9912 8678
rect 9936 8676 9992 8678
rect 10016 8676 10072 8678
rect 10436 9274 10492 9276
rect 10516 9274 10572 9276
rect 10596 9274 10652 9276
rect 10676 9274 10732 9276
rect 10436 9222 10482 9274
rect 10482 9222 10492 9274
rect 10516 9222 10546 9274
rect 10546 9222 10558 9274
rect 10558 9222 10572 9274
rect 10596 9222 10610 9274
rect 10610 9222 10622 9274
rect 10622 9222 10652 9274
rect 10676 9222 10686 9274
rect 10686 9222 10732 9274
rect 10436 9220 10492 9222
rect 10516 9220 10572 9222
rect 10596 9220 10652 9222
rect 10676 9220 10732 9222
rect 10436 8186 10492 8188
rect 10516 8186 10572 8188
rect 10596 8186 10652 8188
rect 10676 8186 10732 8188
rect 10436 8134 10482 8186
rect 10482 8134 10492 8186
rect 10516 8134 10546 8186
rect 10546 8134 10558 8186
rect 10558 8134 10572 8186
rect 10596 8134 10610 8186
rect 10610 8134 10622 8186
rect 10622 8134 10652 8186
rect 10676 8134 10686 8186
rect 10686 8134 10732 8186
rect 10436 8132 10492 8134
rect 10516 8132 10572 8134
rect 10596 8132 10652 8134
rect 10676 8132 10732 8134
rect 9776 7642 9832 7644
rect 9856 7642 9912 7644
rect 9936 7642 9992 7644
rect 10016 7642 10072 7644
rect 9776 7590 9822 7642
rect 9822 7590 9832 7642
rect 9856 7590 9886 7642
rect 9886 7590 9898 7642
rect 9898 7590 9912 7642
rect 9936 7590 9950 7642
rect 9950 7590 9962 7642
rect 9962 7590 9992 7642
rect 10016 7590 10026 7642
rect 10026 7590 10072 7642
rect 9776 7588 9832 7590
rect 9856 7588 9912 7590
rect 9936 7588 9992 7590
rect 10016 7588 10072 7590
rect 10436 7098 10492 7100
rect 10516 7098 10572 7100
rect 10596 7098 10652 7100
rect 10676 7098 10732 7100
rect 10436 7046 10482 7098
rect 10482 7046 10492 7098
rect 10516 7046 10546 7098
rect 10546 7046 10558 7098
rect 10558 7046 10572 7098
rect 10596 7046 10610 7098
rect 10610 7046 10622 7098
rect 10622 7046 10652 7098
rect 10676 7046 10686 7098
rect 10686 7046 10732 7098
rect 10436 7044 10492 7046
rect 10516 7044 10572 7046
rect 10596 7044 10652 7046
rect 10676 7044 10732 7046
rect 9776 6554 9832 6556
rect 9856 6554 9912 6556
rect 9936 6554 9992 6556
rect 10016 6554 10072 6556
rect 9776 6502 9822 6554
rect 9822 6502 9832 6554
rect 9856 6502 9886 6554
rect 9886 6502 9898 6554
rect 9898 6502 9912 6554
rect 9936 6502 9950 6554
rect 9950 6502 9962 6554
rect 9962 6502 9992 6554
rect 10016 6502 10026 6554
rect 10026 6502 10072 6554
rect 9776 6500 9832 6502
rect 9856 6500 9912 6502
rect 9936 6500 9992 6502
rect 10016 6500 10072 6502
rect 10436 6010 10492 6012
rect 10516 6010 10572 6012
rect 10596 6010 10652 6012
rect 10676 6010 10732 6012
rect 10436 5958 10482 6010
rect 10482 5958 10492 6010
rect 10516 5958 10546 6010
rect 10546 5958 10558 6010
rect 10558 5958 10572 6010
rect 10596 5958 10610 6010
rect 10610 5958 10622 6010
rect 10622 5958 10652 6010
rect 10676 5958 10686 6010
rect 10686 5958 10732 6010
rect 10436 5956 10492 5958
rect 10516 5956 10572 5958
rect 10596 5956 10652 5958
rect 10676 5956 10732 5958
rect 10874 5888 10930 5944
rect 9776 5466 9832 5468
rect 9856 5466 9912 5468
rect 9936 5466 9992 5468
rect 10016 5466 10072 5468
rect 9776 5414 9822 5466
rect 9822 5414 9832 5466
rect 9856 5414 9886 5466
rect 9886 5414 9898 5466
rect 9898 5414 9912 5466
rect 9936 5414 9950 5466
rect 9950 5414 9962 5466
rect 9962 5414 9992 5466
rect 10016 5414 10026 5466
rect 10026 5414 10072 5466
rect 9776 5412 9832 5414
rect 9856 5412 9912 5414
rect 9936 5412 9992 5414
rect 10016 5412 10072 5414
rect 13709 9818 13765 9820
rect 13789 9818 13845 9820
rect 13869 9818 13925 9820
rect 13949 9818 14005 9820
rect 13709 9766 13755 9818
rect 13755 9766 13765 9818
rect 13789 9766 13819 9818
rect 13819 9766 13831 9818
rect 13831 9766 13845 9818
rect 13869 9766 13883 9818
rect 13883 9766 13895 9818
rect 13895 9766 13925 9818
rect 13949 9766 13959 9818
rect 13959 9766 14005 9818
rect 13709 9764 13765 9766
rect 13789 9764 13845 9766
rect 13869 9764 13925 9766
rect 13949 9764 14005 9766
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14609 12538 14665 12540
rect 14369 12486 14415 12538
rect 14415 12486 14425 12538
rect 14449 12486 14479 12538
rect 14479 12486 14491 12538
rect 14491 12486 14505 12538
rect 14529 12486 14543 12538
rect 14543 12486 14555 12538
rect 14555 12486 14585 12538
rect 14609 12486 14619 12538
rect 14619 12486 14665 12538
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 14609 12484 14665 12486
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14609 11450 14665 11452
rect 14369 11398 14415 11450
rect 14415 11398 14425 11450
rect 14449 11398 14479 11450
rect 14479 11398 14491 11450
rect 14491 11398 14505 11450
rect 14529 11398 14543 11450
rect 14543 11398 14555 11450
rect 14555 11398 14585 11450
rect 14609 11398 14619 11450
rect 14619 11398 14665 11450
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 14609 11396 14665 11398
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14609 10362 14665 10364
rect 14369 10310 14415 10362
rect 14415 10310 14425 10362
rect 14449 10310 14479 10362
rect 14479 10310 14491 10362
rect 14491 10310 14505 10362
rect 14529 10310 14543 10362
rect 14543 10310 14555 10362
rect 14555 10310 14585 10362
rect 14609 10310 14619 10362
rect 14619 10310 14665 10362
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 14609 10308 14665 10310
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14609 9274 14665 9276
rect 14369 9222 14415 9274
rect 14415 9222 14425 9274
rect 14449 9222 14479 9274
rect 14479 9222 14491 9274
rect 14491 9222 14505 9274
rect 14529 9222 14543 9274
rect 14543 9222 14555 9274
rect 14555 9222 14585 9274
rect 14609 9222 14619 9274
rect 14619 9222 14665 9274
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 14609 9220 14665 9222
rect 13709 8730 13765 8732
rect 13789 8730 13845 8732
rect 13869 8730 13925 8732
rect 13949 8730 14005 8732
rect 13709 8678 13755 8730
rect 13755 8678 13765 8730
rect 13789 8678 13819 8730
rect 13819 8678 13831 8730
rect 13831 8678 13845 8730
rect 13869 8678 13883 8730
rect 13883 8678 13895 8730
rect 13895 8678 13925 8730
rect 13949 8678 13959 8730
rect 13959 8678 14005 8730
rect 13709 8676 13765 8678
rect 13789 8676 13845 8678
rect 13869 8676 13925 8678
rect 13949 8676 14005 8678
rect 13709 7642 13765 7644
rect 13789 7642 13845 7644
rect 13869 7642 13925 7644
rect 13949 7642 14005 7644
rect 13709 7590 13755 7642
rect 13755 7590 13765 7642
rect 13789 7590 13819 7642
rect 13819 7590 13831 7642
rect 13831 7590 13845 7642
rect 13869 7590 13883 7642
rect 13883 7590 13895 7642
rect 13895 7590 13925 7642
rect 13949 7590 13959 7642
rect 13959 7590 14005 7642
rect 13709 7588 13765 7590
rect 13789 7588 13845 7590
rect 13869 7588 13925 7590
rect 13949 7588 14005 7590
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14609 8186 14665 8188
rect 14369 8134 14415 8186
rect 14415 8134 14425 8186
rect 14449 8134 14479 8186
rect 14479 8134 14491 8186
rect 14491 8134 14505 8186
rect 14529 8134 14543 8186
rect 14543 8134 14555 8186
rect 14555 8134 14585 8186
rect 14609 8134 14619 8186
rect 14619 8134 14665 8186
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 14609 8132 14665 8134
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14609 7098 14665 7100
rect 14369 7046 14415 7098
rect 14415 7046 14425 7098
rect 14449 7046 14479 7098
rect 14479 7046 14491 7098
rect 14491 7046 14505 7098
rect 14529 7046 14543 7098
rect 14543 7046 14555 7098
rect 14555 7046 14585 7098
rect 14609 7046 14619 7098
rect 14619 7046 14665 7098
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14609 7044 14665 7046
rect 9586 4684 9642 4720
rect 9586 4664 9588 4684
rect 9588 4664 9640 4684
rect 9640 4664 9642 4684
rect 9776 4378 9832 4380
rect 9856 4378 9912 4380
rect 9936 4378 9992 4380
rect 10016 4378 10072 4380
rect 9776 4326 9822 4378
rect 9822 4326 9832 4378
rect 9856 4326 9886 4378
rect 9886 4326 9898 4378
rect 9898 4326 9912 4378
rect 9936 4326 9950 4378
rect 9950 4326 9962 4378
rect 9962 4326 9992 4378
rect 10016 4326 10026 4378
rect 10026 4326 10072 4378
rect 9776 4324 9832 4326
rect 9856 4324 9912 4326
rect 9936 4324 9992 4326
rect 10016 4324 10072 4326
rect 10436 4922 10492 4924
rect 10516 4922 10572 4924
rect 10596 4922 10652 4924
rect 10676 4922 10732 4924
rect 10436 4870 10482 4922
rect 10482 4870 10492 4922
rect 10516 4870 10546 4922
rect 10546 4870 10558 4922
rect 10558 4870 10572 4922
rect 10596 4870 10610 4922
rect 10610 4870 10622 4922
rect 10622 4870 10652 4922
rect 10676 4870 10686 4922
rect 10686 4870 10732 4922
rect 10436 4868 10492 4870
rect 10516 4868 10572 4870
rect 10596 4868 10652 4870
rect 10676 4868 10732 4870
rect 10506 4528 10562 4584
rect 10874 4020 10876 4040
rect 10876 4020 10928 4040
rect 10928 4020 10930 4040
rect 10874 3984 10930 4020
rect 10436 3834 10492 3836
rect 10516 3834 10572 3836
rect 10596 3834 10652 3836
rect 10676 3834 10732 3836
rect 10436 3782 10482 3834
rect 10482 3782 10492 3834
rect 10516 3782 10546 3834
rect 10546 3782 10558 3834
rect 10558 3782 10572 3834
rect 10596 3782 10610 3834
rect 10610 3782 10622 3834
rect 10622 3782 10652 3834
rect 10676 3782 10686 3834
rect 10686 3782 10732 3834
rect 10436 3780 10492 3782
rect 10516 3780 10572 3782
rect 10596 3780 10652 3782
rect 10676 3780 10732 3782
rect 9776 3290 9832 3292
rect 9856 3290 9912 3292
rect 9936 3290 9992 3292
rect 10016 3290 10072 3292
rect 9776 3238 9822 3290
rect 9822 3238 9832 3290
rect 9856 3238 9886 3290
rect 9886 3238 9898 3290
rect 9898 3238 9912 3290
rect 9936 3238 9950 3290
rect 9950 3238 9962 3290
rect 9962 3238 9992 3290
rect 10016 3238 10026 3290
rect 10026 3238 10072 3290
rect 9776 3236 9832 3238
rect 9856 3236 9912 3238
rect 9936 3236 9992 3238
rect 10016 3236 10072 3238
rect 10436 2746 10492 2748
rect 10516 2746 10572 2748
rect 10596 2746 10652 2748
rect 10676 2746 10732 2748
rect 10436 2694 10482 2746
rect 10482 2694 10492 2746
rect 10516 2694 10546 2746
rect 10546 2694 10558 2746
rect 10558 2694 10572 2746
rect 10596 2694 10610 2746
rect 10610 2694 10622 2746
rect 10622 2694 10652 2746
rect 10676 2694 10686 2746
rect 10686 2694 10732 2746
rect 10436 2692 10492 2694
rect 10516 2692 10572 2694
rect 10596 2692 10652 2694
rect 10676 2692 10732 2694
rect 9776 2202 9832 2204
rect 9856 2202 9912 2204
rect 9936 2202 9992 2204
rect 10016 2202 10072 2204
rect 9776 2150 9822 2202
rect 9822 2150 9832 2202
rect 9856 2150 9886 2202
rect 9886 2150 9898 2202
rect 9898 2150 9912 2202
rect 9936 2150 9950 2202
rect 9950 2150 9962 2202
rect 9962 2150 9992 2202
rect 10016 2150 10026 2202
rect 10026 2150 10072 2202
rect 9776 2148 9832 2150
rect 9856 2148 9912 2150
rect 9936 2148 9992 2150
rect 10016 2148 10072 2150
rect 10436 1658 10492 1660
rect 10516 1658 10572 1660
rect 10596 1658 10652 1660
rect 10676 1658 10732 1660
rect 10436 1606 10482 1658
rect 10482 1606 10492 1658
rect 10516 1606 10546 1658
rect 10546 1606 10558 1658
rect 10558 1606 10572 1658
rect 10596 1606 10610 1658
rect 10610 1606 10622 1658
rect 10622 1606 10652 1658
rect 10676 1606 10686 1658
rect 10686 1606 10732 1658
rect 10436 1604 10492 1606
rect 10516 1604 10572 1606
rect 10596 1604 10652 1606
rect 10676 1604 10732 1606
rect 11242 3984 11298 4040
rect 9776 1114 9832 1116
rect 9856 1114 9912 1116
rect 9936 1114 9992 1116
rect 10016 1114 10072 1116
rect 9776 1062 9822 1114
rect 9822 1062 9832 1114
rect 9856 1062 9886 1114
rect 9886 1062 9898 1114
rect 9898 1062 9912 1114
rect 9936 1062 9950 1114
rect 9950 1062 9962 1114
rect 9962 1062 9992 1114
rect 10016 1062 10026 1114
rect 10026 1062 10072 1114
rect 9776 1060 9832 1062
rect 9856 1060 9912 1062
rect 9936 1060 9992 1062
rect 10016 1060 10072 1062
rect 13709 6554 13765 6556
rect 13789 6554 13845 6556
rect 13869 6554 13925 6556
rect 13949 6554 14005 6556
rect 13709 6502 13755 6554
rect 13755 6502 13765 6554
rect 13789 6502 13819 6554
rect 13819 6502 13831 6554
rect 13831 6502 13845 6554
rect 13869 6502 13883 6554
rect 13883 6502 13895 6554
rect 13895 6502 13925 6554
rect 13949 6502 13959 6554
rect 13959 6502 14005 6554
rect 13709 6500 13765 6502
rect 13789 6500 13845 6502
rect 13869 6500 13925 6502
rect 13949 6500 14005 6502
rect 13726 5888 13782 5944
rect 13709 5466 13765 5468
rect 13789 5466 13845 5468
rect 13869 5466 13925 5468
rect 13949 5466 14005 5468
rect 13709 5414 13755 5466
rect 13755 5414 13765 5466
rect 13789 5414 13819 5466
rect 13819 5414 13831 5466
rect 13831 5414 13845 5466
rect 13869 5414 13883 5466
rect 13883 5414 13895 5466
rect 13895 5414 13925 5466
rect 13949 5414 13959 5466
rect 13959 5414 14005 5466
rect 13709 5412 13765 5414
rect 13789 5412 13845 5414
rect 13869 5412 13925 5414
rect 13949 5412 14005 5414
rect 13709 4378 13765 4380
rect 13789 4378 13845 4380
rect 13869 4378 13925 4380
rect 13949 4378 14005 4380
rect 13709 4326 13755 4378
rect 13755 4326 13765 4378
rect 13789 4326 13819 4378
rect 13819 4326 13831 4378
rect 13831 4326 13845 4378
rect 13869 4326 13883 4378
rect 13883 4326 13895 4378
rect 13895 4326 13925 4378
rect 13949 4326 13959 4378
rect 13959 4326 14005 4378
rect 13709 4324 13765 4326
rect 13789 4324 13845 4326
rect 13869 4324 13925 4326
rect 13949 4324 14005 4326
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14609 6010 14665 6012
rect 14369 5958 14415 6010
rect 14415 5958 14425 6010
rect 14449 5958 14479 6010
rect 14479 5958 14491 6010
rect 14491 5958 14505 6010
rect 14529 5958 14543 6010
rect 14543 5958 14555 6010
rect 14555 5958 14585 6010
rect 14609 5958 14619 6010
rect 14619 5958 14665 6010
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 14609 5956 14665 5958
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14609 4922 14665 4924
rect 14369 4870 14415 4922
rect 14415 4870 14425 4922
rect 14449 4870 14479 4922
rect 14479 4870 14491 4922
rect 14491 4870 14505 4922
rect 14529 4870 14543 4922
rect 14543 4870 14555 4922
rect 14555 4870 14585 4922
rect 14609 4870 14619 4922
rect 14619 4870 14665 4922
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 14609 4868 14665 4870
rect 14646 4528 14702 4584
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14609 3834 14665 3836
rect 14369 3782 14415 3834
rect 14415 3782 14425 3834
rect 14449 3782 14479 3834
rect 14479 3782 14491 3834
rect 14491 3782 14505 3834
rect 14529 3782 14543 3834
rect 14543 3782 14555 3834
rect 14555 3782 14585 3834
rect 14609 3782 14619 3834
rect 14619 3782 14665 3834
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 14609 3780 14665 3782
rect 13709 3290 13765 3292
rect 13789 3290 13845 3292
rect 13869 3290 13925 3292
rect 13949 3290 14005 3292
rect 13709 3238 13755 3290
rect 13755 3238 13765 3290
rect 13789 3238 13819 3290
rect 13819 3238 13831 3290
rect 13831 3238 13845 3290
rect 13869 3238 13883 3290
rect 13883 3238 13895 3290
rect 13895 3238 13925 3290
rect 13949 3238 13959 3290
rect 13959 3238 14005 3290
rect 13709 3236 13765 3238
rect 13789 3236 13845 3238
rect 13869 3236 13925 3238
rect 13949 3236 14005 3238
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14609 2746 14665 2748
rect 14369 2694 14415 2746
rect 14415 2694 14425 2746
rect 14449 2694 14479 2746
rect 14479 2694 14491 2746
rect 14491 2694 14505 2746
rect 14529 2694 14543 2746
rect 14543 2694 14555 2746
rect 14555 2694 14585 2746
rect 14609 2694 14619 2746
rect 14619 2694 14665 2746
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 14609 2692 14665 2694
rect 13709 2202 13765 2204
rect 13789 2202 13845 2204
rect 13869 2202 13925 2204
rect 13949 2202 14005 2204
rect 13709 2150 13755 2202
rect 13755 2150 13765 2202
rect 13789 2150 13819 2202
rect 13819 2150 13831 2202
rect 13831 2150 13845 2202
rect 13869 2150 13883 2202
rect 13883 2150 13895 2202
rect 13895 2150 13925 2202
rect 13949 2150 13959 2202
rect 13959 2150 14005 2202
rect 13709 2148 13765 2150
rect 13789 2148 13845 2150
rect 13869 2148 13925 2150
rect 13949 2148 14005 2150
rect 15382 11872 15438 11928
rect 15382 10920 15438 10976
rect 15382 9696 15438 9752
rect 15382 8608 15438 8664
rect 15382 7520 15438 7576
rect 15474 6432 15530 6488
rect 15382 5344 15438 5400
rect 15290 4256 15346 4312
rect 15474 3188 15530 3224
rect 15474 3168 15476 3188
rect 15476 3168 15528 3188
rect 15528 3168 15530 3188
rect 13709 1114 13765 1116
rect 13789 1114 13845 1116
rect 13869 1114 13925 1116
rect 13949 1114 14005 1116
rect 13709 1062 13755 1114
rect 13755 1062 13765 1114
rect 13789 1062 13819 1114
rect 13819 1062 13831 1114
rect 13831 1062 13845 1114
rect 13869 1062 13883 1114
rect 13883 1062 13895 1114
rect 13895 1062 13925 1114
rect 13949 1062 13959 1114
rect 13959 1062 14005 1114
rect 13709 1060 13765 1062
rect 13789 1060 13845 1062
rect 13869 1060 13925 1062
rect 13949 1060 14005 1062
rect 14369 1658 14425 1660
rect 14449 1658 14505 1660
rect 14529 1658 14585 1660
rect 14609 1658 14665 1660
rect 14369 1606 14415 1658
rect 14415 1606 14425 1658
rect 14449 1606 14479 1658
rect 14479 1606 14491 1658
rect 14491 1606 14505 1658
rect 14529 1606 14543 1658
rect 14543 1606 14555 1658
rect 14555 1606 14585 1658
rect 14609 1606 14619 1658
rect 14619 1606 14665 1658
rect 14369 1604 14425 1606
rect 14449 1604 14505 1606
rect 14529 1604 14585 1606
rect 14609 1604 14665 1606
rect 15382 2080 15438 2136
rect 15382 992 15438 1048
rect 386 756 388 776
rect 388 756 440 776
rect 440 756 442 776
rect 386 720 442 756
rect 2570 570 2626 572
rect 2650 570 2706 572
rect 2730 570 2786 572
rect 2810 570 2866 572
rect 2570 518 2616 570
rect 2616 518 2626 570
rect 2650 518 2680 570
rect 2680 518 2692 570
rect 2692 518 2706 570
rect 2730 518 2744 570
rect 2744 518 2756 570
rect 2756 518 2786 570
rect 2810 518 2820 570
rect 2820 518 2866 570
rect 2570 516 2626 518
rect 2650 516 2706 518
rect 2730 516 2786 518
rect 2810 516 2866 518
rect 6503 570 6559 572
rect 6583 570 6639 572
rect 6663 570 6719 572
rect 6743 570 6799 572
rect 6503 518 6549 570
rect 6549 518 6559 570
rect 6583 518 6613 570
rect 6613 518 6625 570
rect 6625 518 6639 570
rect 6663 518 6677 570
rect 6677 518 6689 570
rect 6689 518 6719 570
rect 6743 518 6753 570
rect 6753 518 6799 570
rect 6503 516 6559 518
rect 6583 516 6639 518
rect 6663 516 6719 518
rect 6743 516 6799 518
rect 10436 570 10492 572
rect 10516 570 10572 572
rect 10596 570 10652 572
rect 10676 570 10732 572
rect 10436 518 10482 570
rect 10482 518 10492 570
rect 10516 518 10546 570
rect 10546 518 10558 570
rect 10558 518 10572 570
rect 10596 518 10610 570
rect 10610 518 10622 570
rect 10622 518 10652 570
rect 10676 518 10686 570
rect 10686 518 10732 570
rect 10436 516 10492 518
rect 10516 516 10572 518
rect 10596 516 10652 518
rect 10676 516 10732 518
rect 10782 312 10838 368
rect 14369 570 14425 572
rect 14449 570 14505 572
rect 14529 570 14585 572
rect 14609 570 14665 572
rect 14369 518 14415 570
rect 14415 518 14425 570
rect 14449 518 14479 570
rect 14479 518 14491 570
rect 14491 518 14505 570
rect 14529 518 14543 570
rect 14543 518 14555 570
rect 14555 518 14585 570
rect 14609 518 14619 570
rect 14619 518 14665 570
rect 14369 516 14425 518
rect 14449 516 14505 518
rect 14529 516 14585 518
rect 14609 516 14665 518
rect 1306 40 1362 96
rect 3238 40 3294 96
rect 5262 40 5318 96
rect 7102 40 7158 96
rect 8942 40 8998 96
rect 12806 40 12862 96
rect 14738 40 14794 96
<< metal3 >>
rect 1096 13834 1216 14000
rect 982 13800 1216 13834
rect 3000 13834 3120 14000
rect 3233 13834 3299 13837
rect 3000 13832 3299 13834
rect 3000 13800 3238 13832
rect 982 13774 1156 13800
rect 3036 13776 3238 13800
rect 3294 13776 3299 13832
rect 4904 13834 5024 14000
rect 5257 13834 5323 13837
rect 4904 13832 5323 13834
rect 4904 13800 5262 13832
rect 3036 13774 3299 13776
rect 4968 13776 5262 13800
rect 5318 13776 5323 13832
rect 4968 13774 5323 13776
rect 982 13698 1042 13774
rect 3233 13771 3299 13774
rect 5257 13771 5323 13774
rect 6637 13834 6703 13837
rect 6808 13834 6928 14000
rect 6637 13832 6928 13834
rect 6637 13776 6642 13832
rect 6698 13800 6928 13832
rect 8712 13834 8832 14000
rect 8937 13834 9003 13837
rect 8712 13832 9003 13834
rect 8712 13800 8942 13832
rect 6698 13776 6868 13800
rect 6637 13774 6868 13776
rect 8772 13776 8942 13800
rect 8998 13776 9003 13832
rect 10616 13834 10736 14000
rect 12520 13970 12640 14000
rect 12801 13970 12867 13973
rect 12520 13968 12867 13970
rect 12520 13912 12806 13968
rect 12862 13912 12867 13968
rect 12520 13910 12867 13912
rect 10869 13834 10935 13837
rect 10616 13832 10935 13834
rect 10616 13800 10874 13832
rect 8772 13774 9003 13776
rect 10672 13776 10874 13800
rect 10930 13776 10935 13832
rect 12520 13800 12640 13910
rect 12801 13907 12867 13910
rect 14424 13834 14544 14000
rect 14641 13834 14707 13837
rect 14424 13832 14707 13834
rect 14424 13800 14646 13832
rect 10672 13774 10935 13776
rect 14484 13776 14646 13800
rect 14702 13776 14707 13832
rect 14484 13774 14707 13776
rect 6637 13771 6703 13774
rect 8937 13771 9003 13774
rect 10869 13771 10935 13774
rect 14641 13771 14707 13774
rect 982 13638 1186 13698
rect 1126 13293 1186 13638
rect 1117 13288 1186 13293
rect 1117 13232 1122 13288
rect 1178 13232 1186 13288
rect 1117 13230 1186 13232
rect 1117 13227 1183 13230
rect 841 13154 907 13157
rect 0 13152 907 13154
rect 0 13096 846 13152
rect 902 13096 907 13152
rect 0 13094 907 13096
rect 841 13091 907 13094
rect 1900 13088 2216 13089
rect 1900 13024 1906 13088
rect 1970 13024 1986 13088
rect 2050 13024 2066 13088
rect 2130 13024 2146 13088
rect 2210 13024 2216 13088
rect 1900 13023 2216 13024
rect 5833 13088 6149 13089
rect 5833 13024 5839 13088
rect 5903 13024 5919 13088
rect 5983 13024 5999 13088
rect 6063 13024 6079 13088
rect 6143 13024 6149 13088
rect 5833 13023 6149 13024
rect 9766 13088 10082 13089
rect 9766 13024 9772 13088
rect 9836 13024 9852 13088
rect 9916 13024 9932 13088
rect 9996 13024 10012 13088
rect 10076 13024 10082 13088
rect 9766 13023 10082 13024
rect 13699 13088 14015 13089
rect 13699 13024 13705 13088
rect 13769 13024 13785 13088
rect 13849 13024 13865 13088
rect 13929 13024 13945 13088
rect 14009 13024 14015 13088
rect 13699 13023 14015 13024
rect 15469 13018 15535 13021
rect 15469 13016 16000 13018
rect 15469 12960 15474 13016
rect 15530 12960 16000 13016
rect 15469 12958 16000 12960
rect 15469 12955 15535 12958
rect 2560 12544 2876 12545
rect 2560 12480 2566 12544
rect 2630 12480 2646 12544
rect 2710 12480 2726 12544
rect 2790 12480 2806 12544
rect 2870 12480 2876 12544
rect 2560 12479 2876 12480
rect 6493 12544 6809 12545
rect 6493 12480 6499 12544
rect 6563 12480 6579 12544
rect 6643 12480 6659 12544
rect 6723 12480 6739 12544
rect 6803 12480 6809 12544
rect 6493 12479 6809 12480
rect 10426 12544 10742 12545
rect 10426 12480 10432 12544
rect 10496 12480 10512 12544
rect 10576 12480 10592 12544
rect 10656 12480 10672 12544
rect 10736 12480 10742 12544
rect 10426 12479 10742 12480
rect 14359 12544 14675 12545
rect 14359 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14605 12544
rect 14669 12480 14675 12544
rect 14359 12479 14675 12480
rect 381 12202 447 12205
rect 0 12200 447 12202
rect 0 12144 386 12200
rect 442 12144 447 12200
rect 0 12142 447 12144
rect 381 12139 447 12142
rect 1900 12000 2216 12001
rect 1900 11936 1906 12000
rect 1970 11936 1986 12000
rect 2050 11936 2066 12000
rect 2130 11936 2146 12000
rect 2210 11936 2216 12000
rect 1900 11935 2216 11936
rect 5833 12000 6149 12001
rect 5833 11936 5839 12000
rect 5903 11936 5919 12000
rect 5983 11936 5999 12000
rect 6063 11936 6079 12000
rect 6143 11936 6149 12000
rect 5833 11935 6149 11936
rect 9766 12000 10082 12001
rect 9766 11936 9772 12000
rect 9836 11936 9852 12000
rect 9916 11936 9932 12000
rect 9996 11936 10012 12000
rect 10076 11936 10082 12000
rect 9766 11935 10082 11936
rect 13699 12000 14015 12001
rect 13699 11936 13705 12000
rect 13769 11936 13785 12000
rect 13849 11936 13865 12000
rect 13929 11936 13945 12000
rect 14009 11936 14015 12000
rect 13699 11935 14015 11936
rect 15377 11930 15443 11933
rect 15377 11928 16000 11930
rect 15377 11872 15382 11928
rect 15438 11872 16000 11928
rect 15377 11870 16000 11872
rect 15377 11867 15443 11870
rect 2560 11456 2876 11457
rect 2560 11392 2566 11456
rect 2630 11392 2646 11456
rect 2710 11392 2726 11456
rect 2790 11392 2806 11456
rect 2870 11392 2876 11456
rect 2560 11391 2876 11392
rect 6493 11456 6809 11457
rect 6493 11392 6499 11456
rect 6563 11392 6579 11456
rect 6643 11392 6659 11456
rect 6723 11392 6739 11456
rect 6803 11392 6809 11456
rect 6493 11391 6809 11392
rect 10426 11456 10742 11457
rect 10426 11392 10432 11456
rect 10496 11392 10512 11456
rect 10576 11392 10592 11456
rect 10656 11392 10672 11456
rect 10736 11392 10742 11456
rect 10426 11391 10742 11392
rect 14359 11456 14675 11457
rect 14359 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14605 11456
rect 14669 11392 14675 11456
rect 14359 11391 14675 11392
rect 473 11250 539 11253
rect 0 11248 539 11250
rect 0 11192 478 11248
rect 534 11192 539 11248
rect 0 11190 539 11192
rect 473 11187 539 11190
rect 15377 10978 15443 10981
rect 15377 10976 15578 10978
rect 15377 10920 15382 10976
rect 15438 10920 15578 10976
rect 15377 10918 15578 10920
rect 15377 10915 15443 10918
rect 1900 10912 2216 10913
rect 1900 10848 1906 10912
rect 1970 10848 1986 10912
rect 2050 10848 2066 10912
rect 2130 10848 2146 10912
rect 2210 10848 2216 10912
rect 1900 10847 2216 10848
rect 5833 10912 6149 10913
rect 5833 10848 5839 10912
rect 5903 10848 5919 10912
rect 5983 10848 5999 10912
rect 6063 10848 6079 10912
rect 6143 10848 6149 10912
rect 5833 10847 6149 10848
rect 9766 10912 10082 10913
rect 9766 10848 9772 10912
rect 9836 10848 9852 10912
rect 9916 10848 9932 10912
rect 9996 10848 10012 10912
rect 10076 10848 10082 10912
rect 9766 10847 10082 10848
rect 13699 10912 14015 10913
rect 13699 10848 13705 10912
rect 13769 10848 13785 10912
rect 13849 10848 13865 10912
rect 13929 10848 13945 10912
rect 14009 10848 14015 10912
rect 13699 10847 14015 10848
rect 15518 10842 15578 10918
rect 15518 10782 16000 10842
rect 2560 10368 2876 10369
rect 2560 10304 2566 10368
rect 2630 10304 2646 10368
rect 2710 10304 2726 10368
rect 2790 10304 2806 10368
rect 2870 10304 2876 10368
rect 2560 10303 2876 10304
rect 6493 10368 6809 10369
rect 6493 10304 6499 10368
rect 6563 10304 6579 10368
rect 6643 10304 6659 10368
rect 6723 10304 6739 10368
rect 6803 10304 6809 10368
rect 6493 10303 6809 10304
rect 10426 10368 10742 10369
rect 10426 10304 10432 10368
rect 10496 10304 10512 10368
rect 10576 10304 10592 10368
rect 10656 10304 10672 10368
rect 10736 10304 10742 10368
rect 10426 10303 10742 10304
rect 14359 10368 14675 10369
rect 14359 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14605 10368
rect 14669 10304 14675 10368
rect 14359 10303 14675 10304
rect 473 10298 539 10301
rect 0 10296 539 10298
rect 0 10240 478 10296
rect 534 10240 539 10296
rect 0 10238 539 10240
rect 473 10235 539 10238
rect 1900 9824 2216 9825
rect 1900 9760 1906 9824
rect 1970 9760 1986 9824
rect 2050 9760 2066 9824
rect 2130 9760 2146 9824
rect 2210 9760 2216 9824
rect 1900 9759 2216 9760
rect 5833 9824 6149 9825
rect 5833 9760 5839 9824
rect 5903 9760 5919 9824
rect 5983 9760 5999 9824
rect 6063 9760 6079 9824
rect 6143 9760 6149 9824
rect 5833 9759 6149 9760
rect 9766 9824 10082 9825
rect 9766 9760 9772 9824
rect 9836 9760 9852 9824
rect 9916 9760 9932 9824
rect 9996 9760 10012 9824
rect 10076 9760 10082 9824
rect 9766 9759 10082 9760
rect 13699 9824 14015 9825
rect 13699 9760 13705 9824
rect 13769 9760 13785 9824
rect 13849 9760 13865 9824
rect 13929 9760 13945 9824
rect 14009 9760 14015 9824
rect 13699 9759 14015 9760
rect 15377 9754 15443 9757
rect 15377 9752 16000 9754
rect 15377 9696 15382 9752
rect 15438 9696 16000 9752
rect 15377 9694 16000 9696
rect 15377 9691 15443 9694
rect 473 9346 539 9349
rect 0 9344 539 9346
rect 0 9288 478 9344
rect 534 9288 539 9344
rect 0 9286 539 9288
rect 473 9283 539 9286
rect 2560 9280 2876 9281
rect 2560 9216 2566 9280
rect 2630 9216 2646 9280
rect 2710 9216 2726 9280
rect 2790 9216 2806 9280
rect 2870 9216 2876 9280
rect 2560 9215 2876 9216
rect 6493 9280 6809 9281
rect 6493 9216 6499 9280
rect 6563 9216 6579 9280
rect 6643 9216 6659 9280
rect 6723 9216 6739 9280
rect 6803 9216 6809 9280
rect 6493 9215 6809 9216
rect 10426 9280 10742 9281
rect 10426 9216 10432 9280
rect 10496 9216 10512 9280
rect 10576 9216 10592 9280
rect 10656 9216 10672 9280
rect 10736 9216 10742 9280
rect 10426 9215 10742 9216
rect 14359 9280 14675 9281
rect 14359 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14605 9280
rect 14669 9216 14675 9280
rect 14359 9215 14675 9216
rect 1900 8736 2216 8737
rect 1900 8672 1906 8736
rect 1970 8672 1986 8736
rect 2050 8672 2066 8736
rect 2130 8672 2146 8736
rect 2210 8672 2216 8736
rect 1900 8671 2216 8672
rect 5833 8736 6149 8737
rect 5833 8672 5839 8736
rect 5903 8672 5919 8736
rect 5983 8672 5999 8736
rect 6063 8672 6079 8736
rect 6143 8672 6149 8736
rect 5833 8671 6149 8672
rect 9766 8736 10082 8737
rect 9766 8672 9772 8736
rect 9836 8672 9852 8736
rect 9916 8672 9932 8736
rect 9996 8672 10012 8736
rect 10076 8672 10082 8736
rect 9766 8671 10082 8672
rect 13699 8736 14015 8737
rect 13699 8672 13705 8736
rect 13769 8672 13785 8736
rect 13849 8672 13865 8736
rect 13929 8672 13945 8736
rect 14009 8672 14015 8736
rect 13699 8671 14015 8672
rect 15377 8666 15443 8669
rect 15377 8664 16000 8666
rect 15377 8608 15382 8664
rect 15438 8608 16000 8664
rect 15377 8606 16000 8608
rect 15377 8603 15443 8606
rect 381 8394 447 8397
rect 0 8392 447 8394
rect 0 8336 386 8392
rect 442 8336 447 8392
rect 0 8334 447 8336
rect 381 8331 447 8334
rect 2560 8192 2876 8193
rect 2560 8128 2566 8192
rect 2630 8128 2646 8192
rect 2710 8128 2726 8192
rect 2790 8128 2806 8192
rect 2870 8128 2876 8192
rect 2560 8127 2876 8128
rect 6493 8192 6809 8193
rect 6493 8128 6499 8192
rect 6563 8128 6579 8192
rect 6643 8128 6659 8192
rect 6723 8128 6739 8192
rect 6803 8128 6809 8192
rect 6493 8127 6809 8128
rect 10426 8192 10742 8193
rect 10426 8128 10432 8192
rect 10496 8128 10512 8192
rect 10576 8128 10592 8192
rect 10656 8128 10672 8192
rect 10736 8128 10742 8192
rect 10426 8127 10742 8128
rect 14359 8192 14675 8193
rect 14359 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14605 8192
rect 14669 8128 14675 8192
rect 14359 8127 14675 8128
rect 1900 7648 2216 7649
rect 1900 7584 1906 7648
rect 1970 7584 1986 7648
rect 2050 7584 2066 7648
rect 2130 7584 2146 7648
rect 2210 7584 2216 7648
rect 1900 7583 2216 7584
rect 5833 7648 6149 7649
rect 5833 7584 5839 7648
rect 5903 7584 5919 7648
rect 5983 7584 5999 7648
rect 6063 7584 6079 7648
rect 6143 7584 6149 7648
rect 5833 7583 6149 7584
rect 9766 7648 10082 7649
rect 9766 7584 9772 7648
rect 9836 7584 9852 7648
rect 9916 7584 9932 7648
rect 9996 7584 10012 7648
rect 10076 7584 10082 7648
rect 9766 7583 10082 7584
rect 13699 7648 14015 7649
rect 13699 7584 13705 7648
rect 13769 7584 13785 7648
rect 13849 7584 13865 7648
rect 13929 7584 13945 7648
rect 14009 7584 14015 7648
rect 13699 7583 14015 7584
rect 15377 7578 15443 7581
rect 15377 7576 16000 7578
rect 15377 7520 15382 7576
rect 15438 7520 16000 7576
rect 15377 7518 16000 7520
rect 15377 7515 15443 7518
rect 473 7442 539 7445
rect 0 7440 539 7442
rect 0 7384 478 7440
rect 534 7384 539 7440
rect 0 7382 539 7384
rect 473 7379 539 7382
rect 2560 7104 2876 7105
rect 2560 7040 2566 7104
rect 2630 7040 2646 7104
rect 2710 7040 2726 7104
rect 2790 7040 2806 7104
rect 2870 7040 2876 7104
rect 2560 7039 2876 7040
rect 6493 7104 6809 7105
rect 6493 7040 6499 7104
rect 6563 7040 6579 7104
rect 6643 7040 6659 7104
rect 6723 7040 6739 7104
rect 6803 7040 6809 7104
rect 6493 7039 6809 7040
rect 10426 7104 10742 7105
rect 10426 7040 10432 7104
rect 10496 7040 10512 7104
rect 10576 7040 10592 7104
rect 10656 7040 10672 7104
rect 10736 7040 10742 7104
rect 10426 7039 10742 7040
rect 14359 7104 14675 7105
rect 14359 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14605 7104
rect 14669 7040 14675 7104
rect 14359 7039 14675 7040
rect 1900 6560 2216 6561
rect 1900 6496 1906 6560
rect 1970 6496 1986 6560
rect 2050 6496 2066 6560
rect 2130 6496 2146 6560
rect 2210 6496 2216 6560
rect 1900 6495 2216 6496
rect 5833 6560 6149 6561
rect 5833 6496 5839 6560
rect 5903 6496 5919 6560
rect 5983 6496 5999 6560
rect 6063 6496 6079 6560
rect 6143 6496 6149 6560
rect 5833 6495 6149 6496
rect 9766 6560 10082 6561
rect 9766 6496 9772 6560
rect 9836 6496 9852 6560
rect 9916 6496 9932 6560
rect 9996 6496 10012 6560
rect 10076 6496 10082 6560
rect 9766 6495 10082 6496
rect 13699 6560 14015 6561
rect 13699 6496 13705 6560
rect 13769 6496 13785 6560
rect 13849 6496 13865 6560
rect 13929 6496 13945 6560
rect 14009 6496 14015 6560
rect 13699 6495 14015 6496
rect 473 6490 539 6493
rect 0 6488 539 6490
rect 0 6432 478 6488
rect 534 6432 539 6488
rect 0 6430 539 6432
rect 473 6427 539 6430
rect 15469 6490 15535 6493
rect 15469 6488 16000 6490
rect 15469 6432 15474 6488
rect 15530 6432 16000 6488
rect 15469 6430 16000 6432
rect 15469 6427 15535 6430
rect 3601 6218 3667 6221
rect 4613 6218 4679 6221
rect 6177 6218 6243 6221
rect 3601 6216 6243 6218
rect 3601 6160 3606 6216
rect 3662 6160 4618 6216
rect 4674 6160 6182 6216
rect 6238 6160 6243 6216
rect 3601 6158 6243 6160
rect 3601 6155 3667 6158
rect 4613 6155 4679 6158
rect 6177 6155 6243 6158
rect 2560 6016 2876 6017
rect 2560 5952 2566 6016
rect 2630 5952 2646 6016
rect 2710 5952 2726 6016
rect 2790 5952 2806 6016
rect 2870 5952 2876 6016
rect 2560 5951 2876 5952
rect 6493 6016 6809 6017
rect 6493 5952 6499 6016
rect 6563 5952 6579 6016
rect 6643 5952 6659 6016
rect 6723 5952 6739 6016
rect 6803 5952 6809 6016
rect 6493 5951 6809 5952
rect 10426 6016 10742 6017
rect 10426 5952 10432 6016
rect 10496 5952 10512 6016
rect 10576 5952 10592 6016
rect 10656 5952 10672 6016
rect 10736 5952 10742 6016
rect 10426 5951 10742 5952
rect 14359 6016 14675 6017
rect 14359 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14605 6016
rect 14669 5952 14675 6016
rect 14359 5951 14675 5952
rect 10869 5946 10935 5949
rect 13721 5946 13787 5949
rect 10869 5944 13787 5946
rect 10869 5888 10874 5944
rect 10930 5888 13726 5944
rect 13782 5888 13787 5944
rect 10869 5886 13787 5888
rect 10869 5883 10935 5886
rect 13721 5883 13787 5886
rect 473 5538 539 5541
rect 0 5536 539 5538
rect 0 5480 478 5536
rect 534 5480 539 5536
rect 0 5478 539 5480
rect 473 5475 539 5478
rect 4061 5538 4127 5541
rect 5533 5538 5599 5541
rect 4061 5536 5599 5538
rect 4061 5480 4066 5536
rect 4122 5480 5538 5536
rect 5594 5480 5599 5536
rect 4061 5478 5599 5480
rect 4061 5475 4127 5478
rect 5533 5475 5599 5478
rect 1900 5472 2216 5473
rect 1900 5408 1906 5472
rect 1970 5408 1986 5472
rect 2050 5408 2066 5472
rect 2130 5408 2146 5472
rect 2210 5408 2216 5472
rect 1900 5407 2216 5408
rect 5833 5472 6149 5473
rect 5833 5408 5839 5472
rect 5903 5408 5919 5472
rect 5983 5408 5999 5472
rect 6063 5408 6079 5472
rect 6143 5408 6149 5472
rect 5833 5407 6149 5408
rect 9766 5472 10082 5473
rect 9766 5408 9772 5472
rect 9836 5408 9852 5472
rect 9916 5408 9932 5472
rect 9996 5408 10012 5472
rect 10076 5408 10082 5472
rect 9766 5407 10082 5408
rect 13699 5472 14015 5473
rect 13699 5408 13705 5472
rect 13769 5408 13785 5472
rect 13849 5408 13865 5472
rect 13929 5408 13945 5472
rect 14009 5408 14015 5472
rect 13699 5407 14015 5408
rect 15377 5402 15443 5405
rect 15377 5400 16000 5402
rect 15377 5344 15382 5400
rect 15438 5344 16000 5400
rect 15377 5342 16000 5344
rect 15377 5339 15443 5342
rect 2560 4928 2876 4929
rect 2560 4864 2566 4928
rect 2630 4864 2646 4928
rect 2710 4864 2726 4928
rect 2790 4864 2806 4928
rect 2870 4864 2876 4928
rect 2560 4863 2876 4864
rect 6493 4928 6809 4929
rect 6493 4864 6499 4928
rect 6563 4864 6579 4928
rect 6643 4864 6659 4928
rect 6723 4864 6739 4928
rect 6803 4864 6809 4928
rect 6493 4863 6809 4864
rect 10426 4928 10742 4929
rect 10426 4864 10432 4928
rect 10496 4864 10512 4928
rect 10576 4864 10592 4928
rect 10656 4864 10672 4928
rect 10736 4864 10742 4928
rect 10426 4863 10742 4864
rect 14359 4928 14675 4929
rect 14359 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14605 4928
rect 14669 4864 14675 4928
rect 14359 4863 14675 4864
rect 5809 4722 5875 4725
rect 9581 4722 9647 4725
rect 5809 4720 9647 4722
rect 5809 4664 5814 4720
rect 5870 4664 9586 4720
rect 9642 4664 9647 4720
rect 5809 4662 9647 4664
rect 5809 4659 5875 4662
rect 9581 4659 9647 4662
rect 10501 4586 10567 4589
rect 14641 4586 14707 4589
rect 0 4526 306 4586
rect 246 4450 306 4526
rect 10501 4584 14707 4586
rect 10501 4528 10506 4584
rect 10562 4528 14646 4584
rect 14702 4528 14707 4584
rect 10501 4526 14707 4528
rect 10501 4523 10567 4526
rect 14641 4523 14707 4526
rect 62 4390 306 4450
rect 62 4178 122 4390
rect 1900 4384 2216 4385
rect 1900 4320 1906 4384
rect 1970 4320 1986 4384
rect 2050 4320 2066 4384
rect 2130 4320 2146 4384
rect 2210 4320 2216 4384
rect 1900 4319 2216 4320
rect 5833 4384 6149 4385
rect 5833 4320 5839 4384
rect 5903 4320 5919 4384
rect 5983 4320 5999 4384
rect 6063 4320 6079 4384
rect 6143 4320 6149 4384
rect 5833 4319 6149 4320
rect 9766 4384 10082 4385
rect 9766 4320 9772 4384
rect 9836 4320 9852 4384
rect 9916 4320 9932 4384
rect 9996 4320 10012 4384
rect 10076 4320 10082 4384
rect 9766 4319 10082 4320
rect 13699 4384 14015 4385
rect 13699 4320 13705 4384
rect 13769 4320 13785 4384
rect 13849 4320 13865 4384
rect 13929 4320 13945 4384
rect 14009 4320 14015 4384
rect 13699 4319 14015 4320
rect 15285 4314 15351 4317
rect 15285 4312 16000 4314
rect 15285 4256 15290 4312
rect 15346 4256 16000 4312
rect 15285 4254 16000 4256
rect 15285 4251 15351 4254
rect 473 4178 539 4181
rect 62 4176 539 4178
rect 62 4120 478 4176
rect 534 4120 539 4176
rect 62 4118 539 4120
rect 473 4115 539 4118
rect 10869 4042 10935 4045
rect 11237 4042 11303 4045
rect 10869 4040 11303 4042
rect 10869 3984 10874 4040
rect 10930 3984 11242 4040
rect 11298 3984 11303 4040
rect 10869 3982 11303 3984
rect 10869 3979 10935 3982
rect 11237 3979 11303 3982
rect 2560 3840 2876 3841
rect 2560 3776 2566 3840
rect 2630 3776 2646 3840
rect 2710 3776 2726 3840
rect 2790 3776 2806 3840
rect 2870 3776 2876 3840
rect 2560 3775 2876 3776
rect 6493 3840 6809 3841
rect 6493 3776 6499 3840
rect 6563 3776 6579 3840
rect 6643 3776 6659 3840
rect 6723 3776 6739 3840
rect 6803 3776 6809 3840
rect 6493 3775 6809 3776
rect 10426 3840 10742 3841
rect 10426 3776 10432 3840
rect 10496 3776 10512 3840
rect 10576 3776 10592 3840
rect 10656 3776 10672 3840
rect 10736 3776 10742 3840
rect 10426 3775 10742 3776
rect 14359 3840 14675 3841
rect 14359 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14605 3840
rect 14669 3776 14675 3840
rect 14359 3775 14675 3776
rect 1117 3634 1183 3637
rect 0 3632 1183 3634
rect 0 3576 1122 3632
rect 1178 3576 1183 3632
rect 0 3574 1183 3576
rect 1117 3571 1183 3574
rect 1900 3296 2216 3297
rect 1900 3232 1906 3296
rect 1970 3232 1986 3296
rect 2050 3232 2066 3296
rect 2130 3232 2146 3296
rect 2210 3232 2216 3296
rect 1900 3231 2216 3232
rect 5833 3296 6149 3297
rect 5833 3232 5839 3296
rect 5903 3232 5919 3296
rect 5983 3232 5999 3296
rect 6063 3232 6079 3296
rect 6143 3232 6149 3296
rect 5833 3231 6149 3232
rect 9766 3296 10082 3297
rect 9766 3232 9772 3296
rect 9836 3232 9852 3296
rect 9916 3232 9932 3296
rect 9996 3232 10012 3296
rect 10076 3232 10082 3296
rect 9766 3231 10082 3232
rect 13699 3296 14015 3297
rect 13699 3232 13705 3296
rect 13769 3232 13785 3296
rect 13849 3232 13865 3296
rect 13929 3232 13945 3296
rect 14009 3232 14015 3296
rect 13699 3231 14015 3232
rect 15469 3226 15535 3229
rect 15469 3224 16000 3226
rect 15469 3168 15474 3224
rect 15530 3168 16000 3224
rect 15469 3166 16000 3168
rect 15469 3163 15535 3166
rect 2560 2752 2876 2753
rect 2560 2688 2566 2752
rect 2630 2688 2646 2752
rect 2710 2688 2726 2752
rect 2790 2688 2806 2752
rect 2870 2688 2876 2752
rect 2560 2687 2876 2688
rect 6493 2752 6809 2753
rect 6493 2688 6499 2752
rect 6563 2688 6579 2752
rect 6643 2688 6659 2752
rect 6723 2688 6739 2752
rect 6803 2688 6809 2752
rect 6493 2687 6809 2688
rect 10426 2752 10742 2753
rect 10426 2688 10432 2752
rect 10496 2688 10512 2752
rect 10576 2688 10592 2752
rect 10656 2688 10672 2752
rect 10736 2688 10742 2752
rect 10426 2687 10742 2688
rect 14359 2752 14675 2753
rect 14359 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14605 2752
rect 14669 2688 14675 2752
rect 14359 2687 14675 2688
rect 381 2682 447 2685
rect 0 2680 447 2682
rect 0 2624 386 2680
rect 442 2624 447 2680
rect 0 2622 447 2624
rect 381 2619 447 2622
rect 1900 2208 2216 2209
rect 1900 2144 1906 2208
rect 1970 2144 1986 2208
rect 2050 2144 2066 2208
rect 2130 2144 2146 2208
rect 2210 2144 2216 2208
rect 1900 2143 2216 2144
rect 5833 2208 6149 2209
rect 5833 2144 5839 2208
rect 5903 2144 5919 2208
rect 5983 2144 5999 2208
rect 6063 2144 6079 2208
rect 6143 2144 6149 2208
rect 5833 2143 6149 2144
rect 9766 2208 10082 2209
rect 9766 2144 9772 2208
rect 9836 2144 9852 2208
rect 9916 2144 9932 2208
rect 9996 2144 10012 2208
rect 10076 2144 10082 2208
rect 9766 2143 10082 2144
rect 13699 2208 14015 2209
rect 13699 2144 13705 2208
rect 13769 2144 13785 2208
rect 13849 2144 13865 2208
rect 13929 2144 13945 2208
rect 14009 2144 14015 2208
rect 13699 2143 14015 2144
rect 15377 2138 15443 2141
rect 15377 2136 16000 2138
rect 15377 2080 15382 2136
rect 15438 2080 16000 2136
rect 15377 2078 16000 2080
rect 15377 2075 15443 2078
rect 4061 1866 4127 1869
rect 2270 1864 4127 1866
rect 2270 1808 4066 1864
rect 4122 1808 4127 1864
rect 2270 1806 4127 1808
rect 2270 1730 2330 1806
rect 4061 1803 4127 1806
rect 0 1670 2330 1730
rect 2560 1664 2876 1665
rect 2560 1600 2566 1664
rect 2630 1600 2646 1664
rect 2710 1600 2726 1664
rect 2790 1600 2806 1664
rect 2870 1600 2876 1664
rect 2560 1599 2876 1600
rect 6493 1664 6809 1665
rect 6493 1600 6499 1664
rect 6563 1600 6579 1664
rect 6643 1600 6659 1664
rect 6723 1600 6739 1664
rect 6803 1600 6809 1664
rect 6493 1599 6809 1600
rect 10426 1664 10742 1665
rect 10426 1600 10432 1664
rect 10496 1600 10512 1664
rect 10576 1600 10592 1664
rect 10656 1600 10672 1664
rect 10736 1600 10742 1664
rect 10426 1599 10742 1600
rect 14359 1664 14675 1665
rect 14359 1600 14365 1664
rect 14429 1600 14445 1664
rect 14509 1600 14525 1664
rect 14589 1600 14605 1664
rect 14669 1600 14675 1664
rect 14359 1599 14675 1600
rect 1900 1120 2216 1121
rect 1900 1056 1906 1120
rect 1970 1056 1986 1120
rect 2050 1056 2066 1120
rect 2130 1056 2146 1120
rect 2210 1056 2216 1120
rect 1900 1055 2216 1056
rect 5833 1120 6149 1121
rect 5833 1056 5839 1120
rect 5903 1056 5919 1120
rect 5983 1056 5999 1120
rect 6063 1056 6079 1120
rect 6143 1056 6149 1120
rect 5833 1055 6149 1056
rect 9766 1120 10082 1121
rect 9766 1056 9772 1120
rect 9836 1056 9852 1120
rect 9916 1056 9932 1120
rect 9996 1056 10012 1120
rect 10076 1056 10082 1120
rect 9766 1055 10082 1056
rect 13699 1120 14015 1121
rect 13699 1056 13705 1120
rect 13769 1056 13785 1120
rect 13849 1056 13865 1120
rect 13929 1056 13945 1120
rect 14009 1056 14015 1120
rect 13699 1055 14015 1056
rect 15377 1050 15443 1053
rect 15377 1048 16000 1050
rect 15377 992 15382 1048
rect 15438 992 16000 1048
rect 15377 990 16000 992
rect 15377 987 15443 990
rect 381 778 447 781
rect 0 776 447 778
rect 0 720 386 776
rect 442 720 447 776
rect 0 718 447 720
rect 381 715 447 718
rect 2560 576 2876 577
rect 2560 512 2566 576
rect 2630 512 2646 576
rect 2710 512 2726 576
rect 2790 512 2806 576
rect 2870 512 2876 576
rect 2560 511 2876 512
rect 6493 576 6809 577
rect 6493 512 6499 576
rect 6563 512 6579 576
rect 6643 512 6659 576
rect 6723 512 6739 576
rect 6803 512 6809 576
rect 6493 511 6809 512
rect 10426 576 10742 577
rect 10426 512 10432 576
rect 10496 512 10512 576
rect 10576 512 10592 576
rect 10656 512 10672 576
rect 10736 512 10742 576
rect 10426 511 10742 512
rect 14359 576 14675 577
rect 14359 512 14365 576
rect 14429 512 14445 576
rect 14509 512 14525 576
rect 14589 512 14605 576
rect 14669 512 14675 576
rect 14359 511 14675 512
rect 10777 370 10843 373
rect 10642 368 10843 370
rect 10642 312 10782 368
rect 10838 312 10843 368
rect 10642 310 10843 312
rect 10642 234 10702 310
rect 10777 307 10843 310
rect 10642 200 10794 234
rect 1096 98 1216 200
rect 1301 98 1367 101
rect 1096 96 1367 98
rect 1096 40 1306 96
rect 1362 40 1367 96
rect 1096 38 1367 40
rect 1096 0 1216 38
rect 1301 35 1367 38
rect 3000 98 3120 200
rect 3233 98 3299 101
rect 3000 96 3299 98
rect 3000 40 3238 96
rect 3294 40 3299 96
rect 3000 38 3299 40
rect 3000 0 3120 38
rect 3233 35 3299 38
rect 4904 98 5024 200
rect 5257 98 5323 101
rect 4904 96 5323 98
rect 4904 40 5262 96
rect 5318 40 5323 96
rect 4904 38 5323 40
rect 4904 0 5024 38
rect 5257 35 5323 38
rect 6808 98 6928 200
rect 7097 98 7163 101
rect 6808 96 7163 98
rect 6808 40 7102 96
rect 7158 40 7163 96
rect 6808 38 7163 40
rect 6808 0 6928 38
rect 7097 35 7163 38
rect 8712 98 8832 200
rect 8937 98 9003 101
rect 8712 96 9003 98
rect 8712 40 8942 96
rect 8998 40 9003 96
rect 8712 38 9003 40
rect 8712 0 8832 38
rect 8937 35 9003 38
rect 10616 38 10794 200
rect 12520 98 12640 200
rect 12801 98 12867 101
rect 12520 96 12867 98
rect 12520 40 12806 96
rect 12862 40 12867 96
rect 12520 38 12867 40
rect 10616 0 10736 38
rect 12520 0 12640 38
rect 12801 35 12867 38
rect 14424 98 14544 200
rect 14733 98 14799 101
rect 14424 96 14799 98
rect 14424 40 14738 96
rect 14794 40 14799 96
rect 14424 38 14799 40
rect 14424 0 14544 38
rect 14733 35 14799 38
<< via3 >>
rect 1906 13084 1970 13088
rect 1906 13028 1910 13084
rect 1910 13028 1966 13084
rect 1966 13028 1970 13084
rect 1906 13024 1970 13028
rect 1986 13084 2050 13088
rect 1986 13028 1990 13084
rect 1990 13028 2046 13084
rect 2046 13028 2050 13084
rect 1986 13024 2050 13028
rect 2066 13084 2130 13088
rect 2066 13028 2070 13084
rect 2070 13028 2126 13084
rect 2126 13028 2130 13084
rect 2066 13024 2130 13028
rect 2146 13084 2210 13088
rect 2146 13028 2150 13084
rect 2150 13028 2206 13084
rect 2206 13028 2210 13084
rect 2146 13024 2210 13028
rect 5839 13084 5903 13088
rect 5839 13028 5843 13084
rect 5843 13028 5899 13084
rect 5899 13028 5903 13084
rect 5839 13024 5903 13028
rect 5919 13084 5983 13088
rect 5919 13028 5923 13084
rect 5923 13028 5979 13084
rect 5979 13028 5983 13084
rect 5919 13024 5983 13028
rect 5999 13084 6063 13088
rect 5999 13028 6003 13084
rect 6003 13028 6059 13084
rect 6059 13028 6063 13084
rect 5999 13024 6063 13028
rect 6079 13084 6143 13088
rect 6079 13028 6083 13084
rect 6083 13028 6139 13084
rect 6139 13028 6143 13084
rect 6079 13024 6143 13028
rect 9772 13084 9836 13088
rect 9772 13028 9776 13084
rect 9776 13028 9832 13084
rect 9832 13028 9836 13084
rect 9772 13024 9836 13028
rect 9852 13084 9916 13088
rect 9852 13028 9856 13084
rect 9856 13028 9912 13084
rect 9912 13028 9916 13084
rect 9852 13024 9916 13028
rect 9932 13084 9996 13088
rect 9932 13028 9936 13084
rect 9936 13028 9992 13084
rect 9992 13028 9996 13084
rect 9932 13024 9996 13028
rect 10012 13084 10076 13088
rect 10012 13028 10016 13084
rect 10016 13028 10072 13084
rect 10072 13028 10076 13084
rect 10012 13024 10076 13028
rect 13705 13084 13769 13088
rect 13705 13028 13709 13084
rect 13709 13028 13765 13084
rect 13765 13028 13769 13084
rect 13705 13024 13769 13028
rect 13785 13084 13849 13088
rect 13785 13028 13789 13084
rect 13789 13028 13845 13084
rect 13845 13028 13849 13084
rect 13785 13024 13849 13028
rect 13865 13084 13929 13088
rect 13865 13028 13869 13084
rect 13869 13028 13925 13084
rect 13925 13028 13929 13084
rect 13865 13024 13929 13028
rect 13945 13084 14009 13088
rect 13945 13028 13949 13084
rect 13949 13028 14005 13084
rect 14005 13028 14009 13084
rect 13945 13024 14009 13028
rect 2566 12540 2630 12544
rect 2566 12484 2570 12540
rect 2570 12484 2626 12540
rect 2626 12484 2630 12540
rect 2566 12480 2630 12484
rect 2646 12540 2710 12544
rect 2646 12484 2650 12540
rect 2650 12484 2706 12540
rect 2706 12484 2710 12540
rect 2646 12480 2710 12484
rect 2726 12540 2790 12544
rect 2726 12484 2730 12540
rect 2730 12484 2786 12540
rect 2786 12484 2790 12540
rect 2726 12480 2790 12484
rect 2806 12540 2870 12544
rect 2806 12484 2810 12540
rect 2810 12484 2866 12540
rect 2866 12484 2870 12540
rect 2806 12480 2870 12484
rect 6499 12540 6563 12544
rect 6499 12484 6503 12540
rect 6503 12484 6559 12540
rect 6559 12484 6563 12540
rect 6499 12480 6563 12484
rect 6579 12540 6643 12544
rect 6579 12484 6583 12540
rect 6583 12484 6639 12540
rect 6639 12484 6643 12540
rect 6579 12480 6643 12484
rect 6659 12540 6723 12544
rect 6659 12484 6663 12540
rect 6663 12484 6719 12540
rect 6719 12484 6723 12540
rect 6659 12480 6723 12484
rect 6739 12540 6803 12544
rect 6739 12484 6743 12540
rect 6743 12484 6799 12540
rect 6799 12484 6803 12540
rect 6739 12480 6803 12484
rect 10432 12540 10496 12544
rect 10432 12484 10436 12540
rect 10436 12484 10492 12540
rect 10492 12484 10496 12540
rect 10432 12480 10496 12484
rect 10512 12540 10576 12544
rect 10512 12484 10516 12540
rect 10516 12484 10572 12540
rect 10572 12484 10576 12540
rect 10512 12480 10576 12484
rect 10592 12540 10656 12544
rect 10592 12484 10596 12540
rect 10596 12484 10652 12540
rect 10652 12484 10656 12540
rect 10592 12480 10656 12484
rect 10672 12540 10736 12544
rect 10672 12484 10676 12540
rect 10676 12484 10732 12540
rect 10732 12484 10736 12540
rect 10672 12480 10736 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 14605 12540 14669 12544
rect 14605 12484 14609 12540
rect 14609 12484 14665 12540
rect 14665 12484 14669 12540
rect 14605 12480 14669 12484
rect 1906 11996 1970 12000
rect 1906 11940 1910 11996
rect 1910 11940 1966 11996
rect 1966 11940 1970 11996
rect 1906 11936 1970 11940
rect 1986 11996 2050 12000
rect 1986 11940 1990 11996
rect 1990 11940 2046 11996
rect 2046 11940 2050 11996
rect 1986 11936 2050 11940
rect 2066 11996 2130 12000
rect 2066 11940 2070 11996
rect 2070 11940 2126 11996
rect 2126 11940 2130 11996
rect 2066 11936 2130 11940
rect 2146 11996 2210 12000
rect 2146 11940 2150 11996
rect 2150 11940 2206 11996
rect 2206 11940 2210 11996
rect 2146 11936 2210 11940
rect 5839 11996 5903 12000
rect 5839 11940 5843 11996
rect 5843 11940 5899 11996
rect 5899 11940 5903 11996
rect 5839 11936 5903 11940
rect 5919 11996 5983 12000
rect 5919 11940 5923 11996
rect 5923 11940 5979 11996
rect 5979 11940 5983 11996
rect 5919 11936 5983 11940
rect 5999 11996 6063 12000
rect 5999 11940 6003 11996
rect 6003 11940 6059 11996
rect 6059 11940 6063 11996
rect 5999 11936 6063 11940
rect 6079 11996 6143 12000
rect 6079 11940 6083 11996
rect 6083 11940 6139 11996
rect 6139 11940 6143 11996
rect 6079 11936 6143 11940
rect 9772 11996 9836 12000
rect 9772 11940 9776 11996
rect 9776 11940 9832 11996
rect 9832 11940 9836 11996
rect 9772 11936 9836 11940
rect 9852 11996 9916 12000
rect 9852 11940 9856 11996
rect 9856 11940 9912 11996
rect 9912 11940 9916 11996
rect 9852 11936 9916 11940
rect 9932 11996 9996 12000
rect 9932 11940 9936 11996
rect 9936 11940 9992 11996
rect 9992 11940 9996 11996
rect 9932 11936 9996 11940
rect 10012 11996 10076 12000
rect 10012 11940 10016 11996
rect 10016 11940 10072 11996
rect 10072 11940 10076 11996
rect 10012 11936 10076 11940
rect 13705 11996 13769 12000
rect 13705 11940 13709 11996
rect 13709 11940 13765 11996
rect 13765 11940 13769 11996
rect 13705 11936 13769 11940
rect 13785 11996 13849 12000
rect 13785 11940 13789 11996
rect 13789 11940 13845 11996
rect 13845 11940 13849 11996
rect 13785 11936 13849 11940
rect 13865 11996 13929 12000
rect 13865 11940 13869 11996
rect 13869 11940 13925 11996
rect 13925 11940 13929 11996
rect 13865 11936 13929 11940
rect 13945 11996 14009 12000
rect 13945 11940 13949 11996
rect 13949 11940 14005 11996
rect 14005 11940 14009 11996
rect 13945 11936 14009 11940
rect 2566 11452 2630 11456
rect 2566 11396 2570 11452
rect 2570 11396 2626 11452
rect 2626 11396 2630 11452
rect 2566 11392 2630 11396
rect 2646 11452 2710 11456
rect 2646 11396 2650 11452
rect 2650 11396 2706 11452
rect 2706 11396 2710 11452
rect 2646 11392 2710 11396
rect 2726 11452 2790 11456
rect 2726 11396 2730 11452
rect 2730 11396 2786 11452
rect 2786 11396 2790 11452
rect 2726 11392 2790 11396
rect 2806 11452 2870 11456
rect 2806 11396 2810 11452
rect 2810 11396 2866 11452
rect 2866 11396 2870 11452
rect 2806 11392 2870 11396
rect 6499 11452 6563 11456
rect 6499 11396 6503 11452
rect 6503 11396 6559 11452
rect 6559 11396 6563 11452
rect 6499 11392 6563 11396
rect 6579 11452 6643 11456
rect 6579 11396 6583 11452
rect 6583 11396 6639 11452
rect 6639 11396 6643 11452
rect 6579 11392 6643 11396
rect 6659 11452 6723 11456
rect 6659 11396 6663 11452
rect 6663 11396 6719 11452
rect 6719 11396 6723 11452
rect 6659 11392 6723 11396
rect 6739 11452 6803 11456
rect 6739 11396 6743 11452
rect 6743 11396 6799 11452
rect 6799 11396 6803 11452
rect 6739 11392 6803 11396
rect 10432 11452 10496 11456
rect 10432 11396 10436 11452
rect 10436 11396 10492 11452
rect 10492 11396 10496 11452
rect 10432 11392 10496 11396
rect 10512 11452 10576 11456
rect 10512 11396 10516 11452
rect 10516 11396 10572 11452
rect 10572 11396 10576 11452
rect 10512 11392 10576 11396
rect 10592 11452 10656 11456
rect 10592 11396 10596 11452
rect 10596 11396 10652 11452
rect 10652 11396 10656 11452
rect 10592 11392 10656 11396
rect 10672 11452 10736 11456
rect 10672 11396 10676 11452
rect 10676 11396 10732 11452
rect 10732 11396 10736 11452
rect 10672 11392 10736 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 14605 11452 14669 11456
rect 14605 11396 14609 11452
rect 14609 11396 14665 11452
rect 14665 11396 14669 11452
rect 14605 11392 14669 11396
rect 1906 10908 1970 10912
rect 1906 10852 1910 10908
rect 1910 10852 1966 10908
rect 1966 10852 1970 10908
rect 1906 10848 1970 10852
rect 1986 10908 2050 10912
rect 1986 10852 1990 10908
rect 1990 10852 2046 10908
rect 2046 10852 2050 10908
rect 1986 10848 2050 10852
rect 2066 10908 2130 10912
rect 2066 10852 2070 10908
rect 2070 10852 2126 10908
rect 2126 10852 2130 10908
rect 2066 10848 2130 10852
rect 2146 10908 2210 10912
rect 2146 10852 2150 10908
rect 2150 10852 2206 10908
rect 2206 10852 2210 10908
rect 2146 10848 2210 10852
rect 5839 10908 5903 10912
rect 5839 10852 5843 10908
rect 5843 10852 5899 10908
rect 5899 10852 5903 10908
rect 5839 10848 5903 10852
rect 5919 10908 5983 10912
rect 5919 10852 5923 10908
rect 5923 10852 5979 10908
rect 5979 10852 5983 10908
rect 5919 10848 5983 10852
rect 5999 10908 6063 10912
rect 5999 10852 6003 10908
rect 6003 10852 6059 10908
rect 6059 10852 6063 10908
rect 5999 10848 6063 10852
rect 6079 10908 6143 10912
rect 6079 10852 6083 10908
rect 6083 10852 6139 10908
rect 6139 10852 6143 10908
rect 6079 10848 6143 10852
rect 9772 10908 9836 10912
rect 9772 10852 9776 10908
rect 9776 10852 9832 10908
rect 9832 10852 9836 10908
rect 9772 10848 9836 10852
rect 9852 10908 9916 10912
rect 9852 10852 9856 10908
rect 9856 10852 9912 10908
rect 9912 10852 9916 10908
rect 9852 10848 9916 10852
rect 9932 10908 9996 10912
rect 9932 10852 9936 10908
rect 9936 10852 9992 10908
rect 9992 10852 9996 10908
rect 9932 10848 9996 10852
rect 10012 10908 10076 10912
rect 10012 10852 10016 10908
rect 10016 10852 10072 10908
rect 10072 10852 10076 10908
rect 10012 10848 10076 10852
rect 13705 10908 13769 10912
rect 13705 10852 13709 10908
rect 13709 10852 13765 10908
rect 13765 10852 13769 10908
rect 13705 10848 13769 10852
rect 13785 10908 13849 10912
rect 13785 10852 13789 10908
rect 13789 10852 13845 10908
rect 13845 10852 13849 10908
rect 13785 10848 13849 10852
rect 13865 10908 13929 10912
rect 13865 10852 13869 10908
rect 13869 10852 13925 10908
rect 13925 10852 13929 10908
rect 13865 10848 13929 10852
rect 13945 10908 14009 10912
rect 13945 10852 13949 10908
rect 13949 10852 14005 10908
rect 14005 10852 14009 10908
rect 13945 10848 14009 10852
rect 2566 10364 2630 10368
rect 2566 10308 2570 10364
rect 2570 10308 2626 10364
rect 2626 10308 2630 10364
rect 2566 10304 2630 10308
rect 2646 10364 2710 10368
rect 2646 10308 2650 10364
rect 2650 10308 2706 10364
rect 2706 10308 2710 10364
rect 2646 10304 2710 10308
rect 2726 10364 2790 10368
rect 2726 10308 2730 10364
rect 2730 10308 2786 10364
rect 2786 10308 2790 10364
rect 2726 10304 2790 10308
rect 2806 10364 2870 10368
rect 2806 10308 2810 10364
rect 2810 10308 2866 10364
rect 2866 10308 2870 10364
rect 2806 10304 2870 10308
rect 6499 10364 6563 10368
rect 6499 10308 6503 10364
rect 6503 10308 6559 10364
rect 6559 10308 6563 10364
rect 6499 10304 6563 10308
rect 6579 10364 6643 10368
rect 6579 10308 6583 10364
rect 6583 10308 6639 10364
rect 6639 10308 6643 10364
rect 6579 10304 6643 10308
rect 6659 10364 6723 10368
rect 6659 10308 6663 10364
rect 6663 10308 6719 10364
rect 6719 10308 6723 10364
rect 6659 10304 6723 10308
rect 6739 10364 6803 10368
rect 6739 10308 6743 10364
rect 6743 10308 6799 10364
rect 6799 10308 6803 10364
rect 6739 10304 6803 10308
rect 10432 10364 10496 10368
rect 10432 10308 10436 10364
rect 10436 10308 10492 10364
rect 10492 10308 10496 10364
rect 10432 10304 10496 10308
rect 10512 10364 10576 10368
rect 10512 10308 10516 10364
rect 10516 10308 10572 10364
rect 10572 10308 10576 10364
rect 10512 10304 10576 10308
rect 10592 10364 10656 10368
rect 10592 10308 10596 10364
rect 10596 10308 10652 10364
rect 10652 10308 10656 10364
rect 10592 10304 10656 10308
rect 10672 10364 10736 10368
rect 10672 10308 10676 10364
rect 10676 10308 10732 10364
rect 10732 10308 10736 10364
rect 10672 10304 10736 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 14605 10364 14669 10368
rect 14605 10308 14609 10364
rect 14609 10308 14665 10364
rect 14665 10308 14669 10364
rect 14605 10304 14669 10308
rect 1906 9820 1970 9824
rect 1906 9764 1910 9820
rect 1910 9764 1966 9820
rect 1966 9764 1970 9820
rect 1906 9760 1970 9764
rect 1986 9820 2050 9824
rect 1986 9764 1990 9820
rect 1990 9764 2046 9820
rect 2046 9764 2050 9820
rect 1986 9760 2050 9764
rect 2066 9820 2130 9824
rect 2066 9764 2070 9820
rect 2070 9764 2126 9820
rect 2126 9764 2130 9820
rect 2066 9760 2130 9764
rect 2146 9820 2210 9824
rect 2146 9764 2150 9820
rect 2150 9764 2206 9820
rect 2206 9764 2210 9820
rect 2146 9760 2210 9764
rect 5839 9820 5903 9824
rect 5839 9764 5843 9820
rect 5843 9764 5899 9820
rect 5899 9764 5903 9820
rect 5839 9760 5903 9764
rect 5919 9820 5983 9824
rect 5919 9764 5923 9820
rect 5923 9764 5979 9820
rect 5979 9764 5983 9820
rect 5919 9760 5983 9764
rect 5999 9820 6063 9824
rect 5999 9764 6003 9820
rect 6003 9764 6059 9820
rect 6059 9764 6063 9820
rect 5999 9760 6063 9764
rect 6079 9820 6143 9824
rect 6079 9764 6083 9820
rect 6083 9764 6139 9820
rect 6139 9764 6143 9820
rect 6079 9760 6143 9764
rect 9772 9820 9836 9824
rect 9772 9764 9776 9820
rect 9776 9764 9832 9820
rect 9832 9764 9836 9820
rect 9772 9760 9836 9764
rect 9852 9820 9916 9824
rect 9852 9764 9856 9820
rect 9856 9764 9912 9820
rect 9912 9764 9916 9820
rect 9852 9760 9916 9764
rect 9932 9820 9996 9824
rect 9932 9764 9936 9820
rect 9936 9764 9992 9820
rect 9992 9764 9996 9820
rect 9932 9760 9996 9764
rect 10012 9820 10076 9824
rect 10012 9764 10016 9820
rect 10016 9764 10072 9820
rect 10072 9764 10076 9820
rect 10012 9760 10076 9764
rect 13705 9820 13769 9824
rect 13705 9764 13709 9820
rect 13709 9764 13765 9820
rect 13765 9764 13769 9820
rect 13705 9760 13769 9764
rect 13785 9820 13849 9824
rect 13785 9764 13789 9820
rect 13789 9764 13845 9820
rect 13845 9764 13849 9820
rect 13785 9760 13849 9764
rect 13865 9820 13929 9824
rect 13865 9764 13869 9820
rect 13869 9764 13925 9820
rect 13925 9764 13929 9820
rect 13865 9760 13929 9764
rect 13945 9820 14009 9824
rect 13945 9764 13949 9820
rect 13949 9764 14005 9820
rect 14005 9764 14009 9820
rect 13945 9760 14009 9764
rect 2566 9276 2630 9280
rect 2566 9220 2570 9276
rect 2570 9220 2626 9276
rect 2626 9220 2630 9276
rect 2566 9216 2630 9220
rect 2646 9276 2710 9280
rect 2646 9220 2650 9276
rect 2650 9220 2706 9276
rect 2706 9220 2710 9276
rect 2646 9216 2710 9220
rect 2726 9276 2790 9280
rect 2726 9220 2730 9276
rect 2730 9220 2786 9276
rect 2786 9220 2790 9276
rect 2726 9216 2790 9220
rect 2806 9276 2870 9280
rect 2806 9220 2810 9276
rect 2810 9220 2866 9276
rect 2866 9220 2870 9276
rect 2806 9216 2870 9220
rect 6499 9276 6563 9280
rect 6499 9220 6503 9276
rect 6503 9220 6559 9276
rect 6559 9220 6563 9276
rect 6499 9216 6563 9220
rect 6579 9276 6643 9280
rect 6579 9220 6583 9276
rect 6583 9220 6639 9276
rect 6639 9220 6643 9276
rect 6579 9216 6643 9220
rect 6659 9276 6723 9280
rect 6659 9220 6663 9276
rect 6663 9220 6719 9276
rect 6719 9220 6723 9276
rect 6659 9216 6723 9220
rect 6739 9276 6803 9280
rect 6739 9220 6743 9276
rect 6743 9220 6799 9276
rect 6799 9220 6803 9276
rect 6739 9216 6803 9220
rect 10432 9276 10496 9280
rect 10432 9220 10436 9276
rect 10436 9220 10492 9276
rect 10492 9220 10496 9276
rect 10432 9216 10496 9220
rect 10512 9276 10576 9280
rect 10512 9220 10516 9276
rect 10516 9220 10572 9276
rect 10572 9220 10576 9276
rect 10512 9216 10576 9220
rect 10592 9276 10656 9280
rect 10592 9220 10596 9276
rect 10596 9220 10652 9276
rect 10652 9220 10656 9276
rect 10592 9216 10656 9220
rect 10672 9276 10736 9280
rect 10672 9220 10676 9276
rect 10676 9220 10732 9276
rect 10732 9220 10736 9276
rect 10672 9216 10736 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 14605 9276 14669 9280
rect 14605 9220 14609 9276
rect 14609 9220 14665 9276
rect 14665 9220 14669 9276
rect 14605 9216 14669 9220
rect 1906 8732 1970 8736
rect 1906 8676 1910 8732
rect 1910 8676 1966 8732
rect 1966 8676 1970 8732
rect 1906 8672 1970 8676
rect 1986 8732 2050 8736
rect 1986 8676 1990 8732
rect 1990 8676 2046 8732
rect 2046 8676 2050 8732
rect 1986 8672 2050 8676
rect 2066 8732 2130 8736
rect 2066 8676 2070 8732
rect 2070 8676 2126 8732
rect 2126 8676 2130 8732
rect 2066 8672 2130 8676
rect 2146 8732 2210 8736
rect 2146 8676 2150 8732
rect 2150 8676 2206 8732
rect 2206 8676 2210 8732
rect 2146 8672 2210 8676
rect 5839 8732 5903 8736
rect 5839 8676 5843 8732
rect 5843 8676 5899 8732
rect 5899 8676 5903 8732
rect 5839 8672 5903 8676
rect 5919 8732 5983 8736
rect 5919 8676 5923 8732
rect 5923 8676 5979 8732
rect 5979 8676 5983 8732
rect 5919 8672 5983 8676
rect 5999 8732 6063 8736
rect 5999 8676 6003 8732
rect 6003 8676 6059 8732
rect 6059 8676 6063 8732
rect 5999 8672 6063 8676
rect 6079 8732 6143 8736
rect 6079 8676 6083 8732
rect 6083 8676 6139 8732
rect 6139 8676 6143 8732
rect 6079 8672 6143 8676
rect 9772 8732 9836 8736
rect 9772 8676 9776 8732
rect 9776 8676 9832 8732
rect 9832 8676 9836 8732
rect 9772 8672 9836 8676
rect 9852 8732 9916 8736
rect 9852 8676 9856 8732
rect 9856 8676 9912 8732
rect 9912 8676 9916 8732
rect 9852 8672 9916 8676
rect 9932 8732 9996 8736
rect 9932 8676 9936 8732
rect 9936 8676 9992 8732
rect 9992 8676 9996 8732
rect 9932 8672 9996 8676
rect 10012 8732 10076 8736
rect 10012 8676 10016 8732
rect 10016 8676 10072 8732
rect 10072 8676 10076 8732
rect 10012 8672 10076 8676
rect 13705 8732 13769 8736
rect 13705 8676 13709 8732
rect 13709 8676 13765 8732
rect 13765 8676 13769 8732
rect 13705 8672 13769 8676
rect 13785 8732 13849 8736
rect 13785 8676 13789 8732
rect 13789 8676 13845 8732
rect 13845 8676 13849 8732
rect 13785 8672 13849 8676
rect 13865 8732 13929 8736
rect 13865 8676 13869 8732
rect 13869 8676 13925 8732
rect 13925 8676 13929 8732
rect 13865 8672 13929 8676
rect 13945 8732 14009 8736
rect 13945 8676 13949 8732
rect 13949 8676 14005 8732
rect 14005 8676 14009 8732
rect 13945 8672 14009 8676
rect 2566 8188 2630 8192
rect 2566 8132 2570 8188
rect 2570 8132 2626 8188
rect 2626 8132 2630 8188
rect 2566 8128 2630 8132
rect 2646 8188 2710 8192
rect 2646 8132 2650 8188
rect 2650 8132 2706 8188
rect 2706 8132 2710 8188
rect 2646 8128 2710 8132
rect 2726 8188 2790 8192
rect 2726 8132 2730 8188
rect 2730 8132 2786 8188
rect 2786 8132 2790 8188
rect 2726 8128 2790 8132
rect 2806 8188 2870 8192
rect 2806 8132 2810 8188
rect 2810 8132 2866 8188
rect 2866 8132 2870 8188
rect 2806 8128 2870 8132
rect 6499 8188 6563 8192
rect 6499 8132 6503 8188
rect 6503 8132 6559 8188
rect 6559 8132 6563 8188
rect 6499 8128 6563 8132
rect 6579 8188 6643 8192
rect 6579 8132 6583 8188
rect 6583 8132 6639 8188
rect 6639 8132 6643 8188
rect 6579 8128 6643 8132
rect 6659 8188 6723 8192
rect 6659 8132 6663 8188
rect 6663 8132 6719 8188
rect 6719 8132 6723 8188
rect 6659 8128 6723 8132
rect 6739 8188 6803 8192
rect 6739 8132 6743 8188
rect 6743 8132 6799 8188
rect 6799 8132 6803 8188
rect 6739 8128 6803 8132
rect 10432 8188 10496 8192
rect 10432 8132 10436 8188
rect 10436 8132 10492 8188
rect 10492 8132 10496 8188
rect 10432 8128 10496 8132
rect 10512 8188 10576 8192
rect 10512 8132 10516 8188
rect 10516 8132 10572 8188
rect 10572 8132 10576 8188
rect 10512 8128 10576 8132
rect 10592 8188 10656 8192
rect 10592 8132 10596 8188
rect 10596 8132 10652 8188
rect 10652 8132 10656 8188
rect 10592 8128 10656 8132
rect 10672 8188 10736 8192
rect 10672 8132 10676 8188
rect 10676 8132 10732 8188
rect 10732 8132 10736 8188
rect 10672 8128 10736 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 14605 8188 14669 8192
rect 14605 8132 14609 8188
rect 14609 8132 14665 8188
rect 14665 8132 14669 8188
rect 14605 8128 14669 8132
rect 1906 7644 1970 7648
rect 1906 7588 1910 7644
rect 1910 7588 1966 7644
rect 1966 7588 1970 7644
rect 1906 7584 1970 7588
rect 1986 7644 2050 7648
rect 1986 7588 1990 7644
rect 1990 7588 2046 7644
rect 2046 7588 2050 7644
rect 1986 7584 2050 7588
rect 2066 7644 2130 7648
rect 2066 7588 2070 7644
rect 2070 7588 2126 7644
rect 2126 7588 2130 7644
rect 2066 7584 2130 7588
rect 2146 7644 2210 7648
rect 2146 7588 2150 7644
rect 2150 7588 2206 7644
rect 2206 7588 2210 7644
rect 2146 7584 2210 7588
rect 5839 7644 5903 7648
rect 5839 7588 5843 7644
rect 5843 7588 5899 7644
rect 5899 7588 5903 7644
rect 5839 7584 5903 7588
rect 5919 7644 5983 7648
rect 5919 7588 5923 7644
rect 5923 7588 5979 7644
rect 5979 7588 5983 7644
rect 5919 7584 5983 7588
rect 5999 7644 6063 7648
rect 5999 7588 6003 7644
rect 6003 7588 6059 7644
rect 6059 7588 6063 7644
rect 5999 7584 6063 7588
rect 6079 7644 6143 7648
rect 6079 7588 6083 7644
rect 6083 7588 6139 7644
rect 6139 7588 6143 7644
rect 6079 7584 6143 7588
rect 9772 7644 9836 7648
rect 9772 7588 9776 7644
rect 9776 7588 9832 7644
rect 9832 7588 9836 7644
rect 9772 7584 9836 7588
rect 9852 7644 9916 7648
rect 9852 7588 9856 7644
rect 9856 7588 9912 7644
rect 9912 7588 9916 7644
rect 9852 7584 9916 7588
rect 9932 7644 9996 7648
rect 9932 7588 9936 7644
rect 9936 7588 9992 7644
rect 9992 7588 9996 7644
rect 9932 7584 9996 7588
rect 10012 7644 10076 7648
rect 10012 7588 10016 7644
rect 10016 7588 10072 7644
rect 10072 7588 10076 7644
rect 10012 7584 10076 7588
rect 13705 7644 13769 7648
rect 13705 7588 13709 7644
rect 13709 7588 13765 7644
rect 13765 7588 13769 7644
rect 13705 7584 13769 7588
rect 13785 7644 13849 7648
rect 13785 7588 13789 7644
rect 13789 7588 13845 7644
rect 13845 7588 13849 7644
rect 13785 7584 13849 7588
rect 13865 7644 13929 7648
rect 13865 7588 13869 7644
rect 13869 7588 13925 7644
rect 13925 7588 13929 7644
rect 13865 7584 13929 7588
rect 13945 7644 14009 7648
rect 13945 7588 13949 7644
rect 13949 7588 14005 7644
rect 14005 7588 14009 7644
rect 13945 7584 14009 7588
rect 2566 7100 2630 7104
rect 2566 7044 2570 7100
rect 2570 7044 2626 7100
rect 2626 7044 2630 7100
rect 2566 7040 2630 7044
rect 2646 7100 2710 7104
rect 2646 7044 2650 7100
rect 2650 7044 2706 7100
rect 2706 7044 2710 7100
rect 2646 7040 2710 7044
rect 2726 7100 2790 7104
rect 2726 7044 2730 7100
rect 2730 7044 2786 7100
rect 2786 7044 2790 7100
rect 2726 7040 2790 7044
rect 2806 7100 2870 7104
rect 2806 7044 2810 7100
rect 2810 7044 2866 7100
rect 2866 7044 2870 7100
rect 2806 7040 2870 7044
rect 6499 7100 6563 7104
rect 6499 7044 6503 7100
rect 6503 7044 6559 7100
rect 6559 7044 6563 7100
rect 6499 7040 6563 7044
rect 6579 7100 6643 7104
rect 6579 7044 6583 7100
rect 6583 7044 6639 7100
rect 6639 7044 6643 7100
rect 6579 7040 6643 7044
rect 6659 7100 6723 7104
rect 6659 7044 6663 7100
rect 6663 7044 6719 7100
rect 6719 7044 6723 7100
rect 6659 7040 6723 7044
rect 6739 7100 6803 7104
rect 6739 7044 6743 7100
rect 6743 7044 6799 7100
rect 6799 7044 6803 7100
rect 6739 7040 6803 7044
rect 10432 7100 10496 7104
rect 10432 7044 10436 7100
rect 10436 7044 10492 7100
rect 10492 7044 10496 7100
rect 10432 7040 10496 7044
rect 10512 7100 10576 7104
rect 10512 7044 10516 7100
rect 10516 7044 10572 7100
rect 10572 7044 10576 7100
rect 10512 7040 10576 7044
rect 10592 7100 10656 7104
rect 10592 7044 10596 7100
rect 10596 7044 10652 7100
rect 10652 7044 10656 7100
rect 10592 7040 10656 7044
rect 10672 7100 10736 7104
rect 10672 7044 10676 7100
rect 10676 7044 10732 7100
rect 10732 7044 10736 7100
rect 10672 7040 10736 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 14605 7100 14669 7104
rect 14605 7044 14609 7100
rect 14609 7044 14665 7100
rect 14665 7044 14669 7100
rect 14605 7040 14669 7044
rect 1906 6556 1970 6560
rect 1906 6500 1910 6556
rect 1910 6500 1966 6556
rect 1966 6500 1970 6556
rect 1906 6496 1970 6500
rect 1986 6556 2050 6560
rect 1986 6500 1990 6556
rect 1990 6500 2046 6556
rect 2046 6500 2050 6556
rect 1986 6496 2050 6500
rect 2066 6556 2130 6560
rect 2066 6500 2070 6556
rect 2070 6500 2126 6556
rect 2126 6500 2130 6556
rect 2066 6496 2130 6500
rect 2146 6556 2210 6560
rect 2146 6500 2150 6556
rect 2150 6500 2206 6556
rect 2206 6500 2210 6556
rect 2146 6496 2210 6500
rect 5839 6556 5903 6560
rect 5839 6500 5843 6556
rect 5843 6500 5899 6556
rect 5899 6500 5903 6556
rect 5839 6496 5903 6500
rect 5919 6556 5983 6560
rect 5919 6500 5923 6556
rect 5923 6500 5979 6556
rect 5979 6500 5983 6556
rect 5919 6496 5983 6500
rect 5999 6556 6063 6560
rect 5999 6500 6003 6556
rect 6003 6500 6059 6556
rect 6059 6500 6063 6556
rect 5999 6496 6063 6500
rect 6079 6556 6143 6560
rect 6079 6500 6083 6556
rect 6083 6500 6139 6556
rect 6139 6500 6143 6556
rect 6079 6496 6143 6500
rect 9772 6556 9836 6560
rect 9772 6500 9776 6556
rect 9776 6500 9832 6556
rect 9832 6500 9836 6556
rect 9772 6496 9836 6500
rect 9852 6556 9916 6560
rect 9852 6500 9856 6556
rect 9856 6500 9912 6556
rect 9912 6500 9916 6556
rect 9852 6496 9916 6500
rect 9932 6556 9996 6560
rect 9932 6500 9936 6556
rect 9936 6500 9992 6556
rect 9992 6500 9996 6556
rect 9932 6496 9996 6500
rect 10012 6556 10076 6560
rect 10012 6500 10016 6556
rect 10016 6500 10072 6556
rect 10072 6500 10076 6556
rect 10012 6496 10076 6500
rect 13705 6556 13769 6560
rect 13705 6500 13709 6556
rect 13709 6500 13765 6556
rect 13765 6500 13769 6556
rect 13705 6496 13769 6500
rect 13785 6556 13849 6560
rect 13785 6500 13789 6556
rect 13789 6500 13845 6556
rect 13845 6500 13849 6556
rect 13785 6496 13849 6500
rect 13865 6556 13929 6560
rect 13865 6500 13869 6556
rect 13869 6500 13925 6556
rect 13925 6500 13929 6556
rect 13865 6496 13929 6500
rect 13945 6556 14009 6560
rect 13945 6500 13949 6556
rect 13949 6500 14005 6556
rect 14005 6500 14009 6556
rect 13945 6496 14009 6500
rect 2566 6012 2630 6016
rect 2566 5956 2570 6012
rect 2570 5956 2626 6012
rect 2626 5956 2630 6012
rect 2566 5952 2630 5956
rect 2646 6012 2710 6016
rect 2646 5956 2650 6012
rect 2650 5956 2706 6012
rect 2706 5956 2710 6012
rect 2646 5952 2710 5956
rect 2726 6012 2790 6016
rect 2726 5956 2730 6012
rect 2730 5956 2786 6012
rect 2786 5956 2790 6012
rect 2726 5952 2790 5956
rect 2806 6012 2870 6016
rect 2806 5956 2810 6012
rect 2810 5956 2866 6012
rect 2866 5956 2870 6012
rect 2806 5952 2870 5956
rect 6499 6012 6563 6016
rect 6499 5956 6503 6012
rect 6503 5956 6559 6012
rect 6559 5956 6563 6012
rect 6499 5952 6563 5956
rect 6579 6012 6643 6016
rect 6579 5956 6583 6012
rect 6583 5956 6639 6012
rect 6639 5956 6643 6012
rect 6579 5952 6643 5956
rect 6659 6012 6723 6016
rect 6659 5956 6663 6012
rect 6663 5956 6719 6012
rect 6719 5956 6723 6012
rect 6659 5952 6723 5956
rect 6739 6012 6803 6016
rect 6739 5956 6743 6012
rect 6743 5956 6799 6012
rect 6799 5956 6803 6012
rect 6739 5952 6803 5956
rect 10432 6012 10496 6016
rect 10432 5956 10436 6012
rect 10436 5956 10492 6012
rect 10492 5956 10496 6012
rect 10432 5952 10496 5956
rect 10512 6012 10576 6016
rect 10512 5956 10516 6012
rect 10516 5956 10572 6012
rect 10572 5956 10576 6012
rect 10512 5952 10576 5956
rect 10592 6012 10656 6016
rect 10592 5956 10596 6012
rect 10596 5956 10652 6012
rect 10652 5956 10656 6012
rect 10592 5952 10656 5956
rect 10672 6012 10736 6016
rect 10672 5956 10676 6012
rect 10676 5956 10732 6012
rect 10732 5956 10736 6012
rect 10672 5952 10736 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 14605 6012 14669 6016
rect 14605 5956 14609 6012
rect 14609 5956 14665 6012
rect 14665 5956 14669 6012
rect 14605 5952 14669 5956
rect 1906 5468 1970 5472
rect 1906 5412 1910 5468
rect 1910 5412 1966 5468
rect 1966 5412 1970 5468
rect 1906 5408 1970 5412
rect 1986 5468 2050 5472
rect 1986 5412 1990 5468
rect 1990 5412 2046 5468
rect 2046 5412 2050 5468
rect 1986 5408 2050 5412
rect 2066 5468 2130 5472
rect 2066 5412 2070 5468
rect 2070 5412 2126 5468
rect 2126 5412 2130 5468
rect 2066 5408 2130 5412
rect 2146 5468 2210 5472
rect 2146 5412 2150 5468
rect 2150 5412 2206 5468
rect 2206 5412 2210 5468
rect 2146 5408 2210 5412
rect 5839 5468 5903 5472
rect 5839 5412 5843 5468
rect 5843 5412 5899 5468
rect 5899 5412 5903 5468
rect 5839 5408 5903 5412
rect 5919 5468 5983 5472
rect 5919 5412 5923 5468
rect 5923 5412 5979 5468
rect 5979 5412 5983 5468
rect 5919 5408 5983 5412
rect 5999 5468 6063 5472
rect 5999 5412 6003 5468
rect 6003 5412 6059 5468
rect 6059 5412 6063 5468
rect 5999 5408 6063 5412
rect 6079 5468 6143 5472
rect 6079 5412 6083 5468
rect 6083 5412 6139 5468
rect 6139 5412 6143 5468
rect 6079 5408 6143 5412
rect 9772 5468 9836 5472
rect 9772 5412 9776 5468
rect 9776 5412 9832 5468
rect 9832 5412 9836 5468
rect 9772 5408 9836 5412
rect 9852 5468 9916 5472
rect 9852 5412 9856 5468
rect 9856 5412 9912 5468
rect 9912 5412 9916 5468
rect 9852 5408 9916 5412
rect 9932 5468 9996 5472
rect 9932 5412 9936 5468
rect 9936 5412 9992 5468
rect 9992 5412 9996 5468
rect 9932 5408 9996 5412
rect 10012 5468 10076 5472
rect 10012 5412 10016 5468
rect 10016 5412 10072 5468
rect 10072 5412 10076 5468
rect 10012 5408 10076 5412
rect 13705 5468 13769 5472
rect 13705 5412 13709 5468
rect 13709 5412 13765 5468
rect 13765 5412 13769 5468
rect 13705 5408 13769 5412
rect 13785 5468 13849 5472
rect 13785 5412 13789 5468
rect 13789 5412 13845 5468
rect 13845 5412 13849 5468
rect 13785 5408 13849 5412
rect 13865 5468 13929 5472
rect 13865 5412 13869 5468
rect 13869 5412 13925 5468
rect 13925 5412 13929 5468
rect 13865 5408 13929 5412
rect 13945 5468 14009 5472
rect 13945 5412 13949 5468
rect 13949 5412 14005 5468
rect 14005 5412 14009 5468
rect 13945 5408 14009 5412
rect 2566 4924 2630 4928
rect 2566 4868 2570 4924
rect 2570 4868 2626 4924
rect 2626 4868 2630 4924
rect 2566 4864 2630 4868
rect 2646 4924 2710 4928
rect 2646 4868 2650 4924
rect 2650 4868 2706 4924
rect 2706 4868 2710 4924
rect 2646 4864 2710 4868
rect 2726 4924 2790 4928
rect 2726 4868 2730 4924
rect 2730 4868 2786 4924
rect 2786 4868 2790 4924
rect 2726 4864 2790 4868
rect 2806 4924 2870 4928
rect 2806 4868 2810 4924
rect 2810 4868 2866 4924
rect 2866 4868 2870 4924
rect 2806 4864 2870 4868
rect 6499 4924 6563 4928
rect 6499 4868 6503 4924
rect 6503 4868 6559 4924
rect 6559 4868 6563 4924
rect 6499 4864 6563 4868
rect 6579 4924 6643 4928
rect 6579 4868 6583 4924
rect 6583 4868 6639 4924
rect 6639 4868 6643 4924
rect 6579 4864 6643 4868
rect 6659 4924 6723 4928
rect 6659 4868 6663 4924
rect 6663 4868 6719 4924
rect 6719 4868 6723 4924
rect 6659 4864 6723 4868
rect 6739 4924 6803 4928
rect 6739 4868 6743 4924
rect 6743 4868 6799 4924
rect 6799 4868 6803 4924
rect 6739 4864 6803 4868
rect 10432 4924 10496 4928
rect 10432 4868 10436 4924
rect 10436 4868 10492 4924
rect 10492 4868 10496 4924
rect 10432 4864 10496 4868
rect 10512 4924 10576 4928
rect 10512 4868 10516 4924
rect 10516 4868 10572 4924
rect 10572 4868 10576 4924
rect 10512 4864 10576 4868
rect 10592 4924 10656 4928
rect 10592 4868 10596 4924
rect 10596 4868 10652 4924
rect 10652 4868 10656 4924
rect 10592 4864 10656 4868
rect 10672 4924 10736 4928
rect 10672 4868 10676 4924
rect 10676 4868 10732 4924
rect 10732 4868 10736 4924
rect 10672 4864 10736 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 14605 4924 14669 4928
rect 14605 4868 14609 4924
rect 14609 4868 14665 4924
rect 14665 4868 14669 4924
rect 14605 4864 14669 4868
rect 1906 4380 1970 4384
rect 1906 4324 1910 4380
rect 1910 4324 1966 4380
rect 1966 4324 1970 4380
rect 1906 4320 1970 4324
rect 1986 4380 2050 4384
rect 1986 4324 1990 4380
rect 1990 4324 2046 4380
rect 2046 4324 2050 4380
rect 1986 4320 2050 4324
rect 2066 4380 2130 4384
rect 2066 4324 2070 4380
rect 2070 4324 2126 4380
rect 2126 4324 2130 4380
rect 2066 4320 2130 4324
rect 2146 4380 2210 4384
rect 2146 4324 2150 4380
rect 2150 4324 2206 4380
rect 2206 4324 2210 4380
rect 2146 4320 2210 4324
rect 5839 4380 5903 4384
rect 5839 4324 5843 4380
rect 5843 4324 5899 4380
rect 5899 4324 5903 4380
rect 5839 4320 5903 4324
rect 5919 4380 5983 4384
rect 5919 4324 5923 4380
rect 5923 4324 5979 4380
rect 5979 4324 5983 4380
rect 5919 4320 5983 4324
rect 5999 4380 6063 4384
rect 5999 4324 6003 4380
rect 6003 4324 6059 4380
rect 6059 4324 6063 4380
rect 5999 4320 6063 4324
rect 6079 4380 6143 4384
rect 6079 4324 6083 4380
rect 6083 4324 6139 4380
rect 6139 4324 6143 4380
rect 6079 4320 6143 4324
rect 9772 4380 9836 4384
rect 9772 4324 9776 4380
rect 9776 4324 9832 4380
rect 9832 4324 9836 4380
rect 9772 4320 9836 4324
rect 9852 4380 9916 4384
rect 9852 4324 9856 4380
rect 9856 4324 9912 4380
rect 9912 4324 9916 4380
rect 9852 4320 9916 4324
rect 9932 4380 9996 4384
rect 9932 4324 9936 4380
rect 9936 4324 9992 4380
rect 9992 4324 9996 4380
rect 9932 4320 9996 4324
rect 10012 4380 10076 4384
rect 10012 4324 10016 4380
rect 10016 4324 10072 4380
rect 10072 4324 10076 4380
rect 10012 4320 10076 4324
rect 13705 4380 13769 4384
rect 13705 4324 13709 4380
rect 13709 4324 13765 4380
rect 13765 4324 13769 4380
rect 13705 4320 13769 4324
rect 13785 4380 13849 4384
rect 13785 4324 13789 4380
rect 13789 4324 13845 4380
rect 13845 4324 13849 4380
rect 13785 4320 13849 4324
rect 13865 4380 13929 4384
rect 13865 4324 13869 4380
rect 13869 4324 13925 4380
rect 13925 4324 13929 4380
rect 13865 4320 13929 4324
rect 13945 4380 14009 4384
rect 13945 4324 13949 4380
rect 13949 4324 14005 4380
rect 14005 4324 14009 4380
rect 13945 4320 14009 4324
rect 2566 3836 2630 3840
rect 2566 3780 2570 3836
rect 2570 3780 2626 3836
rect 2626 3780 2630 3836
rect 2566 3776 2630 3780
rect 2646 3836 2710 3840
rect 2646 3780 2650 3836
rect 2650 3780 2706 3836
rect 2706 3780 2710 3836
rect 2646 3776 2710 3780
rect 2726 3836 2790 3840
rect 2726 3780 2730 3836
rect 2730 3780 2786 3836
rect 2786 3780 2790 3836
rect 2726 3776 2790 3780
rect 2806 3836 2870 3840
rect 2806 3780 2810 3836
rect 2810 3780 2866 3836
rect 2866 3780 2870 3836
rect 2806 3776 2870 3780
rect 6499 3836 6563 3840
rect 6499 3780 6503 3836
rect 6503 3780 6559 3836
rect 6559 3780 6563 3836
rect 6499 3776 6563 3780
rect 6579 3836 6643 3840
rect 6579 3780 6583 3836
rect 6583 3780 6639 3836
rect 6639 3780 6643 3836
rect 6579 3776 6643 3780
rect 6659 3836 6723 3840
rect 6659 3780 6663 3836
rect 6663 3780 6719 3836
rect 6719 3780 6723 3836
rect 6659 3776 6723 3780
rect 6739 3836 6803 3840
rect 6739 3780 6743 3836
rect 6743 3780 6799 3836
rect 6799 3780 6803 3836
rect 6739 3776 6803 3780
rect 10432 3836 10496 3840
rect 10432 3780 10436 3836
rect 10436 3780 10492 3836
rect 10492 3780 10496 3836
rect 10432 3776 10496 3780
rect 10512 3836 10576 3840
rect 10512 3780 10516 3836
rect 10516 3780 10572 3836
rect 10572 3780 10576 3836
rect 10512 3776 10576 3780
rect 10592 3836 10656 3840
rect 10592 3780 10596 3836
rect 10596 3780 10652 3836
rect 10652 3780 10656 3836
rect 10592 3776 10656 3780
rect 10672 3836 10736 3840
rect 10672 3780 10676 3836
rect 10676 3780 10732 3836
rect 10732 3780 10736 3836
rect 10672 3776 10736 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 14605 3836 14669 3840
rect 14605 3780 14609 3836
rect 14609 3780 14665 3836
rect 14665 3780 14669 3836
rect 14605 3776 14669 3780
rect 1906 3292 1970 3296
rect 1906 3236 1910 3292
rect 1910 3236 1966 3292
rect 1966 3236 1970 3292
rect 1906 3232 1970 3236
rect 1986 3292 2050 3296
rect 1986 3236 1990 3292
rect 1990 3236 2046 3292
rect 2046 3236 2050 3292
rect 1986 3232 2050 3236
rect 2066 3292 2130 3296
rect 2066 3236 2070 3292
rect 2070 3236 2126 3292
rect 2126 3236 2130 3292
rect 2066 3232 2130 3236
rect 2146 3292 2210 3296
rect 2146 3236 2150 3292
rect 2150 3236 2206 3292
rect 2206 3236 2210 3292
rect 2146 3232 2210 3236
rect 5839 3292 5903 3296
rect 5839 3236 5843 3292
rect 5843 3236 5899 3292
rect 5899 3236 5903 3292
rect 5839 3232 5903 3236
rect 5919 3292 5983 3296
rect 5919 3236 5923 3292
rect 5923 3236 5979 3292
rect 5979 3236 5983 3292
rect 5919 3232 5983 3236
rect 5999 3292 6063 3296
rect 5999 3236 6003 3292
rect 6003 3236 6059 3292
rect 6059 3236 6063 3292
rect 5999 3232 6063 3236
rect 6079 3292 6143 3296
rect 6079 3236 6083 3292
rect 6083 3236 6139 3292
rect 6139 3236 6143 3292
rect 6079 3232 6143 3236
rect 9772 3292 9836 3296
rect 9772 3236 9776 3292
rect 9776 3236 9832 3292
rect 9832 3236 9836 3292
rect 9772 3232 9836 3236
rect 9852 3292 9916 3296
rect 9852 3236 9856 3292
rect 9856 3236 9912 3292
rect 9912 3236 9916 3292
rect 9852 3232 9916 3236
rect 9932 3292 9996 3296
rect 9932 3236 9936 3292
rect 9936 3236 9992 3292
rect 9992 3236 9996 3292
rect 9932 3232 9996 3236
rect 10012 3292 10076 3296
rect 10012 3236 10016 3292
rect 10016 3236 10072 3292
rect 10072 3236 10076 3292
rect 10012 3232 10076 3236
rect 13705 3292 13769 3296
rect 13705 3236 13709 3292
rect 13709 3236 13765 3292
rect 13765 3236 13769 3292
rect 13705 3232 13769 3236
rect 13785 3292 13849 3296
rect 13785 3236 13789 3292
rect 13789 3236 13845 3292
rect 13845 3236 13849 3292
rect 13785 3232 13849 3236
rect 13865 3292 13929 3296
rect 13865 3236 13869 3292
rect 13869 3236 13925 3292
rect 13925 3236 13929 3292
rect 13865 3232 13929 3236
rect 13945 3292 14009 3296
rect 13945 3236 13949 3292
rect 13949 3236 14005 3292
rect 14005 3236 14009 3292
rect 13945 3232 14009 3236
rect 2566 2748 2630 2752
rect 2566 2692 2570 2748
rect 2570 2692 2626 2748
rect 2626 2692 2630 2748
rect 2566 2688 2630 2692
rect 2646 2748 2710 2752
rect 2646 2692 2650 2748
rect 2650 2692 2706 2748
rect 2706 2692 2710 2748
rect 2646 2688 2710 2692
rect 2726 2748 2790 2752
rect 2726 2692 2730 2748
rect 2730 2692 2786 2748
rect 2786 2692 2790 2748
rect 2726 2688 2790 2692
rect 2806 2748 2870 2752
rect 2806 2692 2810 2748
rect 2810 2692 2866 2748
rect 2866 2692 2870 2748
rect 2806 2688 2870 2692
rect 6499 2748 6563 2752
rect 6499 2692 6503 2748
rect 6503 2692 6559 2748
rect 6559 2692 6563 2748
rect 6499 2688 6563 2692
rect 6579 2748 6643 2752
rect 6579 2692 6583 2748
rect 6583 2692 6639 2748
rect 6639 2692 6643 2748
rect 6579 2688 6643 2692
rect 6659 2748 6723 2752
rect 6659 2692 6663 2748
rect 6663 2692 6719 2748
rect 6719 2692 6723 2748
rect 6659 2688 6723 2692
rect 6739 2748 6803 2752
rect 6739 2692 6743 2748
rect 6743 2692 6799 2748
rect 6799 2692 6803 2748
rect 6739 2688 6803 2692
rect 10432 2748 10496 2752
rect 10432 2692 10436 2748
rect 10436 2692 10492 2748
rect 10492 2692 10496 2748
rect 10432 2688 10496 2692
rect 10512 2748 10576 2752
rect 10512 2692 10516 2748
rect 10516 2692 10572 2748
rect 10572 2692 10576 2748
rect 10512 2688 10576 2692
rect 10592 2748 10656 2752
rect 10592 2692 10596 2748
rect 10596 2692 10652 2748
rect 10652 2692 10656 2748
rect 10592 2688 10656 2692
rect 10672 2748 10736 2752
rect 10672 2692 10676 2748
rect 10676 2692 10732 2748
rect 10732 2692 10736 2748
rect 10672 2688 10736 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 14605 2748 14669 2752
rect 14605 2692 14609 2748
rect 14609 2692 14665 2748
rect 14665 2692 14669 2748
rect 14605 2688 14669 2692
rect 1906 2204 1970 2208
rect 1906 2148 1910 2204
rect 1910 2148 1966 2204
rect 1966 2148 1970 2204
rect 1906 2144 1970 2148
rect 1986 2204 2050 2208
rect 1986 2148 1990 2204
rect 1990 2148 2046 2204
rect 2046 2148 2050 2204
rect 1986 2144 2050 2148
rect 2066 2204 2130 2208
rect 2066 2148 2070 2204
rect 2070 2148 2126 2204
rect 2126 2148 2130 2204
rect 2066 2144 2130 2148
rect 2146 2204 2210 2208
rect 2146 2148 2150 2204
rect 2150 2148 2206 2204
rect 2206 2148 2210 2204
rect 2146 2144 2210 2148
rect 5839 2204 5903 2208
rect 5839 2148 5843 2204
rect 5843 2148 5899 2204
rect 5899 2148 5903 2204
rect 5839 2144 5903 2148
rect 5919 2204 5983 2208
rect 5919 2148 5923 2204
rect 5923 2148 5979 2204
rect 5979 2148 5983 2204
rect 5919 2144 5983 2148
rect 5999 2204 6063 2208
rect 5999 2148 6003 2204
rect 6003 2148 6059 2204
rect 6059 2148 6063 2204
rect 5999 2144 6063 2148
rect 6079 2204 6143 2208
rect 6079 2148 6083 2204
rect 6083 2148 6139 2204
rect 6139 2148 6143 2204
rect 6079 2144 6143 2148
rect 9772 2204 9836 2208
rect 9772 2148 9776 2204
rect 9776 2148 9832 2204
rect 9832 2148 9836 2204
rect 9772 2144 9836 2148
rect 9852 2204 9916 2208
rect 9852 2148 9856 2204
rect 9856 2148 9912 2204
rect 9912 2148 9916 2204
rect 9852 2144 9916 2148
rect 9932 2204 9996 2208
rect 9932 2148 9936 2204
rect 9936 2148 9992 2204
rect 9992 2148 9996 2204
rect 9932 2144 9996 2148
rect 10012 2204 10076 2208
rect 10012 2148 10016 2204
rect 10016 2148 10072 2204
rect 10072 2148 10076 2204
rect 10012 2144 10076 2148
rect 13705 2204 13769 2208
rect 13705 2148 13709 2204
rect 13709 2148 13765 2204
rect 13765 2148 13769 2204
rect 13705 2144 13769 2148
rect 13785 2204 13849 2208
rect 13785 2148 13789 2204
rect 13789 2148 13845 2204
rect 13845 2148 13849 2204
rect 13785 2144 13849 2148
rect 13865 2204 13929 2208
rect 13865 2148 13869 2204
rect 13869 2148 13925 2204
rect 13925 2148 13929 2204
rect 13865 2144 13929 2148
rect 13945 2204 14009 2208
rect 13945 2148 13949 2204
rect 13949 2148 14005 2204
rect 14005 2148 14009 2204
rect 13945 2144 14009 2148
rect 2566 1660 2630 1664
rect 2566 1604 2570 1660
rect 2570 1604 2626 1660
rect 2626 1604 2630 1660
rect 2566 1600 2630 1604
rect 2646 1660 2710 1664
rect 2646 1604 2650 1660
rect 2650 1604 2706 1660
rect 2706 1604 2710 1660
rect 2646 1600 2710 1604
rect 2726 1660 2790 1664
rect 2726 1604 2730 1660
rect 2730 1604 2786 1660
rect 2786 1604 2790 1660
rect 2726 1600 2790 1604
rect 2806 1660 2870 1664
rect 2806 1604 2810 1660
rect 2810 1604 2866 1660
rect 2866 1604 2870 1660
rect 2806 1600 2870 1604
rect 6499 1660 6563 1664
rect 6499 1604 6503 1660
rect 6503 1604 6559 1660
rect 6559 1604 6563 1660
rect 6499 1600 6563 1604
rect 6579 1660 6643 1664
rect 6579 1604 6583 1660
rect 6583 1604 6639 1660
rect 6639 1604 6643 1660
rect 6579 1600 6643 1604
rect 6659 1660 6723 1664
rect 6659 1604 6663 1660
rect 6663 1604 6719 1660
rect 6719 1604 6723 1660
rect 6659 1600 6723 1604
rect 6739 1660 6803 1664
rect 6739 1604 6743 1660
rect 6743 1604 6799 1660
rect 6799 1604 6803 1660
rect 6739 1600 6803 1604
rect 10432 1660 10496 1664
rect 10432 1604 10436 1660
rect 10436 1604 10492 1660
rect 10492 1604 10496 1660
rect 10432 1600 10496 1604
rect 10512 1660 10576 1664
rect 10512 1604 10516 1660
rect 10516 1604 10572 1660
rect 10572 1604 10576 1660
rect 10512 1600 10576 1604
rect 10592 1660 10656 1664
rect 10592 1604 10596 1660
rect 10596 1604 10652 1660
rect 10652 1604 10656 1660
rect 10592 1600 10656 1604
rect 10672 1660 10736 1664
rect 10672 1604 10676 1660
rect 10676 1604 10732 1660
rect 10732 1604 10736 1660
rect 10672 1600 10736 1604
rect 14365 1660 14429 1664
rect 14365 1604 14369 1660
rect 14369 1604 14425 1660
rect 14425 1604 14429 1660
rect 14365 1600 14429 1604
rect 14445 1660 14509 1664
rect 14445 1604 14449 1660
rect 14449 1604 14505 1660
rect 14505 1604 14509 1660
rect 14445 1600 14509 1604
rect 14525 1660 14589 1664
rect 14525 1604 14529 1660
rect 14529 1604 14585 1660
rect 14585 1604 14589 1660
rect 14525 1600 14589 1604
rect 14605 1660 14669 1664
rect 14605 1604 14609 1660
rect 14609 1604 14665 1660
rect 14665 1604 14669 1660
rect 14605 1600 14669 1604
rect 1906 1116 1970 1120
rect 1906 1060 1910 1116
rect 1910 1060 1966 1116
rect 1966 1060 1970 1116
rect 1906 1056 1970 1060
rect 1986 1116 2050 1120
rect 1986 1060 1990 1116
rect 1990 1060 2046 1116
rect 2046 1060 2050 1116
rect 1986 1056 2050 1060
rect 2066 1116 2130 1120
rect 2066 1060 2070 1116
rect 2070 1060 2126 1116
rect 2126 1060 2130 1116
rect 2066 1056 2130 1060
rect 2146 1116 2210 1120
rect 2146 1060 2150 1116
rect 2150 1060 2206 1116
rect 2206 1060 2210 1116
rect 2146 1056 2210 1060
rect 5839 1116 5903 1120
rect 5839 1060 5843 1116
rect 5843 1060 5899 1116
rect 5899 1060 5903 1116
rect 5839 1056 5903 1060
rect 5919 1116 5983 1120
rect 5919 1060 5923 1116
rect 5923 1060 5979 1116
rect 5979 1060 5983 1116
rect 5919 1056 5983 1060
rect 5999 1116 6063 1120
rect 5999 1060 6003 1116
rect 6003 1060 6059 1116
rect 6059 1060 6063 1116
rect 5999 1056 6063 1060
rect 6079 1116 6143 1120
rect 6079 1060 6083 1116
rect 6083 1060 6139 1116
rect 6139 1060 6143 1116
rect 6079 1056 6143 1060
rect 9772 1116 9836 1120
rect 9772 1060 9776 1116
rect 9776 1060 9832 1116
rect 9832 1060 9836 1116
rect 9772 1056 9836 1060
rect 9852 1116 9916 1120
rect 9852 1060 9856 1116
rect 9856 1060 9912 1116
rect 9912 1060 9916 1116
rect 9852 1056 9916 1060
rect 9932 1116 9996 1120
rect 9932 1060 9936 1116
rect 9936 1060 9992 1116
rect 9992 1060 9996 1116
rect 9932 1056 9996 1060
rect 10012 1116 10076 1120
rect 10012 1060 10016 1116
rect 10016 1060 10072 1116
rect 10072 1060 10076 1116
rect 10012 1056 10076 1060
rect 13705 1116 13769 1120
rect 13705 1060 13709 1116
rect 13709 1060 13765 1116
rect 13765 1060 13769 1116
rect 13705 1056 13769 1060
rect 13785 1116 13849 1120
rect 13785 1060 13789 1116
rect 13789 1060 13845 1116
rect 13845 1060 13849 1116
rect 13785 1056 13849 1060
rect 13865 1116 13929 1120
rect 13865 1060 13869 1116
rect 13869 1060 13925 1116
rect 13925 1060 13929 1116
rect 13865 1056 13929 1060
rect 13945 1116 14009 1120
rect 13945 1060 13949 1116
rect 13949 1060 14005 1116
rect 14005 1060 14009 1116
rect 13945 1056 14009 1060
rect 2566 572 2630 576
rect 2566 516 2570 572
rect 2570 516 2626 572
rect 2626 516 2630 572
rect 2566 512 2630 516
rect 2646 572 2710 576
rect 2646 516 2650 572
rect 2650 516 2706 572
rect 2706 516 2710 572
rect 2646 512 2710 516
rect 2726 572 2790 576
rect 2726 516 2730 572
rect 2730 516 2786 572
rect 2786 516 2790 572
rect 2726 512 2790 516
rect 2806 572 2870 576
rect 2806 516 2810 572
rect 2810 516 2866 572
rect 2866 516 2870 572
rect 2806 512 2870 516
rect 6499 572 6563 576
rect 6499 516 6503 572
rect 6503 516 6559 572
rect 6559 516 6563 572
rect 6499 512 6563 516
rect 6579 572 6643 576
rect 6579 516 6583 572
rect 6583 516 6639 572
rect 6639 516 6643 572
rect 6579 512 6643 516
rect 6659 572 6723 576
rect 6659 516 6663 572
rect 6663 516 6719 572
rect 6719 516 6723 572
rect 6659 512 6723 516
rect 6739 572 6803 576
rect 6739 516 6743 572
rect 6743 516 6799 572
rect 6799 516 6803 572
rect 6739 512 6803 516
rect 10432 572 10496 576
rect 10432 516 10436 572
rect 10436 516 10492 572
rect 10492 516 10496 572
rect 10432 512 10496 516
rect 10512 572 10576 576
rect 10512 516 10516 572
rect 10516 516 10572 572
rect 10572 516 10576 572
rect 10512 512 10576 516
rect 10592 572 10656 576
rect 10592 516 10596 572
rect 10596 516 10652 572
rect 10652 516 10656 572
rect 10592 512 10656 516
rect 10672 572 10736 576
rect 10672 516 10676 572
rect 10676 516 10732 572
rect 10732 516 10736 572
rect 10672 512 10736 516
rect 14365 572 14429 576
rect 14365 516 14369 572
rect 14369 516 14425 572
rect 14425 516 14429 572
rect 14365 512 14429 516
rect 14445 572 14509 576
rect 14445 516 14449 572
rect 14449 516 14505 572
rect 14505 516 14509 572
rect 14445 512 14509 516
rect 14525 572 14589 576
rect 14525 516 14529 572
rect 14529 516 14585 572
rect 14585 516 14589 572
rect 14525 512 14589 516
rect 14605 572 14669 576
rect 14605 516 14609 572
rect 14609 516 14665 572
rect 14665 516 14669 572
rect 14605 512 14669 516
<< metal4 >>
rect 1898 13088 2218 13104
rect 1898 13024 1906 13088
rect 1970 13024 1986 13088
rect 2050 13024 2066 13088
rect 2130 13024 2146 13088
rect 2210 13024 2218 13088
rect 1898 12000 2218 13024
rect 1898 11936 1906 12000
rect 1970 11936 1986 12000
rect 2050 11936 2066 12000
rect 2130 11936 2146 12000
rect 2210 11936 2218 12000
rect 1898 11610 2218 11936
rect 1898 11374 1940 11610
rect 2176 11374 2218 11610
rect 1898 10912 2218 11374
rect 1898 10848 1906 10912
rect 1970 10848 1986 10912
rect 2050 10848 2066 10912
rect 2130 10848 2146 10912
rect 2210 10848 2218 10912
rect 1898 9824 2218 10848
rect 1898 9760 1906 9824
rect 1970 9760 1986 9824
rect 2050 9760 2066 9824
rect 2130 9760 2146 9824
rect 2210 9760 2218 9824
rect 1898 8736 2218 9760
rect 1898 8672 1906 8736
rect 1970 8672 1986 8736
rect 2050 8672 2066 8736
rect 2130 8672 2146 8736
rect 2210 8672 2218 8736
rect 1898 8482 2218 8672
rect 1898 8246 1940 8482
rect 2176 8246 2218 8482
rect 1898 7648 2218 8246
rect 1898 7584 1906 7648
rect 1970 7584 1986 7648
rect 2050 7584 2066 7648
rect 2130 7584 2146 7648
rect 2210 7584 2218 7648
rect 1898 6560 2218 7584
rect 1898 6496 1906 6560
rect 1970 6496 1986 6560
rect 2050 6496 2066 6560
rect 2130 6496 2146 6560
rect 2210 6496 2218 6560
rect 1898 5472 2218 6496
rect 1898 5408 1906 5472
rect 1970 5408 1986 5472
rect 2050 5408 2066 5472
rect 2130 5408 2146 5472
rect 2210 5408 2218 5472
rect 1898 5354 2218 5408
rect 1898 5118 1940 5354
rect 2176 5118 2218 5354
rect 1898 4384 2218 5118
rect 1898 4320 1906 4384
rect 1970 4320 1986 4384
rect 2050 4320 2066 4384
rect 2130 4320 2146 4384
rect 2210 4320 2218 4384
rect 1898 3296 2218 4320
rect 1898 3232 1906 3296
rect 1970 3232 1986 3296
rect 2050 3232 2066 3296
rect 2130 3232 2146 3296
rect 2210 3232 2218 3296
rect 1898 2226 2218 3232
rect 1898 2208 1940 2226
rect 2176 2208 2218 2226
rect 1898 2144 1906 2208
rect 2210 2144 2218 2208
rect 1898 1990 1940 2144
rect 2176 1990 2218 2144
rect 1898 1120 2218 1990
rect 1898 1056 1906 1120
rect 1970 1056 1986 1120
rect 2050 1056 2066 1120
rect 2130 1056 2146 1120
rect 2210 1056 2218 1120
rect 1898 496 2218 1056
rect 2558 12544 2878 13104
rect 2558 12480 2566 12544
rect 2630 12480 2646 12544
rect 2710 12480 2726 12544
rect 2790 12480 2806 12544
rect 2870 12480 2878 12544
rect 2558 12270 2878 12480
rect 2558 12034 2600 12270
rect 2836 12034 2878 12270
rect 2558 11456 2878 12034
rect 2558 11392 2566 11456
rect 2630 11392 2646 11456
rect 2710 11392 2726 11456
rect 2790 11392 2806 11456
rect 2870 11392 2878 11456
rect 2558 10368 2878 11392
rect 2558 10304 2566 10368
rect 2630 10304 2646 10368
rect 2710 10304 2726 10368
rect 2790 10304 2806 10368
rect 2870 10304 2878 10368
rect 2558 9280 2878 10304
rect 2558 9216 2566 9280
rect 2630 9216 2646 9280
rect 2710 9216 2726 9280
rect 2790 9216 2806 9280
rect 2870 9216 2878 9280
rect 2558 9142 2878 9216
rect 2558 8906 2600 9142
rect 2836 8906 2878 9142
rect 2558 8192 2878 8906
rect 2558 8128 2566 8192
rect 2630 8128 2646 8192
rect 2710 8128 2726 8192
rect 2790 8128 2806 8192
rect 2870 8128 2878 8192
rect 2558 7104 2878 8128
rect 2558 7040 2566 7104
rect 2630 7040 2646 7104
rect 2710 7040 2726 7104
rect 2790 7040 2806 7104
rect 2870 7040 2878 7104
rect 2558 6016 2878 7040
rect 2558 5952 2566 6016
rect 2630 6014 2646 6016
rect 2710 6014 2726 6016
rect 2790 6014 2806 6016
rect 2870 5952 2878 6016
rect 2558 5778 2600 5952
rect 2836 5778 2878 5952
rect 2558 4928 2878 5778
rect 2558 4864 2566 4928
rect 2630 4864 2646 4928
rect 2710 4864 2726 4928
rect 2790 4864 2806 4928
rect 2870 4864 2878 4928
rect 2558 3840 2878 4864
rect 2558 3776 2566 3840
rect 2630 3776 2646 3840
rect 2710 3776 2726 3840
rect 2790 3776 2806 3840
rect 2870 3776 2878 3840
rect 2558 2886 2878 3776
rect 2558 2752 2600 2886
rect 2836 2752 2878 2886
rect 2558 2688 2566 2752
rect 2870 2688 2878 2752
rect 2558 2650 2600 2688
rect 2836 2650 2878 2688
rect 2558 1664 2878 2650
rect 2558 1600 2566 1664
rect 2630 1600 2646 1664
rect 2710 1600 2726 1664
rect 2790 1600 2806 1664
rect 2870 1600 2878 1664
rect 2558 576 2878 1600
rect 2558 512 2566 576
rect 2630 512 2646 576
rect 2710 512 2726 576
rect 2790 512 2806 576
rect 2870 512 2878 576
rect 2558 496 2878 512
rect 5831 13088 6151 13104
rect 5831 13024 5839 13088
rect 5903 13024 5919 13088
rect 5983 13024 5999 13088
rect 6063 13024 6079 13088
rect 6143 13024 6151 13088
rect 5831 12000 6151 13024
rect 5831 11936 5839 12000
rect 5903 11936 5919 12000
rect 5983 11936 5999 12000
rect 6063 11936 6079 12000
rect 6143 11936 6151 12000
rect 5831 11610 6151 11936
rect 5831 11374 5873 11610
rect 6109 11374 6151 11610
rect 5831 10912 6151 11374
rect 5831 10848 5839 10912
rect 5903 10848 5919 10912
rect 5983 10848 5999 10912
rect 6063 10848 6079 10912
rect 6143 10848 6151 10912
rect 5831 9824 6151 10848
rect 5831 9760 5839 9824
rect 5903 9760 5919 9824
rect 5983 9760 5999 9824
rect 6063 9760 6079 9824
rect 6143 9760 6151 9824
rect 5831 8736 6151 9760
rect 5831 8672 5839 8736
rect 5903 8672 5919 8736
rect 5983 8672 5999 8736
rect 6063 8672 6079 8736
rect 6143 8672 6151 8736
rect 5831 8482 6151 8672
rect 5831 8246 5873 8482
rect 6109 8246 6151 8482
rect 5831 7648 6151 8246
rect 5831 7584 5839 7648
rect 5903 7584 5919 7648
rect 5983 7584 5999 7648
rect 6063 7584 6079 7648
rect 6143 7584 6151 7648
rect 5831 6560 6151 7584
rect 5831 6496 5839 6560
rect 5903 6496 5919 6560
rect 5983 6496 5999 6560
rect 6063 6496 6079 6560
rect 6143 6496 6151 6560
rect 5831 5472 6151 6496
rect 5831 5408 5839 5472
rect 5903 5408 5919 5472
rect 5983 5408 5999 5472
rect 6063 5408 6079 5472
rect 6143 5408 6151 5472
rect 5831 5354 6151 5408
rect 5831 5118 5873 5354
rect 6109 5118 6151 5354
rect 5831 4384 6151 5118
rect 5831 4320 5839 4384
rect 5903 4320 5919 4384
rect 5983 4320 5999 4384
rect 6063 4320 6079 4384
rect 6143 4320 6151 4384
rect 5831 3296 6151 4320
rect 5831 3232 5839 3296
rect 5903 3232 5919 3296
rect 5983 3232 5999 3296
rect 6063 3232 6079 3296
rect 6143 3232 6151 3296
rect 5831 2226 6151 3232
rect 5831 2208 5873 2226
rect 6109 2208 6151 2226
rect 5831 2144 5839 2208
rect 6143 2144 6151 2208
rect 5831 1990 5873 2144
rect 6109 1990 6151 2144
rect 5831 1120 6151 1990
rect 5831 1056 5839 1120
rect 5903 1056 5919 1120
rect 5983 1056 5999 1120
rect 6063 1056 6079 1120
rect 6143 1056 6151 1120
rect 5831 496 6151 1056
rect 6491 12544 6811 13104
rect 6491 12480 6499 12544
rect 6563 12480 6579 12544
rect 6643 12480 6659 12544
rect 6723 12480 6739 12544
rect 6803 12480 6811 12544
rect 6491 12270 6811 12480
rect 6491 12034 6533 12270
rect 6769 12034 6811 12270
rect 6491 11456 6811 12034
rect 6491 11392 6499 11456
rect 6563 11392 6579 11456
rect 6643 11392 6659 11456
rect 6723 11392 6739 11456
rect 6803 11392 6811 11456
rect 6491 10368 6811 11392
rect 6491 10304 6499 10368
rect 6563 10304 6579 10368
rect 6643 10304 6659 10368
rect 6723 10304 6739 10368
rect 6803 10304 6811 10368
rect 6491 9280 6811 10304
rect 6491 9216 6499 9280
rect 6563 9216 6579 9280
rect 6643 9216 6659 9280
rect 6723 9216 6739 9280
rect 6803 9216 6811 9280
rect 6491 9142 6811 9216
rect 6491 8906 6533 9142
rect 6769 8906 6811 9142
rect 6491 8192 6811 8906
rect 6491 8128 6499 8192
rect 6563 8128 6579 8192
rect 6643 8128 6659 8192
rect 6723 8128 6739 8192
rect 6803 8128 6811 8192
rect 6491 7104 6811 8128
rect 6491 7040 6499 7104
rect 6563 7040 6579 7104
rect 6643 7040 6659 7104
rect 6723 7040 6739 7104
rect 6803 7040 6811 7104
rect 6491 6016 6811 7040
rect 6491 5952 6499 6016
rect 6563 6014 6579 6016
rect 6643 6014 6659 6016
rect 6723 6014 6739 6016
rect 6803 5952 6811 6016
rect 6491 5778 6533 5952
rect 6769 5778 6811 5952
rect 6491 4928 6811 5778
rect 6491 4864 6499 4928
rect 6563 4864 6579 4928
rect 6643 4864 6659 4928
rect 6723 4864 6739 4928
rect 6803 4864 6811 4928
rect 6491 3840 6811 4864
rect 6491 3776 6499 3840
rect 6563 3776 6579 3840
rect 6643 3776 6659 3840
rect 6723 3776 6739 3840
rect 6803 3776 6811 3840
rect 6491 2886 6811 3776
rect 6491 2752 6533 2886
rect 6769 2752 6811 2886
rect 6491 2688 6499 2752
rect 6803 2688 6811 2752
rect 6491 2650 6533 2688
rect 6769 2650 6811 2688
rect 6491 1664 6811 2650
rect 6491 1600 6499 1664
rect 6563 1600 6579 1664
rect 6643 1600 6659 1664
rect 6723 1600 6739 1664
rect 6803 1600 6811 1664
rect 6491 576 6811 1600
rect 6491 512 6499 576
rect 6563 512 6579 576
rect 6643 512 6659 576
rect 6723 512 6739 576
rect 6803 512 6811 576
rect 6491 496 6811 512
rect 9764 13088 10084 13104
rect 9764 13024 9772 13088
rect 9836 13024 9852 13088
rect 9916 13024 9932 13088
rect 9996 13024 10012 13088
rect 10076 13024 10084 13088
rect 9764 12000 10084 13024
rect 9764 11936 9772 12000
rect 9836 11936 9852 12000
rect 9916 11936 9932 12000
rect 9996 11936 10012 12000
rect 10076 11936 10084 12000
rect 9764 11610 10084 11936
rect 9764 11374 9806 11610
rect 10042 11374 10084 11610
rect 9764 10912 10084 11374
rect 9764 10848 9772 10912
rect 9836 10848 9852 10912
rect 9916 10848 9932 10912
rect 9996 10848 10012 10912
rect 10076 10848 10084 10912
rect 9764 9824 10084 10848
rect 9764 9760 9772 9824
rect 9836 9760 9852 9824
rect 9916 9760 9932 9824
rect 9996 9760 10012 9824
rect 10076 9760 10084 9824
rect 9764 8736 10084 9760
rect 9764 8672 9772 8736
rect 9836 8672 9852 8736
rect 9916 8672 9932 8736
rect 9996 8672 10012 8736
rect 10076 8672 10084 8736
rect 9764 8482 10084 8672
rect 9764 8246 9806 8482
rect 10042 8246 10084 8482
rect 9764 7648 10084 8246
rect 9764 7584 9772 7648
rect 9836 7584 9852 7648
rect 9916 7584 9932 7648
rect 9996 7584 10012 7648
rect 10076 7584 10084 7648
rect 9764 6560 10084 7584
rect 9764 6496 9772 6560
rect 9836 6496 9852 6560
rect 9916 6496 9932 6560
rect 9996 6496 10012 6560
rect 10076 6496 10084 6560
rect 9764 5472 10084 6496
rect 9764 5408 9772 5472
rect 9836 5408 9852 5472
rect 9916 5408 9932 5472
rect 9996 5408 10012 5472
rect 10076 5408 10084 5472
rect 9764 5354 10084 5408
rect 9764 5118 9806 5354
rect 10042 5118 10084 5354
rect 9764 4384 10084 5118
rect 9764 4320 9772 4384
rect 9836 4320 9852 4384
rect 9916 4320 9932 4384
rect 9996 4320 10012 4384
rect 10076 4320 10084 4384
rect 9764 3296 10084 4320
rect 9764 3232 9772 3296
rect 9836 3232 9852 3296
rect 9916 3232 9932 3296
rect 9996 3232 10012 3296
rect 10076 3232 10084 3296
rect 9764 2226 10084 3232
rect 9764 2208 9806 2226
rect 10042 2208 10084 2226
rect 9764 2144 9772 2208
rect 10076 2144 10084 2208
rect 9764 1990 9806 2144
rect 10042 1990 10084 2144
rect 9764 1120 10084 1990
rect 9764 1056 9772 1120
rect 9836 1056 9852 1120
rect 9916 1056 9932 1120
rect 9996 1056 10012 1120
rect 10076 1056 10084 1120
rect 9764 496 10084 1056
rect 10424 12544 10744 13104
rect 10424 12480 10432 12544
rect 10496 12480 10512 12544
rect 10576 12480 10592 12544
rect 10656 12480 10672 12544
rect 10736 12480 10744 12544
rect 10424 12270 10744 12480
rect 10424 12034 10466 12270
rect 10702 12034 10744 12270
rect 10424 11456 10744 12034
rect 10424 11392 10432 11456
rect 10496 11392 10512 11456
rect 10576 11392 10592 11456
rect 10656 11392 10672 11456
rect 10736 11392 10744 11456
rect 10424 10368 10744 11392
rect 10424 10304 10432 10368
rect 10496 10304 10512 10368
rect 10576 10304 10592 10368
rect 10656 10304 10672 10368
rect 10736 10304 10744 10368
rect 10424 9280 10744 10304
rect 10424 9216 10432 9280
rect 10496 9216 10512 9280
rect 10576 9216 10592 9280
rect 10656 9216 10672 9280
rect 10736 9216 10744 9280
rect 10424 9142 10744 9216
rect 10424 8906 10466 9142
rect 10702 8906 10744 9142
rect 10424 8192 10744 8906
rect 10424 8128 10432 8192
rect 10496 8128 10512 8192
rect 10576 8128 10592 8192
rect 10656 8128 10672 8192
rect 10736 8128 10744 8192
rect 10424 7104 10744 8128
rect 10424 7040 10432 7104
rect 10496 7040 10512 7104
rect 10576 7040 10592 7104
rect 10656 7040 10672 7104
rect 10736 7040 10744 7104
rect 10424 6016 10744 7040
rect 10424 5952 10432 6016
rect 10496 6014 10512 6016
rect 10576 6014 10592 6016
rect 10656 6014 10672 6016
rect 10736 5952 10744 6016
rect 10424 5778 10466 5952
rect 10702 5778 10744 5952
rect 10424 4928 10744 5778
rect 10424 4864 10432 4928
rect 10496 4864 10512 4928
rect 10576 4864 10592 4928
rect 10656 4864 10672 4928
rect 10736 4864 10744 4928
rect 10424 3840 10744 4864
rect 10424 3776 10432 3840
rect 10496 3776 10512 3840
rect 10576 3776 10592 3840
rect 10656 3776 10672 3840
rect 10736 3776 10744 3840
rect 10424 2886 10744 3776
rect 10424 2752 10466 2886
rect 10702 2752 10744 2886
rect 10424 2688 10432 2752
rect 10736 2688 10744 2752
rect 10424 2650 10466 2688
rect 10702 2650 10744 2688
rect 10424 1664 10744 2650
rect 10424 1600 10432 1664
rect 10496 1600 10512 1664
rect 10576 1600 10592 1664
rect 10656 1600 10672 1664
rect 10736 1600 10744 1664
rect 10424 576 10744 1600
rect 10424 512 10432 576
rect 10496 512 10512 576
rect 10576 512 10592 576
rect 10656 512 10672 576
rect 10736 512 10744 576
rect 10424 496 10744 512
rect 13697 13088 14017 13104
rect 13697 13024 13705 13088
rect 13769 13024 13785 13088
rect 13849 13024 13865 13088
rect 13929 13024 13945 13088
rect 14009 13024 14017 13088
rect 13697 12000 14017 13024
rect 13697 11936 13705 12000
rect 13769 11936 13785 12000
rect 13849 11936 13865 12000
rect 13929 11936 13945 12000
rect 14009 11936 14017 12000
rect 13697 11610 14017 11936
rect 13697 11374 13739 11610
rect 13975 11374 14017 11610
rect 13697 10912 14017 11374
rect 13697 10848 13705 10912
rect 13769 10848 13785 10912
rect 13849 10848 13865 10912
rect 13929 10848 13945 10912
rect 14009 10848 14017 10912
rect 13697 9824 14017 10848
rect 13697 9760 13705 9824
rect 13769 9760 13785 9824
rect 13849 9760 13865 9824
rect 13929 9760 13945 9824
rect 14009 9760 14017 9824
rect 13697 8736 14017 9760
rect 13697 8672 13705 8736
rect 13769 8672 13785 8736
rect 13849 8672 13865 8736
rect 13929 8672 13945 8736
rect 14009 8672 14017 8736
rect 13697 8482 14017 8672
rect 13697 8246 13739 8482
rect 13975 8246 14017 8482
rect 13697 7648 14017 8246
rect 13697 7584 13705 7648
rect 13769 7584 13785 7648
rect 13849 7584 13865 7648
rect 13929 7584 13945 7648
rect 14009 7584 14017 7648
rect 13697 6560 14017 7584
rect 13697 6496 13705 6560
rect 13769 6496 13785 6560
rect 13849 6496 13865 6560
rect 13929 6496 13945 6560
rect 14009 6496 14017 6560
rect 13697 5472 14017 6496
rect 13697 5408 13705 5472
rect 13769 5408 13785 5472
rect 13849 5408 13865 5472
rect 13929 5408 13945 5472
rect 14009 5408 14017 5472
rect 13697 5354 14017 5408
rect 13697 5118 13739 5354
rect 13975 5118 14017 5354
rect 13697 4384 14017 5118
rect 13697 4320 13705 4384
rect 13769 4320 13785 4384
rect 13849 4320 13865 4384
rect 13929 4320 13945 4384
rect 14009 4320 14017 4384
rect 13697 3296 14017 4320
rect 13697 3232 13705 3296
rect 13769 3232 13785 3296
rect 13849 3232 13865 3296
rect 13929 3232 13945 3296
rect 14009 3232 14017 3296
rect 13697 2226 14017 3232
rect 13697 2208 13739 2226
rect 13975 2208 14017 2226
rect 13697 2144 13705 2208
rect 14009 2144 14017 2208
rect 13697 1990 13739 2144
rect 13975 1990 14017 2144
rect 13697 1120 14017 1990
rect 13697 1056 13705 1120
rect 13769 1056 13785 1120
rect 13849 1056 13865 1120
rect 13929 1056 13945 1120
rect 14009 1056 14017 1120
rect 13697 496 14017 1056
rect 14357 12544 14677 13104
rect 14357 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14605 12544
rect 14669 12480 14677 12544
rect 14357 12270 14677 12480
rect 14357 12034 14399 12270
rect 14635 12034 14677 12270
rect 14357 11456 14677 12034
rect 14357 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14605 11456
rect 14669 11392 14677 11456
rect 14357 10368 14677 11392
rect 14357 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14605 10368
rect 14669 10304 14677 10368
rect 14357 9280 14677 10304
rect 14357 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14605 9280
rect 14669 9216 14677 9280
rect 14357 9142 14677 9216
rect 14357 8906 14399 9142
rect 14635 8906 14677 9142
rect 14357 8192 14677 8906
rect 14357 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14605 8192
rect 14669 8128 14677 8192
rect 14357 7104 14677 8128
rect 14357 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14605 7104
rect 14669 7040 14677 7104
rect 14357 6016 14677 7040
rect 14357 5952 14365 6016
rect 14429 6014 14445 6016
rect 14509 6014 14525 6016
rect 14589 6014 14605 6016
rect 14669 5952 14677 6016
rect 14357 5778 14399 5952
rect 14635 5778 14677 5952
rect 14357 4928 14677 5778
rect 14357 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14605 4928
rect 14669 4864 14677 4928
rect 14357 3840 14677 4864
rect 14357 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14605 3840
rect 14669 3776 14677 3840
rect 14357 2886 14677 3776
rect 14357 2752 14399 2886
rect 14635 2752 14677 2886
rect 14357 2688 14365 2752
rect 14669 2688 14677 2752
rect 14357 2650 14399 2688
rect 14635 2650 14677 2688
rect 14357 1664 14677 2650
rect 14357 1600 14365 1664
rect 14429 1600 14445 1664
rect 14509 1600 14525 1664
rect 14589 1600 14605 1664
rect 14669 1600 14677 1664
rect 14357 576 14677 1600
rect 14357 512 14365 576
rect 14429 512 14445 576
rect 14509 512 14525 576
rect 14589 512 14605 576
rect 14669 512 14677 576
rect 14357 496 14677 512
<< via4 >>
rect 1940 11374 2176 11610
rect 1940 8246 2176 8482
rect 1940 5118 2176 5354
rect 1940 2208 2176 2226
rect 1940 2144 1970 2208
rect 1970 2144 1986 2208
rect 1986 2144 2050 2208
rect 2050 2144 2066 2208
rect 2066 2144 2130 2208
rect 2130 2144 2146 2208
rect 2146 2144 2176 2208
rect 1940 1990 2176 2144
rect 2600 12034 2836 12270
rect 2600 8906 2836 9142
rect 2600 5952 2630 6014
rect 2630 5952 2646 6014
rect 2646 5952 2710 6014
rect 2710 5952 2726 6014
rect 2726 5952 2790 6014
rect 2790 5952 2806 6014
rect 2806 5952 2836 6014
rect 2600 5778 2836 5952
rect 2600 2752 2836 2886
rect 2600 2688 2630 2752
rect 2630 2688 2646 2752
rect 2646 2688 2710 2752
rect 2710 2688 2726 2752
rect 2726 2688 2790 2752
rect 2790 2688 2806 2752
rect 2806 2688 2836 2752
rect 2600 2650 2836 2688
rect 5873 11374 6109 11610
rect 5873 8246 6109 8482
rect 5873 5118 6109 5354
rect 5873 2208 6109 2226
rect 5873 2144 5903 2208
rect 5903 2144 5919 2208
rect 5919 2144 5983 2208
rect 5983 2144 5999 2208
rect 5999 2144 6063 2208
rect 6063 2144 6079 2208
rect 6079 2144 6109 2208
rect 5873 1990 6109 2144
rect 6533 12034 6769 12270
rect 6533 8906 6769 9142
rect 6533 5952 6563 6014
rect 6563 5952 6579 6014
rect 6579 5952 6643 6014
rect 6643 5952 6659 6014
rect 6659 5952 6723 6014
rect 6723 5952 6739 6014
rect 6739 5952 6769 6014
rect 6533 5778 6769 5952
rect 6533 2752 6769 2886
rect 6533 2688 6563 2752
rect 6563 2688 6579 2752
rect 6579 2688 6643 2752
rect 6643 2688 6659 2752
rect 6659 2688 6723 2752
rect 6723 2688 6739 2752
rect 6739 2688 6769 2752
rect 6533 2650 6769 2688
rect 9806 11374 10042 11610
rect 9806 8246 10042 8482
rect 9806 5118 10042 5354
rect 9806 2208 10042 2226
rect 9806 2144 9836 2208
rect 9836 2144 9852 2208
rect 9852 2144 9916 2208
rect 9916 2144 9932 2208
rect 9932 2144 9996 2208
rect 9996 2144 10012 2208
rect 10012 2144 10042 2208
rect 9806 1990 10042 2144
rect 10466 12034 10702 12270
rect 10466 8906 10702 9142
rect 10466 5952 10496 6014
rect 10496 5952 10512 6014
rect 10512 5952 10576 6014
rect 10576 5952 10592 6014
rect 10592 5952 10656 6014
rect 10656 5952 10672 6014
rect 10672 5952 10702 6014
rect 10466 5778 10702 5952
rect 10466 2752 10702 2886
rect 10466 2688 10496 2752
rect 10496 2688 10512 2752
rect 10512 2688 10576 2752
rect 10576 2688 10592 2752
rect 10592 2688 10656 2752
rect 10656 2688 10672 2752
rect 10672 2688 10702 2752
rect 10466 2650 10702 2688
rect 13739 11374 13975 11610
rect 13739 8246 13975 8482
rect 13739 5118 13975 5354
rect 13739 2208 13975 2226
rect 13739 2144 13769 2208
rect 13769 2144 13785 2208
rect 13785 2144 13849 2208
rect 13849 2144 13865 2208
rect 13865 2144 13929 2208
rect 13929 2144 13945 2208
rect 13945 2144 13975 2208
rect 13739 1990 13975 2144
rect 14399 12034 14635 12270
rect 14399 8906 14635 9142
rect 14399 5952 14429 6014
rect 14429 5952 14445 6014
rect 14445 5952 14509 6014
rect 14509 5952 14525 6014
rect 14525 5952 14589 6014
rect 14589 5952 14605 6014
rect 14605 5952 14635 6014
rect 14399 5778 14635 5952
rect 14399 2752 14635 2886
rect 14399 2688 14429 2752
rect 14429 2688 14445 2752
rect 14445 2688 14509 2752
rect 14509 2688 14525 2752
rect 14525 2688 14589 2752
rect 14589 2688 14605 2752
rect 14605 2688 14635 2752
rect 14399 2650 14635 2688
<< metal5 >>
rect 44 12270 15872 12312
rect 44 12034 2600 12270
rect 2836 12034 6533 12270
rect 6769 12034 10466 12270
rect 10702 12034 14399 12270
rect 14635 12034 15872 12270
rect 44 11992 15872 12034
rect 44 11610 15872 11652
rect 44 11374 1940 11610
rect 2176 11374 5873 11610
rect 6109 11374 9806 11610
rect 10042 11374 13739 11610
rect 13975 11374 15872 11610
rect 44 11332 15872 11374
rect 44 9142 15872 9184
rect 44 8906 2600 9142
rect 2836 8906 6533 9142
rect 6769 8906 10466 9142
rect 10702 8906 14399 9142
rect 14635 8906 15872 9142
rect 44 8864 15872 8906
rect 44 8482 15872 8524
rect 44 8246 1940 8482
rect 2176 8246 5873 8482
rect 6109 8246 9806 8482
rect 10042 8246 13739 8482
rect 13975 8246 15872 8482
rect 44 8204 15872 8246
rect 44 6014 15872 6056
rect 44 5778 2600 6014
rect 2836 5778 6533 6014
rect 6769 5778 10466 6014
rect 10702 5778 14399 6014
rect 14635 5778 15872 6014
rect 44 5736 15872 5778
rect 44 5354 15872 5396
rect 44 5118 1940 5354
rect 2176 5118 5873 5354
rect 6109 5118 9806 5354
rect 10042 5118 13739 5354
rect 13975 5118 15872 5354
rect 44 5076 15872 5118
rect 44 2886 15872 2928
rect 44 2650 2600 2886
rect 2836 2650 6533 2886
rect 6769 2650 10466 2886
rect 10702 2650 14399 2886
rect 14635 2650 15872 2886
rect 44 2608 15872 2650
rect 44 2226 15872 2268
rect 44 1990 1940 2226
rect 2176 1990 5873 2226
rect 6109 1990 9806 2226
rect 10042 1990 13739 2226
rect 13975 1990 15872 2226
rect 44 1948 15872 1990
use sky130_fd_sc_hd__or2_1  _137_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 2668 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _138_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 1748 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 1472 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _140_
timestamp 1693170804
transform 1 0 2024 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp 1693170804
transform -1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1693170804
transform -1 0 3220 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _143_
timestamp 1693170804
transform 1 0 3772 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _144_
timestamp 1693170804
transform 1 0 13892 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 1693170804
transform 1 0 14352 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _146_
timestamp 1693170804
transform 1 0 2300 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _147_
timestamp 1693170804
transform 1 0 11776 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148_
timestamp 1693170804
transform 1 0 12328 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _149_
timestamp 1693170804
transform 1 0 8924 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _150_
timestamp 1693170804
transform 1 0 9844 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _151_
timestamp 1693170804
transform 1 0 11040 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _152_
timestamp 1693170804
transform 1 0 8004 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _153_
timestamp 1693170804
transform 1 0 8740 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1693170804
transform -1 0 8832 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _155_
timestamp 1693170804
transform 1 0 5428 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _156_
timestamp 1693170804
transform 1 0 6164 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _157_
timestamp 1693170804
transform 1 0 6716 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _158_
timestamp 1693170804
transform 1 0 2760 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _159_
timestamp 1693170804
transform 1 0 4140 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1693170804
transform 1 0 4784 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _161_
timestamp 1693170804
transform 1 0 14904 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _162_
timestamp 1693170804
transform -1 0 15180 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1693170804
transform 1 0 14996 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 4416 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1693170804
transform -1 0 8280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _166_
timestamp 1693170804
transform -1 0 6440 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _167_
timestamp 1693170804
transform 1 0 3772 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 8188 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4600 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 7544 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 7912 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _172_
timestamp 1693170804
transform 1 0 14536 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _173_
timestamp 1693170804
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1693170804
transform -1 0 15456 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _175_
timestamp 1693170804
transform 1 0 14536 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _176_
timestamp 1693170804
transform 1 0 14996 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1693170804
transform -1 0 14996 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _178_
timestamp 1693170804
transform 1 0 11224 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _179_
timestamp 1693170804
transform 1 0 14904 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1693170804
transform -1 0 14996 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _181_
timestamp 1693170804
transform 1 0 10120 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _182_
timestamp 1693170804
transform 1 0 14628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1693170804
transform -1 0 14996 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1693170804
transform 1 0 4968 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _185_
timestamp 1693170804
transform 1 0 4508 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5428 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 14352 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _188_
timestamp 1693170804
transform 1 0 14996 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 8004 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_2  _190_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8280 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9568 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 4784 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _193_
timestamp 1693170804
transform 1 0 11316 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _194_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 10396 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9384 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1693170804
transform -1 0 8924 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _197_
timestamp 1693170804
transform 1 0 9844 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 9844 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9568 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8740 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8004 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 8096 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 6440 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 5888 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5520 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp 1693170804
transform -1 0 6348 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 1693170804
transform 1 0 5980 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 5980 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _210_
timestamp 1693170804
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _211_
timestamp 1693170804
transform -1 0 1288 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _212_
timestamp 1693170804
transform 1 0 1012 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _213_
timestamp 1693170804
transform 1 0 736 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _214_
timestamp 1693170804
transform 1 0 2576 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _215_
timestamp 1693170804
transform -1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _216_
timestamp 1693170804
transform 1 0 1564 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _217_
timestamp 1693170804
transform -1 0 1196 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _218_
timestamp 1693170804
transform -1 0 6348 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _219_
timestamp 1693170804
transform -1 0 5980 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _220_
timestamp 1693170804
transform -1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _221_
timestamp 1693170804
transform -1 0 6348 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _222_
timestamp 1693170804
transform 1 0 3312 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _223_
timestamp 1693170804
transform 1 0 3404 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _224_
timestamp 1693170804
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _225_
timestamp 1693170804
transform -1 0 1288 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5428 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 8096 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _228_
timestamp 1693170804
transform 1 0 6440 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _229_
timestamp 1693170804
transform -1 0 6348 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _230_
timestamp 1693170804
transform 1 0 9384 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _231_
timestamp 1693170804
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 5244 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 828 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _234_
timestamp 1693170804
transform -1 0 3680 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _235_
timestamp 1693170804
transform 1 0 4784 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _236_
timestamp 1693170804
transform -1 0 4876 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _237_
timestamp 1693170804
transform 1 0 3312 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1693170804
transform 1 0 2208 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_2  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 7176 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _240_
timestamp 1693170804
transform -1 0 6348 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _241_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 2760 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _242_
timestamp 1693170804
transform 1 0 6440 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _243_
timestamp 1693170804
transform -1 0 5060 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _244_
timestamp 1693170804
transform 1 0 5336 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _245_
timestamp 1693170804
transform 1 0 2116 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _246_
timestamp 1693170804
transform 1 0 2944 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _247_
timestamp 1693170804
transform -1 0 3404 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _248_
timestamp 1693170804
transform -1 0 5244 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _249_
timestamp 1693170804
transform 1 0 6072 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _250_
timestamp 1693170804
transform 1 0 5888 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _251_
timestamp 1693170804
transform 1 0 2760 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1693170804
transform -1 0 2760 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _253_
timestamp 1693170804
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _254_
timestamp 1693170804
transform -1 0 7544 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8280 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _256_
timestamp 1693170804
transform 1 0 10948 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _257_
timestamp 1693170804
transform 1 0 10672 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _258_
timestamp 1693170804
transform 1 0 11040 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _259_
timestamp 1693170804
transform -1 0 11132 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _260_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 7636 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _261_
timestamp 1693170804
transform -1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8280 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _263_
timestamp 1693170804
transform -1 0 5888 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9476 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _265_
timestamp 1693170804
transform 1 0 13616 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _266_
timestamp 1693170804
transform 1 0 9016 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _267_
timestamp 1693170804
transform -1 0 13432 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp 1693170804
transform -1 0 12972 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _269_
timestamp 1693170804
transform 1 0 13800 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _270_
timestamp 1693170804
transform -1 0 13892 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp 1693170804
transform -1 0 13432 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _272_
timestamp 1693170804
transform 1 0 13800 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _273_
timestamp 1693170804
transform 1 0 13248 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1693170804
transform 1 0 13340 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _275_
timestamp 1693170804
transform 1 0 10488 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _276_
timestamp 1693170804
transform 1 0 9660 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1693170804
transform 1 0 10120 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _278_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 10396 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_4  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 10028 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp 1693170804
transform 1 0 10580 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 3864 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _282_
timestamp 1693170804
transform 1 0 3680 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _283_
timestamp 1693170804
transform -1 0 4416 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _284_
timestamp 1693170804
transform 1 0 10948 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _285_
timestamp 1693170804
transform 1 0 10764 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _286_
timestamp 1693170804
transform 1 0 11040 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _287_
timestamp 1693170804
transform 1 0 10672 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _288_
timestamp 1693170804
transform -1 0 15180 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _289_
timestamp 1693170804
transform 1 0 14168 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _290_
timestamp 1693170804
transform -1 0 15456 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 14904 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 13064 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _293_
timestamp 1693170804
transform 1 0 14168 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _294_
timestamp 1693170804
transform 1 0 14720 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _295_
timestamp 1693170804
transform 1 0 13708 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _296_
timestamp 1693170804
transform -1 0 15456 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _297_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 14904 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _298_
timestamp 1693170804
transform 1 0 13064 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 14720 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _300_
timestamp 1693170804
transform 1 0 13064 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _301_
timestamp 1693170804
transform -1 0 14352 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _302_
timestamp 1693170804
transform 1 0 10672 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_2  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8188 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 12144 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _305_
timestamp 1693170804
transform 1 0 6808 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _306_
timestamp 1693170804
transform 1 0 5980 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _307_
timestamp 1693170804
transform 1 0 368 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _308_
timestamp 1693170804
transform 1 0 368 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _309_
timestamp 1693170804
transform 1 0 736 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _310_
timestamp 1693170804
transform 1 0 368 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _311_
timestamp 1693170804
transform 1 0 6440 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _312_
timestamp 1693170804
transform 1 0 6348 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _313_
timestamp 1693170804
transform 1 0 3404 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _314_
timestamp 1693170804
transform 1 0 552 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _315_
timestamp 1693170804
transform 1 0 368 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _316_
timestamp 1693170804
transform 1 0 1840 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _317_
timestamp 1693170804
transform 1 0 2116 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _318_
timestamp 1693170804
transform 1 0 4416 0 1 1632
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _319_
timestamp 1693170804
transform 1 0 2760 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _320_
timestamp 1693170804
transform 1 0 3588 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _321_
timestamp 1693170804
transform 1 0 2760 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 1693170804
transform 1 0 4416 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _323_
timestamp 1693170804
transform 1 0 7912 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _324_
timestamp 1693170804
transform 1 0 6716 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _325_
timestamp 1693170804
transform 1 0 3404 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1693170804
transform 1 0 552 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _327_
timestamp 1693170804
transform 1 0 11040 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _328_
timestamp 1693170804
transform 1 0 11316 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _329_
timestamp 1693170804
transform 1 0 11408 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _330_
timestamp 1693170804
transform 1 0 8464 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _331_
timestamp 1693170804
transform -1 0 8464 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _332_
timestamp 1693170804
transform 1 0 13064 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _333_
timestamp 1693170804
transform 1 0 13432 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _334_
timestamp 1693170804
transform 1 0 13064 0 -1 1632
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _335_
timestamp 1693170804
transform 1 0 9568 0 1 1632
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _336_
timestamp 1693170804
transform 1 0 8556 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _337_
timestamp 1693170804
transform 1 0 4232 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 10212 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _339_
timestamp 1693170804
transform 1 0 11960 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _340_
timestamp 1693170804
transform 1 0 11868 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _341_
timestamp 1693170804
transform 1 0 10948 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 7912 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1693170804
transform -1 0 4600 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1693170804
transform -1 0 4600 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1693170804
transform 1 0 8188 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1693170804
transform 1 0 8188 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  clone1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 6992 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clone7
timestamp 1693170804
transform 1 0 5060 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 1693170804
transform -1 0 1932 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1693170804
transform 1 0 4968 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 1693170804
transform 1 0 3312 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1693170804
transform 1 0 10028 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 1693170804
transform -1 0 9752 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 644 0 1 544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 1564 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 2760 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_36
timestamp 1693170804
transform 1 0 3404 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4508 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_63
timestamp 1693170804
transform 1 0 5888 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_71
timestamp 1693170804
transform 1 0 6624 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_80 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 7452 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1693170804
transform 1 0 7912 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8648 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_98
timestamp 1693170804
transform 1 0 9108 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 10212 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1693170804
transform 1 0 10488 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_122
timestamp 1693170804
transform 1 0 11316 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_134
timestamp 1693170804
transform 1 0 12420 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1693170804
transform 1 0 13064 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_153
timestamp 1693170804
transform 1 0 14168 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_160
timestamp 1693170804
transform 1 0 14812 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_164
timestamp 1693170804
transform 1 0 15180 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3
timestamp 1693170804
transform 1 0 368 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_11
timestamp 1693170804
transform 1 0 1104 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1693170804
transform 1 0 1472 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_27
timestamp 1693170804
transform 1 0 2576 0 -1 1632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_34
timestamp 1693170804
transform 1 0 3220 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_46
timestamp 1693170804
transform 1 0 4324 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1693170804
transform 1 0 5060 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1693170804
transform 1 0 5336 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1693170804
transform 1 0 6440 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_81
timestamp 1693170804
transform 1 0 7544 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_89
timestamp 1693170804
transform 1 0 8280 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_95
timestamp 1693170804
transform 1 0 8832 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_103
timestamp 1693170804
transform 1 0 9568 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_119
timestamp 1693170804
transform 1 0 11040 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_126
timestamp 1693170804
transform 1 0 11684 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_138
timestamp 1693170804
transform 1 0 12788 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_161
timestamp 1693170804
transform 1 0 14904 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1693170804
transform 1 0 368 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1693170804
transform 1 0 1472 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1693170804
transform 1 0 2576 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1693170804
transform 1 0 2760 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_41
timestamp 1693170804
transform 1 0 3864 0 1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_67
timestamp 1693170804
transform 1 0 6256 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_79
timestamp 1693170804
transform 1 0 7360 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1693170804
transform 1 0 7728 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1693170804
transform 1 0 7912 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_97
timestamp 1693170804
transform 1 0 9016 0 1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_123
timestamp 1693170804
transform 1 0 11408 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_135
timestamp 1693170804
transform 1 0 12512 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1693170804
transform 1 0 12880 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_141
timestamp 1693170804
transform 1 0 13064 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_148
timestamp 1693170804
transform 1 0 13708 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_158
timestamp 1693170804
transform 1 0 14628 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_165
timestamp 1693170804
transform 1 0 15272 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1693170804
transform 1 0 368 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_15
timestamp 1693170804
transform 1 0 1472 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_21
timestamp 1693170804
transform 1 0 2024 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_42
timestamp 1693170804
transform 1 0 3956 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1693170804
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1693170804
transform 1 0 5336 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_69
timestamp 1693170804
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1693170804
transform 1 0 10304 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_120
timestamp 1693170804
transform 1 0 11132 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_143
timestamp 1693170804
transform 1 0 13248 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_147
timestamp 1693170804
transform 1 0 13616 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_153
timestamp 1693170804
transform 1 0 14168 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 1693170804
transform 1 0 644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1693170804
transform 1 0 1748 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1693170804
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_29
timestamp 1693170804
transform 1 0 2760 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_39
timestamp 1693170804
transform 1 0 3680 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_57
timestamp 1693170804
transform 1 0 5336 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_69
timestamp 1693170804
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 1693170804
transform 1 0 7544 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_85
timestamp 1693170804
transform 1 0 7912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_117
timestamp 1693170804
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_126
timestamp 1693170804
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1693170804
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_141
timestamp 1693170804
transform 1 0 13064 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_155
timestamp 1693170804
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_12
timestamp 1693170804
transform 1 0 1196 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_18
timestamp 1693170804
transform 1 0 1748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_39
timestamp 1693170804
transform 1 0 3680 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_47
timestamp 1693170804
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_53
timestamp 1693170804
transform 1 0 4968 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1693170804
transform 1 0 5336 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_69
timestamp 1693170804
transform 1 0 6440 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_73
timestamp 1693170804
transform 1 0 6808 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_88
timestamp 1693170804
transform 1 0 8188 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 1693170804
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1693170804
transform 1 0 368 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_7
timestamp 1693170804
transform 1 0 736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_15
timestamp 1693170804
transform 1 0 1472 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1693170804
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1693170804
transform 1 0 2760 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_37
timestamp 1693170804
transform 1 0 3496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_61
timestamp 1693170804
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_68
timestamp 1693170804
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 1693170804
transform 1 0 7544 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_89
timestamp 1693170804
transform 1 0 8280 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_95
timestamp 1693170804
transform 1 0 8832 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_108
timestamp 1693170804
transform 1 0 10028 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_114
timestamp 1693170804
transform 1 0 10580 0 1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_125
timestamp 1693170804
transform 1 0 11592 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 1693170804
transform 1 0 12696 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_141
timestamp 1693170804
transform 1 0 13064 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_150
timestamp 1693170804
transform 1 0 13892 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_157
timestamp 1693170804
transform 1 0 14536 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_167
timestamp 1693170804
transform 1 0 15456 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_23
timestamp 1693170804
transform 1 0 2208 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_44
timestamp 1693170804
transform 1 0 4140 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_63
timestamp 1693170804
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_68
timestamp 1693170804
transform 1 0 6348 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_79
timestamp 1693170804
transform 1 0 7360 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_87
timestamp 1693170804
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_94
timestamp 1693170804
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1693170804
transform 1 0 10304 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_113
timestamp 1693170804
transform 1 0 10488 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_145
timestamp 1693170804
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_153
timestamp 1693170804
transform 1 0 14168 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_157
timestamp 1693170804
transform 1 0 14536 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_161
timestamp 1693170804
transform 1 0 14904 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1693170804
transform 1 0 368 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1693170804
transform 1 0 1472 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1693170804
transform 1 0 2576 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1693170804
transform 1 0 2760 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_33
timestamp 1693170804
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_57
timestamp 1693170804
transform 1 0 5336 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_77
timestamp 1693170804
transform 1 0 7176 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1693170804
transform 1 0 7912 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_100
timestamp 1693170804
transform 1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_112
timestamp 1693170804
transform 1 0 10396 0 1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1693170804
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_133
timestamp 1693170804
transform 1 0 12328 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_166
timestamp 1693170804
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 1693170804
transform 1 0 920 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_13
timestamp 1693170804
transform 1 0 1288 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_18
timestamp 1693170804
transform 1 0 1748 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_26
timestamp 1693170804
transform 1 0 2484 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_52
timestamp 1693170804
transform 1 0 4876 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 1693170804
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_64
timestamp 1693170804
transform 1 0 5980 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_76
timestamp 1693170804
transform 1 0 7084 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_86
timestamp 1693170804
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1693170804
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1693170804
transform 1 0 11592 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1693170804
transform 1 0 12696 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_149
timestamp 1693170804
transform 1 0 13800 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_157
timestamp 1693170804
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_29
timestamp 1693170804
transform 1 0 2760 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_35
timestamp 1693170804
transform 1 0 3312 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_44
timestamp 1693170804
transform 1 0 4140 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_68
timestamp 1693170804
transform 1 0 6348 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1693170804
transform 1 0 7452 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1693170804
transform 1 0 7912 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_93
timestamp 1693170804
transform 1 0 8648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_115
timestamp 1693170804
transform 1 0 10672 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1693170804
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_165
timestamp 1693170804
transform 1 0 15272 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_7
timestamp 1693170804
transform 1 0 736 0 -1 7072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1693170804
transform 1 0 1748 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_30
timestamp 1693170804
transform 1 0 2852 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_42
timestamp 1693170804
transform 1 0 3956 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_47
timestamp 1693170804
transform 1 0 4416 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1693170804
transform 1 0 5152 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1693170804
transform 1 0 5336 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_72
timestamp 1693170804
transform 1 0 6716 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_80
timestamp 1693170804
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_87
timestamp 1693170804
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1693170804
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_113
timestamp 1693170804
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_117
timestamp 1693170804
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_123
timestamp 1693170804
transform 1 0 11408 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_135
timestamp 1693170804
transform 1 0 12512 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_147
timestamp 1693170804
transform 1 0 13616 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_159
timestamp 1693170804
transform 1 0 14720 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_23
timestamp 1693170804
transform 1 0 2208 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1693170804
transform 1 0 2576 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_49
timestamp 1693170804
transform 1 0 4600 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_62
timestamp 1693170804
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_105
timestamp 1693170804
transform 1 0 9752 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_131
timestamp 1693170804
transform 1 0 12144 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1693170804
transform 1 0 12880 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_167
timestamp 1693170804
transform 1 0 15456 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_20
timestamp 1693170804
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_52
timestamp 1693170804
transform 1 0 4876 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_57
timestamp 1693170804
transform 1 0 5336 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_69
timestamp 1693170804
transform 1 0 6440 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_96
timestamp 1693170804
transform 1 0 8924 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_100
timestamp 1693170804
transform 1 0 9292 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1693170804
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_113
timestamp 1693170804
transform 1 0 10488 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_119
timestamp 1693170804
transform 1 0 11040 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_127
timestamp 1693170804
transform 1 0 11776 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_149
timestamp 1693170804
transform 1 0 13800 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_153
timestamp 1693170804
transform 1 0 14168 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_161
timestamp 1693170804
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_9
timestamp 1693170804
transform 1 0 920 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_14
timestamp 1693170804
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_20
timestamp 1693170804
transform 1 0 1932 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1693170804
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1693170804
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_76
timestamp 1693170804
transform 1 0 7084 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1693170804
transform 1 0 7912 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_92
timestamp 1693170804
transform 1 0 8556 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_100
timestamp 1693170804
transform 1 0 9292 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_107
timestamp 1693170804
transform 1 0 9936 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_119
timestamp 1693170804
transform 1 0 11040 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_131
timestamp 1693170804
transform 1 0 12144 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1693170804
transform 1 0 12880 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_148
timestamp 1693170804
transform 1 0 13708 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_152
timestamp 1693170804
transform 1 0 14076 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_158
timestamp 1693170804
transform 1 0 14628 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_164
timestamp 1693170804
transform 1 0 15180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_3
timestamp 1693170804
transform 1 0 368 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_31
timestamp 1693170804
transform 1 0 2944 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_39
timestamp 1693170804
transform 1 0 3680 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_45
timestamp 1693170804
transform 1 0 4232 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1693170804
transform 1 0 4968 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_63
timestamp 1693170804
transform 1 0 5888 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_71
timestamp 1693170804
transform 1 0 6624 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_75
timestamp 1693170804
transform 1 0 6992 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_87
timestamp 1693170804
transform 1 0 8096 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_96
timestamp 1693170804
transform 1 0 8924 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_100
timestamp 1693170804
transform 1 0 9292 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1693170804
transform 1 0 9752 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1693170804
transform 1 0 10304 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1693170804
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_118
timestamp 1693170804
transform 1 0 10948 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_128
timestamp 1693170804
transform 1 0 11868 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_159
timestamp 1693170804
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_7
timestamp 1693170804
transform 1 0 736 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_12
timestamp 1693170804
transform 1 0 1196 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_20
timestamp 1693170804
transform 1 0 1932 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_36
timestamp 1693170804
transform 1 0 3404 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_44
timestamp 1693170804
transform 1 0 4140 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_67
timestamp 1693170804
transform 1 0 6256 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_79
timestamp 1693170804
transform 1 0 7360 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1693170804
transform 1 0 7728 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_85
timestamp 1693170804
transform 1 0 7912 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_109
timestamp 1693170804
transform 1 0 10120 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_131
timestamp 1693170804
transform 1 0 12144 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1693170804
transform 1 0 12880 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1693170804
transform 1 0 13064 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_153
timestamp 1693170804
transform 1 0 14168 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_167
timestamp 1693170804
transform 1 0 15456 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_23
timestamp 1693170804
transform 1 0 2208 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1693170804
transform 1 0 5336 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_68
timestamp 1693170804
transform 1 0 6348 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_89
timestamp 1693170804
transform 1 0 8280 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_95
timestamp 1693170804
transform 1 0 8832 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_101
timestamp 1693170804
transform 1 0 9384 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1693170804
transform 1 0 10120 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1693170804
transform 1 0 10488 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1693170804
transform 1 0 11592 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1693170804
transform 1 0 12696 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1693170804
transform 1 0 13800 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_161
timestamp 1693170804
transform 1 0 14904 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_7
timestamp 1693170804
transform 1 0 736 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_13
timestamp 1693170804
transform 1 0 1288 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_20
timestamp 1693170804
transform 1 0 1932 0 1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1693170804
transform 1 0 2760 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1693170804
transform 1 0 3864 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1693170804
transform 1 0 4968 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_72
timestamp 1693170804
transform 1 0 6716 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_105
timestamp 1693170804
transform 1 0 9752 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1693170804
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_121
timestamp 1693170804
transform 1 0 11224 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_130
timestamp 1693170804
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_136
timestamp 1693170804
transform 1 0 12604 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1693170804
transform 1 0 13064 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_153
timestamp 1693170804
transform 1 0 14168 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_161
timestamp 1693170804
transform 1 0 14904 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_165
timestamp 1693170804
transform 1 0 15272 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_3
timestamp 1693170804
transform 1 0 368 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_25
timestamp 1693170804
transform 1 0 2392 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_57
timestamp 1693170804
transform 1 0 5336 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_70
timestamp 1693170804
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_92
timestamp 1693170804
transform 1 0 8556 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_104
timestamp 1693170804
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1693170804
transform 1 0 10488 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1693170804
transform 1 0 11592 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1693170804
transform 1 0 12696 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_149
timestamp 1693170804
transform 1 0 13800 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_157
timestamp 1693170804
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_7
timestamp 1693170804
transform 1 0 736 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_13
timestamp 1693170804
transform 1 0 1288 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_18
timestamp 1693170804
transform 1 0 1748 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 1693170804
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_29
timestamp 1693170804
transform 1 0 2760 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_39
timestamp 1693170804
transform 1 0 3680 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_43
timestamp 1693170804
transform 1 0 4048 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_47
timestamp 1693170804
transform 1 0 4416 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_54
timestamp 1693170804
transform 1 0 5060 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_62
timestamp 1693170804
transform 1 0 5796 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_67
timestamp 1693170804
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_71
timestamp 1693170804
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_75
timestamp 1693170804
transform 1 0 6992 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1693170804
transform 1 0 7728 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1693170804
transform 1 0 7912 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_91
timestamp 1693170804
transform 1 0 8464 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1693170804
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1693170804
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1693170804
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1693170804
transform 1 0 12328 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1693170804
transform 1 0 12880 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1693170804
transform 1 0 13064 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1693170804
transform 1 0 14168 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_165
timestamp 1693170804
transform 1 0 15272 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1693170804
transform 1 0 368 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_25
timestamp 1693170804
transform 1 0 2392 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_34
timestamp 1693170804
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_57
timestamp 1693170804
transform 1 0 5336 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_63
timestamp 1693170804
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_88
timestamp 1693170804
transform 1 0 8188 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_100
timestamp 1693170804
transform 1 0 9292 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1693170804
transform 1 0 10488 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1693170804
transform 1 0 11592 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1693170804
transform 1 0 12696 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_149
timestamp 1693170804
transform 1 0 13800 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_157
timestamp 1693170804
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_9
timestamp 1693170804
transform 1 0 920 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_20
timestamp 1693170804
transform 1 0 1932 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 1693170804
transform 1 0 2760 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_39
timestamp 1693170804
transform 1 0 3680 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_51
timestamp 1693170804
transform 1 0 4784 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_55
timestamp 1693170804
transform 1 0 5152 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_63
timestamp 1693170804
transform 1 0 5888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_69
timestamp 1693170804
transform 1 0 6440 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_73
timestamp 1693170804
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_80
timestamp 1693170804
transform 1 0 7452 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1693170804
transform 1 0 7912 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_93
timestamp 1693170804
transform 1 0 8648 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_98
timestamp 1693170804
transform 1 0 9108 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_110
timestamp 1693170804
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_113
timestamp 1693170804
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_119
timestamp 1693170804
transform 1 0 11040 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_131
timestamp 1693170804
transform 1 0 12144 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_135
timestamp 1693170804
transform 1 0 12512 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1693170804
transform 1 0 13064 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_153
timestamp 1693170804
transform 1 0 14168 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_160
timestamp 1693170804
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1693170804
transform 1 0 920 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1693170804
transform -1 0 15548 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1693170804
transform -1 0 644 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1693170804
transform 1 0 368 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1693170804
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1693170804
transform -1 0 1564 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1693170804
transform 1 0 3036 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1693170804
transform 1 0 14444 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1693170804
transform 1 0 12604 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1693170804
transform -1 0 11040 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1693170804
transform 1 0 8740 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 1693170804
transform 1 0 6900 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1693170804
transform 1 0 5336 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1693170804
transform -1 0 1564 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1693170804
transform -1 0 3404 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1693170804
transform 1 0 14444 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1693170804
transform 1 0 12604 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1693170804
transform -1 0 11040 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1693170804
transform -1 0 9108 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1693170804
transform 1 0 6900 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1693170804
transform 1 0 5336 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1693170804
transform -1 0 736 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1693170804
transform -1 0 736 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1693170804
transform -1 0 920 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1693170804
transform -1 0 736 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1693170804
transform -1 0 736 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1693170804
transform -1 0 736 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 1693170804
transform -1 0 920 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1693170804
transform -1 0 1932 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1693170804
transform -1 0 920 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1693170804
transform 1 0 14996 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1693170804
transform -1 0 15548 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1693170804
transform 1 0 14996 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1693170804
transform 1 0 14996 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1693170804
transform 1 0 14996 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1693170804
transform 1 0 14996 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1693170804
transform 1 0 14996 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 1693170804
transform 1 0 14996 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1693170804
transform 1 0 14996 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1693170804
transform 1 0 14996 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1693170804
transform -1 0 920 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_23
timestamp 1693170804
transform 1 0 92 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1693170804
transform -1 0 15824 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_24
timestamp 1693170804
transform 1 0 92 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1693170804
transform -1 0 15824 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_25
timestamp 1693170804
transform 1 0 92 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1693170804
transform -1 0 15824 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_26
timestamp 1693170804
transform 1 0 92 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1693170804
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_27
timestamp 1693170804
transform 1 0 92 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1693170804
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_28
timestamp 1693170804
transform 1 0 92 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1693170804
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_29
timestamp 1693170804
transform 1 0 92 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1693170804
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_30
timestamp 1693170804
transform 1 0 92 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1693170804
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_31
timestamp 1693170804
transform 1 0 92 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1693170804
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_32
timestamp 1693170804
transform 1 0 92 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1693170804
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_33
timestamp 1693170804
transform 1 0 92 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1693170804
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_34
timestamp 1693170804
transform 1 0 92 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1693170804
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_35
timestamp 1693170804
transform 1 0 92 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1693170804
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_36
timestamp 1693170804
transform 1 0 92 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1693170804
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_37
timestamp 1693170804
transform 1 0 92 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1693170804
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_38
timestamp 1693170804
transform 1 0 92 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1693170804
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_39
timestamp 1693170804
transform 1 0 92 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1693170804
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_40
timestamp 1693170804
transform 1 0 92 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1693170804
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_41
timestamp 1693170804
transform 1 0 92 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1693170804
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_42
timestamp 1693170804
transform 1 0 92 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1693170804
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_43
timestamp 1693170804
transform 1 0 92 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1693170804
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_44
timestamp 1693170804
transform 1 0 92 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1693170804
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_45
timestamp 1693170804
transform 1 0 92 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1693170804
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer1
timestamp 1693170804
transform 1 0 14260 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer2
timestamp 1693170804
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer3
timestamp 1693170804
transform 1 0 10948 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  rebuffer4
timestamp 1693170804
transform -1 0 7084 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  rebuffer5
timestamp 1693170804
transform -1 0 6440 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  rebuffer6
timestamp 1693170804
transform -1 0 6992 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 2668 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_47
timestamp 1693170804
transform 1 0 5244 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_48
timestamp 1693170804
transform 1 0 7820 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_49
timestamp 1693170804
transform 1 0 10396 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_50
timestamp 1693170804
transform 1 0 12972 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_51
timestamp 1693170804
transform 1 0 5244 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_52
timestamp 1693170804
transform 1 0 10396 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp 1693170804
transform 1 0 2668 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_54
timestamp 1693170804
transform 1 0 7820 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_55
timestamp 1693170804
transform 1 0 12972 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp 1693170804
transform 1 0 5244 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp 1693170804
transform 1 0 10396 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_58
timestamp 1693170804
transform 1 0 2668 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp 1693170804
transform 1 0 7820 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp 1693170804
transform 1 0 12972 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_61
timestamp 1693170804
transform 1 0 5244 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_62
timestamp 1693170804
transform 1 0 10396 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_63
timestamp 1693170804
transform 1 0 2668 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_64
timestamp 1693170804
transform 1 0 7820 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_65
timestamp 1693170804
transform 1 0 12972 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_66
timestamp 1693170804
transform 1 0 5244 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_67
timestamp 1693170804
transform 1 0 10396 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_68
timestamp 1693170804
transform 1 0 2668 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_69
timestamp 1693170804
transform 1 0 7820 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_70
timestamp 1693170804
transform 1 0 12972 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_71
timestamp 1693170804
transform 1 0 5244 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_72
timestamp 1693170804
transform 1 0 10396 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_73
timestamp 1693170804
transform 1 0 2668 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_74
timestamp 1693170804
transform 1 0 7820 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_75
timestamp 1693170804
transform 1 0 12972 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_76
timestamp 1693170804
transform 1 0 5244 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_77
timestamp 1693170804
transform 1 0 10396 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_78
timestamp 1693170804
transform 1 0 2668 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_79
timestamp 1693170804
transform 1 0 7820 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_80
timestamp 1693170804
transform 1 0 12972 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_81
timestamp 1693170804
transform 1 0 5244 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_82
timestamp 1693170804
transform 1 0 10396 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_83
timestamp 1693170804
transform 1 0 2668 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_84
timestamp 1693170804
transform 1 0 7820 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_85
timestamp 1693170804
transform 1 0 12972 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_86
timestamp 1693170804
transform 1 0 5244 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_87
timestamp 1693170804
transform 1 0 10396 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_88
timestamp 1693170804
transform 1 0 2668 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_89
timestamp 1693170804
transform 1 0 7820 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_90
timestamp 1693170804
transform 1 0 12972 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_91
timestamp 1693170804
transform 1 0 5244 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_92
timestamp 1693170804
transform 1 0 10396 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_93
timestamp 1693170804
transform 1 0 2668 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_94
timestamp 1693170804
transform 1 0 7820 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_95
timestamp 1693170804
transform 1 0 12972 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_96
timestamp 1693170804
transform 1 0 5244 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_97
timestamp 1693170804
transform 1 0 10396 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_98
timestamp 1693170804
transform 1 0 2668 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_99
timestamp 1693170804
transform 1 0 7820 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_100
timestamp 1693170804
transform 1 0 12972 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_101
timestamp 1693170804
transform 1 0 5244 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_102
timestamp 1693170804
transform 1 0 10396 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_103
timestamp 1693170804
transform 1 0 2668 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_104
timestamp 1693170804
transform 1 0 5244 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_105
timestamp 1693170804
transform 1 0 7820 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_106
timestamp 1693170804
transform 1 0 10396 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_107
timestamp 1693170804
transform 1 0 12972 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire42
timestamp 1693170804
transform -1 0 7820 0 1 4896
box -38 -48 314 592
<< labels >>
flabel metal4 s 2558 496 2878 13104 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6491 496 6811 13104 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10424 496 10744 13104 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14357 496 14677 13104 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 44 2608 15872 2928 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 44 5736 15872 6056 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 44 8864 15872 9184 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 44 11992 15872 12312 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1898 496 2218 13104 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5831 496 6151 13104 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9764 496 10084 13104 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13697 496 14017 13104 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 44 1948 15872 2268 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 44 5076 15872 5396 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 44 8204 15872 8524 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 44 11332 15872 11652 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 3574 200 3634 0 FreeSans 480 0 0 0 cal
port 2 nsew signal input
flabel metal3 s 0 1670 200 1730 0 FreeSans 480 0 0 0 clk
port 3 nsew signal input
flabel metal3 s 15800 6430 16000 6490 0 FreeSans 480 0 0 0 clkc
port 4 nsew signal tristate
flabel metal3 s 15800 7518 16000 7578 0 FreeSans 480 0 0 0 comp
port 5 nsew signal input
flabel metal3 s 1096 0 1216 200 0 FreeSans 960 0 0 0 ctln[0]
port 6 nsew signal tristate
flabel metal3 s 3000 0 3120 200 0 FreeSans 960 0 0 0 ctln[1]
port 7 nsew signal tristate
flabel metal3 s 14424 0 14544 200 0 FreeSans 960 0 0 0 ctln[2]
port 8 nsew signal tristate
flabel metal3 s 12520 0 12640 200 0 FreeSans 960 0 0 0 ctln[3]
port 9 nsew signal tristate
flabel metal3 s 10616 0 10736 200 0 FreeSans 960 0 0 0 ctln[4]
port 10 nsew signal tristate
flabel metal3 s 8712 0 8832 200 0 FreeSans 960 0 0 0 ctln[5]
port 11 nsew signal tristate
flabel metal3 s 6808 0 6928 200 0 FreeSans 960 0 0 0 ctln[6]
port 12 nsew signal tristate
flabel metal3 s 4904 0 5024 200 0 FreeSans 960 0 0 0 ctln[7]
port 13 nsew signal tristate
flabel metal3 s 1096 13800 1216 14000 0 FreeSans 960 0 0 0 ctlp[0]
port 14 nsew signal tristate
flabel metal3 s 3000 13800 3120 14000 0 FreeSans 960 0 0 0 ctlp[1]
port 15 nsew signal tristate
flabel metal3 s 14424 13800 14544 14000 0 FreeSans 960 0 0 0 ctlp[2]
port 16 nsew signal tristate
flabel metal3 s 12520 13800 12640 14000 0 FreeSans 960 0 0 0 ctlp[3]
port 17 nsew signal tristate
flabel metal3 s 10616 13800 10736 14000 0 FreeSans 960 0 0 0 ctlp[4]
port 18 nsew signal tristate
flabel metal3 s 8712 13800 8832 14000 0 FreeSans 960 0 0 0 ctlp[5]
port 19 nsew signal tristate
flabel metal3 s 6808 13800 6928 14000 0 FreeSans 960 0 0 0 ctlp[6]
port 20 nsew signal tristate
flabel metal3 s 4904 13800 5024 14000 0 FreeSans 960 0 0 0 ctlp[7]
port 21 nsew signal tristate
flabel metal3 s 0 2622 200 2682 0 FreeSans 480 0 0 0 en
port 22 nsew signal input
flabel metal3 s 0 6430 200 6490 0 FreeSans 480 0 0 0 result[0]
port 23 nsew signal tristate
flabel metal3 s 0 7382 200 7442 0 FreeSans 480 0 0 0 result[1]
port 24 nsew signal tristate
flabel metal3 s 0 8334 200 8394 0 FreeSans 480 0 0 0 result[2]
port 25 nsew signal tristate
flabel metal3 s 0 9286 200 9346 0 FreeSans 480 0 0 0 result[3]
port 26 nsew signal tristate
flabel metal3 s 0 10238 200 10298 0 FreeSans 480 0 0 0 result[4]
port 27 nsew signal tristate
flabel metal3 s 0 11190 200 11250 0 FreeSans 480 0 0 0 result[5]
port 28 nsew signal tristate
flabel metal3 s 0 12142 200 12202 0 FreeSans 480 0 0 0 result[6]
port 29 nsew signal tristate
flabel metal3 s 0 13094 200 13154 0 FreeSans 480 0 0 0 result[7]
port 30 nsew signal tristate
flabel metal3 s 0 718 200 778 0 FreeSans 480 0 0 0 rstn
port 31 nsew signal input
flabel metal3 s 0 5478 200 5538 0 FreeSans 480 0 0 0 sample
port 32 nsew signal tristate
flabel metal3 s 15800 3166 16000 3226 0 FreeSans 480 0 0 0 trim[0]
port 33 nsew signal tristate
flabel metal3 s 15800 4254 16000 4314 0 FreeSans 480 0 0 0 trim[1]
port 34 nsew signal tristate
flabel metal3 s 15800 2078 16000 2138 0 FreeSans 480 0 0 0 trim[2]
port 35 nsew signal tristate
flabel metal3 s 15800 990 16000 1050 0 FreeSans 480 0 0 0 trim[3]
port 36 nsew signal tristate
flabel metal3 s 15800 5342 16000 5402 0 FreeSans 480 0 0 0 trim[4]
port 37 nsew signal tristate
flabel metal3 s 15800 10782 16000 10842 0 FreeSans 480 0 0 0 trimb[0]
port 38 nsew signal tristate
flabel metal3 s 15800 9694 16000 9754 0 FreeSans 480 0 0 0 trimb[1]
port 39 nsew signal tristate
flabel metal3 s 15800 11870 16000 11930 0 FreeSans 480 0 0 0 trimb[2]
port 40 nsew signal tristate
flabel metal3 s 15800 12958 16000 13018 0 FreeSans 480 0 0 0 trimb[3]
port 41 nsew signal tristate
flabel metal3 s 15800 8606 16000 8666 0 FreeSans 480 0 0 0 trimb[4]
port 42 nsew signal tristate
flabel metal3 s 0 4526 200 4586 0 FreeSans 480 0 0 0 valid
port 43 nsew signal tristate
rlabel metal1 7958 12512 7958 12512 0 VGND
rlabel metal1 7958 13056 7958 13056 0 VPWR
rlabel metal1 8648 9146 8648 9146 0 _000_
rlabel metal1 11684 7242 11684 7242 0 _001_
rlabel metal1 7130 8024 7130 8024 0 _002_
rlabel metal1 6394 6970 6394 6970 0 _003_
rlabel metal1 920 5882 920 5882 0 _004_
rlabel metal1 736 7378 736 7378 0 _005_
rlabel metal1 1196 8602 1196 8602 0 _006_
rlabel metal1 920 9690 920 9690 0 _007_
rlabel metal1 6440 10030 6440 10030 0 _008_
rlabel metal1 6440 12342 6440 12342 0 _009_
rlabel metal2 3542 12517 3542 12517 0 _010_
rlabel metal1 1058 11866 1058 11866 0 _011_
rlabel metal1 1058 4250 1058 4250 0 _012_
rlabel metal1 2208 3638 2208 3638 0 _013_
rlabel metal2 2438 3536 2438 3536 0 _014_
rlabel metal2 4738 2349 4738 2349 0 _015_
rlabel metal2 2714 7616 2714 7616 0 _016_
rlabel metal1 3726 8466 3726 8466 0 _017_
rlabel metal2 2806 9758 2806 9758 0 _018_
rlabel metal2 4738 9724 4738 9724 0 _019_
rlabel metal1 7452 10506 7452 10506 0 _020_
rlabel metal1 6762 11254 6762 11254 0 _021_
rlabel metal1 3634 11118 3634 11118 0 _022_
rlabel metal1 1150 10778 1150 10778 0 _023_
rlabel metal1 11500 4250 11500 4250 0 _024_
rlabel metal1 11454 3638 11454 3638 0 _025_
rlabel metal2 11684 2550 11684 2550 0 _026_
rlabel metal1 9660 2414 9660 2414 0 _027_
rlabel metal1 7866 2414 7866 2414 0 _028_
rlabel metal1 13156 5066 13156 5066 0 _029_
rlabel metal1 13662 3502 13662 3502 0 _030_
rlabel metal2 13386 1870 13386 1870 0 _031_
rlabel metal1 10028 1530 10028 1530 0 _032_
rlabel metal1 9752 3094 9752 3094 0 _033_
rlabel metal1 4452 6426 4452 6426 0 _034_
rlabel metal1 10764 9146 10764 9146 0 _035_
rlabel metal2 12374 8772 12374 8772 0 _036_
rlabel metal2 12282 7684 12282 7684 0 _037_
rlabel metal1 11362 5610 11362 5610 0 _038_
rlabel metal1 1978 6426 1978 6426 0 _039_
rlabel metal1 3082 8296 3082 8296 0 _040_
rlabel metal1 13938 9078 13938 9078 0 _041_
rlabel metal1 2714 9656 2714 9656 0 _042_
rlabel metal1 9614 10234 9614 10234 0 _043_
rlabel metal1 8602 11662 8602 11662 0 _044_
rlabel metal1 6026 12750 6026 12750 0 _045_
rlabel metal1 4186 11696 4186 11696 0 _046_
rlabel metal1 15180 4046 15180 4046 0 _047_
rlabel metal2 3726 4352 3726 4352 0 _048_
rlabel metal1 6256 6222 6256 6222 0 _049_
rlabel metal1 7176 5134 7176 5134 0 _050_
rlabel metal2 7774 3128 7774 3128 0 _051_
rlabel metal1 6900 4114 6900 4114 0 _052_
rlabel metal2 7314 3604 7314 3604 0 _053_
rlabel metal1 7774 3978 7774 3978 0 _054_
rlabel metal1 15134 3162 15134 3162 0 _055_
rlabel metal1 14996 1870 14996 1870 0 _056_
rlabel metal1 14950 816 14950 816 0 _057_
rlabel metal2 10534 4369 10534 4369 0 _058_
rlabel metal2 5474 5100 5474 5100 0 _059_
rlabel metal1 5520 4046 5520 4046 0 _060_
rlabel metal1 14950 6222 14950 6222 0 _061_
rlabel metal1 10120 5134 10120 5134 0 _062_
rlabel metal1 10810 7888 10810 7888 0 _063_
rlabel metal2 10902 2655 10902 2655 0 _064_
rlabel metal1 10994 6800 10994 6800 0 _065_
rlabel metal1 11132 5746 11132 5746 0 _066_
rlabel metal1 10120 6970 10120 6970 0 _067_
rlabel metal1 9154 6630 9154 6630 0 _068_
rlabel metal2 9890 8092 9890 8092 0 _069_
rlabel metal1 9614 8432 9614 8432 0 _070_
rlabel metal1 8740 6426 8740 6426 0 _071_
rlabel metal1 8326 7718 8326 7718 0 _072_
rlabel metal1 7176 6834 7176 6834 0 _073_
rlabel metal1 3634 12682 3634 12682 0 _074_
rlabel metal1 6026 5882 6026 5882 0 _075_
rlabel metal1 6394 8466 6394 8466 0 _076_
rlabel metal1 5980 8398 5980 8398 0 _077_
rlabel metal1 1334 7888 1334 7888 0 _078_
rlabel metal1 1242 5814 1242 5814 0 _079_
rlabel metal1 782 7888 782 7888 0 _080_
rlabel metal1 1978 8398 1978 8398 0 _081_
rlabel metal1 1380 9486 1380 9486 0 _082_
rlabel metal2 5934 10166 5934 10166 0 _083_
rlabel metal1 6302 12240 6302 12240 0 _084_
rlabel metal1 3450 12716 3450 12716 0 _085_
rlabel metal1 1242 11730 1242 11730 0 _086_
rlabel metal1 6072 4658 6072 4658 0 _087_
rlabel metal1 7176 4250 7176 4250 0 _088_
rlabel metal1 6118 4080 6118 4080 0 _089_
rlabel metal1 5060 4488 5060 4488 0 _090_
rlabel metal1 9890 6222 9890 6222 0 _091_
rlabel metal1 10764 5746 10764 5746 0 _092_
rlabel metal1 1242 4080 1242 4080 0 _093_
rlabel metal2 5198 5712 5198 5712 0 _094_
rlabel metal1 3450 5100 3450 5100 0 _095_
rlabel metal2 4830 4794 4830 4794 0 _096_
rlabel metal2 3358 4250 3358 4250 0 _097_
rlabel metal1 7038 5032 7038 5032 0 _098_
rlabel metal1 3082 4726 3082 4726 0 _099_
rlabel metal1 5014 4080 5014 4080 0 _100_
rlabel metal1 2346 7888 2346 7888 0 _101_
rlabel metal1 2254 10574 2254 10574 0 _102_
rlabel metal1 7866 4658 7866 4658 0 _103_
rlabel metal1 10534 2482 10534 2482 0 _104_
rlabel metal1 8602 5100 8602 5100 0 _105_
rlabel metal1 9016 4726 9016 4726 0 _106_
rlabel via2 5842 4675 5842 4675 0 _107_
rlabel metal1 9430 4012 9430 4012 0 _108_
rlabel metal1 13524 4590 13524 4590 0 _109_
rlabel metal1 12880 1938 12880 1938 0 _110_
rlabel metal1 12880 4794 12880 4794 0 _111_
rlabel metal1 13708 3162 13708 3162 0 _112_
rlabel metal1 13294 3570 13294 3570 0 _113_
rlabel metal1 13662 1870 13662 1870 0 _114_
rlabel metal1 13616 2074 13616 2074 0 _115_
rlabel metal1 9890 1360 9890 1360 0 _116_
rlabel metal1 10212 1394 10212 1394 0 _117_
rlabel metal1 9614 4080 9614 4080 0 _118_
rlabel metal1 9890 2958 9890 2958 0 _119_
rlabel metal1 3772 5338 3772 5338 0 _120_
rlabel metal1 4140 6426 4140 6426 0 _121_
rlabel metal2 13570 7106 13570 7106 0 _122_
rlabel metal2 13386 7854 13386 7854 0 _123_
rlabel metal1 10994 9010 10994 9010 0 _124_
rlabel metal1 14398 9078 14398 9078 0 _125_
rlabel metal1 14858 9010 14858 9010 0 _126_
rlabel metal1 14858 9554 14858 9554 0 _127_
rlabel metal1 13294 8432 13294 8432 0 _128_
rlabel metal1 14444 7922 14444 7922 0 _129_
rlabel metal1 14674 7378 14674 7378 0 _130_
rlabel metal1 14306 7174 14306 7174 0 _131_
rlabel metal1 15042 7514 15042 7514 0 _132_
rlabel metal1 13294 7378 13294 7378 0 _133_
rlabel metal2 14122 6528 14122 6528 0 _134_
rlabel metal1 13846 6290 13846 6290 0 _135_
rlabel metal2 10902 5831 10902 5831 0 _136_
rlabel metal3 636 3604 636 3604 0 cal
rlabel metal1 14582 8976 14582 8976 0 cal_count\[0\]
rlabel metal1 13662 8466 13662 8466 0 cal_count\[1\]
rlabel metal1 13754 7276 13754 7276 0 cal_count\[2\]
rlabel metal1 9246 5236 9246 5236 0 cal_count\[3\]
rlabel metal1 10120 8058 10120 8058 0 cal_itt\[0\]
rlabel metal1 9108 6834 9108 6834 0 cal_itt\[1\]
rlabel metal1 8556 8058 8556 8058 0 cal_itt\[2\]
rlabel metal1 7912 6766 7912 6766 0 cal_itt\[3\]
rlabel metal1 1656 4454 1656 4454 0 calibrate
rlabel metal3 1211 1700 1211 1700 0 clk
rlabel metal3 15694 6460 15694 6460 0 clkc
rlabel metal1 4508 5746 4508 5746 0 clknet_0_clk
rlabel metal1 2208 2414 2208 2414 0 clknet_2_0__leaf_clk
rlabel metal1 3772 9554 3772 9554 0 clknet_2_1__leaf_clk
rlabel metal1 13294 3502 13294 3502 0 clknet_2_2__leaf_clk
rlabel metal1 12650 6120 12650 6120 0 clknet_2_3__leaf_clk
rlabel metal3 15648 7548 15648 7548 0 comp
rlabel metal3 1260 68 1260 68 0 ctln[0]
rlabel metal3 3166 68 3166 68 0 ctln[1]
rlabel metal3 14640 68 14640 68 0 ctln[2]
rlabel metal3 12734 68 12734 68 0 ctln[3]
rlabel metal3 10733 68 10733 68 0 ctln[4]
rlabel metal3 8886 68 8886 68 0 ctln[5]
rlabel metal3 7014 68 7014 68 0 ctln[6]
rlabel metal3 5144 68 5144 68 0 ctln[7]
rlabel metal3 1069 13804 1069 13804 0 ctlp[0]
rlabel metal1 3220 12954 3220 12954 0 ctlp[1]
rlabel metal2 14674 13379 14674 13379 0 ctlp[2]
rlabel metal2 12834 13447 12834 13447 0 ctlp[3]
rlabel metal1 10856 12954 10856 12954 0 ctlp[4]
rlabel metal1 8924 12954 8924 12954 0 ctlp[5]
rlabel metal2 6670 13379 6670 13379 0 ctlp[6]
rlabel metal3 5144 13804 5144 13804 0 ctlp[7]
rlabel metal3 268 2652 268 2652 0 en
rlabel metal1 7452 6358 7452 6358 0 en_co_clk
rlabel metal1 2484 6222 2484 6222 0 mask\[0\]
rlabel metal1 1840 7990 1840 7990 0 mask\[1\]
rlabel metal1 4278 9078 4278 9078 0 mask\[2\]
rlabel metal2 2530 9758 2530 9758 0 mask\[3\]
rlabel metal1 9154 10200 9154 10200 0 mask\[4\]
rlabel metal2 8510 11458 8510 11458 0 mask\[5\]
rlabel metal1 3542 11628 3542 11628 0 mask\[6\]
rlabel metal2 2438 11798 2438 11798 0 mask\[7\]
rlabel metal1 920 4046 920 4046 0 net1
rlabel metal1 10994 748 10994 748 0 net10
rlabel metal1 8740 782 8740 782 0 net11
rlabel metal1 6716 782 6716 782 0 net12
rlabel metal1 5244 782 5244 782 0 net13
rlabel metal1 1472 6630 1472 6630 0 net14
rlabel metal1 3312 12750 3312 12750 0 net15
rlabel metal1 14306 12750 14306 12750 0 net16
rlabel metal1 12512 12750 12512 12750 0 net17
rlabel metal1 10580 10438 10580 10438 0 net18
rlabel metal1 8924 1394 8924 1394 0 net19
rlabel metal1 15134 8364 15134 8364 0 net2
rlabel metal1 6647 12614 6647 12614 0 net20
rlabel metal1 5152 11662 5152 11662 0 net21
rlabel metal1 1380 5814 1380 5814 0 net22
rlabel metal1 2300 8330 2300 8330 0 net23
rlabel metal1 1656 8806 1656 8806 0 net24
rlabel metal1 1150 9418 1150 9418 0 net25
rlabel metal1 690 10540 690 10540 0 net26
rlabel metal1 1334 11662 1334 11662 0 net27
rlabel metal1 1058 12682 1058 12682 0 net28
rlabel metal1 2116 12750 2116 12750 0 net29
rlabel metal1 1679 3162 1679 3162 0 net3
rlabel metal1 782 5712 782 5712 0 net30
rlabel metal1 14950 3944 14950 3944 0 net31
rlabel metal1 15456 3706 15456 3706 0 net32
rlabel metal1 15042 2550 15042 2550 0 net33
rlabel metal2 15134 1224 15134 1224 0 net34
rlabel metal1 14904 5746 14904 5746 0 net35
rlabel metal2 15134 10982 15134 10982 0 net36
rlabel metal1 15226 3910 15226 3910 0 net37
rlabel metal1 14996 11322 14996 11322 0 net38
rlabel metal1 14996 12410 14996 12410 0 net39
rlabel metal2 9522 4318 9522 4318 0 net4
rlabel metal2 14858 6919 14858 6919 0 net40
rlabel metal1 1288 3638 1288 3638 0 net41
rlabel metal1 8050 5270 8050 5270 0 net42
rlabel metal2 1518 11798 1518 11798 0 net43
rlabel metal2 7774 11764 7774 11764 0 net44
rlabel metal1 2077 4658 2077 4658 0 net45
rlabel metal1 13163 2482 13163 2482 0 net46
rlabel metal2 13110 8534 13110 8534 0 net47
rlabel metal1 14306 1972 14306 1972 0 net48
rlabel metal1 14352 2958 14352 2958 0 net49
rlabel metal1 15272 6426 15272 6426 0 net5
rlabel metal2 10994 3196 10994 3196 0 net50
rlabel metal1 6302 7888 6302 7888 0 net51
rlabel metal1 2714 11152 2714 11152 0 net52
rlabel metal1 6670 10574 6670 10574 0 net53
rlabel metal2 5290 3774 5290 3774 0 net54
rlabel metal1 5244 5134 5244 5134 0 net55
rlabel metal1 1426 782 1426 782 0 net6
rlabel metal2 3082 986 3082 986 0 net7
rlabel metal1 14398 782 14398 782 0 net8
rlabel metal2 12558 6596 12558 6596 0 net9
rlabel metal3 314 6460 314 6460 0 result[0]
rlabel metal3 314 7412 314 7412 0 result[1]
rlabel metal3 268 8364 268 8364 0 result[2]
rlabel metal3 314 9316 314 9316 0 result[3]
rlabel metal3 314 10268 314 10268 0 result[4]
rlabel metal3 314 11220 314 11220 0 result[5]
rlabel metal3 268 12172 268 12172 0 result[6]
rlabel metal1 1288 12886 1288 12886 0 result[7]
rlabel metal3 268 748 268 748 0 rstn
rlabel metal3 314 5508 314 5508 0 sample
rlabel metal1 4646 3570 4646 3570 0 state\[0\]
rlabel metal1 4922 2958 4922 2958 0 state\[1\]
rlabel metal1 6670 2958 6670 2958 0 state\[2\]
rlabel metal1 15456 3162 15456 3162 0 trim[0]
rlabel metal3 15602 4284 15602 4284 0 trim[1]
rlabel metal3 15648 2108 15648 2108 0 trim[2]
rlabel metal3 15648 1020 15648 1020 0 trim[3]
rlabel metal3 15648 5372 15648 5372 0 trim[4]
rlabel metal2 8878 5236 8878 5236 0 trim_mask\[0\]
rlabel metal1 13846 2822 13846 2822 0 trim_mask\[1\]
rlabel metal1 13892 2550 13892 2550 0 trim_mask\[2\]
rlabel metal1 10902 2482 10902 2482 0 trim_mask\[3\]
rlabel metal1 11178 2482 11178 2482 0 trim_mask\[4\]
rlabel metal1 14812 4998 14812 4998 0 trim_val\[0\]
rlabel metal1 14812 2958 14812 2958 0 trim_val\[1\]
rlabel metal1 14812 2482 14812 2482 0 trim_val\[2\]
rlabel metal1 11408 1462 11408 1462 0 trim_val\[3\]
rlabel metal1 10028 4046 10028 4046 0 trim_val\[4\]
rlabel metal3 15717 10812 15717 10812 0 trimb[0]
rlabel metal3 15648 9724 15648 9724 0 trimb[1]
rlabel metal3 15648 11900 15648 11900 0 trimb[2]
rlabel metal1 15456 12954 15456 12954 0 trimb[3]
rlabel metal3 15648 8636 15648 8636 0 trimb[4]
rlabel metal3 199 4556 199 4556 0 valid
<< properties >>
string FIXED_BBOX 0 0 16000 14000
<< end >>
