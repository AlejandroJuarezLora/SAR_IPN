* NGSPICE file created from comparator.ext - technology: sky130B

.subckt sky130_fd_pr__cap_mim_m3_1_FJFAMD m3_n386_n240# c1_n346_n200#
X0 c1_n346_n200# m3_n386_n240# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt trimcap m1_179_405# m1_176_1185#
XXC2 m1_179_405# m1_176_1185# sky130_fd_pr__cap_mim_m3_1_FJFAMD
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_E33R59 D S G B
X0 S G D B sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt trim DRAIN VSS d0 d1 d2 d3 d4
Xtrimcap_12 DRAIN sky130_fd_pr__nfet_01v8_lvt_E33R59_2/D trimcap
Xtrimcap_11 DRAIN sky130_fd_pr__nfet_01v8_lvt_E33R59_2/D trimcap
Xtrimcap_13 DRAIN sky130_fd_pr__nfet_01v8_lvt_E33R59_2/D trimcap
Xtrimcap_14 DRAIN sky130_fd_pr__nfet_01v8_lvt_E33R59_2/D trimcap
Xtrimcap_15 DRAIN sky130_fd_pr__nfet_01v8_lvt_E33R59_2/D trimcap
Xtrimcap_0 DRAIN sky130_fd_pr__nfet_01v8_lvt_E33R59_2/D trimcap
Xtrimcap_1 sky130_fd_pr__nfet_01v8_lvt_E33R59_1/D DRAIN trimcap
Xtrimcap_2 sky130_fd_pr__nfet_01v8_lvt_E33R59_3/D DRAIN trimcap
Xsky130_fd_pr__nfet_01v8_lvt_E33R59_0 sky130_fd_pr__nfet_01v8_lvt_E33R59_0/D VSS d2
+ VSS sky130_fd_pr__nfet_01v8_lvt_E33R59
Xsky130_fd_pr__nfet_01v8_lvt_E33R59_1 sky130_fd_pr__nfet_01v8_lvt_E33R59_1/D VSS d0
+ VSS sky130_fd_pr__nfet_01v8_lvt_E33R59
Xtrimcap_3 sky130_fd_pr__nfet_01v8_lvt_E33R59_0/D DRAIN trimcap
Xtrimcap_4 sky130_fd_pr__nfet_01v8_lvt_E33R59_0/D DRAIN trimcap
Xsky130_fd_pr__nfet_01v8_lvt_E33R59_2 sky130_fd_pr__nfet_01v8_lvt_E33R59_2/D VSS d4
+ VSS sky130_fd_pr__nfet_01v8_lvt_E33R59
Xsky130_fd_pr__nfet_01v8_lvt_E33R59_3 sky130_fd_pr__nfet_01v8_lvt_E33R59_3/D VSS d1
+ VSS sky130_fd_pr__nfet_01v8_lvt_E33R59
Xtrimcap_5 sky130_fd_pr__nfet_01v8_lvt_E33R59_4/D DRAIN trimcap
Xtrimcap_6 sky130_fd_pr__nfet_01v8_lvt_E33R59_4/D DRAIN trimcap
Xsky130_fd_pr__nfet_01v8_lvt_E33R59_4 sky130_fd_pr__nfet_01v8_lvt_E33R59_4/D VSS d3
+ VSS sky130_fd_pr__nfet_01v8_lvt_E33R59
Xtrimcap_7 sky130_fd_pr__nfet_01v8_lvt_E33R59_4/D DRAIN trimcap
Xtrimcap_8 sky130_fd_pr__nfet_01v8_lvt_E33R59_4/D DRAIN trimcap
Xtrimcap_9 DRAIN sky130_fd_pr__nfet_01v8_lvt_E33R59_2/D trimcap
Xtrimcap_10 DRAIN sky130_fd_pr__nfet_01v8_lvt_E33R59_2/D trimcap
.ends

.subckt sky130_fd_pr__nfet_01v8_96AECY D S G B
X0 S G D B sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt sky130_fd_pr__pfet_01v8_7G6J3C D S G B
X0 S G D B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
.ends

.subckt comparator vdd vss vn vp outn outp clk trim0 trim1 trim2 trim3 trim4 trimb0
+ trimb1 trimb2 trimb3 trimb4
Xtrim_0 IP vss trimb0 trimb1 trimb2 trimb3 trimb4 trim
Xtrim_1 IN vss trim0 trim1 trim2 trim3 trim4 trim
Xsky130_fd_pr__nfet_01v8_96AECY_0 IN diff vn vss sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__nfet_01v8_96AECY_1 IP diff vp vss sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__nfet_01v8_96AECY_2 outn IN outp vss sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__nfet_01v8_96AECY_3 outp IP outn vss sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__nfet_01v8_96AECY_5 diff vss clk vss sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__nfet_01v8_96AECY_4 diff vss clk vss sky130_fd_pr__nfet_01v8_96AECY
Xsky130_fd_pr__pfet_01v8_7G6J3C_0 outp vdd outn sky130_fd_pr__pfet_01v8_7G6J3C_0/B
+ sky130_fd_pr__pfet_01v8_7G6J3C
Xsky130_fd_pr__pfet_01v8_7G6J3C_1 outn vdd outp sky130_fd_pr__pfet_01v8_7G6J3C_1/B
+ sky130_fd_pr__pfet_01v8_7G6J3C
Xsky130_fd_pr__pfet_01v8_7G6J3C_2 outp vdd clk sky130_fd_pr__pfet_01v8_7G6J3C_2/B
+ sky130_fd_pr__pfet_01v8_7G6J3C
Xsky130_fd_pr__pfet_01v8_7G6J3C_3 outn vdd clk sky130_fd_pr__pfet_01v8_7G6J3C_3/B
+ sky130_fd_pr__pfet_01v8_7G6J3C
Xsky130_fd_pr__pfet_01v8_7G6J3C_4 IN vdd clk sky130_fd_pr__pfet_01v8_7G6J3C_4/B sky130_fd_pr__pfet_01v8_7G6J3C
Xsky130_fd_pr__pfet_01v8_7G6J3C_5 IP vdd clk sky130_fd_pr__pfet_01v8_7G6J3C_5/B sky130_fd_pr__pfet_01v8_7G6J3C
.ends

