magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 682 542
<< pwell >>
rect 1 -19 643 163
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 109 137
rect 265 7 295 137
rect 349 7 379 137
rect 451 7 481 137
rect 535 7 565 137
<< scpmoshvt >>
rect 83 257 113 457
rect 265 257 295 457
rect 343 257 373 457
rect 463 257 493 457
rect 535 257 565 457
<< ndiff >>
rect 27 96 79 137
rect 27 62 35 96
rect 69 62 79 96
rect 27 7 79 62
rect 109 65 159 137
rect 213 123 265 137
rect 213 89 221 123
rect 255 89 265 123
rect 213 83 265 89
rect 109 55 161 65
rect 109 21 119 55
rect 153 21 161 55
rect 109 7 161 21
rect 215 7 265 83
rect 295 55 349 137
rect 295 21 305 55
rect 339 21 349 55
rect 295 7 349 21
rect 379 109 451 137
rect 379 75 389 109
rect 423 75 451 109
rect 379 7 451 75
rect 481 49 535 137
rect 481 15 491 49
rect 525 15 535 49
rect 481 7 535 15
rect 565 123 617 137
rect 565 89 575 123
rect 609 89 617 123
rect 565 55 617 89
rect 565 21 575 55
rect 609 21 617 55
rect 565 7 617 21
<< pdiff >>
rect 27 437 83 457
rect 27 403 39 437
rect 73 403 83 437
rect 27 369 83 403
rect 27 335 39 369
rect 73 335 83 369
rect 27 301 83 335
rect 27 267 39 301
rect 73 267 83 301
rect 27 257 83 267
rect 113 437 265 457
rect 113 403 126 437
rect 160 403 218 437
rect 252 403 265 437
rect 113 369 265 403
rect 113 335 126 369
rect 160 335 218 369
rect 252 335 265 369
rect 113 257 265 335
rect 295 257 343 457
rect 373 445 463 457
rect 373 411 383 445
rect 417 411 463 445
rect 373 377 463 411
rect 373 343 383 377
rect 417 343 463 377
rect 373 309 463 343
rect 373 275 383 309
rect 417 275 463 309
rect 373 257 463 275
rect 493 257 535 457
rect 565 445 617 457
rect 565 411 575 445
rect 609 411 617 445
rect 565 377 617 411
rect 565 343 575 377
rect 609 343 617 377
rect 565 309 617 343
rect 565 275 575 309
rect 609 275 617 309
rect 565 257 617 275
<< ndiffc >>
rect 35 62 69 96
rect 221 89 255 123
rect 119 21 153 55
rect 305 21 339 55
rect 389 75 423 109
rect 491 15 525 49
rect 575 89 609 123
rect 575 21 609 55
<< pdiffc >>
rect 39 403 73 437
rect 39 335 73 369
rect 39 267 73 301
rect 126 403 160 437
rect 218 403 252 437
rect 126 335 160 369
rect 218 335 252 369
rect 383 411 417 445
rect 383 343 417 377
rect 383 275 417 309
rect 575 411 609 445
rect 575 343 609 377
rect 575 275 609 309
<< poly >>
rect 83 457 113 483
rect 265 457 295 483
rect 343 457 373 483
rect 463 457 493 483
rect 535 457 565 483
rect 83 225 113 257
rect 265 225 295 257
rect 49 209 113 225
rect 49 175 59 209
rect 93 175 113 209
rect 49 173 113 175
rect 227 209 295 225
rect 227 175 237 209
rect 271 175 295 209
rect 49 159 109 173
rect 227 159 295 175
rect 343 225 373 257
rect 463 225 493 257
rect 343 209 397 225
rect 343 175 353 209
rect 387 175 397 209
rect 343 159 397 175
rect 439 209 493 225
rect 439 175 449 209
rect 483 175 493 209
rect 439 159 493 175
rect 535 225 565 257
rect 535 209 620 225
rect 535 175 570 209
rect 604 175 620 209
rect 535 159 620 175
rect 79 137 109 159
rect 265 137 295 159
rect 349 137 379 159
rect 451 137 481 159
rect 535 137 565 159
rect 79 -19 109 7
rect 265 -19 295 7
rect 349 -19 379 7
rect 451 -19 481 7
rect 535 -19 565 7
<< polycont >>
rect 59 175 93 209
rect 237 175 271 209
rect 353 175 387 209
rect 449 175 483 209
rect 570 175 604 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 644 521
rect 17 437 73 453
rect 17 403 39 437
rect 17 369 73 403
rect 17 335 39 369
rect 110 437 268 487
rect 110 403 126 437
rect 160 403 218 437
rect 252 403 268 437
rect 110 369 268 403
rect 110 335 126 369
rect 160 335 218 369
rect 252 335 268 369
rect 347 445 449 453
rect 347 411 383 445
rect 417 411 449 445
rect 575 445 627 487
rect 347 377 449 411
rect 347 343 383 377
rect 417 343 449 377
rect 17 301 73 335
rect 347 317 449 343
rect 347 309 425 317
rect 347 301 383 309
rect 17 267 39 301
rect 73 275 383 301
rect 417 275 425 309
rect 493 283 535 441
rect 73 267 425 275
rect 17 259 425 267
rect 17 209 93 225
rect 17 175 59 209
rect 17 159 93 175
rect 127 125 168 259
rect 459 249 535 283
rect 609 411 627 445
rect 575 377 627 411
rect 609 343 627 377
rect 575 309 627 343
rect 609 275 627 309
rect 575 251 627 275
rect 202 209 271 225
rect 202 175 237 209
rect 202 159 271 175
rect 305 209 397 225
rect 459 209 501 249
rect 305 175 353 209
rect 387 175 397 209
rect 433 175 449 209
rect 483 175 501 209
rect 535 209 627 215
rect 535 175 570 209
rect 604 175 627 209
rect 305 159 397 175
rect 421 125 627 133
rect 17 96 168 125
rect 17 62 35 96
rect 69 89 168 96
rect 202 123 627 125
rect 202 89 221 123
rect 255 109 575 123
rect 255 89 389 109
rect 17 33 69 62
rect 423 99 575 109
rect 423 75 444 99
rect 103 21 119 55
rect 153 21 305 55
rect 339 21 355 55
rect 389 16 444 75
rect 559 89 575 99
rect 609 89 627 123
rect 491 49 525 65
rect 559 55 627 89
rect 559 21 575 55
rect 609 21 627 55
rect 559 16 627 21
rect 491 -23 525 15
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 644 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
<< metal1 >>
rect 0 521 644 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 644 521
rect 0 456 644 487
rect 0 -23 644 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 644 -23
rect 0 -88 644 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 o221ai_1
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 497 317 531 351 0 FreeSans 400 0 0 0 A2
port 8 nsew
flabel locali s 397 385 431 419 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel locali s 213 181 247 215 0 FreeSans 400 0 0 0 B1
port 12 nsew
flabel locali s 29 181 63 215 0 FreeSans 400 0 0 0 C1
port 11 nsew
flabel locali s 581 181 615 215 0 FreeSans 400 0 0 0 A1
port 7 nsew
flabel locali s 397 317 431 351 0 FreeSans 400 0 0 0 Y
port 9 nsew
flabel locali s 341 181 375 215 0 FreeSans 400 0 0 0 B2
port 10 nsew
<< properties >>
string FIXED_BBOX 0 -40 644 504
string path 0.000 -1.000 16.100 -1.000 
<< end >>
