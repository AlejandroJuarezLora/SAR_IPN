* NGSPICE file created from DAC.ext - technology: sky130B

.subckt inv2 w_0_269# a_67_305# a_59_207# a_149_55# a_67_55# VSUBS
X0 a_67_55# a_59_207# a_149_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_149_55# a_59_207# a_67_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_67_305# a_59_207# a_149_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_149_55# a_59_207# a_67_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt decap_8 a_65_55# a_65_331# w_0_269# VSUBS
X0 a_65_55# a_65_331# a_65_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=2.89
X1 a_65_331# a_65_55# a_65_331# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=2.89
.ends

.subckt M1_3 a_207_n176# a_n29_n176# a_26_55# a_n328_55# a_89_n176# a_n446_55# a_n564_55#
+ a_n210_55# a_n501_n176# a_561_n176# a_n383_n176# a_498_55# a_144_55# a_443_n176#
+ a_n265_n176# a_262_55# a_380_55# a_n619_n176# a_n92_55# w_n757_n324# a_325_n176#
+ a_n147_n176#
X0 a_n383_n176# a_n446_55# a_n501_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 a_n29_n176# a_n92_55# a_n147_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 a_325_n176# a_262_55# a_207_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 a_561_n176# a_498_55# a_443_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X4 a_n265_n176# a_n328_55# a_n383_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X5 a_89_n176# a_26_55# a_n29_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 a_207_n176# a_144_55# a_89_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_n501_n176# a_n564_55# a_n619_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X8 a_n147_n176# a_n210_55# a_n265_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X9 a_443_n176# a_380_55# a_325_n176# w_n757_n324# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt M2_2 a_26_51# a_89_n171# a_n328_51# a_n446_51# a_n564_51# a_n501_n171# a_n210_51#
+ a_561_n171# a_n383_n171# a_498_51# a_443_n171# a_144_51# a_n265_n171# a_262_51#
+ a_n619_n171# a_380_51# a_n92_51# a_n721_n283# a_325_n171# a_n147_n171# a_207_n171#
+ a_n29_n171#
X0 a_89_n171# a_26_51# a_n29_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X1 a_207_n171# a_144_51# a_89_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 a_n147_n171# a_n210_51# a_n265_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 a_n501_n171# a_n564_51# a_n619_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X4 a_443_n171# a_380_51# a_325_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X5 a_n383_n171# a_n446_51# a_n501_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 a_n29_n171# a_n92_51# a_n147_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 a_325_n171# a_262_51# a_207_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X8 a_561_n171# a_498_51# a_443_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X9 a_n265_n171# a_n328_51# a_n383_n171# a_n721_n283# sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
.ends

.subckt inv_4 w_0_269# a_59_207# a_75_55# a_75_305# a_157_55# VSUBS
X0 a_75_55# a_59_207# a_157_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_75_305# a_59_207# a_157_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_157_55# a_59_207# a_75_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 a_157_55# a_59_207# a_75_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_157_55# a_59_207# a_75_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_75_305# a_59_207# a_157_55# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_75_55# a_59_207# a_157_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_157_55# a_59_207# a_75_305# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt decap_3 a_65_55# a_65_331# w_0_269# VSUBS
X0 a_65_55# a_65_331# a_65_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=0.59
X1 a_65_331# a_65_55# a_65_331# w_0_269# sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=0.59
.ends

.subckt sw_top out en m2_1158_361# m2_990_200# inv_4_1/w_0_269# vdd in vss
Xdecap_8_0 vss vdd inv_4_1/w_0_269# vss decap_8
XM1_3_0 out out m2_1158_361# m2_1158_361# in m2_1158_361# m2_1158_361# m2_1158_361#
+ out in in m2_1158_361# m2_1158_361# out out m2_1158_361# m2_1158_361# in m2_1158_361#
+ vdd in in M1_3
XM2_2_0 m2_990_200# in m2_990_200# m2_990_200# m2_990_200# out m2_990_200# in in m2_990_200#
+ out m2_990_200# out m2_990_200# in m2_990_200# m2_990_200# vss in in out out M2_2
Xinv_4_0 inv_4_1/w_0_269# m2_1158_361# vss vdd m2_990_200# vss inv_4
Xinv_4_1 inv_4_1/w_0_269# en vss vdd m2_1158_361# vss inv_4
Xdecap_3_0 vss vdd inv_4_1/w_0_269# vss decap_3
.ends

.subckt C7 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt DUMMY m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C6 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt CDUM m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C4 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C2 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C5 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C3 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C1 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt C0_1 m3_n450_n340# c1_n250_n240#
X0 c1_n250_n240# m3_n450_n340# sky130_fd_pr__cap_mim_m3_1 l=2 w=2
.ends

.subckt carray n5 n7 n6 n2 n3 n4 n1 n0 ndum top
XC7_121 n7 top C7
XC7_110 n7 top C7
XDUMMY_80 via23_4_712/m2_1_40# top DUMMY
XC6_20 n6 top C6
XC6_53 n6 top C6
XC6_31 n6 top C6
XC6_42 n6 top C6
XC7_122 n7 top C7
XC7_100 n7 top C7
XC7_111 n7 top C7
XDUMMY_81 via23_4_709/m2_1_40# top DUMMY
XDUMMY_70 via23_4_642/m2_1_40# top DUMMY
XC6_21 n6 top C6
XC6_10 n6 top C6
XC6_54 n6 top C6
XC6_32 n6 top C6
XC6_43 n6 top C6
XC6_0 n6 top C6
XC7_123 n7 top C7
XC7_101 n7 top C7
XC7_112 n7 top C7
XDUMMY_71 via23_4_641/m2_1_40# top DUMMY
XDUMMY_82 via23_4_439/m2_1_40# top DUMMY
XDUMMY_60 via23_4_448/m2_1_40# top DUMMY
XC6_44 n6 top C6
XC6_22 n6 top C6
XC6_55 n6 top C6
XC6_11 n6 top C6
XC6_33 n6 top C6
XC6_1 n6 top C6
XC7_124 n7 top C7
XC7_102 n7 top C7
XC7_113 n7 top C7
XDUMMY_72 via23_4_676/m2_1_40# top DUMMY
XDUMMY_83 via23_4_675/m2_1_40# top DUMMY
XDUMMY_61 via23_4_588/m2_1_40# top DUMMY
XDUMMY_50 via23_4_429/m2_1_40# top DUMMY
XC6_56 n6 top C6
XC6_12 n6 top C6
XC6_45 n6 top C6
XC6_23 n6 top C6
XC6_34 n6 top C6
XC6_2 n6 top C6
XCDUM_0 ndum top CDUM
XC7_103 n7 top C7
XC7_125 n7 top C7
XC7_114 n7 top C7
XDUMMY_73 via23_4_677/m2_1_40# top DUMMY
XDUMMY_62 via23_4_589/m2_1_40# top DUMMY
XDUMMY_40 via23_4_326/m2_1_40# top DUMMY
XDUMMY_51 via23_4_414/m2_1_40# top DUMMY
XC6_57 n6 top C6
XC6_24 n6 top C6
XC6_46 n6 top C6
XC6_13 n6 top C6
XC6_35 n6 top C6
XDUMMY_0 via23_4_3/m2_1_40# top DUMMY
XC6_3 n6 top C6
XC4_0 n4 top C4
XC7_104 n7 top C7
XC7_115 n7 top C7
XC7_126 n7 top C7
XDUMMY_74 via23_4_678/m2_1_40# top DUMMY
XDUMMY_63 via23_4_590/m2_1_40# top DUMMY
XDUMMY_30 via23_4_251/m2_1_40# top DUMMY
XDUMMY_52 via23_4_381/m2_1_40# top DUMMY
XDUMMY_41 via23_4_89/m2_1_40# top DUMMY
XC6_47 n6 top C6
XC6_14 n6 top C6
XC6_58 n6 top C6
XC6_25 n6 top C6
XC6_36 n6 top C6
XDUMMY_1 via23_4_9/m2_1_40# top DUMMY
XC7_90 n7 top C7
XC6_4 n6 top C6
XC4_1 n4 top C4
XC7_116 n7 top C7
XC7_105 n7 top C7
XC7_127 n7 top C7
XDUMMY_20 via23_4_199/m2_1_40# top DUMMY
XDUMMY_64 via23_4_584/m2_1_40# top DUMMY
XDUMMY_31 via23_4_245/m2_1_40# top DUMMY
XDUMMY_75 via23_4_704/m2_1_40# top DUMMY
XDUMMY_42 via23_4_366/m2_1_40# top DUMMY
XDUMMY_53 via23_4_449/m2_1_40# top DUMMY
XC6_26 n6 top C6
XC6_15 n6 top C6
XC6_59 n6 top C6
XC6_48 n6 top C6
XDUMMY_2 via23_4_1/m2_1_40# top DUMMY
XC6_37 n6 top C6
XC7_91 n7 top C7
XC7_80 n7 top C7
XC6_5 n6 top C6
XC4_2 n4 top C4
XC7_117 n7 top C7
XC7_106 n7 top C7
XDUMMY_76 via23_4_702/m2_1_40# top DUMMY
XDUMMY_65 via23_4_600/m2_1_40# top DUMMY
XDUMMY_32 via23_4_331/m2_1_40# top DUMMY
XDUMMY_21 via23_4_198/m2_1_40# top DUMMY
XDUMMY_43 via23_4_367/m2_1_40# top DUMMY
XDUMMY_54 via23_4_446/m2_1_40# top DUMMY
XDUMMY_10 via23_4_90/m2_1_40# top DUMMY
XC6_27 n6 top C6
XC6_16 n6 top C6
XC6_49 n6 top C6
XC6_38 n6 top C6
XDUMMY_3 via23_4_2/m2_1_40# top DUMMY
XC7_92 n7 top C7
XC7_81 n7 top C7
XC7_70 n7 top C7
XC6_6 n6 top C6
XC4_3 n4 top C4
XC7_118 n7 top C7
XC7_107 n7 top C7
XC2_0 n2 top C2
XDUMMY_66 via23_4_601/m2_1_40# top DUMMY
XDUMMY_33 via23_4_332/m2_1_40# top DUMMY
XDUMMY_22 via23_4_220/m2_1_40# top DUMMY
XDUMMY_77 via23_4_705/m2_1_40# top DUMMY
XDUMMY_44 via23_4_368/m2_1_40# top DUMMY
XDUMMY_55 via23_4_447/m2_1_40# top DUMMY
XDUMMY_11 via23_4_96/m2_1_40# top DUMMY
XC6_28 n6 top C6
XC6_17 n6 top C6
XC6_39 n6 top C6
XDUMMY_4 via23_4_20/m2_1_40# top DUMMY
XC7_60 n7 top C7
XC7_93 n7 top C7
XC7_82 n7 top C7
XC7_71 n7 top C7
XC6_7 n6 top C6
XC4_4 n4 top C4
XC7_119 n7 top C7
XC7_108 n7 top C7
XC2_1 n2 top C2
XDUMMY_78 via23_4_710/m2_1_40# top DUMMY
XDUMMY_67 via23_4_599/m2_1_40# top DUMMY
XDUMMY_34 via23_4_333/m2_1_40# top DUMMY
XDUMMY_23 via23_4_213/m2_1_40# top DUMMY
XDUMMY_45 via23_4_369/m2_1_40# top DUMMY
XDUMMY_56 via23_4_458/m2_1_40# top DUMMY
XDUMMY_12 via23_4_103/m2_1_40# top DUMMY
XC6_18 n6 top C6
XC6_29 n6 top C6
XDUMMY_5 via23_4_21/m2_1_40# top DUMMY
XC7_61 n7 top C7
XC7_94 n7 top C7
XC7_50 n7 top C7
XC7_72 n7 top C7
XC7_83 n7 top C7
XC6_8 n6 top C6
XC4_5 n4 top C4
XC7_109 n7 top C7
XC2_2 n2 top C2
XDUMMY_79 via23_4_711/m2_1_40# top DUMMY
XDUMMY_68 via23_4_598/m2_1_40# top DUMMY
XDUMMY_35 via23_4_347/m2_1_40# top DUMMY
XDUMMY_24 via23_4_229/m2_1_40# top DUMMY
XDUMMY_46 via23_4_378/m2_1_40# top DUMMY
XDUMMY_57 via23_4_455/m2_1_40# top DUMMY
XDUMMY_13 via23_4_91/m2_1_40# top DUMMY
XC6_19 n6 top C6
XDUMMY_6 via23_4_22/m2_1_40# top DUMMY
XC7_62 n7 top C7
XC7_40 n7 top C7
XC7_95 n7 top C7
XC7_51 n7 top C7
XC7_73 n7 top C7
XC7_84 n7 top C7
XC6_9 n6 top C6
XC4_6 n4 top C4
XC2_3 n2 top C2
XDUMMY_36 via23_4_354/m2_1_40# top DUMMY
XDUMMY_25 via23_4_228/m2_1_40# top DUMMY
XDUMMY_14 via23_4_94/m2_1_40# top DUMMY
XDUMMY_69 via23_4_635/m2_1_40# top DUMMY
XDUMMY_47 via23_4_379/m2_1_40# top DUMMY
XDUMMY_58 via23_4_459/m2_1_40# top DUMMY
XDUMMY_7 via23_4_23/m2_1_40# top DUMMY
XC7_41 n7 top C7
XC7_63 n7 top C7
XC7_96 n7 top C7
XC7_52 n7 top C7
XC7_30 n7 top C7
XC7_74 n7 top C7
XC7_85 n7 top C7
XC4_7 n4 top C4
XDUMMY_37 via23_4_345/m2_1_40# top DUMMY
XDUMMY_26 via23_4_230/m2_1_40# top DUMMY
XDUMMY_48 via23_4_380/m2_1_40# top DUMMY
XDUMMY_59 via23_4_460/m2_1_40# top DUMMY
XDUMMY_15 via23_4_117/m2_1_40# top DUMMY
XDUMMY_8 via23_4_87/m2_1_40# top DUMMY
XC7_97 n7 top C7
XC7_42 n7 top C7
XC7_53 n7 top C7
XC7_31 n7 top C7
XC7_86 n7 top C7
XC7_20 n7 top C7
XC7_64 n7 top C7
XC7_75 n7 top C7
XC4_10 n4 top C4
XC4_8 n4 top C4
XDUMMY_38 via23_4_346/m2_1_40# top DUMMY
XDUMMY_27 via23_4_218/m2_1_40# top DUMMY
XDUMMY_16 via23_4_111/m2_1_40# top DUMMY
XDUMMY_49 via23_4_419/m2_1_40# top DUMMY
XDUMMY_9 via23_4_88/m2_1_40# top DUMMY
XC7_98 n7 top C7
XC7_43 n7 top C7
XC7_54 n7 top C7
XC7_32 n7 top C7
XC7_87 n7 top C7
XC7_65 n7 top C7
XC7_10 n7 top C7
XC7_21 n7 top C7
XC7_76 n7 top C7
XC4_11 n4 top C4
XC4_9 n4 top C4
XDUMMY_39 via23_4_334/m2_1_40# top DUMMY
XDUMMY_28 via23_4_249/m2_1_40# top DUMMY
XDUMMY_17 via23_4_128/m2_1_40# top DUMMY
XC7_99 n7 top C7
XC7_33 n7 top C7
XC7_88 n7 top C7
XC7_55 n7 top C7
XC7_44 n7 top C7
XC7_66 n7 top C7
XC7_11 n7 top C7
XC7_77 n7 top C7
XC7_22 n7 top C7
XC4_12 n4 top C4
XDUMMY_29 via23_4_250/m2_1_40# top DUMMY
XDUMMY_18 via23_4_95/m2_1_40# top DUMMY
XC7_45 n7 top C7
XC7_56 n7 top C7
XC7_34 n7 top C7
XC7_89 n7 top C7
XC7_12 n7 top C7
XC7_23 n7 top C7
XC7_78 n7 top C7
XC7_67 n7 top C7
XC4_13 n4 top C4
XDUMMY_19 via23_4_200/m2_1_40# top DUMMY
XC7_46 n7 top C7
XC7_57 n7 top C7
XC7_24 n7 top C7
XC7_35 n7 top C7
XC7_13 n7 top C7
XC7_79 n7 top C7
XC7_68 n7 top C7
XC4_14 n4 top C4
XC7_36 n7 top C7
XC7_58 n7 top C7
XC7_47 n7 top C7
XC7_25 n7 top C7
XC7_14 n7 top C7
XC7_69 n7 top C7
XC4_15 n4 top C4
XC7_0 n7 top C7
XC7_37 n7 top C7
XC7_59 n7 top C7
XC7_26 n7 top C7
XC7_48 n7 top C7
XC7_15 n7 top C7
XC7_1 n7 top C7
XC7_38 n7 top C7
XC7_27 n7 top C7
XC7_49 n7 top C7
XC7_16 n7 top C7
XC7_2 n7 top C7
XC7_39 n7 top C7
XC7_28 n7 top C7
XC7_17 n7 top C7
XC7_3 n7 top C7
XC5_0 n5 top C5
XC7_29 n7 top C7
XC7_18 n7 top C7
XC7_4 n7 top C7
XC5_1 n5 top C5
XC7_19 n7 top C7
XC5_30 n5 top C5
XC7_5 n7 top C7
XC5_2 n5 top C5
XC5_31 n5 top C5
XC5_20 n5 top C5
XC7_6 n7 top C7
XC5_3 n5 top C5
XC3_0 n3 top C3
XC5_10 n5 top C5
XC5_21 n5 top C5
XC7_7 n7 top C7
XC5_4 n5 top C5
XC3_1 n3 top C3
XC5_22 n5 top C5
XC5_11 n5 top C5
XC7_8 n7 top C7
XC5_5 n5 top C5
XC3_2 n3 top C3
XC5_23 n5 top C5
XC7_9 n7 top C7
XC5_12 n5 top C5
XC5_6 n5 top C5
XC3_3 n3 top C3
XC1_0 n1 top C1
XC5_24 n5 top C5
XC5_13 n5 top C5
XC5_7 n5 top C5
XC3_4 n3 top C3
XC1_1 n1 top C1
XC5_25 n5 top C5
XC5_14 n5 top C5
XC5_8 n5 top C5
XC3_5 n3 top C3
XC5_15 n5 top C5
XC5_26 n5 top C5
XC5_9 n5 top C5
XC3_6 n3 top C3
XC5_16 n5 top C5
XC5_27 n5 top C5
XC3_7 n3 top C3
XC0_1_0 n0 top C0_1
XC5_28 n5 top C5
XC5_17 n5 top C5
XC6_60 n6 top C6
XC5_29 n5 top C5
XC5_18 n5 top C5
XC6_61 n6 top C6
XC6_50 n6 top C6
XC5_19 n5 top C5
XC6_51 n6 top C6
XC6_62 n6 top C6
XC6_40 n6 top C6
XC7_120 n7 top C7
XC6_63 n6 top C6
XC6_52 n6 top C6
XC6_30 n6 top C6
XC6_41 n6 top C6
.ends

.subckt DAC enb en_buf ctl1 ctl0 dum ctl3 ctl4 ctl5 ctl6 ctl7 ctl2 vdd vss sample
+ out vin
Xinv2_0 vdd vdd ctl7 carray_0/n7 vss vss inv2
Xinv2_1 vdd vdd ctl6 carray_0/n6 vss vss inv2
Xinv2_2 vdd vdd dum carray_0/ndum vss vss inv2
Xinv2_3 vdd vdd ctl0 carray_0/n0 vss vss inv2
Xinv2_4 vdd vdd ctl1 carray_0/n1 vss vss inv2
Xinv2_5 vdd vdd ctl5 carray_0/n5 vss vss inv2
Xinv2_6 vdd vdd ctl4 carray_0/n4 vss vss inv2
Xinv2_7 vdd vdd ctl2 carray_0/n2 vss vss inv2
Xinv2_8 vdd vdd ctl3 carray_0/n3 vss vss inv2
Xsw_top_0 out sample sw_top_0/m2_1158_361# sw_top_0/m2_990_200# vdd vdd vin vss sw_top
Xcarray_0 carray_0/n5 carray_0/n7 carray_0/n6 carray_0/n2 carray_0/n3 carray_0/n4
+ carray_0/n1 carray_0/n0 carray_0/ndum out carray
Xsw_top_1 out sample enb en_buf vdd vdd vin vss sw_top
Xsw_top_2 out sample enb en_buf vdd vdd vin vss sw_top
Xsw_top_3 out sample sw_top_3/m2_1158_361# sw_top_3/m2_990_200# vdd vdd vin vss sw_top
.ends

