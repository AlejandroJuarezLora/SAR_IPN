* NGSPICE file created from comparator_temp.ext - technology: sky130B

.subckt comparator trimb_4 trimb_1 trimb_0 trimb_2 trimb_3 clk vdd vp vn outp
+ outn vss trim_4 trim_3 trim_2 trim_1 trim_0
X0 trim_1.n3.t3 trimb_3.t0 vss.t29 vss.t28 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X1 vss.t1 trim_3.t0 trim_0.n3.t3 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X2 vss.t41 trim_4.t0 trim_0.n4.t7 vss.t40 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X3 vss.t27 trimb_3.t1 trim_1.n3.t2 vss.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X4 vss.t31 trim_4.t1 trim_0.n4.t6 vss.t30 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X5 vss.t69 trimb_4.t0 trim_1.n4.t7 vss.t68 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X6 trim_0.n3.t2 trim_3.t1 vss.t43 vss.t42 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X7 vss.t5 trim_4.t2 trim_0.n4.t5 vss.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X8 trim_1.n3.t1 trimb_3.t2 vss.t25 vss.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X9 vss.t14 trimb_4.t1 trim_1.n4.t6 vss.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X10 vss.t48 trim_2.t0 trim_0.n2 vss.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X11 comparator_core_0.diff vn.t0 trim_0.drain.t0 vss.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X12 trim_1.drain.t1 vp.t0 comparator_core_0.diff vss.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X13 vss.t62 trimb_2.t0 trim_1.n2 vss.t61 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X14 trim_0.n4.t4 trim_4.t3 vss.t35 vss.t34 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X15 trim_1.n4.t5 trimb_4.t2 vss.t39 vss.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X16 trim_1.drain.t2 clk.t0 vdd.t3 w_4048_2972# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X17 comparator_core_0.diff clk.t1 vss.t63 vss.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X18 trim_1.n4.t4 trimb_4.t3 vss.t21 vss.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X19 vdd.t0 outp.t3 outn.t1 w_4048_2972# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X20 outp.t2 outn.t3 vdd.t5 w_4048_2972# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X21 trim_0.n4.t3 trim_4.t4 vss.t60 vss.t59 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X22 outn.t0 clk.t2 vdd.t4 w_4048_2972# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X23 vss.t10 trim_3.t2 trim_0.n3.t1 vss.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X24 trim_0.drain.t1 outp.t4 outn.t2 vss.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X25 vss.t23 trimb_3.t3 trim_1.n3.t0 vss.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X26 vss.t50 trim_1.t0 trim_0.n1 vss.t49 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X27 trim_0.n2 trim_2.t1 vss.t54 vss.t53 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X28 outp.t0 outn.t4 trim_1.drain.t0 vss.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X29 vss.t52 trimb_1.t0 trim_1.n1 vss.t51 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X30 trim_1.n2 trimb_2.t1 vss.t65 vss.t64 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X31 vss.t12 trim_4.t5 trim_0.n4.t2 vss.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X32 vdd.t1 clk.t3 outp.t1 w_4048_2972# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X33 vss.t17 trimb_4.t4 trim_1.n4.t3 vss.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X34 trim_0.n4.t1 trim_4.t6 vss.t37 vss.t36 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X35 trim_1.n4.t2 trimb_4.t5 vss.t33 vss.t32 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X36 vdd.t2 clk.t4 trim_0.drain.t2 w_4048_2972# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X37 trim_1.n4.t1 trimb_4.t6 vss.t7 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X38 vss.t46 clk.t5 comparator_core_0.diff vss.t44 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X39 trim_0.n4.t0 trim_4.t7 vss.t19 vss.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X40 vss.t67 trimb_4.t7 trim_1.n4.t0 vss.t66 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X41 trim_0.n0 trim_0.t0 vss.t56 vss.t55 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X42 trim_0.n3.t0 trim_3.t3 vss.t3 vss.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X43 trim_1.n0 trimb_0.t0 vss.t58 vss.t57 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
R0 trimb_3.n0 trimb_3.t0 135.841
R1 trimb_3.n1 trimb_3.t1 135.841
R2 trimb_3.n1 trimb_3.t2 135.52
R3 trimb_3.n0 trimb_3.t3 135.52
R4 trimb_3 trimb_3.n2 2.48064
R5 trimb_3.n2 trimb_3.n0 0.0793043
R6 trimb_3.n2 trimb_3.n1 0.0793043
R7 vss.n143 vss.n142 1096.98
R8 vss.n505 vss.n504 1084.91
R9 vss.n109 vss.n108 292.5
R10 vss.n107 vss.n106 292.5
R11 vss.n105 vss.n104 292.5
R12 vss.n103 vss.n102 292.5
R13 vss.n101 vss.n100 292.5
R14 vss.n99 vss.n98 292.5
R15 vss.n97 vss.n96 292.5
R16 vss.n95 vss.n94 292.5
R17 vss.n93 vss.n92 292.5
R18 vss.n91 vss.n90 292.5
R19 vss.n89 vss.n88 292.5
R20 vss.n88 vss.n87 292.5
R21 vss.n86 vss.n85 292.5
R22 vss.n85 vss.n84 292.5
R23 vss.n83 vss.n82 292.5
R24 vss.n82 vss.n81 292.5
R25 vss.n80 vss.n79 292.5
R26 vss.n79 vss.n78 292.5
R27 vss.n77 vss.n76 292.5
R28 vss.n76 vss.n75 292.5
R29 vss.n74 vss.n73 292.5
R30 vss.n73 vss.n72 292.5
R31 vss.n71 vss.n70 292.5
R32 vss.n70 vss.n69 292.5
R33 vss.n68 vss.n67 292.5
R34 vss.n67 vss.n66 292.5
R35 vss.n533 vss.n532 292.5
R36 vss.n532 vss.n531 292.5
R37 vss.n536 vss.n535 292.5
R38 vss.n535 vss.n534 292.5
R39 vss.n539 vss.n538 292.5
R40 vss.n538 vss.n537 292.5
R41 vss.n542 vss.n541 292.5
R42 vss.n541 vss.n540 292.5
R43 vss.n545 vss.n544 292.5
R44 vss.n544 vss.n543 292.5
R45 vss.n548 vss.n547 292.5
R46 vss.n547 vss.n546 292.5
R47 vss.n551 vss.n550 292.5
R48 vss.n550 vss.n549 292.5
R49 vss.n553 vss.n552 292.5
R50 vss.n555 vss.n554 292.5
R51 vss.n557 vss.n556 292.5
R52 vss.n559 vss.n558 292.5
R53 vss.n561 vss.n560 292.5
R54 vss.n563 vss.n562 292.5
R55 vss.n565 vss.n564 292.5
R56 vss.n567 vss.n566 292.5
R57 vss.n569 vss.n568 292.5
R58 vss.n571 vss.n570 292.5
R59 vss.n416 vss.n415 292.5
R60 vss.n414 vss.n413 292.5
R61 vss.n412 vss.n411 292.5
R62 vss.n410 vss.n409 292.5
R63 vss.n408 vss.n407 292.5
R64 vss.n406 vss.n405 292.5
R65 vss.n404 vss.n403 292.5
R66 vss.n402 vss.n401 292.5
R67 vss.n400 vss.n399 292.5
R68 vss.n398 vss.n397 292.5
R69 vss.n396 vss.n395 292.5
R70 vss.n394 vss.n393 292.5
R71 vss.n392 vss.n391 292.5
R72 vss.n390 vss.n389 292.5
R73 vss.n388 vss.n387 292.5
R74 vss.n386 vss.n385 292.5
R75 vss.n384 vss.n383 292.5
R76 vss.n1 vss.n0 292.5
R77 vss.n3 vss.n2 292.5
R78 vss.n5 vss.n4 292.5
R79 vss.n7 vss.n6 292.5
R80 vss.n9 vss.n8 292.5
R81 vss.n11 vss.n10 292.5
R82 vss.n13 vss.n12 292.5
R83 vss.n15 vss.n14 292.5
R84 vss.n17 vss.n16 292.5
R85 vss.n19 vss.n18 292.5
R86 vss.n21 vss.n20 292.5
R87 vss.n23 vss.n22 292.5
R88 vss.n25 vss.n24 292.5
R89 vss.n27 vss.n26 292.5
R90 vss.n29 vss.n28 292.5
R91 vss.n31 vss.n30 292.5
R92 vss.n33 vss.n32 292.5
R93 vss.n494 vss.n493 292.5
R94 vss.n492 vss.n491 292.5
R95 vss.n450 vss.n449 292.5
R96 vss.n443 vss.n442 292.5
R97 vss.n436 vss.n435 292.5
R98 vss.n438 vss.n437 292.5
R99 vss.n133 vss.n132 292.5
R100 vss.n131 vss.n130 292.5
R101 vss.n460 vss.n459 292.5
R102 vss.n475 vss.n474 292.5
R103 vss.n428 vss.n427 292.5
R104 vss.n430 vss.n429 292.5
R105 vss.n485 vss.n484 292.5
R106 vss.n483 vss.n482 292.5
R107 vss.n481 vss.n480 292.5
R108 vss.n454 vss.n453 292.5
R109 vss.n456 vss.n455 292.5
R110 vss.n458 vss.n457 292.5
R111 vss.n372 vss.n371 292.5
R112 vss.n370 vss.n369 292.5
R113 vss.n368 vss.n367 292.5
R114 vss.n366 vss.n365 292.5
R115 vss.n364 vss.n363 292.5
R116 vss.n362 vss.n361 292.5
R117 vss.n360 vss.n359 292.5
R118 vss.n358 vss.n357 292.5
R119 vss.n356 vss.n355 292.5
R120 vss.n354 vss.n353 292.5
R121 vss.n352 vss.n351 292.5
R122 vss.n351 vss.n350 292.5
R123 vss.n349 vss.n348 292.5
R124 vss.n348 vss.n347 292.5
R125 vss.n346 vss.n345 292.5
R126 vss.n345 vss.n344 292.5
R127 vss.n343 vss.n342 292.5
R128 vss.n342 vss.n341 292.5
R129 vss.n340 vss.n339 292.5
R130 vss.n339 vss.n338 292.5
R131 vss.n337 vss.n336 292.5
R132 vss.n336 vss.n335 292.5
R133 vss.n334 vss.n333 292.5
R134 vss.n333 vss.n332 292.5
R135 vss.n331 vss.n330 292.5
R136 vss.n330 vss.n329 292.5
R137 vss.n328 vss.n327 292.5
R138 vss.n327 vss.n326 292.5
R139 vss.n325 vss.n324 292.5
R140 vss.n324 vss.n323 292.5
R141 vss.n322 vss.n321 292.5
R142 vss.n321 vss.n320 292.5
R143 vss.n319 vss.n318 292.5
R144 vss.n318 vss.n317 292.5
R145 vss.n316 vss.n315 292.5
R146 vss.n315 vss.n314 292.5
R147 vss.n313 vss.n312 292.5
R148 vss.n312 vss.n311 292.5
R149 vss.n310 vss.n309 292.5
R150 vss.n309 vss.n308 292.5
R151 vss.n307 vss.n306 292.5
R152 vss.n306 vss.n305 292.5
R153 vss.n304 vss.n303 292.5
R154 vss.n303 vss.n302 292.5
R155 vss.n301 vss.n300 292.5
R156 vss.n300 vss.n299 292.5
R157 vss.n298 vss.n297 292.5
R158 vss.n297 vss.n296 292.5
R159 vss.n295 vss.n294 292.5
R160 vss.n294 vss.n293 292.5
R161 vss.n292 vss.n291 292.5
R162 vss.n291 vss.n290 292.5
R163 vss.n289 vss.n288 292.5
R164 vss.n288 vss.n287 292.5
R165 vss.n286 vss.n285 292.5
R166 vss.n284 vss.n283 292.5
R167 vss.n282 vss.n281 292.5
R168 vss.n239 vss.n238 292.5
R169 vss.n161 vss.n160 292.5
R170 vss.n163 vss.n162 292.5
R171 vss.n165 vss.n164 292.5
R172 vss.n167 vss.n166 292.5
R173 vss.n169 vss.n168 292.5
R174 vss.n171 vss.n170 292.5
R175 vss.n173 vss.n172 292.5
R176 vss.n175 vss.n174 292.5
R177 vss.n177 vss.n176 292.5
R178 vss.n179 vss.n178 292.5
R179 vss.n181 vss.n180 292.5
R180 vss.n183 vss.n182 292.5
R181 vss.n185 vss.n184 292.5
R182 vss.n187 vss.n186 292.5
R183 vss.n189 vss.n188 292.5
R184 vss.n191 vss.n190 292.5
R185 vss.n193 vss.n192 292.5
R186 vss.n195 vss.n194 292.5
R187 vss.n197 vss.n196 292.5
R188 vss.n199 vss.n198 292.5
R189 vss.n201 vss.n200 292.5
R190 vss.n203 vss.n202 292.5
R191 vss.n205 vss.n204 292.5
R192 vss.n207 vss.n206 292.5
R193 vss.n209 vss.n208 292.5
R194 vss.n211 vss.n210 292.5
R195 vss.n213 vss.n212 292.5
R196 vss.n215 vss.n214 292.5
R197 vss.n217 vss.n216 292.5
R198 vss.n219 vss.n218 292.5
R199 vss.n221 vss.n220 292.5
R200 vss.n223 vss.n222 292.5
R201 vss.n225 vss.n224 292.5
R202 vss.n227 vss.n226 292.5
R203 vss.n154 vss.t18 197.065
R204 vss.n516 vss.t6 196.667
R205 vss.n251 vss.t2 195.952
R206 vss.n54 vss.t28 195.556
R207 vss.n34 vss.n33 163.766
R208 vss.n518 vss.n517 157.778
R209 vss.n56 vss.n55 157.778
R210 vss.n156 vss.n155 156.576
R211 vss.n444 vss.n443 155.482
R212 vss.n439 vss.n438 150.213
R213 vss.n504 vss.n500 147.875
R214 vss.n500 vss.t8 147.875
R215 vss.n138 vss.t15 147.875
R216 vss.n142 vss.n138 147.875
R217 vss.n463 vss.n462 146.447
R218 vss.n478 vss.n477 144.189
R219 vss.n417 vss.n416 144.189
R220 vss.n228 vss.n227 144.189
R221 vss.n451 vss.n450 140.968
R222 vss.n495 vss.n494 135.697
R223 vss.n572 vss.n571 131.766
R224 vss.n373 vss.n372 131.766
R225 vss.n110 vss.n109 125.742
R226 vss.n282 vss.n280 125.742
R227 vss.n141 vss.n139 117.719
R228 vss.n503 vss.n502 117.719
R229 vss.n503 vss.n501 117.719
R230 vss.n141 vss.n140 117.719
R231 vss.n430 vss.n428 102.606
R232 vss.n133 vss.n131 102.606
R233 vss.n486 vss.n479 100.216
R234 vss.n465 vss.n464 100.216
R235 vss.n504 vss.n503 87.3927
R236 vss.n142 vss.n141 87.3927
R237 vss.n250 vss.n249 75.709
R238 vss.n146 vss.n145 75.709
R239 vss.n148 vss.n147 75.709
R240 vss.n151 vss.n150 75.709
R241 vss.n153 vss.n152 75.709
R242 vss.n53 vss.n52 75.5561
R243 vss.n51 vss.n50 75.5561
R244 vss.n49 vss.n48 75.5561
R245 vss.n47 vss.n46 75.5561
R246 vss.n46 vss.n45 75.5561
R247 vss.n45 vss.n44 75.5561
R248 vss.n508 vss.n507 75.5561
R249 vss.n510 vss.n509 75.5561
R250 vss.n513 vss.n512 75.5561
R251 vss.n515 vss.n514 75.5561
R252 vss.t26 vss.n47 68.8894
R253 vss.n149 vss.t30 65.6888
R254 vss.t59 vss.n149 65.6888
R255 vss.n511 vss.t68 65.5561
R256 vss.t20 vss.n511 65.5561
R257 vss.n137 vss.n136 63.7358
R258 vss.n499 vss.n433 63.7358
R259 vss.n131 vss.n129 57.3393
R260 vss.n247 vss.n246 52.1476
R261 vss.t11 vss.n144 50.1017
R262 vss.t16 vss.n506 50.0005
R263 vss.n290 vss.t42 48.9884
R264 vss.t24 vss.n49 48.8894
R265 vss.n314 vss.t47 47.875
R266 vss.n44 vss.t64 47.7783
R267 vss.n249 vss.t9 46.7616
R268 vss.n52 vss.t22 46.6672
R269 vss.n157 vss.n127 46.3534
R270 vss.n147 vss.t34 45.6483
R271 vss.t40 vss.n151 45.6483
R272 vss.n509 vss.t38 45.5561
R273 vss.t66 vss.n513 45.5561
R274 vss.n428 vss.n426 45.268
R275 vss.n425 vss.n424 45.268
R276 vss.n252 vss.n247 42.3273
R277 vss.t45 vss.n128 42.2502
R278 vss.n522 vss.n521 40.5593
R279 vss.n57 vss.n43 40.5593
R280 vss.t44 vss.n425 33.1967
R281 vss.n465 vss.n458 30.5684
R282 vss.t34 vss.n146 30.0612
R283 vss.n152 vss.t40 30.0612
R284 vss.t38 vss.n508 30.0005
R285 vss.n514 vss.t66 30.0005
R286 vss.t9 vss.n248 28.9479
R287 vss.t22 vss.n51 28.8894
R288 vss.n486 vss.n485 28.3093
R289 vss.n308 vss.t53 27.8345
R290 vss.n84 vss.t61 27.7783
R291 vss.n520 vss.n519 27.6046
R292 vss.n42 vss.n41 27.6046
R293 vss.n521 vss.n520 27.6046
R294 vss.n43 vss.n42 27.6046
R295 vss.n332 vss.t49 26.7211
R296 vss.n50 vss.t24 26.6672
R297 vss.n531 vss.t51 26.6672
R298 vss.n582 vss.t14 26.601
R299 vss.n578 vss.t7 26.601
R300 vss.n264 vss.t5 26.5994
R301 vss.n122 vss.t19 26.5994
R302 vss.n145 vss.t11 25.6078
R303 vss.t18 vss.n153 25.6078
R304 vss.n479 vss.n478 25.6005
R305 vss.n477 vss.n476 25.6005
R306 vss.n476 vss.n475 25.6005
R307 vss.n461 vss.n460 25.6005
R308 vss.n462 vss.n461 25.6005
R309 vss.n464 vss.n463 25.6005
R310 vss.n485 vss.n483 25.6005
R311 vss.n483 vss.n481 25.6005
R312 vss.n456 vss.n454 25.6005
R313 vss.n458 vss.n456 25.6005
R314 vss.n494 vss.n492 25.6005
R315 vss.n438 vss.n436 25.6005
R316 vss.n109 vss.n107 25.6005
R317 vss.n107 vss.n105 25.6005
R318 vss.n105 vss.n103 25.6005
R319 vss.n103 vss.n101 25.6005
R320 vss.n101 vss.n99 25.6005
R321 vss.n99 vss.n97 25.6005
R322 vss.n97 vss.n95 25.6005
R323 vss.n95 vss.n93 25.6005
R324 vss.n93 vss.n91 25.6005
R325 vss.n91 vss.n89 25.6005
R326 vss.n89 vss.n86 25.6005
R327 vss.n86 vss.n83 25.6005
R328 vss.n83 vss.n80 25.6005
R329 vss.n80 vss.n77 25.6005
R330 vss.n77 vss.n74 25.6005
R331 vss.n74 vss.n71 25.6005
R332 vss.n71 vss.n68 25.6005
R333 vss.n536 vss.n533 25.6005
R334 vss.n539 vss.n536 25.6005
R335 vss.n542 vss.n539 25.6005
R336 vss.n545 vss.n542 25.6005
R337 vss.n548 vss.n545 25.6005
R338 vss.n551 vss.n548 25.6005
R339 vss.n553 vss.n551 25.6005
R340 vss.n555 vss.n553 25.6005
R341 vss.n557 vss.n555 25.6005
R342 vss.n559 vss.n557 25.6005
R343 vss.n561 vss.n559 25.6005
R344 vss.n563 vss.n561 25.6005
R345 vss.n565 vss.n563 25.6005
R346 vss.n567 vss.n565 25.6005
R347 vss.n569 vss.n567 25.6005
R348 vss.n571 vss.n569 25.6005
R349 vss.n33 vss.n31 25.6005
R350 vss.n31 vss.n29 25.6005
R351 vss.n29 vss.n27 25.6005
R352 vss.n27 vss.n25 25.6005
R353 vss.n25 vss.n23 25.6005
R354 vss.n23 vss.n21 25.6005
R355 vss.n21 vss.n19 25.6005
R356 vss.n19 vss.n17 25.6005
R357 vss.n17 vss.n15 25.6005
R358 vss.n15 vss.n13 25.6005
R359 vss.n13 vss.n11 25.6005
R360 vss.n11 vss.n9 25.6005
R361 vss.n9 vss.n7 25.6005
R362 vss.n7 vss.n5 25.6005
R363 vss.n5 vss.n3 25.6005
R364 vss.n3 vss.n1 25.6005
R365 vss.n386 vss.n384 25.6005
R366 vss.n388 vss.n386 25.6005
R367 vss.n390 vss.n388 25.6005
R368 vss.n392 vss.n390 25.6005
R369 vss.n394 vss.n392 25.6005
R370 vss.n396 vss.n394 25.6005
R371 vss.n398 vss.n396 25.6005
R372 vss.n400 vss.n398 25.6005
R373 vss.n402 vss.n400 25.6005
R374 vss.n404 vss.n402 25.6005
R375 vss.n406 vss.n404 25.6005
R376 vss.n408 vss.n406 25.6005
R377 vss.n410 vss.n408 25.6005
R378 vss.n412 vss.n410 25.6005
R379 vss.n414 vss.n412 25.6005
R380 vss.n416 vss.n414 25.6005
R381 vss.n284 vss.n282 25.6005
R382 vss.n286 vss.n284 25.6005
R383 vss.n289 vss.n286 25.6005
R384 vss.n292 vss.n289 25.6005
R385 vss.n295 vss.n292 25.6005
R386 vss.n298 vss.n295 25.6005
R387 vss.n301 vss.n298 25.6005
R388 vss.n304 vss.n301 25.6005
R389 vss.n307 vss.n304 25.6005
R390 vss.n310 vss.n307 25.6005
R391 vss.n313 vss.n310 25.6005
R392 vss.n316 vss.n313 25.6005
R393 vss.n319 vss.n316 25.6005
R394 vss.n322 vss.n319 25.6005
R395 vss.n325 vss.n322 25.6005
R396 vss.n328 vss.n325 25.6005
R397 vss.n331 vss.n328 25.6005
R398 vss.n334 vss.n331 25.6005
R399 vss.n337 vss.n334 25.6005
R400 vss.n340 vss.n337 25.6005
R401 vss.n343 vss.n340 25.6005
R402 vss.n346 vss.n343 25.6005
R403 vss.n349 vss.n346 25.6005
R404 vss.n352 vss.n349 25.6005
R405 vss.n354 vss.n352 25.6005
R406 vss.n356 vss.n354 25.6005
R407 vss.n358 vss.n356 25.6005
R408 vss.n360 vss.n358 25.6005
R409 vss.n362 vss.n360 25.6005
R410 vss.n364 vss.n362 25.6005
R411 vss.n366 vss.n364 25.6005
R412 vss.n368 vss.n366 25.6005
R413 vss.n370 vss.n368 25.6005
R414 vss.n372 vss.n370 25.6005
R415 vss.n163 vss.n161 25.6005
R416 vss.n165 vss.n163 25.6005
R417 vss.n167 vss.n165 25.6005
R418 vss.n169 vss.n167 25.6005
R419 vss.n171 vss.n169 25.6005
R420 vss.n173 vss.n171 25.6005
R421 vss.n175 vss.n173 25.6005
R422 vss.n177 vss.n175 25.6005
R423 vss.n179 vss.n177 25.6005
R424 vss.n181 vss.n179 25.6005
R425 vss.n183 vss.n181 25.6005
R426 vss.n185 vss.n183 25.6005
R427 vss.n187 vss.n185 25.6005
R428 vss.n189 vss.n187 25.6005
R429 vss.n191 vss.n189 25.6005
R430 vss.n193 vss.n191 25.6005
R431 vss.n195 vss.n193 25.6005
R432 vss.n197 vss.n195 25.6005
R433 vss.n199 vss.n197 25.6005
R434 vss.n201 vss.n199 25.6005
R435 vss.n203 vss.n201 25.6005
R436 vss.n205 vss.n203 25.6005
R437 vss.n207 vss.n205 25.6005
R438 vss.n209 vss.n207 25.6005
R439 vss.n211 vss.n209 25.6005
R440 vss.n213 vss.n211 25.6005
R441 vss.n215 vss.n213 25.6005
R442 vss.n217 vss.n215 25.6005
R443 vss.n219 vss.n217 25.6005
R444 vss.n221 vss.n219 25.6005
R445 vss.n223 vss.n221 25.6005
R446 vss.n225 vss.n223 25.6005
R447 vss.n227 vss.n225 25.6005
R448 vss.n507 vss.t16 25.5561
R449 vss.t6 vss.n515 25.5561
R450 vss.n126 vss.n125 24.962
R451 vss.n127 vss.n126 24.962
R452 vss.n426 vss.t44 24.1432
R453 vss.n441 vss.t63 23.9627
R454 vss.n440 vss.t46 23.9618
R455 vss.n280 vss.n237 18.0711
R456 vss.n271 vss.t3 17.4005
R457 vss.n271 vss.t10 17.4005
R458 vss.n269 vss.t43 17.4005
R459 vss.n269 vss.t1 17.4005
R460 vss.n267 vss.t54 17.4005
R461 vss.n267 vss.t48 17.4005
R462 vss.n265 vss.t56 17.4005
R463 vss.n265 vss.t50 17.4005
R464 vss.n262 vss.t37 17.4005
R465 vss.n262 vss.t12 17.4005
R466 vss.n260 vss.t35 17.4005
R467 vss.n260 vss.t31 17.4005
R468 vss.n258 vss.t60 17.4005
R469 vss.n258 vss.t41 17.4005
R470 vss.n121 vss.t21 17.4005
R471 vss.n121 vss.t67 17.4005
R472 vss.n120 vss.t39 17.4005
R473 vss.n120 vss.t69 17.4005
R474 vss.n119 vss.t33 17.4005
R475 vss.n119 vss.t17 17.4005
R476 vss.n118 vss.t58 17.4005
R477 vss.n118 vss.t52 17.4005
R478 vss.n117 vss.t65 17.4005
R479 vss.n117 vss.t62 17.4005
R480 vss.n116 vss.t25 17.4005
R481 vss.n116 vss.t27 17.4005
R482 vss.n115 vss.t29 17.4005
R483 vss.n115 vss.t23 17.4005
R484 vss.n135 vss.n134 16.8818
R485 vss.n432 vss.n431 16.8818
R486 vss.n136 vss.n135 16.8818
R487 vss.n433 vss.n432 16.8818
R488 vss.n418 vss.n417 16.5652
R489 vss.n35 vss.n34 16.5652
R490 vss.n240 vss.n239 16.1887
R491 vss.n229 vss.n228 16.1887
R492 vss.t15 vss.n133 15.0897
R493 vss.n344 vss.t4 14.4742
R494 vss.n543 vss.t13 14.4449
R495 vss.n144 vss.n143 13.3608
R496 vss.n506 vss.n505 13.3338
R497 vss.t30 vss.n148 10.0207
R498 vss.n150 vss.t59 10.0207
R499 vss.t68 vss.n510 10.0005
R500 vss.n512 vss.t20 10.0005
R501 vss.n241 vss.n240 9.31144
R502 vss.n230 vss.n229 9.31144
R503 vss.n36 vss.n35 9.31039
R504 vss.n419 vss.n418 9.31039
R505 vss.n524 vss.n523 9.3005
R506 vss.n523 vss.n522 9.3005
R507 vss.n59 vss.n58 9.3005
R508 vss.n58 vss.n57 9.3005
R509 vss.n138 vss.n137 9.3005
R510 vss.n499 vss.n498 9.3005
R511 vss.n500 vss.n499 9.3005
R512 vss.n255 vss.n254 9.3005
R513 vss.n254 vss.n253 9.3005
R514 vss.n159 vss.n158 9.3005
R515 vss.n158 vss.n157 9.3005
R516 vss.n586 vss.n115 9.20119
R517 vss.n585 vss.n116 9.20119
R518 vss.n584 vss.n117 9.20119
R519 vss.n583 vss.n118 9.20119
R520 vss.n581 vss.n119 9.20119
R521 vss.n580 vss.n120 9.20119
R522 vss.n579 vss.n121 9.20119
R523 vss.n272 vss.n271 9.19943
R524 vss.n270 vss.n269 9.19943
R525 vss.n268 vss.n267 9.19943
R526 vss.n266 vss.n265 9.19943
R527 vss.n263 vss.n262 9.19943
R528 vss.n261 vss.n260 9.19943
R529 vss.n259 vss.n258 9.19943
R530 vss.n421 vss.n420 9.0005
R531 vss.n38 vss.n37 9.0005
R532 vss.n243 vss.n242 9.0005
R533 vss.n232 vss.n231 9.0005
R534 vss.t2 vss.n250 8.90738
R535 vss.t28 vss.n53 8.88939
R536 vss.n252 vss.n251 8.49312
R537 vss.n293 vss.t0 6.68066
R538 vss.n326 vss.t55 6.68066
R539 vss.n48 vss.t26 6.66717
R540 vss.n69 vss.t57 6.66717
R541 vss.t8 vss.n430 6.03617
R542 vss.n350 vss.t36 5.5673
R543 vss.n549 vss.t32 5.55606
R544 vss.n522 vss.n518 5.01811
R545 vss.n57 vss.n56 5.01748
R546 vss.n157 vss.n156 4.97926
R547 vss.n452 vss.n444 4.57427
R548 vss.n490 vss.n439 4.57427
R549 vss.n573 vss.n572 4.57427
R550 vss.n111 vss.n110 4.57427
R551 vss.n280 vss.n279 4.57427
R552 vss.n374 vss.n373 4.57427
R553 vss.n156 vss.n154 4.18956
R554 vss.n518 vss.n516 4.15288
R555 vss.n56 vss.n54 4.15252
R556 vss.n448 vss.n447 4.14168
R557 vss.n498 vss.n497 4.14168
R558 vss.n577 vss.n382 4.02849
R559 vss.n423 vss.n422 3.76521
R560 vss.n40 vss.n39 3.76521
R561 vss.n124 vss.n123 3.38874
R562 vss.n129 vss.t45 3.01833
R563 vss.n254 vss.n245 3.01226
R564 vss.n158 vss.n124 3.01226
R565 vss.n278 vss.n277 3.0005
R566 vss.n61 vss.n60 3.0005
R567 vss.n113 vss.n112 3.0005
R568 vss.n526 vss.n525 3.0005
R569 vss.n575 vss.n574 3.0005
R570 vss.n234 vss.n233 3.0005
R571 vss.n378 vss.n377 3.0005
R572 vss.n451 vss.n448 2.65111
R573 vss.n498 vss.n495 2.65111
R574 vss.n523 vss.n423 2.63579
R575 vss.n58 vss.n40 2.63579
R576 vss.n447 vss.n446 2.25932
R577 vss.n497 vss.n496 2.25932
R578 vss.n382 vss.n381 2.21752
R579 vss.n452 vss.n451 2.05223
R580 vss.n495 vss.n490 2.05223
R581 vss.n487 vss.n486 1.84239
R582 vss.n466 vss.n465 1.84237
R583 vss.n381 vss.n380 1.81065
R584 vss.n490 vss.n489 1.77862
R585 vss.n468 vss.n452 1.4761
R586 vss vss.n382 1.47472
R587 vss.n268 vss.n266 0.80675
R588 vss.n270 vss.n268 0.80675
R589 vss.n585 vss.n584 0.80675
R590 vss.n584 vss.n583 0.80675
R591 vss.n381 vss 0.752104
R592 vss.n472 vss.n471 0.673937
R593 vss.n471 vss.n470 0.673937
R594 vss.n253 vss.n252 0.67388
R595 vss.n266 vss.n264 0.560917
R596 vss.n583 vss.n582 0.560917
R597 vss vss.n272 0.448417
R598 vss.n471 vss 0.41925
R599 vss.n259 vss.n122 0.408833
R600 vss.n261 vss.n259 0.408833
R601 vss.n263 vss.n261 0.408833
R602 vss.n264 vss.n263 0.408833
R603 vss.n272 vss.n270 0.408833
R604 vss.n586 vss.n585 0.408833
R605 vss.n582 vss.n581 0.408833
R606 vss.n581 vss.n580 0.408833
R607 vss.n580 vss.n579 0.408833
R608 vss.n579 vss.n578 0.408833
R609 vss.n587 vss.n586 0.385917
R610 vss.n380 vss.n379 0.359081
R611 vss.n587 vss.n114 0.358301
R612 vss.n577 vss.n576 0.358301
R613 vss.n273 vss 0.296581
R614 vss.n380 vss.n122 0.142167
R615 vss.n578 vss.n577 0.142167
R616 vss.n489 vss.n488 0.0697748
R617 vss vss.n587 0.063
R618 vss.n468 vss.n467 0.0589808
R619 vss.n469 vss.n468 0.0581328
R620 vss.n257 vss.n256 0.0525833
R621 vss.n65 vss.n64 0.0525833
R622 vss.n530 vss.n529 0.0525833
R623 vss.n376 vss.n375 0.0525833
R624 vss.n489 vss.n473 0.0467812
R625 vss.n278 vss.n257 0.0421667
R626 vss.n377 vss.n376 0.0421667
R627 vss.n112 vss.n65 0.0400833
R628 vss.n574 vss.n530 0.0400833
R629 vss.n276 vss.n275 0.0395625
R630 vss.n63 vss.n62 0.0395625
R631 vss.n528 vss.n527 0.0395625
R632 vss.n236 vss.n235 0.0395625
R633 vss.n256 vss.n255 0.0338333
R634 vss.n277 vss.n276 0.03175
R635 vss.n473 vss.n472 0.03175
R636 vss.n470 vss.n469 0.03175
R637 vss.n62 vss.n61 0.03175
R638 vss.n527 vss.n526 0.03175
R639 vss.n378 vss.n236 0.03175
R640 vss.n275 vss.n274 0.0301875
R641 vss.n488 vss.n487 0.0301875
R642 vss.n467 vss.n466 0.0301875
R643 vss.n113 vss.n63 0.0301875
R644 vss.n575 vss.n528 0.0301875
R645 vss.n235 vss.n234 0.0301875
R646 vss.n114 vss.n113 0.022812
R647 vss.n576 vss.n575 0.022812
R648 vss.n277 vss.n273 0.0220368
R649 vss.n379 vss.n378 0.0220368
R650 vss.n490 vss.n440 0.0201429
R651 vss.n452 vss.n445 0.0201429
R652 vss.n452 vss.n441 0.01925
R653 vss.n243 vss.n241 0.0113746
R654 vss.n232 vss.n230 0.0113746
R655 vss.n490 vss.n434 0.0103652
R656 vss.n38 vss.n36 0.0103391
R657 vss.n421 vss.n419 0.0103391
R658 vss.n279 vss.n278 0.00883333
R659 vss.n244 vss.n243 0.00883333
R660 vss.n60 vss.n38 0.00883333
R661 vss.n60 vss.n59 0.00883333
R662 vss.n112 vss.n111 0.00883333
R663 vss.n525 vss.n421 0.00883333
R664 vss.n525 vss.n524 0.00883333
R665 vss.n574 vss.n573 0.00883333
R666 vss.n377 vss.n374 0.00883333
R667 vss.n233 vss.n232 0.00883333
R668 vss.n255 vss.n244 0.00675
R669 vss.n233 vss.n159 0.00675
R670 trim_1.n3.n1 trim_1.n3.t2 25.4402
R671 trim_1.n3.n2 trim_1.n3.t3 24.9249
R672 trim_1.n3.n0 trim_1.n3.t0 17.4005
R673 trim_1.n3.n0 trim_1.n3.t1 17.4005
R674 trim_1.n3.n1 trim_1.n3.n0 7.52492
R675 trim_1.n3 trim_1.n3.n2 1.4543
R676 trim_1.n3.n2 trim_1.n3.n1 0.516804
R677 trim_3.n0 trim_3.t3 135.841
R678 trim_3.n1 trim_3.t0 135.841
R679 trim_3.n1 trim_3.t1 135.52
R680 trim_3.n0 trim_3.t2 135.52
R681 trim_3 trim_3.n2 2.56687
R682 trim_3.n2 trim_3.n0 0.0793043
R683 trim_3.n2 trim_3.n1 0.0793043
R684 trim_0.n3.n1 trim_0.n3.t3 25.4412
R685 trim_0.n3.n2 trim_0.n3.t0 24.9249
R686 trim_0.n3.n0 trim_0.n3.t1 17.4005
R687 trim_0.n3.n0 trim_0.n3.t2 17.4005
R688 trim_0.n3.n1 trim_0.n3.n0 7.52464
R689 trim_0.n3 trim_0.n3.n2 1.3293
R690 trim_0.n3.n2 trim_0.n3.n1 0.516804
R691 trim_4.n0 trim_4.t2 135.841
R692 trim_4.n3 trim_4.t7 135.841
R693 trim_4.n3 trim_4.t0 135.52
R694 trim_4.n4 trim_4.t4 135.52
R695 trim_4.n5 trim_4.t1 135.52
R696 trim_4.n2 trim_4.t3 135.52
R697 trim_4.n1 trim_4.t5 135.52
R698 trim_4.n0 trim_4.t6 135.52
R699 trim_4 trim_4.n6 2.56687
R700 trim_4.n1 trim_4.n0 0.321152
R701 trim_4.n2 trim_4.n1 0.321152
R702 trim_4.n5 trim_4.n4 0.321152
R703 trim_4.n4 trim_4.n3 0.321152
R704 trim_4.n6 trim_4.n2 0.0793043
R705 trim_4.n6 trim_4.n5 0.0793043
R706 trim_0.n4.n5 trim_0.n4.t7 17.4005
R707 trim_0.n4.n5 trim_0.n4.t0 17.4005
R708 trim_0.n4.n0 trim_0.n4.t5 17.4005
R709 trim_0.n4.n0 trim_0.n4.t1 17.4005
R710 trim_0.n4.n1 trim_0.n4.t2 17.4005
R711 trim_0.n4.n1 trim_0.n4.t4 17.4005
R712 trim_0.n4.n3 trim_0.n4.t6 17.4005
R713 trim_0.n4.n3 trim_0.n4.t3 17.4005
R714 trim_0.n4.n2 trim_0.n4.n0 8.04122
R715 trim_0.n4.n2 trim_0.n4.n1 7.52492
R716 trim_0.n4.n4 trim_0.n4.n3 7.52464
R717 trim_0.n4 trim_0.n4.n5 7.46242
R718 trim_0.n4 trim_0.n4.n4 0.579304
R719 trim_0.n4.n4 trim_0.n4.n2 0.516804
R720 trimb_4.n0 trimb_4.t1 135.841
R721 trimb_4.n3 trimb_4.t6 135.841
R722 trimb_4.n3 trimb_4.t7 135.52
R723 trimb_4.n4 trimb_4.t3 135.52
R724 trimb_4.n5 trimb_4.t0 135.52
R725 trimb_4.n2 trimb_4.t2 135.52
R726 trimb_4.n1 trimb_4.t4 135.52
R727 trimb_4.n0 trimb_4.t5 135.52
R728 trimb_4 trimb_4.n6 2.48064
R729 trimb_4.n1 trimb_4.n0 0.321152
R730 trimb_4.n2 trimb_4.n1 0.321152
R731 trimb_4.n5 trimb_4.n4 0.321152
R732 trimb_4.n4 trimb_4.n3 0.321152
R733 trimb_4.n6 trimb_4.n2 0.0793043
R734 trimb_4.n6 trimb_4.n5 0.0793043
R735 trim_1.n4.n0 trim_1.n4.t0 17.4005
R736 trim_1.n4.n0 trim_1.n4.t1 17.4005
R737 trim_1.n4.n1 trim_1.n4.t7 17.4005
R738 trim_1.n4.n1 trim_1.n4.t4 17.4005
R739 trim_1.n4.n2 trim_1.n4.t3 17.4005
R740 trim_1.n4.n2 trim_1.n4.t5 17.4005
R741 trim_1.n4.n3 trim_1.n4.t6 17.4005
R742 trim_1.n4.n3 trim_1.n4.t2 17.4005
R743 trim_1.n4.n4 trim_1.n4.n3 8.04069
R744 trim_1.n4.n6 trim_1.n4.n0 7.52492
R745 trim_1.n4.n5 trim_1.n4.n1 7.52492
R746 trim_1.n4.n4 trim_1.n4.n2 7.52492
R747 trim_1.n4.n6 trim_1.n4.n5 0.516804
R748 trim_1.n4.n5 trim_1.n4.n4 0.516804
R749 trim_1.n4 trim_1.n4.n6 0.063
R750 trim_2.n0 trim_2.t1 135.6
R751 trim_2.n0 trim_2.t0 135.6
R752 trim_2 trim_2.n0 2.56687
R753 vn.n1 vn.t0 138.87
R754 vn vn.n7 1.64973
R755 vn.n5 vn.n1 0.750898
R756 vn.n6 vn.n5 0.513756
R757 vn.n1 vn.n0 0.0589632
R758 vn.n5 vn.n4 0.0392964
R759 vn.n7 vn.n6 0.0146
R760 vn.n3 vn.n2 0.00434178
R761 vn.n4 vn.n3 0.0034375
R762 trim_0.drain.n1 trim_0.drain.t2 41.0976
R763 trim_0.drain.n0 trim_0.drain.t0 17.4005
R764 trim_0.drain.n0 trim_0.drain.t1 17.4005
R765 trim_0.drain trim_0.drain.n0 7.1934
R766 trim_0.drain.n1 trim_0.drain 4.54309
R767 trim_0.drain trim_0.drain.n1 2.78583
R768 vp.n1 vp.t0 138.87
R769 vp vp.n7 1.64973
R770 vp.n5 vp.n1 0.751481
R771 vp.n6 vp.n5 0.512485
R772 vp.n1 vp.n0 0.0589631
R773 vp.n5 vp.n4 0.0390429
R774 vp.n7 vp.n6 0.0146
R775 vp.n3 vp.n2 0.00458983
R776 vp.n4 vp.n3 0.0034375
R777 trim_1.drain.n1 trim_1.drain.t2 41.1194
R778 trim_1.drain.n0 trim_1.drain.t0 17.4005
R779 trim_1.drain.n0 trim_1.drain.t1 17.4005
R780 trim_1.drain.n2 trim_1.drain.n0 7.1309
R781 trim_1.drain.n1 trim_1.drain 4.54309
R782 trim_1.drain.n2 trim_1.drain.n1 2.84833
R783 trim_1.drain trim_1.drain.n2 0.063
R784 trimb_2.n0 trimb_2.t1 135.6
R785 trimb_2.n0 trimb_2.t0 135.6
R786 trimb_2 trimb_2.n0 2.48064
R787 clk.n2 clk.t3 142.917
R788 clk.n0 clk.t2 142.911
R789 clk.n0 clk.t4 142.911
R790 clk.n2 clk.t0 142.905
R791 clk.n3 clk.t5 135.52
R792 clk.n1 clk.t1 135.52
R793 clk.n3 clk.n2 12.4888
R794 clk.n1 clk.n0 12.4715
R795 clk clk.n4 0.84425
R796 clk.n4 clk.n1 0.0793043
R797 clk.n4 clk.n3 0.0793043
R798 vdd.n5 vdd.t5 28.5655
R799 vdd.n5 vdd.t0 28.5655
R800 vdd.n0 vdd.t3 28.5655
R801 vdd.n0 vdd.t1 28.5655
R802 vdd.n18 vdd.t4 28.5655
R803 vdd.n18 vdd.t2 28.5655
R804 vdd.n1 vdd.n0 10.885
R805 vdd.n19 vdd.n18 10.3327
R806 vdd.n6 vdd.n5 9.04359
R807 vdd.n13 vdd.n12 4.91552
R808 vdd.n15 vdd.n14 1.13717
R809 vdd.n19 vdd.n17 0.580105
R810 vdd.n2 vdd.n1 0.567646
R811 vdd.n17 vdd.n16 0.555146
R812 vdd vdd.n19 0.0942085
R813 vdd.n6 vdd.n4 0.0565253
R814 vdd.n7 vdd.n6 0.0565253
R815 vdd.n11 vdd.n10 0.041625
R816 vdd.n3 vdd.n2 0.0364375
R817 vdd.n16 vdd.n15 0.0364375
R818 vdd.n12 vdd 0.024
R819 vdd.n9 vdd.n8 0.0140125
R820 vdd.n14 vdd.n13 0.0140125
R821 vdd.n4 vdd.n3 0.0083125
R822 vdd.n15 vdd.n7 0.0083125
R823 vdd.n10 vdd.n9 0.0034375
R824 vdd.n14 vdd.n11 0.0034375
R825 outp.n1 outp.t3 146.688
R826 outp.n1 outp.t4 138.821
R827 outp.n0 outp.t2 36.1754
R828 outp.n0 outp.t1 35.8981
R829 outp.n3 outp.t0 26.2669
R830 outp.n2 outp.n1 6.69396
R831 outp.n2 outp.n0 3.51216
R832 outp outp.n3 1.81295
R833 outp.n3 outp.n2 1.14368
R834 outn.n1 outn.t3 146.68
R835 outn.n1 outn.t4 138.822
R836 outn.n0 outn.t1 36.1794
R837 outn.n0 outn.t0 35.915
R838 outn.n3 outn.t2 26.2669
R839 outn.n2 outn.n1 6.69758
R840 outn.n2 outn.n0 3.51216
R841 outn outn.n3 1.81295
R842 outn.n3 outn.n2 1.14368
R843 trim_1 trim_1.t0 138.256
R844 trimb_1 trimb_1.t0 138.169
R845 trim_0 trim_0.t0 138.256
R846 trimb_0 trimb_0.t0 138.169
C0 trimb_1 trimb_0 0.934f
C1 trim_1.n2 trim_1.n4 0.551f
C2 outn clk 0.265f
C3 trim_1.drain w_4048_2972# 0.0387f
C4 trim_1.n2 trim_1.n1 0.0775f
C5 trim_1.drain clk 0.505f
C6 trim_1.n4 vdd 0.0293f
C7 vdd trim_1.n1 0.00179f
C8 trim_0.n3 vdd 0.0253f
C9 trim_0.drain vdd 0.263f
C10 a_3988_2912# vdd 0.252f
C11 outn trim_1.drain 0.0249f
C12 trim_0.n1 vdd 0.00179f
C13 trim_1.drain trim_1.n3 3.41f
C14 trim_0.n0 vdd 0.00143f
C15 trimb_3 trim_1.n4 6.08e-20
C16 w_3952_2876# vdd 0.0479f
C17 trimb_4 trim_1.n4 0.262f
C18 trim_0.n4 trim_0.n3 1.35f
C19 trim_0.drain comparator_core_0.diff 0.202f
C20 trim_0.n4 trim_0.drain 6.89f
C21 trimb_4 trim_1.n1 1.67e-19
C22 trim_0.n4 trim_0.n1 0.164f
C23 trimb_1 trim_1.n3 4.93e-20
C24 trim_1.n4 trimb_0 2.85e-20
C25 trim_1.n1 trimb_0 2.97e-19
C26 trim_0.n4 trim_0.n0 0.138f
C27 trim_1.n0 trim_1.n4 0.138f
C28 trim_0.n3 trim_0.n2 0.671f
C29 trim_1.n0 trim_1.n1 0.507f
C30 trim_0.n3 trim_0 4.93e-20
C31 trim_0.drain trim_0.n2 1.71f
C32 trim_0.n1 trim_0.n2 0.0775f
C33 trim_0.n1 trim_0 2.97e-19
C34 trim_4 trim_0.n3 4.9e-19
C35 vdd trim_2 0.12f
C36 trim_4 trim_0.drain 2.61e-20
C37 trim_0.n0 trim_0.n2 0.247f
C38 trim_4 trim_0.n1 1.67e-19
C39 trim_0.n0 trim_0 0.0508f
C40 trim_1.n4 clk 2.01e-19
C41 trim_0.drain w_4048_2972# 0.039f
C42 trim_0.n3 trim_1 4.93e-20
C43 trim_0.drain clk 0.527f
C44 trim_0.n3 trim_3 0.114f
C45 trim_0.drain trim_3 1.1e-19
C46 trim_0.n1 trim_1 0.0505f
C47 outn trim_1.n4 3.12e-21
C48 trim_1.n4 trim_1.n3 1.35f
C49 trim_0.n4 trim_2 1.61e-19
C50 trim_1.drain trim_1.n4 6.89f
C51 trim_1.n3 trim_1.n1 0.0769f
C52 outn trim_0.drain 0.24f
C53 trim_1.drain trim_1.n1 0.851f
C54 w_3952_2876# clk 0.0102f
C55 trim_1.n2 trimb_2 0.0413f
C56 trim_2 trim_0.n2 0.0413f
C57 vdd trimb_2 0.12f
C58 trim_0 trim_2 1.04f
C59 outn w_3952_2876# 0.00854f
C60 outp vdd 0.566f
C61 trim_1.drain w_3952_2876# 0.00574f
C62 trim_4 trim_2 0.00265f
C63 trim_1.n4 trimb_1 0.00218f
C64 trimb_1 trim_1.n1 0.0505f
C65 trim_1 trim_2 4.8e-19
C66 trimb_3 trimb_2 1.11f
C67 trim_3 trim_2 1.11f
C68 trimb_4 trimb_2 0.00265f
C69 outp comparator_core_0.diff 0.00669f
C70 trim_0.n4 outp 3.12e-21
C71 trim_1.n2 vdd 0.00772f
C72 trimb_0 trimb_2 1.04f
C73 trim_1.n0 trimb_2 1.67e-19
C74 trimb_3 trim_1.n2 7.7e-19
C75 trim_1.n4 trim_1.n1 0.164f
C76 trimb_4 trim_1.n2 0.00497f
C77 trim_0.n3 trim_0.drain 3.41f
C78 trimb_3 vdd 0.435f
C79 trim_0.n1 trim_0.n3 0.0769f
C80 comparator_core_0.diff vdd 0.0019f
C81 trim_0.n4 vdd 0.0293f
C82 trim_0.n1 trim_0.drain 0.851f
C83 trim_1.n2 trimb_0 0.00237f
C84 trimb_4 vdd 0.103f
C85 outp w_4048_2972# 0.32f
C86 trim_0.n3 trim_0.n0 0.077f
C87 outp clk 0.224f
C88 trim_0.drain trim_0.n0 0.851f
C89 vdd trimb_0 0.0784f
C90 trim_0.n1 trim_0.n0 0.507f
C91 trim_1.n0 trim_1.n2 0.247f
C92 trim_1.n3 trimb_2 2.66e-19
C93 w_3952_2876# trim_0.drain 0.00577f
C94 trim_1.drain trimb_2 2.61e-20
C95 outp outn 1.07f
C96 vdd trim_0.n2 0.00772f
C97 trim_1.n0 vdd 0.00143f
C98 trim_0 vdd 0.0784f
C99 outp trim_1.drain 0.24f
C100 trimb_3 trimb_4 0.00191f
C101 trim_4 vdd 0.103f
C102 trimb_3 trimb_0 3.33e-19
C103 vdd w_4048_2972# 0.74f
C104 trimb_4 trimb_0 0.0039f
C105 vdd clk 0.426f
C106 trim_1 vdd 0.0649f
C107 trimb_1 trimb_2 4.8e-19
C108 trim_0.n4 trim_0.n2 0.551f
C109 trim_3 vdd 0.435f
C110 trim_0.n3 trim_2 2.66e-19
C111 trim_0.n4 trim_0 2.85e-20
C112 trim_1.n2 trim_1.n3 0.671f
C113 trim_0.drain trim_2 2.61e-20
C114 trim_1.drain trim_1.n2 1.71f
C115 trim_0.n4 trim_4 0.262f
C116 outn vdd 0.573f
C117 vdd trim_1.n3 0.0253f
C118 trim_1.n0 trimb_0 0.0508f
C119 trim_1.drain vdd 0.262f
C120 trim_0.n0 trim_2 1.67e-19
C121 trim_0 trim_0.n2 0.00237f
C122 comparator_core_0.diff clk 0.0546f
C123 trim_0.n4 clk 2.01e-19
C124 trim_0.n4 trim_1 0.00218f
C125 trim_4 trim_0.n2 0.00497f
C126 trim_0.n4 trim_3 6.08e-20
C127 trim_4 trim_0 0.0039f
C128 trim_1.n2 trimb_1 0.00221f
C129 trimb_3 trim_1.n3 0.114f
C130 outn comparator_core_0.diff 0.00221f
C131 trim_1.drain trimb_3 1.1e-19
C132 trim_1.drain comparator_core_0.diff 0.202f
C133 vdd trimb_1 0.0649f
C134 trimb_4 trim_1.n3 4.9e-19
C135 trim_1.drain trimb_4 2.61e-20
C136 trim_1 trim_0.n2 0.00221f
C137 trim_3 trim_0.n2 7.7e-19
C138 trim_1 trim_0 0.934f
C139 trim_1.n4 trimb_2 1.61e-19
C140 trim_3 trim_0 3.33e-19
C141 trim_1.n3 trimb_0 4.93e-20
C142 trim_4 trim_1 0.592f
C143 trim_4 trim_3 0.00191f
C144 outp trim_0.drain 0.0249f
C145 trim_1.n0 trim_1.n3 0.077f
C146 trim_1.n0 trim_1.drain 0.851f
C147 trimb_3 trimb_1 3.33e-19
C148 w_4048_2972# clk 0.397f
C149 trimb_4 trimb_1 0.592f
C150 trim_1 trim_3 3.33e-19
C151 outn w_4048_2972# 0.328f
C152 outp w_3952_2876# 0.00774f
.ends

