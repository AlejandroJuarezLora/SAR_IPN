magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 866 542
<< pwell >>
rect 1 117 187 163
rect 1 -19 781 117
rect 84 -57 118 -19
<< scnmos >>
rect 79 7 109 137
rect 188 7 218 91
rect 284 7 314 91
rect 409 7 439 91
rect 505 7 535 91
rect 673 7 703 91
<< scpmoshvt >>
rect 79 257 109 457
rect 188 334 218 418
rect 291 334 321 418
rect 505 334 535 418
rect 577 334 607 418
rect 673 334 703 418
<< ndiff >>
rect 27 72 79 137
rect 27 38 35 72
rect 69 38 79 72
rect 27 7 79 38
rect 109 91 161 137
rect 109 53 188 91
rect 109 19 119 53
rect 153 19 188 53
rect 109 7 188 19
rect 218 7 284 91
rect 314 68 409 91
rect 314 34 326 68
rect 360 34 409 68
rect 314 7 409 34
rect 439 7 505 91
rect 535 68 673 91
rect 535 34 561 68
rect 595 34 629 68
rect 663 34 673 68
rect 535 7 673 34
rect 703 68 755 91
rect 703 34 713 68
rect 747 34 755 68
rect 703 7 755 34
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 377 79 411
rect 27 343 35 377
rect 69 343 79 377
rect 27 309 79 343
rect 27 275 35 309
rect 69 275 79 309
rect 27 257 79 275
rect 109 445 161 457
rect 109 411 119 445
rect 153 418 161 445
rect 153 411 188 418
rect 109 377 188 411
rect 109 343 119 377
rect 153 343 188 377
rect 109 334 188 343
rect 218 334 291 418
rect 321 385 505 418
rect 321 351 355 385
rect 389 351 430 385
rect 464 351 505 385
rect 321 334 505 351
rect 535 334 577 418
rect 607 385 673 418
rect 607 351 627 385
rect 661 351 673 385
rect 607 334 673 351
rect 703 385 759 418
rect 703 351 713 385
rect 747 351 759 385
rect 703 334 759 351
rect 109 309 161 334
rect 109 275 119 309
rect 153 275 161 309
rect 109 257 161 275
<< ndiffc >>
rect 35 38 69 72
rect 119 19 153 53
rect 326 34 360 68
rect 561 34 595 68
rect 629 34 663 68
rect 713 34 747 68
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 35 275 69 309
rect 119 411 153 445
rect 119 343 153 377
rect 355 351 389 385
rect 430 351 464 385
rect 627 351 661 385
rect 713 351 747 385
rect 119 275 153 309
<< poly >>
rect 79 457 109 483
rect 188 418 218 444
rect 291 418 321 444
rect 505 418 535 444
rect 577 418 607 444
rect 673 418 703 444
rect 79 225 109 257
rect 188 225 218 334
rect 291 319 321 334
rect 291 289 439 319
rect 505 302 535 334
rect 76 209 130 225
rect 76 175 86 209
rect 120 175 130 209
rect 76 159 130 175
rect 172 209 226 225
rect 172 175 182 209
rect 216 175 226 209
rect 409 189 439 289
rect 481 286 535 302
rect 481 252 491 286
rect 525 252 535 286
rect 481 236 535 252
rect 172 159 226 175
rect 284 173 367 189
rect 79 137 109 159
rect 188 91 218 159
rect 284 139 323 173
rect 357 139 367 173
rect 284 123 367 139
rect 409 173 463 189
rect 577 183 607 334
rect 673 302 703 334
rect 649 286 703 302
rect 649 252 659 286
rect 693 252 703 286
rect 649 236 703 252
rect 409 139 419 173
rect 453 139 463 173
rect 565 173 631 183
rect 565 159 581 173
rect 409 123 463 139
rect 505 139 581 159
rect 615 139 631 173
rect 505 129 631 139
rect 284 91 314 123
rect 409 91 439 123
rect 505 91 535 129
rect 673 91 703 236
rect 79 -19 109 7
rect 188 -19 218 7
rect 284 -19 314 7
rect 409 -19 439 7
rect 505 -19 535 7
rect 673 -19 703 7
<< polycont >>
rect 86 175 120 209
rect 182 175 216 209
rect 491 252 525 286
rect 323 139 357 173
rect 659 252 693 286
rect 419 139 453 173
rect 581 139 615 173
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 828 521
rect 18 445 85 453
rect 18 411 35 445
rect 69 411 85 445
rect 18 377 85 411
rect 18 343 35 377
rect 69 343 85 377
rect 18 309 85 343
rect 18 275 35 309
rect 69 275 85 309
rect 18 259 85 275
rect 119 445 153 487
rect 119 377 153 411
rect 119 309 153 343
rect 119 259 153 275
rect 187 419 593 453
rect 18 125 52 259
rect 187 225 221 419
rect 86 209 137 225
rect 120 175 137 209
rect 86 159 137 175
rect 182 209 221 225
rect 216 175 221 209
rect 182 159 221 175
rect 255 351 355 385
rect 389 351 430 385
rect 464 351 480 385
rect 103 125 137 159
rect 255 125 289 351
rect 18 72 69 125
rect 103 91 289 125
rect 323 286 525 317
rect 323 283 491 286
rect 323 173 357 283
rect 487 252 491 283
rect 323 123 357 139
rect 398 173 453 243
rect 398 139 419 173
rect 18 38 35 72
rect 254 84 289 91
rect 254 68 360 84
rect 18 11 69 38
rect 103 53 169 57
rect 103 19 119 53
rect 153 19 169 53
rect 103 -23 169 19
rect 254 34 326 68
rect 254 11 360 34
rect 398 11 453 139
rect 487 11 525 252
rect 559 286 593 419
rect 627 385 661 487
rect 627 335 661 351
rect 708 385 811 417
rect 708 351 713 385
rect 747 351 811 385
rect 708 335 811 351
rect 559 252 659 286
rect 693 252 709 286
rect 559 248 709 252
rect 743 173 811 335
rect 565 139 581 173
rect 615 139 811 173
rect 561 68 663 84
rect 595 34 629 68
rect 561 -23 663 34
rect 707 68 756 139
rect 707 34 713 68
rect 747 34 756 68
rect 707 18 756 34
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 828 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
<< metal1 >>
rect 0 521 828 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 828 521
rect 0 456 828 487
rect 0 -23 828 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 828 -23
rect 0 -88 828 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 mux2_1
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 74 487 108 521 0 FreeSans 250 0 0 0 VPB
port 5 nsew
flabel pwell s 84 -57 118 -23 0 FreeSans 250 0 0 0 VNB
port 6 nsew
flabel locali s 674 249 708 283 0 FreeSans 250 0 0 0 S
port 9 nsew
flabel locali s 582 249 616 283 0 FreeSans 250 0 0 0 S
port 9 nsew
flabel locali s 490 113 524 147 0 FreeSans 250 0 0 0 A1
port 8 nsew
flabel locali s 490 181 524 215 0 FreeSans 250 0 0 0 A1
port 8 nsew
flabel locali s 398 181 432 215 0 FreeSans 250 0 0 0 A0
port 10 nsew
flabel locali s 30 45 64 79 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 30 317 64 351 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 30 385 64 419 0 FreeSans 250 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 828 504
string path 0.000 -1.000 20.700 -1.000 
<< end >>
