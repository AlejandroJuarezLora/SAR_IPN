magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< pwell >>
rect -671 -365 1615 -279
rect -671 -847 -585 -365
rect 1529 -847 1615 -365
rect -671 -933 1615 -847
<< psubdiff >>
rect -645 -339 -481 -305
rect -447 -339 -413 -305
rect -379 -339 -345 -305
rect -311 -339 -277 -305
rect -243 -339 -209 -305
rect -175 -339 -141 -305
rect -107 -339 -73 -305
rect -39 -339 -5 -305
rect 29 -339 63 -305
rect 97 -339 131 -305
rect 165 -339 199 -305
rect 233 -339 267 -305
rect 301 -339 335 -305
rect 369 -339 403 -305
rect 437 -339 471 -305
rect 505 -339 539 -305
rect 573 -339 607 -305
rect 641 -339 675 -305
rect 709 -339 743 -305
rect 777 -339 811 -305
rect 845 -339 879 -305
rect 913 -339 947 -305
rect 981 -339 1015 -305
rect 1049 -339 1083 -305
rect 1117 -339 1151 -305
rect 1185 -339 1219 -305
rect 1253 -339 1287 -305
rect 1321 -339 1355 -305
rect 1389 -339 1589 -305
rect -645 -537 -611 -339
rect -645 -605 -611 -571
rect -645 -673 -611 -639
rect -645 -873 -611 -707
rect 1555 -537 1589 -339
rect 1555 -605 1589 -571
rect 1555 -673 1589 -639
rect 1555 -873 1589 -707
rect -645 -907 -413 -873
rect -379 -907 -345 -873
rect -311 -907 -277 -873
rect -243 -907 -209 -873
rect -175 -907 -141 -873
rect -107 -907 -73 -873
rect -39 -907 -5 -873
rect 29 -907 63 -873
rect 97 -907 131 -873
rect 165 -907 199 -873
rect 233 -907 267 -873
rect 301 -907 335 -873
rect 369 -907 403 -873
rect 437 -907 471 -873
rect 505 -907 539 -873
rect 573 -907 607 -873
rect 641 -907 675 -873
rect 709 -907 743 -873
rect 777 -907 811 -873
rect 845 -907 879 -873
rect 913 -907 947 -873
rect 981 -907 1015 -873
rect 1049 -907 1083 -873
rect 1117 -907 1151 -873
rect 1185 -907 1219 -873
rect 1253 -907 1287 -873
rect 1321 -907 1355 -873
rect 1389 -907 1589 -873
<< psubdiffcont >>
rect -481 -339 -447 -305
rect -413 -339 -379 -305
rect -345 -339 -311 -305
rect -277 -339 -243 -305
rect -209 -339 -175 -305
rect -141 -339 -107 -305
rect -73 -339 -39 -305
rect -5 -339 29 -305
rect 63 -339 97 -305
rect 131 -339 165 -305
rect 199 -339 233 -305
rect 267 -339 301 -305
rect 335 -339 369 -305
rect 403 -339 437 -305
rect 471 -339 505 -305
rect 539 -339 573 -305
rect 607 -339 641 -305
rect 675 -339 709 -305
rect 743 -339 777 -305
rect 811 -339 845 -305
rect 879 -339 913 -305
rect 947 -339 981 -305
rect 1015 -339 1049 -305
rect 1083 -339 1117 -305
rect 1151 -339 1185 -305
rect 1219 -339 1253 -305
rect 1287 -339 1321 -305
rect 1355 -339 1389 -305
rect -645 -571 -611 -537
rect -645 -639 -611 -605
rect -645 -707 -611 -673
rect 1555 -571 1589 -537
rect 1555 -639 1589 -605
rect 1555 -707 1589 -673
rect -413 -907 -379 -873
rect -345 -907 -311 -873
rect -277 -907 -243 -873
rect -209 -907 -175 -873
rect -141 -907 -107 -873
rect -73 -907 -39 -873
rect -5 -907 29 -873
rect 63 -907 97 -873
rect 131 -907 165 -873
rect 199 -907 233 -873
rect 267 -907 301 -873
rect 335 -907 369 -873
rect 403 -907 437 -873
rect 471 -907 505 -873
rect 539 -907 573 -873
rect 607 -907 641 -873
rect 675 -907 709 -873
rect 743 -907 777 -873
rect 811 -907 845 -873
rect 879 -907 913 -873
rect 947 -907 981 -873
rect 1015 -907 1049 -873
rect 1083 -907 1117 -873
rect 1151 -907 1185 -873
rect 1219 -907 1253 -873
rect 1287 -907 1321 -873
rect 1355 -907 1389 -873
<< locali >>
rect -645 -339 -481 -305
rect -447 -339 -413 -305
rect -379 -339 -345 -305
rect -311 -339 -277 -305
rect -243 -339 -209 -305
rect -175 -339 -141 -305
rect -107 -339 -73 -305
rect -39 -339 -5 -305
rect 29 -339 63 -305
rect 97 -339 131 -305
rect 165 -339 199 -305
rect 233 -339 267 -305
rect 301 -339 335 -305
rect 369 -339 403 -305
rect 437 -339 471 -305
rect 505 -339 539 -305
rect 573 -339 607 -305
rect 641 -339 675 -305
rect 709 -339 743 -305
rect 777 -339 811 -305
rect 845 -339 879 -305
rect 913 -339 947 -305
rect 981 -339 1015 -305
rect 1049 -339 1083 -305
rect 1117 -339 1151 -305
rect 1185 -339 1219 -305
rect 1253 -339 1287 -305
rect 1321 -339 1355 -305
rect 1389 -339 1589 -305
rect -645 -537 -611 -339
rect -645 -605 -611 -571
rect -645 -673 -611 -639
rect -645 -873 -611 -707
rect 1555 -537 1589 -339
rect 1555 -605 1589 -571
rect 1555 -673 1589 -639
rect 1555 -873 1589 -707
rect -645 -907 -413 -873
rect -379 -907 -345 -873
rect -311 -907 -277 -873
rect -243 -907 -209 -873
rect -175 -907 -141 -873
rect -107 -907 -73 -873
rect -39 -907 -5 -873
rect 29 -907 63 -873
rect 97 -907 131 -873
rect 165 -907 199 -873
rect 233 -907 267 -873
rect 301 -907 335 -873
rect 369 -907 403 -873
rect 437 -907 471 -873
rect 505 -907 539 -873
rect 573 -907 607 -873
rect 641 -907 675 -873
rect 709 -907 743 -873
rect 777 -907 811 -873
rect 845 -907 879 -873
rect 913 -907 947 -873
rect 981 -907 1015 -873
rect 1049 -907 1083 -873
rect 1117 -907 1151 -873
rect 1185 -907 1219 -873
rect 1253 -907 1287 -873
rect 1321 -907 1355 -873
rect 1389 -907 1589 -873
<< properties >>
string path -16.125 -8.050 39.300 -8.050 39.300 -22.250 -15.700 -22.250 -15.700 -8.050 
<< end >>
