magic
tech sky130B
magscale 1 2
timestamp 1695772279
<< nmoslvt >>
rect -30 -131 30 69
<< ndiff >>
rect -94 39 -30 69
rect -94 -101 -76 39
rect -42 -101 -30 39
rect -94 -131 -30 -101
rect 30 39 88 69
rect 30 -101 42 39
rect 76 -101 88 39
rect 30 -131 88 -101
<< ndiffc >>
rect -76 -101 -42 39
rect 42 -101 76 39
<< psubdiff >>
rect -166 39 -94 69
rect -166 -101 -150 39
rect -116 -101 -94 39
rect -166 -131 -94 -101
<< psubdiffcont >>
rect -150 -101 -116 39
<< poly >>
rect -33 141 33 157
rect -33 107 -17 141
rect 17 107 33 141
rect -33 91 33 107
rect -30 69 30 91
rect -30 -157 30 -131
<< polycont >>
rect -17 107 17 141
<< locali >>
rect -33 107 -17 141
rect 17 107 33 141
rect -160 57 -62 58
rect -160 39 -76 57
rect -160 -101 -150 39
rect -116 -101 -76 39
rect -160 -119 -76 -101
<< viali >>
rect -17 107 17 141
rect -76 39 -42 57
rect -76 -101 -42 39
rect -76 -119 -42 -101
rect 42 39 76 57
rect 42 -101 76 39
rect 42 -119 76 -101
<< metal1 >>
rect -38 141 40 150
rect -38 107 -17 141
rect 17 107 40 141
rect -38 98 40 107
rect -82 57 -36 69
rect -82 -119 -76 57
rect -42 -119 -36 57
rect -82 -131 -36 -119
rect 36 57 82 69
rect 36 -119 42 57
rect 76 -119 82 57
rect 36 -131 82 -119
<< labels >>
rlabel metal1 -82 -131 -36 -119 7 S
rlabel metal1 36 57 82 69 7 D
rlabel metal1 17 98 40 150 7 G
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 1 l 0.3 m 1 nf 1 diffcov 80 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
