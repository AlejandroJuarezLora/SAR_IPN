magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 498 542
<< pwell >>
rect 1 -19 459 163
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 109 137
rect 166 7 196 137
rect 267 7 297 137
rect 351 7 381 137
<< scpmoshvt >>
rect 79 257 109 457
rect 154 257 184 457
rect 277 257 307 457
rect 349 257 379 457
<< ndiff >>
rect 27 55 79 137
rect 27 21 35 55
rect 69 21 79 55
rect 27 7 79 21
rect 109 123 166 137
rect 109 89 119 123
rect 153 89 166 123
rect 109 7 166 89
rect 196 123 267 137
rect 196 89 219 123
rect 253 89 267 123
rect 196 55 267 89
rect 196 21 219 55
rect 253 21 267 55
rect 196 7 267 21
rect 297 49 351 137
rect 297 15 307 49
rect 341 15 351 49
rect 297 7 351 15
rect 381 123 433 137
rect 381 89 391 123
rect 425 89 433 123
rect 381 55 433 89
rect 381 21 391 55
rect 425 21 433 55
rect 381 7 433 21
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 257 79 411
rect 109 257 154 457
rect 184 437 277 457
rect 184 403 194 437
rect 228 403 277 437
rect 184 369 277 403
rect 184 335 194 369
rect 228 335 277 369
rect 184 257 277 335
rect 307 257 349 457
rect 379 441 433 457
rect 379 407 389 441
rect 423 407 433 441
rect 379 373 433 407
rect 379 339 389 373
rect 423 339 433 373
rect 379 305 433 339
rect 379 271 389 305
rect 423 271 433 305
rect 379 257 433 271
<< ndiffc >>
rect 35 21 69 55
rect 119 89 153 123
rect 219 89 253 123
rect 219 21 253 55
rect 307 15 341 49
rect 391 89 425 123
rect 391 21 425 55
<< pdiffc >>
rect 35 411 69 445
rect 194 403 228 437
rect 194 335 228 369
rect 389 407 423 441
rect 389 339 423 373
rect 389 271 423 305
<< poly >>
rect 79 457 109 483
rect 154 457 184 483
rect 277 457 307 483
rect 349 457 379 483
rect 79 225 109 257
rect 21 209 109 225
rect 21 175 31 209
rect 65 175 109 209
rect 21 159 109 175
rect 154 225 184 257
rect 277 225 307 257
rect 154 209 211 225
rect 154 175 167 209
rect 201 175 211 209
rect 154 159 211 175
rect 253 209 307 225
rect 253 175 263 209
rect 297 175 307 209
rect 253 159 307 175
rect 349 225 379 257
rect 349 209 415 225
rect 349 175 367 209
rect 401 175 415 209
rect 349 159 415 175
rect 79 137 109 159
rect 166 137 196 159
rect 267 137 297 159
rect 351 137 381 159
rect 79 -19 109 7
rect 166 -19 196 7
rect 267 -19 297 7
rect 351 -19 381 7
<< polycont >>
rect 31 175 65 209
rect 167 175 201 209
rect 263 175 297 209
rect 367 175 401 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 27 445 69 487
rect 27 411 35 445
rect 27 395 69 411
rect 167 437 267 453
rect 379 441 443 487
rect 167 403 194 437
rect 228 403 267 437
rect 167 369 267 403
rect 17 209 65 358
rect 17 175 31 209
rect 17 93 65 175
rect 99 335 194 369
rect 228 335 267 369
rect 99 327 267 335
rect 99 125 133 327
rect 167 243 247 293
rect 305 283 345 441
rect 281 249 345 283
rect 379 407 389 441
rect 423 407 443 441
rect 379 373 443 407
rect 379 339 389 373
rect 423 339 443 373
rect 379 305 443 339
rect 379 271 389 305
rect 423 271 443 305
rect 379 251 443 271
rect 167 209 201 243
rect 281 209 317 249
rect 244 175 263 209
rect 297 175 317 209
rect 351 209 443 215
rect 351 175 367 209
rect 401 175 443 209
rect 167 159 201 175
rect 237 125 443 133
rect 99 123 169 125
rect 99 89 119 123
rect 153 89 169 123
rect 203 123 443 125
rect 203 89 219 123
rect 253 99 391 123
rect 253 89 269 99
rect 203 55 269 89
rect 375 89 391 99
rect 425 89 443 123
rect 17 21 35 55
rect 69 21 219 55
rect 253 21 269 55
rect 17 19 269 21
rect 307 49 341 65
rect 375 55 443 89
rect 375 21 391 55
rect 425 21 443 55
rect 375 16 443 21
rect 307 -23 341 15
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
<< metal1 >>
rect 0 521 460 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 0 456 460 487
rect 0 -23 460 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
rect 0 -88 460 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 o22ai_1
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 305 317 339 351 0 FreeSans 400 0 0 0 A2
port 8 nsew
flabel locali s 29 113 63 147 0 FreeSans 400 0 0 0 B1
port 9 nsew
flabel locali s 213 385 247 419 0 FreeSans 400 0 0 0 Y
port 11 nsew
flabel locali s 397 181 431 215 0 FreeSans 400 0 0 0 A1
port 7 nsew
flabel locali s 213 249 247 283 0 FreeSans 400 0 0 0 B2
port 10 nsew
<< properties >>
string FIXED_BBOX 0 -40 460 504
string path 0.000 -1.000 11.500 -1.000 
<< end >>
