magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 1970 542
<< pwell >>
rect 1 -19 1907 163
rect 30 -57 64 -19
<< scnmos >>
rect 83 7 113 137
rect 167 7 197 137
rect 251 7 281 137
rect 335 7 365 137
rect 523 7 553 137
rect 607 7 637 137
rect 691 7 721 137
rect 775 7 805 137
rect 859 7 889 137
rect 943 7 973 137
rect 1027 7 1057 137
rect 1111 7 1141 137
rect 1211 7 1241 137
rect 1295 7 1325 137
rect 1379 7 1409 137
rect 1463 7 1493 137
rect 1547 7 1577 137
rect 1631 7 1661 137
rect 1715 7 1745 137
rect 1799 7 1829 137
<< scpmoshvt >>
rect 83 257 113 457
rect 167 257 197 457
rect 251 257 281 457
rect 335 257 365 457
rect 523 257 553 457
rect 607 257 637 457
rect 691 257 721 457
rect 775 257 805 457
rect 859 257 889 457
rect 943 257 973 457
rect 1027 257 1057 457
rect 1111 257 1141 457
rect 1211 257 1241 457
rect 1295 257 1325 457
rect 1379 257 1409 457
rect 1463 257 1493 457
rect 1547 257 1577 457
rect 1631 257 1661 457
rect 1715 257 1745 457
rect 1799 257 1829 457
<< ndiff >>
rect 27 123 83 137
rect 27 89 39 123
rect 73 89 83 123
rect 27 55 83 89
rect 27 21 39 55
rect 73 21 83 55
rect 27 7 83 21
rect 113 123 167 137
rect 113 89 123 123
rect 157 89 167 123
rect 113 7 167 89
rect 197 55 251 137
rect 197 21 207 55
rect 241 21 251 55
rect 197 7 251 21
rect 281 123 335 137
rect 281 89 291 123
rect 325 89 335 123
rect 281 7 335 89
rect 365 55 417 137
rect 365 21 375 55
rect 409 21 417 55
rect 365 7 417 21
rect 471 123 523 137
rect 471 89 479 123
rect 513 89 523 123
rect 471 7 523 89
rect 553 55 607 137
rect 553 21 563 55
rect 597 21 607 55
rect 553 7 607 21
rect 637 123 691 137
rect 637 89 647 123
rect 681 89 691 123
rect 637 7 691 89
rect 721 55 775 137
rect 721 21 731 55
rect 765 21 775 55
rect 721 7 775 21
rect 805 123 859 137
rect 805 89 815 123
rect 849 89 859 123
rect 805 7 859 89
rect 889 55 943 137
rect 889 21 899 55
rect 933 21 943 55
rect 889 7 943 21
rect 973 123 1027 137
rect 973 89 983 123
rect 1017 89 1027 123
rect 973 7 1027 89
rect 1057 55 1111 137
rect 1057 21 1067 55
rect 1101 21 1111 55
rect 1057 7 1111 21
rect 1141 123 1211 137
rect 1141 89 1167 123
rect 1201 89 1211 123
rect 1141 55 1211 89
rect 1141 21 1167 55
rect 1201 21 1211 55
rect 1141 7 1211 21
rect 1241 55 1295 137
rect 1241 21 1251 55
rect 1285 21 1295 55
rect 1241 7 1295 21
rect 1325 123 1379 137
rect 1325 89 1335 123
rect 1369 89 1379 123
rect 1325 55 1379 89
rect 1325 21 1335 55
rect 1369 21 1379 55
rect 1325 7 1379 21
rect 1409 55 1463 137
rect 1409 21 1419 55
rect 1453 21 1463 55
rect 1409 7 1463 21
rect 1493 123 1547 137
rect 1493 89 1503 123
rect 1537 89 1547 123
rect 1493 55 1547 89
rect 1493 21 1503 55
rect 1537 21 1547 55
rect 1493 7 1547 21
rect 1577 55 1631 137
rect 1577 21 1587 55
rect 1621 21 1631 55
rect 1577 7 1631 21
rect 1661 123 1715 137
rect 1661 89 1671 123
rect 1705 89 1715 123
rect 1661 55 1715 89
rect 1661 21 1671 55
rect 1705 21 1715 55
rect 1661 7 1715 21
rect 1745 55 1799 137
rect 1745 21 1755 55
rect 1789 21 1799 55
rect 1745 7 1799 21
rect 1829 123 1881 137
rect 1829 89 1839 123
rect 1873 89 1881 123
rect 1829 55 1881 89
rect 1829 21 1839 55
rect 1873 21 1881 55
rect 1829 7 1881 21
<< pdiff >>
rect 27 443 83 457
rect 27 409 39 443
rect 73 409 83 443
rect 27 375 83 409
rect 27 341 39 375
rect 73 341 83 375
rect 27 307 83 341
rect 27 273 39 307
rect 73 273 83 307
rect 27 257 83 273
rect 113 437 167 457
rect 113 403 123 437
rect 157 403 167 437
rect 113 369 167 403
rect 113 335 123 369
rect 157 335 167 369
rect 113 301 167 335
rect 113 267 123 301
rect 157 267 167 301
rect 113 257 167 267
rect 197 443 251 457
rect 197 409 207 443
rect 241 409 251 443
rect 197 375 251 409
rect 197 341 207 375
rect 241 341 251 375
rect 197 257 251 341
rect 281 437 335 457
rect 281 403 291 437
rect 325 403 335 437
rect 281 369 335 403
rect 281 335 291 369
rect 325 335 335 369
rect 281 301 335 335
rect 281 267 291 301
rect 325 267 335 301
rect 281 257 335 267
rect 365 437 523 457
rect 365 403 375 437
rect 409 403 479 437
rect 513 403 523 437
rect 365 257 523 403
rect 553 437 607 457
rect 553 403 563 437
rect 597 403 607 437
rect 553 369 607 403
rect 553 335 563 369
rect 597 335 607 369
rect 553 257 607 335
rect 637 437 691 457
rect 637 403 647 437
rect 681 403 691 437
rect 637 257 691 403
rect 721 437 775 457
rect 721 403 731 437
rect 765 403 775 437
rect 721 369 775 403
rect 721 335 731 369
rect 765 335 775 369
rect 721 257 775 335
rect 805 369 859 457
rect 805 335 815 369
rect 849 335 859 369
rect 805 257 859 335
rect 889 447 943 457
rect 889 413 899 447
rect 933 413 943 447
rect 889 257 943 413
rect 973 369 1027 457
rect 973 335 983 369
rect 1017 335 1027 369
rect 973 257 1027 335
rect 1057 447 1111 457
rect 1057 413 1067 447
rect 1101 413 1111 447
rect 1057 257 1111 413
rect 1141 447 1211 457
rect 1141 413 1159 447
rect 1193 413 1211 447
rect 1141 257 1211 413
rect 1241 447 1295 457
rect 1241 413 1251 447
rect 1285 413 1295 447
rect 1241 257 1295 413
rect 1325 369 1379 457
rect 1325 335 1335 369
rect 1369 335 1379 369
rect 1325 257 1379 335
rect 1409 437 1463 457
rect 1409 403 1419 437
rect 1453 403 1463 437
rect 1409 257 1463 403
rect 1493 369 1547 457
rect 1493 335 1503 369
rect 1537 335 1547 369
rect 1493 257 1547 335
rect 1577 437 1631 457
rect 1577 403 1587 437
rect 1621 403 1631 437
rect 1577 369 1631 403
rect 1577 335 1587 369
rect 1621 335 1631 369
rect 1577 257 1631 335
rect 1661 437 1715 457
rect 1661 403 1671 437
rect 1705 403 1715 437
rect 1661 257 1715 403
rect 1745 437 1799 457
rect 1745 403 1755 437
rect 1789 403 1799 437
rect 1745 369 1799 403
rect 1745 335 1755 369
rect 1789 335 1799 369
rect 1745 301 1799 335
rect 1745 267 1755 301
rect 1789 267 1799 301
rect 1745 257 1799 267
rect 1829 437 1888 457
rect 1829 403 1839 437
rect 1873 403 1888 437
rect 1829 369 1888 403
rect 1829 335 1839 369
rect 1873 335 1888 369
rect 1829 301 1888 335
rect 1829 267 1839 301
rect 1873 267 1888 301
rect 1829 257 1888 267
<< ndiffc >>
rect 39 89 73 123
rect 39 21 73 55
rect 123 89 157 123
rect 207 21 241 55
rect 291 89 325 123
rect 375 21 409 55
rect 479 89 513 123
rect 563 21 597 55
rect 647 89 681 123
rect 731 21 765 55
rect 815 89 849 123
rect 899 21 933 55
rect 983 89 1017 123
rect 1067 21 1101 55
rect 1167 89 1201 123
rect 1167 21 1201 55
rect 1251 21 1285 55
rect 1335 89 1369 123
rect 1335 21 1369 55
rect 1419 21 1453 55
rect 1503 89 1537 123
rect 1503 21 1537 55
rect 1587 21 1621 55
rect 1671 89 1705 123
rect 1671 21 1705 55
rect 1755 21 1789 55
rect 1839 89 1873 123
rect 1839 21 1873 55
<< pdiffc >>
rect 39 409 73 443
rect 39 341 73 375
rect 39 273 73 307
rect 123 403 157 437
rect 123 335 157 369
rect 123 267 157 301
rect 207 409 241 443
rect 207 341 241 375
rect 291 403 325 437
rect 291 335 325 369
rect 291 267 325 301
rect 375 403 409 437
rect 479 403 513 437
rect 563 403 597 437
rect 563 335 597 369
rect 647 403 681 437
rect 731 403 765 437
rect 731 335 765 369
rect 815 335 849 369
rect 899 413 933 447
rect 983 335 1017 369
rect 1067 413 1101 447
rect 1159 413 1193 447
rect 1251 413 1285 447
rect 1335 335 1369 369
rect 1419 403 1453 437
rect 1503 335 1537 369
rect 1587 403 1621 437
rect 1587 335 1621 369
rect 1671 403 1705 437
rect 1755 403 1789 437
rect 1755 335 1789 369
rect 1755 267 1789 301
rect 1839 403 1873 437
rect 1839 335 1873 369
rect 1839 267 1873 301
<< poly >>
rect 83 457 113 483
rect 167 457 197 483
rect 251 457 281 483
rect 335 457 365 483
rect 523 457 553 483
rect 607 457 637 483
rect 691 457 721 483
rect 775 457 805 483
rect 859 457 889 483
rect 943 457 973 483
rect 1027 457 1057 483
rect 1111 457 1141 483
rect 1211 457 1241 483
rect 1295 457 1325 483
rect 1379 457 1409 483
rect 1463 457 1493 483
rect 1547 457 1577 483
rect 1631 457 1661 483
rect 1715 457 1745 483
rect 1799 457 1829 483
rect 83 225 113 257
rect 167 225 197 257
rect 251 225 281 257
rect 335 225 365 257
rect 523 225 553 257
rect 607 225 637 257
rect 691 225 721 257
rect 65 209 365 225
rect 65 175 81 209
rect 115 175 149 209
rect 183 175 217 209
rect 251 175 285 209
rect 319 175 365 209
rect 65 159 365 175
rect 514 209 721 225
rect 514 175 530 209
rect 564 175 598 209
rect 632 175 666 209
rect 700 175 721 209
rect 514 159 721 175
rect 83 137 113 159
rect 167 137 197 159
rect 251 137 281 159
rect 335 137 365 159
rect 523 137 553 159
rect 607 137 637 159
rect 691 137 721 159
rect 775 225 805 257
rect 859 225 889 257
rect 943 225 973 257
rect 1027 225 1057 257
rect 1111 225 1141 257
rect 1211 225 1241 257
rect 1295 225 1325 257
rect 1379 225 1409 257
rect 1463 225 1493 257
rect 1547 225 1577 257
rect 775 209 1057 225
rect 775 175 945 209
rect 979 175 1013 209
rect 1047 175 1057 209
rect 775 159 1057 175
rect 1099 209 1153 225
rect 1099 175 1109 209
rect 1143 175 1153 209
rect 1099 159 1153 175
rect 1199 209 1253 225
rect 1199 175 1209 209
rect 1243 175 1253 209
rect 1199 159 1253 175
rect 1295 209 1577 225
rect 1295 175 1311 209
rect 1345 175 1379 209
rect 1413 175 1447 209
rect 1481 175 1515 209
rect 1549 175 1577 209
rect 1295 159 1577 175
rect 775 137 805 159
rect 859 137 889 159
rect 943 137 973 159
rect 1027 137 1057 159
rect 1111 137 1141 159
rect 1211 137 1241 159
rect 1295 137 1325 159
rect 1379 137 1409 159
rect 1463 137 1493 159
rect 1547 137 1577 159
rect 1631 225 1661 257
rect 1715 225 1745 257
rect 1799 225 1829 257
rect 1631 209 1838 225
rect 1631 175 1647 209
rect 1681 175 1715 209
rect 1749 175 1783 209
rect 1817 175 1838 209
rect 1631 159 1838 175
rect 1631 137 1661 159
rect 1715 137 1745 159
rect 1799 137 1829 159
rect 83 -19 113 7
rect 167 -19 197 7
rect 251 -19 281 7
rect 335 -19 365 7
rect 523 -19 553 7
rect 607 -19 637 7
rect 691 -19 721 7
rect 775 -19 805 7
rect 859 -19 889 7
rect 943 -19 973 7
rect 1027 -19 1057 7
rect 1111 -19 1141 7
rect 1211 -19 1241 7
rect 1295 -19 1325 7
rect 1379 -19 1409 7
rect 1463 -19 1493 7
rect 1547 -19 1577 7
rect 1631 -19 1661 7
rect 1715 -19 1745 7
rect 1799 -19 1829 7
<< polycont >>
rect 81 175 115 209
rect 149 175 183 209
rect 217 175 251 209
rect 285 175 319 209
rect 530 175 564 209
rect 598 175 632 209
rect 666 175 700 209
rect 945 175 979 209
rect 1013 175 1047 209
rect 1109 175 1143 209
rect 1209 175 1243 209
rect 1311 175 1345 209
rect 1379 175 1413 209
rect 1447 175 1481 209
rect 1515 175 1549 209
rect 1647 175 1681 209
rect 1715 175 1749 209
rect 1783 175 1817 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1133 521
rect 1167 487 1225 521
rect 1259 487 1317 521
rect 1351 487 1409 521
rect 1443 487 1501 521
rect 1535 487 1593 521
rect 1627 487 1685 521
rect 1719 487 1777 521
rect 1811 487 1869 521
rect 1903 487 1932 521
rect 31 443 81 487
rect 31 409 39 443
rect 73 409 81 443
rect 31 375 81 409
rect 31 341 39 375
rect 73 341 81 375
rect 31 307 81 341
rect 31 273 39 307
rect 73 273 81 307
rect 31 257 81 273
rect 115 437 165 453
rect 115 403 123 437
rect 157 403 165 437
rect 115 369 165 403
rect 115 335 123 369
rect 157 335 165 369
rect 115 301 165 335
rect 199 443 249 487
rect 199 409 207 443
rect 241 409 249 443
rect 199 375 249 409
rect 199 341 207 375
rect 241 341 249 375
rect 199 325 249 341
rect 283 437 333 453
rect 283 403 291 437
rect 325 403 333 437
rect 283 369 333 403
rect 367 437 521 487
rect 367 403 375 437
rect 409 403 479 437
rect 513 403 521 437
rect 367 385 521 403
rect 555 437 605 453
rect 555 403 563 437
rect 597 403 605 437
rect 283 335 291 369
rect 325 351 333 369
rect 555 369 605 403
rect 639 437 689 487
rect 639 403 647 437
rect 681 403 689 437
rect 639 385 689 403
rect 723 447 1117 453
rect 723 437 899 447
rect 723 403 731 437
rect 765 419 899 437
rect 325 335 425 351
rect 115 267 123 301
rect 157 283 165 301
rect 283 301 425 335
rect 555 335 563 369
rect 597 351 605 369
rect 723 369 765 403
rect 891 413 899 419
rect 933 419 1067 447
rect 933 413 941 419
rect 891 395 941 413
rect 1051 413 1067 419
rect 1101 413 1117 447
rect 1051 395 1117 413
rect 1151 447 1201 487
rect 1151 413 1159 447
rect 1193 413 1201 447
rect 1151 395 1201 413
rect 1235 447 1629 453
rect 1235 413 1251 447
rect 1285 437 1629 447
rect 1285 419 1419 437
rect 1285 413 1301 419
rect 1235 395 1301 413
rect 1411 403 1419 419
rect 1453 419 1587 437
rect 1453 403 1461 419
rect 1411 385 1461 403
rect 1579 403 1587 419
rect 1621 403 1629 437
rect 723 351 731 369
rect 597 335 731 351
rect 555 317 765 335
rect 799 369 857 385
rect 799 335 815 369
rect 849 361 857 369
rect 975 369 1017 385
rect 975 361 983 369
rect 849 335 983 361
rect 1335 369 1377 385
rect 1017 335 1335 361
rect 1369 351 1377 369
rect 1495 369 1545 385
rect 1495 351 1503 369
rect 1369 335 1503 351
rect 1537 335 1545 369
rect 799 327 1545 335
rect 283 283 291 301
rect 157 267 291 283
rect 325 283 425 301
rect 799 283 833 327
rect 1193 317 1545 327
rect 1579 369 1629 403
rect 1663 437 1713 487
rect 1663 403 1671 437
rect 1705 403 1713 437
rect 1663 385 1713 403
rect 1747 437 1797 453
rect 1747 403 1755 437
rect 1789 403 1797 437
rect 1579 335 1587 369
rect 1621 351 1629 369
rect 1747 369 1797 403
rect 1747 351 1755 369
rect 1621 335 1755 351
rect 1789 335 1797 369
rect 1579 317 1797 335
rect 1747 301 1797 317
rect 325 267 833 283
rect 115 249 833 267
rect 867 259 1159 293
rect 18 209 350 215
rect 18 175 81 209
rect 115 175 149 209
rect 183 175 217 209
rect 251 175 285 209
rect 319 175 350 209
rect 23 123 73 139
rect 384 133 425 249
rect 867 215 901 259
rect 472 209 901 215
rect 472 175 530 209
rect 564 175 598 209
rect 632 175 666 209
rect 700 175 901 209
rect 935 209 1057 225
rect 935 175 945 209
rect 979 175 1013 209
rect 1047 175 1057 209
rect 1093 209 1159 259
rect 1093 175 1109 209
rect 1143 175 1159 209
rect 1193 249 1684 283
rect 1747 267 1755 301
rect 1789 267 1797 301
rect 1747 249 1797 267
rect 1831 437 1881 487
rect 1831 403 1839 437
rect 1873 403 1881 437
rect 1831 369 1881 403
rect 1831 335 1839 369
rect 1873 335 1881 369
rect 1831 301 1881 335
rect 1831 267 1839 301
rect 1873 267 1881 301
rect 1831 249 1881 267
rect 1193 209 1259 249
rect 1631 215 1684 249
rect 1193 175 1209 209
rect 1243 175 1259 209
rect 1295 209 1577 215
rect 1295 175 1311 209
rect 1345 175 1379 209
rect 1413 175 1447 209
rect 1481 175 1515 209
rect 1549 175 1577 209
rect 1631 209 1915 215
rect 1631 175 1647 209
rect 1681 175 1715 209
rect 1749 175 1783 209
rect 1817 175 1915 209
rect 935 159 1057 175
rect 23 89 39 123
rect 107 123 425 133
rect 1093 124 1889 141
rect 107 89 123 123
rect 157 89 291 123
rect 325 89 425 123
rect 463 123 1889 124
rect 463 89 479 123
rect 513 89 647 123
rect 681 89 815 123
rect 849 89 983 123
rect 1017 89 1167 123
rect 1201 107 1335 123
rect 1201 89 1217 107
rect 23 55 73 89
rect 1151 55 1217 89
rect 1319 89 1335 107
rect 1369 105 1503 123
rect 1369 89 1385 105
rect 23 21 39 55
rect 73 21 207 55
rect 241 21 375 55
rect 409 21 563 55
rect 597 21 731 55
rect 765 21 899 55
rect 933 21 1067 55
rect 1101 21 1117 55
rect 23 11 1117 21
rect 1151 21 1167 55
rect 1201 21 1217 55
rect 1151 11 1217 21
rect 1251 55 1285 71
rect 1251 -23 1285 21
rect 1319 55 1385 89
rect 1487 89 1503 105
rect 1537 107 1671 123
rect 1537 89 1553 107
rect 1319 21 1335 55
rect 1369 21 1385 55
rect 1319 11 1385 21
rect 1419 55 1453 71
rect 1419 -23 1453 21
rect 1487 55 1553 89
rect 1655 89 1671 107
rect 1705 105 1839 123
rect 1705 89 1721 105
rect 1487 21 1503 55
rect 1537 21 1553 55
rect 1487 11 1553 21
rect 1587 55 1621 71
rect 1587 -23 1621 21
rect 1655 55 1721 89
rect 1823 89 1839 105
rect 1873 89 1889 123
rect 1655 21 1671 55
rect 1705 21 1721 55
rect 1655 11 1721 21
rect 1755 55 1789 71
rect 1755 -23 1789 21
rect 1823 55 1889 89
rect 1823 21 1839 55
rect 1873 21 1889 55
rect 1823 11 1889 21
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1133 -23
rect 1167 -57 1225 -23
rect 1259 -57 1317 -23
rect 1351 -57 1409 -23
rect 1443 -57 1501 -23
rect 1535 -57 1593 -23
rect 1627 -57 1685 -23
rect 1719 -57 1777 -23
rect 1811 -57 1869 -23
rect 1903 -57 1932 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 857 487 891 521
rect 949 487 983 521
rect 1041 487 1075 521
rect 1133 487 1167 521
rect 1225 487 1259 521
rect 1317 487 1351 521
rect 1409 487 1443 521
rect 1501 487 1535 521
rect 1593 487 1627 521
rect 1685 487 1719 521
rect 1777 487 1811 521
rect 1869 487 1903 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
rect 857 -57 891 -23
rect 949 -57 983 -23
rect 1041 -57 1075 -23
rect 1133 -57 1167 -23
rect 1225 -57 1259 -23
rect 1317 -57 1351 -23
rect 1409 -57 1443 -23
rect 1501 -57 1535 -23
rect 1593 -57 1627 -23
rect 1685 -57 1719 -23
rect 1777 -57 1811 -23
rect 1869 -57 1903 -23
<< metal1 >>
rect 0 521 1932 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1133 521
rect 1167 487 1225 521
rect 1259 487 1317 521
rect 1351 487 1409 521
rect 1443 487 1501 521
rect 1535 487 1593 521
rect 1627 487 1685 521
rect 1719 487 1777 521
rect 1811 487 1869 521
rect 1903 487 1932 521
rect 0 456 1932 487
rect 0 -23 1932 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1133 -23
rect 1167 -57 1225 -23
rect 1259 -57 1317 -23
rect 1351 -57 1409 -23
rect 1443 -57 1501 -23
rect 1535 -57 1593 -23
rect 1627 -57 1685 -23
rect 1719 -57 1777 -23
rect 1811 -57 1869 -23
rect 1903 -57 1932 -23
rect 0 -88 1932 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 o221ai_4
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 586 181 620 215 0 FreeSans 400 0 0 0 B1
port 11 nsew
flabel locali s 954 181 988 215 0 FreeSans 400 0 0 0 B2
port 7 nsew
flabel locali s 1414 181 1448 215 0 FreeSans 400 180 0 0 A2
port 9 nsew
flabel locali s 214 181 248 215 0 FreeSans 400 0 0 0 C1
port 12 nsew
flabel locali s 1230 317 1264 351 0 FreeSans 400 180 0 0 Y
port 8 nsew
flabel locali s 1690 181 1724 215 0 FreeSans 400 180 0 0 A1
port 10 nsew
<< properties >>
string FIXED_BBOX 0 -40 1932 504
string path 0.000 -1.000 48.300 -1.000 
<< end >>
