magic
tech sky130B
magscale 1 2
timestamp 1696279433
<< nwell >>
rect 1946 1054 2036 1114
<< locali >>
rect 1638 345 1672 453
rect 1638 338 2375 345
rect 3021 338 3055 444
rect 1638 311 3055 338
rect 2341 304 3055 311
rect 2341 -17 2375 304
rect 2085 -51 2599 -17
rect 2341 -529 2375 -51
rect 2316 -532 2375 -529
rect 2308 -681 2410 -532
rect 2287 -715 2435 -681
rect 2345 -910 2379 -715
<< viali >>
rect 2345 -944 2379 -910
<< metal1 >>
rect -443 1552 -375 1625
rect -431 1116 -387 1552
rect 1416 1518 1444 1560
rect 3223 1518 3252 1555
rect 1398 1466 1404 1518
rect 1456 1466 1462 1518
rect 250 1405 278 1406
rect 2286 1405 2314 1501
rect 3204 1466 3210 1518
rect 3262 1466 3268 1518
rect 250 1377 4445 1405
rect 250 1141 278 1377
rect -435 1110 -383 1116
rect -435 1052 -383 1058
rect 55 1114 115 1120
rect 430 1106 458 1377
rect 1068 1124 1096 1377
rect 874 1114 934 1120
rect 55 1048 115 1054
rect 1251 1087 1279 1377
rect 1620 1104 1648 1377
rect 1835 1121 1863 1377
rect 1963 1090 2023 1120
rect 2846 1113 2874 1377
rect 2436 1090 2464 1094
rect 874 1048 934 1054
rect 1963 1062 2177 1090
rect 1963 1048 2023 1062
rect 244 730 272 1031
rect 1063 844 1091 1025
rect 1404 856 1456 862
rect 1063 816 1404 844
rect 1796 849 1824 1028
rect 1913 849 1919 861
rect 1796 844 1919 849
rect 1456 821 1919 844
rect 1456 816 1824 821
rect 1404 798 1456 804
rect 1796 552 1824 816
rect 1913 809 1919 821
rect 1971 809 1977 861
rect 2149 785 2177 1062
rect 2436 1062 2706 1090
rect 2436 867 2464 1062
rect 2664 1048 2720 1054
rect 3039 1052 3067 1377
rect 3408 1057 3436 1377
rect 3602 1116 3630 1377
rect 3747 1114 3807 1120
rect 4226 1063 4254 1377
rect 4417 1125 4445 1377
rect 4576 1114 4636 1120
rect 3747 1048 3807 1054
rect 4576 1048 4636 1054
rect 2420 861 2472 867
rect 2420 803 2472 809
rect 2882 813 2910 1028
rect 3210 939 3262 945
rect 3210 881 3262 887
rect 3222 813 3250 881
rect 3601 813 3629 1018
rect 2131 733 2137 785
rect 2189 733 2195 785
rect 2149 502 2177 733
rect 2002 474 2177 502
rect 2436 515 2464 803
rect 2882 791 3629 813
rect 2870 785 3629 791
rect 2870 727 2922 733
rect 2882 552 2910 727
rect 4423 712 4451 1027
rect 2436 487 2692 515
rect 2436 478 2464 487
rect 1840 264 1869 448
rect 1502 235 1869 264
rect 1840 49 1869 235
rect 2810 250 2839 446
rect 2810 221 3289 250
rect 2810 47 2839 221
rect 1738 -3715 1768 -12
rect 1896 -220 1926 -74
rect 2719 -220 2749 -73
rect 1896 -250 2749 -220
rect 2169 -333 2199 -250
rect 2169 -363 2563 -333
rect 2169 -579 2199 -363
rect 2533 -581 2563 -363
rect 2742 -588 2802 -582
rect 1922 -594 1982 -588
rect 2742 -654 2754 -648
rect 2784 -654 2802 -648
rect 1922 -660 1982 -654
rect 2141 -912 2171 -667
rect 2339 -910 2385 -898
rect 2339 -912 2345 -910
rect 2141 -942 2345 -912
rect 1727 -3721 1779 -3715
rect 1727 -3779 1779 -3773
rect 1738 -3926 1768 -3925
rect 2144 -3926 2174 -942
rect 2339 -944 2345 -942
rect 2379 -912 2385 -910
rect 2585 -912 2615 -679
rect 2379 -942 2618 -912
rect 2379 -944 2385 -942
rect 2339 -956 2385 -944
rect 2922 -1037 2952 -10
rect 2755 -1067 2952 -1037
rect 2755 -3586 2785 -1067
rect 2743 -3592 2795 -3586
rect 2743 -3650 2795 -3644
rect 2754 -3926 2784 -3925
rect 252 -3947 284 -3936
rect 25 -3975 59 -3947
rect 87 -3975 121 -3947
rect 162 -3975 196 -3947
rect 251 -3975 285 -3947
rect 395 -3974 429 -3946
rect 524 -3956 4281 -3926
rect 1721 -4069 1727 -4017
rect 1779 -4069 1785 -4017
rect 2140 -4059 2170 -3956
rect 4364 -3990 4398 -3962
rect 4506 -3985 4540 -3957
rect 4596 -3985 4630 -3957
rect 4671 -3985 4705 -3957
rect 4733 -3985 4767 -3957
rect 2737 -4071 2743 -4019
rect 2795 -4071 2801 -4019
<< via1 >>
rect 1404 1466 1456 1518
rect 3210 1466 3262 1518
rect -435 1058 -383 1110
rect 55 1054 115 1114
rect 874 1054 934 1114
rect 1404 804 1456 856
rect 1919 809 1971 861
rect 3747 1054 3807 1114
rect 4576 1054 4636 1114
rect 2420 809 2472 861
rect 3210 887 3262 939
rect 2137 733 2189 785
rect 2870 733 2922 785
rect 1922 -654 1982 -594
rect 2742 -648 2802 -588
rect 1727 -3773 1779 -3721
rect 2743 -3644 2795 -3592
rect 1727 -4069 1779 -4017
rect 2743 -4071 2795 -4019
<< metal2 >>
rect 1404 1518 1456 1524
rect 1404 1460 1456 1466
rect 3210 1518 3262 1524
rect 3210 1460 3262 1466
rect 57 1114 113 1121
rect 876 1114 932 1121
rect -448 1054 -439 1114
rect -379 1054 -370 1114
rect 49 1054 55 1114
rect 115 1054 121 1114
rect 868 1054 874 1114
rect 934 1054 940 1114
rect 57 1047 113 1054
rect 876 1047 932 1054
rect 1416 856 1444 1460
rect 3222 939 3250 1460
rect 3749 1114 3805 1121
rect 4578 1114 4634 1121
rect 3741 1054 3747 1114
rect 3807 1054 3813 1114
rect 4570 1054 4576 1114
rect 4636 1054 4642 1114
rect 3749 1047 3805 1054
rect 4578 1047 4634 1054
rect 3204 887 3210 939
rect 3262 887 3268 939
rect 1919 861 1971 867
rect 1398 804 1404 856
rect 1456 804 1462 856
rect 2414 849 2420 861
rect 1971 821 2420 849
rect 2414 809 2420 821
rect 2472 809 2478 861
rect 1919 803 1971 809
rect 2137 785 2189 791
rect 2864 773 2870 785
rect 2189 745 2870 773
rect 2864 733 2870 745
rect 2922 733 2928 785
rect 2137 727 2189 733
rect 1924 -594 1980 -587
rect 2744 -588 2800 -581
rect 1916 -654 1922 -594
rect 1982 -654 1988 -594
rect 2736 -648 2742 -588
rect 2802 -648 2808 -588
rect 1924 -661 1980 -654
rect 2744 -655 2800 -648
rect 2737 -3644 2743 -3592
rect 2795 -3644 2801 -3592
rect 1721 -3773 1727 -3721
rect 1779 -3773 1785 -3721
rect 1738 -4011 1768 -3773
rect 1727 -4017 1779 -4011
rect 2754 -4013 2784 -3644
rect 1727 -4075 1779 -4069
rect 2743 -4019 2795 -4013
rect 2743 -4077 2795 -4071
<< via2 >>
rect -439 1110 -379 1114
rect -439 1058 -435 1110
rect -435 1058 -383 1110
rect -383 1058 -379 1110
rect -439 1054 -379 1058
rect 57 1056 113 1112
rect 876 1056 932 1112
rect 3749 1056 3805 1112
rect 4578 1056 4634 1112
rect 1924 -652 1980 -596
rect 2744 -646 2800 -590
<< metal3 >>
rect -444 1114 -374 1119
rect 52 1114 118 1117
rect 871 1114 937 1117
rect 3744 1114 3810 1117
rect 4573 1114 4639 1117
rect -444 1054 -439 1114
rect -379 1112 4639 1114
rect -379 1056 57 1112
rect 113 1056 876 1112
rect 932 1056 3749 1112
rect 3805 1056 4578 1112
rect 4634 1056 4639 1112
rect -379 1054 4639 1056
rect -444 1049 -374 1054
rect 52 1051 118 1054
rect 871 1051 937 1054
rect 2226 -588 2286 1054
rect 3744 1051 3810 1054
rect 4573 1051 4639 1054
rect 2739 -588 2805 -585
rect 2226 -590 2805 -588
rect 1919 -594 1985 -591
rect 2226 -594 2744 -590
rect 1919 -596 2744 -594
rect 1919 -652 1924 -596
rect 1980 -646 2744 -596
rect 2800 -646 2805 -590
rect 1980 -648 2805 -646
rect 1980 -652 2286 -648
rect 2739 -651 2805 -648
rect 1919 -654 2286 -652
rect 1919 -657 1985 -654
use sky130_fd_pr__nfet_01v8  sky130_fd_pr__nfet_01v8_0
timestamp 1696114978
transform 0 -1 1878 -1 0 -14
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8  sky130_fd_pr__nfet_01v8_1
timestamp 1696114978
transform 0 1 2811 -1 0 -19
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8  sky130_fd_pr__nfet_01v8_2
timestamp 1696114978
transform 0 1 1882 -1 0 498
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8  sky130_fd_pr__nfet_01v8_3
timestamp 1696114978
transform 0 -1 2814 -1 0 502
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8  sky130_fd_pr__nfet_01v8_4
timestamp 1696114978
transform 0 1 2643 -1 0 -624
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8  sky130_fd_pr__nfet_01v8_5
timestamp 1696114978
transform 0 -1 2077 -1 0 -620
box -226 -279 226 279
use sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_0
timestamp 1696114596
transform 0 -1 2820 1 0 1068
box -226 -284 226 284
use sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_1
timestamp 1696114596
transform 0 1 1864 1 0 1076
box -226 -284 226 284
use sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_2
timestamp 1696114596
transform 0 1 3650 1 0 1068
box -226 -284 226 284
use sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_3
timestamp 1696114596
transform 0 -1 1034 1 0 1076
box -226 -284 226 284
use sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_4
timestamp 1696114596
transform 0 -1 212 1 0 1080
box -226 -284 226 284
use sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_5
timestamp 1696114596
transform 0 1 4472 1 0 1072
box -226 -284 226 284
use trim  trim_0
timestamp 1696279213
transform 0 -1 8203 -1 0 697
box -43 2464 4673 5034
use trim  trim_1
timestamp 1696279213
transform 0 1 -3412 -1 0 715
box -43 2464 4673 5034
<< labels >>
flabel metal1 1840 49 1869 448 0 FreeSans 640 0 0 0 IN
flabel metal1 2810 47 2839 446 0 FreeSans 640 0 0 0 IP
flabel metal1 1416 1532 1444 1560 0 FreeSans 640 0 0 0 outn
port 4 nsew
flabel metal1 3223 1518 3252 1555 0 FreeSans 640 0 0 0 outp
port 5 nsew
flabel metal1 2169 -319 2199 -289 0 FreeSans 640 0 0 0 diff
flabel via1 1727 -4069 1779 -4017 0 FreeSans 640 0 0 0 vn
port 2 nsew
flabel via1 2743 -4071 2795 -4019 0 FreeSans 640 0 0 0 vp
port 3 nsew
flabel metal1 2140 -4059 2170 -4029 0 FreeSans 640 0 0 0 vss
port 1 nsew
flabel metal1 2286 1473 2314 1501 0 FreeSans 640 0 0 0 vdd
port 0 nsew
flabel metal1 -443 1552 -375 1625 0 FreeSans 640 0 0 0 clk
port 6 nsew
flabel metal1 395 -3974 429 -3946 0 FreeSans 160 0 0 0 trim0
port 7 nsew
flabel metal1 251 -3975 285 -3947 0 FreeSans 160 0 0 0 trim1
port 8 nsew
flabel metal1 162 -3975 196 -3947 0 FreeSans 160 0 0 0 trim2
port 9 nsew
flabel metal1 87 -3975 121 -3947 0 FreeSans 160 0 0 0 trim3
port 10 nsew
flabel metal1 25 -3975 59 -3947 0 FreeSans 160 0 0 0 trim4
port 11 nsew
flabel metal1 4364 -3990 4398 -3962 0 FreeSans 160 0 0 0 trimb0
port 12 nsew
flabel metal1 4506 -3985 4540 -3957 0 FreeSans 160 0 0 0 trimb1
port 13 nsew
flabel metal1 4596 -3985 4630 -3957 0 FreeSans 160 0 0 0 trimb2
port 14 nsew
flabel metal1 4671 -3985 4705 -3957 0 FreeSans 160 0 0 0 trimb3
port 15 nsew
flabel metal1 4733 -3985 4767 -3957 0 FreeSans 160 0 0 0 trimb4
port 16 nsew
<< end >>
