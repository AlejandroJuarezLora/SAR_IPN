magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< pwell >>
rect 8130 1576 8766 1662
rect 8130 1197 8216 1576
rect 8680 1197 8766 1576
rect 8130 1111 8766 1197
<< psubdiff >>
rect 8156 1602 8370 1636
rect 8404 1602 8438 1636
rect 8472 1602 8506 1636
rect 8540 1602 8740 1636
rect 8156 1436 8190 1602
rect 8156 1171 8190 1402
rect 8706 1436 8740 1602
rect 8706 1171 8740 1402
rect 8156 1137 8370 1171
rect 8404 1137 8438 1171
rect 8472 1137 8506 1171
rect 8540 1137 8740 1171
<< psubdiffcont >>
rect 8370 1602 8404 1636
rect 8438 1602 8472 1636
rect 8506 1602 8540 1636
rect 8156 1402 8190 1436
rect 8706 1402 8740 1436
rect 8370 1137 8404 1171
rect 8438 1137 8472 1171
rect 8506 1137 8540 1171
<< locali >>
rect 8156 1602 8370 1636
rect 8404 1602 8438 1636
rect 8472 1602 8506 1636
rect 8540 1602 8740 1636
rect 8156 1436 8190 1602
rect 8156 1171 8190 1402
rect 8706 1436 8740 1602
rect 8706 1171 8740 1402
rect 8156 1137 8370 1171
rect 8404 1137 8438 1171
rect 8472 1137 8506 1171
rect 8540 1137 8740 1171
<< properties >>
string path 40.780 8.095 43.615 8.095 43.615 5.770 40.865 5.770 40.865 8.095 
<< end >>
