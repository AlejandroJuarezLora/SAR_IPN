magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_p >>
rect -29 105 29 111
rect -29 71 -17 105
rect -29 65 29 71
<< nwell >>
rect -124 -238 124 124
<< pmos >>
rect -30 -176 30 24
<< pdiff >>
rect -88 9 -30 24
rect -88 -25 -76 9
rect -42 -25 -30 9
rect -88 -59 -30 -25
rect -88 -93 -76 -59
rect -42 -93 -30 -59
rect -88 -127 -30 -93
rect -88 -161 -76 -127
rect -42 -161 -30 -127
rect -88 -176 -30 -161
rect 30 9 88 24
rect 30 -25 42 9
rect 76 -25 88 9
rect 30 -59 88 -25
rect 30 -93 42 -59
rect 76 -93 88 -59
rect 30 -127 88 -93
rect 30 -161 42 -127
rect 76 -161 88 -127
rect 30 -176 88 -161
<< pdiffc >>
rect -76 -25 -42 9
rect -76 -93 -42 -59
rect -76 -161 -42 -127
rect 42 -25 76 9
rect 42 -93 76 -59
rect 42 -161 76 -127
<< poly >>
rect -33 105 33 121
rect -33 71 -17 105
rect 17 71 33 105
rect -33 55 33 71
rect -30 24 30 55
rect -30 -202 30 -176
<< polycont >>
rect -17 71 17 105
<< locali >>
rect -33 71 -17 105
rect 17 71 33 105
rect -76 9 -42 28
rect -76 -59 -42 -57
rect -76 -95 -42 -93
rect -76 -180 -42 -161
rect 42 9 76 28
rect 42 -59 76 -57
rect 42 -95 76 -93
rect 42 -180 76 -161
<< viali >>
rect -17 71 17 105
rect -76 -25 -42 -23
rect -76 -57 -42 -25
rect -76 -127 -42 -95
rect -76 -129 -42 -127
rect 42 -25 76 -23
rect 42 -57 76 -25
rect 42 -127 76 -95
rect 42 -129 76 -127
<< metal1 >>
rect -29 105 29 111
rect -29 71 -17 105
rect 17 71 29 105
rect -29 65 29 71
rect -82 -23 -36 24
rect -82 -57 -76 -23
rect -42 -57 -36 -23
rect -82 -95 -36 -57
rect -82 -129 -76 -95
rect -42 -129 -36 -95
rect -82 -176 -36 -129
rect 36 -23 82 24
rect 36 -57 42 -23
rect 76 -57 82 -23
rect 36 -95 82 -57
rect 36 -129 42 -95
rect 76 -129 82 -95
rect 36 -176 82 -129
<< end >>
