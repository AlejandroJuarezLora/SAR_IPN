magic
tech sky130B
magscale 1 2
timestamp 1696114978
<< pwell >>
rect -226 -279 226 279
<< nmos >>
rect -30 -131 30 69
<< ndiff >>
rect -88 39 -30 69
rect -88 -101 -76 39
rect -42 -101 -30 39
rect -88 -131 -30 -101
rect 30 39 88 69
rect 30 -101 42 39
rect 76 -101 88 39
rect 30 -131 88 -101
<< ndiffc >>
rect -76 -101 -42 39
rect 42 -101 76 39
<< psubdiff >>
rect -190 209 190 243
rect -190 -209 -156 209
rect 156 -209 190 209
rect -190 -243 -75 -209
rect 75 -243 190 -209
<< psubdiffcont >>
rect -75 -243 75 -209
<< poly >>
rect -33 141 33 157
rect -33 107 -17 141
rect 17 107 33 141
rect -33 91 33 107
rect -30 69 30 91
rect -30 -157 30 -131
<< polycont >>
rect -17 107 17 141
<< locali >>
rect -33 107 -17 141
rect 17 107 33 141
rect -76 39 -42 55
rect -76 -117 -42 -101
rect 42 39 76 55
rect 42 -117 76 -101
rect -91 -243 -75 -209
rect 75 -243 91 -209
<< viali >>
rect -17 107 17 141
rect -76 -101 -42 39
rect 42 -84 76 22
<< metal1 >>
rect -30 141 30 154
rect -30 107 -17 141
rect 17 107 30 141
rect -30 96 30 107
rect -82 39 -36 51
rect -82 -101 -76 39
rect -42 -101 -36 39
rect 36 22 82 34
rect 36 -84 42 22
rect 76 -84 82 22
rect 36 -96 82 -84
rect -82 -113 -36 -101
<< labels >>
flabel metal1 -82 -113 -76 51 0 FreeSans 480 0 0 0 D
port 0 nsew
flabel metal1 76 -96 82 34 0 FreeSans 480 0 0 0 S
port 1 nsew
flabel metal1 -30 141 30 154 0 FreeSans 480 0 0 0 G
port 2 nsew
flabel locali -91 -243 -75 -209 0 FreeSans 480 0 0 0 B
port 3 nsew
<< properties >>
string FIXED_BBOX -173 -226 173 226
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.3 m 1 nf 1 diffcov 80 polycov 80 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 80 rlcov 80 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 60 viadrn 80 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
