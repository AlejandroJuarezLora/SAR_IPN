magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< pwell >>
rect 2250 -495 5032 -409
rect 2250 -901 2336 -495
rect 4946 -901 5032 -495
rect 2250 -987 5032 -901
<< psubdiff >>
rect 2276 -469 2460 -435
rect 2494 -469 2528 -435
rect 2562 -469 2596 -435
rect 2630 -469 2664 -435
rect 2698 -469 2732 -435
rect 2766 -469 2800 -435
rect 2834 -469 2868 -435
rect 2902 -469 2936 -435
rect 2970 -469 3004 -435
rect 3038 -469 3072 -435
rect 3106 -469 3140 -435
rect 3174 -469 3208 -435
rect 3242 -469 3276 -435
rect 3310 -469 3344 -435
rect 3378 -469 3412 -435
rect 3446 -469 3480 -435
rect 3514 -469 3548 -435
rect 3582 -469 3616 -435
rect 3650 -469 3684 -435
rect 3718 -469 3752 -435
rect 3786 -469 3820 -435
rect 3854 -469 3888 -435
rect 3922 -469 3956 -435
rect 3990 -469 4024 -435
rect 4058 -469 4092 -435
rect 4126 -469 4160 -435
rect 4194 -469 4228 -435
rect 4262 -469 4296 -435
rect 4330 -469 4364 -435
rect 4398 -469 4432 -435
rect 4466 -469 4500 -435
rect 4534 -469 4568 -435
rect 4602 -469 4636 -435
rect 4670 -469 4704 -435
rect 4738 -469 4772 -435
rect 4806 -469 5006 -435
rect 2276 -659 2310 -469
rect 2276 -727 2310 -693
rect 2276 -927 2310 -761
rect 4972 -659 5006 -469
rect 4972 -727 5006 -693
rect 4972 -927 5006 -761
rect 2276 -961 2528 -927
rect 2562 -961 2596 -927
rect 2630 -961 2664 -927
rect 2698 -961 2732 -927
rect 2766 -961 2800 -927
rect 2834 -961 2868 -927
rect 2902 -961 2936 -927
rect 2970 -961 3004 -927
rect 3038 -961 3072 -927
rect 3106 -961 3140 -927
rect 3174 -961 3208 -927
rect 3242 -961 3276 -927
rect 3310 -961 3344 -927
rect 3378 -961 3412 -927
rect 3446 -961 3480 -927
rect 3514 -961 3548 -927
rect 3582 -961 3616 -927
rect 3650 -961 3684 -927
rect 3718 -961 3752 -927
rect 3786 -961 3820 -927
rect 3854 -961 3888 -927
rect 3922 -961 3956 -927
rect 3990 -961 4024 -927
rect 4058 -961 4092 -927
rect 4126 -961 4160 -927
rect 4194 -961 4228 -927
rect 4262 -961 4296 -927
rect 4330 -961 4364 -927
rect 4398 -961 4432 -927
rect 4466 -961 4500 -927
rect 4534 -961 4568 -927
rect 4602 -961 4636 -927
rect 4670 -961 4704 -927
rect 4738 -961 4772 -927
rect 4806 -961 5006 -927
<< psubdiffcont >>
rect 2460 -469 2494 -435
rect 2528 -469 2562 -435
rect 2596 -469 2630 -435
rect 2664 -469 2698 -435
rect 2732 -469 2766 -435
rect 2800 -469 2834 -435
rect 2868 -469 2902 -435
rect 2936 -469 2970 -435
rect 3004 -469 3038 -435
rect 3072 -469 3106 -435
rect 3140 -469 3174 -435
rect 3208 -469 3242 -435
rect 3276 -469 3310 -435
rect 3344 -469 3378 -435
rect 3412 -469 3446 -435
rect 3480 -469 3514 -435
rect 3548 -469 3582 -435
rect 3616 -469 3650 -435
rect 3684 -469 3718 -435
rect 3752 -469 3786 -435
rect 3820 -469 3854 -435
rect 3888 -469 3922 -435
rect 3956 -469 3990 -435
rect 4024 -469 4058 -435
rect 4092 -469 4126 -435
rect 4160 -469 4194 -435
rect 4228 -469 4262 -435
rect 4296 -469 4330 -435
rect 4364 -469 4398 -435
rect 4432 -469 4466 -435
rect 4500 -469 4534 -435
rect 4568 -469 4602 -435
rect 4636 -469 4670 -435
rect 4704 -469 4738 -435
rect 4772 -469 4806 -435
rect 2276 -693 2310 -659
rect 2276 -761 2310 -727
rect 4972 -693 5006 -659
rect 4972 -761 5006 -727
rect 2528 -961 2562 -927
rect 2596 -961 2630 -927
rect 2664 -961 2698 -927
rect 2732 -961 2766 -927
rect 2800 -961 2834 -927
rect 2868 -961 2902 -927
rect 2936 -961 2970 -927
rect 3004 -961 3038 -927
rect 3072 -961 3106 -927
rect 3140 -961 3174 -927
rect 3208 -961 3242 -927
rect 3276 -961 3310 -927
rect 3344 -961 3378 -927
rect 3412 -961 3446 -927
rect 3480 -961 3514 -927
rect 3548 -961 3582 -927
rect 3616 -961 3650 -927
rect 3684 -961 3718 -927
rect 3752 -961 3786 -927
rect 3820 -961 3854 -927
rect 3888 -961 3922 -927
rect 3956 -961 3990 -927
rect 4024 -961 4058 -927
rect 4092 -961 4126 -927
rect 4160 -961 4194 -927
rect 4228 -961 4262 -927
rect 4296 -961 4330 -927
rect 4364 -961 4398 -927
rect 4432 -961 4466 -927
rect 4500 -961 4534 -927
rect 4568 -961 4602 -927
rect 4636 -961 4670 -927
rect 4704 -961 4738 -927
rect 4772 -961 4806 -927
<< locali >>
rect 2276 -469 2460 -435
rect 2494 -469 2528 -435
rect 2562 -469 2596 -435
rect 2630 -469 2664 -435
rect 2698 -469 2732 -435
rect 2766 -469 2800 -435
rect 2834 -469 2868 -435
rect 2902 -469 2936 -435
rect 2970 -469 3004 -435
rect 3038 -469 3072 -435
rect 3106 -469 3140 -435
rect 3174 -469 3208 -435
rect 3242 -469 3276 -435
rect 3310 -469 3344 -435
rect 3378 -469 3412 -435
rect 3446 -469 3480 -435
rect 3514 -469 3548 -435
rect 3582 -469 3616 -435
rect 3650 -469 3684 -435
rect 3718 -469 3752 -435
rect 3786 -469 3820 -435
rect 3854 -469 3888 -435
rect 3922 -469 3956 -435
rect 3990 -469 4024 -435
rect 4058 -469 4092 -435
rect 4126 -469 4160 -435
rect 4194 -469 4228 -435
rect 4262 -469 4296 -435
rect 4330 -469 4364 -435
rect 4398 -469 4432 -435
rect 4466 -469 4500 -435
rect 4534 -469 4568 -435
rect 4602 -469 4636 -435
rect 4670 -469 4704 -435
rect 4738 -469 4772 -435
rect 4806 -469 5006 -435
rect 2276 -659 2310 -469
rect 2276 -727 2310 -693
rect 2276 -927 2310 -761
rect 4972 -659 5006 -469
rect 4972 -727 5006 -693
rect 4972 -927 5006 -761
rect 2276 -961 2528 -927
rect 2562 -961 2596 -927
rect 2630 -961 2664 -927
rect 2698 -961 2732 -927
rect 2766 -961 2800 -927
rect 2834 -961 2868 -927
rect 2902 -961 2936 -927
rect 2970 -961 3004 -927
rect 3038 -961 3072 -927
rect 3106 -961 3140 -927
rect 3174 -961 3208 -927
rect 3242 -961 3276 -927
rect 3310 -961 3344 -927
rect 3378 -961 3412 -927
rect 3446 -961 3480 -927
rect 3514 -961 3548 -927
rect 3582 -961 3616 -927
rect 3650 -961 3684 -927
rect 3718 -961 3752 -927
rect 3786 -961 3820 -927
rect 3854 -961 3888 -927
rect 3922 -961 3956 -927
rect 3990 -961 4024 -927
rect 4058 -961 4092 -927
rect 4126 -961 4160 -927
rect 4194 -961 4228 -927
rect 4262 -961 4296 -927
rect 4330 -961 4364 -927
rect 4398 -961 4432 -927
rect 4466 -961 4500 -927
rect 4534 -961 4568 -927
rect 4602 -961 4636 -927
rect 4670 -961 4704 -927
rect 4738 -961 4772 -927
rect 4806 -961 5006 -927
<< properties >>
string path 11.380 -2.260 24.945 -2.260 24.945 -4.720 11.465 -4.720 11.465 -2.260 
<< end >>
