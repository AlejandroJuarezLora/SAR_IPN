magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 590 542
<< pwell >>
rect 1 -19 551 163
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 109 137
rect 267 7 297 137
rect 359 7 389 137
rect 443 7 473 137
<< scpmoshvt >>
rect 83 257 113 457
rect 244 257 274 457
rect 352 257 382 457
rect 443 257 473 457
<< ndiff >>
rect 27 124 79 137
rect 27 90 35 124
rect 69 90 79 124
rect 27 56 79 90
rect 27 22 35 56
rect 69 22 79 56
rect 27 7 79 22
rect 109 53 161 137
rect 109 19 119 53
rect 153 19 161 53
rect 109 7 161 19
rect 215 125 267 137
rect 215 91 223 125
rect 257 91 267 125
rect 215 57 267 91
rect 215 23 223 57
rect 257 23 267 57
rect 215 7 267 23
rect 297 121 359 137
rect 297 87 315 121
rect 349 87 359 121
rect 297 7 359 87
rect 389 53 443 137
rect 389 19 399 53
rect 433 19 443 53
rect 389 7 443 19
rect 473 125 525 137
rect 473 91 483 125
rect 517 91 525 125
rect 473 57 525 91
rect 473 23 483 57
rect 517 23 525 57
rect 473 7 525 23
<< pdiff >>
rect 27 437 83 457
rect 27 403 39 437
rect 73 403 83 437
rect 27 369 83 403
rect 27 335 39 369
rect 73 335 83 369
rect 27 301 83 335
rect 27 267 39 301
rect 73 267 83 301
rect 27 257 83 267
rect 113 445 244 457
rect 113 411 125 445
rect 159 411 199 445
rect 233 411 244 445
rect 113 377 244 411
rect 113 343 125 377
rect 159 343 199 377
rect 233 343 244 377
rect 113 257 244 343
rect 274 445 352 457
rect 274 411 299 445
rect 333 411 352 445
rect 274 377 352 411
rect 274 343 299 377
rect 333 343 352 377
rect 274 309 352 343
rect 274 275 299 309
rect 333 275 352 309
rect 274 257 352 275
rect 382 257 443 457
rect 473 445 525 457
rect 473 411 483 445
rect 517 411 525 445
rect 473 377 525 411
rect 473 343 483 377
rect 517 343 525 377
rect 473 257 525 343
<< ndiffc >>
rect 35 90 69 124
rect 35 22 69 56
rect 119 19 153 53
rect 223 91 257 125
rect 223 23 257 57
rect 315 87 349 121
rect 399 19 433 53
rect 483 91 517 125
rect 483 23 517 57
<< pdiffc >>
rect 39 403 73 437
rect 39 335 73 369
rect 39 267 73 301
rect 125 411 159 445
rect 199 411 233 445
rect 125 343 159 377
rect 199 343 233 377
rect 299 411 333 445
rect 299 343 333 377
rect 299 275 333 309
rect 483 411 517 445
rect 483 343 517 377
<< poly >>
rect 83 457 113 483
rect 244 457 274 483
rect 352 457 382 483
rect 443 457 473 483
rect 83 225 113 257
rect 244 225 274 257
rect 352 225 382 257
rect 443 229 473 257
rect 79 209 163 225
rect 79 175 119 209
rect 153 175 163 209
rect 79 159 163 175
rect 244 209 301 225
rect 244 175 257 209
rect 291 175 301 209
rect 244 159 301 175
rect 347 209 401 225
rect 347 175 357 209
rect 391 175 401 209
rect 347 159 401 175
rect 443 209 529 229
rect 443 175 485 209
rect 519 175 529 209
rect 443 159 529 175
rect 79 137 109 159
rect 267 137 297 159
rect 359 137 389 159
rect 443 137 473 159
rect 79 -19 109 7
rect 267 -19 297 7
rect 359 -19 389 7
rect 443 -19 473 7
<< polycont >>
rect 119 175 153 209
rect 257 175 291 209
rect 357 175 391 209
rect 485 175 519 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 552 521
rect 17 437 73 453
rect 17 403 39 437
rect 17 369 73 403
rect 17 335 39 369
rect 17 301 73 335
rect 107 445 249 487
rect 107 411 125 445
rect 159 411 199 445
rect 233 411 249 445
rect 107 377 249 411
rect 107 343 125 377
rect 159 343 199 377
rect 233 343 249 377
rect 107 332 249 343
rect 283 445 349 453
rect 283 411 299 445
rect 333 411 349 445
rect 467 445 533 487
rect 283 377 349 411
rect 283 343 299 377
rect 333 343 349 377
rect 17 267 39 301
rect 283 309 349 343
rect 283 298 299 309
rect 17 166 73 267
rect 119 275 299 298
rect 333 275 349 309
rect 119 255 349 275
rect 119 209 176 255
rect 153 175 176 209
rect 213 209 307 221
rect 388 215 431 438
rect 467 411 483 445
rect 517 411 533 445
rect 467 377 533 411
rect 467 343 483 377
rect 517 343 533 377
rect 489 215 535 283
rect 213 175 257 209
rect 291 175 307 209
rect 341 209 431 215
rect 341 175 357 209
rect 391 179 431 209
rect 469 209 535 215
rect 391 175 407 179
rect 469 175 485 209
rect 519 175 535 209
rect 17 124 85 166
rect 17 90 35 124
rect 69 90 85 124
rect 119 141 176 175
rect 119 125 261 141
rect 119 103 223 125
rect 17 56 85 90
rect 201 91 223 103
rect 257 91 261 125
rect 201 75 261 91
rect 299 125 535 141
rect 299 121 483 125
rect 299 87 315 121
rect 349 103 483 121
rect 349 87 365 103
rect 467 91 483 103
rect 517 91 535 125
rect 201 73 264 75
rect 201 71 266 73
rect 201 70 268 71
rect 17 22 35 56
rect 69 22 85 56
rect 17 11 85 22
rect 119 53 153 69
rect 119 -23 153 19
rect 201 68 269 70
rect 201 67 270 68
rect 201 65 271 67
rect 201 64 272 65
rect 201 57 273 64
rect 201 23 223 57
rect 257 23 273 57
rect 201 11 273 23
rect 399 53 433 69
rect 399 -23 433 19
rect 467 57 535 91
rect 467 23 483 57
rect 517 23 535 57
rect 467 11 535 23
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 552 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
<< metal1 >>
rect 0 521 552 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 552 521
rect 0 456 552 487
rect 0 -23 552 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 552 -23
rect 0 -88 552 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 o21a_1
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 29 317 63 351 0 FreeSans 340 0 0 0 X
port 10 nsew
flabel locali s 489 249 523 283 0 FreeSans 340 0 0 0 A1
port 7 nsew
flabel locali s 213 181 247 215 0 FreeSans 340 0 0 0 B1
port 9 nsew
flabel locali s 397 181 431 215 0 FreeSans 340 0 0 0 A2
port 8 nsew
<< properties >>
string FIXED_BBOX 0 -40 552 504
string path 0.000 -1.000 13.800 -1.000 
<< end >>
