magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 682 542
<< pwell >>
rect 1 -19 643 163
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 109 137
rect 155 7 185 137
rect 343 7 373 137
rect 443 7 473 137
rect 535 7 565 137
<< scpmoshvt >>
rect 79 257 109 457
rect 163 257 193 457
rect 349 257 379 457
rect 443 257 473 457
rect 535 257 565 457
<< ndiff >>
rect 27 125 79 137
rect 27 91 35 125
rect 69 91 79 125
rect 27 57 79 91
rect 27 23 35 57
rect 69 23 79 57
rect 27 7 79 23
rect 109 7 155 137
rect 185 53 237 137
rect 185 19 195 53
rect 229 19 237 53
rect 185 7 237 19
rect 291 53 343 137
rect 291 19 299 53
rect 333 19 343 53
rect 291 7 343 19
rect 373 7 443 137
rect 473 49 535 137
rect 473 15 491 49
rect 525 15 535 49
rect 473 7 535 15
rect 565 61 617 137
rect 565 27 575 61
rect 609 27 617 61
rect 565 7 617 27
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 377 79 411
rect 27 343 35 377
rect 69 343 79 377
rect 27 309 79 343
rect 27 275 35 309
rect 69 275 79 309
rect 27 257 79 275
rect 109 369 163 457
rect 109 335 119 369
rect 153 335 163 369
rect 109 257 163 335
rect 193 314 243 457
rect 297 445 349 457
rect 297 411 305 445
rect 339 411 349 445
rect 297 399 349 411
rect 193 303 245 314
rect 193 269 203 303
rect 237 269 245 303
rect 193 257 245 269
rect 299 257 349 399
rect 379 437 443 457
rect 379 403 391 437
rect 425 403 443 437
rect 379 369 443 403
rect 379 335 391 369
rect 425 335 443 369
rect 379 257 443 335
rect 473 449 535 457
rect 473 415 491 449
rect 525 415 535 449
rect 473 381 535 415
rect 473 347 491 381
rect 525 347 535 381
rect 473 257 535 347
rect 565 437 617 457
rect 565 403 575 437
rect 609 403 617 437
rect 565 369 617 403
rect 565 335 575 369
rect 609 335 617 369
rect 565 257 617 335
<< ndiffc >>
rect 35 91 69 125
rect 35 23 69 57
rect 195 19 229 53
rect 299 19 333 53
rect 491 15 525 49
rect 575 27 609 61
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 35 275 69 309
rect 119 335 153 369
rect 305 411 339 445
rect 203 269 237 303
rect 391 403 425 437
rect 391 335 425 369
rect 491 415 525 449
rect 491 347 525 381
rect 575 403 609 437
rect 575 335 609 369
<< poly >>
rect 79 457 109 483
rect 163 457 193 483
rect 349 457 379 483
rect 443 457 473 483
rect 535 457 565 483
rect 79 225 109 257
rect 163 225 193 257
rect 349 242 379 257
rect 327 231 379 242
rect 299 228 377 231
rect 299 227 376 228
rect 299 225 375 227
rect 443 225 473 257
rect 535 225 565 257
rect 55 209 109 225
rect 55 175 65 209
rect 99 175 109 209
rect 55 159 109 175
rect 79 137 109 159
rect 155 209 213 225
rect 155 175 169 209
rect 203 175 213 209
rect 155 159 213 175
rect 299 224 374 225
rect 423 224 473 225
rect 299 209 373 224
rect 421 221 473 224
rect 420 218 473 221
rect 419 215 473 218
rect 418 213 473 215
rect 299 175 313 209
rect 347 175 373 209
rect 299 159 373 175
rect 155 137 185 159
rect 343 137 373 159
rect 417 209 473 213
rect 417 175 429 209
rect 463 175 473 209
rect 417 152 473 175
rect 515 209 589 225
rect 515 175 525 209
rect 559 175 589 209
rect 515 159 589 175
rect 443 137 473 152
rect 535 137 565 159
rect 79 -19 109 7
rect 155 -19 185 7
rect 343 -19 373 7
rect 443 -19 473 7
rect 535 -19 565 7
<< polycont >>
rect 65 175 99 209
rect 169 175 203 209
rect 313 175 347 209
rect 429 175 463 209
rect 525 175 559 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 644 521
rect 18 445 85 453
rect 18 411 35 445
rect 69 411 85 445
rect 286 445 357 487
rect 286 411 305 445
rect 339 411 357 445
rect 391 437 441 453
rect 18 409 85 411
rect 18 377 69 409
rect 425 403 441 437
rect 18 343 35 377
rect 18 309 69 343
rect 119 377 165 385
rect 391 377 441 403
rect 119 369 441 377
rect 153 337 391 369
rect 153 335 156 337
rect 274 335 391 337
rect 425 335 441 369
rect 491 449 541 487
rect 525 415 541 449
rect 491 381 541 415
rect 525 347 541 381
rect 119 319 156 335
rect 491 331 541 347
rect 575 437 627 453
rect 609 403 627 437
rect 575 369 627 403
rect 609 335 627 369
rect 575 317 627 335
rect 18 275 35 309
rect 187 285 203 303
rect 69 275 203 285
rect 18 269 203 275
rect 237 297 253 303
rect 237 285 547 297
rect 237 269 559 285
rect 18 263 559 269
rect 18 251 253 263
rect 519 256 559 263
rect 17 209 115 215
rect 17 175 65 209
rect 99 175 115 209
rect 153 209 248 217
rect 153 175 169 209
rect 203 175 248 209
rect 18 125 109 130
rect 18 91 35 125
rect 69 91 109 125
rect 204 95 248 175
rect 297 209 363 217
rect 297 175 313 209
rect 347 175 363 209
rect 397 209 479 229
rect 397 175 429 209
rect 463 175 479 209
rect 297 95 339 175
rect 397 168 479 175
rect 525 209 559 256
rect 525 141 559 175
rect 505 117 559 141
rect 390 108 559 117
rect 18 57 109 91
rect 18 23 35 57
rect 69 23 109 57
rect 390 83 541 108
rect 390 53 424 83
rect 593 77 627 317
rect 18 -23 109 23
rect 164 19 195 53
rect 229 19 299 53
rect 333 19 424 53
rect 575 61 627 77
rect 164 11 424 19
rect 475 15 491 49
rect 525 15 541 49
rect 475 -23 541 15
rect 609 27 627 61
rect 575 11 627 27
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 644 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
<< metal1 >>
rect 0 521 644 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 644 521
rect 0 456 644 487
rect 0 -23 644 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 644 -23
rect 0 -88 644 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 a22o_1
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 305 181 339 215 0 FreeSans 200 0 0 0 A1
port 8 nsew
flabel locali s 397 181 431 215 0 FreeSans 200 0 0 0 A2
port 9 nsew
flabel locali s 581 385 615 419 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel locali s 30 181 64 215 0 FreeSans 200 0 0 0 B2
port 11 nsew
flabel locali s 214 181 248 215 0 FreeSans 200 0 0 0 B1
port 7 nsew
flabel locali s 305 113 339 147 0 FreeSans 200 0 0 0 A1
port 8 nsew
flabel locali s 214 113 248 147 0 FreeSans 200 0 0 0 B1
port 7 nsew
flabel locali s 581 317 615 351 0 FreeSans 200 0 0 0 X
port 10 nsew
<< properties >>
string FIXED_BBOX 0 -40 644 504
string path 0.000 -1.000 16.100 -1.000 
<< end >>
