magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 498 542
<< pwell >>
rect 268 123 459 163
rect 3 -13 459 123
rect 28 -57 62 -13
rect 268 -19 459 -13
<< scnmos >>
rect 81 13 111 97
rect 165 13 195 97
rect 249 13 279 97
rect 347 7 377 137
<< scpmoshvt >>
rect 81 257 111 341
rect 153 257 183 341
rect 249 257 279 341
rect 347 257 377 457
<< ndiff >>
rect 294 97 347 137
rect 29 71 81 97
rect 29 37 37 71
rect 71 37 81 71
rect 29 13 81 37
rect 111 57 165 97
rect 111 23 121 57
rect 155 23 165 57
rect 111 13 165 23
rect 195 71 249 97
rect 195 37 205 71
rect 239 37 249 71
rect 195 13 249 37
rect 279 57 347 97
rect 279 23 299 57
rect 333 23 347 57
rect 279 13 347 23
rect 294 7 347 13
rect 377 95 433 137
rect 377 61 387 95
rect 421 61 433 95
rect 377 7 433 61
<< pdiff >>
rect 294 445 347 457
rect 294 411 302 445
rect 336 411 347 445
rect 294 377 347 411
rect 294 343 302 377
rect 336 343 347 377
rect 294 341 347 343
rect 29 314 81 341
rect 29 280 37 314
rect 71 280 81 314
rect 29 257 81 280
rect 111 257 153 341
rect 183 257 249 341
rect 279 257 347 341
rect 377 414 433 457
rect 377 380 387 414
rect 421 380 433 414
rect 377 346 433 380
rect 377 312 387 346
rect 421 312 433 346
rect 377 257 433 312
<< ndiffc >>
rect 37 37 71 71
rect 121 23 155 57
rect 205 37 239 71
rect 299 23 333 57
rect 387 61 421 95
<< pdiffc >>
rect 302 411 336 445
rect 302 343 336 377
rect 37 280 71 314
rect 387 380 421 414
rect 387 312 421 346
<< poly >>
rect 347 457 377 483
rect 147 433 213 443
rect 147 399 163 433
rect 197 399 213 433
rect 147 389 213 399
rect 81 341 111 367
rect 153 341 183 389
rect 249 341 279 367
rect 81 225 111 257
rect 24 209 111 225
rect 24 175 34 209
rect 68 175 111 209
rect 24 159 111 175
rect 81 97 111 159
rect 153 142 183 257
rect 249 225 279 257
rect 347 225 377 257
rect 234 209 288 225
rect 234 175 244 209
rect 278 175 288 209
rect 234 159 288 175
rect 330 209 384 225
rect 330 175 340 209
rect 374 175 384 209
rect 330 159 384 175
rect 153 112 195 142
rect 165 97 195 112
rect 249 97 279 159
rect 347 137 377 159
rect 81 -13 111 13
rect 165 -13 195 13
rect 249 -13 279 13
rect 347 -19 377 7
<< polycont >>
rect 163 399 197 433
rect 34 175 68 209
rect 244 175 278 209
rect 340 175 374 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 289 445 345 487
rect 17 433 255 443
rect 17 399 163 433
rect 197 399 255 433
rect 17 385 255 399
rect 289 411 302 445
rect 336 411 345 445
rect 289 377 345 411
rect 21 317 255 351
rect 289 343 302 377
rect 336 343 345 377
rect 289 327 345 343
rect 387 414 442 453
rect 421 380 442 414
rect 387 346 442 380
rect 21 314 86 317
rect 21 280 37 314
rect 71 280 86 314
rect 221 293 255 317
rect 421 312 442 346
rect 21 259 86 280
rect 120 225 159 283
rect 221 259 353 293
rect 387 259 442 312
rect 319 225 353 259
rect 17 209 86 225
rect 17 175 34 209
rect 68 175 86 209
rect 17 159 86 175
rect 120 209 285 225
rect 120 175 244 209
rect 278 175 285 209
rect 120 159 285 175
rect 319 209 374 225
rect 319 175 340 209
rect 319 159 374 175
rect 319 125 353 159
rect 20 91 353 125
rect 408 112 442 259
rect 387 95 442 112
rect 20 71 71 91
rect 20 37 37 71
rect 205 71 239 91
rect 20 21 71 37
rect 105 23 121 57
rect 155 23 171 57
rect 105 -23 171 23
rect 421 61 442 95
rect 205 21 239 37
rect 273 23 299 57
rect 333 23 349 57
rect 387 43 442 61
rect 273 -23 349 23
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
<< metal1 >>
rect 0 521 460 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 460 521
rect 0 456 460 487
rect 0 -23 460 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 460 -23
rect 0 -88 460 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 or3_1
flabel metal1 s 28 487 62 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 28 -57 62 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 28 487 62 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 28 -57 62 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 212 181 246 215 0 FreeSans 400 0 0 0 A
port 9 nsew
flabel locali s 120 181 154 215 0 FreeSans 400 0 0 0 A
port 9 nsew
flabel locali s 396 317 430 351 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel locali s 120 249 154 283 0 FreeSans 400 0 0 0 A
port 9 nsew
flabel locali s 28 385 62 419 0 FreeSans 400 0 0 0 B
port 7 nsew
flabel locali s 120 385 154 419 0 FreeSans 400 0 0 0 B
port 7 nsew
flabel locali s 28 181 62 215 0 FreeSans 400 0 0 0 C
port 8 nsew
<< properties >>
string FIXED_BBOX 0 -40 460 504
string path 0.000 -1.000 11.500 -1.000 
<< end >>
