magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect 0 269 352 590
<< pwell >>
rect 41 29 311 211
<< scnmos >>
rect 119 55 149 185
rect 203 55 233 185
<< scpmoshvt >>
rect 119 305 149 505
rect 203 305 233 505
<< ndiff >>
rect 67 173 119 185
rect 67 139 75 173
rect 109 139 119 173
rect 67 101 119 139
rect 67 67 75 101
rect 109 67 119 101
rect 67 55 119 67
rect 149 173 203 185
rect 149 139 159 173
rect 193 139 203 173
rect 149 101 203 139
rect 149 67 159 101
rect 193 67 203 101
rect 149 55 203 67
rect 233 173 285 185
rect 233 139 243 173
rect 277 139 285 173
rect 233 101 285 139
rect 233 67 243 101
rect 277 67 285 101
rect 233 55 285 67
<< pdiff >>
rect 67 493 119 505
rect 67 459 75 493
rect 109 459 119 493
rect 67 425 119 459
rect 67 391 75 425
rect 109 391 119 425
rect 67 357 119 391
rect 67 323 75 357
rect 109 323 119 357
rect 67 305 119 323
rect 149 493 203 505
rect 149 459 159 493
rect 193 459 203 493
rect 149 425 203 459
rect 149 391 159 425
rect 193 391 203 425
rect 149 357 203 391
rect 149 323 159 357
rect 193 323 203 357
rect 149 305 203 323
rect 233 493 285 505
rect 233 459 243 493
rect 277 459 285 493
rect 233 425 285 459
rect 233 391 243 425
rect 277 391 285 425
rect 233 357 285 391
rect 233 323 243 357
rect 277 323 285 357
rect 233 305 285 323
<< ndiffc >>
rect 75 139 109 173
rect 75 67 109 101
rect 159 139 193 173
rect 159 67 193 101
rect 243 139 277 173
rect 243 67 277 101
<< pdiffc >>
rect 75 459 109 493
rect 75 391 109 425
rect 75 323 109 357
rect 159 459 193 493
rect 159 391 193 425
rect 159 323 193 357
rect 243 459 277 493
rect 243 391 277 425
rect 243 323 277 357
<< poly >>
rect 119 505 149 531
rect 203 505 233 531
rect 119 273 149 305
rect 203 273 233 305
rect 59 257 233 273
rect 59 223 75 257
rect 109 223 233 257
rect 59 207 233 223
rect 119 185 149 207
rect 203 185 233 207
rect 119 29 149 55
rect 203 29 233 55
<< polycont >>
rect 75 223 109 257
<< locali >>
rect 38 535 67 569
rect 101 535 159 569
rect 193 535 251 569
rect 285 535 314 569
rect 63 493 109 535
rect 63 459 75 493
rect 63 425 109 459
rect 63 391 75 425
rect 63 357 109 391
rect 63 323 75 357
rect 63 307 109 323
rect 143 493 209 501
rect 143 459 159 493
rect 193 459 209 493
rect 143 425 209 459
rect 143 391 159 425
rect 193 391 209 425
rect 143 357 209 391
rect 143 323 159 357
rect 193 323 209 357
rect 143 305 209 323
rect 243 493 285 535
rect 277 459 285 493
rect 243 425 285 459
rect 277 391 285 425
rect 243 357 285 391
rect 277 323 285 357
rect 243 307 285 323
rect 59 257 125 273
rect 59 223 75 257
rect 109 223 125 257
rect 63 173 109 189
rect 159 185 209 305
rect 63 139 75 173
rect 63 101 109 139
rect 63 67 75 101
rect 63 25 109 67
rect 143 173 209 185
rect 143 139 159 173
rect 193 139 209 173
rect 143 101 209 139
rect 143 67 159 101
rect 193 67 209 101
rect 143 59 209 67
rect 243 173 285 189
rect 277 139 285 173
rect 243 101 285 139
rect 277 67 285 101
rect 243 25 285 67
rect 38 -9 67 25
rect 101 -9 159 25
rect 193 -9 251 25
rect 285 -9 314 25
<< viali >>
rect 67 535 101 569
rect 159 535 193 569
rect 251 535 285 569
rect 67 -9 101 25
rect 159 -9 193 25
rect 251 -9 285 25
<< metal1 >>
rect 38 569 314 600
rect 38 535 67 569
rect 101 535 159 569
rect 193 535 251 569
rect 285 535 314 569
rect 38 504 314 535
rect 38 25 314 56
rect 38 -9 67 25
rect 101 -9 159 25
rect 193 -9 251 25
rect 285 -9 314 25
rect 38 -40 314 -9
<< labels >>
rlabel comment s 38 8 38 8 4 inv_2
flabel comment s 84 246 84 246 0 FreeSans 340 0 0 0 A
flabel comment s 176 178 176 178 0 FreeSans 340 0 0 0 Y
flabel comment s 176 314 176 314 0 FreeSans 340 0 0 0 Y
flabel comment s 176 246 176 246 0 FreeSans 340 0 0 0 Y
<< properties >>
string FIXED_BBOX 38 8 314 552
string path 0.950 0.200 7.850 0.200 
<< end >>
