magic
tech sky130B
magscale 1 2
timestamp 1697152928
<< nwell >>
rect -410 -198 1590 -100
rect -410 -202 -237 -198
rect 878 -519 1590 -198
<< nsubdiff >>
rect -199 -166 78 -165
rect -199 -200 -171 -166
rect -137 -200 78 -166
rect -199 -211 78 -200
<< nsubdiffcont >>
rect -171 -200 -137 -166
<< locali >>
rect -196 754 -161 755
rect -162 720 -161 754
rect -196 644 -161 720
rect 36 474 71 651
rect 273 476 308 697
rect 507 476 542 685
rect 742 476 777 685
rect 273 474 777 476
rect 978 474 1013 701
rect 36 439 1318 474
rect 36 216 71 439
rect 273 241 308 439
rect 507 252 542 439
rect 742 236 777 439
rect 978 252 1013 439
rect -200 -166 82 -142
rect -200 -200 -171 -166
rect -137 -200 82 -166
rect -200 -229 82 -200
rect 759 -496 761 -456
rect 795 -496 798 -456
rect 397 -521 560 -520
rect 437 -561 560 -521
rect 759 -616 798 -496
rect 978 -564 1074 -525
rect 1207 -628 1246 -567
<< viali >>
rect -196 720 -162 754
rect 1206 135 1240 169
rect 761 -496 795 -456
rect 397 -561 437 -521
rect 938 -565 978 -525
rect 1206 -567 1246 -527
<< metal1 >>
rect 898 898 950 904
rect -34 852 898 891
rect 950 852 1080 891
rect 898 840 950 846
rect -354 754 -319 759
rect -208 754 -150 760
rect -354 720 -196 754
rect -162 720 -150 754
rect -354 719 -150 720
rect -354 -195 -319 719
rect -208 714 -150 719
rect -85 477 -49 687
rect 150 477 186 719
rect -85 476 186 477
rect 387 476 423 707
rect 622 476 658 722
rect 862 476 898 665
rect 1095 476 1131 668
rect -85 475 1131 476
rect -251 439 1131 475
rect -85 237 -49 439
rect 150 224 186 439
rect 387 141 423 439
rect 622 224 658 439
rect 862 232 898 439
rect 1095 201 1131 439
rect 1423 178 1475 184
rect 1194 169 1252 175
rect 1194 135 1206 169
rect 1240 135 1423 169
rect 1194 134 1423 135
rect 1194 129 1252 134
rect 1475 134 1484 169
rect 1423 120 1475 126
rect 1077 73 1083 80
rect -36 34 1083 73
rect 1077 28 1083 34
rect 1135 28 1141 80
rect 743 -502 749 -450
rect 801 -502 807 -450
rect 385 -567 391 -515
rect 443 -567 449 -515
rect 932 -519 984 -513
rect 932 -577 984 -571
rect 1194 -573 1200 -521
rect 1252 -573 1258 -521
rect 1418 -807 1424 -755
rect 1476 -807 1482 -755
<< via1 >>
rect 898 846 950 898
rect 1423 126 1475 178
rect 1083 28 1135 80
rect 749 -456 801 -450
rect 749 -496 761 -456
rect 761 -496 795 -456
rect 795 -496 801 -456
rect 749 -502 801 -496
rect 391 -521 443 -515
rect 391 -561 397 -521
rect 397 -561 437 -521
rect 437 -561 443 -521
rect 391 -567 443 -561
rect 932 -525 984 -519
rect 932 -565 938 -525
rect 938 -565 978 -525
rect 978 -565 984 -525
rect 932 -571 984 -565
rect 1200 -527 1252 -521
rect 1200 -567 1206 -527
rect 1206 -567 1246 -527
rect 1246 -567 1252 -527
rect 1200 -573 1252 -567
rect 1424 -807 1476 -755
<< metal2 >>
rect 892 846 898 898
rect 950 846 956 898
rect 905 -346 944 846
rect 1417 126 1423 178
rect 1475 126 1481 178
rect 1083 80 1135 86
rect 1135 35 1245 74
rect 1083 22 1135 28
rect 899 -347 944 -346
rect 755 -386 944 -347
rect 755 -444 794 -386
rect 749 -450 801 -444
rect 749 -508 801 -502
rect 391 -515 443 -509
rect 899 -519 938 -386
rect 1206 -515 1245 35
rect 899 -565 932 -519
rect 391 -573 443 -567
rect 926 -571 932 -565
rect 984 -571 990 -519
rect 1200 -521 1252 -515
rect 396 -892 437 -573
rect 1200 -579 1252 -573
rect 1432 -749 1467 126
rect 1424 -755 1476 -749
rect 1424 -813 1476 -807
use sky130_fd_pr__nfet_01v8_JJRV6Y  sky130_fd_pr__nfet_01v8_JJRV6Y_0
timestamp 1696895721
transform 1 0 523 0 -1 179
box -757 -279 757 279
use sky130_fd_pr__pfet_01v8_VVAZD4  sky130_fd_pr__pfet_01v8_VVAZD4_0
timestamp 1696984848
transform 1 0 525 0 1 743
box -757 -284 757 284
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0
timestamp 1693170804
transform 1 0 1275 0 1 -780
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_0
timestamp 1693170804
transform 1 0 -372 0 1 -780
box -38 -48 774 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1693170804
transform 1 0 815 0 1 -780
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_1
timestamp 1693170804
transform 1 0 362 0 1 -780
box -38 -48 498 592
<< labels >>
flabel metal2 905 -369 944 846 0 FreeSans 640 0 0 0 en_buf
flabel locali 1283 439 1318 474 0 FreeSans 640 0 0 0 out
port 0 nsew
flabel metal2 396 -892 437 -567 0 FreeSans 640 0 0 0 en
port 1 nsew
flabel metal1 -251 439 -215 475 0 FreeSans 640 0 0 0 in
port 4 nsew
flabel metal2 1206 -521 1245 74 0 FreeSans 640 0 0 0 net1
flabel metal2 1432 -755 1467 126 0 FreeSans 640 0 0 0 vss
port 2 nsew
flabel metal1 -354 -195 -319 759 0 FreeSans 640 0 0 0 vdd
port 3 nsew
<< end >>
