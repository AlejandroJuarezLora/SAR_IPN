magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect 0 309 260 630
<< pwell >>
rect 41 86 219 243
<< psubdiff >>
rect 67 193 193 217
rect 101 159 159 193
rect 67 112 193 159
<< nsubdiff >>
rect 67 495 193 528
rect 101 461 159 495
rect 67 411 193 461
rect 101 377 159 411
rect 67 353 193 377
<< psubdiffcont >>
rect 67 159 101 193
rect 159 159 193 193
<< nsubdiffcont >>
rect 67 461 101 495
rect 159 461 193 495
rect 67 377 101 411
rect 159 377 193 411
<< locali >>
rect 38 575 67 609
rect 101 575 159 609
rect 193 575 222 609
rect 55 495 205 575
rect 55 461 67 495
rect 101 461 159 495
rect 193 461 205 495
rect 55 411 205 461
rect 55 377 67 411
rect 101 377 159 411
rect 193 377 205 411
rect 55 342 205 377
rect 55 193 205 210
rect 55 159 67 193
rect 101 159 159 193
rect 193 159 205 193
rect 55 65 205 159
rect 38 31 67 65
rect 101 31 159 65
rect 193 31 222 65
<< viali >>
rect 67 575 101 609
rect 159 575 193 609
rect 67 31 101 65
rect 159 31 193 65
<< metal1 >>
rect 38 609 222 640
rect 38 575 67 609
rect 101 575 159 609
rect 193 575 222 609
rect 38 544 222 575
rect 38 65 222 96
rect 38 31 67 65
rect 101 31 159 65
rect 193 31 222 65
rect 38 0 222 31
<< labels >>
rlabel comment s 38 48 38 48 4 tap_2
<< properties >>
string FIXED_BBOX 38 48 222 592
string path 0.950 1.200 5.550 1.200 
<< end >>
