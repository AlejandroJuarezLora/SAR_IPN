magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_p >>
rect -560 105 -502 111
rect -442 105 -384 111
rect -324 105 -266 111
rect -206 105 -148 111
rect -88 105 -30 111
rect 30 105 88 111
rect 148 105 206 111
rect 266 105 324 111
rect 384 105 442 111
rect 502 105 560 111
rect -560 71 -548 105
rect -442 71 -430 105
rect -324 71 -312 105
rect -206 71 -194 105
rect -88 71 -76 105
rect 30 71 42 105
rect 148 71 160 105
rect 266 71 278 105
rect 384 71 396 105
rect 502 71 514 105
rect -560 65 -502 71
rect -442 65 -384 71
rect -324 65 -266 71
rect -206 65 -148 71
rect -88 65 -30 71
rect 30 65 88 71
rect 148 65 206 71
rect 266 65 324 71
rect 384 65 442 71
rect 502 65 560 71
<< nwell >>
rect -757 -324 757 244
<< pmos >>
rect -561 -176 -501 24
rect -443 -176 -383 24
rect -325 -176 -265 24
rect -207 -176 -147 24
rect -89 -176 -29 24
rect 29 -176 89 24
rect 147 -176 207 24
rect 265 -176 325 24
rect 383 -176 443 24
rect 501 -176 561 24
<< pdiff >>
rect -619 9 -561 24
rect -619 -25 -607 9
rect -573 -25 -561 9
rect -619 -59 -561 -25
rect -619 -93 -607 -59
rect -573 -93 -561 -59
rect -619 -127 -561 -93
rect -619 -161 -607 -127
rect -573 -161 -561 -127
rect -619 -176 -561 -161
rect -501 9 -443 24
rect -501 -25 -489 9
rect -455 -25 -443 9
rect -501 -59 -443 -25
rect -501 -93 -489 -59
rect -455 -93 -443 -59
rect -501 -127 -443 -93
rect -501 -161 -489 -127
rect -455 -161 -443 -127
rect -501 -176 -443 -161
rect -383 9 -325 24
rect -383 -25 -371 9
rect -337 -25 -325 9
rect -383 -59 -325 -25
rect -383 -93 -371 -59
rect -337 -93 -325 -59
rect -383 -127 -325 -93
rect -383 -161 -371 -127
rect -337 -161 -325 -127
rect -383 -176 -325 -161
rect -265 9 -207 24
rect -265 -25 -253 9
rect -219 -25 -207 9
rect -265 -59 -207 -25
rect -265 -93 -253 -59
rect -219 -93 -207 -59
rect -265 -127 -207 -93
rect -265 -161 -253 -127
rect -219 -161 -207 -127
rect -265 -176 -207 -161
rect -147 9 -89 24
rect -147 -25 -135 9
rect -101 -25 -89 9
rect -147 -59 -89 -25
rect -147 -93 -135 -59
rect -101 -93 -89 -59
rect -147 -127 -89 -93
rect -147 -161 -135 -127
rect -101 -161 -89 -127
rect -147 -176 -89 -161
rect -29 9 29 24
rect -29 -25 -17 9
rect 17 -25 29 9
rect -29 -59 29 -25
rect -29 -93 -17 -59
rect 17 -93 29 -59
rect -29 -127 29 -93
rect -29 -161 -17 -127
rect 17 -161 29 -127
rect -29 -176 29 -161
rect 89 9 147 24
rect 89 -25 101 9
rect 135 -25 147 9
rect 89 -59 147 -25
rect 89 -93 101 -59
rect 135 -93 147 -59
rect 89 -127 147 -93
rect 89 -161 101 -127
rect 135 -161 147 -127
rect 89 -176 147 -161
rect 207 9 265 24
rect 207 -25 219 9
rect 253 -25 265 9
rect 207 -59 265 -25
rect 207 -93 219 -59
rect 253 -93 265 -59
rect 207 -127 265 -93
rect 207 -161 219 -127
rect 253 -161 265 -127
rect 207 -176 265 -161
rect 325 9 383 24
rect 325 -25 337 9
rect 371 -25 383 9
rect 325 -59 383 -25
rect 325 -93 337 -59
rect 371 -93 383 -59
rect 325 -127 383 -93
rect 325 -161 337 -127
rect 371 -161 383 -127
rect 325 -176 383 -161
rect 443 9 501 24
rect 443 -25 455 9
rect 489 -25 501 9
rect 443 -59 501 -25
rect 443 -93 455 -59
rect 489 -93 501 -59
rect 443 -127 501 -93
rect 443 -161 455 -127
rect 489 -161 501 -127
rect 443 -176 501 -161
rect 561 9 619 24
rect 561 -25 573 9
rect 607 -25 619 9
rect 561 -59 619 -25
rect 561 -93 573 -59
rect 607 -93 619 -59
rect 561 -127 619 -93
rect 561 -161 573 -127
rect 607 -161 619 -127
rect 561 -176 619 -161
<< pdiffc >>
rect -607 -25 -573 9
rect -607 -93 -573 -59
rect -607 -161 -573 -127
rect -489 -25 -455 9
rect -489 -93 -455 -59
rect -489 -161 -455 -127
rect -371 -25 -337 9
rect -371 -93 -337 -59
rect -371 -161 -337 -127
rect -253 -25 -219 9
rect -253 -93 -219 -59
rect -253 -161 -219 -127
rect -135 -25 -101 9
rect -135 -93 -101 -59
rect -135 -161 -101 -127
rect -17 -25 17 9
rect -17 -93 17 -59
rect -17 -161 17 -127
rect 101 -25 135 9
rect 101 -93 135 -59
rect 101 -161 135 -127
rect 219 -25 253 9
rect 219 -93 253 -59
rect 219 -161 253 -127
rect 337 -25 371 9
rect 337 -93 371 -59
rect 337 -161 371 -127
rect 455 -25 489 9
rect 455 -93 489 -59
rect 455 -161 489 -127
rect 573 -25 607 9
rect 573 -93 607 -59
rect 573 -161 607 -127
<< nsubdiff >>
rect -721 174 -595 208
rect -561 174 -527 208
rect -493 174 -459 208
rect -425 174 -391 208
rect -357 174 -323 208
rect -289 174 -255 208
rect -221 174 -187 208
rect -153 174 -119 208
rect -85 174 -51 208
rect -17 174 17 208
rect 51 174 85 208
rect 119 174 153 208
rect 187 174 221 208
rect 255 174 289 208
rect 323 174 357 208
rect 391 174 425 208
rect 459 174 493 208
rect 527 174 561 208
rect 595 174 721 208
rect -721 79 -687 174
rect 687 79 721 174
rect -721 11 -687 45
rect -721 -57 -687 -23
rect -721 -125 -687 -91
rect -721 -254 -687 -159
rect 687 11 721 45
rect 687 -57 721 -23
rect 687 -125 721 -91
rect 687 -254 721 -159
rect -721 -288 -595 -254
rect -561 -288 -527 -254
rect -493 -288 -459 -254
rect -425 -288 -391 -254
rect -357 -288 -323 -254
rect -289 -288 -255 -254
rect -221 -288 -187 -254
rect -153 -288 -119 -254
rect -85 -288 -51 -254
rect -17 -288 17 -254
rect 51 -288 85 -254
rect 119 -288 153 -254
rect 187 -288 221 -254
rect 255 -288 289 -254
rect 323 -288 357 -254
rect 391 -288 425 -254
rect 459 -288 493 -254
rect 527 -288 561 -254
rect 595 -288 721 -254
<< nsubdiffcont >>
rect -595 174 -561 208
rect -527 174 -493 208
rect -459 174 -425 208
rect -391 174 -357 208
rect -323 174 -289 208
rect -255 174 -221 208
rect -187 174 -153 208
rect -119 174 -85 208
rect -51 174 -17 208
rect 17 174 51 208
rect 85 174 119 208
rect 153 174 187 208
rect 221 174 255 208
rect 289 174 323 208
rect 357 174 391 208
rect 425 174 459 208
rect 493 174 527 208
rect 561 174 595 208
rect -721 45 -687 79
rect 687 45 721 79
rect -721 -23 -687 11
rect -721 -91 -687 -57
rect -721 -159 -687 -125
rect 687 -23 721 11
rect 687 -91 721 -57
rect 687 -159 721 -125
rect -595 -288 -561 -254
rect -527 -288 -493 -254
rect -459 -288 -425 -254
rect -391 -288 -357 -254
rect -323 -288 -289 -254
rect -255 -288 -221 -254
rect -187 -288 -153 -254
rect -119 -288 -85 -254
rect -51 -288 -17 -254
rect 17 -288 51 -254
rect 85 -288 119 -254
rect 153 -288 187 -254
rect 221 -288 255 -254
rect 289 -288 323 -254
rect 357 -288 391 -254
rect 425 -288 459 -254
rect 493 -288 527 -254
rect 561 -288 595 -254
<< poly >>
rect -564 105 -498 121
rect -564 71 -548 105
rect -514 71 -498 105
rect -564 55 -498 71
rect -446 105 -380 121
rect -446 71 -430 105
rect -396 71 -380 105
rect -446 55 -380 71
rect -328 105 -262 121
rect -328 71 -312 105
rect -278 71 -262 105
rect -328 55 -262 71
rect -210 105 -144 121
rect -210 71 -194 105
rect -160 71 -144 105
rect -210 55 -144 71
rect -92 105 -26 121
rect -92 71 -76 105
rect -42 71 -26 105
rect -92 55 -26 71
rect 26 105 92 121
rect 26 71 42 105
rect 76 71 92 105
rect 26 55 92 71
rect 144 105 210 121
rect 144 71 160 105
rect 194 71 210 105
rect 144 55 210 71
rect 262 105 328 121
rect 262 71 278 105
rect 312 71 328 105
rect 262 55 328 71
rect 380 105 446 121
rect 380 71 396 105
rect 430 71 446 105
rect 380 55 446 71
rect 498 105 564 121
rect 498 71 514 105
rect 548 71 564 105
rect 498 55 564 71
rect -561 24 -501 55
rect -443 24 -383 55
rect -325 24 -265 55
rect -207 24 -147 55
rect -89 24 -29 55
rect 29 24 89 55
rect 147 24 207 55
rect 265 24 325 55
rect 383 24 443 55
rect 501 24 561 55
rect -561 -202 -501 -176
rect -443 -202 -383 -176
rect -325 -202 -265 -176
rect -207 -202 -147 -176
rect -89 -202 -29 -176
rect 29 -202 89 -176
rect 147 -202 207 -176
rect 265 -202 325 -176
rect 383 -202 443 -176
rect 501 -202 561 -176
<< polycont >>
rect -548 71 -514 105
rect -430 71 -396 105
rect -312 71 -278 105
rect -194 71 -160 105
rect -76 71 -42 105
rect 42 71 76 105
rect 160 71 194 105
rect 278 71 312 105
rect 396 71 430 105
rect 514 71 548 105
<< locali >>
rect -721 174 -595 208
rect -561 174 -527 208
rect -493 174 -459 208
rect -425 174 -391 208
rect -357 174 -323 208
rect -289 174 -255 208
rect -221 174 -187 208
rect -153 174 -119 208
rect -85 174 -51 208
rect -17 174 17 208
rect 51 174 85 208
rect 119 174 153 208
rect 187 174 221 208
rect 255 174 289 208
rect 323 174 357 208
rect 391 174 425 208
rect 459 174 493 208
rect 527 174 561 208
rect 595 174 721 208
rect -721 79 -687 174
rect -564 71 -548 105
rect -514 71 -498 105
rect -446 71 -430 105
rect -396 71 -380 105
rect -328 71 -312 105
rect -278 71 -262 105
rect -210 71 -194 105
rect -160 71 -144 105
rect -92 71 -76 105
rect -42 71 -26 105
rect 26 71 42 105
rect 76 71 92 105
rect 144 71 160 105
rect 194 71 210 105
rect 262 71 278 105
rect 312 71 328 105
rect 380 71 396 105
rect 430 71 446 105
rect 498 71 514 105
rect 548 71 564 105
rect 687 79 721 174
rect -721 11 -687 45
rect -721 -57 -687 -23
rect -721 -125 -687 -91
rect -721 -254 -687 -159
rect -607 9 -573 28
rect -607 -59 -573 -57
rect -607 -95 -573 -93
rect -607 -180 -573 -161
rect -489 9 -455 28
rect -489 -59 -455 -57
rect -489 -95 -455 -93
rect -489 -180 -455 -161
rect -371 9 -337 28
rect -371 -59 -337 -57
rect -371 -95 -337 -93
rect -371 -180 -337 -161
rect -253 9 -219 28
rect -253 -59 -219 -57
rect -253 -95 -219 -93
rect -253 -180 -219 -161
rect -135 9 -101 28
rect -135 -59 -101 -57
rect -135 -95 -101 -93
rect -135 -180 -101 -161
rect -17 9 17 28
rect -17 -59 17 -57
rect -17 -95 17 -93
rect -17 -180 17 -161
rect 101 9 135 28
rect 101 -59 135 -57
rect 101 -95 135 -93
rect 101 -180 135 -161
rect 219 9 253 28
rect 219 -59 253 -57
rect 219 -95 253 -93
rect 219 -180 253 -161
rect 337 9 371 28
rect 337 -59 371 -57
rect 337 -95 371 -93
rect 337 -180 371 -161
rect 455 9 489 28
rect 455 -59 489 -57
rect 455 -95 489 -93
rect 455 -180 489 -161
rect 573 9 607 28
rect 573 -59 607 -57
rect 573 -95 607 -93
rect 573 -180 607 -161
rect 687 11 721 45
rect 687 -57 721 -23
rect 687 -125 721 -91
rect 687 -254 721 -159
rect -721 -288 -595 -254
rect -561 -288 -527 -254
rect -493 -288 -459 -254
rect -425 -288 -391 -254
rect -357 -288 -323 -254
rect -289 -288 -255 -254
rect -221 -288 -187 -254
rect -153 -288 -119 -254
rect -85 -288 -51 -254
rect -17 -288 17 -254
rect 51 -288 85 -254
rect 119 -288 153 -254
rect 187 -288 221 -254
rect 255 -288 289 -254
rect 323 -288 357 -254
rect 391 -288 425 -254
rect 459 -288 493 -254
rect 527 -288 561 -254
rect 595 -288 721 -254
<< viali >>
rect -548 71 -514 105
rect -430 71 -396 105
rect -312 71 -278 105
rect -194 71 -160 105
rect -76 71 -42 105
rect 42 71 76 105
rect 160 71 194 105
rect 278 71 312 105
rect 396 71 430 105
rect 514 71 548 105
rect -607 -25 -573 -23
rect -607 -57 -573 -25
rect -607 -127 -573 -95
rect -607 -129 -573 -127
rect -489 -25 -455 -23
rect -489 -57 -455 -25
rect -489 -127 -455 -95
rect -489 -129 -455 -127
rect -371 -25 -337 -23
rect -371 -57 -337 -25
rect -371 -127 -337 -95
rect -371 -129 -337 -127
rect -253 -25 -219 -23
rect -253 -57 -219 -25
rect -253 -127 -219 -95
rect -253 -129 -219 -127
rect -135 -25 -101 -23
rect -135 -57 -101 -25
rect -135 -127 -101 -95
rect -135 -129 -101 -127
rect -17 -25 17 -23
rect -17 -57 17 -25
rect -17 -127 17 -95
rect -17 -129 17 -127
rect 101 -25 135 -23
rect 101 -57 135 -25
rect 101 -127 135 -95
rect 101 -129 135 -127
rect 219 -25 253 -23
rect 219 -57 253 -25
rect 219 -127 253 -95
rect 219 -129 253 -127
rect 337 -25 371 -23
rect 337 -57 371 -25
rect 337 -127 371 -95
rect 337 -129 371 -127
rect 455 -25 489 -23
rect 455 -57 489 -25
rect 455 -127 489 -95
rect 455 -129 489 -127
rect 573 -25 607 -23
rect 573 -57 607 -25
rect 573 -127 607 -95
rect 573 -129 607 -127
<< metal1 >>
rect -560 105 -502 111
rect -560 71 -548 105
rect -514 71 -502 105
rect -560 65 -502 71
rect -442 105 -384 111
rect -442 71 -430 105
rect -396 71 -384 105
rect -442 65 -384 71
rect -324 105 -266 111
rect -324 71 -312 105
rect -278 71 -266 105
rect -324 65 -266 71
rect -206 105 -148 111
rect -206 71 -194 105
rect -160 71 -148 105
rect -206 65 -148 71
rect -88 105 -30 111
rect -88 71 -76 105
rect -42 71 -30 105
rect -88 65 -30 71
rect 30 105 88 111
rect 30 71 42 105
rect 76 71 88 105
rect 30 65 88 71
rect 148 105 206 111
rect 148 71 160 105
rect 194 71 206 105
rect 148 65 206 71
rect 266 105 324 111
rect 266 71 278 105
rect 312 71 324 105
rect 266 65 324 71
rect 384 105 442 111
rect 384 71 396 105
rect 430 71 442 105
rect 384 65 442 71
rect 502 105 560 111
rect 502 71 514 105
rect 548 71 560 105
rect 502 65 560 71
rect -613 -23 -567 24
rect -613 -57 -607 -23
rect -573 -57 -567 -23
rect -613 -95 -567 -57
rect -613 -129 -607 -95
rect -573 -129 -567 -95
rect -613 -176 -567 -129
rect -495 -23 -449 24
rect -495 -57 -489 -23
rect -455 -57 -449 -23
rect -495 -95 -449 -57
rect -495 -129 -489 -95
rect -455 -129 -449 -95
rect -495 -176 -449 -129
rect -377 -23 -331 24
rect -377 -57 -371 -23
rect -337 -57 -331 -23
rect -377 -95 -331 -57
rect -377 -129 -371 -95
rect -337 -129 -331 -95
rect -377 -176 -331 -129
rect -259 -23 -213 24
rect -259 -57 -253 -23
rect -219 -57 -213 -23
rect -259 -95 -213 -57
rect -259 -129 -253 -95
rect -219 -129 -213 -95
rect -259 -176 -213 -129
rect -141 -23 -95 24
rect -141 -57 -135 -23
rect -101 -57 -95 -23
rect -141 -95 -95 -57
rect -141 -129 -135 -95
rect -101 -129 -95 -95
rect -141 -176 -95 -129
rect -23 -23 23 24
rect -23 -57 -17 -23
rect 17 -57 23 -23
rect -23 -95 23 -57
rect -23 -129 -17 -95
rect 17 -129 23 -95
rect -23 -176 23 -129
rect 95 -23 141 24
rect 95 -57 101 -23
rect 135 -57 141 -23
rect 95 -95 141 -57
rect 95 -129 101 -95
rect 135 -129 141 -95
rect 95 -176 141 -129
rect 213 -23 259 24
rect 213 -57 219 -23
rect 253 -57 259 -23
rect 213 -95 259 -57
rect 213 -129 219 -95
rect 253 -129 259 -95
rect 213 -176 259 -129
rect 331 -23 377 24
rect 331 -57 337 -23
rect 371 -57 377 -23
rect 331 -95 377 -57
rect 331 -129 337 -95
rect 371 -129 377 -95
rect 331 -176 377 -129
rect 449 -23 495 24
rect 449 -57 455 -23
rect 489 -57 495 -23
rect 449 -95 495 -57
rect 449 -129 455 -95
rect 489 -129 495 -95
rect 449 -176 495 -129
rect 567 -23 613 24
rect 567 -57 573 -23
rect 607 -57 613 -23
rect 567 -95 613 -57
rect 567 -129 573 -95
rect 607 -129 613 -95
rect 567 -176 613 -129
<< properties >>
string FIXED_BBOX -704 -271 704 191
<< end >>
