magic
tech sky130B
magscale 1 2
timestamp 1696111957
<< metal1 >>
rect 1376 1286 3106 1314
rect 1380 490 3110 518
rect 2180 242 2208 490
rect 2314 164 2372 224
rect 2150 124 2220 144
use sky130_fd_pr__nfet_01v8_lvt_E33R59  sky130_fd_pr__nfet_01v8_lvt_E33R59_0
timestamp 1696108744
transform 0 1 2219 -1 0 194
box -226 -279 226 279
use trimcap  trimcap_0
timestamp 1696109480
transform 1 0 1140 0 1 60
box 0 376 476 1324
use trimcap  trimcap_1
timestamp 1696109480
transform 1 0 2852 0 1 66
box 0 376 476 1324
use trimcap  trimcap_2
timestamp 1696109480
transform 1 0 1710 0 1 60
box 0 376 476 1324
use trimcap  trimcap_3
timestamp 1696109480
transform 1 0 2280 0 1 64
box 0 376 476 1324
<< labels >>
flabel metal1 1376 1286 3106 1314 0 FreeSans 800 0 0 0 todrain
flabel metal1 2314 164 2372 224 0 FreeSans 800 0 0 0 d_i
flabel metal1 2150 124 2220 144 0 FreeSans 480 0 0 0 tovss
<< end >>
