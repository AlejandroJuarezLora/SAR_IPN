magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 1050 542
<< pwell >>
rect 1 27 1010 163
rect 29 -19 1010 27
rect 29 -57 63 -19
<< scnmos >>
rect 79 53 109 137
rect 267 7 297 137
rect 373 7 403 137
rect 457 7 487 137
rect 541 7 571 137
rect 647 7 677 137
rect 731 7 761 137
rect 815 7 845 137
rect 899 7 929 137
<< scpmoshvt >>
rect 79 373 109 457
rect 267 257 297 457
rect 373 257 403 457
rect 457 257 487 457
rect 541 257 571 457
rect 647 257 677 457
rect 731 257 761 457
rect 815 257 845 457
rect 899 257 929 457
<< ndiff >>
rect 27 109 79 137
rect 27 75 35 109
rect 69 75 79 109
rect 27 53 79 75
rect 109 125 161 137
rect 109 91 119 125
rect 153 91 161 125
rect 109 80 161 91
rect 109 53 159 80
rect 217 64 267 137
rect 215 53 267 64
rect 215 19 223 53
rect 257 19 267 53
rect 215 7 267 19
rect 297 75 373 137
rect 297 41 323 75
rect 357 41 373 75
rect 297 7 373 41
rect 403 57 457 137
rect 403 23 413 57
rect 447 23 457 57
rect 403 7 457 23
rect 487 75 541 137
rect 487 41 497 75
rect 531 41 541 75
rect 487 7 541 41
rect 571 57 647 137
rect 571 23 601 57
rect 635 23 647 57
rect 571 7 647 23
rect 677 74 731 137
rect 677 40 687 74
rect 721 40 731 74
rect 677 7 731 40
rect 761 55 815 137
rect 761 21 771 55
rect 805 21 815 55
rect 761 7 815 21
rect 845 123 899 137
rect 845 89 855 123
rect 889 89 899 123
rect 845 55 899 89
rect 845 21 855 55
rect 889 21 899 55
rect 845 7 899 21
rect 929 55 984 137
rect 929 21 939 55
rect 973 21 984 55
rect 929 7 984 21
<< pdiff >>
rect 27 437 79 457
rect 27 403 35 437
rect 69 403 79 437
rect 27 373 79 403
rect 109 432 161 457
rect 109 398 119 432
rect 153 398 161 432
rect 109 373 161 398
rect 215 445 267 457
rect 215 411 223 445
rect 257 411 267 445
rect 215 377 267 411
rect 215 343 223 377
rect 257 343 267 377
rect 215 309 267 343
rect 215 275 223 309
rect 257 275 267 309
rect 215 257 267 275
rect 297 257 373 457
rect 403 257 457 457
rect 487 257 541 457
rect 571 437 647 457
rect 571 403 592 437
rect 626 403 647 437
rect 571 369 647 403
rect 571 335 592 369
rect 626 335 647 369
rect 571 257 647 335
rect 677 437 731 457
rect 677 403 687 437
rect 721 403 731 437
rect 677 369 731 403
rect 677 335 687 369
rect 721 335 731 369
rect 677 301 731 335
rect 677 267 687 301
rect 721 267 731 301
rect 677 257 731 267
rect 761 437 815 457
rect 761 403 771 437
rect 805 403 815 437
rect 761 369 815 403
rect 761 335 771 369
rect 805 335 815 369
rect 761 257 815 335
rect 845 437 899 457
rect 845 403 855 437
rect 889 403 899 437
rect 845 369 899 403
rect 845 335 855 369
rect 889 335 899 369
rect 845 301 899 335
rect 845 267 855 301
rect 889 267 899 301
rect 845 257 899 267
rect 929 437 981 457
rect 929 403 939 437
rect 973 403 981 437
rect 929 369 981 403
rect 929 335 939 369
rect 973 335 981 369
rect 929 257 981 335
<< ndiffc >>
rect 35 75 69 109
rect 119 91 153 125
rect 223 19 257 53
rect 323 41 357 75
rect 413 23 447 57
rect 497 41 531 75
rect 601 23 635 57
rect 687 40 721 74
rect 771 21 805 55
rect 855 89 889 123
rect 855 21 889 55
rect 939 21 973 55
<< pdiffc >>
rect 35 403 69 437
rect 119 398 153 432
rect 223 411 257 445
rect 223 343 257 377
rect 223 275 257 309
rect 592 403 626 437
rect 592 335 626 369
rect 687 403 721 437
rect 687 335 721 369
rect 687 267 721 301
rect 771 403 805 437
rect 771 335 805 369
rect 855 403 889 437
rect 855 335 889 369
rect 855 267 889 301
rect 939 403 973 437
rect 939 335 973 369
<< poly >>
rect 79 457 109 483
rect 267 457 297 483
rect 373 457 403 483
rect 457 457 487 483
rect 541 457 571 483
rect 647 457 677 483
rect 731 457 761 483
rect 815 457 845 483
rect 899 457 929 483
rect 79 225 109 373
rect 267 225 297 257
rect 373 225 403 257
rect 457 225 487 257
rect 541 225 571 257
rect 647 225 677 257
rect 731 225 761 257
rect 815 225 845 257
rect 899 225 929 257
rect 45 209 113 225
rect 45 175 55 209
rect 89 175 113 209
rect 45 159 113 175
rect 199 209 297 225
rect 199 175 209 209
rect 243 175 297 209
rect 199 159 297 175
rect 349 209 403 225
rect 349 175 359 209
rect 393 175 403 209
rect 349 159 403 175
rect 445 209 499 225
rect 445 175 455 209
rect 489 175 499 209
rect 445 159 499 175
rect 541 209 595 225
rect 541 175 551 209
rect 585 175 595 209
rect 541 159 595 175
rect 647 209 929 225
rect 647 175 657 209
rect 691 175 725 209
rect 759 175 793 209
rect 827 175 861 209
rect 895 175 929 209
rect 647 159 929 175
rect 79 137 109 159
rect 267 137 297 159
rect 373 137 403 159
rect 457 137 487 159
rect 541 137 571 159
rect 647 137 677 159
rect 731 137 761 159
rect 815 137 845 159
rect 899 137 929 159
rect 79 27 109 53
rect 267 -19 297 7
rect 373 -19 403 7
rect 457 -19 487 7
rect 541 -19 571 7
rect 647 -19 677 7
rect 731 -19 761 7
rect 815 -19 845 7
rect 899 -19 929 7
<< polycont >>
rect 55 175 89 209
rect 209 175 243 209
rect 359 175 393 209
rect 455 175 489 209
rect 551 175 585 209
rect 657 175 691 209
rect 725 175 759 209
rect 793 175 827 209
rect 861 175 895 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1012 521
rect 17 437 73 487
rect 17 403 35 437
rect 69 403 73 437
rect 17 387 73 403
rect 119 432 157 451
rect 153 398 157 432
rect 119 373 157 398
rect 21 209 89 351
rect 21 175 55 209
rect 21 159 89 175
rect 123 225 157 373
rect 207 445 273 450
rect 207 411 223 445
rect 257 411 273 445
rect 584 437 634 487
rect 207 377 273 411
rect 207 343 223 377
rect 257 343 273 377
rect 207 309 273 343
rect 207 275 223 309
rect 257 275 325 309
rect 123 209 243 225
rect 123 175 209 209
rect 123 159 243 175
rect 123 141 157 159
rect 119 125 157 141
rect 17 109 69 125
rect 17 75 35 109
rect 17 -23 69 75
rect 153 91 157 125
rect 291 125 325 275
rect 359 284 431 435
rect 467 317 527 435
rect 584 403 592 437
rect 626 403 634 437
rect 584 369 634 403
rect 584 335 592 369
rect 626 335 634 369
rect 584 319 634 335
rect 679 437 729 453
rect 679 403 687 437
rect 721 403 729 437
rect 679 369 729 403
rect 679 335 687 369
rect 721 335 729 369
rect 359 209 393 284
rect 467 250 505 317
rect 679 301 729 335
rect 763 437 813 487
rect 763 403 771 437
rect 805 403 813 437
rect 763 369 813 403
rect 763 335 771 369
rect 805 335 813 369
rect 763 319 813 335
rect 847 437 897 453
rect 847 403 855 437
rect 889 403 897 437
rect 847 369 897 403
rect 847 335 855 369
rect 889 335 897 369
rect 359 159 393 175
rect 439 209 505 250
rect 439 175 455 209
rect 489 175 505 209
rect 439 159 505 175
rect 551 249 638 283
rect 679 267 687 301
rect 721 285 729 301
rect 847 301 897 335
rect 931 437 981 487
rect 931 403 939 437
rect 973 403 981 437
rect 931 369 981 403
rect 931 335 939 369
rect 973 335 981 369
rect 931 319 981 335
rect 847 285 855 301
rect 721 267 855 285
rect 889 285 897 301
rect 889 267 993 285
rect 679 251 993 267
rect 551 209 585 249
rect 551 159 585 175
rect 619 175 657 209
rect 691 175 725 209
rect 759 175 793 209
rect 827 175 861 209
rect 895 175 911 209
rect 619 125 653 175
rect 945 141 993 251
rect 291 91 653 125
rect 687 123 993 141
rect 687 105 855 123
rect 119 47 157 91
rect 207 53 257 77
rect 207 19 223 53
rect 323 75 357 91
rect 497 75 531 91
rect 323 21 357 41
rect 397 23 413 57
rect 447 23 463 57
rect 207 -23 257 19
rect 397 -23 463 23
rect 687 74 737 105
rect 497 21 531 41
rect 575 23 601 57
rect 635 23 651 57
rect 575 -23 651 23
rect 721 40 737 74
rect 839 89 855 105
rect 889 105 993 123
rect 889 89 905 105
rect 687 11 737 40
rect 771 55 805 71
rect 771 -23 805 21
rect 839 55 905 89
rect 839 21 855 55
rect 889 21 905 55
rect 839 11 905 21
rect 939 55 973 71
rect 939 -23 973 21
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1012 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 857 487 891 521
rect 949 487 983 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
rect 857 -57 891 -23
rect 949 -57 983 -23
<< metal1 >>
rect 0 521 1012 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1012 521
rect 0 456 1012 487
rect 0 -23 1012 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1012 -23
rect 0 -88 1012 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 or4b_4
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 29 181 63 215 0 FreeSans 400 0 0 0 D_N
port 8 nsew
flabel locali s 489 385 523 419 0 FreeSans 400 0 0 0 B
port 10 nsew
flabel locali s 489 317 523 351 0 FreeSans 400 0 0 0 B
port 10 nsew
flabel locali s 397 317 431 351 0 FreeSans 400 0 0 0 C
port 9 nsew
flabel locali s 581 249 615 283 0 FreeSans 400 0 0 0 A
port 11 nsew
flabel locali s 397 385 431 419 0 FreeSans 400 0 0 0 C
port 9 nsew
flabel locali s 949 113 983 147 0 FreeSans 400 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 1012 504
string path 0.000 -1.000 25.300 -1.000 
<< end >>
