magic
tech sky130B
magscale 1 2
timestamp 1696034456
<< nwell >>
rect 1992 -2 2354 366
rect 2608 -3 2970 365
rect 3226 0 3588 368
<< pmos >>
rect 2092 92 2292 152
rect 2670 91 2870 151
rect 3288 94 3488 154
<< pdiff >>
rect 2092 198 2292 210
rect 2092 164 2104 198
rect 2280 164 2292 198
rect 2092 152 2292 164
rect 2670 197 2870 209
rect 2670 163 2682 197
rect 2858 163 2870 197
rect 2670 151 2870 163
rect 3288 200 3488 212
rect 3288 166 3300 200
rect 3476 166 3488 200
rect 3288 154 3488 166
rect 2092 80 2292 92
rect 2092 46 2104 80
rect 2280 46 2292 80
rect 2092 34 2292 46
rect 2670 79 2870 91
rect 2670 45 2682 79
rect 2858 45 2870 79
rect 2670 33 2870 45
rect 3288 82 3488 94
rect 3288 48 3300 82
rect 3476 48 3488 82
rect 3288 36 3488 48
<< pdiffc >>
rect 2104 164 2280 198
rect 2682 163 2858 197
rect 3300 166 3476 200
rect 2104 46 2280 80
rect 2682 45 2858 79
rect 3300 48 3476 82
<< nsubdiff >>
rect 2092 312 2292 324
rect 2092 278 2131 312
rect 2253 278 2292 312
rect 2092 267 2292 278
rect 2670 311 2870 323
rect 2670 277 2709 311
rect 2831 277 2870 311
rect 2670 266 2870 277
rect 3288 314 3488 326
rect 3288 280 3327 314
rect 3449 280 3488 314
rect 3288 269 3488 280
<< nsubdiffcont >>
rect 2131 278 2253 312
rect 2709 277 2831 311
rect 3327 280 3449 314
<< poly >>
rect 1995 152 2061 155
rect 1995 139 2092 152
rect 1995 105 2011 139
rect 2045 105 2092 139
rect 1995 92 2092 105
rect 2292 92 2318 152
rect 3519 154 3585 157
rect 2901 151 2967 154
rect 1995 89 2061 92
rect 2644 91 2670 151
rect 2870 138 2967 151
rect 2870 104 2917 138
rect 2951 104 2967 138
rect 2870 91 2967 104
rect 3262 94 3288 154
rect 3488 141 3585 154
rect 3488 107 3535 141
rect 3569 107 3585 141
rect 3488 94 3585 107
rect 2901 88 2967 91
rect 3519 91 3585 94
<< polycont >>
rect 2011 105 2045 139
rect 2917 104 2951 138
rect 3535 107 3569 141
<< locali >>
rect 2088 278 2104 312
rect 2280 278 2296 312
rect 2666 277 2682 311
rect 2858 277 2874 311
rect 3284 280 3300 314
rect 3476 280 3492 314
rect 2088 164 2104 198
rect 2280 164 2296 198
rect 2666 163 2682 197
rect 2858 163 2874 197
rect 3284 166 3300 200
rect 3476 166 3492 200
rect 2011 139 2045 155
rect 2011 89 2045 105
rect 2917 138 2951 154
rect 2917 88 2951 104
rect 3535 141 3569 157
rect 3535 91 3569 107
rect 2088 46 2104 80
rect 2280 46 2296 80
rect 2666 45 2682 79
rect 2858 45 2874 79
rect 3284 48 3300 82
rect 3476 48 3492 82
<< viali >>
rect 2104 278 2131 312
rect 2131 278 2253 312
rect 2253 278 2280 312
rect 2682 277 2709 311
rect 2709 277 2831 311
rect 2831 277 2858 311
rect 3300 280 3327 314
rect 3327 280 3449 314
rect 3449 280 3476 314
rect 2104 164 2280 198
rect 2682 163 2858 197
rect 3300 166 3476 200
rect 2011 105 2045 139
rect 2917 104 2951 138
rect 3535 107 3569 141
rect 2104 46 2280 80
rect 2682 45 2858 79
rect 3300 48 3476 82
<< metal1 >>
rect 1099 572 1127 623
rect 1081 520 1087 572
rect 1139 520 1145 572
rect 2461 568 2489 624
rect 2443 516 2449 568
rect 2501 516 2507 568
rect -635 146 -605 485
rect -46 395 3644 423
rect 192 185 220 395
rect 804 180 832 395
rect 1087 206 1139 212
rect 1396 177 1424 395
rect 2174 318 2202 395
rect 2092 312 2292 318
rect 2766 317 2794 395
rect 3378 320 3406 395
rect 2092 278 2104 312
rect 2280 278 2292 312
rect 2092 272 2292 278
rect 2670 311 2870 317
rect 2670 277 2682 311
rect 2858 277 2870 311
rect 2174 230 2202 272
rect 2670 271 2870 277
rect 3288 314 3488 320
rect 3288 280 3300 314
rect 3476 280 3488 314
rect 3288 274 3488 280
rect 2116 204 2202 230
rect 2449 206 2501 212
rect 2092 198 2292 204
rect 2092 164 2104 198
rect 2280 164 2292 198
rect 2092 158 2292 164
rect -646 140 -594 146
rect -646 82 -594 88
rect 18 144 78 150
rect -635 78 -605 82
rect 18 78 78 84
rect 636 144 696 150
rect 1087 148 1139 154
rect 636 78 696 84
rect -635 -172 -605 -142
rect 191 -165 221 76
rect 802 9 831 63
rect 1099 9 1127 148
rect 1998 139 2058 152
rect 1998 137 2011 139
rect 1566 108 1701 136
rect 1462 60 1490 71
rect 1450 40 1502 60
rect 1441 34 1506 40
rect 1441 22 1507 34
rect 1441 9 1447 22
rect 802 -19 1447 9
rect 1441 -30 1447 -19
rect 1501 -30 1507 22
rect 1441 -36 1507 -30
rect 1462 -103 1490 -36
rect 1673 -47 1701 108
rect 1869 109 2011 137
rect 1869 64 1897 109
rect 1998 105 2011 109
rect 2045 105 2058 139
rect 1998 92 2058 105
rect 2116 86 2176 158
rect 2766 203 2794 271
rect 3378 206 3406 274
rect 2670 197 2870 203
rect 2670 163 2682 197
rect 2858 163 2870 197
rect 2670 157 2870 163
rect 3288 200 3488 206
rect 3288 166 3300 200
rect 3476 166 3488 200
rect 3288 160 3488 166
rect 2449 148 2501 154
rect 2904 150 2964 151
rect 2092 80 2292 86
rect 1844 52 1920 64
rect 1844 -1 1857 52
rect 1909 -1 1920 52
rect 2092 46 2104 80
rect 2280 46 2292 80
rect 2092 40 2292 46
rect 1844 -12 1920 -1
rect 2102 9 2130 40
rect 2461 9 2489 148
rect 2902 144 2964 150
rect 2670 79 2870 85
rect 2670 45 2682 79
rect 2858 45 2870 79
rect 2962 91 2964 144
rect 3522 150 3582 154
rect 3522 144 3586 150
rect 3522 94 3526 144
rect 2902 78 2962 84
rect 3288 82 3488 88
rect 2670 39 2870 45
rect 3288 48 3300 82
rect 3476 48 3488 82
rect 3526 78 3586 84
rect 3288 42 3488 48
rect 2710 9 2738 39
rect 1673 -58 1749 -47
rect 1079 -136 1259 -106
rect 1229 -203 1259 -136
rect 1673 -112 1685 -58
rect 1738 -112 1749 -58
rect 1673 -123 1749 -112
rect 1673 -143 1701 -123
rect 1576 -171 1701 -143
rect 1869 -145 1897 -12
rect 2102 -14 2748 9
rect 2102 -67 2115 -14
rect 2167 -19 2748 -14
rect 2167 -67 2179 -19
rect 2102 -79 2179 -67
rect 2102 -98 2130 -79
rect 1869 -173 2022 -145
rect 2477 -172 2656 -142
rect 3375 -164 3405 42
rect 1869 -174 1897 -173
rect 1229 -232 1398 -203
rect 2477 -206 2507 -172
rect 1434 -232 1465 -211
rect 1229 -411 1259 -232
rect 1434 -240 1435 -232
rect 2219 -234 2507 -206
rect 2313 -236 2507 -234
rect 1504 -347 2181 -319
rect 1229 -440 1454 -411
rect 1763 -440 1792 -347
rect 2313 -400 2342 -236
rect 2133 -428 2342 -400
rect 1229 -442 1259 -440
rect 1426 -479 1454 -440
rect 1738 -450 1814 -440
rect 1738 -504 1749 -450
rect 1801 -504 1814 -450
rect 2133 -477 2161 -428
rect 2313 -429 2342 -428
rect 1738 -516 1814 -504
rect 1560 -616 2034 -588
rect 1647 -690 1726 -678
rect 1647 -701 1661 -690
rect 1576 -731 1661 -701
rect 1647 -743 1661 -731
rect 1713 -704 1726 -690
rect 1777 -704 1805 -616
rect 1864 -687 1943 -677
rect 1864 -704 1881 -687
rect 1713 -736 1881 -704
rect 1713 -743 1726 -736
rect 1647 -757 1726 -743
rect 1777 -827 1805 -736
rect 1864 -740 1881 -736
rect 1933 -699 1943 -687
rect 1933 -729 2021 -699
rect 1933 -740 1943 -729
rect 1864 -756 1943 -740
rect 1570 -855 2044 -827
rect 1478 -1087 1511 -939
rect 1738 -1050 1819 -1036
rect 1738 -1061 1751 -1050
rect 1571 -1089 1751 -1061
rect 1680 -1090 1708 -1089
rect 1738 -1104 1751 -1089
rect 1808 -1061 1819 -1050
rect 1808 -1089 2045 -1061
rect 1808 -1104 1851 -1089
rect 2052 -1090 2085 -942
rect 1738 -1115 1851 -1104
rect 1821 -5061 1851 -1115
rect 1108 -5091 2590 -5061
rect -218 -5406 -196 -5386
rect -679 -5440 -650 -5418
rect -550 -5439 -521 -5417
rect -450 -5435 -421 -5413
rect -335 -5437 -306 -5415
rect -218 -5418 -190 -5406
rect -218 -5429 -186 -5418
rect -215 -5440 -186 -5429
rect 1818 -5459 1848 -5091
rect 3923 -5437 3953 -5417
rect 4043 -5436 4073 -5416
rect 4151 -5437 4181 -5417
rect 4265 -5435 4295 -5415
rect 4382 -5438 4412 -5418
<< via1 >>
rect 1087 520 1139 572
rect 2449 516 2501 568
rect 1087 154 1139 206
rect -646 88 -594 140
rect 18 84 78 144
rect 636 84 696 144
rect 1447 -30 1501 22
rect 2449 154 2501 206
rect 1857 -1 1909 52
rect 2902 138 2962 144
rect 2902 104 2917 138
rect 2917 104 2951 138
rect 2951 104 2962 138
rect 2902 84 2962 104
rect 3526 141 3586 144
rect 3526 107 3535 141
rect 3535 107 3569 141
rect 3569 107 3586 141
rect 3526 84 3586 107
rect 1685 -112 1738 -58
rect 2115 -67 2167 -14
rect 1749 -504 1801 -450
rect 1661 -743 1713 -690
rect 1881 -740 1933 -687
rect 1751 -1104 1808 -1050
<< metal2 >>
rect 1087 572 1139 578
rect 1087 514 1139 520
rect 2449 568 2501 574
rect 1099 206 1127 514
rect 2449 510 2501 516
rect 2461 206 2489 510
rect 1081 154 1087 206
rect 1139 154 1145 206
rect 2443 154 2449 206
rect 2501 154 2507 206
rect 20 144 76 151
rect 638 144 694 151
rect 2904 144 2960 151
rect 3528 144 3584 151
rect -659 84 -650 144
rect -590 84 -581 144
rect 12 84 18 144
rect 78 84 84 144
rect 630 84 636 144
rect 696 84 702 144
rect 2896 84 2902 144
rect 2962 84 2968 144
rect 3520 84 3526 144
rect 3586 84 3592 144
rect 20 77 76 84
rect 638 77 694 84
rect 2904 77 2960 84
rect 3528 77 3584 84
rect 1844 52 1920 64
rect 1441 22 1507 34
rect 1441 -30 1447 22
rect 1501 16 1507 22
rect 1844 16 1857 52
rect 1501 -1 1857 16
rect 1909 -1 1920 52
rect 1501 -12 1920 -1
rect 1501 -30 1507 -12
rect 1441 -36 1507 -30
rect 2102 -14 2179 -3
rect 2102 -47 2115 -14
rect 1673 -58 2115 -47
rect 1673 -112 1685 -58
rect 1738 -67 2115 -58
rect 2167 -67 2179 -14
rect 1738 -75 2179 -67
rect 1738 -112 1749 -75
rect 2102 -79 2179 -75
rect 1673 -123 1749 -112
rect 1738 -450 1814 -440
rect 1738 -504 1749 -450
rect 1801 -504 1814 -450
rect 1738 -516 1814 -504
rect 1647 -690 1726 -678
rect 1647 -743 1661 -690
rect 1713 -704 1726 -690
rect 1764 -704 1797 -516
rect 1864 -687 1943 -677
rect 1864 -704 1881 -687
rect 1713 -736 1881 -704
rect 1713 -743 1726 -736
rect 1647 -757 1726 -743
rect 1764 -904 1797 -736
rect 1864 -740 1881 -736
rect 1933 -740 1943 -687
rect 1864 -756 1943 -740
rect 1763 -1036 1797 -904
rect 1738 -1050 1819 -1036
rect 1738 -1104 1751 -1050
rect 1808 -1104 1819 -1050
rect 1738 -1115 1819 -1104
<< via2 >>
rect -650 140 -590 144
rect -650 88 -646 140
rect -646 88 -594 140
rect -594 88 -590 140
rect -650 84 -590 88
rect 20 86 76 142
rect 638 86 694 142
rect 2904 86 2960 142
rect 3528 86 3584 142
<< metal3 >>
rect -655 144 -585 149
rect 15 144 81 147
rect 633 144 699 147
rect 2899 144 2965 147
rect 3523 144 3589 147
rect -655 84 -650 144
rect -590 142 3598 144
rect -590 86 20 142
rect 76 86 638 142
rect 694 86 2904 142
rect 2960 86 3528 142
rect 3584 86 3598 142
rect -590 84 3598 86
rect -655 79 -585 84
rect 15 81 81 84
rect 633 81 699 84
rect 2899 81 2965 84
rect 3523 81 3589 84
use sky130_fd_pr__nfet_01v8_96AECY  sky130_fd_pr__nfet_01v8_96AECY_0
timestamp 1695862321
transform 0 1 1455 1 0 -158
box -200 -157 88 157
use sky130_fd_pr__nfet_01v8_96AECY  sky130_fd_pr__nfet_01v8_96AECY_1
timestamp 1695862321
transform 0 1 2110 1 0 -541
box -200 -157 88 157
use sky130_fd_pr__nfet_01v8_96AECY  sky130_fd_pr__nfet_01v8_96AECY_2
timestamp 1695862321
transform 0 -1 2150 1 0 -161
box -200 -157 88 157
use sky130_fd_pr__nfet_01v8_96AECY  sky130_fd_pr__nfet_01v8_96AECY_3
timestamp 1695862321
transform 0 -1 1477 1 0 -545
box -200 -157 88 157
use sky130_fd_pr__nfet_01v8_96AECY  sky130_fd_pr__nfet_01v8_96AECY_4
timestamp 1695862321
transform 0 1 2108 1 0 -902
box -200 -157 88 157
use sky130_fd_pr__nfet_01v8_96AECY  sky130_fd_pr__nfet_01v8_96AECY_5
timestamp 1695862321
transform 0 -1 1476 1 0 -900
box -200 -157 88 157
use sky130_fd_pr__pfet_01v8_7G6J3C  sky130_fd_pr__pfet_01v8_7G6J3C_0
timestamp 1695925836
transform 0 -1 174 -1 0 124
box -244 -198 124 164
use sky130_fd_pr__pfet_01v8_7G6J3C  sky130_fd_pr__pfet_01v8_7G6J3C_1
timestamp 1695925836
transform 0 1 1442 -1 0 122
box -244 -198 124 164
use sky130_fd_pr__pfet_01v8_7G6J3C  sky130_fd_pr__pfet_01v8_7G6J3C_2
timestamp 1695925836
transform 0 -1 792 -1 0 121
box -244 -198 124 164
use trim  trim_0
timestamp 1696032376
transform 0 1 -1972 -1 0 -127
box -10 60 5302 3118
use trim  trim_1
timestamp 1696032376
transform 0 -1 5707 -1 0 -126
box -10 60 5302 3118
<< labels >>
rlabel viali 2766 291 2766 291 5 B
rlabel polycont 2936 121 2936 121 5 G
rlabel viali 2766 181 2766 181 5 S
rlabel viali 2766 61 2766 61 5 D
rlabel viali 2196 292 2196 292 5 B
rlabel viali 2026 122 2026 122 5 G
rlabel viali 2196 182 2196 182 5 S
rlabel viali 2196 62 2196 62 5 D
rlabel viali 3384 294 3384 294 5 B
rlabel polycont 3554 124 3554 124 5 G
rlabel viali 3384 184 3384 184 5 S
rlabel viali 3384 64 3384 64 5 D
rlabel metal1 1230 -137 1258 -106 1 IN
rlabel metal1 2477 -173 2507 -143 1 IP
rlabel metal1 -46 395 3644 423 1 vdd
port 1 n
rlabel metal1 1821 -5091 1851 -1061 5 vss
port 2 s
rlabel metal1 -201 -5440 -201 -5438 5 trim0
port 4 s
rlabel metal1 -320 -5437 -319 -5436 5 trim1
port 5 s
rlabel metal1 -436 -5435 -435 -5434 5 trim2
port 6 s
rlabel metal1 -537 -5437 -536 -5436 5 trim3
port 7 s
rlabel metal1 -664 -5437 -663 -5436 5 trim4
port 8 s
rlabel metal1 3938 -5435 3938 -5435 5 trimb0
port 9 s
rlabel metal1 4059 -5434 4059 -5434 5 trimb1
port 10 s
rlabel metal1 4165 -5435 4165 -5435 5 trimb2
port 11 s
rlabel metal1 4280 -5434 4280 -5434 5 trimb3
port 12 s
rlabel metal1 4396 -5436 4396 -5436 5 trimb4
port 13 s
rlabel metal1 1099 595 1127 623 1 outn
rlabel metal1 2461 596 2489 624 1 outp
rlabel metal1 -620 476 -620 476 1 clk
port 3 n
<< end >>
