magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 866 542
<< pwell >>
rect 1 -19 827 163
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 109 137
rect 276 7 306 137
rect 379 7 409 137
rect 482 7 512 137
rect 634 7 664 137
rect 718 7 748 137
<< scpmoshvt >>
rect 79 257 109 457
rect 262 257 292 457
rect 379 257 409 457
rect 531 257 561 457
rect 646 257 676 457
rect 718 257 748 457
<< ndiff >>
rect 27 61 79 137
rect 27 27 35 61
rect 69 27 79 61
rect 27 7 79 27
rect 109 53 161 137
rect 109 19 119 53
rect 153 19 161 53
rect 109 7 161 19
rect 215 121 276 137
rect 215 87 223 121
rect 257 87 276 121
rect 215 53 276 87
rect 215 19 223 53
rect 257 19 276 53
rect 215 7 276 19
rect 306 7 379 137
rect 409 7 482 137
rect 512 129 634 137
rect 512 95 590 129
rect 624 95 634 129
rect 512 61 634 95
rect 512 27 590 61
rect 624 27 634 61
rect 512 7 634 27
rect 664 51 718 137
rect 664 17 674 51
rect 708 17 718 51
rect 664 7 718 17
rect 748 61 801 137
rect 748 27 758 61
rect 792 27 801 61
rect 748 7 801 27
<< pdiff >>
rect 27 437 79 457
rect 27 403 35 437
rect 69 403 79 437
rect 27 369 79 403
rect 27 335 35 369
rect 69 335 79 369
rect 27 257 79 335
rect 109 445 262 457
rect 109 411 121 445
rect 155 411 217 445
rect 251 411 262 445
rect 109 377 262 411
rect 109 343 121 377
rect 155 343 217 377
rect 251 343 262 377
rect 109 257 262 343
rect 292 437 379 457
rect 292 403 317 437
rect 351 403 379 437
rect 292 369 379 403
rect 292 335 317 369
rect 351 335 379 369
rect 292 257 379 335
rect 409 445 531 457
rect 409 343 419 445
rect 521 343 531 445
rect 409 257 531 343
rect 561 437 646 457
rect 561 403 602 437
rect 636 403 646 437
rect 561 309 646 403
rect 561 275 602 309
rect 636 275 646 309
rect 561 257 646 275
rect 676 257 718 457
rect 748 445 801 457
rect 748 411 758 445
rect 792 411 801 445
rect 748 377 801 411
rect 748 343 758 377
rect 792 343 801 377
rect 748 257 801 343
<< ndiffc >>
rect 35 27 69 61
rect 119 19 153 53
rect 223 87 257 121
rect 223 19 257 53
rect 590 95 624 129
rect 590 27 624 61
rect 674 17 708 51
rect 758 27 792 61
<< pdiffc >>
rect 35 403 69 437
rect 35 335 69 369
rect 121 411 155 445
rect 217 411 251 445
rect 121 343 155 377
rect 217 343 251 377
rect 317 403 351 437
rect 317 335 351 369
rect 419 343 521 445
rect 602 403 636 437
rect 602 275 636 309
rect 758 411 792 445
rect 758 343 792 377
<< poly >>
rect 79 457 109 483
rect 262 457 292 483
rect 379 457 409 483
rect 531 457 561 483
rect 646 457 676 483
rect 718 457 748 483
rect 79 225 109 257
rect 79 209 149 225
rect 262 219 292 257
rect 379 219 409 257
rect 531 219 561 257
rect 646 219 676 257
rect 79 175 105 209
rect 139 175 149 209
rect 79 159 149 175
rect 253 209 319 219
rect 253 175 269 209
rect 303 175 319 209
rect 253 165 319 175
rect 373 209 439 219
rect 373 175 389 209
rect 423 175 439 209
rect 373 165 439 175
rect 482 209 561 219
rect 482 175 507 209
rect 541 175 561 209
rect 482 165 561 175
rect 610 209 676 219
rect 610 175 626 209
rect 660 175 676 209
rect 610 165 676 175
rect 718 221 748 257
rect 718 209 807 221
rect 718 175 757 209
rect 791 175 807 209
rect 79 137 109 159
rect 276 137 306 165
rect 379 137 409 165
rect 482 137 512 165
rect 634 137 664 165
rect 718 163 807 175
rect 718 137 748 163
rect 79 -19 109 7
rect 276 -19 306 7
rect 379 -19 409 7
rect 482 -19 512 7
rect 634 -19 664 7
rect 718 -19 748 7
<< polycont >>
rect 105 175 139 209
rect 269 175 303 209
rect 389 175 423 209
rect 507 175 541 209
rect 626 175 660 209
rect 757 175 791 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 828 521
rect 19 437 71 453
rect 19 403 35 437
rect 69 403 71 437
rect 19 369 71 403
rect 19 335 35 369
rect 69 335 71 369
rect 19 61 71 335
rect 105 445 267 487
rect 105 411 121 445
rect 155 411 217 445
rect 251 411 267 445
rect 105 377 267 411
rect 105 343 121 377
rect 155 343 217 377
rect 251 343 267 377
rect 105 327 267 343
rect 301 437 367 453
rect 301 403 317 437
rect 351 403 367 437
rect 301 369 367 403
rect 301 335 317 369
rect 351 335 367 369
rect 301 293 367 335
rect 404 445 552 487
rect 404 343 419 445
rect 521 343 552 445
rect 404 327 552 343
rect 586 437 636 453
rect 746 445 811 487
rect 586 403 602 437
rect 586 309 636 403
rect 586 293 602 309
rect 139 275 602 293
rect 139 259 636 275
rect 139 225 173 259
rect 670 225 707 443
rect 746 411 758 445
rect 792 411 811 445
rect 746 377 811 411
rect 746 343 758 377
rect 792 343 811 377
rect 746 327 811 343
rect 105 209 173 225
rect 139 175 173 209
rect 253 209 349 225
rect 253 175 269 209
rect 303 175 349 209
rect 105 159 173 175
rect 139 141 173 159
rect 139 121 273 141
rect 139 107 223 121
rect 205 87 223 107
rect 257 87 273 121
rect 19 27 35 61
rect 69 27 71 61
rect 19 11 71 27
rect 107 53 169 73
rect 107 19 119 53
rect 153 19 169 53
rect 107 -23 169 19
rect 205 53 273 87
rect 205 19 223 53
rect 257 19 273 53
rect 307 38 349 175
rect 385 209 439 225
rect 385 175 389 209
rect 423 175 439 209
rect 385 38 439 175
rect 489 209 541 225
rect 489 175 507 209
rect 610 209 707 225
rect 610 175 626 209
rect 660 175 707 209
rect 741 209 807 292
rect 741 175 757 209
rect 791 175 807 209
rect 489 159 541 175
rect 489 38 538 159
rect 574 129 811 135
rect 574 95 590 129
rect 624 101 811 129
rect 624 95 632 101
rect 574 61 632 95
rect 205 11 273 19
rect 574 27 590 61
rect 624 27 632 61
rect 574 11 632 27
rect 666 51 724 67
rect 666 17 674 51
rect 708 17 724 51
rect 666 -23 724 17
rect 758 61 811 101
rect 792 27 811 61
rect 758 11 811 27
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 828 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
<< metal1 >>
rect 0 521 828 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 828 521
rect 0 456 828 487
rect 0 -23 828 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 828 -23
rect 0 -88 828 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 o2111a_1
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 29 385 63 419 0 FreeSans 400 0 0 0 X
port 8 nsew
flabel locali s 29 317 63 351 0 FreeSans 400 0 0 0 X
port 8 nsew
flabel locali s 29 181 63 215 0 FreeSans 400 0 0 0 X
port 8 nsew
flabel locali s 29 113 63 147 0 FreeSans 400 0 0 0 X
port 8 nsew
flabel locali s 29 45 63 79 0 FreeSans 400 0 0 0 X
port 8 nsew
flabel locali s 305 181 339 215 0 FreeSans 400 0 0 0 D1
port 9 nsew
flabel locali s 397 181 431 215 0 FreeSans 400 0 0 0 C1
port 10 nsew
flabel locali s 397 113 431 147 0 FreeSans 400 0 0 0 C1
port 10 nsew
flabel locali s 397 45 431 79 0 FreeSans 400 0 0 0 C1
port 10 nsew
flabel locali s 489 181 523 215 0 FreeSans 400 0 0 0 B1
port 11 nsew
flabel locali s 673 181 707 215 0 FreeSans 400 0 0 0 A2
port 12 nsew
flabel locali s 765 249 799 283 0 FreeSans 400 0 0 0 A1
port 13 nsew
flabel locali s 765 181 799 215 0 FreeSans 400 0 0 0 A1
port 13 nsew
flabel locali s 29 249 63 283 0 FreeSans 400 0 0 0 X
port 8 nsew
<< properties >>
string FIXED_BBOX 0 -40 828 504
string path 0.000 -1.000 20.700 -1.000 
<< end >>
