magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_p >>
rect -36 -147 36 -141
rect -36 -181 -17 -147
rect -36 -187 36 -181
<< pwell >>
rect -124 -135 124 117
<< nmoslvt >>
rect -40 -109 40 91
<< ndiff >>
rect -98 76 -40 91
rect -98 42 -86 76
rect -52 42 -40 76
rect -98 8 -40 42
rect -98 -26 -86 8
rect -52 -26 -40 8
rect -98 -60 -40 -26
rect -98 -94 -86 -60
rect -52 -94 -40 -60
rect -98 -109 -40 -94
rect 40 76 98 91
rect 40 42 52 76
rect 86 42 98 76
rect 40 8 98 42
rect 40 -26 52 8
rect 86 -26 98 8
rect 40 -60 98 -26
rect 40 -94 52 -60
rect 86 -94 98 -60
rect 40 -109 98 -94
<< ndiffc >>
rect -86 42 -52 76
rect -86 -26 -52 8
rect -86 -94 -52 -60
rect 52 42 86 76
rect 52 -26 86 8
rect 52 -94 86 -60
<< poly >>
rect -40 91 40 117
rect -40 -147 40 -109
rect -40 -181 -17 -147
rect 17 -181 40 -147
rect -40 -197 40 -181
<< polycont >>
rect -17 -181 17 -147
<< locali >>
rect -86 76 -52 95
rect -86 8 -52 10
rect -86 -28 -52 -26
rect -86 -113 -52 -94
rect 52 76 86 95
rect 52 8 86 10
rect 52 -28 86 -26
rect 52 -113 86 -94
rect -40 -181 -17 -147
rect 17 -181 40 -147
<< viali >>
rect -86 42 -52 44
rect -86 10 -52 42
rect -86 -60 -52 -28
rect -86 -62 -52 -60
rect 52 42 86 44
rect 52 10 86 42
rect 52 -60 86 -28
rect 52 -62 86 -60
rect -17 -181 17 -147
<< metal1 >>
rect -92 44 -46 91
rect -92 10 -86 44
rect -52 10 -46 44
rect -92 -28 -46 10
rect -92 -62 -86 -28
rect -52 -62 -46 -28
rect -92 -109 -46 -62
rect 46 44 92 91
rect 46 10 52 44
rect 86 10 92 44
rect 46 -28 92 10
rect 46 -62 52 -28
rect 86 -62 92 -28
rect 46 -109 92 -62
rect -36 -147 36 -141
rect -36 -181 -17 -147
rect 17 -181 36 -147
rect -36 -187 36 -181
<< end >>
