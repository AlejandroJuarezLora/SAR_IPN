magic
tech sky130B
magscale 1 2
timestamp 1697155012
<< locali >>
rect 7759 4366 7922 4367
rect 3925 4329 4006 4364
rect 5819 4362 6019 4363
rect 5819 4328 5984 4362
rect 6018 4328 6019 4362
rect 7759 4332 7887 4366
rect 7921 4332 7922 4366
rect 9697 4364 9900 4365
rect 9697 4330 9865 4364
rect 9899 4330 9900 4364
<< viali >>
rect 27918 5394 27958 5434
rect 28100 5306 28140 5346
rect 27920 5127 27960 5167
rect 28079 5029 28119 5069
rect 27926 4847 27966 4887
rect 28082 4757 28122 4797
rect 27926 4577 27966 4617
rect 28081 4481 28121 4521
rect 4006 4329 4041 4364
rect 5984 4328 6018 4362
rect 7887 4332 7921 4366
rect 9865 4330 9899 4364
rect 27920 4290 27964 4334
rect 28078 4210 28118 4250
rect 28081 3935 28121 3975
rect 27918 3838 27958 3878
rect 28084 3661 28124 3701
rect 27920 3576 27960 3616
rect 28086 3386 28126 3426
rect 27922 3298 27958 3334
rect 28082 3112 28122 3152
rect 27922 3032 27957 3067
<< metal1 >>
rect 4953 5309 4988 7085
rect 28235 5611 28269 5747
rect 10557 5577 28269 5611
rect 4945 5303 4997 5309
rect 4945 5245 4997 5251
rect 4953 4963 4988 5245
rect 4006 4928 9899 4963
rect 2383 4373 2435 4379
rect 4006 4376 4041 4928
rect 2383 4315 2435 4321
rect 4000 4364 4047 4376
rect 4000 4329 4006 4364
rect 4041 4329 4047 4364
rect 4000 4317 4047 4329
rect 4302 4320 4308 4372
rect 4360 4320 4366 4372
rect 5983 4368 6018 4928
rect 7886 4378 7921 4928
rect 5972 4362 6030 4368
rect 5972 4328 5984 4362
rect 6018 4328 6030 4362
rect 5972 4322 6030 4328
rect 6222 4320 6228 4372
rect 6280 4320 6286 4372
rect 7881 4366 7927 4378
rect 7881 4332 7887 4366
rect 7921 4332 7927 4366
rect 7881 4320 7927 4332
rect 8151 4325 8157 4377
rect 8209 4325 8215 4377
rect 9864 4376 9899 4928
rect 9859 4364 9905 4376
rect 9859 4330 9865 4364
rect 9899 4330 9905 4364
rect 9859 4318 9905 4330
rect 10557 3663 10591 5577
rect 27671 5417 27705 5465
rect 27912 5440 27964 5446
rect 27912 5382 27964 5388
rect 28235 5380 28269 5577
rect 28094 5352 28146 5358
rect 27418 5248 27482 5311
rect 27545 5248 27551 5311
rect 28094 5294 28146 5300
rect 27914 5173 27966 5179
rect 27914 5115 27966 5121
rect 28073 5075 28125 5081
rect 28073 5017 28125 5023
rect 27920 4893 27972 4899
rect 27920 4835 27972 4841
rect 28076 4803 28128 4809
rect 28076 4745 28128 4751
rect 27423 4647 27504 4731
rect 27562 4647 27568 4731
rect 27920 4623 27972 4629
rect 27920 4565 27972 4571
rect 28075 4527 28127 4533
rect 28075 4469 28127 4475
rect 27914 4340 27970 4346
rect 27914 4278 27970 4284
rect 28072 4256 28124 4262
rect 28072 4198 28124 4204
rect 27409 4028 27458 4112
rect 27542 4028 27548 4112
rect 28075 3981 28127 3987
rect 28075 3923 28127 3929
rect 27912 3884 27964 3890
rect 27912 3826 27964 3832
rect 9893 3629 10591 3663
rect 28078 3707 28130 3713
rect 28078 3649 28130 3655
rect 27914 3622 27966 3628
rect 27908 3570 27914 3622
rect 27966 3570 27972 3622
rect 27914 3564 27966 3570
rect 28080 3432 28132 3438
rect 28080 3374 28132 3380
rect 27802 3334 27970 3340
rect 27802 3298 27922 3334
rect 27958 3298 27970 3334
rect 27802 3292 27970 3298
rect 9749 2804 9796 3119
rect 27674 2804 27721 3208
rect 9749 2757 27721 2804
rect 27674 1581 27721 2757
rect 27802 2385 27850 3292
rect 28076 3158 28128 3164
rect 28076 3100 28128 3106
rect 27916 3067 27963 3079
rect 27916 3032 27922 3067
rect 27957 3032 27963 3067
rect 27779 2303 27852 2385
rect 27779 2224 27852 2230
rect 27916 1730 27963 3032
rect 27901 1724 27964 1730
rect 27901 1655 27964 1661
rect 27669 1473 27721 1581
rect 27669 1171 27716 1473
<< via1 >>
rect 4945 5251 4997 5303
rect 2383 4321 2435 4373
rect 4308 4320 4360 4372
rect 6228 4320 6280 4372
rect 8157 4325 8209 4377
rect 27912 5434 27964 5440
rect 27912 5394 27918 5434
rect 27918 5394 27958 5434
rect 27958 5394 27964 5434
rect 27912 5388 27964 5394
rect 28094 5346 28146 5352
rect 27482 5248 27545 5311
rect 28094 5306 28100 5346
rect 28100 5306 28140 5346
rect 28140 5306 28146 5346
rect 28094 5300 28146 5306
rect 27914 5167 27966 5173
rect 27914 5127 27920 5167
rect 27920 5127 27960 5167
rect 27960 5127 27966 5167
rect 27914 5121 27966 5127
rect 28073 5069 28125 5075
rect 28073 5029 28079 5069
rect 28079 5029 28119 5069
rect 28119 5029 28125 5069
rect 28073 5023 28125 5029
rect 27920 4887 27972 4893
rect 27920 4847 27926 4887
rect 27926 4847 27966 4887
rect 27966 4847 27972 4887
rect 27920 4841 27972 4847
rect 28076 4797 28128 4803
rect 28076 4757 28082 4797
rect 28082 4757 28122 4797
rect 28122 4757 28128 4797
rect 28076 4751 28128 4757
rect 27504 4647 27562 4731
rect 27920 4617 27972 4623
rect 27920 4577 27926 4617
rect 27926 4577 27966 4617
rect 27966 4577 27972 4617
rect 27920 4571 27972 4577
rect 28075 4521 28127 4527
rect 28075 4481 28081 4521
rect 28081 4481 28121 4521
rect 28121 4481 28127 4521
rect 28075 4475 28127 4481
rect 27914 4334 27970 4340
rect 27914 4290 27920 4334
rect 27920 4290 27964 4334
rect 27964 4290 27970 4334
rect 27914 4284 27970 4290
rect 28072 4250 28124 4256
rect 28072 4210 28078 4250
rect 28078 4210 28118 4250
rect 28118 4210 28124 4250
rect 28072 4204 28124 4210
rect 27458 4028 27542 4112
rect 28075 3975 28127 3981
rect 28075 3935 28081 3975
rect 28081 3935 28121 3975
rect 28121 3935 28127 3975
rect 28075 3929 28127 3935
rect 27912 3878 27964 3884
rect 27912 3838 27918 3878
rect 27918 3838 27958 3878
rect 27958 3838 27964 3878
rect 27912 3832 27964 3838
rect 28078 3701 28130 3707
rect 28078 3661 28084 3701
rect 28084 3661 28124 3701
rect 28124 3661 28130 3701
rect 28078 3655 28130 3661
rect 27914 3616 27966 3622
rect 27914 3576 27920 3616
rect 27920 3576 27960 3616
rect 27960 3576 27966 3616
rect 27914 3570 27966 3576
rect 28080 3426 28132 3432
rect 28080 3386 28086 3426
rect 28086 3386 28126 3426
rect 28126 3386 28132 3426
rect 28080 3380 28132 3386
rect 28076 3152 28128 3158
rect 28076 3112 28082 3152
rect 28082 3112 28122 3152
rect 28122 3112 28128 3152
rect 28076 3106 28128 3112
rect 27779 2230 27852 2303
rect 27901 1661 27964 1724
<< metal2 >>
rect 27397 6446 27403 6535
rect 27492 6514 27498 6535
rect 27492 6466 27968 6514
rect 27492 6446 27498 6466
rect 27411 5893 27709 5908
rect 27411 5850 27808 5893
rect 27411 5832 27709 5850
rect 4941 5307 5001 5316
rect 27482 5311 27545 5317
rect 4939 5251 4941 5303
rect 5001 5251 5003 5303
rect 4941 5238 5001 5247
rect 27482 5242 27545 5248
rect 212 5032 8200 5068
rect 2391 4373 2427 5032
rect 4316 4378 4352 5032
rect 6236 4378 6272 5032
rect 8165 4383 8200 5032
rect 27500 4886 27539 5242
rect 27765 5165 27808 5850
rect 27920 5440 27968 6466
rect 27906 5388 27912 5440
rect 27964 5388 27970 5440
rect 28088 5300 28094 5352
rect 28146 5348 28152 5352
rect 28146 5304 28378 5348
rect 28146 5300 28152 5304
rect 27908 5165 27914 5173
rect 27765 5122 27914 5165
rect 27908 5121 27914 5122
rect 27966 5121 27972 5173
rect 28067 5023 28073 5075
rect 28125 5069 28131 5075
rect 28125 5029 28378 5069
rect 28125 5023 28131 5029
rect 27914 4886 27920 4893
rect 27500 4847 27920 4886
rect 27914 4841 27920 4847
rect 27972 4841 27978 4893
rect 28070 4751 28076 4803
rect 28128 4797 28134 4803
rect 28128 4757 28378 4797
rect 28128 4751 28134 4757
rect 27504 4731 27562 4737
rect 27504 4614 27562 4647
rect 27914 4614 27920 4623
rect 27504 4579 27920 4614
rect 27504 4567 27562 4579
rect 27914 4571 27920 4579
rect 27972 4571 27978 4623
rect 28069 4475 28075 4527
rect 28127 4521 28133 4527
rect 28127 4481 28378 4521
rect 28127 4475 28133 4481
rect 2377 4321 2383 4373
rect 2435 4321 2441 4373
rect 4308 4372 4360 4378
rect 4308 4314 4360 4320
rect 6228 4372 6280 4378
rect 6228 4314 6280 4320
rect 8157 4377 8209 4383
rect 8157 4319 8209 4325
rect 27472 4284 27914 4340
rect 27970 4284 27976 4340
rect 27472 4118 27528 4284
rect 28066 4204 28072 4256
rect 28124 4250 28130 4256
rect 28124 4210 28378 4250
rect 28124 4204 28130 4210
rect 27458 4112 27542 4118
rect 27458 4022 27542 4028
rect 28069 3929 28075 3981
rect 28127 3975 28133 3981
rect 28127 3934 28378 3975
rect 28127 3929 28133 3934
rect 27906 3883 27912 3884
rect 27506 3832 27912 3883
rect 27964 3832 27970 3884
rect 27506 3537 27557 3832
rect 28072 3655 28078 3707
rect 28130 3701 28136 3707
rect 28130 3660 28378 3701
rect 28130 3655 28136 3660
rect 27505 3531 27557 3537
rect 27416 3449 27557 3531
rect 27505 3443 27557 3449
rect 27914 3622 27966 3628
rect 3038 2887 3079 3039
rect 4963 2887 5004 3040
rect 6882 2887 6923 3032
rect 8807 2887 8848 3042
rect 198 2846 8848 2887
rect 27423 2913 27599 2937
rect 27914 2913 27966 3570
rect 28074 3380 28080 3432
rect 28132 3426 28138 3432
rect 28132 3386 28378 3426
rect 28132 3380 28138 3386
rect 28070 3106 28076 3158
rect 28128 3152 28134 3158
rect 28128 3112 28378 3152
rect 28128 3106 28134 3112
rect 27423 2861 27966 2913
rect 27423 2856 27599 2861
rect 27542 2855 27594 2856
rect 27422 2230 27779 2303
rect 27852 2230 27858 2303
rect 27419 1661 27901 1724
rect 27964 1661 27970 1724
<< via2 >>
rect 4941 5303 5001 5307
rect 4941 5251 4945 5303
rect 4945 5251 4997 5303
rect 4997 5251 5001 5303
rect 4941 5247 5001 5251
<< metal3 >>
rect 4920 5312 5018 5328
rect 4920 5248 4936 5312
rect 5006 5248 5018 5312
rect 4920 5247 4941 5248
rect 5001 5247 5018 5248
rect 4920 5228 5018 5247
<< via3 >>
rect 4936 5307 5006 5312
rect 4936 5248 4941 5307
rect 4941 5248 5001 5307
rect 5001 5248 5006 5307
<< metal4 >>
rect 4941 5313 5001 5512
rect 4935 5312 5007 5313
rect 4935 5248 4936 5312
rect 5006 5248 5007 5312
rect 4935 5247 5007 5248
use carray  carray_0
timestamp 1697065033
transform 1 0 270 0 1 6536
box 62 -5400 27238 480
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1693170804
transform 0 1 27702 -1 0 5189
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_2
timestamp 1693170804
transform 0 1 27702 1 0 2990
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_3
timestamp 1693170804
transform 0 1 27702 1 0 3540
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_4
timestamp 1693170804
transform 0 1 27702 -1 0 4637
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_5
timestamp 1693170804
transform 0 1 27702 -1 0 4913
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_6
timestamp 1693170804
transform 0 1 27702 1 0 3812
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_7
timestamp 1693170804
transform 0 1 27702 -1 0 4364
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_8
timestamp 1693170804
transform 0 1 27702 1 0 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_9
timestamp 1693170804
transform 0 1 27702 -1 0 5465
box -38 -48 314 592
use sw_top  sw_top_0
timestamp 1697152928
transform 1 0 8411 0 1 3890
box -410 -892 1590 1027
use sw_top  sw_top_1
timestamp 1697152928
transform 1 0 6488 0 1 3890
box -410 -892 1590 1027
use sw_top  sw_top_2
timestamp 1697152928
transform 1 0 4565 0 1 3890
box -410 -892 1590 1027
use sw_top  sw_top_3
timestamp 1697152928
transform 1 0 2642 0 1 3890
box -410 -892 1590 1027
<< labels >>
flabel metal1 s 28235 5713 28269 5747 0 FreeSans 640 0 0 0 vdd
port 12 nsew
flabel metal1 s 27669 1171 27716 1218 0 FreeSans 640 0 0 0 vss
port 13 nsew
flabel metal2 s 28338 3112 28378 3152 0 FreeSans 800 0 0 0 dum
port 11 nsew
flabel metal2 s 28338 3386 28378 3426 0 FreeSans 800 0 0 0 ctl_0_
port 10 nsew
flabel metal2 s 28337 3660 28378 3701 0 FreeSans 800 0 0 0 ctl_1_
port 9 nsew
flabel metal2 s 28337 3934 28378 3975 0 FreeSans 800 0 0 0 ctl_2_
port 8 nsew
flabel metal2 s 28338 4210 28378 4250 0 FreeSans 800 0 0 0 ctl_3_
port 7 nsew
flabel metal2 s 28338 4481 28378 4521 0 FreeSans 800 0 0 0 ctl_4_
port 6 nsew
flabel metal2 s 28338 4757 28378 4797 0 FreeSans 800 0 0 0 ctl_5_
port 5 nsew
flabel metal2 s 28338 5029 28378 5069 0 FreeSans 800 0 0 0 ctl_6_
port 4 nsew
flabel metal2 s 28334 5304 28378 5348 0 FreeSans 800 0 0 0 ctl_7_
port 3 nsew
flabel metal2 216 5032 252 5068 0 FreeSans 800 0 0 0 vin
port 0 nsew
flabel metal2 216 2846 263 2887 0 FreeSans 800 0 0 0 sample
port 1 nsew
flabel metal1 4953 7050 4988 7085 0 FreeSans 800 0 0 0 out
port 2 nsew
<< end >>
