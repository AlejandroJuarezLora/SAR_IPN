magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 682 542
<< pwell >>
rect 1 -19 643 163
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 109 137
rect 163 7 193 137
rect 367 7 397 137
rect 451 7 481 137
rect 535 7 565 137
<< scpmoshvt >>
rect 79 257 109 457
rect 151 257 181 457
rect 367 257 397 457
rect 451 257 481 457
rect 535 257 565 457
<< ndiff >>
rect 27 121 79 137
rect 27 87 35 121
rect 69 87 79 121
rect 27 53 79 87
rect 27 19 35 53
rect 69 19 79 53
rect 27 7 79 19
rect 109 89 163 137
rect 109 55 119 89
rect 153 55 163 89
rect 109 7 163 55
rect 193 53 367 137
rect 193 19 203 53
rect 237 19 271 53
rect 305 19 367 53
rect 193 7 367 19
rect 397 89 451 137
rect 397 55 407 89
rect 441 55 451 89
rect 397 7 451 55
rect 481 7 535 137
rect 565 121 617 137
rect 565 87 575 121
rect 609 87 617 121
rect 565 53 617 87
rect 565 19 575 53
rect 609 19 617 53
rect 565 7 617 19
<< pdiff >>
rect 27 443 79 457
rect 27 409 35 443
rect 69 409 79 443
rect 27 375 79 409
rect 27 341 35 375
rect 69 341 79 375
rect 27 257 79 341
rect 109 257 151 457
rect 181 441 233 457
rect 181 407 191 441
rect 225 407 233 441
rect 181 373 233 407
rect 181 339 191 373
rect 225 339 233 373
rect 181 305 233 339
rect 181 271 191 305
rect 225 271 233 305
rect 181 257 233 271
rect 299 441 367 457
rect 299 407 307 441
rect 341 407 367 441
rect 299 373 367 407
rect 299 339 323 373
rect 357 339 367 373
rect 299 257 367 339
rect 397 441 451 457
rect 397 407 407 441
rect 441 407 451 441
rect 397 257 451 407
rect 481 449 535 457
rect 481 415 491 449
rect 525 415 535 449
rect 481 257 535 415
rect 565 437 617 457
rect 565 403 575 437
rect 609 403 617 437
rect 565 351 617 403
rect 565 317 575 351
rect 609 317 617 351
rect 565 257 617 317
<< ndiffc >>
rect 35 87 69 121
rect 35 19 69 53
rect 119 55 153 89
rect 203 19 237 53
rect 271 19 305 53
rect 407 55 441 89
rect 575 87 609 121
rect 575 19 609 53
<< pdiffc >>
rect 35 409 69 443
rect 35 341 69 375
rect 191 407 225 441
rect 191 339 225 373
rect 191 271 225 305
rect 307 407 341 441
rect 323 339 357 373
rect 407 407 441 441
rect 491 415 525 449
rect 575 403 609 437
rect 575 317 609 351
<< poly >>
rect 79 457 109 483
rect 151 457 181 483
rect 367 457 397 483
rect 451 457 481 483
rect 535 457 565 483
rect 79 225 109 257
rect 55 209 109 225
rect 55 175 65 209
rect 99 175 109 209
rect 55 159 109 175
rect 151 225 181 257
rect 367 225 397 257
rect 451 225 481 257
rect 535 225 565 257
rect 151 209 205 225
rect 151 175 161 209
rect 195 175 205 209
rect 151 159 205 175
rect 271 209 397 225
rect 271 175 282 209
rect 316 175 397 209
rect 271 159 397 175
rect 439 209 493 225
rect 439 175 449 209
rect 483 175 493 209
rect 439 159 493 175
rect 535 209 600 225
rect 535 175 556 209
rect 590 175 600 209
rect 535 159 600 175
rect 79 137 109 159
rect 163 137 193 159
rect 367 137 397 159
rect 451 137 481 159
rect 535 137 565 159
rect 79 -19 109 7
rect 163 -19 193 7
rect 367 -19 397 7
rect 451 -19 481 7
rect 535 -19 565 7
<< polycont >>
rect 65 175 99 209
rect 161 175 195 209
rect 282 175 316 209
rect 449 175 483 209
rect 556 175 590 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 644 521
rect 19 443 85 487
rect 19 409 35 443
rect 69 409 85 443
rect 19 375 85 409
rect 19 341 35 375
rect 69 341 85 375
rect 19 321 85 341
rect 175 441 241 453
rect 175 407 191 441
rect 225 407 241 441
rect 175 373 241 407
rect 175 339 191 373
rect 225 339 241 373
rect 175 305 241 339
rect 284 441 357 453
rect 284 407 307 441
rect 341 407 357 441
rect 391 441 457 453
rect 391 407 407 441
rect 441 407 457 441
rect 284 373 357 407
rect 284 339 323 373
rect 423 351 457 407
rect 491 449 541 487
rect 525 415 541 449
rect 491 387 541 415
rect 575 437 626 453
rect 609 403 626 437
rect 575 351 626 403
rect 357 339 389 351
rect 284 317 389 339
rect 423 317 575 351
rect 609 317 626 351
rect 30 209 104 283
rect 175 271 191 305
rect 225 283 241 305
rect 225 271 316 283
rect 175 249 316 271
rect 30 175 65 209
rect 99 175 104 209
rect 30 159 104 175
rect 145 209 248 215
rect 145 175 161 209
rect 195 175 248 209
rect 145 162 248 175
rect 282 209 316 249
rect 282 126 316 175
rect 19 121 85 125
rect 19 87 35 121
rect 69 87 85 121
rect 19 53 85 87
rect 19 19 35 53
rect 69 19 85 53
rect 19 -23 85 19
rect 119 92 316 126
rect 355 125 389 317
rect 449 209 522 283
rect 483 175 522 209
rect 449 159 522 175
rect 556 209 614 283
rect 590 175 614 209
rect 556 159 614 175
rect 119 89 153 92
rect 355 89 441 125
rect 119 11 153 55
rect 187 53 321 58
rect 187 19 203 53
rect 237 19 271 53
rect 305 19 321 53
rect 187 -23 321 19
rect 355 55 407 89
rect 355 11 441 55
rect 488 45 522 159
rect 559 121 625 125
rect 559 87 575 121
rect 609 87 625 121
rect 559 53 625 87
rect 559 19 575 53
rect 609 19 625 53
rect 559 -23 625 19
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 644 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
<< metal1 >>
rect 0 521 644 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 644 521
rect 0 456 644 487
rect 0 -23 644 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 644 -23
rect 0 -88 644 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 a2bb2oi_1
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 30 249 64 283 0 FreeSans 200 0 0 0 A1_N
port 9 nsew
flabel locali s 30 181 64 215 0 FreeSans 200 0 0 0 A1_N
port 9 nsew
flabel locali s 304 385 338 419 0 FreeSans 200 0 0 0 Y
port 7 nsew
flabel locali s 304 317 338 351 0 FreeSans 200 0 0 0 Y
port 7 nsew
flabel locali s 396 45 430 79 0 FreeSans 200 0 0 0 Y
port 7 nsew
flabel locali s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel locali s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel locali s 488 45 522 79 0 FreeSans 200 0 0 0 B2
port 10 nsew
flabel locali s 488 113 522 147 0 FreeSans 200 0 0 0 B2
port 10 nsew
flabel locali s 488 181 522 215 0 FreeSans 200 0 0 0 B2
port 10 nsew
flabel locali s 488 249 522 283 0 FreeSans 200 0 0 0 B2
port 10 nsew
flabel locali s 580 181 614 215 0 FreeSans 200 0 0 0 B1
port 11 nsew
flabel locali s 214 181 248 215 0 FreeSans 200 0 0 0 A2_N
port 8 nsew
<< properties >>
string FIXED_BBOX 0 -40 644 504
string path 0.000 -1.000 16.100 -1.000 
<< end >>
