magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 590 542
<< pwell >>
rect 269 123 551 163
rect 4 -13 551 123
rect 29 -57 63 -13
rect 272 -19 551 -13
<< scnmos >>
rect 82 13 112 97
rect 154 13 184 97
rect 235 13 265 97
rect 356 7 386 137
rect 440 7 470 137
<< scpmoshvt >>
rect 81 271 111 355
rect 165 271 195 355
rect 260 257 290 341
rect 359 257 389 457
rect 443 257 473 457
<< ndiff >>
rect 295 97 356 137
rect 30 71 82 97
rect 30 37 38 71
rect 72 37 82 71
rect 30 13 82 37
rect 112 13 154 97
rect 184 13 235 97
rect 265 76 356 97
rect 265 42 311 76
rect 345 42 356 76
rect 265 13 356 42
rect 298 7 356 13
rect 386 83 440 137
rect 386 49 396 83
rect 430 49 440 83
rect 386 7 440 49
rect 470 80 525 137
rect 470 46 480 80
rect 514 46 525 80
rect 470 7 525 46
<< pdiff >>
rect 305 437 359 457
rect 305 403 315 437
rect 349 403 359 437
rect 305 368 359 403
rect 29 329 81 355
rect 29 295 37 329
rect 71 295 81 329
rect 29 271 81 295
rect 111 347 165 355
rect 111 313 121 347
rect 155 313 165 347
rect 111 271 165 313
rect 195 341 245 355
rect 305 341 315 368
rect 195 322 260 341
rect 195 288 216 322
rect 250 288 260 322
rect 195 271 260 288
rect 210 257 260 271
rect 290 334 315 341
rect 349 334 359 368
rect 290 257 359 334
rect 389 437 443 457
rect 389 403 399 437
rect 433 403 443 437
rect 389 369 443 403
rect 389 335 399 369
rect 433 335 443 369
rect 389 257 443 335
rect 473 437 525 457
rect 473 403 483 437
rect 517 403 525 437
rect 473 369 525 403
rect 473 335 483 369
rect 517 335 525 369
rect 473 257 525 335
<< ndiffc >>
rect 38 37 72 71
rect 311 42 345 76
rect 396 49 430 83
rect 480 46 514 80
<< pdiffc >>
rect 315 403 349 437
rect 37 295 71 329
rect 121 313 155 347
rect 216 288 250 322
rect 315 334 349 368
rect 399 403 433 437
rect 399 335 433 369
rect 483 403 517 437
rect 483 335 517 369
<< poly >>
rect 165 437 223 460
rect 359 457 389 483
rect 443 457 473 483
rect 165 403 179 437
rect 213 403 223 437
rect 165 387 223 403
rect 81 355 111 385
rect 165 355 195 387
rect 260 341 290 367
rect 81 225 111 271
rect 165 256 195 271
rect 154 239 195 256
rect 154 230 193 239
rect 28 209 112 225
rect 28 175 38 209
rect 72 175 112 209
rect 28 159 112 175
rect 82 97 112 159
rect 154 212 192 230
rect 260 225 290 257
rect 359 225 389 257
rect 443 225 473 257
rect 154 97 184 212
rect 235 209 292 225
rect 235 175 245 209
rect 279 175 292 209
rect 235 159 292 175
rect 334 209 474 225
rect 334 175 344 209
rect 378 175 474 209
rect 334 159 474 175
rect 235 97 265 159
rect 356 137 386 159
rect 440 137 470 159
rect 82 -13 112 13
rect 154 -13 184 13
rect 235 -13 265 13
rect 356 -19 386 7
rect 440 -19 470 7
<< polycont >>
rect 179 403 213 437
rect 38 175 72 209
rect 245 175 279 209
rect 344 175 378 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 552 521
rect 17 386 143 487
rect 20 329 71 352
rect 20 295 37 329
rect 105 351 143 386
rect 179 437 274 453
rect 213 403 274 437
rect 179 385 274 403
rect 311 437 354 487
rect 311 403 315 437
rect 349 403 354 437
rect 311 368 354 403
rect 105 347 171 351
rect 105 313 121 347
rect 155 313 171 347
rect 216 322 266 338
rect 20 279 71 295
rect 250 288 266 322
rect 311 334 315 368
rect 349 334 354 368
rect 311 318 354 334
rect 394 437 449 453
rect 394 403 399 437
rect 433 403 449 437
rect 394 369 449 403
rect 394 335 399 369
rect 433 335 449 369
rect 394 319 449 335
rect 216 279 266 288
rect 20 245 378 279
rect 415 249 449 319
rect 483 437 535 487
rect 517 403 535 437
rect 483 369 535 403
rect 517 335 535 369
rect 483 285 535 335
rect 17 175 38 209
rect 72 175 94 209
rect 17 113 94 175
rect 128 74 179 245
rect 332 209 378 245
rect 21 71 179 74
rect 21 37 38 71
rect 72 37 179 71
rect 21 21 179 37
rect 213 175 245 209
rect 279 175 295 209
rect 213 110 295 175
rect 332 175 344 209
rect 332 159 378 175
rect 412 145 535 249
rect 213 21 259 110
rect 412 103 446 145
rect 396 83 446 103
rect 295 42 311 76
rect 345 42 361 76
rect 295 -23 361 42
rect 430 49 446 83
rect 396 11 446 49
rect 480 80 535 109
rect 514 46 535 80
rect 480 -23 535 46
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 552 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
<< metal1 >>
rect 0 521 552 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 552 521
rect 0 456 552 487
rect 0 -23 552 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 552 -23
rect 0 -88 552 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 and3_2
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 46 504 46 504 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 46 -40 46 -40 0 FreeSans 200 0 0 0 VGND
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 213 385 247 419 0 FreeSans 400 0 0 0 B
port 9 nsew
flabel locali s 397 45 431 79 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 397 385 431 419 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 29 113 63 147 0 FreeSans 400 0 0 0 A
port 10 nsew
flabel locali s 213 113 247 147 0 FreeSans 400 0 0 0 C
port 8 nsew
flabel locali s 489 181 523 215 0 FreeSans 200 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 552 504
<< end >>
