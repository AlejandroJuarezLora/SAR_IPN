magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 866 542
<< pwell >>
rect 1 117 269 163
rect 1 -19 827 117
rect 30 -57 64 -19
<< scnmos >>
rect 79 7 109 137
rect 163 7 193 137
rect 258 7 288 91
rect 353 7 383 91
rect 548 7 578 91
rect 633 7 663 91
rect 717 7 747 91
<< scpmoshvt >>
rect 79 257 109 457
rect 163 257 193 457
rect 276 329 306 457
rect 449 329 479 457
rect 561 329 591 457
rect 633 329 663 457
rect 717 329 747 457
<< ndiff >>
rect 27 121 79 137
rect 27 87 35 121
rect 69 87 79 121
rect 27 53 79 87
rect 27 19 35 53
rect 69 19 79 53
rect 27 7 79 19
rect 109 61 163 137
rect 109 27 119 61
rect 153 27 163 61
rect 109 7 163 27
rect 193 91 243 137
rect 193 53 258 91
rect 193 19 203 53
rect 237 19 258 53
rect 193 7 258 19
rect 288 7 353 91
rect 383 53 548 91
rect 383 19 393 53
rect 427 19 496 53
rect 530 19 548 53
rect 383 7 548 19
rect 578 7 633 91
rect 663 61 717 91
rect 663 27 673 61
rect 707 27 717 61
rect 663 7 717 27
rect 747 61 801 91
rect 747 27 759 61
rect 793 27 801 61
rect 747 7 801 27
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 377 79 411
rect 27 343 35 377
rect 69 343 79 377
rect 27 309 79 343
rect 27 275 35 309
rect 69 275 79 309
rect 27 257 79 275
rect 109 437 163 457
rect 109 403 119 437
rect 153 403 163 437
rect 109 369 163 403
rect 109 335 119 369
rect 153 335 163 369
rect 109 257 163 335
rect 193 445 276 457
rect 193 411 213 445
rect 247 411 276 445
rect 193 329 276 411
rect 306 329 449 457
rect 479 445 561 457
rect 479 411 509 445
rect 543 411 561 445
rect 479 329 561 411
rect 591 329 633 457
rect 663 445 717 457
rect 663 411 673 445
rect 707 411 717 445
rect 663 329 717 411
rect 747 445 801 457
rect 747 411 759 445
rect 793 411 801 445
rect 747 377 801 411
rect 747 343 759 377
rect 793 343 801 377
rect 747 329 801 343
rect 193 257 243 329
<< ndiffc >>
rect 35 87 69 121
rect 35 19 69 53
rect 119 27 153 61
rect 203 19 237 53
rect 393 19 427 53
rect 496 19 530 53
rect 673 27 707 61
rect 759 27 793 61
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 35 275 69 309
rect 119 403 153 437
rect 119 335 153 369
rect 213 411 247 445
rect 509 411 543 445
rect 673 411 707 445
rect 759 411 793 445
rect 759 343 793 377
<< poly >>
rect 79 457 109 483
rect 163 457 193 483
rect 276 457 306 483
rect 449 457 479 483
rect 561 457 591 483
rect 633 457 663 483
rect 717 457 747 483
rect 79 225 109 257
rect 163 225 193 257
rect 276 225 306 329
rect 79 209 215 225
rect 79 175 171 209
rect 205 175 215 209
rect 79 159 215 175
rect 257 209 311 225
rect 257 175 267 209
rect 301 175 311 209
rect 257 159 311 175
rect 353 163 407 179
rect 79 137 109 159
rect 163 137 193 159
rect 258 91 288 159
rect 353 129 363 163
rect 397 129 407 163
rect 449 175 479 329
rect 561 271 591 329
rect 525 261 591 271
rect 525 227 541 261
rect 575 227 591 261
rect 525 217 591 227
rect 633 225 663 329
rect 717 225 747 329
rect 633 209 747 225
rect 633 175 674 209
rect 708 175 747 209
rect 449 165 591 175
rect 449 145 541 165
rect 353 113 407 129
rect 525 131 541 145
rect 575 131 591 165
rect 525 121 591 131
rect 633 159 747 175
rect 353 91 383 113
rect 548 91 578 121
rect 633 91 663 159
rect 717 91 747 159
rect 79 -19 109 7
rect 163 -19 193 7
rect 258 -19 288 7
rect 353 -19 383 7
rect 548 -19 578 7
rect 633 -19 663 7
rect 717 -19 747 7
<< polycont >>
rect 171 175 205 209
rect 267 175 301 209
rect 363 129 397 163
rect 541 227 575 261
rect 674 175 708 209
rect 541 131 575 165
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 828 521
rect 18 445 69 487
rect 18 411 35 445
rect 18 377 69 411
rect 18 343 35 377
rect 18 309 69 343
rect 18 275 35 309
rect 18 259 69 275
rect 103 437 165 453
rect 103 403 119 437
rect 153 403 165 437
rect 103 369 165 403
rect 205 445 263 487
rect 665 445 709 487
rect 205 411 213 445
rect 247 411 263 445
rect 205 395 263 411
rect 297 411 509 445
rect 543 411 559 445
rect 665 411 673 445
rect 707 411 709 445
rect 103 335 119 369
rect 153 335 165 369
rect 297 361 331 411
rect 665 395 709 411
rect 743 445 810 453
rect 743 411 759 445
rect 793 411 810 445
rect 743 377 810 411
rect 743 361 759 377
rect 103 279 165 335
rect 199 327 331 361
rect 365 343 759 361
rect 793 343 810 377
rect 365 327 810 343
rect 18 121 69 137
rect 18 87 35 121
rect 18 53 69 87
rect 18 19 35 53
rect 18 -23 69 19
rect 103 110 137 279
rect 199 225 233 327
rect 365 293 399 327
rect 171 209 233 225
rect 205 175 233 209
rect 171 159 233 175
rect 267 259 399 293
rect 455 261 618 285
rect 267 209 301 259
rect 455 227 541 261
rect 575 227 618 261
rect 455 223 618 227
rect 455 216 489 223
rect 267 159 301 175
rect 363 163 489 216
rect 672 209 710 285
rect 672 175 674 209
rect 708 175 710 209
rect 199 121 233 159
rect 397 129 489 163
rect 103 61 153 110
rect 199 87 321 121
rect 363 113 489 129
rect 525 131 541 165
rect 575 131 618 165
rect 525 107 618 131
rect 672 111 710 175
rect 103 27 119 61
rect 287 53 321 87
rect 103 11 153 27
rect 187 19 203 53
rect 237 19 253 53
rect 287 19 393 53
rect 427 19 496 53
rect 530 19 546 53
rect 580 44 618 107
rect 670 61 710 77
rect 670 27 673 61
rect 707 27 710 61
rect 187 -23 253 19
rect 670 -23 710 27
rect 744 61 810 327
rect 744 27 759 61
rect 793 27 810 61
rect 744 11 810 27
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 828 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
<< metal1 >>
rect 0 521 828 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 828 521
rect 0 456 828 487
rect 0 -23 828 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 828 -23
rect 0 -88 828 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 mux2_2
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 582 113 616 147 0 FreeSans 200 0 0 0 A1
port 8 nsew
flabel locali s 490 249 524 283 0 FreeSans 200 0 0 0 A0
port 9 nsew
flabel locali s 398 181 432 215 0 FreeSans 200 0 0 0 A0
port 9 nsew
flabel locali s 398 113 432 147 0 FreeSans 200 0 0 0 A0
port 9 nsew
flabel locali s 674 113 708 147 0 FreeSans 200 0 0 0 S
port 7 nsew
flabel locali s 582 45 616 79 0 FreeSans 200 0 0 0 A1
port 8 nsew
flabel locali s 122 385 156 419 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel locali s 122 317 156 351 0 FreeSans 200 0 0 0 X
port 10 nsew
flabel locali s 582 249 616 283 0 FreeSans 200 0 0 0 A0
port 9 nsew
flabel locali s 674 249 708 283 0 FreeSans 200 0 0 0 S
port 7 nsew
flabel locali s 674 181 708 215 0 FreeSans 200 0 0 0 S
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 828 504
string path 0.000 -1.000 20.700 -1.000 
<< end >>
