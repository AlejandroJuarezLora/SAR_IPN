* SPICE3 file created from sarlogic.ext - technology: sky130B

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.05
C0 VGND VPWR 0.546f
C1 VPB VPWR 0.0787f
C2 VPB VGND 0.116f
C3 VPWR VNB 0.619f
C4 VGND VNB 0.554f
C5 VPB VNB 0.428f
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=2.89
C0 VPB VGND 0.22f
C1 VPWR VGND 1.27f
C2 VPWR VPB 0.105f
C3 VPWR VNB 1.14f
C4 VGND VNB 0.992f
C5 VPB VNB 0.782f
.ends

.subckt sky130_fd_sc_hd__inv_2 VPWR VGND VPB VNB Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 Y VGND 0.155f
C1 VGND A 0.0638f
C2 VGND VPB 0.00649f
C3 VPWR VGND 0.0423f
C4 Y A 0.0894f
C5 Y VPB 0.0061f
C6 VPWR Y 0.209f
C7 VPB A 0.0742f
C8 VPWR A 0.0631f
C9 VPWR VPB 0.0521f
C10 VGND VNB 0.266f
C11 Y VNB 0.0332f
C12 VPWR VNB 0.246f
C13 A VNB 0.263f
C14 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__dfstp_1 VPWR VGND VPB VNB Q SET_B D CLK a_652_n19# a_1602_7#
+ a_562_373# a_1032_373# a_1296_7# a_796_7# a_586_7# a_1056_7# a_381_7# a_193_7# a_1140_373#
+ a_27_7# a_956_373# a_476_7# a_1224_7# a_1182_221#
X0 VPWR a_1032_373# a_1602_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1 a_1032_373# a_193_7# a_1056_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 VPWR SET_B a_1032_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_476_7# a_27_7# a_381_7# VNB sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X4 a_1296_7# a_1182_221# a_1224_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 a_1032_373# a_27_7# a_956_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X6 a_1182_221# a_1032_373# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X7 Q a_1602_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X8 a_652_n19# a_476_7# a_796_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X9 a_1140_373# a_193_7# a_1032_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X10 a_586_7# a_193_7# a_476_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X11 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_381_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X14 a_1224_7# a_27_7# a_1032_373# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X15 a_1182_221# a_1032_373# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X16 VGND a_1032_373# a_1602_7# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X17 a_956_373# a_476_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 Q a_1602_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X19 a_796_7# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X20 VPWR a_476_7# a_652_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VGND SET_B a_1296_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
X22 VGND a_652_n19# a_586_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X23 a_381_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X24 a_652_n19# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X25 a_562_373# a_27_7# a_476_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X27 VPWR a_1182_221# a_1140_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X28 a_476_7# a_193_7# a_381_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X29 a_1056_7# a_476_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X30 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X31 VPWR a_652_n19# a_562_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
C0 a_1032_373# a_1602_7# 0.111f
C1 Q a_193_7# 6.4e-20
C2 CLK VGND 0.0194f
C3 VPB Q 0.0174f
C4 D VPWR 0.0158f
C5 a_956_373# a_652_n19# 3.11e-19
C6 a_1224_7# a_652_n19# 1.57e-19
C7 a_1032_373# a_1140_373# 0.00523f
C8 a_1032_373# a_1296_7# 0.00384f
C9 a_1602_7# a_193_7# 4.3e-19
C10 SET_B a_27_7# 0.0407f
C11 a_1602_7# VPB 0.0453f
C12 D VGND 0.014f
C13 a_1182_221# a_1602_7# 0.144f
C14 a_476_7# a_381_7# 0.0356f
C15 SET_B VPWR 0.0807f
C16 a_652_n19# a_381_7# 7.79e-20
C17 a_193_7# a_381_7# 0.157f
C18 VPB a_381_7# 0.0101f
C19 VPWR a_27_7# 0.438f
C20 a_1182_221# a_1296_7# 1.84e-19
C21 a_796_7# SET_B 0.00149f
C22 a_586_7# a_476_7# 0.00807f
C23 SET_B VGND 0.338f
C24 a_586_7# a_193_7# 0.00206f
C25 VGND a_27_7# 0.164f
C26 a_1056_7# SET_B 0.00152f
C27 a_1032_373# a_476_7# 0.00329f
C28 a_1032_373# a_652_n19# 0.00971f
C29 SET_B Q 4.58e-19
C30 VPWR VGND 0.0687f
C31 a_1032_373# a_193_7# 0.0573f
C32 a_562_373# a_27_7# 0.0018f
C33 a_1056_7# a_27_7# 0.00248f
C34 a_1032_373# VPB 0.177f
C35 D a_381_7# 0.14f
C36 a_1182_221# a_1032_373# 0.344f
C37 Q a_27_7# 1.08e-19
C38 a_562_373# VPWR 0.0041f
C39 a_1224_7# SET_B 8.75e-19
C40 a_796_7# VGND 0.00583f
C41 a_652_n19# a_476_7# 0.26f
C42 a_193_7# a_476_7# 0.215f
C43 a_1602_7# SET_B 0.00213f
C44 VPB a_476_7# 0.146f
C45 VPWR Q 0.0704f
C46 a_193_7# a_652_n19# 0.0849f
C47 VPB a_652_n19# 0.0992f
C48 a_956_373# a_27_7# 0.00294f
C49 a_1224_7# a_27_7# 1.63e-19
C50 VPB a_193_7# 0.179f
C51 a_1602_7# a_27_7# 2.39e-19
C52 a_1182_221# a_193_7# 0.0728f
C53 a_1140_373# SET_B 6.31e-19
C54 a_956_373# VPWR 0.00457f
C55 a_1182_221# VPB 0.112f
C56 a_1296_7# SET_B 0.00167f
C57 a_1056_7# VGND 0.00386f
C58 a_1602_7# VPWR 0.135f
C59 VGND Q 0.0595f
C60 a_27_7# a_381_7# 0.0729f
C61 CLK a_193_7# 0.00156f
C62 VPB CLK 0.0702f
C63 a_1140_373# VPWR 0.00334f
C64 a_956_373# VGND 3.4e-19
C65 VPWR a_381_7# 0.0942f
C66 a_1224_7# VGND 0.00169f
C67 a_1602_7# VGND 0.0942f
C68 D a_476_7# 1.36e-19
C69 D a_193_7# 0.0606f
C70 VPB D 0.0485f
C71 a_1032_373# SET_B 0.215f
C72 VGND a_381_7# 0.0787f
C73 a_1296_7# VGND 0.00523f
C74 a_1602_7# Q 0.0715f
C75 a_1032_373# a_27_7# 0.183f
C76 a_562_373# a_381_7# 8.75e-19
C77 SET_B a_476_7# 0.203f
C78 SET_B a_652_n19# 0.157f
C79 a_1032_373# VPWR 0.257f
C80 SET_B a_193_7# 0.202f
C81 a_586_7# VGND 0.00172f
C82 VPB SET_B 0.143f
C83 a_27_7# a_476_7# 0.223f
C84 a_1182_221# SET_B 0.12f
C85 a_27_7# a_652_n19# 0.19f
C86 a_27_7# a_193_7# 0.797f
C87 VPB a_27_7# 0.226f
C88 VPWR a_476_7# 0.12f
C89 VPWR a_652_n19# 0.144f
C90 a_1182_221# a_27_7# 0.0608f
C91 a_1032_373# VGND 0.157f
C92 VPWR a_193_7# 0.101f
C93 VPB VPWR 0.218f
C94 a_796_7# a_476_7# 0.00184f
C95 a_1182_221# VPWR 0.123f
C96 a_796_7# a_652_n19# 0.00196f
C97 a_1032_373# a_1056_7# 0.0016f
C98 CLK a_27_7# 0.214f
C99 VGND a_476_7# 0.178f
C100 VGND a_652_n19# 0.0761f
C101 a_1032_373# Q 0.00365f
C102 VGND a_193_7# 0.219f
C103 VPB VGND 0.0173f
C104 CLK VPWR 0.0194f
C105 a_562_373# a_476_7# 0.00972f
C106 a_1182_221# VGND 0.0628f
C107 a_562_373# a_652_n19# 9.35e-20
C108 a_1056_7# a_652_n19# 3.94e-19
C109 a_1032_373# a_956_373# 0.00212f
C110 a_562_373# a_193_7# 4.45e-20
C111 a_1032_373# a_1224_7# 0.00536f
C112 D a_27_7# 0.103f
C113 a_586_7# a_381_7# 3.7e-19
C114 Q VNB 0.0834f
C115 VGND VNB 1.08f
C116 VPWR VNB 0.875f
C117 SET_B VNB 0.247f
C118 D VNB 0.107f
C119 CLK VNB 0.196f
C120 VPB VNB 1.93f
C121 a_381_7# VNB 0.0203f
C122 a_1602_7# VNB 0.126f
C123 a_1032_373# VNB 0.305f
C124 a_1182_221# VNB 0.128f
C125 a_476_7# VNB 0.286f
C126 a_652_n19# VNB 0.119f
C127 a_193_7# VNB 0.322f
C128 a_27_7# VNB 0.437f
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=1.97
C0 VPB VPWR 0.0858f
C1 VGND VPWR 0.903f
C2 VPB VGND 0.161f
C3 VPWR VNB 0.867f
C4 VGND VNB 0.761f
C5 VPB VNB 0.605f
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 B2 a_584_7# a_346_7#
+ a_256_7# a_250_257# a_93_n19#
X0 a_346_7# A2 a_256_7# VNB sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X1 a_250_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2 a_93_n19# A1 a_346_7# VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.146 ps=1.1 w=0.65 l=0.15
X3 a_93_n19# B1 a_250_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X4 VGND B2 a_584_7# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0683 ps=0.86 w=0.65 l=0.15
X5 VPWR a_93_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.33 ps=2.66 w=1 l=0.15
X6 VGND a_93_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.214 ps=1.96 w=0.65 l=0.15
X7 a_250_257# B2 a_93_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_256_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167 ps=1.16 w=0.65 l=0.15
X9 a_250_257# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.243 ps=1.49 w=1 l=0.15
X10 a_584_7# B1 a_93_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X11 VPWR A2 a_250_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
C0 A2 A3 0.0788f
C1 VGND a_256_7# 0.00394f
C2 A1 B1 0.0965f
C3 A3 a_250_257# 0.00602f
C4 a_346_7# VPWR 0.00109f
C5 A1 B2 3.14e-19
C6 VGND a_346_7# 0.00514f
C7 A3 a_256_7# 4.42e-19
C8 a_93_n19# B1 0.0774f
C9 a_584_7# VPWR 9.47e-19
C10 A2 B1 1.44e-20
C11 X VPWR 0.0849f
C12 VGND VPWR 0.076f
C13 B2 a_93_n19# 0.0147f
C14 A2 B2 1.46e-19
C15 VPB VPWR 0.0756f
C16 VGND a_584_7# 0.00683f
C17 VGND X 0.06f
C18 a_250_257# B1 0.0125f
C19 VPB X 0.0108f
C20 B2 a_250_257# 0.0344f
C21 VPB VGND 0.00788f
C22 A3 VPWR 0.0158f
C23 A1 a_93_n19# 0.0641f
C24 a_256_7# B1 2.07e-20
C25 A2 A1 0.0971f
C26 A3 X 2.45e-19
C27 A3 VGND 0.00974f
C28 A1 a_250_257# 0.0129f
C29 A3 VPB 0.0291f
C30 A2 a_93_n19# 0.0747f
C31 a_346_7# B1 5.39e-20
C32 VPWR B1 0.01f
C33 a_93_n19# a_250_257# 0.188f
C34 A2 a_250_257# 0.0129f
C35 a_584_7# B1 0.00143f
C36 B2 VPWR 0.0108f
C37 X B1 3.83e-20
C38 VGND B1 0.0344f
C39 VPB B1 0.0276f
C40 a_93_n19# a_256_7# 0.0114f
C41 B2 VGND 0.0469f
C42 A1 a_346_7# 0.00465f
C43 A2 a_256_7# 0.00256f
C44 B2 VPB 0.0355f
C45 A1 VPWR 0.016f
C46 A3 B1 7.88e-22
C47 A1 X 6.03e-20
C48 a_93_n19# a_346_7# 0.0119f
C49 B2 A3 9.12e-20
C50 A1 VGND 0.0133f
C51 A2 a_346_7# 0.00252f
C52 A1 VPB 0.0296f
C53 a_93_n19# VPWR 0.0907f
C54 A2 VPWR 0.0133f
C55 a_93_n19# a_584_7# 0.00278f
C56 a_93_n19# X 0.0841f
C57 VGND a_93_n19# 0.251f
C58 A2 X 1.19e-19
C59 A2 VGND 0.0114f
C60 a_250_257# VPWR 0.313f
C61 VPB a_93_n19# 0.0485f
C62 A2 VPB 0.0287f
C63 a_250_257# a_584_7# 2.43e-19
C64 a_250_257# X 5.42e-19
C65 B2 B1 0.0823f
C66 VGND a_250_257# 0.0072f
C67 a_256_7# VPWR 9.47e-19
C68 A3 a_93_n19# 0.124f
C69 VPB a_250_257# 0.00616f
C70 VGND VNB 0.465f
C71 VPWR VNB 0.365f
C72 X VNB 0.0937f
C73 B2 VNB 0.14f
C74 B1 VNB 0.101f
C75 A1 VNB 0.0951f
C76 A2 VNB 0.0921f
C77 A3 VNB 0.0929f
C78 VPB VNB 0.782f
C79 a_250_257# VNB 0.0278f
C80 a_93_n19# VNB 0.151f
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR VPB VNB CLK D RESET_B Q a_639_7# a_805_7#
+ a_448_7# a_543_7# a_1283_n19# a_1462_7# a_1270_373# a_193_7# a_1217_7# a_761_249#
+ a_27_7# a_1108_7# a_651_373#
X0 VGND a_1283_n19# a_1217_7# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1 a_543_7# a_193_7# a_448_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2 VPWR a_1283_n19# a_1270_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR a_1108_7# a_1283_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1108_7# a_193_7# a_761_249# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 a_1270_373# a_193_7# a_1108_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1283_n19# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7 VPWR a_761_249# a_651_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X8 a_543_7# a_27_7# a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X9 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X10 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X11 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X12 a_651_373# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X13 a_761_249# a_543_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X14 VGND RESET_B a_805_7# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_651_373# a_27_7# a_543_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X16 a_1217_7# a_27_7# a_1108_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X17 a_448_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X18 a_639_7# a_193_7# a_543_7# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X19 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X20 a_448_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X21 a_1283_n19# a_1108_7# a_1462_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X22 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X23 a_805_7# a_761_249# a_639_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X24 a_1462_7# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X25 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X26 a_1108_7# a_27_7# a_761_249# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X27 a_761_249# a_543_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
C0 a_543_7# RESET_B 0.153f
C1 a_193_7# Q 1.81e-19
C2 a_193_7# a_761_249# 0.186f
C3 a_639_7# a_761_249# 3.16e-19
C4 Q VPWR 0.0997f
C5 a_193_7# a_543_7# 0.23f
C6 VGND a_1108_7# 0.148f
C7 a_193_7# RESET_B 0.0269f
C8 a_543_7# a_639_7# 0.0138f
C9 VPWR a_761_249# 0.105f
C10 RESET_B a_639_7# 9.54e-19
C11 a_27_7# Q 2.63e-20
C12 VGND a_1217_7# 9.68e-19
C13 VGND a_1283_n19# 0.24f
C14 a_543_7# VPWR 0.1f
C15 VPB VGND 0.00999f
C16 VGND a_448_7# 0.0661f
C17 a_1217_7# a_1108_7# 0.00742f
C18 RESET_B VPWR 0.0652f
C19 a_27_7# a_761_249# 0.0701f
C20 a_1283_n19# a_1108_7# 0.234f
C21 VPB a_1108_7# 0.113f
C22 a_27_7# a_543_7# 0.115f
C23 a_27_7# RESET_B 0.296f
C24 VPB a_1283_n19# 0.137f
C25 a_193_7# a_639_7# 2.28e-19
C26 CLK VGND 0.0172f
C27 VPB a_448_7# 0.0141f
C28 VGND D 0.0516f
C29 a_193_7# VPWR 0.396f
C30 VPB a_651_373# 0.0135f
C31 a_1270_373# a_1108_7# 0.00645f
C32 VGND a_1462_7# 0.00221f
C33 VPB CLK 0.0693f
C34 VPB D 0.138f
C35 a_27_7# a_193_7# 0.906f
C36 a_448_7# D 0.156f
C37 a_27_7# a_639_7# 0.00188f
C38 a_1462_7# a_1283_n19# 0.0074f
C39 a_27_7# VPWR 0.152f
C40 VGND Q 0.0616f
C41 Q a_1108_7# 9.8e-19
C42 VGND a_761_249# 0.0734f
C43 VGND a_805_7# 0.00579f
C44 a_1108_7# a_761_249# 0.0512f
C45 Q a_1283_n19# 0.0598f
C46 a_543_7# VGND 0.123f
C47 VPB Q 0.011f
C48 VGND RESET_B 0.288f
C49 a_1217_7# a_761_249# 4.2e-19
C50 a_543_7# a_1108_7# 7.99e-20
C51 RESET_B a_1108_7# 0.237f
C52 VPB a_761_249# 0.0994f
C53 RESET_B a_1217_7# 6.03e-19
C54 a_651_373# a_761_249# 0.0977f
C55 a_543_7# VPB 0.0958f
C56 RESET_B a_1283_n19# 0.278f
C57 a_543_7# a_448_7# 0.0498f
C58 VPB RESET_B 0.138f
C59 a_448_7# RESET_B 2.45e-19
C60 a_543_7# a_651_373# 0.0572f
C61 a_193_7# VGND 0.0631f
C62 a_651_373# RESET_B 0.0122f
C63 VGND a_639_7# 0.00863f
C64 a_193_7# a_1108_7# 0.125f
C65 a_1270_373# a_761_249# 2.6e-19
C66 a_543_7# D 7.35e-20
C67 CLK RESET_B 1.09e-19
C68 a_193_7# a_1217_7# 2.36e-20
C69 VGND VPWR 0.0502f
C70 D RESET_B 4.72e-19
C71 a_193_7# a_1283_n19# 0.0424f
C72 a_193_7# VPB 0.171f
C73 a_193_7# a_448_7# 0.0642f
C74 VPWR a_1108_7# 0.173f
C75 a_1270_373# RESET_B 2.06e-19
C76 a_448_7# a_639_7# 4.61e-19
C77 a_193_7# a_651_373# 0.0346f
C78 a_27_7# VGND 0.254f
C79 RESET_B a_1462_7# 0.00288f
C80 VPWR a_1283_n19# 0.209f
C81 a_27_7# a_1108_7# 0.102f
C82 VPB VPWR 0.216f
C83 a_448_7# VPWR 0.0681f
C84 a_193_7# CLK 7.94e-19
C85 a_193_7# D 0.218f
C86 a_27_7# a_1217_7# 2.56e-19
C87 a_651_373# VPWR 0.129f
C88 a_27_7# a_1283_n19# 0.0436f
C89 a_27_7# VPB 0.262f
C90 a_193_7# a_1270_373# 1.46e-19
C91 a_27_7# a_448_7# 0.0931f
C92 CLK VPWR 0.0174f
C93 Q RESET_B 9.12e-19
C94 a_805_7# a_761_249# 3.69e-19
C95 D VPWR 0.0812f
C96 a_27_7# a_651_373# 9.73e-19
C97 a_543_7# a_761_249# 0.21f
C98 a_1270_373# VPWR 7.19e-19
C99 RESET_B a_761_249# 0.166f
C100 a_543_7# a_805_7# 0.00171f
C101 a_27_7# CLK 0.234f
C102 a_27_7# D 0.133f
C103 RESET_B a_805_7# 0.00316f
C104 Q VNB 0.0899f
C105 VGND VNB 1.02f
C106 VPWR VNB 0.831f
C107 RESET_B VNB 0.264f
C108 D VNB 0.16f
C109 CLK VNB 0.195f
C110 VPB VNB 1.85f
C111 a_651_373# VNB 0.00469f
C112 a_448_7# VNB 0.0139f
C113 a_1108_7# VNB 0.139f
C114 a_1283_n19# VNB 0.299f
C115 a_543_7# VNB 0.158f
C116 a_761_249# VNB 0.121f
C117 a_193_7# VNB 0.274f
C118 a_27_7# VNB 0.496f
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR VPB VNB A X a_27_7#
X0 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X2 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X4 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 X A 0.0123f
C1 VGND A 0.0453f
C2 a_27_7# VPWR 0.167f
C3 VPB A 0.0335f
C4 VPWR X 0.139f
C5 VPWR VGND 0.0381f
C6 a_27_7# X 0.165f
C7 VPWR VPB 0.0438f
C8 a_27_7# VGND 0.105f
C9 a_27_7# VPB 0.0686f
C10 VPWR A 0.022f
C11 a_27_7# A 0.209f
C12 X VGND 0.115f
C13 X VPB 0.00837f
C14 VPB VGND 0.00461f
C15 VGND VNB 0.263f
C16 X VNB 0.0731f
C17 VPWR VNB 0.221f
C18 A VNB 0.148f
C19 VPB VNB 0.428f
C20 a_27_7# VNB 0.32f
.ends

.subckt sky130_fd_sc_hd__or2_2 VPWR VGND VPB VNB X A B a_121_257# a_39_257#
X0 a_121_257# B a_39_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1 X a_39_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=1 w=0.65 l=0.15
X2 VGND a_39_257# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND A a_39_257# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=1 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 VPWR a_39_257# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 X a_39_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.156 ps=1.36 w=1 l=0.15
X6 VPWR A a_121_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.156 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 a_39_257# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VPWR a_39_257# 0.0899f
C1 a_121_257# VPWR 0.00132f
C2 a_121_257# a_39_257# 0.00477f
C3 X VPWR 0.165f
C4 X a_39_257# 0.148f
C5 X a_121_257# 4.62e-19
C6 VPWR B 0.00593f
C7 B a_39_257# 0.0955f
C8 X B 1.51e-19
C9 VPWR A 0.00734f
C10 a_39_257# A 0.176f
C11 VPWR VPB 0.0714f
C12 VPB a_39_257# 0.0809f
C13 VGND VPWR 0.0475f
C14 VGND a_39_257# 0.14f
C15 a_121_257# VGND 4.62e-19
C16 X A 0.014f
C17 X VPB 0.0108f
C18 X VGND 0.0981f
C19 B A 0.0751f
C20 B VPB 0.0416f
C21 VGND B 0.0362f
C22 VPB A 0.0318f
C23 VGND A 0.0509f
C24 VGND VPB 0.00955f
C25 VGND VNB 0.323f
C26 X VNB 0.0724f
C27 A VNB 0.112f
C28 B VNB 0.178f
C29 VPWR VNB 0.284f
C30 VPB VNB 0.516f
C31 a_39_257# VNB 0.229f
.ends

.subckt sky130_fd_sc_hd__or2_1 VGND VPWR VPB VNB X A B a_68_257# a_150_257#
X0 a_68_257# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 a_150_257# B a_68_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 VGND A a_68_257# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 X a_68_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X4 VPWR A a_150_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 X a_68_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
C0 B VPB 0.0462f
C1 VPWR a_150_257# 0.00193f
C2 A X 0.0131f
C3 A VGND 0.0347f
C4 VGND X 0.114f
C5 VPWR VPB 0.0805f
C6 A a_68_257# 0.158f
C7 a_68_257# X 0.105f
C8 VPWR B 0.00855f
C9 a_68_257# VGND 0.118f
C10 X a_150_257# 4.96e-19
C11 VGND a_150_257# 4.62e-19
C12 a_68_257# a_150_257# 0.00477f
C13 A VPB 0.031f
C14 X VPB 0.0209f
C15 B A 0.0751f
C16 B X 1.65e-19
C17 VGND VPB 0.0112f
C18 B VGND 0.0437f
C19 a_68_257# VPB 0.0611f
C20 B a_68_257# 0.0984f
C21 VPWR A 0.00846f
C22 VPWR X 0.129f
C23 VPWR VGND 0.0464f
C24 VPWR a_68_257# 0.089f
C25 VGND VNB 0.32f
C26 X VNB 0.101f
C27 A VNB 0.111f
C28 B VNB 0.183f
C29 VPWR VNB 0.269f
C30 VPB VNB 0.516f
C31 a_68_257# VNB 0.154f
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND VPB VNB A2 A1 B1 Y a_199_7# a_113_257#
X0 VGND A2 a_199_7# VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X1 a_113_257# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2 a_199_7# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X4 VPWR A1 a_113_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X5 a_113_257# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
C0 VPWR VPB 0.0424f
C1 VPWR A2 0.0147f
C2 VPWR a_113_257# 0.177f
C3 a_199_7# VPWR 4.76e-19
C4 VPB A2 0.0373f
C5 a_113_257# VPB 0.0108f
C6 a_113_257# A2 0.0476f
C7 a_199_7# a_113_257# 2.42e-19
C8 VPWR B1 0.0134f
C9 VPB B1 0.0389f
C10 a_113_257# B1 0.00758f
C11 VPWR A1 0.0154f
C12 VPWR VGND 0.037f
C13 VPWR Y 0.0447f
C14 VPB A1 0.0264f
C15 A2 A1 0.0912f
C16 a_113_257# A1 0.05f
C17 VGND VPB 0.00548f
C18 VGND A2 0.0495f
C19 Y VPB 0.0146f
C20 a_199_7# A1 0.00917f
C21 a_113_257# VGND 0.00882f
C22 Y A2 0.00122f
C23 a_113_257# Y 0.0909f
C24 a_199_7# VGND 0.00428f
C25 a_199_7# Y 0.00151f
C26 B1 A1 0.0518f
C27 VGND B1 0.0436f
C28 Y B1 0.113f
C29 VGND A1 0.078f
C30 Y A1 0.0813f
C31 Y VGND 0.0654f
C32 VGND VNB 0.286f
C33 VPWR VNB 0.211f
C34 Y VNB 0.0544f
C35 A2 VNB 0.144f
C36 A1 VNB 0.0981f
C37 B1 VNB 0.162f
C38 VPB VNB 0.428f
C39 a_113_257# VNB 0.034f
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VPB VNB X A1 S A0 a_505_n19# a_535_334#
+ a_76_159# a_218_334# a_439_7# a_218_7#
X0 VPWR a_76_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1 VPWR a_505_n19# a_535_334# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 a_505_n19# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3 a_76_159# A1 a_218_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_505_n19# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X5 a_439_7# A0 a_76_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X6 a_218_334# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X7 a_76_159# A0 a_218_334# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X8 a_535_334# A1 a_76_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X9 VGND a_505_n19# a_439_7# VNB sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 VGND a_76_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_218_7# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
C0 a_439_7# A1 0.00498f
C1 a_535_334# VPWR 8.63e-19
C2 a_439_7# VPWR 4.69e-19
C3 VPWR X 0.128f
C4 a_76_159# a_535_334# 6.64e-19
C5 a_76_159# X 0.0776f
C6 a_505_n19# S 0.198f
C7 a_505_n19# VGND 0.124f
C8 a_218_7# VPWR 4.95e-19
C9 VPB a_505_n19# 0.0781f
C10 S VGND 0.033f
C11 a_218_7# a_76_159# 0.00783f
C12 VPB S 0.168f
C13 VPB VGND 0.0134f
C14 a_505_n19# A0 0.0383f
C15 a_218_7# X 2.88e-19
C16 S A0 0.0341f
C17 A0 VGND 0.0432f
C18 VPB A0 0.107f
C19 a_505_n19# A1 0.0993f
C20 a_505_n19# VPWR 0.0818f
C21 S A1 0.0872f
C22 VGND A1 0.0752f
C23 S VPWR 0.392f
C24 VPWR VGND 0.0804f
C25 a_218_334# S 0.00688f
C26 a_218_334# VGND 7.29e-19
C27 a_76_159# S 0.318f
C28 VPB A1 0.0721f
C29 a_76_159# VGND 0.16f
C30 VPB VPWR 0.11f
C31 VPB a_76_159# 0.0481f
C32 S a_535_334# 0.00526f
C33 a_535_334# VGND 6.38e-19
C34 a_439_7# VGND 0.00354f
C35 A0 A1 0.267f
C36 S X 0.00823f
C37 VGND X 0.0586f
C38 A0 VPWR 0.00732f
C39 a_76_159# A0 0.0544f
C40 VPB X 0.012f
C41 a_218_7# VGND 0.00328f
C42 a_439_7# A0 0.00369f
C43 VPWR A1 0.0114f
C44 a_76_159# A1 0.187f
C45 a_218_334# VPWR 0.00177f
C46 a_76_159# VPWR 0.0542f
C47 a_76_159# a_218_334# 0.00557f
C48 VGND VNB 0.499f
C49 A1 VNB 0.14f
C50 A0 VNB 0.134f
C51 S VNB 0.268f
C52 VPWR VNB 0.419f
C53 X VNB 0.0924f
C54 VPB VNB 0.871f
C55 a_505_n19# VNB 0.247f
C56 a_76_159# VNB 0.139f
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=4.73
C0 VGND VPWR 2.01f
C1 VGND VPB 0.336f
C2 VPWR VPB 0.142f
C3 VPWR VNB 1.69f
C4 VGND VNB 1.45f
C5 VPB VNB 1.14f
.ends

.subckt sky130_fd_sc_hd__o21ba_1 VGND VPWR VPB VNB B1_N A1 A2 X a_448_7# a_544_257#
+ a_79_159# a_222_53#
X0 VGND A2 a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1 VPWR a_79_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.186 pd=1.41 as=0.26 ps=2.52 w=1 l=0.15
X2 a_222_53# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.1 ps=0.985 w=0.42 l=0.15
X3 a_448_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VPWR A1 a_544_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X5 a_448_7# a_222_53# a_79_159# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_222_53# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.186 ps=1.41 w=0.42 l=0.15
X7 a_79_159# a_222_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X8 a_544_257# A2 a_79_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X9 VGND a_79_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPWR B1_N 0.00448f
C1 VPWR a_222_53# 0.0224f
C2 X VPB 0.0132f
C3 VGND a_544_257# 0.00166f
C4 a_79_159# X 0.11f
C5 VGND VPWR 0.0742f
C6 a_448_7# VPB 6.33e-19
C7 B1_N a_222_53# 0.106f
C8 VGND A1 0.017f
C9 a_79_159# a_448_7# 0.0461f
C10 a_79_159# VPB 0.0676f
C11 A2 a_448_7# 0.0581f
C12 A2 VPB 0.0259f
C13 VGND B1_N 0.0161f
C14 VGND a_222_53# 0.0731f
C15 A2 a_79_159# 0.0609f
C16 X VPWR 0.0729f
C17 a_448_7# a_544_257# 0.00203f
C18 VPWR a_448_7# 0.00501f
C19 VPWR VPB 0.11f
C20 A1 a_448_7# 0.0574f
C21 A1 VPB 0.0384f
C22 a_79_159# a_544_257# 0.00594f
C23 X B1_N 0.00114f
C24 a_79_159# VPWR 0.263f
C25 a_79_159# A1 0.00575f
C26 X a_222_53# 0.00374f
C27 A2 a_544_257# 0.0012f
C28 A2 VPWR 0.0227f
C29 a_448_7# B1_N 2.55e-19
C30 B1_N VPB 0.0419f
C31 A2 A1 0.0793f
C32 a_448_7# a_222_53# 0.00596f
C33 VPB a_222_53# 0.0639f
C34 a_79_159# B1_N 0.0833f
C35 VGND X 0.0609f
C36 a_79_159# a_222_53# 0.221f
C37 A2 a_222_53# 0.0562f
C38 VGND a_448_7# 0.168f
C39 VGND VPB 0.0116f
C40 VGND a_79_159# 0.0836f
C41 VPWR a_544_257# 0.0132f
C42 VGND A2 0.0157f
C43 A1 VPWR 0.0508f
C44 VGND VNB 0.468f
C45 B1_N VNB 0.105f
C46 VPWR VNB 0.4f
C47 X VNB 0.0865f
C48 A1 VNB 0.136f
C49 A2 VNB 0.0904f
C50 VPB VNB 0.782f
C51 a_448_7# VNB 0.0324f
C52 a_222_53# VNB 0.159f
C53 a_79_159# VNB 0.148f
.ends

.subckt sky130_fd_sc_hd__buf_8 VGND VPWR VPB VNB A X a_27_7#
X0 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X5 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_27_7# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 a_27_7# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X20 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
C0 a_27_7# VPB 0.266f
C1 VPWR a_27_7# 0.465f
C2 VPWR VPB 0.13f
C3 A a_27_7# 0.366f
C4 A VPB 0.0995f
C5 X VGND 0.486f
C6 A VPWR 0.0492f
C7 X a_27_7# 0.63f
C8 VGND a_27_7# 0.355f
C9 X VPB 0.0164f
C10 VPWR X 0.664f
C11 VGND VPB 0.0142f
C12 VPWR VGND 0.13f
C13 A X 6.16e-19
C14 A VGND 0.0543f
C15 VGND VNB 0.654f
C16 X VNB 0.0597f
C17 VPWR VNB 0.556f
C18 A VNB 0.322f
C19 VPB VNB 1.14f
C20 a_27_7# VNB 0.839f
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 VGND VPWR VPB VNB CLK D RESET_B Q a_639_7# a_805_7#
+ a_448_7# a_543_7# a_1283_n19# a_1462_7# a_1270_373# a_193_7# a_1217_7# a_761_249#
+ a_27_7# a_1108_7# a_651_373#
X0 VGND a_1283_n19# a_1217_7# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1 a_543_7# a_193_7# a_448_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2 VPWR a_1283_n19# a_1270_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR a_1108_7# a_1283_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1108_7# a_193_7# a_761_249# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 a_1270_373# a_193_7# a_1108_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1283_n19# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7 VGND a_1283_n19# Q VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR a_761_249# a_651_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X9 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 a_543_7# a_27_7# a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X11 VGND a_1283_n19# Q VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VPWR a_1283_n19# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X14 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_651_373# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X16 a_761_249# a_543_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X17 VGND RESET_B a_805_7# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 a_651_373# a_27_7# a_543_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X20 VPWR a_1283_n19# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 a_1217_7# a_27_7# a_1108_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X22 a_448_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X23 a_639_7# a_193_7# a_543_7# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 a_448_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_1283_n19# a_1108_7# a_1462_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X26 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X28 a_805_7# a_761_249# a_639_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X29 a_1462_7# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X30 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X31 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X32 a_1108_7# a_27_7# a_761_249# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X33 a_761_249# a_543_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
C0 RESET_B a_193_7# 0.0269f
C1 VPWR a_1108_7# 0.173f
C2 RESET_B VGND 0.288f
C3 a_761_249# VPWR 0.105f
C4 a_1462_7# a_1283_n19# 0.0074f
C5 a_1283_n19# Q 0.367f
C6 a_1217_7# a_1108_7# 0.00742f
C7 a_1270_373# VPWR 7.19e-19
C8 a_193_7# a_1108_7# 0.125f
C9 a_1217_7# a_761_249# 4.2e-19
C10 RESET_B D 4.72e-19
C11 a_761_249# a_193_7# 0.186f
C12 VGND a_1108_7# 0.148f
C13 a_1462_7# RESET_B 0.00288f
C14 RESET_B Q 0.00188f
C15 a_761_249# VGND 0.0734f
C16 a_1270_373# a_193_7# 1.46e-19
C17 a_805_7# VGND 0.00579f
C18 a_639_7# a_543_7# 0.0138f
C19 a_639_7# a_448_7# 4.61e-19
C20 Q a_1108_7# 0.0027f
C21 a_193_7# VPWR 0.396f
C22 a_27_7# a_639_7# 0.00188f
C23 VPWR VGND 0.0779f
C24 a_543_7# a_448_7# 0.0498f
C25 a_1217_7# a_193_7# 2.36e-20
C26 a_1217_7# VGND 9.68e-19
C27 VPWR D 0.0812f
C28 a_543_7# VPB 0.0958f
C29 VPB a_448_7# 0.0141f
C30 a_27_7# a_543_7# 0.115f
C31 a_27_7# a_448_7# 0.0931f
C32 a_193_7# VGND 0.0631f
C33 VPWR Q 0.368f
C34 a_651_373# a_543_7# 0.0572f
C35 a_27_7# VPB 0.262f
C36 a_193_7# D 0.218f
C37 VGND D 0.0516f
C38 a_193_7# Q 2.64e-19
C39 a_651_373# VPB 0.0135f
C40 a_651_373# a_27_7# 9.73e-19
C41 a_1462_7# VGND 0.00223f
C42 VGND Q 0.296f
C43 a_639_7# RESET_B 9.54e-19
C44 a_1283_n19# VPB 0.228f
C45 a_27_7# a_1283_n19# 0.0436f
C46 VPB CLK 0.0693f
C47 a_27_7# CLK 0.234f
C48 RESET_B a_543_7# 0.153f
C49 RESET_B a_448_7# 2.45e-19
C50 a_639_7# a_761_249# 3.16e-19
C51 RESET_B VPB 0.138f
C52 a_27_7# RESET_B 0.296f
C53 a_543_7# a_1108_7# 7.99e-20
C54 a_543_7# a_761_249# 0.21f
C55 a_805_7# a_543_7# 0.00171f
C56 a_651_373# RESET_B 0.0122f
C57 VPB a_1108_7# 0.115f
C58 a_27_7# a_1108_7# 0.102f
C59 VPB a_761_249# 0.0994f
C60 a_27_7# a_761_249# 0.0701f
C61 RESET_B a_1283_n19# 0.28f
C62 RESET_B CLK 1.09e-19
C63 a_639_7# a_193_7# 2.28e-19
C64 a_543_7# VPWR 0.1f
C65 a_448_7# VPWR 0.0681f
C66 a_651_373# a_761_249# 0.0977f
C67 a_639_7# VGND 0.00863f
C68 VPB VPWR 0.242f
C69 a_27_7# VPWR 0.152f
C70 a_1283_n19# a_1108_7# 0.234f
C71 a_543_7# a_193_7# 0.23f
C72 a_448_7# a_193_7# 0.0642f
C73 a_543_7# VGND 0.123f
C74 a_448_7# VGND 0.0661f
C75 a_27_7# a_1217_7# 2.56e-19
C76 a_651_373# VPWR 0.129f
C77 VPB a_193_7# 0.171f
C78 a_27_7# a_193_7# 0.906f
C79 RESET_B a_1108_7# 0.237f
C80 a_543_7# D 7.35e-20
C81 VPB VGND 0.0123f
C82 a_448_7# D 0.156f
C83 a_27_7# VGND 0.254f
C84 RESET_B a_761_249# 0.166f
C85 a_651_373# a_193_7# 0.0346f
C86 a_805_7# RESET_B 0.00316f
C87 a_1283_n19# VPWR 0.234f
C88 CLK VPWR 0.0174f
C89 a_1270_373# RESET_B 2.06e-19
C90 VPB D 0.138f
C91 a_27_7# D 0.133f
C92 a_761_249# a_1108_7# 0.0512f
C93 VPB Q 0.0176f
C94 a_27_7# Q 4.52e-20
C95 a_1283_n19# a_193_7# 0.0427f
C96 a_193_7# CLK 7.94e-19
C97 RESET_B VPWR 0.0652f
C98 a_1270_373# a_1108_7# 0.00645f
C99 a_805_7# a_761_249# 3.69e-19
C100 a_1283_n19# VGND 0.299f
C101 CLK VGND 0.0172f
C102 a_1270_373# a_761_249# 2.6e-19
C103 RESET_B a_1217_7# 6.03e-19
C104 Q VNB 0.0615f
C105 VGND VNB 1.18f
C106 VPWR VNB 0.977f
C107 RESET_B VNB 0.26f
C108 D VNB 0.16f
C109 CLK VNB 0.195f
C110 VPB VNB 2.11f
C111 a_651_373# VNB 0.00469f
C112 a_448_7# VNB 0.0139f
C113 a_1108_7# VNB 0.135f
C114 a_1283_n19# VNB 0.564f
C115 a_543_7# VNB 0.158f
C116 a_761_249# VNB 0.121f
C117 a_193_7# VNB 0.273f
C118 a_27_7# VNB 0.496f
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR VPB VNB X A a_27_7#
X0 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
C0 VPB VPWR 0.0355f
C1 VPB X 0.0128f
C2 A VPWR 0.0215f
C3 VGND a_27_7# 0.105f
C4 A X 8.48e-19
C5 VPWR X 0.0897f
C6 VGND VPB 0.00505f
C7 VPB a_27_7# 0.0592f
C8 VGND A 0.0184f
C9 a_27_7# A 0.181f
C10 VGND VPWR 0.029f
C11 a_27_7# VPWR 0.135f
C12 VGND X 0.0546f
C13 a_27_7# X 0.107f
C14 VPB A 0.0524f
C15 VGND VNB 0.207f
C16 X VNB 0.0941f
C17 VPWR VNB 0.175f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_27_7# VNB 0.208f
.ends

.subckt sky130_fd_sc_hd__a31o_1 VGND VPWR VPB VNB X A3 A2 A1 B1 a_209_7# a_209_257#
+ a_303_7# a_80_n19#
X0 VPWR A2 a_209_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1 a_80_n19# B1 a_209_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X2 a_209_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3 VPWR a_80_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND B1 a_80_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X5 a_209_257# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X6 VGND a_80_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X7 a_209_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X8 a_303_7# A2 a_209_7# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X9 a_80_n19# A1 a_303_7# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
C0 X A2 3.42e-19
C1 a_303_7# A2 3.38e-19
C2 VPB X 0.0108f
C3 a_209_257# A2 0.0366f
C4 VPB a_209_257# 0.00284f
C5 a_209_257# B1 0.00622f
C6 a_209_7# VPWR 0.00102f
C7 a_209_7# A3 3.56e-19
C8 VPB A2 0.0285f
C9 VPWR A3 0.0403f
C10 VPB B1 0.0342f
C11 a_80_n19# a_209_7# 0.0101f
C12 A1 VPWR 0.018f
C13 a_80_n19# VPWR 0.0992f
C14 a_80_n19# A3 0.117f
C15 a_209_7# VGND 0.00696f
C16 a_80_n19# A1 0.0367f
C17 VPWR VGND 0.0662f
C18 VGND A3 0.0169f
C19 A1 VGND 0.0135f
C20 a_209_7# X 9.76e-19
C21 a_80_n19# VGND 0.216f
C22 a_209_7# a_209_257# 6.96e-20
C23 VPWR X 0.117f
C24 X A3 0.00625f
C25 a_303_7# VPWR 0.00105f
C26 a_209_257# VPWR 0.205f
C27 a_209_257# A3 0.0268f
C28 A1 X 1.56e-19
C29 A1 a_209_257# 0.0378f
C30 a_80_n19# X 0.0765f
C31 VPWR A2 0.0227f
C32 A3 A2 0.109f
C33 a_80_n19# a_303_7# 0.0115f
C34 a_80_n19# a_209_257# 0.0626f
C35 VPB VPWR 0.0715f
C36 VPB A3 0.0297f
C37 VPWR B1 0.0177f
C38 A1 A2 0.104f
C39 VGND X 0.0572f
C40 a_303_7# VGND 0.00661f
C41 VPB A1 0.0287f
C42 a_209_257# VGND 0.0043f
C43 A1 B1 0.101f
C44 a_80_n19# A2 0.0357f
C45 VPB a_80_n19# 0.051f
C46 a_80_n19# B1 0.111f
C47 VGND A2 0.0148f
C48 VPB VGND 0.00769f
C49 VGND B1 0.0172f
C50 a_303_7# X 6.01e-19
C51 a_209_257# a_303_7# 1.26e-19
C52 VGND VNB 0.41f
C53 VPWR VNB 0.332f
C54 X VNB 0.0895f
C55 B1 VNB 0.115f
C56 A1 VNB 0.0897f
C57 A2 VNB 0.0896f
C58 A3 VNB 0.0899f
C59 VPB VNB 0.693f
C60 a_209_257# VNB 0.00621f
C61 a_80_n19# VNB 0.211f
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR VPB VNB CLK D RESET_B Q a_639_7# a_805_7#
+ a_448_7# a_543_7# a_1283_n19# a_1462_7# a_1270_373# a_193_7# a_1217_7# a_761_249#
+ a_27_7# a_1108_7# a_651_373#
X0 VGND a_1283_n19# a_1217_7# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1 a_543_7# a_193_7# a_448_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2 VPWR a_1283_n19# a_1270_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR a_1108_7# a_1283_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_1108_7# a_193_7# a_761_249# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 a_1270_373# a_193_7# a_1108_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 a_1283_n19# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X7 VPWR a_761_249# a_651_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X8 a_543_7# a_27_7# a_448_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X9 VPWR a_1283_n19# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 Q a_1283_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X11 VPWR CLK a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X12 a_193_7# a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_651_373# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X14 a_761_249# a_543_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X15 VGND RESET_B a_805_7# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X16 a_651_373# a_27_7# a_543_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X17 a_1217_7# a_27_7# a_1108_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X18 a_448_7# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X19 a_639_7# a_193_7# a_543_7# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X20 Q a_1283_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X21 VGND a_1283_n19# Q VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 a_448_7# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X23 a_1283_n19# a_1108_7# a_1462_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X24 VGND CLK a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X25 a_805_7# a_761_249# a_639_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X26 a_1462_7# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X27 a_193_7# a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X28 a_1108_7# a_27_7# a_761_249# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X29 a_761_249# a_543_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
C0 a_27_7# a_448_7# 0.0931f
C1 a_1270_373# a_1108_7# 0.00645f
C2 VPB a_448_7# 0.0141f
C3 a_543_7# a_27_7# 0.115f
C4 a_639_7# a_448_7# 4.61e-19
C5 VGND a_27_7# 0.254f
C6 VPB a_543_7# 0.0958f
C7 VGND VPB 0.0122f
C8 a_639_7# a_543_7# 0.0138f
C9 RESET_B a_27_7# 0.296f
C10 a_639_7# VGND 0.00863f
C11 a_543_7# a_761_249# 0.21f
C12 RESET_B VPB 0.138f
C13 VGND a_761_249# 0.0734f
C14 a_639_7# RESET_B 9.54e-19
C15 RESET_B a_761_249# 0.166f
C16 VPWR a_1283_n19# 0.23f
C17 a_651_373# VPWR 0.129f
C18 VPB a_27_7# 0.262f
C19 a_639_7# a_27_7# 0.00188f
C20 a_761_249# a_27_7# 0.0701f
C21 a_193_7# VPWR 0.396f
C22 VPB a_761_249# 0.0994f
C23 a_1270_373# RESET_B 2.06e-19
C24 a_639_7# a_761_249# 3.16e-19
C25 D VPWR 0.0812f
C26 a_193_7# a_1283_n19# 0.0425f
C27 VPWR Q 0.169f
C28 a_651_373# a_193_7# 0.0346f
C29 a_193_7# a_1217_7# 2.36e-20
C30 VPWR a_1108_7# 0.174f
C31 Q a_1283_n19# 0.0963f
C32 a_1270_373# a_761_249# 2.6e-19
C33 D a_193_7# 0.218f
C34 a_1283_n19# a_1108_7# 0.234f
C35 a_1283_n19# a_1462_7# 0.0074f
C36 a_193_7# Q 1.79e-19
C37 VPWR CLK 0.0174f
C38 a_1108_7# a_1217_7# 0.00742f
C39 a_193_7# a_1108_7# 0.125f
C40 VPWR a_448_7# 0.0681f
C41 VPWR a_543_7# 0.1f
C42 VPWR VGND 0.0719f
C43 Q a_1108_7# 9.64e-19
C44 a_193_7# CLK 7.94e-19
C45 VPWR RESET_B 0.0652f
C46 a_543_7# a_805_7# 0.00171f
C47 VGND a_1283_n19# 0.259f
C48 VGND a_805_7# 0.00579f
C49 a_651_373# a_543_7# 0.0572f
C50 RESET_B a_1283_n19# 0.279f
C51 a_193_7# a_448_7# 0.0642f
C52 RESET_B a_805_7# 0.00316f
C53 VPWR a_27_7# 0.152f
C54 a_651_373# RESET_B 0.0122f
C55 a_193_7# a_543_7# 0.23f
C56 VGND a_1217_7# 9.68e-19
C57 VPWR VPB 0.234f
C58 a_193_7# VGND 0.0631f
C59 D a_448_7# 0.156f
C60 RESET_B a_1217_7# 6.03e-19
C61 a_193_7# RESET_B 0.0269f
C62 VPWR a_761_249# 0.105f
C63 D a_543_7# 7.35e-20
C64 a_1283_n19# a_27_7# 0.0436f
C65 D VGND 0.0516f
C66 a_651_373# a_27_7# 9.73e-19
C67 a_1283_n19# VPB 0.168f
C68 D RESET_B 4.72e-19
C69 VGND Q 0.11f
C70 a_651_373# VPB 0.0135f
C71 a_805_7# a_761_249# 3.69e-19
C72 RESET_B Q 8.96e-19
C73 a_1217_7# a_27_7# 2.56e-19
C74 a_193_7# a_27_7# 0.906f
C75 a_651_373# a_761_249# 0.0977f
C76 a_1108_7# a_543_7# 7.99e-20
C77 VGND a_1108_7# 0.148f
C78 a_193_7# VPB 0.171f
C79 VGND a_1462_7# 0.00221f
C80 a_1270_373# VPWR 7.19e-19
C81 a_639_7# a_193_7# 2.28e-19
C82 RESET_B a_1108_7# 0.237f
C83 a_1217_7# a_761_249# 4.2e-19
C84 RESET_B a_1462_7# 0.00288f
C85 a_193_7# a_761_249# 0.186f
C86 D a_27_7# 0.133f
C87 D VPB 0.138f
C88 Q a_27_7# 2.57e-20
C89 Q VPB 0.00555f
C90 VGND CLK 0.0172f
C91 RESET_B CLK 1.09e-19
C92 a_1108_7# a_27_7# 0.102f
C93 a_1108_7# VPB 0.115f
C94 a_543_7# a_448_7# 0.0498f
C95 a_1270_373# a_193_7# 1.46e-19
C96 VGND a_448_7# 0.0661f
C97 a_1108_7# a_761_249# 0.0512f
C98 RESET_B a_448_7# 2.45e-19
C99 VGND a_543_7# 0.123f
C100 CLK a_27_7# 0.234f
C101 RESET_B a_543_7# 0.153f
C102 CLK VPB 0.0693f
C103 RESET_B VGND 0.288f
C104 Q VNB 0.0296f
C105 VGND VNB 1.1f
C106 VPWR VNB 0.902f
C107 RESET_B VNB 0.263f
C108 D VNB 0.16f
C109 CLK VNB 0.195f
C110 VPB VNB 1.93f
C111 a_651_373# VNB 0.00469f
C112 a_448_7# VNB 0.0139f
C113 a_1108_7# VNB 0.137f
C114 a_1283_n19# VNB 0.389f
C115 a_543_7# VNB 0.158f
C116 a_761_249# VNB 0.121f
C117 a_193_7# VNB 0.273f
C118 a_27_7# VNB 0.496f
.ends

.subckt sky130_fd_sc_hd__or3_2 VGND VPWR VPB VNB B C A X a_184_257# a_112_257# a_30_13#
X0 VPWR A a_184_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1 a_184_257# B a_112_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 X a_30_13# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X3 VPWR a_30_13# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND a_30_13# X VNB sky130_fd_pr__nfet_01v8 ad=0.185 pd=1.87 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 X a_30_13# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.148 ps=1.34 w=1 l=0.15
X6 a_112_257# C a_30_13# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_30_13# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_30_13# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VGND C a_30_13# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
C0 A VPWR 0.00982f
C1 VPB B 0.0972f
C2 VPB a_30_13# 0.0791f
C3 X VPB 0.00385f
C4 A a_112_257# 0.00223f
C5 a_30_13# B 0.121f
C6 X B 6.52e-19
C7 X a_30_13# 0.137f
C8 A VPB 0.0382f
C9 C VGND 0.0163f
C10 A B 0.0788f
C11 a_184_257# VGND 5.47e-19
C12 A a_30_13# 0.244f
C13 A X 0.00129f
C14 VPWR VGND 0.0712f
C15 C VPWR 0.00459f
C16 a_184_257# VPWR 7.72e-19
C17 a_112_257# VGND 3.96e-19
C18 VPB VGND 0.00844f
C19 C VPB 0.0399f
C20 a_112_257# VPWR 5.94e-19
C21 VGND B 0.0151f
C22 C B 0.0802f
C23 a_30_13# VGND 0.236f
C24 VPB VPWR 0.0818f
C25 X VGND 0.0786f
C26 C a_30_13# 0.0862f
C27 VPWR B 0.148f
C28 a_184_257# a_30_13# 0.00863f
C29 VPWR a_30_13# 0.101f
C30 A VGND 0.0192f
C31 X VPWR 0.176f
C32 A C 0.0343f
C33 A a_184_257# 0.00228f
C34 a_112_257# a_30_13# 0.00501f
C35 VGND VNB 0.38f
C36 X VNB 0.0245f
C37 A VNB 0.117f
C38 C VNB 0.161f
C39 B VNB 0.116f
C40 VPWR VNB 0.33f
C41 VPB VNB 0.605f
C42 a_30_13# VNB 0.267f
.ends

.subckt sky130_fd_sc_hd__o21a_1 VGND VPWR VPB VNB A1 A2 B1 X a_382_257# a_79_n19#
+ a_297_7#
X0 a_297_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_79_n19# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X2 a_382_257# A2 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X3 VPWR A1 a_382_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X4 a_297_7# B1 a_79_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X7 VGND A2 a_297_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
C0 A1 A2 0.102f
C1 VPB B1 0.0328f
C2 a_297_7# A2 0.048f
C3 VGND A2 0.0171f
C4 B1 A2 0.0665f
C5 a_297_7# A1 0.0492f
C6 a_382_257# A2 0.0145f
C7 VGND A1 0.0157f
C8 VGND X 0.0736f
C9 a_297_7# VGND 0.125f
C10 B1 X 3.56e-19
C11 a_79_n19# VPWR 0.201f
C12 a_382_257# A1 2.25e-19
C13 a_297_7# B1 0.00637f
C14 VGND B1 0.0182f
C15 a_382_257# a_297_7# 8.13e-19
C16 a_382_257# VGND 8.23e-19
C17 a_79_n19# VPB 0.0489f
C18 VPWR VPB 0.0624f
C19 a_79_n19# A2 0.0889f
C20 VPWR A2 0.0835f
C21 a_79_n19# A1 7.71e-19
C22 a_79_n19# X 0.104f
C23 VPWR A1 0.0449f
C24 VPB A2 0.0334f
C25 a_297_7# a_79_n19# 0.0326f
C26 VPWR X 0.0958f
C27 a_79_n19# VGND 0.129f
C28 a_297_7# VPWR 0.0056f
C29 VPWR VGND 0.0588f
C30 a_79_n19# B1 0.134f
C31 VPB A1 0.0412f
C32 a_382_257# a_79_n19# 0.00145f
C33 VPWR B1 0.0213f
C34 VPB X 0.011f
C35 a_382_257# VPWR 0.00566f
C36 a_297_7# VPB 7.6e-19
C37 VGND VPB 0.0049f
C38 VGND VNB 0.352f
C39 VPWR VNB 0.304f
C40 X VNB 0.0935f
C41 A1 VNB 0.152f
C42 A2 VNB 0.0981f
C43 B1 VNB 0.101f
C44 VPB VNB 0.605f
C45 a_297_7# VNB 0.0348f
C46 a_79_n19# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VPB VNB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.452 ps=4.52 w=0.87 l=0.59
C0 VPWR VGND 0.353f
C1 VPB VPWR 0.0625f
C2 VPB VGND 0.0797f
C3 VPWR VNB 0.47f
C4 VGND VNB 0.427f
C5 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__nor2_1 VGND VPWR VPB VNB A B Y a_109_257#
X0 a_109_257# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 VPWR A a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VPWR a_109_257# 0.00638f
C1 B VPB 0.0367f
C2 VPWR VPB 0.0449f
C3 A Y 0.0471f
C4 A VGND 0.0486f
C5 A B 0.0584f
C6 VPWR A 0.0528f
C7 Y VGND 0.154f
C8 A VPB 0.0415f
C9 Y B 0.0877f
C10 B VGND 0.0451f
C11 VPWR Y 0.0995f
C12 VPWR VGND 0.0314f
C13 Y a_109_257# 0.0113f
C14 VGND a_109_257# 0.00128f
C15 Y VPB 0.0139f
C16 VPB VGND 0.00456f
C17 VPWR B 0.0148f
C18 VGND VNB 0.263f
C19 VPWR VNB 0.214f
C20 Y VNB 0.0605f
C21 A VNB 0.149f
C22 B VNB 0.143f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__a2bb2oi_1 VGND VPWR VPB VNB Y A2_N A1_N B2 B1 a_109_257#
+ a_397_257# a_109_7# a_481_7#
X0 a_109_257# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A2_N a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.283 pd=1.52 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 Y a_109_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.283 ps=1.52 w=0.65 l=0.15
X3 a_109_7# A2_N a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4 a_397_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_481_7# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND B1 a_481_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR B2 a_397_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_397_257# a_109_7# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.34 ps=2.68 w=1 l=0.15
X9 a_109_7# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_109_7# a_109_257# 0.00765f
C1 Y B2 0.0778f
C2 Y a_109_7# 0.192f
C3 a_481_7# a_397_257# 4.76e-19
C4 VGND a_397_257# 0.00847f
C5 VGND B1 0.0479f
C6 VPB A2_N 0.0308f
C7 VPWR VPB 0.0778f
C8 Y a_397_257# 0.0601f
C9 VPB A1_N 0.0331f
C10 VGND a_481_7# 0.00561f
C11 Y B1 0.00112f
C12 VPWR A2_N 0.0192f
C13 A2_N A1_N 0.0842f
C14 VPWR A1_N 0.0498f
C15 VGND a_109_257# 0.00196f
C16 VPB B2 0.0272f
C17 VPB a_109_7# 0.0663f
C18 Y a_481_7# 0.00154f
C19 Y VGND 0.0978f
C20 A2_N a_109_7# 0.147f
C21 VPWR B2 0.0184f
C22 VPWR a_109_7# 0.0963f
C23 A1_N a_109_7# 0.0213f
C24 VPB a_397_257# 0.00776f
C25 VPB B1 0.035f
C26 VPWR a_397_257# 0.174f
C27 B2 a_109_7# 0.0577f
C28 VPWR B1 0.018f
C29 VGND VPB 0.00833f
C30 VGND A2_N 0.0187f
C31 VPWR a_481_7# 6.39e-19
C32 B2 a_397_257# 0.0458f
C33 a_109_7# a_397_257# 0.00647f
C34 VGND VPWR 0.0681f
C35 B1 B2 0.118f
C36 VGND A1_N 0.0492f
C37 Y VPB 0.0105f
C38 A2_N a_109_257# 5.93e-19
C39 VPWR a_109_257# 0.00889f
C40 Y A2_N 5.53e-19
C41 Y VPWR 0.0595f
C42 A1_N a_109_257# 8.3e-19
C43 B2 a_481_7# 0.00732f
C44 VGND B2 0.0678f
C45 VGND a_109_7# 0.185f
C46 B1 a_397_257# 0.0427f
C47 VGND VNB 0.438f
C48 Y VNB 0.0102f
C49 VPWR VNB 0.354f
C50 B1 VNB 0.145f
C51 B2 VNB 0.0969f
C52 A2_N VNB 0.0969f
C53 A1_N VNB 0.141f
C54 VPB VNB 0.693f
C55 a_397_257# VNB 0.0287f
C56 a_109_7# VNB 0.148f
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR VPB VNB X A a_75_172#
X0 a_75_172# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1 VPWR a_75_172# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2 VGND a_75_172# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3 a_75_172# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
C0 X VGND 0.0545f
C1 a_75_172# VPWR 0.134f
C2 VPB a_75_172# 0.0571f
C3 VPB VPWR 0.0355f
C4 A VGND 0.0184f
C5 A X 8.48e-19
C6 a_75_172# VGND 0.105f
C7 VPWR VGND 0.0289f
C8 VPB VGND 0.00507f
C9 X a_75_172# 0.107f
C10 X VPWR 0.0896f
C11 X VPB 0.0128f
C12 A a_75_172# 0.178f
C13 A VPWR 0.0217f
C14 A VPB 0.0525f
C15 VGND VNB 0.207f
C16 VPWR VNB 0.176f
C17 X VNB 0.0942f
C18 A VNB 0.164f
C19 VPB VNB 0.339f
C20 a_75_172# VNB 0.21f
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND VPB VNB B1 A1 A2 X B2 a_27_257# a_109_257#
+ a_373_7# a_109_7#
X0 VGND A2 a_373_7# VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1 a_109_257# B2 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR A2 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3 X a_27_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X4 X a_27_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X5 a_109_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X6 a_27_257# B1 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_7# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_27_257# B1 a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X9 a_373_7# A1 a_27_257# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
C0 B1 a_27_257# 0.0838f
C1 B2 a_27_257# 0.0567f
C2 VPWR B1 0.0139f
C3 VPWR B2 0.0126f
C4 X a_109_257# 0.00169f
C5 X A1 2.98e-19
C6 a_27_257# a_109_257# 0.171f
C7 VPWR a_109_257# 0.187f
C8 A1 a_27_257# 0.0839f
C9 VPWR A1 0.0168f
C10 A2 VGND 0.0162f
C11 VPB VGND 0.00746f
C12 A2 VPB 0.0284f
C13 a_109_7# a_27_257# 0.00393f
C14 X a_27_257# 0.108f
C15 a_373_7# VGND 0.00344f
C16 VPWR a_109_7# 0.00104f
C17 A2 a_373_7# 6.81e-19
C18 VPWR X 0.0914f
C19 B1 VGND 0.0267f
C20 VGND B2 0.0538f
C21 A2 B1 1.81e-19
C22 A2 B2 8.94e-20
C23 VPWR a_27_257# 0.13f
C24 B1 VPB 0.0317f
C25 VPB B2 0.0299f
C26 VGND a_109_257# 0.00426f
C27 A2 a_109_257# 0.00625f
C28 B1 B2 0.0739f
C29 A1 VGND 0.0137f
C30 A2 A1 0.0738f
C31 VPB a_109_257# 0.00882f
C32 A1 VPB 0.0387f
C33 a_373_7# A1 0.00122f
C34 a_109_7# VGND 0.00792f
C35 X VGND 0.0543f
C36 B1 a_109_257# 0.0106f
C37 B2 a_109_257# 0.0015f
C38 X A2 0.0011f
C39 A1 B1 0.0657f
C40 X VPB 0.011f
C41 VGND a_27_257# 0.257f
C42 X a_373_7# 1.97e-19
C43 A2 a_27_257# 0.161f
C44 VPWR VGND 0.0641f
C45 VPWR A2 0.0178f
C46 VPB a_27_257# 0.0591f
C47 B1 a_109_7# 0.00145f
C48 a_109_7# B2 4.58e-19
C49 VPWR VPB 0.0714f
C50 X B1 8.38e-20
C51 X B2 3.26e-20
C52 A1 a_109_257# 0.0105f
C53 a_373_7# a_27_257# 0.0134f
C54 VPWR a_373_7# 7.36e-19
C55 VGND VNB 0.421f
C56 X VNB 0.0917f
C57 VPWR VNB 0.328f
C58 A2 VNB 0.0927f
C59 A1 VNB 0.112f
C60 B1 VNB 0.112f
C61 B2 VNB 0.126f
C62 VPB VNB 0.693f
C63 a_109_257# VNB 0.00274f
C64 a_27_257# VNB 0.19f
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VGND VPWR VPB VNB A X a_110_7#
X0 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VPWR A a_110_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X11 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X12 a_110_7# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X13 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VGND A a_110_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 a_110_7# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X20 VGND A a_110_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X21 a_110_7# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X22 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X25 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X26 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X27 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X29 VPWR a_110_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X30 VPWR A a_110_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X34 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X35 VGND a_110_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 a_110_7# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X39 X a_110_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
C0 VPB a_110_7# 0.528f
C1 VPB VGND 0.0114f
C2 A X 0.00292f
C3 VPB X 0.0315f
C4 VPB A 0.133f
C5 a_110_7# VPWR 0.67f
C6 VPWR VGND 0.187f
C7 a_110_7# VGND 0.512f
C8 VPWR X 1.36f
C9 A VPWR 0.112f
C10 VPB VPWR 0.184f
C11 a_110_7# X 1.62f
C12 VGND X 0.977f
C13 A a_110_7# 0.307f
C14 A VGND 0.115f
C15 VGND VNB 1.01f
C16 X VNB 0.111f
C17 VPWR VNB 0.835f
C18 A VNB 0.495f
C19 VPB VNB 1.85f
C20 a_110_7# VNB 1.73f
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR VPB VNB A2 B1 Y A1 a_109_257# a_27_7#
X0 a_109_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1 Y A2 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X3 VGND A1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4 a_27_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X5 Y B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 VPWR a_109_257# 0.00401f
C1 a_109_257# a_27_7# 5.37e-19
C2 VGND A1 0.0163f
C3 Y a_109_257# 5.24e-19
C4 A1 A2 0.0986f
C5 VGND A2 0.0183f
C6 A1 VPWR 0.0497f
C7 VGND VPWR 0.0381f
C8 VGND B1 0.016f
C9 VPWR A2 0.109f
C10 A2 B1 0.0472f
C11 A1 a_27_7# 0.037f
C12 A1 Y 8.9e-19
C13 A1 VPB 0.0327f
C14 VGND a_27_7# 0.142f
C15 VPWR B1 0.0433f
C16 VGND Y 0.0289f
C17 A2 a_27_7# 0.0388f
C18 VGND VPB 0.00462f
C19 Y A2 0.124f
C20 VPB A2 0.0305f
C21 VPWR a_27_7# 0.00663f
C22 B1 a_27_7# 0.00471f
C23 Y VPWR 0.105f
C24 Y B1 0.0811f
C25 VPB VPWR 0.056f
C26 VPB B1 0.0741f
C27 VGND a_109_257# 4.56e-19
C28 A2 a_109_257# 0.00993f
C29 Y a_27_7# 0.0517f
C30 VPB a_27_7# 8.4e-19
C31 VPB Y 0.00672f
C32 VGND VNB 0.254f
C33 Y VNB 0.0545f
C34 VPWR VNB 0.271f
C35 B1 VNB 0.152f
C36 A2 VNB 0.0962f
C37 A1 VNB 0.138f
C38 VPB VNB 0.428f
C39 a_27_7# VNB 0.0311f
.ends

.subckt sky130_fd_sc_hd__o221ai_4 VGND VPWR VPB VNB B2 Y A2 A1 B1 C1 a_553_257# a_1241_257#
+ a_471_7# a_27_7#
X0 a_1241_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_471_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2 a_553_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Y A2 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_27_7# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.395 pd=1.79 as=0.135 ps=1.27 w=1 l=0.15
X6 Y C1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_27_7# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A1 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X10 a_27_7# B1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_471_7# B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_471_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_1241_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X16 a_471_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 VPWR B1 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND A2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_553_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.395 ps=1.79 w=1 l=0.15
X20 a_471_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND A1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 Y C1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X23 a_1241_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 a_27_7# B2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VPWR B1 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X26 VPWR A1 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_471_7# B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 Y B2 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X30 a_553_257# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 a_1241_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 a_27_7# B1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 a_471_7# B2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X34 a_27_7# B2 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 VGND A1 a_471_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X36 Y A2 a_1241_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_553_257# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 a_471_7# B2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 Y B2 a_553_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
C0 a_553_257# B1 0.0481f
C1 VPB B2 0.114f
C2 C1 B1 0.0183f
C3 a_471_7# a_553_257# 7.04e-20
C4 a_471_7# C1 8.47e-20
C5 a_1241_257# VPB 0.00652f
C6 A1 B2 5.11e-19
C7 VPWR VPB 0.196f
C8 a_1241_257# A1 0.154f
C9 VPWR A1 0.111f
C10 B1 B2 0.254f
C11 A1 VPB 0.133f
C12 a_27_7# Y 0.176f
C13 a_471_7# B2 0.0835f
C14 a_1241_257# B1 9.99e-19
C15 Y VGND 0.0339f
C16 VPWR B1 0.0731f
C17 a_471_7# VPWR 0.0133f
C18 A2 Y 0.0321f
C19 VPB B1 0.129f
C20 a_27_7# VGND 0.598f
C21 a_471_7# VPB 0.00266f
C22 A1 B1 0.093f
C23 Y a_553_257# 0.286f
C24 Y C1 0.324f
C25 a_471_7# A1 0.214f
C26 A2 VGND 0.0584f
C27 a_27_7# C1 0.0594f
C28 a_471_7# B1 0.215f
C29 a_553_257# VGND 0.00615f
C30 VGND C1 0.0373f
C31 Y B2 0.0466f
C32 A2 a_553_257# 3e-20
C33 Y a_1241_257# 0.172f
C34 Y VPWR 0.498f
C35 a_27_7# B2 0.0264f
C36 a_553_257# C1 3.36e-19
C37 VGND B2 0.0278f
C38 Y VPB 0.0189f
C39 a_27_7# VPWR 0.00762f
C40 a_1241_257# VGND 0.00647f
C41 Y A1 0.161f
C42 A2 B2 5.76e-19
C43 VPWR VGND 0.188f
C44 a_27_7# VPB 3.53e-19
C45 A2 a_1241_257# 0.0414f
C46 A2 VPWR 0.0341f
C47 VGND VPB 0.0124f
C48 a_553_257# B2 0.035f
C49 Y B1 0.36f
C50 A1 VGND 0.0628f
C51 a_1241_257# a_553_257# 6.98e-19
C52 a_471_7# Y 0.0206f
C53 A2 VPB 0.115f
C54 VPWR a_553_257# 0.409f
C55 VPWR C1 0.112f
C56 A2 A1 0.291f
C57 a_27_7# B1 0.0242f
C58 a_553_257# VPB 0.00497f
C59 C1 VPB 0.131f
C60 a_471_7# a_27_7# 0.33f
C61 VGND B1 0.0414f
C62 a_553_257# A1 2.35e-20
C63 a_471_7# VGND 0.591f
C64 a_1241_257# B2 1.52e-19
C65 A2 B1 3.11e-19
C66 VPWR B2 0.0281f
C67 a_471_7# A2 0.182f
C68 VPWR a_1241_257# 0.465f
C69 VGND VNB 1.03f
C70 Y VNB 0.0292f
C71 VPWR VNB 0.917f
C72 A2 VNB 0.352f
C73 A1 VNB 0.403f
C74 B2 VNB 0.351f
C75 B1 VNB 0.373f
C76 C1 VNB 0.41f
C77 VPB VNB 1.93f
C78 a_471_7# VNB 0.0538f
C79 a_27_7# VNB 0.0485f
C80 a_553_257# VNB 0.00146f
.ends

.subckt sky130_fd_sc_hd__mux2_2 VGND VPWR VPB VNB S A1 A0 X a_257_159# a_306_329#
+ a_79_n19# a_578_7# a_591_329# a_288_7#
X0 a_288_7# a_257_159# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.097 ps=0.975 w=0.42 l=0.15
X1 X a_79_n19# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 a_257_159# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.173 pd=1.82 as=0.0864 ps=0.91 w=0.64 l=0.15
X3 VPWR S a_591_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.0672 ps=0.85 w=0.64 l=0.15
X4 a_591_329# A0 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.85 as=0.131 ps=1.05 w=0.64 l=0.15
X5 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND S a_578_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0578 ps=0.695 w=0.42 l=0.15
X7 a_257_159# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_79_n19# A1 a_306_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.05 as=0.229 ps=1.36 w=0.64 l=0.15
X9 a_578_7# A1 a_79_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.173 ps=1.25 w=0.42 l=0.15
X10 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.41 as=0.135 ps=1.27 w=1 l=0.15
X11 X a_79_n19# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_79_n19# A0 a_288_7# VNB sky130_fd_pr__nfet_01v8 ad=0.173 pd=1.25 as=0.0683 ps=0.745 w=0.42 l=0.15
X13 a_306_329# a_257_159# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.36 as=0.178 ps=1.41 w=0.64 l=0.15
C0 VPB a_79_n19# 0.0731f
C1 VGND a_257_159# 0.0996f
C2 S VPB 0.0987f
C3 A1 VGND 0.0497f
C4 a_306_329# a_257_159# 0.0102f
C5 VPWR a_257_159# 0.149f
C6 a_288_7# VGND 0.00186f
C7 VPWR A1 0.00994f
C8 VPWR a_288_7# 3.13e-19
C9 a_79_n19# a_257_159# 0.285f
C10 a_306_329# VGND 0.00149f
C11 VPWR VGND 0.0922f
C12 S a_257_159# 0.146f
C13 A1 a_79_n19# 0.0307f
C14 a_288_7# a_79_n19# 0.00727f
C15 VPWR a_306_329# 0.00634f
C16 S A1 0.0662f
C17 VGND a_79_n19# 0.231f
C18 S VGND 0.0569f
C19 a_306_329# a_79_n19# 0.021f
C20 VPWR a_79_n19# 0.25f
C21 S VPWR 0.033f
C22 VPB X 0.00457f
C23 A0 VPB 0.0729f
C24 S a_79_n19# 0.00187f
C25 a_578_7# a_257_159# 4.09e-19
C26 a_578_7# A1 0.00429f
C27 X a_257_159# 0.00258f
C28 A0 a_257_159# 0.159f
C29 A0 A1 0.158f
C30 a_578_7# VGND 0.00424f
C31 VPWR a_578_7# 4.32e-19
C32 a_591_329# a_257_159# 0.00548f
C33 X VGND 0.109f
C34 A0 VGND 0.0185f
C35 VPWR X 0.149f
C36 VPB a_257_159# 0.108f
C37 VPWR A0 0.0177f
C38 a_578_7# a_79_n19# 9.96e-19
C39 A1 VPB 0.0585f
C40 a_591_329# VGND 6.57e-19
C41 X a_79_n19# 0.168f
C42 VPWR a_591_329# 0.00489f
C43 A0 a_79_n19# 0.0671f
C44 VPB VGND 0.011f
C45 S A0 0.0842f
C46 VPWR VPB 0.0953f
C47 A1 a_257_159# 0.0371f
C48 a_591_329# a_79_n19# 0.0015f
C49 a_288_7# a_257_159# 4.59e-19
C50 a_288_7# A1 3.38e-19
C51 VGND VNB 0.516f
C52 X VNB 0.0244f
C53 VPWR VNB 0.441f
C54 S VNB 0.244f
C55 A0 VNB 0.129f
C56 A1 VNB 0.162f
C57 VPB VNB 0.871f
C58 a_257_159# VNB 0.216f
C59 a_79_n19# VNB 0.227f
.ends

.subckt sky130_fd_sc_hd__o211a_1 VGND VPWR VPB VNB X A1 A2 B1 C1 a_510_7# a_79_n19#
+ a_215_7# a_297_257#
X0 a_79_n19# C1 a_510_7# VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.114 ps=1 w=0.65 l=0.15
X1 a_297_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2 a_215_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.106 ps=0.975 w=0.65 l=0.15
X3 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4 VGND A1 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X5 a_79_n19# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X6 VPWR B1 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X7 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_510_7# B1 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X9 a_79_n19# A2 a_297_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.162 ps=1.33 w=1 l=0.15
C0 a_79_n19# A2 0.0474f
C1 VPB B1 0.0298f
C2 A1 A2 0.0693f
C3 a_510_7# a_79_n19# 0.00844f
C4 C1 B1 0.0495f
C5 VPWR VPB 0.0944f
C6 VPWR C1 0.0203f
C7 A2 B1 0.0611f
C8 C1 VPB 0.0553f
C9 a_215_7# VGND 0.226f
C10 a_510_7# B1 0.00122f
C11 VPWR A2 0.0143f
C12 a_510_7# VPWR 0.00153f
C13 X VGND 0.0993f
C14 VPB A2 0.034f
C15 VGND a_79_n19# 0.126f
C16 VGND A1 0.017f
C17 a_215_7# X 5.57e-19
C18 a_215_7# a_79_n19# 0.0458f
C19 a_215_7# A1 0.0493f
C20 VGND B1 0.0186f
C21 X a_79_n19# 0.0491f
C22 X A1 3.68e-19
C23 VGND a_297_257# 0.002f
C24 VGND VPWR 0.0732f
C25 a_215_7# B1 0.00549f
C26 a_79_n19# A1 0.0844f
C27 a_215_7# a_297_257# 1.98e-20
C28 VGND VPB 0.0108f
C29 a_215_7# VPWR 0.00318f
C30 VGND C1 0.0133f
C31 X B1 1.2e-19
C32 a_215_7# VPB 9.29e-19
C33 X VPWR 0.129f
C34 a_79_n19# B1 0.0649f
C35 VGND A2 0.0159f
C36 a_297_257# a_79_n19# 0.0174f
C37 a_297_257# A1 6.93e-20
C38 a_510_7# VGND 0.00833f
C39 X VPB 0.0125f
C40 VPWR a_79_n19# 0.361f
C41 VPWR A1 0.0184f
C42 a_215_7# A2 0.0461f
C43 a_79_n19# VPB 0.0755f
C44 A1 VPB 0.0322f
C45 a_510_7# a_215_7# 0.00529f
C46 a_79_n19# C1 0.0965f
C47 X A2 2.44e-19
C48 VPWR B1 0.0185f
C49 VPWR a_297_257# 0.0107f
C50 VGND VNB 0.45f
C51 VPWR VNB 0.377f
C52 X VNB 0.0951f
C53 C1 VNB 0.167f
C54 B1 VNB 0.095f
C55 A2 VNB 0.101f
C56 A1 VNB 0.0989f
C57 VPB VNB 0.782f
C58 a_215_7# VNB 0.0101f
C59 a_79_n19# VNB 0.225f
.ends

.subckt sky130_fd_sc_hd__o22a_1 VGND VPWR VPB VNB B2 A2 A1 B1 X a_78_159# a_493_257#
+ a_292_257# a_215_7#
X0 a_292_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X1 a_78_159# B1 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_215_7# B2 a_78_159# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR A1 a_493_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4 VGND A2 a_215_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X5 a_215_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 a_493_257# A2 a_78_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X7 VGND a_78_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VPWR a_78_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X9 a_78_159# B2 a_292_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
C0 B2 a_78_159# 0.0816f
C1 B1 a_78_159# 0.148f
C2 X B2 1.65e-19
C3 X B1 6.11e-19
C4 VPWR a_292_257# 0.00854f
C5 A2 a_493_257# 0.0105f
C6 VPWR A2 0.12f
C7 a_78_159# a_292_257# 0.013f
C8 X a_292_257# 4.46e-19
C9 A2 a_78_159# 0.0707f
C10 VPWR a_493_257# 0.00283f
C11 A1 VGND 0.0146f
C12 VPB VGND 0.00596f
C13 A1 VPB 0.0319f
C14 a_493_257# a_78_159# 3.15e-19
C15 VPWR a_78_159# 0.211f
C16 a_215_7# VGND 0.258f
C17 A1 a_215_7# 0.0498f
C18 X VPWR 0.0911f
C19 a_215_7# VPB 9.85e-19
C20 B2 VGND 0.0103f
C21 VGND B1 0.0119f
C22 X a_78_159# 0.105f
C23 B2 VPB 0.0281f
C24 VPB B1 0.0388f
C25 a_215_7# B2 0.0207f
C26 a_215_7# B1 0.00758f
C27 VGND a_292_257# 0.00136f
C28 B2 B1 0.0815f
C29 A2 VGND 0.0153f
C30 A1 A2 0.0879f
C31 A2 VPB 0.0341f
C32 a_215_7# A2 0.0439f
C33 a_493_257# VGND 3.15e-19
C34 VPWR VGND 0.0668f
C35 A1 a_493_257# 9.88e-20
C36 B2 a_292_257# 4.98e-20
C37 VPWR A1 0.057f
C38 A2 B2 0.0676f
C39 A2 B1 3.91e-19
C40 VPWR VPB 0.0744f
C41 a_215_7# a_493_257# 3.25e-19
C42 VGND a_78_159# 0.0684f
C43 VPWR a_215_7# 0.00435f
C44 A1 a_78_159# 4.58e-19
C45 X VGND 0.0472f
C46 VPB a_78_159# 0.0517f
C47 X VPB 0.0107f
C48 VPWR B2 0.0104f
C49 VPWR B1 0.0227f
C50 A2 a_292_257# 4.41e-20
C51 a_215_7# a_78_159# 0.0907f
C52 X a_215_7# 0.00228f
C53 VGND VNB 0.403f
C54 VPWR VNB 0.359f
C55 X VNB 0.0884f
C56 A1 VNB 0.132f
C57 A2 VNB 0.0971f
C58 B2 VNB 0.0913f
C59 B1 VNB 0.11f
C60 VPB VNB 0.693f
C61 a_215_7# VNB 0.0357f
C62 a_78_159# VNB 0.154f
.ends

.subckt sky130_fd_sc_hd__o32a_1 VPWR VGND VPB VNB X A1 A2 A3 B2 B1 a_323_257# a_227_7#
+ a_227_257# a_77_159# a_539_257#
X0 a_227_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_227_7# B1 a_77_159# VNB sky130_fd_pr__nfet_01v8 ad=0.189 pd=1.88 as=0.133 ps=1.06 w=0.65 l=0.15
X2 a_539_257# B2 a_77_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X3 VGND A2 a_227_7# VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.107 ps=0.98 w=0.65 l=0.15
X4 a_77_159# B2 a_227_7# VNB sky130_fd_pr__nfet_01v8 ad=0.133 pd=1.06 as=0.127 ps=1.04 w=0.65 l=0.15
X5 VGND a_77_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_227_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X7 a_323_257# A2 a_227_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X8 a_227_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.127 ps=1.04 w=0.65 l=0.15
X9 VPWR B1 a_539_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X10 VPWR a_77_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X11 a_77_159# A3 a_323_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
C0 a_227_7# VGND 0.326f
C1 a_77_159# A1 0.124f
C2 VPB A1 0.029f
C3 a_539_257# a_77_159# 0.0229f
C4 A3 A2 0.106f
C5 a_227_7# A2 0.0413f
C6 VGND A1 0.0197f
C7 a_227_7# a_227_257# 0.00166f
C8 a_539_257# VGND 0.00177f
C9 a_227_7# B1 0.0341f
C10 A1 A2 0.0751f
C11 a_539_257# A2 6.51e-19
C12 a_227_257# A1 3.62e-20
C13 X VPWR 0.102f
C14 a_227_7# A3 0.0376f
C15 B2 X 7.64e-20
C16 a_323_257# VPWR 0.00357f
C17 a_227_7# A1 0.0151f
C18 X a_77_159# 0.0928f
C19 X VPB 0.0157f
C20 B2 VPWR 0.0122f
C21 X VGND 0.103f
C22 a_323_257# a_77_159# 0.0143f
C23 a_77_159# VPWR 0.36f
C24 VPWR VPB 0.0832f
C25 X A2 2.33e-19
C26 a_323_257# VGND 0.00153f
C27 B2 a_77_159# 0.116f
C28 B2 VPB 0.0338f
C29 X a_227_257# 2.01e-21
C30 VPWR VGND 0.0721f
C31 a_323_257# A2 0.0116f
C32 B2 VGND 0.0105f
C33 a_77_159# VPB 0.0477f
C34 VPWR A2 0.0135f
C35 a_227_257# VPWR 0.00277f
C36 X A3 1.25e-19
C37 a_227_7# X 0.0071f
C38 B2 A2 4.92e-19
C39 B1 VPWR 0.0467f
C40 a_77_159# VGND 0.0387f
C41 VPB VGND 0.00632f
C42 B2 B1 0.044f
C43 a_323_257# A3 0.00159f
C44 a_77_159# A2 0.113f
C45 VPB A2 0.0335f
C46 a_227_7# a_323_257# 0.00186f
C47 X A1 0.00148f
C48 A3 VPWR 0.00881f
C49 a_227_257# a_77_159# 0.0187f
C50 a_227_7# VPWR 0.00742f
C51 B1 a_77_159# 0.0468f
C52 B1 VPB 0.0411f
C53 VGND A2 0.0164f
C54 B2 A3 0.102f
C55 a_227_7# B2 0.0275f
C56 a_227_257# VGND 0.00113f
C57 B1 VGND 0.0107f
C58 VPWR A1 0.0187f
C59 a_77_159# A3 0.0306f
C60 A3 VPB 0.033f
C61 a_539_257# VPWR 0.00916f
C62 a_227_7# a_77_159# 0.0851f
C63 a_227_7# VPB 0.00182f
C64 a_227_257# A2 0.003f
C65 a_539_257# B2 0.00242f
C66 A3 VGND 0.0131f
C67 VGND VNB 0.438f
C68 VPWR VNB 0.404f
C69 X VNB 0.101f
C70 B1 VNB 0.15f
C71 B2 VNB 0.0977f
C72 A3 VNB 0.0965f
C73 A2 VNB 0.0962f
C74 A1 VNB 0.0946f
C75 VPB VNB 0.782f
C76 a_227_7# VNB 0.0309f
C77 a_77_159# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND VPB VNB B C A X a_111_257# a_29_13# a_183_257#
X0 VGND A a_29_13# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_29_13# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X2 a_111_257# C a_29_13# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3 X a_29_13# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X4 a_183_257# B a_111_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 a_29_13# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VPWR A a_183_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VGND C a_29_13# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
C0 VGND VPWR 0.0459f
C1 a_111_257# a_29_13# 0.005f
C2 VGND a_29_13# 0.217f
C3 VPWR B 0.147f
C4 VGND C 0.0161f
C5 X VPWR 0.0885f
C6 B a_29_13# 0.121f
C7 X a_29_13# 0.0991f
C8 C B 0.0802f
C9 VGND a_111_257# 3.96e-19
C10 A VPB 0.0377f
C11 VGND B 0.0152f
C12 A a_183_257# 0.00239f
C13 X VGND 0.036f
C14 X B 6.52e-19
C15 A VPWR 0.00936f
C16 VPB VPWR 0.0649f
C17 A a_29_13# 0.242f
C18 a_183_257# VPWR 8.13e-19
C19 A C 0.0343f
C20 VPB a_29_13# 0.0491f
C21 C VPB 0.0396f
C22 a_183_257# a_29_13# 0.00868f
C23 A a_111_257# 0.00223f
C24 VGND A 0.0187f
C25 VGND VPB 0.00724f
C26 VPWR a_29_13# 0.0833f
C27 VGND a_183_257# 5.75e-19
C28 A B 0.0787f
C29 C VPWR 0.00457f
C30 X A 0.00127f
C31 VPB B 0.0962f
C32 X VPB 0.0109f
C33 C a_29_13# 0.0857f
C34 a_111_257# VPWR 5.94e-19
C35 VGND VNB 0.306f
C36 X VNB 0.0882f
C37 A VNB 0.117f
C38 C VNB 0.16f
C39 B VNB 0.117f
C40 VPWR VNB 0.253f
C41 VPB VNB 0.516f
C42 a_29_13# VNB 0.18f
.ends

.subckt sky130_fd_sc_hd__o221a_1 VGND VPWR VPB VNB B1 B2 A2 A1 X C1 a_149_7# a_245_257#
+ a_240_7# a_51_257# a_512_257#
X0 a_245_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1 VPWR C1 a_51_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X2 a_512_257# A2 a_51_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.83 w=1 l=0.15
X3 a_149_7# B2 a_240_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_240_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X5 VGND A1 a_240_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 X a_51_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 a_51_257# B2 a_245_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.83 as=0.105 ps=1.21 w=1 l=0.15
X8 a_240_7# B1 a_149_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X9 a_149_7# C1 a_51_257# VNB sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.201 ps=1.92 w=0.65 l=0.15
X10 VPWR A1 a_512_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X11 X a_51_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
C0 VPB X 0.0262f
C1 B1 C1 0.052f
C2 a_240_7# VGND 0.164f
C3 a_149_7# C1 0.00154f
C4 a_245_257# VGND 0.001f
C5 a_51_257# B1 0.0669f
C6 a_149_7# a_51_257# 0.0249f
C7 VPWR VGND 0.0799f
C8 B2 VGND 0.0107f
C9 A1 a_240_7# 0.023f
C10 a_51_257# X 0.101f
C11 A1 VPWR 0.0215f
C12 A2 X 3.43e-19
C13 a_149_7# B1 0.017f
C14 a_512_257# a_51_257# 0.0116f
C15 VPB VGND 0.00816f
C16 a_245_257# a_240_7# 7.75e-19
C17 VPWR a_240_7# 0.00289f
C18 a_245_257# VPWR 0.00619f
C19 B1 X 8.13e-20
C20 B2 a_240_7# 0.0408f
C21 A1 VPB 0.0255f
C22 a_245_257# B2 7.41e-19
C23 VGND C1 0.0141f
C24 B2 VPWR 0.0135f
C25 VPB a_240_7# 0.0014f
C26 a_51_257# VGND 0.0874f
C27 A2 VGND 0.0159f
C28 a_512_257# X 1.12e-19
C29 VPB VPWR 0.0879f
C30 B2 VPB 0.0366f
C31 A1 a_51_257# 0.125f
C32 B1 VGND 0.00794f
C33 A1 A2 0.0801f
C34 a_149_7# VGND 0.123f
C35 a_240_7# C1 6.33e-20
C36 a_51_257# a_240_7# 0.0314f
C37 a_245_257# a_51_257# 0.0122f
C38 VPWR C1 0.0201f
C39 A2 a_240_7# 0.0566f
C40 a_51_257# VPWR 0.414f
C41 VGND X 0.144f
C42 A2 VPWR 0.0151f
C43 a_512_257# VGND 7.75e-19
C44 B2 a_51_257# 0.0773f
C45 B1 a_240_7# 0.0119f
C46 B2 A2 0.0746f
C47 a_149_7# a_240_7# 0.0687f
C48 VPB C1 0.0515f
C49 A1 X 9.4e-19
C50 B1 VPWR 0.0115f
C51 a_51_257# VPB 0.0632f
C52 a_149_7# VPWR 0.00235f
C53 A2 VPB 0.0386f
C54 B2 B1 0.0797f
C55 a_149_7# B2 0.00653f
C56 VPWR X 0.143f
C57 VPB B1 0.0251f
C58 a_512_257# VPWR 0.00729f
C59 a_149_7# VPB 1.39e-19
C60 a_51_257# C1 0.102f
C61 B2 X 1.41e-19
C62 A1 VGND 0.0277f
C63 A2 a_51_257# 0.0889f
C64 VGND VNB 0.494f
C65 X VNB 0.107f
C66 VPWR VNB 0.409f
C67 A1 VNB 0.0908f
C68 A2 VNB 0.107f
C69 B2 VNB 0.103f
C70 B1 VNB 0.0897f
C71 C1 VNB 0.164f
C72 VPB VNB 0.871f
C73 a_240_7# VNB 0.0138f
C74 a_149_7# VNB 0.00821f
C75 a_51_257# VNB 0.207f
.ends

.subckt sky130_fd_sc_hd__and3_2 VPWR VGND VPB VNB X C B A a_184_13# a_29_271# a_112_13#
X0 VGND C a_184_13# VNB sky130_fd_pr__nfet_01v8 ad=0.13 pd=1.11 as=0.0536 ps=0.675 w=0.42 l=0.15
X1 VPWR a_29_271# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_29_271# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 X a_29_271# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.151 ps=1.35 w=1 l=0.15
X4 VPWR A a_29_271# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X5 a_184_13# B a_112_13# VNB sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 VPWR C a_29_271# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.35 as=0.0744 ps=0.815 w=0.42 l=0.15
X7 X a_29_271# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.13 ps=1.11 w=0.65 l=0.15
X8 a_112_13# A a_29_271# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND a_29_271# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 a_29_271# VPWR 0.178f
C1 VGND B 0.00756f
C2 X VPWR 0.193f
C3 A B 0.0835f
C4 a_184_13# a_29_271# 0.0026f
C5 VPB VPWR 0.0929f
C6 C VPWR 0.00883f
C7 X a_29_271# 0.125f
C8 C a_184_13# 0.00415f
C9 A VGND 0.0127f
C10 a_29_271# VPB 0.0835f
C11 X VPB 0.00641f
C12 a_112_13# VGND 5.13e-19
C13 C a_29_271# 0.189f
C14 C X 0.0158f
C15 B VPWR 0.13f
C16 C VPB 0.0352f
C17 a_29_271# B 0.0596f
C18 X B 8.26e-19
C19 VGND VPWR 0.0591f
C20 A VPWR 0.0156f
C21 a_184_13# VGND 0.00302f
C22 B VPB 0.0923f
C23 a_112_13# VPWR 1.15e-19
C24 C B 0.0649f
C25 a_29_271# VGND 0.143f
C26 X VGND 0.14f
C27 A a_29_271# 0.134f
C28 a_112_13# a_29_271# 0.0049f
C29 VGND VPB 0.00661f
C30 A VPB 0.0443f
C31 C VGND 0.0714f
C32 a_184_13# VPWR 4.26e-19
C33 VGND VNB 0.369f
C34 X VNB 0.04f
C35 C VNB 0.116f
C36 A VNB 0.17f
C37 VPWR VNB 0.336f
C38 B VNB 0.103f
C39 VPB VNB 0.605f
C40 a_29_271# VNB 0.271f
.ends

.subckt sky130_fd_sc_hd__o2111a_1 VPWR VGND VPB VNB X D1 C1 B1 A2 A1 a_306_7# a_79_n19#
+ a_512_7# a_409_7# a_676_257#
X0 VPWR A1 a_676_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A2 a_512_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.198 ps=1.26 w=0.65 l=0.15
X2 a_512_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VPWR a_79_n19# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.382 pd=1.76 as=0.26 ps=2.52 w=1 l=0.15
X4 a_79_n19# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=1.43 as=0.382 ps=1.76 w=1 l=0.15
X5 a_512_7# B1 a_409_7# VNB sky130_fd_pr__nfet_01v8 ad=0.198 pd=1.26 as=0.119 ps=1.01 w=0.65 l=0.15
X6 a_676_257# A2 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.213 ps=1.42 w=1 l=0.15
X7 a_306_7# D1 a_79_n19# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.198 ps=1.91 w=0.65 l=0.15
X8 VGND a_79_n19# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 a_409_7# C1 a_306_7# VNB sky130_fd_pr__nfet_01v8 ad=0.119 pd=1.01 as=0.119 ps=1.01 w=0.65 l=0.15
X10 VPWR C1 a_79_n19# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.218 ps=1.43 w=1 l=0.15
X11 a_79_n19# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.305 ps=1.61 w=1 l=0.15
C0 a_512_7# VPWR 0.00613f
C1 VPB a_512_7# 9.45e-19
C2 D1 VPWR 0.0233f
C3 a_409_7# VGND 0.00662f
C4 a_306_7# VPWR 8.85e-19
C5 a_79_n19# VGND 0.142f
C6 B1 a_512_7# 0.0468f
C7 VPB D1 0.0365f
C8 A1 VGND 0.0184f
C9 X VPWR 0.0949f
C10 C1 VGND 0.0342f
C11 D1 a_512_7# 1.56e-19
C12 a_79_n19# A2 0.0969f
C13 a_306_7# a_512_7# 5.86e-19
C14 a_676_257# VPWR 0.00372f
C15 VPB X 0.0108f
C16 A2 A1 0.121f
C17 a_306_7# D1 0.0092f
C18 a_79_n19# a_409_7# 0.00296f
C19 C1 A2 2.05e-19
C20 a_79_n19# A1 2.4e-19
C21 a_676_257# a_512_7# 7.22e-19
C22 D1 X 3.34e-19
C23 C1 a_409_7# 0.00808f
C24 a_79_n19# C1 0.0401f
C25 VGND VPWR 0.0865f
C26 VPB VGND 0.00797f
C27 B1 VGND 0.0325f
C28 A2 VPWR 0.0848f
C29 a_512_7# VGND 0.17f
C30 A2 VPB 0.0353f
C31 D1 VGND 0.0387f
C32 A2 B1 0.0534f
C33 a_306_7# VGND 0.00515f
C34 a_409_7# VPWR 0.0011f
C35 a_79_n19# VPWR 0.44f
C36 a_79_n19# VPB 0.0534f
C37 A1 VPWR 0.055f
C38 A2 a_512_7# 0.0516f
C39 B1 a_409_7# 0.00322f
C40 a_79_n19# B1 0.0351f
C41 VPB A1 0.04f
C42 VGND X 0.0654f
C43 A2 D1 1.08e-19
C44 C1 VPWR 0.0217f
C45 B1 A1 6.19e-19
C46 a_676_257# VGND 4.92e-19
C47 a_409_7# a_512_7# 0.00102f
C48 a_79_n19# a_512_7# 0.0103f
C49 C1 VPB 0.0347f
C50 C1 B1 0.104f
C51 A1 a_512_7# 0.0432f
C52 a_79_n19# D1 0.155f
C53 a_306_7# a_79_n19# 0.00291f
C54 C1 a_512_7# 3.26e-19
C55 a_676_257# A2 0.0099f
C56 C1 D1 0.118f
C57 a_306_7# C1 0.00228f
C58 a_79_n19# X 0.091f
C59 a_676_257# a_79_n19# 2.93e-19
C60 a_676_257# A1 2.93e-19
C61 VPB VPWR 0.0881f
C62 B1 VPWR 0.0218f
C63 A2 VGND 0.0191f
C64 B1 VPB 0.0377f
C65 VGND VNB 0.491f
C66 VPWR VNB 0.414f
C67 X VNB 0.0907f
C68 A1 VNB 0.154f
C69 A2 VNB 0.104f
C70 B1 VNB 0.114f
C71 C1 VNB 0.0988f
C72 D1 VNB 0.112f
C73 VPB VNB 0.871f
C74 a_512_7# VNB 0.0326f
C75 a_79_n19# VNB 0.158f
.ends

.subckt sky130_fd_sc_hd__a221oi_2 VGND VPWR VPB VNB A2 A1 B1 B2 Y C1 a_27_257# a_301_257#
+ a_383_7# a_735_7#
X0 a_27_257# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_301_257# B2 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.135 ps=1.27 w=1 l=0.15
X2 a_735_7# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X3 a_27_257# B1 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.176 ps=1.84 w=0.65 l=0.15
X5 a_301_257# B1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_301_257# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.135 ps=1.27 w=1 l=0.15
X7 a_27_257# B2 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X8 VPWR A1 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_301_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y C1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X11 Y A1 a_735_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 a_735_7# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 VGND A2 a_735_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 VPWR A2 a_301_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.175 ps=1.35 w=1 l=0.15
X15 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_383_7# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.257 ps=1.44 w=0.65 l=0.15
X17 Y B1 a_383_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 a_383_7# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 VGND B2 a_383_7# VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 B2 VPWR 0.0224f
C1 B2 Y 0.118f
C2 VGND A1 0.0175f
C3 A2 VPB 0.0709f
C4 a_301_257# A1 0.0293f
C5 VGND C1 0.0632f
C6 B1 VGND 0.0184f
C7 a_735_7# VPB 2.96e-19
C8 B1 a_301_257# 0.0185f
C9 a_27_257# VPB 0.0204f
C10 a_383_7# a_735_7# 2.58e-19
C11 B2 VGND 0.0325f
C12 VPWR VPB 0.108f
C13 Y VPB 0.00812f
C14 B2 a_301_257# 0.0418f
C15 a_735_7# A2 0.0309f
C16 a_27_257# A2 1.13e-19
C17 a_383_7# VPWR 0.00192f
C18 a_383_7# Y 0.0983f
C19 B2 C1 0.0205f
C20 B2 B1 0.213f
C21 VPWR A2 0.0455f
C22 A2 Y 0.0455f
C23 VGND VPB 0.00991f
C24 a_301_257# VPB 0.0181f
C25 VPWR a_735_7# 0.00213f
C26 a_735_7# Y 0.0886f
C27 A1 VPB 0.051f
C28 a_27_257# VPWR 0.164f
C29 a_27_257# Y 0.128f
C30 a_383_7# VGND 0.165f
C31 C1 VPB 0.078f
C32 B1 VPB 0.051f
C33 VPWR Y 0.0129f
C34 VGND A2 0.0568f
C35 a_301_257# A2 0.186f
C36 VGND a_735_7# 0.206f
C37 B1 a_383_7# 0.0137f
C38 B2 VPB 0.0679f
C39 A2 A1 0.207f
C40 a_27_257# VGND 0.00854f
C41 a_27_257# a_301_257# 0.191f
C42 a_735_7# A1 0.0216f
C43 C1 a_735_7# 1.39e-20
C44 VGND VPWR 0.106f
C45 VGND Y 0.258f
C46 B1 a_735_7# 1.04e-19
C47 a_27_257# A1 1.01e-19
C48 B2 a_383_7# 0.00622f
C49 a_301_257# VPWR 0.48f
C50 a_301_257# Y 0.00522f
C51 a_27_257# C1 0.0611f
C52 B1 a_27_257# 0.0195f
C53 B2 A2 0.0926f
C54 VPWR A1 0.0298f
C55 Y A1 0.0483f
C56 VPWR C1 0.0192f
C57 C1 Y 0.106f
C58 B2 a_735_7# 1.28e-19
C59 B1 VPWR 0.0152f
C60 B1 Y 0.0643f
C61 B2 a_27_257# 0.153f
C62 a_301_257# VGND 0.00922f
C63 VGND VNB 0.682f
C64 VPWR VNB 0.52f
C65 Y VNB 0.0379f
C66 A1 VNB 0.166f
C67 A2 VNB 0.23f
C68 B1 VNB 0.166f
C69 B2 VNB 0.195f
C70 C1 VNB 0.255f
C71 VPB VNB 1.14f
C72 a_735_7# VNB 0.00532f
C73 a_383_7# VNB 0.00406f
C74 a_301_257# VNB 0.0376f
C75 a_27_257# VNB 0.0292f
.ends

.subckt sky130_fd_sc_hd__nand2_1 VGND VPWR VPB VNB A Y B a_113_7#
X0 Y A a_113_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_113_7# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
C0 VPWR VPB 0.0509f
C1 VPWR Y 0.211f
C2 Y VPB 0.00618f
C3 a_113_7# VPWR 1.78e-19
C4 a_113_7# Y 0.00937f
C5 VGND A 0.00949f
C6 VGND B 0.0544f
C7 A B 0.051f
C8 VGND VPWR 0.0322f
C9 VPWR A 0.0444f
C10 VPWR B 0.0478f
C11 VGND VPB 0.0044f
C12 VGND Y 0.139f
C13 A VPB 0.0379f
C14 B VPB 0.0391f
C15 A Y 0.0855f
C16 Y B 0.0481f
C17 a_113_7# VGND 0.0019f
C18 VGND VNB 0.232f
C19 Y VNB 0.0557f
C20 VPWR VNB 0.245f
C21 A VNB 0.143f
C22 B VNB 0.146f
C23 VPB VNB 0.339f
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR VPB VNB X C B A a_27_7# a_109_7# a_181_7#
X0 a_27_7# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_181_7# B a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X3 VPWR A a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X4 VPWR C a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X5 VGND C a_181_7# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_109_7# A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X7 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
C0 X VPB 0.0121f
C1 C B 0.0746f
C2 A VPB 0.0426f
C3 a_181_7# VPWR 3.97e-19
C4 A a_109_7# 6.45e-19
C5 C VPWR 0.00464f
C6 a_27_7# B 0.0625f
C7 a_181_7# C 0.00151f
C8 VGND B 0.00714f
C9 a_27_7# VPWR 0.145f
C10 a_27_7# a_181_7# 0.00401f
C11 VGND VPWR 0.0475f
C12 a_27_7# C 0.186f
C13 a_181_7# VGND 0.00261f
C14 B VPB 0.0836f
C15 C VGND 0.0703f
C16 VPWR VPB 0.0795f
C17 X B 0.00111f
C18 a_27_7# VGND 0.134f
C19 a_109_7# VPWR 3.29e-19
C20 A B 0.0869f
C21 C VPB 0.0347f
C22 X VPWR 0.0766f
C23 A VPWR 0.0185f
C24 a_27_7# VPB 0.0501f
C25 C X 0.0149f
C26 a_27_7# a_109_7# 0.00517f
C27 VGND VPB 0.00604f
C28 a_27_7# X 0.087f
C29 a_109_7# VGND 0.00123f
C30 A a_27_7# 0.157f
C31 VGND X 0.0708f
C32 A VGND 0.0154f
C33 B VPWR 0.128f
C34 VGND VNB 0.3f
C35 X VNB 0.0923f
C36 C VNB 0.12f
C37 A VNB 0.174f
C38 VPWR VNB 0.274f
C39 B VNB 0.102f
C40 VPB VNB 0.516f
C41 a_27_7# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__o22ai_1 VGND VPWR VPB VNB A1 A2 B1 B2 Y a_109_257# a_307_257#
+ a_27_7#
X0 Y B2 a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.233 pd=1.47 as=0.112 ps=1.23 w=1 l=0.15
X1 a_109_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.112 pd=1.23 as=0.26 ps=2.52 w=1 l=0.15
X2 VGND A2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.115 ps=1 w=0.65 l=0.15
X3 a_27_7# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_27_7# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0.115 pd=1 as=0.0926 ps=0.935 w=0.65 l=0.15
X5 VPWR A1 a_307_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.105 ps=1.21 w=1 l=0.15
X6 Y B1 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0926 pd=0.935 as=0.169 ps=1.82 w=0.65 l=0.15
X7 a_307_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.233 ps=1.47 w=1 l=0.15
C0 a_27_7# VGND 0.244f
C1 VPB a_27_7# 9.43e-19
C2 B1 VGND 0.0142f
C3 a_109_257# VGND 9.92e-19
C4 A2 a_27_7# 0.046f
C5 VPB B1 0.0427f
C6 a_109_257# A2 3.1e-19
C7 Y VGND 0.00968f
C8 B1 a_27_7# 0.0334f
C9 B2 VGND 0.0105f
C10 VPB Y 0.00499f
C11 A1 VPWR 0.0569f
C12 A2 Y 0.063f
C13 B2 VPB 0.0302f
C14 B2 A2 0.091f
C15 a_27_7# Y 0.0527f
C16 VPWR a_307_257# 0.00219f
C17 B2 a_27_7# 0.0266f
C18 B1 Y 0.132f
C19 a_109_257# Y 0.0135f
C20 B2 B1 0.0576f
C21 B2 a_109_257# 5.79e-19
C22 B2 Y 0.12f
C23 A1 VGND 0.0147f
C24 A1 VPB 0.0315f
C25 A1 A2 0.089f
C26 a_307_257# VGND 2.4e-19
C27 VPWR VGND 0.0459f
C28 A1 a_27_7# 0.0495f
C29 A2 a_307_257# 0.0107f
C30 VPB VPWR 0.0612f
C31 A2 VPWR 0.119f
C32 a_307_257# a_27_7# 2.6e-19
C33 VPWR a_27_7# 0.00678f
C34 A1 Y 5.15e-19
C35 B1 VPWR 0.0451f
C36 a_109_257# VPWR 0.00394f
C37 B2 A1 4.27e-19
C38 a_307_257# Y 3.52e-19
C39 VPWR Y 0.102f
C40 B2 VPWR 0.0114f
C41 VPB VGND 0.0047f
C42 A2 VGND 0.0158f
C43 A2 VPB 0.0309f
C44 VGND VNB 0.298f
C45 Y VNB 0.0144f
C46 VPWR VNB 0.298f
C47 A1 VNB 0.131f
C48 A2 VNB 0.0973f
C49 B2 VNB 0.0939f
C50 B1 VNB 0.184f
C51 VPB VNB 0.516f
C52 a_27_7# VNB 0.0465f
.ends

.subckt sky130_fd_sc_hd__or3_4 VPWR VGND VPB VNB B C A X a_109_257# a_27_7# a_193_257#
X0 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_109_257# C a_27_7# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_7# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.4 ps=1.8 w=1 l=0.15
X4 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.205 pd=1.93 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_27_7# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VGND A a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 VPWR A a_193_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=1.8 as=0.135 ps=1.27 w=1 l=0.15
X8 a_193_257# B a_109_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR a_27_7# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND C a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.26 ps=1.45 w=0.65 l=0.15
X12 VGND a_27_7# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_27_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
C0 B VGND 0.0163f
C1 VPWR VPB 0.0867f
C2 a_27_7# X 0.397f
C3 A a_27_7# 0.159f
C4 VPWR C 0.00921f
C5 a_109_257# VPWR 0.00187f
C6 A X 5.59e-19
C7 VGND VPB 0.00698f
C8 B a_27_7# 0.19f
C9 a_193_257# VPWR 8.05e-19
C10 VGND C 0.0149f
C11 a_109_257# VGND 7.33e-19
C12 B A 0.0783f
C13 VPWR VGND 0.0864f
C14 a_27_7# VPB 0.158f
C15 a_193_257# VGND 2.86e-19
C16 X VPB 0.0146f
C17 a_27_7# C 0.0996f
C18 a_109_257# a_27_7# 0.0105f
C19 A VPB 0.0324f
C20 a_27_7# VPWR 0.363f
C21 a_27_7# a_193_257# 0.015f
C22 B VPB 0.0302f
C23 VPWR X 0.365f
C24 A VPWR 0.0196f
C25 B C 0.0864f
C26 A a_193_257# 3.02e-21
C27 B a_109_257# 0.00939f
C28 a_27_7# VGND 0.352f
C29 B VPWR 0.0132f
C30 VGND X 0.265f
C31 B a_193_257# 0.00132f
C32 A VGND 0.0164f
C33 VPB C 0.0369f
C34 VGND VNB 0.493f
C35 X VNB 0.0611f
C36 VPWR VNB 0.418f
C37 A VNB 0.0987f
C38 B VNB 0.0938f
C39 C VNB 0.141f
C40 VPB VNB 0.871f
C41 a_27_7# VNB 0.499f
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VGND VPWR VPB VNB B1 B2 A2_N A1_N X a_226_257# a_76_159#
+ a_556_7# a_226_7# a_489_373#
X0 VPWR a_76_159# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.43 as=0.26 ps=2.52 w=1 l=0.15
X1 a_226_7# A2_N a_226_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X2 a_76_159# a_226_7# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.139 ps=1.08 w=0.42 l=0.15
X3 a_556_7# B2 a_76_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_226_7# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.12 ps=1.09 w=0.42 l=0.15
X5 VGND B1 a_556_7# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_226_257# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.167 ps=1.43 w=0.42 l=0.15
X7 VGND A2_N a_226_7# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_489_373# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 VPWR B2 a_489_373# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 VGND a_76_159# X VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.09 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_489_373# a_226_7# a_76_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
C0 a_556_7# VPWR 7.24e-19
C1 a_226_257# VPWR 8.54e-19
C2 a_226_7# A2_N 0.141f
C3 a_76_159# A1_N 0.119f
C4 B2 a_489_373# 0.0541f
C5 B1 VGND 0.0471f
C6 X A2_N 2.55e-19
C7 a_76_159# B2 0.0626f
C8 a_226_7# VGND 0.149f
C9 VPWR A1_N 0.00672f
C10 a_76_159# a_489_373# 0.0473f
C11 VPB A1_N 0.0339f
C12 X VGND 0.0627f
C13 B2 VPWR 0.0161f
C14 VPB B2 0.0645f
C15 a_489_373# VPWR 0.143f
C16 X a_226_7# 0.0108f
C17 VPB a_489_373# 0.015f
C18 a_556_7# VGND 0.00639f
C19 a_226_257# VGND 5.63e-19
C20 a_76_159# VPWR 0.2f
C21 VPB a_76_159# 0.0817f
C22 A2_N A1_N 0.11f
C23 a_226_7# a_226_257# 0.00128f
C24 VPB VPWR 0.0951f
C25 VGND A1_N 0.0261f
C26 B2 VGND 0.0335f
C27 B1 B2 0.182f
C28 a_76_159# A2_N 0.0125f
C29 a_226_7# A1_N 0.0209f
C30 a_489_373# VGND 0.0058f
C31 X A1_N 0.00211f
C32 B1 a_489_373# 0.0382f
C33 B2 a_226_7# 0.0975f
C34 a_76_159# VGND 0.108f
C35 A2_N VPWR 0.00449f
C36 a_76_159# B1 0.00185f
C37 VPB A2_N 0.0327f
C38 a_226_7# a_489_373# 0.00579f
C39 a_76_159# a_226_7# 0.188f
C40 VGND VPWR 0.0743f
C41 a_226_257# A1_N 0.00184f
C42 B1 VPWR 0.0188f
C43 VPB VGND 0.0128f
C44 a_76_159# X 0.0995f
C45 VPB B1 0.0803f
C46 B2 a_556_7# 0.00291f
C47 a_226_7# VPWR 0.0187f
C48 VPB a_226_7# 0.111f
C49 X VPWR 0.0589f
C50 VPB X 0.0113f
C51 a_76_159# a_556_7# 0.0017f
C52 a_76_159# a_226_257# 0.00354f
C53 A2_N VGND 0.0174f
C54 VGND VNB 0.462f
C55 A2_N VNB 0.103f
C56 A1_N VNB 0.111f
C57 VPWR VNB 0.369f
C58 X VNB 0.0975f
C59 B1 VNB 0.206f
C60 B2 VNB 0.106f
C61 VPB VNB 0.782f
C62 a_489_373# VNB 0.0254f
C63 a_226_7# VNB 0.162f
C64 a_76_159# VNB 0.141f
.ends

.subckt sky130_fd_sc_hd__nor2_2 VGND VPWR VPB VNB B Y A a_27_257#
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 a_27_257# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 Y B a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_257# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X7 VPWR A a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
C0 VGND A 0.0597f
C1 VGND a_27_257# 0.00726f
C2 VPB A 0.0563f
C3 Y A 0.0523f
C4 a_27_257# VPB 0.0203f
C5 Y a_27_257# 0.152f
C6 VGND VPB 0.00613f
C7 Y VGND 0.289f
C8 B A 0.0712f
C9 a_27_257# B 0.0451f
C10 Y VPB 0.00961f
C11 VPWR A 0.0418f
C12 a_27_257# VPWR 0.321f
C13 VGND B 0.0294f
C14 VGND VPWR 0.0467f
C15 B VPB 0.0566f
C16 Y B 0.179f
C17 VPWR VPB 0.05f
C18 Y VPWR 0.0127f
C19 a_27_257# A 0.0889f
C20 B VPWR 0.0174f
C21 VGND VNB 0.343f
C22 Y VNB 0.0641f
C23 VPWR VNB 0.249f
C24 B VNB 0.198f
C25 A VNB 0.207f
C26 VPB VNB 0.516f
C27 a_27_257# VNB 0.0647f
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND VPB VNB X A B a_145_35# a_59_35#
X0 a_145_35# A a_59_35# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1 VPWR B a_59_35# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 X a_59_35# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X3 VGND B a_145_35# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 a_59_35# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X5 X a_59_35# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
C0 B VPB 0.0629f
C1 VPWR A 0.0362f
C2 a_59_35# VPWR 0.15f
C3 X A 1.68e-19
C4 a_59_35# X 0.109f
C5 VGND a_145_35# 0.00468f
C6 a_59_35# A 0.0809f
C7 B VPWR 0.0117f
C8 B X 0.00276f
C9 VGND VPB 0.008f
C10 B A 0.0971f
C11 B a_59_35# 0.143f
C12 VGND VPWR 0.0461f
C13 VGND X 0.0993f
C14 VPWR a_145_35# 6.31e-19
C15 X a_145_35# 5.76e-19
C16 VGND A 0.0147f
C17 a_59_35# VGND 0.116f
C18 a_59_35# a_145_35# 0.00658f
C19 VPWR VPB 0.0729f
C20 B VGND 0.0115f
C21 X VPB 0.0127f
C22 VPB A 0.0806f
C23 a_59_35# VPB 0.0563f
C24 X VPWR 0.111f
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_35# VNB 0.177f
.ends

.subckt sky130_fd_sc_hd__or4b_4 VGND VPWR VPB VNB X D_N C B A a_403_257# a_215_257#
+ a_487_257# a_109_53# a_297_257#
X0 a_297_257# a_109_53# a_215_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X1 X a_215_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X2 X a_215_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 VGND a_215_257# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_215_257# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VPWR a_215_257# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X7 a_215_257# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.165 ps=1.82 w=0.65 l=0.15
X8 X a_215_257# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X9 VPWR A a_487_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X10 VGND a_215_257# X VNB sky130_fd_pr__nfet_01v8 ad=0.179 pd=1.85 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 a_487_257# B a_403_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 VGND C a_215_257# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X13 a_215_257# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_403_257# C a_297_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X15 VGND A a_215_257# VNB sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X17 VPWR a_215_257# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
C0 B a_403_257# 0.00615f
C1 VGND A 0.0184f
C2 VGND B 0.0177f
C3 VPWR C 0.0452f
C4 X a_487_257# 5.61e-19
C5 a_109_53# C 0.046f
C6 VPWR X 0.358f
C7 a_215_257# D_N 0.00255f
C8 VGND a_487_257# 1e-18
C9 VPWR a_403_257# 0.00597f
C10 a_215_257# a_297_257# 0.0145f
C11 a_109_53# a_403_257# 1.29e-20
C12 VGND VPWR 0.103f
C13 VGND a_109_53# 0.0965f
C14 a_215_257# VPB 0.133f
C15 C a_403_257# 0.011f
C16 VGND C 0.017f
C17 D_N VPB 0.107f
C18 a_215_257# A 0.111f
C19 a_215_257# B 0.0415f
C20 VGND X 0.245f
C21 A D_N 7.84e-20
C22 D_N B 3.04e-19
C23 VGND a_403_257# 0.00131f
C24 a_215_257# a_487_257# 0.00167f
C25 A VPB 0.031f
C26 B VPB 0.0282f
C27 a_215_257# VPWR 0.154f
C28 a_215_257# a_109_53# 0.152f
C29 A B 0.108f
C30 VPWR D_N 0.0486f
C31 a_215_257# C 0.126f
C32 a_109_53# D_N 0.119f
C33 VPWR a_297_257# 0.00828f
C34 a_215_257# X 0.366f
C35 a_109_53# a_297_257# 3.03e-20
C36 D_N C 6.87e-19
C37 VPWR VPB 0.117f
C38 a_109_53# VPB 0.0623f
C39 X D_N 3.65e-19
C40 a_297_257# C 0.0109f
C41 A a_487_257# 7.1e-19
C42 B a_487_257# 0.0126f
C43 a_215_257# a_403_257# 0.00122f
C44 C VPB 0.0292f
C45 VPWR A 0.0526f
C46 VPWR B 0.0819f
C47 VGND a_215_257# 0.294f
C48 a_109_53# A 3.09e-21
C49 a_109_53# B 4.77e-21
C50 X VPB 0.0127f
C51 VGND D_N 0.0426f
C52 B C 0.161f
C53 A X 0.0157f
C54 X B 0.0046f
C55 VGND a_297_257# 0.00213f
C56 VPWR a_487_257# 0.0056f
C57 a_109_53# a_487_257# 8.62e-21
C58 VGND VPB 0.0105f
C59 a_109_53# VPWR 0.0693f
C60 VGND VNB 0.631f
C61 X VNB 0.0581f
C62 VPWR VNB 0.515f
C63 A VNB 0.0911f
C64 B VNB 0.0892f
C65 C VNB 0.0908f
C66 D_N VNB 0.186f
C67 VPB VNB 1.05f
C68 a_215_257# VNB 0.414f
C69 a_109_53# VNB 0.148f
.ends

.subckt sky130_fd_sc_hd__a31oi_2 VPWR VGND VPB VNB B1 Y A1 A2 A3 a_27_257# a_27_7#
+ a_277_7#
X0 VPWR A3 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X2 VPWR A1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X3 a_27_7# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 a_277_7# A2 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_277_7# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X7 a_27_257# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 a_27_257# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X9 a_27_7# A2 a_277_7# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VPWR A2 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 a_27_257# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A1 a_277_7# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X13 a_27_257# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X14 VGND A3 a_27_7# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 Y B1 a_27_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
C0 a_27_7# VGND 0.0907f
C1 a_277_7# Y 0.086f
C2 A3 a_277_7# 7.39e-19
C3 VPB VGND 0.00575f
C4 A1 a_27_7# 0.0129f
C5 A1 VPB 0.0971f
C6 Y VGND 0.168f
C7 B1 a_27_257# 0.045f
C8 VPB a_27_7# 9.31e-19
C9 A3 VGND 0.0355f
C10 B1 VPWR 0.0218f
C11 A1 Y 0.118f
C12 a_27_7# Y 0.0142f
C13 VPWR a_27_257# 0.558f
C14 A3 a_27_7# 0.0773f
C15 VPB Y 0.00779f
C16 a_27_257# A2 0.0837f
C17 A3 VPB 0.0731f
C18 VPWR A2 0.0396f
C19 a_27_257# a_277_7# 1.45e-19
C20 A3 Y 3.4e-19
C21 VPWR a_277_7# 0.00227f
C22 B1 VGND 0.0344f
C23 a_277_7# A2 0.0093f
C24 B1 A1 0.0382f
C25 a_27_257# VGND 0.0107f
C26 VPWR VGND 0.0914f
C27 A1 a_27_257# 0.0972f
C28 B1 VPB 0.0808f
C29 A2 VGND 0.0246f
C30 A1 VPWR 0.0475f
C31 a_27_257# a_27_7# 0.0108f
C32 A1 A2 0.0965f
C33 VPB a_27_257# 0.0116f
C34 VPWR a_27_7# 0.00469f
C35 a_277_7# VGND 0.169f
C36 B1 Y 0.177f
C37 VPB VPWR 0.0885f
C38 a_27_7# A2 0.074f
C39 A1 a_277_7# 0.0176f
C40 VPB A2 0.0568f
C41 a_27_257# Y 0.13f
C42 A3 a_27_257# 0.083f
C43 a_277_7# a_27_7# 0.0683f
C44 VPWR Y 0.0196f
C45 A3 VPWR 0.0415f
C46 A2 Y 7.37e-19
C47 A1 VGND 0.0281f
C48 A3 A2 0.106f
C49 VGND VNB 0.538f
C50 Y VNB 0.06f
C51 VPWR VNB 0.436f
C52 B1 VNB 0.258f
C53 A1 VNB 0.24f
C54 A2 VNB 0.179f
C55 A3 VNB 0.246f
C56 VPB VNB 0.959f
C57 a_277_7# VNB 0.00976f
C58 a_27_7# VNB 0.0193f
C59 a_27_257# VNB 0.0672f
.ends

.subckt sky130_fd_sc_hd__o221ai_1 VGND VPWR VPB VNB A1 A2 Y B2 C1 B1 a_213_83# a_295_257#
+ a_493_257# a_109_7#
X0 a_213_83# B2 a_109_7# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 Y B2 a_295_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.12 ps=1.24 w=1 l=0.15
X2 VPWR A1 a_493_257# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3 VGND A2 a_213_83# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X4 a_213_83# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 a_295_257# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12 pd=1.24 as=0.38 ps=1.76 w=1 l=0.15
X6 a_493_257# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.225 ps=1.45 w=1 l=0.15
X7 a_109_7# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=1.76 as=0.28 ps=2.56 w=1 l=0.15
X9 a_109_7# B1 a_213_83# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.165 ps=1.82 w=0.65 l=0.15
C0 A2 a_213_83# 0.0451f
C1 B2 a_213_83# 0.0489f
C2 VPWR A2 0.115f
C3 VPWR B2 0.00898f
C4 A1 Y 3.82e-19
C5 a_295_257# Y 0.0137f
C6 Y B1 0.0768f
C7 C1 B1 0.0209f
C8 A1 a_213_83# 0.0506f
C9 a_109_7# VPB 4.01e-19
C10 a_295_257# a_213_83# 1.01e-20
C11 C1 Y 0.127f
C12 VPWR A1 0.0503f
C13 VPB VGND 0.0063f
C14 VPWR a_295_257# 0.00875f
C15 a_493_257# VGND 9.1e-20
C16 B1 a_213_83# 0.0383f
C17 VPWR B1 0.0222f
C18 Y a_213_83# 0.0301f
C19 A2 VPB 0.0328f
C20 B2 VPB 0.028f
C21 C1 a_213_83# 1.34e-19
C22 a_493_257# A2 0.0112f
C23 VPWR Y 0.293f
C24 VPWR C1 0.0213f
C25 a_109_7# VGND 0.115f
C26 VPWR a_213_83# 0.004f
C27 a_109_7# B2 0.00286f
C28 A2 VGND 0.0162f
C29 A1 VPB 0.0359f
C30 B2 VGND 0.0119f
C31 B1 VPB 0.0341f
C32 A2 B2 0.0666f
C33 Y VPB 0.0205f
C34 C1 VPB 0.038f
C35 a_493_257# Y 3.47e-19
C36 A1 VGND 0.0151f
C37 a_295_257# VGND 0.00139f
C38 a_109_7# B1 0.00614f
C39 VPB a_213_83# 0.00108f
C40 VPWR VPB 0.0746f
C41 Y a_109_7# 0.0456f
C42 B1 VGND 0.0106f
C43 A1 A2 0.0891f
C44 A1 B2 5.58e-19
C45 C1 a_109_7# 0.00243f
C46 VPWR a_493_257# 8.66e-19
C47 a_295_257# A2 4.69e-20
C48 a_295_257# B2 5.73e-20
C49 Y VGND 0.046f
C50 C1 VGND 0.0128f
C51 A2 B1 4.14e-19
C52 B2 B1 0.0868f
C53 a_109_7# a_213_83# 0.0875f
C54 A2 Y 0.0805f
C55 Y B2 0.0569f
C56 VPWR a_109_7# 0.0018f
C57 VGND a_213_83# 0.167f
C58 VPWR VGND 0.0645f
C59 VGND VNB 0.39f
C60 VPWR VNB 0.362f
C61 Y VNB 0.0858f
C62 A1 VNB 0.14f
C63 A2 VNB 0.0967f
C64 B2 VNB 0.0933f
C65 B1 VNB 0.106f
C66 C1 VNB 0.145f
C67 VPB VNB 0.693f
C68 a_213_83# VNB 0.0371f
C69 a_109_7# VNB 0.0115f
.ends

.subckt sarlogic ctln[0] ctln[1] ctln[2] ctln[3] ctln[4] ctln[5] ctln[6] ctln[7] ctlp[0]
+ ctlp[1] ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6] ctlp[7] cal clk clkc comp en result[0]
+ result[1] result[2] result[3] result[4] result[5] result[6] result[7] rstn sample
+ trim[0] trim[1] trim[2] trim[3] trim[4] trimb[0] trimb[1] trimb[2] trimb[3] trimb[4]
+ valid VPWR VGND
XFILLER_13_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_294_ VPWR VGND VPWR VGND _294_/Y _294_/A sky130_fd_sc_hd__inv_2
X_346_ VPWR VGND VPWR VGND _346_/Q _346_/SET_B _346_/D _297_/B _346_/a_652_n19# _346_/a_1602_7#
+ _346_/a_562_373# _346_/a_1032_373# _346_/a_1296_7# _346_/a_796_7# _346_/a_586_7#
+ _346_/a_1056_7# _346_/a_381_7# _346_/a_193_7# _346_/a_1140_373# _346_/a_27_7# _346_/a_956_373#
+ _346_/a_476_7# _346_/a_1224_7# _346_/a_1182_221# sky130_fd_sc_hd__dfstp_1
X_277_ VPWR VGND VPWR VGND _277_/Y _277_/A sky130_fd_sc_hd__inv_2
XFILLER_5_162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_200_ VGND VPWR VPWR VGND _337_/D _193_/Y _197_/X _338_/Q _337_/Q _194_/X _200_/a_584_7#
+ _200_/a_346_7# _200_/a_256_7# _200_/a_250_257# _200_/a_93_n19# sky130_fd_sc_hd__a32o_1
X_329_ VGND VPWR VPWR VGND _331_/CLK _329_/D _346_/SET_B _329_/Q _329_/a_639_7# _329_/a_805_7#
+ _329_/a_448_7# _329_/a_543_7# _329_/a_1283_n19# _329_/a_1462_7# _329_/a_1270_373#
+ _329_/a_193_7# _329_/a_1217_7# _329_/a_761_249# _329_/a_27_7# _329_/a_1108_7# _329_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_68 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_18_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput20 VGND VPWR VPWR VGND _281_/A ctlp[6] output20/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_16_142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xoutput7 VGND VPWR VPWR VGND _271_/Y ctln[1] output7/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput31 VGND VPWR VPWR VGND _285_/A trim[0] output31/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_22_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_293_ VPWR VGND VPWR VGND _294_/A _340_/Q _313_/Q _293_/a_121_257# _293_/a_39_257#
+ sky130_fd_sc_hd__or2_2
XFILLER_9_138 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_10_126 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_276_ VGND VPWR VPWR VGND _277_/A _328_/Q _319_/Q _276_/a_68_257# _276_/a_150_257#
+ sky130_fd_sc_hd__or2_1
X_345_ VPWR VGND VPWR VGND _345_/Q _346_/SET_B _345_/D _297_/B _345_/a_652_n19# _345_/a_1602_7#
+ _345_/a_562_373# _345_/a_1032_373# _345_/a_1296_7# _345_/a_796_7# _345_/a_586_7#
+ _345_/a_1056_7# _345_/a_381_7# _345_/a_193_7# _345_/a_1140_373# _345_/a_27_7# _345_/a_956_373#
+ _345_/a_476_7# _345_/a_1224_7# _345_/a_1182_221# sky130_fd_sc_hd__dfstp_1
X_328_ VGND VPWR VPWR VGND _297_/B _328_/D _346_/SET_B _328_/Q _328_/a_639_7# _328_/a_805_7#
+ _328_/a_448_7# _328_/a_543_7# _328_/a_1283_n19# _328_/a_1462_7# _328_/a_1270_373#
+ _328_/a_193_7# _328_/a_1217_7# _328_/a_761_249# _328_/a_27_7# _328_/a_1108_7# _328_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_259_ VPWR VGND VPWR VGND _258_/S _339_/Q _312_/Q _261_/A _259_/a_199_7# _259_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
XFILLER_9_67 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_20_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
Xoutput21 VGND VPWR VPWR VGND _283_/A ctlp[7] output21/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_16_154 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput8 VGND VPWR VPWR VGND _273_/Y ctln[2] output8/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput10 VGND VPWR VPWR VGND _277_/Y ctln[4] output10/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput32 VGND VPWR VPWR VGND _288_/A trim[1] output32/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_22_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_292_ VPWR VGND VPWR VGND _292_/Y _292_/A sky130_fd_sc_hd__inv_2
XFILLER_3_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_34 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_109 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_275_ VPWR VGND VPWR VGND _275_/Y _275_/A sky130_fd_sc_hd__inv_2
X_344_ VPWR VGND VPWR VGND _344_/Q _346_/SET_B _344_/D _297_/B _344_/a_652_n19# _344_/a_1602_7#
+ _344_/a_562_373# _344_/a_1032_373# _344_/a_1296_7# _344_/a_796_7# _344_/a_586_7#
+ _344_/a_1056_7# _344_/a_381_7# _344_/a_193_7# _344_/a_1140_373# _344_/a_27_7# _344_/a_956_373#
+ _344_/a_476_7# _344_/a_1224_7# _344_/a_1182_221# sky130_fd_sc_hd__dfstp_1
XFILLER_5_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_59 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_327_ VGND VPWR VPWR VGND _331_/CLK _327_/D _346_/SET_B _327_/Q _327_/a_639_7# _327_/a_805_7#
+ _327_/a_448_7# _327_/a_543_7# _327_/a_1283_n19# _327_/a_1462_7# _327_/a_1270_373#
+ _327_/a_193_7# _327_/a_1217_7# _327_/a_761_249# _327_/a_27_7# _327_/a_1108_7# _327_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_189_ VGND VPWR VPWR VGND _196_/A _190_/A _189_/a_27_7# sky130_fd_sc_hd__clkbuf_2
X_258_ VGND VPWR VPWR VGND _313_/D _306_/X _258_/S _313_/Q _258_/a_505_n19# _258_/a_535_334#
+ _258_/a_76_159# _258_/a_218_334# _258_/a_439_7# _258_/a_218_7# sky130_fd_sc_hd__mux2_1
XFILLER_6_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xoutput22 VGND VPWR VPWR VGND _315_/Q result[0] output22/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput33 VGND VPWR VPWR VGND _290_/A trim[2] output33/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput9 VGND VPWR VPWR VGND _275_/Y ctln[3] output9/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput11 VGND VPWR VPWR VGND _279_/Y ctln[5] output11/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_22_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_291_ VPWR VGND VPWR VGND _292_/A _339_/Q _312_/Q _291_/a_121_257# _291_/a_39_257#
+ sky130_fd_sc_hd__or2_2
XFILLER_12_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_274_ VPWR VGND VPWR VGND _275_/A _327_/Q _318_/Q _274_/a_121_257# _274_/a_39_257#
+ sky130_fd_sc_hd__or2_2
XFILLER_5_154 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_343_ VGND VPWR VPWR VGND _343_/CLK _343_/D repeater43/X _343_/Q _343_/a_639_7# _343_/a_805_7#
+ _343_/a_448_7# _343_/a_543_7# _343_/a_1283_n19# _343_/a_1462_7# _343_/a_1270_373#
+ _343_/a_193_7# _343_/a_1217_7# _343_/a_761_249# _343_/a_27_7# _343_/a_1108_7# _343_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_326_ VGND VPWR VPWR VGND _331_/CLK _326_/D repeater43/X _326_/Q _326_/a_639_7# _326_/a_805_7#
+ _326_/a_448_7# _326_/a_543_7# _326_/a_1283_n19# _326_/a_1462_7# _326_/a_1270_373#
+ _326_/a_193_7# _326_/a_1217_7# _326_/a_761_249# _326_/a_27_7# _326_/a_1108_7# _326_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_257_ VGND VPWR VPWR VGND _260_/B _190_/A _254_/Y _258_/S _257_/a_448_7# _257_/a_544_257#
+ _257_/a_79_159# _257_/a_222_53# sky130_fd_sc_hd__o21ba_1
XFILLER_9_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_188_ VGND VPWR VPWR VGND _341_/D _255_/B _188_/S _307_/X _188_/a_505_n19# _188_/a_535_334#
+ _188_/a_76_159# _188_/a_218_334# _188_/a_439_7# _188_/a_218_7# sky130_fd_sc_hd__mux2_1
XFILLER_18_45 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_309_ VGND VPWR VPWR VGND _340_/CLK _309_/D _346_/SET_B _309_/Q _309_/a_639_7# _309_/a_805_7#
+ _309_/a_448_7# _309_/a_543_7# _309_/a_1283_n19# _309_/a_1462_7# _309_/a_1270_373#
+ _309_/a_193_7# _309_/a_1217_7# _309_/a_761_249# _309_/a_27_7# _309_/a_1108_7# _309_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput23 VGND VPWR VPWR VGND _316_/Q result[1] output23/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput34 VGND VPWR VPWR VGND _292_/A trim[3] output34/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput12 VGND VPWR VPWR VGND _281_/Y ctln[6] output12/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_11_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_290_ VPWR VGND VPWR VGND _290_/Y _290_/A sky130_fd_sc_hd__inv_2
Xrepeater42 VGND VPWR VPWR VGND repeater43/X _346_/SET_B repeater42/a_27_7# sky130_fd_sc_hd__buf_8
XFILLER_9_119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_12_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_273_ VPWR VGND VPWR VGND _273_/Y _273_/A sky130_fd_sc_hd__inv_2
XFILLER_5_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_342_ VGND VPWR VPWR VGND _343_/CLK _342_/D repeater43/X _342_/Q _342_/a_639_7# _342_/a_805_7#
+ _342_/a_448_7# _342_/a_543_7# _342_/a_1283_n19# _342_/a_1462_7# _342_/a_1270_373#
+ _342_/a_193_7# _342_/a_1217_7# _342_/a_761_249# _342_/a_27_7# _342_/a_1108_7# _342_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_4
X_325_ VGND VPWR VPWR VGND _331_/CLK _325_/D repeater43/X _325_/Q _325_/a_639_7# _325_/a_805_7#
+ _325_/a_448_7# _325_/a_543_7# _325_/a_1283_n19# _325_/a_1462_7# _325_/a_1270_373#
+ _325_/a_193_7# _325_/a_1217_7# _325_/a_761_249# _325_/a_27_7# _325_/a_1108_7# _325_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_187_ VGND VPWR VPWR VGND _255_/B _341_/Q _187_/a_27_7# sky130_fd_sc_hd__buf_1
X_256_ VGND VPWR VPWR VGND _260_/B _255_/X _191_/B _196_/A _192_/B _256_/a_209_7#
+ _256_/a_209_257# _256_/a_303_7# _256_/a_80_n19# sky130_fd_sc_hd__a31o_1
X_239_ VPWR VGND VPWR VGND _232_/X _328_/Q _319_/Q _240_/B _239_/a_199_7# _239_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
X_308_ VGND VPWR VPWR VGND _308_/X _227_/A _308_/S _192_/B _308_/a_505_n19# _308_/a_535_334#
+ _308_/a_76_159# _308_/a_218_334# _308_/a_439_7# _308_/a_218_7# sky130_fd_sc_hd__mux2_1
XFILLER_20_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_10_91 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput24 VGND VPWR VPWR VGND _317_/Q result[2] output24/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput13 VGND VPWR VPWR VGND _283_/Y ctln[7] output13/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput35 VGND VPWR VPWR VGND _294_/A trim[4] output35/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_16_135 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_127 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xrepeater43 VGND VPWR VPWR VGND input4/X repeater43/X repeater43/a_27_7# sky130_fd_sc_hd__buf_8
XFILLER_8_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_272_ VPWR VGND VPWR VGND _273_/A _326_/Q _317_/Q _272_/a_121_257# _272_/a_39_257#
+ sky130_fd_sc_hd__or2_2
X_341_ VGND VPWR VPWR VGND _343_/CLK _341_/D repeater43/X _341_/Q _341_/a_639_7# _341_/a_805_7#
+ _341_/a_448_7# _341_/a_543_7# _341_/a_1283_n19# _341_/a_1462_7# _341_/a_1270_373#
+ _341_/a_193_7# _341_/a_1217_7# _341_/a_761_249# _341_/a_27_7# _341_/a_1108_7# _341_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_10_108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_324_ VGND VPWR VPWR VGND _297_/B _324_/D repeater43/X _324_/Q _324_/a_639_7# _324_/a_805_7#
+ _324_/a_448_7# _324_/a_543_7# _324_/a_1283_n19# _324_/a_1462_7# _324_/a_1270_373#
+ _324_/a_193_7# _324_/a_1217_7# _324_/a_761_249# _324_/a_27_7# _324_/a_1108_7# _324_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_2_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_255_ VGND VPWR VPWR VGND _255_/B _298_/C _342_/Q _255_/X _255_/a_184_257# _255_/a_112_257#
+ _255_/a_30_13# sky130_fd_sc_hd__or3_2
X_186_ VGND VPWR VPWR VGND _308_/X _188_/S _172_/A _342_/D _186_/a_382_257# _186_/a_79_n19#
+ _186_/a_297_7# sky130_fd_sc_hd__o21a_1
XFILLER_18_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_238_ VGND VPWR VPWR VGND _242_/A _238_/B _320_/D _238_/a_109_257# sky130_fd_sc_hd__nor2_1
X_307_ VGND VPWR VPWR VGND _307_/X _145_/A _308_/S _296_/Y _307_/a_505_n19# _307_/a_535_334#
+ _307_/a_76_159# _307_/a_218_334# _307_/a_439_7# _307_/a_218_7# sky130_fd_sc_hd__mux2_1
X_169_ VGND VPWR VPWR VGND _172_/A _169_/B _169_/Y _169_/a_109_257# sky130_fd_sc_hd__nor2_1
XFILLER_19_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_13_8 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_28 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput14 VGND VPWR VPWR VGND _269_/A ctlp[0] output14/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_21_80 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xoutput36 VGND VPWR VPWR VGND _285_/Y trimb[0] output36/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput25 VGND VPWR VPWR VGND _318_/Q result[3] output25/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_22_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_0 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_13_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_271_ VPWR VGND VPWR VGND _271_/Y _271_/A sky130_fd_sc_hd__inv_2
X_340_ VGND VPWR VPWR VGND _340_/CLK _340_/D _346_/SET_B _340_/Q _340_/a_639_7# _340_/a_805_7#
+ _340_/a_448_7# _340_/a_543_7# _340_/a_1283_n19# _340_/a_1462_7# _340_/a_1270_373#
+ _340_/a_193_7# _340_/a_1217_7# _340_/a_761_249# _340_/a_27_7# _340_/a_1108_7# _340_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_185_ VPWR VGND VPWR VGND _343_/D _185_/A sky130_fd_sc_hd__inv_2
X_323_ VGND VPWR VPWR VGND _343_/CLK _323_/D repeater43/X _323_/Q _323_/a_639_7# _323_/a_805_7#
+ _323_/a_448_7# _323_/a_543_7# _323_/a_1283_n19# _323_/a_1462_7# _323_/a_1270_373#
+ _323_/a_193_7# _323_/a_1217_7# _323_/a_761_249# _323_/a_27_7# _323_/a_1108_7# _323_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_254_ VGND VPWR VPWR VGND _254_/A _254_/B _254_/Y _254_/a_109_257# sky130_fd_sc_hd__nor2_1
XFILLER_9_17 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_37 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_237_ VPWR VGND VPWR VGND _232_/X _329_/Q _320_/Q _238_/B _237_/a_199_7# _237_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
X_168_ VGND VPWR VPWR VGND _169_/B _167_/X _165_/X _167_/X _165_/X _168_/a_109_257#
+ _168_/a_397_257# _168_/a_109_7# _168_/a_481_7# sky130_fd_sc_hd__a2bb2oi_1
X_306_ VGND VPWR VPWR VGND _306_/X _286_/B _306_/S _294_/A _306_/a_505_n19# _306_/a_535_334#
+ _306_/a_76_159# _306_/a_218_334# _306_/a_439_7# _306_/a_218_7# sky130_fd_sc_hd__mux2_1
XFILLER_20_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_19_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput15 VGND VPWR VPWR VGND _271_/A ctlp[1] output15/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput26 VGND VPWR VPWR VGND _319_/Q result[4] output26/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput37 VGND VPWR VPWR VGND _288_/Y trimb[1] output37/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_16_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_1 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_2_3_0_clk VGND VPWR VPWR VGND _297_/B clkbuf_2_3_0_clk/A clkbuf_2_3_0_clk/a_75_172#
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_92 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_8_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_270_ VPWR VGND VPWR VGND _271_/A _325_/Q _316_/Q _270_/a_121_257# _270_/a_39_257#
+ sky130_fd_sc_hd__or2_2
X_322_ VGND VPWR VPWR VGND _331_/CLK _322_/D repeater43/X _322_/Q _322_/a_639_7# _322_/a_805_7#
+ _322_/a_448_7# _322_/a_543_7# _322_/a_1283_n19# _322_/a_1462_7# _322_/a_1270_373#
+ _322_/a_193_7# _322_/a_1217_7# _322_/a_761_249# _322_/a_27_7# _322_/a_1108_7# _322_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_253_ VPWR VGND VPWR VGND _254_/A _347_/Q sky130_fd_sc_hd__inv_2
XFILLER_13_82 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_184_ VGND VPWR VPWR VGND _185_/A _150_/C _188_/S _182_/X _184_/a_505_n19# _184_/a_535_334#
+ _184_/a_76_159# _184_/a_218_334# _184_/a_439_7# _184_/a_218_7# sky130_fd_sc_hd__mux2_1
X_236_ VGND VPWR VPWR VGND _242_/A _236_/B _321_/D _236_/a_109_257# sky130_fd_sc_hd__nor2_1
X_167_ VPWR VGND VPWR VGND _166_/Y _346_/Q _162_/X _167_/X _160_/X _167_/a_27_257#
+ _167_/a_109_257# _167_/a_373_7# _167_/a_109_7# sky130_fd_sc_hd__a22o_1
X_305_ VGND VPWR VPWR VGND _305_/X _286_/B _306_/S _254_/B _305_/a_505_n19# _305_/a_535_334#
+ _305_/a_76_159# _305_/a_218_334# _305_/a_439_7# _305_/a_218_7# sky130_fd_sc_hd__mux2_1
XFILLER_1_52 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_219_ VGND VPWR VPWR VGND _329_/D _216_/X _330_/Q _212_/X _217_/X _329_/Q _219_/a_584_7#
+ _219_/a_346_7# _219_/a_256_7# _219_/a_250_257# _219_/a_93_n19# sky130_fd_sc_hd__a32o_1
XFILLER_19_70 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput16 VGND VPWR VPWR VGND _273_/A ctlp[2] output16/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput38 VGND VPWR VPWR VGND _290_/Y trimb[2] output38/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput27 VGND VPWR VPWR VGND _320_/Q result[5] output27/a_27_7# sky130_fd_sc_hd__clkbuf_2
XPHY_2 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk VGND VPWR VPWR VGND clk clkbuf_0_clk/X clkbuf_0_clk/a_110_7# sky130_fd_sc_hd__clkbuf_16
XFILLER_7_62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_5_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_129 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_clk VGND VPWR VPWR VGND _340_/CLK clkbuf_2_3_0_clk/A clkbuf_2_2_0_clk/a_75_172#
+ sky130_fd_sc_hd__clkbuf_1
X_321_ VGND VPWR VPWR VGND _331_/CLK _321_/D repeater43/X _321_/Q _321_/a_639_7# _321_/a_805_7#
+ _321_/a_448_7# _321_/a_543_7# _321_/a_1283_n19# _321_/a_1462_7# _321_/a_1270_373#
+ _321_/a_193_7# _321_/a_1217_7# _321_/a_761_249# _321_/a_27_7# _321_/a_1108_7# _321_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_252_ VGND VPWR VPWR VGND _251_/X _228_/A _314_/D _297_/A _252_/a_109_257# _252_/a_27_7#
+ sky130_fd_sc_hd__o21ai_1
X_183_ VGND VPWR VPWR VGND _298_/A _188_/S _181_/X _324_/Q _150_/C _157_/A _183_/a_553_257#
+ _183_/a_1241_257# _183_/a_471_7# _183_/a_27_7# sky130_fd_sc_hd__o221ai_4
X_235_ VPWR VGND VPWR VGND _232_/X _330_/Q _321_/Q _236_/B _235_/a_199_7# _235_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
X_304_ VGND VPWR VPWR VGND _304_/S _227_/A _216_/X _304_/X _304_/a_257_159# _304_/a_306_329#
+ _304_/a_79_n19# _304_/a_578_7# _304_/a_591_329# _304_/a_288_7# sky130_fd_sc_hd__mux2_2
X_166_ VPWR VGND VPWR VGND _166_/Y _346_/Q sky130_fd_sc_hd__inv_2
X_218_ VGND VPWR VPWR VGND _330_/D _216_/X _304_/X _331_/Q _217_/X _330_/Q _218_/a_584_7#
+ _218_/a_346_7# _218_/a_256_7# _218_/a_250_257# _218_/a_93_n19# sky130_fd_sc_hd__a32o_1
XFILLER_19_82 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_149_ VGND VPWR VPWR VGND _149_/A _150_/C _149_/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput39 VGND VPWR VPWR VGND _292_/Y trimb[3] output39/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput17 VGND VPWR VPWR VGND _275_/A ctlp[3] output17/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput28 VGND VPWR VPWR VGND _321_/Q result[6] output28/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_16_128 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_50 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_320_ VGND VPWR VPWR VGND _297_/B _320_/D _346_/SET_B _320_/Q _320_/a_639_7# _320_/a_805_7#
+ _320_/a_448_7# _320_/a_543_7# _320_/a_1283_n19# _320_/a_1462_7# _320_/a_1270_373#
+ _320_/a_193_7# _320_/a_1217_7# _320_/a_761_249# _320_/a_27_7# _320_/a_1108_7# _320_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_73 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_251_ VGND VPWR VPWR VGND _251_/X _324_/Q _181_/X _172_/A _250_/X _251_/a_510_7#
+ _251_/a_79_n19# _251_/a_215_7# _251_/a_297_257# sky130_fd_sc_hd__o211a_1
X_182_ VGND VPWR VPWR VGND _182_/X _175_/Y _286_/B _196_/A _181_/X _182_/a_510_7#
+ _182_/a_79_n19# _182_/a_215_7# _182_/a_297_257# sky130_fd_sc_hd__o211a_1
XFILLER_18_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_234_ VGND VPWR VPWR VGND _242_/A _234_/B _322_/D _234_/a_109_257# sky130_fd_sc_hd__nor2_1
Xclkbuf_2_1_0_clk VGND VPWR VPWR VGND _331_/CLK clkbuf_2_1_0_clk/A clkbuf_2_1_0_clk/a_75_172#
+ sky130_fd_sc_hd__clkbuf_1
X_165_ VGND VPWR VPWR VGND _164_/Y _160_/X _158_/Y _161_/Y _165_/X _165_/a_78_159#
+ _165_/a_493_257# _165_/a_292_257# _165_/a_215_7# sky130_fd_sc_hd__o22a_1
X_303_ VPWR VGND VPWR VGND _347_/D _303_/A sky130_fd_sc_hd__inv_2
XFILLER_1_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_19_126 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_217_ VGND VPWR VPWR VGND _217_/A _217_/X _217_/a_27_7# sky130_fd_sc_hd__clkbuf_2
X_148_ VPWR VGND VPWR VGND _298_/B _341_/Q sky130_fd_sc_hd__inv_2
Xoutput18 VGND VPWR VPWR VGND _277_/A ctlp[4] output18/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput29 VGND VPWR VPWR VGND _322_/Q result[7] output29/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_21_73 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_4 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_12_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_181_ VGND VPWR VPWR VGND _215_/A _181_/X _181_/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_1_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_250_ VGND VPWR VPWR VGND _190_/A _216_/A _260_/A _284_/A _250_/X _250_/a_78_159#
+ _250_/a_493_257# _250_/a_292_257# _250_/a_215_7# sky130_fd_sc_hd__o22a_1
XFILLER_1_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_233_ VPWR VGND VPWR VGND _232_/X _331_/Q _322_/Q _234_/B _233_/a_199_7# _233_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
X_302_ VPWR VGND VPWR VGND _303_/A _157_/A _300_/Y _301_/X _147_/A _254_/A _302_/a_323_257#
+ _302_/a_227_7# _302_/a_227_257# _302_/a_77_159# _302_/a_539_257# sky130_fd_sc_hd__o32a_1
X_164_ VPWR VGND VPWR VGND _164_/Y _164_/A sky130_fd_sc_hd__inv_2
XFILLER_19_138 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_216_ VGND VPWR VPWR VGND _216_/A _216_/X _216_/a_27_7# sky130_fd_sc_hd__clkbuf_2
X_147_ VPWR VGND VPWR VGND _147_/Y _147_/A sky130_fd_sc_hd__inv_2
Xoutput19 VGND VPWR VPWR VGND _279_/A ctlp[5] output19/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_21_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xclkbuf_2_0_0_clk VGND VPWR VPWR VGND _343_/CLK clkbuf_2_1_0_clk/A clkbuf_2_0_0_clk/a_75_172#
+ sky130_fd_sc_hd__clkbuf_1
XPHY_5 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_7_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_21_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_16_85 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_107 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_77 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_180_ VPWR VGND VPWR VGND _298_/A _298_/B _298_/C _215_/A _180_/a_111_257# _180_/a_29_13#
+ _180_/a_183_257# sky130_fd_sc_hd__or3_1
XFILLER_1_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_232_ VGND VPWR VPWR VGND _232_/A _232_/X _232_/a_27_7# sky130_fd_sc_hd__clkbuf_2
X_163_ VGND VPWR VPWR VGND _162_/X _160_/A _158_/Y _345_/Q _164_/A _163_/a_78_159#
+ _163_/a_493_257# _163_/a_292_257# _163_/a_215_7# sky130_fd_sc_hd__o22a_1
X_301_ VGND VPWR VPWR VGND _162_/X _254_/A _347_/Q _160_/X _301_/X _299_/X _301_/a_149_7#
+ _301_/a_245_257# _301_/a_240_7# _301_/a_51_257# _301_/a_512_257# sky130_fd_sc_hd__o221a_1
XFILLER_19_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_146_ VPWR VGND VPWR VGND _147_/A _146_/C _341_/Q _177_/A _146_/a_184_13# _146_/a_29_271#
+ _146_/a_112_13# sky130_fd_sc_hd__and3_2
X_215_ VPWR VGND VPWR VGND _216_/A _215_/A sky130_fd_sc_hd__inv_2
XFILLER_21_42 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_6 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_7_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_21_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_101 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_231_ VPWR VGND VPWR VGND _232_/A _146_/C _255_/B _150_/C _162_/X _298_/A _231_/a_306_7#
+ _231_/a_79_n19# _231_/a_512_7# _231_/a_409_7# _231_/a_676_257# sky130_fd_sc_hd__o2111a_1
X_162_ VGND VPWR VPWR VGND _162_/A _162_/X _162_/a_27_7# sky130_fd_sc_hd__clkbuf_2
X_300_ VGND VPWR VPWR VGND _254_/A _160_/X _162_/X _347_/Q _300_/Y _299_/X _300_/a_27_257#
+ _300_/a_301_257# _300_/a_383_7# _300_/a_735_7# sky130_fd_sc_hd__a221oi_2
XFILLER_1_79 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
Xinput1 VGND VPWR VPWR VGND input1/X cal input1/a_75_172# sky130_fd_sc_hd__clkbuf_1
XFILLER_10_44 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_214_ VPWR VGND VPWR VGND _331_/Q _212_/X _181_/X _331_/D _217_/A _214_/a_27_257#
+ _214_/a_109_257# _214_/a_373_7# _214_/a_109_7# sky130_fd_sc_hd__a22o_1
X_145_ VGND VPWR VPWR VGND _145_/A _146_/C _304_/S _145_/a_113_7# sky130_fd_sc_hd__nand2_1
XFILLER_21_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_7 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_21_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_7_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_8_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_230_ VGND VPWR VPWR VGND _248_/A _242_/A _230_/a_27_7# sky130_fd_sc_hd__clkbuf_2
X_161_ VPWR VGND VPWR VGND _161_/Y _344_/Q sky130_fd_sc_hd__inv_2
XFILLER_1_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xinput2 VGND VPWR VPWR VGND _162_/A comp input2/a_27_7# sky130_fd_sc_hd__buf_1
XFILLER_10_67 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_19_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_213_ VPWR VGND VPWR VGND _217_/A _304_/X sky130_fd_sc_hd__inv_2
X_144_ VGND VPWR VPWR VGND _304_/S _144_/A _144_/a_27_7# sky130_fd_sc_hd__buf_1
XFILLER_21_99 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_8 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_21_136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_16_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_16_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_4_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_69 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_160_ VGND VPWR VPWR VGND _160_/A _160_/X _160_/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xinput3 VGND VPWR VPWR VGND en _227_/A input3/a_27_7# sky130_fd_sc_hd__clkbuf_2
X_289_ VPWR VGND VPWR VGND _290_/A _338_/Q _311_/Q _289_/a_121_257# _289_/a_39_257#
+ sky130_fd_sc_hd__or2_2
XFILLER_19_99 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_19_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_212_ VGND VPWR VPWR VGND _212_/X _304_/X _212_/a_27_7# sky130_fd_sc_hd__buf_1
X_143_ VGND VPWR VPWR VGND _144_/A _149_/A _341_/Q _177_/A _143_/a_27_7# _143_/a_109_7#
+ _143_/a_181_7# sky130_fd_sc_hd__and3_1
XFILLER_18_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_9 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_12_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_130 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_46 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_1_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_288_ VPWR VGND VPWR VGND _288_/Y _288_/A sky130_fd_sc_hd__inv_2
Xinput4 VGND VPWR VPWR VGND input4/X rstn input4/a_27_7# sky130_fd_sc_hd__buf_1
X_211_ VPWR VGND VPWR VGND _153_/B _332_/Q _206_/A _332_/D _197_/X _211_/a_27_257#
+ _211_/a_109_257# _211_/a_373_7# _211_/a_109_7# sky130_fd_sc_hd__a22o_1
X_142_ VPWR VGND VPWR VGND _149_/A _343_/Q sky130_fd_sc_hd__inv_2
XFILLER_10_58 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_15_102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_16_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_13_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_90 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_287_ VPWR VGND VPWR VGND _288_/A _337_/Q _310_/Q _287_/a_121_257# _287_/a_39_257#
+ sky130_fd_sc_hd__or2_2
XFILLER_19_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_210_ VGND VPWR VPWR VGND _153_/A _207_/C _306_/S _209_/X _333_/D _210_/a_109_257#
+ _210_/a_307_257# _210_/a_27_7# sky130_fd_sc_hd__o22ai_1
X_141_ VPWR VGND VPWR VGND _145_/A _227_/A sky130_fd_sc_hd__inv_2
X_339_ VGND VPWR VPWR VGND _340_/CLK _339_/D _346_/SET_B _339_/Q _339_/a_639_7# _339_/a_805_7#
+ _339_/a_448_7# _339_/a_543_7# _339_/a_1283_n19# _339_/a_1462_7# _339_/a_1270_373#
+ _339_/a_193_7# _339_/a_1217_7# _339_/a_761_249# _339_/a_27_7# _339_/a_1108_7# _339_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_12_128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_14_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_5_60 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_286_ VGND VPWR VPWR VGND _306_/S _286_/Y _286_/B _286_/a_113_7# sky130_fd_sc_hd__nand2_1
X_140_ VPWR VGND VPWR VGND _177_/A _342_/Q sky130_fd_sc_hd__inv_2
X_338_ VGND VPWR VPWR VGND _340_/CLK _338_/D _346_/SET_B _338_/Q _338_/a_639_7# _338_/a_805_7#
+ _338_/a_448_7# _338_/a_543_7# _338_/a_1283_n19# _338_/a_1462_7# _338_/a_1270_373#
+ _338_/a_193_7# _338_/a_1217_7# _338_/a_761_249# _338_/a_27_7# _338_/a_1108_7# _338_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_269_ VPWR VGND VPWR VGND _269_/Y _269_/A sky130_fd_sc_hd__inv_2
XFILLER_7_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_7_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_71 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_82 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_29 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_1_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_285_ VPWR VGND VPWR VGND _285_/Y _285_/A sky130_fd_sc_hd__inv_2
XFILLER_4_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_124 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_clk VGND VPWR VPWR VGND clkbuf_2_3_0_clk/A clkbuf_0_clk/X clkbuf_1_1_0_clk/a_75_172#
+ sky130_fd_sc_hd__clkbuf_1
X_268_ VPWR VGND VPWR VGND _269_/A _324_/Q _315_/Q _268_/a_121_257# _268_/a_39_257#
+ sky130_fd_sc_hd__or2_2
XFILLER_2_73 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_84 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_337_ VGND VPWR VPWR VGND _340_/CLK _337_/D _346_/SET_B _337_/Q _337_/a_639_7# _337_/a_805_7#
+ _337_/a_448_7# _337_/a_543_7# _337_/a_1283_n19# _337_/a_1462_7# _337_/a_1270_373#
+ _337_/a_193_7# _337_/a_1217_7# _337_/a_761_249# _337_/a_27_7# _337_/a_1108_7# _337_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_199_ VGND VPWR VPWR VGND _338_/D _193_/Y _197_/X _339_/Q _338_/Q _194_/X _199_/a_584_7#
+ _199_/a_346_7# _199_/a_256_7# _199_/a_250_257# _199_/a_93_n19# sky130_fd_sc_hd__a32o_1
XFILLER_21_49 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_123 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_4_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_13_17 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_40 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_95 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_284_ VPWR VGND VPWR VGND _285_/A _284_/A _309_/Q _284_/a_121_257# _284_/a_39_257#
+ sky130_fd_sc_hd__or2_2
XFILLER_19_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_18_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_198_ VGND VPWR VPWR VGND _339_/D _193_/Y _197_/X _340_/Q _339_/Q _194_/X _198_/a_584_7#
+ _198_/a_346_7# _198_/a_256_7# _198_/a_250_257# _198_/a_93_n19# sky130_fd_sc_hd__a32o_1
X_267_ VGND VPWR VPWR VGND _267_/A _267_/B _309_/D _267_/a_109_257# sky130_fd_sc_hd__nor2_1
X_336_ VGND VPWR VPWR VGND _340_/CLK _336_/D _346_/SET_B _336_/Q _336_/a_639_7# _336_/a_805_7#
+ _336_/a_448_7# _336_/a_543_7# _336_/a_1283_n19# _336_/a_1462_7# _336_/a_1270_373#
+ _336_/a_193_7# _336_/a_1217_7# _336_/a_761_249# _336_/a_27_7# _336_/a_1108_7# _336_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_319_ VGND VPWR VPWR VGND _297_/B _319_/D _346_/SET_B _319_/Q _319_/a_639_7# _319_/a_805_7#
+ _319_/a_448_7# _319_/a_543_7# _319_/a_1283_n19# _319_/a_1462_7# _319_/a_1270_373#
+ _319_/a_193_7# _319_/a_1217_7# _319_/a_761_249# _319_/a_27_7# _319_/a_1108_7# _319_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_0_0_clk VGND VPWR VPWR VGND clkbuf_2_1_0_clk/A clkbuf_0_clk/X clkbuf_1_0_0_clk/a_75_172#
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_4_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_83 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_283_ VPWR VGND VPWR VGND _283_/Y _283_/A sky130_fd_sc_hd__inv_2
XFILLER_18_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_335_ VGND VPWR VPWR VGND _343_/CLK _335_/D repeater43/X _335_/Q _335_/a_639_7# _335_/a_805_7#
+ _335_/a_448_7# _335_/a_543_7# _335_/a_1283_n19# _335_/a_1462_7# _335_/a_1270_373#
+ _335_/a_193_7# _335_/a_1217_7# _335_/a_761_249# _335_/a_27_7# _335_/a_1108_7# _335_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_197_ VGND VPWR VPWR VGND _260_/A _197_/X _197_/a_27_7# sky130_fd_sc_hd__clkbuf_2
X_266_ VPWR VGND VPWR VGND _258_/S _284_/A _309_/Q _267_/B _266_/a_199_7# _266_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
XFILLER_2_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_318_ VGND VPWR VPWR VGND _331_/CLK _318_/D repeater43/X _318_/Q _318_/a_639_7# _318_/a_805_7#
+ _318_/a_448_7# _318_/a_543_7# _318_/a_1283_n19# _318_/a_1462_7# _318_/a_1270_373#
+ _318_/a_193_7# _318_/a_1217_7# _318_/a_761_249# _318_/a_27_7# _318_/a_1108_7# _318_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_249_ VPWR VGND VPWR VGND _297_/A _314_/Q sky130_fd_sc_hd__inv_2
XFILLER_20_165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_20_110 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_114 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_282_ VPWR VGND VPWR VGND _283_/A _331_/Q _322_/Q _282_/a_121_257# _282_/a_39_257#
+ sky130_fd_sc_hd__or2_2
XFILLER_18_138 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_334_ VGND VPWR VPWR VGND _343_/CLK _334_/D repeater43/X _334_/Q _334_/a_639_7# _334_/a_805_7#
+ _334_/a_448_7# _334_/a_543_7# _334_/a_1283_n19# _334_/a_1462_7# _334_/a_1270_373#
+ _334_/a_193_7# _334_/a_1217_7# _334_/a_761_249# _334_/a_27_7# _334_/a_1108_7# _334_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_196_ VPWR VGND VPWR VGND _260_/A _196_/A sky130_fd_sc_hd__inv_2
X_265_ VGND VPWR VPWR VGND _267_/A _265_/B _310_/D _265_/a_109_257# sky130_fd_sc_hd__nor2_1
XFILLER_11_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_248_ VGND VPWR VPWR VGND _248_/A _248_/B _315_/D _248_/a_109_257# sky130_fd_sc_hd__nor2_1
X_317_ VGND VPWR VPWR VGND _331_/CLK _317_/D repeater43/X _317_/Q _317_/a_639_7# _317_/a_805_7#
+ _317_/a_448_7# _317_/a_543_7# _317_/a_1283_n19# _317_/a_1462_7# _317_/a_1270_373#
+ _317_/a_193_7# _317_/a_1217_7# _317_/a_761_249# _317_/a_27_7# _317_/a_1108_7# _317_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_179_ VGND VPWR VPWR VGND _191_/B _286_/B _179_/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_20_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_11_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_281_ VPWR VGND VPWR VGND _281_/Y _281_/A sky130_fd_sc_hd__inv_2
XPHY_40 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_195_ VPWR VGND VPWR VGND _340_/Q _306_/S _193_/Y _340_/D _194_/X _195_/a_27_257#
+ _195_/a_109_257# _195_/a_373_7# _195_/a_109_7# sky130_fd_sc_hd__a22o_1
X_333_ VGND VPWR VPWR VGND _343_/CLK _333_/D repeater43/X _333_/Q _333_/a_639_7# _333_/a_805_7#
+ _333_/a_448_7# _333_/a_543_7# _333_/a_1283_n19# _333_/a_1462_7# _333_/a_1270_373#
+ _333_/a_193_7# _333_/a_1217_7# _333_/a_761_249# _333_/a_27_7# _333_/a_1108_7# _333_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_4
X_264_ VPWR VGND VPWR VGND _258_/S _337_/Q _310_/Q _265_/B _264_/a_199_7# _264_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
X_316_ VGND VPWR VPWR VGND _331_/CLK _316_/D repeater43/X _316_/Q _316_/a_639_7# _316_/a_805_7#
+ _316_/a_448_7# _316_/a_543_7# _316_/a_1283_n19# _316_/a_1462_7# _316_/a_1270_373#
+ _316_/a_193_7# _316_/a_1217_7# _316_/a_761_249# _316_/a_27_7# _316_/a_1108_7# _316_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_247_ VPWR VGND VPWR VGND _232_/A _324_/Q _315_/Q _248_/B _247_/a_199_7# _247_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
XFILLER_11_64 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_134 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
X_178_ VPWR VGND VPWR VGND _298_/A _341_/Q _298_/C _191_/B _178_/a_109_257# _178_/a_27_7#
+ _178_/a_193_257# sky130_fd_sc_hd__or3_4
XFILLER_22_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_96 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_17_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_280_ VGND VPWR VPWR VGND _281_/A _330_/Q _321_/Q _280_/a_68_257# _280_/a_150_257#
+ sky130_fd_sc_hd__or2_1
XFILLER_14_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_332_ VGND VPWR VPWR VGND _340_/CLK _332_/D repeater43/X _332_/Q _332_/a_639_7# _332_/a_805_7#
+ _332_/a_448_7# _332_/a_543_7# _332_/a_1283_n19# _332_/a_1462_7# _332_/a_1270_373#
+ _332_/a_193_7# _332_/a_1217_7# _332_/a_761_249# _332_/a_27_7# _332_/a_1108_7# _332_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_4
X_194_ VGND VPWR VPWR VGND _194_/X _194_/A _194_/a_27_7# sky130_fd_sc_hd__buf_1
X_263_ VGND VPWR VPWR VGND _267_/A _263_/B _311_/D _263_/a_109_257# sky130_fd_sc_hd__nor2_1
XFILLER_11_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_246_ VGND VPWR VPWR VGND _248_/A _246_/B _316_/D _246_/a_109_257# sky130_fd_sc_hd__nor2_1
XFILLER_20_157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_20_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_315_ VGND VPWR VPWR VGND _343_/CLK _315_/D repeater43/X _315_/Q _315_/a_639_7# _315_/a_805_7#
+ _315_/a_448_7# _315_/a_543_7# _315_/a_1283_n19# _315_/a_1462_7# _315_/a_1270_373#
+ _315_/a_193_7# _315_/a_1217_7# _315_/a_761_249# _315_/a_27_7# _315_/a_1108_7# _315_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_177_ VGND VPWR VPWR VGND _177_/A _298_/A _177_/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_7_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_229_ VGND VPWR VPWR VGND input1/X _248_/A _226_/X _175_/Y _323_/D _229_/a_226_257#
+ _229_/a_76_159# _229_/a_556_7# _229_/a_226_7# _229_/a_489_373# sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_3_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_112 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_42 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_331_ VGND VPWR VPWR VGND _331_/CLK _331_/D repeater43/X _331_/Q _331_/a_639_7# _331_/a_805_7#
+ _331_/a_448_7# _331_/a_543_7# _331_/a_1283_n19# _331_/a_1462_7# _331_/a_1270_373#
+ _331_/a_193_7# _331_/a_1217_7# _331_/a_761_249# _331_/a_27_7# _331_/a_1108_7# _331_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
XPHY_31 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_193_ VPWR VGND VPWR VGND _193_/Y _194_/A sky130_fd_sc_hd__inv_2
X_262_ VPWR VGND VPWR VGND _258_/S _338_/Q _311_/Q _263_/B _262_/a_199_7# _262_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
XPHY_20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_2_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_6 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_245_ VPWR VGND VPWR VGND _232_/A _325_/Q _316_/Q _246_/B _245_/a_199_7# _245_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
XFILLER_14_133 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_122 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_314_ VGND VPWR VPWR VGND _297_/B _314_/D _346_/SET_B _314_/Q _314_/a_639_7# _314_/a_805_7#
+ _314_/a_448_7# _314_/a_543_7# _314_/a_1283_n19# _314_/a_1462_7# _314_/a_1270_373#
+ _314_/a_193_7# _314_/a_1217_7# _314_/a_761_249# _314_/a_27_7# _314_/a_1108_7# _314_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_176_ VGND VPWR VPWR VGND _298_/C _343_/Q _176_/a_27_7# sky130_fd_sc_hd__buf_1
XFILLER_22_54 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_0_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_159_ VPWR VGND VPWR VGND _160_/A _162_/A sky130_fd_sc_hd__inv_2
X_228_ VPWR VGND VPWR VGND _248_/A _228_/A sky130_fd_sc_hd__inv_2
XFILLER_17_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_65 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_5_68 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_43 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_330_ VGND VPWR VPWR VGND _331_/CLK _330_/D repeater43/X _330_/Q _330_/a_639_7# _330_/a_805_7#
+ _330_/a_448_7# _330_/a_543_7# _330_/a_1283_n19# _330_/a_1462_7# _330_/a_1270_373#
+ _330_/a_193_7# _330_/a_1217_7# _330_/a_761_249# _330_/a_27_7# _330_/a_1108_7# _330_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
XPHY_32 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_261_ VGND VPWR VPWR VGND _261_/A _267_/A _312_/D _261_/a_109_257# sky130_fd_sc_hd__nor2_1
XPHY_10 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_192_ VGND VPWR VPWR VGND _194_/A _305_/X _192_/B _192_/a_68_257# _192_/a_150_257#
+ sky130_fd_sc_hd__or2_1
XPHY_21 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_120 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_175_ VPWR VGND VPWR VGND _175_/Y _323_/Q sky130_fd_sc_hd__inv_2
X_244_ VGND VPWR VPWR VGND _248_/A _244_/B _317_/D _244_/a_109_257# sky130_fd_sc_hd__nor2_1
X_313_ VGND VPWR VPWR VGND _340_/CLK _313_/D _346_/SET_B _313_/Q _313_/a_639_7# _313_/a_805_7#
+ _313_/a_448_7# _313_/a_543_7# _313_/a_1283_n19# _313_/a_1462_7# _313_/a_1270_373#
+ _313_/a_193_7# _313_/a_1217_7# _313_/a_761_249# _313_/a_27_7# _313_/a_1108_7# _313_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_99 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_66 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_11_115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_158_ VPWR VGND VPWR VGND _158_/Y _345_/Q sky130_fd_sc_hd__inv_2
X_227_ VGND VPWR VPWR VGND _227_/A _228_/A _304_/S _227_/a_113_7# sky130_fd_sc_hd__nand2_1
XFILLER_3_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_125 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_12
XFILLER_5_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_5_47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_22 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_11 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_260_ VGND VPWR VPWR VGND _260_/B _267_/A _260_/A _260_/a_27_257# sky130_fd_sc_hd__nor2_2
XFILLER_2_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_191_ VGND VPWR VPWR VGND _323_/Q _191_/B _192_/B _191_/a_109_257# sky130_fd_sc_hd__nor2_1
X_243_ VPWR VGND VPWR VGND _232_/A _326_/Q _317_/Q _244_/B _243_/a_199_7# _243_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
X_312_ VGND VPWR VPWR VGND _340_/CLK _312_/D _346_/SET_B _312_/Q _312_/a_639_7# _312_/a_805_7#
+ _312_/a_448_7# _312_/a_543_7# _312_/a_1283_n19# _312_/a_1462_7# _312_/a_1270_373#
+ _312_/a_193_7# _312_/a_1217_7# _312_/a_761_249# _312_/a_27_7# _312_/a_1108_7# _312_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_174_ VPWR VGND VPWR VGND _161_/Y _344_/Q _172_/A _344_/D _147_/A _174_/a_27_257#
+ _174_/a_109_257# _174_/a_373_7# _174_/a_109_7# sky130_fd_sc_hd__a22o_1
XFILLER_22_78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_19_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_226_ VGND VPWR VPWR VGND _150_/C _225_/X _147_/A _226_/X _226_/a_382_257# _226_/a_79_n19#
+ _226_/a_297_7# sky130_fd_sc_hd__o21a_1
XFILLER_6_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_157_ VGND VPWR VPWR VGND _157_/A _172_/A _157_/a_27_7# sky130_fd_sc_hd__clkbuf_2
X_209_ VPWR VGND VPWR VGND _153_/A _333_/Q _332_/Q _209_/X _153_/B _209_/a_27_257#
+ _209_/a_109_257# _209_/a_373_7# _209_/a_109_7# sky130_fd_sc_hd__a22o_1
XFILLER_14_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_12 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_45 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_23 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X_190_ VGND VPWR VPWR VGND _190_/A _306_/S _190_/a_27_7# sky130_fd_sc_hd__clkbuf_2
X_242_ VGND VPWR VPWR VGND _242_/A _242_/B _318_/D _242_/a_109_257# sky130_fd_sc_hd__nor2_1
XFILLER_14_158 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_173_ VGND VPWR VPWR VGND _345_/Q _147_/Y _172_/Y _147_/Y _345_/D _173_/a_226_257#
+ _173_/a_76_159# _173_/a_556_7# _173_/a_226_7# _173_/a_489_373# sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_311_ VGND VPWR VPWR VGND _340_/CLK _311_/D _346_/SET_B _311_/Q _311_/a_639_7# _311_/a_805_7#
+ _311_/a_448_7# _311_/a_543_7# _311_/a_1283_n19# _311_/a_1462_7# _311_/a_1270_373#
+ _311_/a_193_7# _311_/a_1217_7# _311_/a_761_249# _311_/a_27_7# _311_/a_1108_7# _311_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_151 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_22_46 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_13 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_81 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_156_ VPWR VGND VPWR VGND _157_/A _196_/A _225_/B _156_/a_121_257# _156_/a_39_257#
+ sky130_fd_sc_hd__or2_2
X_225_ VPWR VGND VPWR VGND _225_/X _336_/Q _225_/B _225_/a_145_35# _225_/a_59_35#
+ sky130_fd_sc_hd__and2_1
X_208_ VGND VPWR VPWR VGND _207_/X _204_/Y _206_/A _334_/Q _334_/D _208_/a_78_159#
+ _208_/a_493_257# _208_/a_292_257# _208_/a_215_7# sky130_fd_sc_hd__o22a_1
XFILLER_0_105 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_58 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_70 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XPHY_35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_24 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_13 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_9_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_156 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_310_ VGND VPWR VPWR VGND _340_/CLK _310_/D _346_/SET_B _310_/Q _310_/a_639_7# _310_/a_805_7#
+ _310_/a_448_7# _310_/a_543_7# _310_/a_1283_n19# _310_/a_1462_7# _310_/a_1270_373#
+ _310_/a_193_7# _310_/a_1217_7# _310_/a_761_249# _310_/a_27_7# _310_/a_1108_7# _310_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
X_241_ VPWR VGND VPWR VGND _232_/X _327_/Q _318_/Q _242_/B _241_/a_199_7# _241_/a_113_257#
+ sky130_fd_sc_hd__a21oi_1
X_172_ VGND VPWR VPWR VGND _172_/A _172_/B _172_/Y _172_/a_109_257# sky130_fd_sc_hd__nor2_1
X_224_ VGND VPWR VPWR VGND _324_/D _216_/A _325_/Q _304_/X _217_/A _324_/Q _224_/a_584_7#
+ _224_/a_346_7# _224_/a_256_7# _224_/a_250_257# _224_/a_93_n19# sky130_fd_sc_hd__a32o_1
XFILLER_6_122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_155 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_8_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_155_ VPWR VGND VPWR VGND _225_/B _254_/B sky130_fd_sc_hd__inv_2
XFILLER_17_25 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_207_ VGND VPWR VPWR VGND _207_/X _207_/C _332_/Q _333_/Q _207_/a_27_7# _207_/a_109_7#
+ _207_/a_181_7# sky130_fd_sc_hd__and3_1
XFILLER_0_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_83 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_26 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_36 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_25 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_14 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_240_ VGND VPWR VPWR VGND _242_/A _240_/B _319_/D _240_/a_109_257# sky130_fd_sc_hd__nor2_1
X_171_ VGND VPWR VPWR VGND _164_/A _164_/Y _161_/Y _344_/Q _172_/B _171_/a_78_159#
+ _171_/a_493_257# _171_/a_292_257# _171_/a_215_7# sky130_fd_sc_hd__o22a_1
XFILLER_9_131 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_59 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_223_ VGND VPWR VPWR VGND _325_/D _216_/A _326_/Q _304_/X _217_/A _325_/Q _223_/a_584_7#
+ _223_/a_346_7# _223_/a_256_7# _223_/a_250_257# _223_/a_93_n19# sky130_fd_sc_hd__a32o_1
XFILLER_8_28 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_154_ VGND VPWR VPWR VGND _254_/B _154_/A _154_/a_27_7# sky130_fd_sc_hd__buf_1
X_206_ VPWR VGND VPWR VGND _207_/C _206_/A sky130_fd_sc_hd__inv_2
XFILLER_5_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_37 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_26 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_15 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_11_39 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_170_ VGND VPWR VPWR VGND _346_/Q _147_/Y _169_/Y _147_/Y _346_/D _170_/a_226_257#
+ _170_/a_76_159# _170_/a_556_7# _170_/a_226_7# _170_/a_489_373# sky130_fd_sc_hd__a2bb2o_1
X_299_ VGND VPWR VPWR VGND _167_/X _160_/X _166_/Y _165_/X _299_/X _299_/a_78_159#
+ _299_/a_493_257# _299_/a_292_257# _299_/a_215_7# sky130_fd_sc_hd__o22a_1
XFILLER_3_73 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_22_38 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_222_ VGND VPWR VPWR VGND _326_/D _216_/A _327_/Q _212_/X _217_/X _326_/Q _222_/a_584_7#
+ _222_/a_346_7# _222_/a_256_7# _222_/a_250_257# _222_/a_93_n19# sky130_fd_sc_hd__a32o_1
X_153_ VGND VPWR VPWR VGND _154_/A _334_/Q _335_/Q _153_/B _153_/A _153_/a_403_257#
+ _153_/a_215_257# _153_/a_487_257# _153_/a_109_53# _153_/a_297_257# sky130_fd_sc_hd__or4b_4
XFILLER_10_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
X_205_ VGND VPWR VPWR VGND _206_/A _204_/Y _335_/Q _335_/D _205_/a_382_257# _205_/a_79_n19#
+ _205_/a_297_7# sky130_fd_sc_hd__o21a_1
XFILLER_0_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_94 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_38 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_27 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_6_51 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_6_84 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_16 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_15_82 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_11_18 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_30 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_298_ VGND VPWR VPWR VGND _298_/X _298_/C _298_/B _298_/A _298_/a_27_7# _298_/a_109_7#
+ _298_/a_181_7# sky130_fd_sc_hd__and3_1
XFILLER_9_144 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_221_ VGND VPWR VPWR VGND _327_/D _216_/X _328_/Q _212_/X _217_/X _327_/Q _221_/a_584_7#
+ _221_/a_346_7# _221_/a_256_7# _221_/a_250_257# _221_/a_93_n19# sky130_fd_sc_hd__a32o_1
X_152_ VPWR VGND VPWR VGND _153_/B _332_/Q sky130_fd_sc_hd__inv_2
X_204_ VPWR VGND VPWR VGND _190_/A _204_/Y _333_/Q _332_/Q _334_/Q _204_/a_27_257#
+ _204_/a_27_7# _204_/a_277_7# sky130_fd_sc_hd__a31oi_2
XFILLER_3_117 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_3_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_0_75 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_18_93 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_3 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XPHY_28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_17 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_39 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_127 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_22_141 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_14_108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_13_163 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_297_ VGND VPWR VPWR VGND _297_/B _297_/Y _297_/A _297_/a_27_257# sky130_fd_sc_hd__nor2_2
X_220_ VGND VPWR VPWR VGND _328_/D _216_/X _329_/Q _212_/X _217_/X _328_/Q _220_/a_584_7#
+ _220_/a_346_7# _220_/a_256_7# _220_/a_250_257# _220_/a_93_n19# sky130_fd_sc_hd__a32o_1
X_151_ VPWR VGND VPWR VGND _153_/A _333_/Q sky130_fd_sc_hd__inv_2
XFILLER_6_115 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_100 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_133 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_10_144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_3_129 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_0_54 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_203_ VGND VPWR VPWR VGND _206_/A _298_/C _225_/B _336_/Q _147_/Y _203_/a_209_7#
+ _203_/a_209_257# _203_/a_303_7# _203_/a_80_n19# sky130_fd_sc_hd__a31o_1
XFILLER_9_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_41 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_6_97 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_17_106 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_29 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XPHY_18 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
XFILLER_17_139 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_95 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_51 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_16_161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_22_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_296_ VGND VPWR VPWR VGND _342_/Q _255_/B _296_/Y _306_/S _286_/B _284_/A _296_/a_213_83#
+ _296_/a_295_257# _296_/a_493_257# _296_/a_109_7# sky130_fd_sc_hd__o221ai_1
XFILLER_3_87 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
X_150_ VPWR VGND VPWR VGND _298_/B _150_/C _342_/Q _196_/A _150_/a_109_257# _150_/a_27_7#
+ _150_/a_193_257# sky130_fd_sc_hd__or3_4
X_279_ VPWR VGND VPWR VGND _279_/Y _279_/A sky130_fd_sc_hd__inv_2
XFILLER_17_7 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_202_ VGND VPWR VPWR VGND _336_/D _193_/Y _197_/X _337_/Q _284_/A _194_/X _202_/a_584_7#
+ _202_/a_346_7# _202_/a_256_7# _202_/a_250_257# _202_/a_93_n19# sky130_fd_sc_hd__a32o_1
XFILLER_0_88 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_8
XFILLER_9_9 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XPHY_19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
Xoutput40 VGND VPWR VPWR VGND _294_/Y trimb[4] output40/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_15_30 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput5 VGND VPWR VPWR VGND clkc _297_/Y output5/a_27_7# sky130_fd_sc_hd__buf_1
XFILLER_3_11 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_295_ VPWR VGND VPWR VGND _308_/S _181_/X _190_/A _286_/B _255_/B _342_/Q _295_/a_306_7#
+ _295_/a_79_n19# _295_/a_512_7# _295_/a_409_7# _295_/a_676_257# sky130_fd_sc_hd__o2111a_1
XFILLER_10_157 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_278_ VGND VPWR VPWR VGND _279_/A _329_/Q _320_/Q _278_/a_68_257# _278_/a_150_257#
+ sky130_fd_sc_hd__or2_1
X_347_ VGND VPWR VPWR VGND _297_/B _347_/D _346_/SET_B _347_/Q _347_/a_639_7# _347_/a_805_7#
+ _347_/a_448_7# _347_/a_543_7# _347_/a_1283_n19# _347_/a_1462_7# _347_/a_1270_373#
+ _347_/a_193_7# _347_/a_1217_7# _347_/a_761_249# _347_/a_27_7# _347_/a_1108_7# _347_/a_651_373#
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_2_153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_6
XFILLER_2_164 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
X_201_ VGND VPWR VPWR VGND _336_/Q _284_/A _201_/a_27_7# sky130_fd_sc_hd__clkbuf_2
XFILLER_9_54 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_9_87 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_86 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_53 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_20_3 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
XFILLER_15_75 VGND VPWR VPWR VGND sky130_fd_sc_hd__decap_4
Xoutput6 VGND VPWR VPWR VGND _269_/Y ctln[0] output6/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput41 VGND VPWR VPWR VGND _298_/X valid output41/a_27_7# sky130_fd_sc_hd__clkbuf_2
Xoutput30 VGND VPWR VPWR VGND _286_/Y sample output30/a_27_7# sky130_fd_sc_hd__clkbuf_2
X0 VGND VPWR.t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=233 ps=2.47k w=0 l=0
X1 VGND VPWR.t372 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X2 VPWR VGND.t249 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=355 ps=3.37k w=0 l=0
X3 VGND VPWR.t345 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X4 VPWR VGND.t87 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X5 VGND VPWR.t298 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X6 VPWR VGND.t74 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X7 VGND VPWR.t14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X8 VGND VPWR.t99 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X9 VPWR VGND.t375 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X10 VPWR VGND.t339 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X11 VGND VPWR.t32 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X12 VPWR VGND.t391 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X13 VGND VPWR.t61 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X14 VPWR VGND.t95 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X15 VGND VPWR.t120 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X16 VPWR VGND.t158 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X17 VGND VPWR.t347 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X18 VGND VPWR.t297 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X19 VGND VPWR.t86 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X20 VPWR VGND.t353 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X21 VPWR VGND.t61 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X22 VGND VPWR.t64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X23 VGND VPWR.t255 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X24 VPWR VGND.t251 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X25 VGND VPWR.t354 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X26 VGND clk.t4 clkbuf_0_clk/a_110_7# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0 l=0
X27 VPWR VGND.t93 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X28 VGND VPWR.t126 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X29 VPWR VGND.t26 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X30 VPWR VGND.t78 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X31 VGND VPWR.t66 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X32 VGND VPWR.t102 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X33 VPWR VGND.t383 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X34 VPWR VGND.t347 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X35 VGND VPWR.t339 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X36 VGND VPWR.t306 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X37 VPWR VGND.t236 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X38 VGND en.t1 input3/a_27_7# VGND sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0 l=0
X39 VGND VPWR.t17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X40 VPWR VGND.t168 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X41 VPWR VGND.t144 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X42 VGND VPWR.t165 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X43 VPWR VGND.t255 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X44 VPWR VGND.t354 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X45 VGND VPWR.t171 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X46 VPWR VGND.t256 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X47 VGND VPWR.t101 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X48 VGND VPWR.t382 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X49 VGND VPWR.t131 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X50 VPWR VGND.t191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X51 VPWR VGND.t308 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X52 VGND VPWR.t254 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X53 VPWR VGND.t17 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X54 VPWR VGND.t341 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X55 VGND VPWR.t114 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X56 VPWR VGND.t133 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X57 VGND VPWR.t344 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X58 VGND VPWR.t278 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X59 VGND VPWR.t141 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X60 VPWR VGND.t320 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X61 VPWR VGND.t187 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X62 VPWR VGND.t254 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X63 VPWR VGND.t245 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X64 VGND VPWR.t173 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X65 VGND VPWR.t276 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X66 VGND VPWR.t41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X67 VPWR VGND.t340 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X68 VPWR VGND.t59 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X69 VPWR VGND.t337 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X70 VPWR VGND.t83 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X71 VPWR VGND.t346 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X72 VGND VPWR.t388 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X73 VPWR VGND.t291 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X74 VGND VPWR.t224 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X75 VGND VPWR.t170 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X76 VPWR VGND.t276 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X77 VGND VPWR.t62 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X78 VGND VPWR.t140 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X79 VGND VPWR.t308 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X80 VGND VPWR.t15 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X81 VPWR VGND.t57 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X82 VPWR VGND.t388 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X83 VGND VPWR.t219 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X84 VGND VPWR.t129 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X85 VGND VPWR.t139 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X86 VPWR VGND.t192 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X87 VGND VPWR.t67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X88 VPWR VGND.t224 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X89 VPWR VGND.t62 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X90 VGND VPWR.t105 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X91 VGND VPWR.t187 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X92 VGND VPWR.t386 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X93 VPWR VGND.t311 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X94 VPWR VGND.t284 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X95 VPWR VGND.t207 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X96 VGND VPWR.t375 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X97 VPWR VGND.t219 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X98 VGND VPWR.t59 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X99 VPWR VGND.t194 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X100 VGND VPWR.t337 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X101 VPWR VGND.t67 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X102 VPWR VGND.t367 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X103 VPWR VGND.t315 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X104 VGND VPWR.t261 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X105 VPWR VGND.t0 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X106 VPWR VGND.t121 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X107 VPWR VGND.t292 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X108 VPWR VGND.t372 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X109 VPWR VGND.t289 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X110 VPWR VGND.t286 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X111 VPWR VGND.t123 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X112 VPWR VGND.t376 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X113 VPWR VGND.t274 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X114 VPWR VGND.t153 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X115 VGND VPWR.t342 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X116 VPWR VGND.t261 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X117 VGND VPWR.t10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X118 VPWR VGND.t81 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X119 VGND VPWR.t182 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X120 VGND VPWR.t317 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X121 VPWR VGND.t230 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X122 VGND VPWR.t98 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X123 VPWR VGND.t235 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X124 VPWR VGND.t225 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X125 VPWR VGND.t32 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X126 VGND VPWR.t289 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X127 VPWR VGND.t82 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X128 VGND VPWR.t383 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X129 VGND VPWR.t284 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X130 VPWR VGND.t10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X131 VGND VPWR.t20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X132 VGND VPWR.t194 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X133 VGND VPWR.t263 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X134 VPWR VGND.t98 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X135 VPWR VGND.t120 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X136 VGND VPWR.t54 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X137 VPWR VGND.t366 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X138 VGND VPWR.t203 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X139 VPWR VGND.t199 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X140 VPWR VGND.t231 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X141 VPWR VGND.t20 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X142 VPWR VGND.t40 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X143 VGND VPWR.t56 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X144 VGND VPWR.t153 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X145 VPWR VGND.t126 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X146 VGND VPWR.t321 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X147 VGND VPWR.t299 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X148 VGND VPWR.t178 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X149 VGND VPWR.t42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X150 VPWR VGND.t54 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X151 VGND VPWR.t336 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X152 VPWR VGND.t294 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X153 VPWR VGND.t58 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X154 VGND VPWR.t353 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X155 VGND VPWR.t269 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X156 VGND VPWR.t212 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X157 VGND VPWR.t162 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X158 VGND VPWR.t124 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X159 VPWR VGND.t171 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X160 VPWR VGND.t299 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X161 VPWR VGND.t252 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X162 VPWR VGND.t97 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X163 VGND VPWR.t319 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X164 VGND VPWR.t83 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X165 VPWR VGND.t101 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X166 VPWR VGND.t132 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X167 VGND VPWR.t346 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X168 VPWR VGND.t269 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X169 VGND VPWR.t378 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X170 VPWR VGND.t212 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X171 VPWR VGND.t107 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X172 VGND VPWR.t356 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X173 VGND VPWR.t366 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X174 VPWR VGND.t162 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X175 VGND VPWR.t12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X176 VGND VPWR.t227 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X177 VPWR VGND.t14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X178 VGND VPWR.t89 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X179 VPWR VGND.t152 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X180 VGND VPWR.t60 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X181 VPWR VGND.t173 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X182 VGND VPWR.t104 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X183 VGND VPWR.t282 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X184 VPWR VGND.t324 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X185 VGND VPWR.t58 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X186 VGND VPWR.t175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X187 VPWR VGND.t227 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X188 VPWR VGND.t183 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X189 VPWR VGND.t297 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X190 VGND VPWR.t207 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X191 VPWR VGND.t92 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X192 VGND VPWR.t312 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X193 VPWR VGND.t312 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X194 VGND VPWR.t201 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X195 VGND VPWR.t127 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X196 VGND VPWR.t179 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X197 VGND VPWR.t34 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X198 VGND VPWR.t43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X199 VGND VPWR.t121 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X200 VPWR VGND.t66 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X201 VPWR VGND.t102 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X202 VGND VPWR.t122 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X203 VGND VPWR.t125 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X204 VPWR VGND.t279 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X205 VGND VPWR.t273 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X206 VGND VPWR.t274 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X207 VPWR VGND.t165 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X208 VPWR VGND.t35 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X209 VGND VPWR.t152 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X210 VPWR VGND.t164 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X211 VGND VPWR.t296 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X212 VGND VPWR.t230 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X213 VPWR VGND.t11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X214 VPWR VGND.t273 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X215 VGND VPWR.t264 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X216 VPWR VGND.t302 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X217 VGND VPWR.t183 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X218 VPWR VGND.t344 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X219 VPWR VGND.t382 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X220 VPWR VGND.t296 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X221 VPWR VGND.t278 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X222 VGND VPWR.t92 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X223 VPWR VGND.t99 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X224 VPWR VGND.t151 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X225 VPWR VGND.t163 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X226 VGND VPWR.t365 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X227 VPWR VGND.t86 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X228 VGND VPWR.t199 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X229 VGND VPWR.t307 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X230 VGND VPWR.t143 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X231 VPWR VGND.t154 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X232 VPWR VGND.t244 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X233 VPWR VGND.t223 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X234 VPWR VGND.t264 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X235 VGND VPWR.t53 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X236 VGND VPWR.t151 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X237 VPWR VGND.t170 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X238 VGND VPWR.t352 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X239 VGND VPWR.t163 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X240 VPWR VGND.t386 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X241 VPWR VGND.t15 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X242 VPWR VGND.t155 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X243 VPWR VGND.t129 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X244 VPWR VGND.t139 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X245 VPWR VGND.t53 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X246 VGND VPWR.t63 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X247 VPWR VGND.t141 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X248 VGND VPWR.t154 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X249 VPWR VGND.t336 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X250 VGND VPWR.t9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X251 VGND VPWR.t303 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X252 VPWR VGND.t105 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X253 VGND VPWR.t268 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X254 VGND VPWR.t324 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X255 VGND VPWR.t313 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X256 VPWR VGND.t184 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X257 VGND VPWR.t72 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X258 VPWR VGND.t342 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X259 VPWR VGND.t9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X260 VGND VPWR.t327 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X261 VPWR VGND.t275 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X262 VGND VPWR.t247 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X263 VPWR VGND.t356 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X264 VPWR VGND.t268 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X265 VPWR VGND.t182 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X266 VPWR VGND.t313 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X267 VPWR VGND.t41 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X268 VGND VPWR.t38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X269 VGND VPWR.t103 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X270 VPWR VGND.t72 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X271 VPWR VGND.t140 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X272 VGND VPWR.t380 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X273 VGND VPWR.t80 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X274 VGND VPWR.t155 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X275 VPWR VGND.t185 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X276 VGND VPWR.t279 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X277 VGND VPWR.t166 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X278 VGND VPWR.t221 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X279 VGND VPWR.t35 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X280 VGND VPWR.t326 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X281 VGND VPWR.t11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X282 VGND VPWR.t184 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X283 VPWR VGND.t203 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X284 VPWR VGND.t332 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X285 VGND VPWR.t116 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X286 VPWR VGND.t169 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X287 VPWR VGND.t263 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X288 VPWR VGND.t309 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X289 VGND VPWR.t300 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X290 VPWR VGND.t323 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X291 VPWR VGND.t321 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X292 VPWR VGND.t204 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X293 VGND VPWR.t21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X294 VGND VPWR.t128 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X295 VPWR VGND.t100 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X296 VPWR VGND.t125 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X297 VGND VPWR.t206 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X298 VGND VPWR.t157 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X299 VGND VPWR.t174 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X300 VGND VPWR.t214 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X301 VGND VPWR.t134 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X302 VPWR VGND.t338 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X303 VGND VPWR.t185 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X304 VGND VPWR.t130 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X305 VGND VPWR.t232 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X306 VGND VPWR.t193 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X307 VGND VPWR.t110 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X308 VPWR VGND.t206 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X309 VPWR VGND.t378 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X310 VGND VPWR.t147 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X311 VGND VPWR.t244 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X312 VPWR VGND.t12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X313 VGND VPWR.t371 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X314 VPWR VGND.t301 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X315 VGND VPWR.t169 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X316 VPWR VGND.t317 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X317 VGND VPWR.t172 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X318 VPWR VGND.t50 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X319 VPWR VGND.t89 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X320 VGND VPWR.t223 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X321 VGND VPWR.t215 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X322 VPWR VGND.t357 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X323 VGND VPWR.t323 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X324 VGND VPWR.t309 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X325 VGND VPWR.t204 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X326 VGND VPWR.t200 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X327 VPWR VGND.t365 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X328 VPWR VGND.t143 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X329 VPWR VGND.t272 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X330 VPWR VGND.t262 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X331 VPWR VGND.t56 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X332 VPWR VGND.t172 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X333 VGND VPWR.t338 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X334 VGND VPWR.t213 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X335 VPWR VGND.t215 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X336 VPWR VGND.t240 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X337 VGND VPWR.t305 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X338 VGND VPWR.t51 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X339 VPWR VGND.t127 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X340 VPWR VGND.t122 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X341 VGND VPWR.t368 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X342 VPWR VGND.t228 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X343 VGND VPWR.t5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X344 VPWR VGND.t213 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X345 VGND VPWR.t348 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X346 VGND VPWR.t301 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X347 VPWR VGND.t178 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X348 VPWR VGND.t42 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X349 VGND VPWR.t50 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X350 VGND VPWR.t384 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X351 VPWR VGND.t201 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X352 VPWR VGND.t195 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X353 VGND VPWR.t357 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X354 VGND VPWR.t275 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X355 VPWR VGND.t5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X356 VGND VPWR.t176 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X357 VPWR VGND.t124 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X358 VPWR VGND.t146 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X359 VPWR VGND.t348 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X360 VGND VPWR.t242 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X361 VPWR VGND.t222 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X362 VGND VPWR.t46 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X363 VPWR VGND.t63 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X364 VPWR VGND.t60 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X365 VPWR VGND.t384 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X366 VPWR VGND.t104 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X367 VGND VPWR.t111 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X368 VPWR VGND.t282 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X369 VGND VPWR.t208 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X370 VPWR VGND.t175 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X371 VPWR VGND.t242 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X372 VPWR VGND.t46 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X373 VGND VPWR.t246 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X374 VGND VPWR.t239 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X375 VGND VPWR.t253 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X376 VGND VPWR.t106 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X377 VGND VPWR.t216 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X378 VPWR VGND.t380 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X379 VGND VPWR.t100 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X380 VGND VPWR.t146 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X381 VGND VPWR.t167 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X382 VGND VPWR.t16 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X383 VGND VPWR.t222 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X384 VPWR VGND.t253 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X385 VPWR VGND.t106 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X386 VPWR VGND.t179 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X387 VPWR VGND.t216 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X388 VPWR VGND.t34 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X389 VPWR VGND.t326 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X390 VPWR VGND.t319 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X391 VPWR VGND.t43 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X392 clkbuf_0_clk/a_110_7# clk.t1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=0 l=0
X393 VGND VPWR.t363 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X394 VPWR VGND.t31 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X395 VPWR VGND.t16 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X396 VGND VPWR.t33 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X397 VGND VPWR.t314 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X398 input1/a_75_172# cal.t1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0 l=0
X399 VPWR VGND.t21 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X400 VGND VPWR.t318 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X401 VGND VPWR.t228 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X402 VPWR VGND.t28 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X403 VPWR rstn.t0 input4/a_27_7# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0 l=0
X404 VGND VPWR.t36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X405 VPWR VGND.t290 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X406 VGND VPWR.t280 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X407 VPWR VGND.t33 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X408 VGND VPWR.t359 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X409 VPWR VGND.t314 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X410 VGND VPWR.t272 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X411 VPWR VGND.t241 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X412 VGND VPWR.t377 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X413 VGND VPWR.t262 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X414 VPWR en.t0 input3/a_27_7# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=0 l=0
X415 VGND VPWR.t8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X416 VPWR VGND.t327 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X417 VGND VPWR.t96 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X418 VGND VPWR.t328 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X419 VPWR VGND.t280 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X420 VGND VPWR.t240 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X421 VGND VPWR.t31 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X422 VGND rstn.t1 input4/a_27_7# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0 l=0
X423 VPWR VGND.t371 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X424 VPWR VGND.t307 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X425 VPWR VGND.t103 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X426 VPWR VGND.t377 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X427 VGND VPWR.t119 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X428 VGND VPWR.t385 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X429 VPWR VGND.t247 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X430 VPWR VGND.t166 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X431 VGND VPWR.t373 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X432 VPWR VGND.t352 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X433 VPWR VGND.t221 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X434 VGND VPWR.t70 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X435 VPWR VGND.t385 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X436 VGND VPWR.t257 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X437 VPWR VGND.t116 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X438 VGND VPWR.t335 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X439 VPWR VGND.t304 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X440 VPWR VGND.t373 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X441 VGND VPWR.t24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X442 VGND VPWR.t325 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X443 VPWR VGND.t128 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X444 VGND VPWR.t18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X445 VPWR VGND.t136 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X446 VPWR VGND.t157 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X447 VPWR VGND.t214 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X448 VGND VPWR.t210 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X449 VPWR VGND.t134 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X450 VPWR VGND.t306 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X451 VGND VPWR.t229 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X452 VPWR VGND.t24 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X453 VPWR VGND.t303 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X454 VGND VPWR.t238 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X455 VPWR VGND.t325 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X456 VPWR VGND.t193 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X457 VPWR VGND.t38 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X458 VPWR VGND.t110 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X459 VGND VPWR.t112 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X460 VGND VPWR.t333 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X461 VPWR VGND.t210 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X462 VGND VPWR.t55 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X463 VGND VPWR.t260 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X464 VPWR VGND.t80 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X465 VGND VPWR.t311 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X466 VPWR VGND.t238 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X467 VGND VPWR.t150 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X468 VGND VPWR.t304 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X469 VGND VPWR.t364 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X470 VGND VPWR.t2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X471 VPWR VGND.t112 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X472 VPWR VGND.t333 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X473 VGND VPWR.t161 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X474 VPWR VGND.t246 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X475 VGND VPWR.t350 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X476 VGND VPWR.t281 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X477 VGND VPWR.t136 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X478 VPWR VGND.t161 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X479 VGND VPWR.t28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X480 VGND VPWR.t69 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X481 VGND VPWR.t160 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X482 VPWR VGND.t167 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X483 VGND VPWR.t360 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X484 VPWR VGND.t305 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X485 VGND VPWR.t197 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X486 VGND VPWR.t379 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X487 VPWR VGND.t281 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X488 VGND VPWR.t73 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X489 VPWR VGND.t27 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X490 VPWR VGND.t300 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X491 VGND VPWR.t90 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X492 VGND VPWR.t241 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X493 VPWR VGND.t130 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X494 VPWR VGND.t51 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X495 VPWR VGND.t73 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X496 VPWR VGND.t174 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X497 VGND VPWR.t94 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X498 VPWR VGND.t147 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X499 VGND VPWR.t195 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X500 VPWR VGND.t229 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X501 VGND VPWR.t1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X502 VGND VPWR.t234 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X503 VPWR VGND.t232 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X504 clkbuf_0_clk/a_110_7# clk.t3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=0 l=0
X505 VPWR VGND.t200 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X506 VGND VPWR.t13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X507 VPWR VGND.t94 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X508 VGND VPWR.t209 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X509 VGND VPWR.t7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X510 VGND VPWR.t148 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X511 VGND VPWR.t322 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X512 VGND VPWR.t47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X513 VPWR VGND.t76 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X514 VGND VPWR.t27 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X515 VPWR VGND.t8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X516 VGND VPWR.t79 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X517 VPWR VGND.t239 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X518 VGND VPWR.t358 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X519 VGND VPWR.t19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X520 VPWR VGND.t7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X521 VPWR VGND.t148 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X522 VPWR VGND.t209 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X523 VPWR VGND.t322 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X524 VGND VPWR.t77 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X525 VPWR VGND.t198 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X526 VGND VPWR.t362 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X527 VGND VPWR.t387 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X528 VGND VPWR.t49 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X529 VGND VPWR.t250 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X530 VGND VPWR.t138 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X531 VGND VPWR.t117 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X532 VGND VPWR.t156 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X533 VPWR VGND.t368 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X534 VPWR VGND.t329 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X535 VPWR VGND.t70 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X536 VPWR VGND.t176 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X537 VPWR VGND.t362 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X538 VPWR VGND.t363 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X539 VGND VPWR.t76 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X540 VPWR VGND.t113 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X541 VPWR VGND.t250 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X542 VGND VPWR.t302 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X543 VPWR VGND.t45 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X544 VGND VPWR.t355 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X545 VPWR VGND.t318 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X546 VPWR VGND.t111 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X547 VGND VPWR.t189 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X548 VPWR comp.t0 input2/a_27_7# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0 l=0
X549 VPWR VGND.t36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X550 VGND VPWR.t39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X551 VPWR VGND.t65 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X552 VGND VPWR.t237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X553 VGND VPWR.t220 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X554 VPWR VGND.t208 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X555 VPWR VGND.t3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X556 clkbuf_0_clk/a_110_7# clk.t5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0 l=0
X557 VGND VPWR.t218 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X558 VPWR VGND.t189 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X559 VGND VPWR.t186 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X560 VPWR VGND.t328 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X561 VPWR VGND.t359 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X562 VGND VPWR.t367 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X563 VGND VPWR.t331 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X564 VGND VPWR.t113 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X565 VPWR VGND.t237 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X566 VPWR clk.t6 clkbuf_0_clk/a_110_7# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=0 l=0
X567 VGND comp.t1 input2/a_27_7# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0 l=0
X568 VPWR VGND.t370 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X569 VPWR VGND.t2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X570 VPWR VGND.t287 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X571 VPWR VGND.t259 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X572 VGND VPWR.t109 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X573 VGND VPWR.t65 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X574 VGND VPWR.t334 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X575 VGND VPWR.t349 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X576 VGND VPWR.t295 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X577 VPWR VGND.t197 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X578 VGND VPWR.t271 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X579 VGND VPWR.t256 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X580 VPWR VGND.t44 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X581 VGND VPWR.t159 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X582 VPWR VGND.t265 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X583 VPWR VGND.t18 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X584 VGND VPWR.t142 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X585 VPWR VGND.t349 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X586 VGND VPWR.t390 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X587 VPWR VGND.t295 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X588 VPWR VGND.t30 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X589 VGND VPWR.t287 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X590 VPWR VGND.t205 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X591 VPWR VGND.t96 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X592 VPWR VGND.t1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X593 VPWR VGND.t390 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X594 VPWR VGND.t115 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X595 VPWR VGND.t142 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X596 VPWR VGND.t234 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X597 VGND VPWR.t332 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X598 VPWR VGND.t55 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X599 VGND VPWR.t198 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X600 VGND VPWR.t217 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X601 VGND VPWR.t88 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X602 VPWR VGND.t119 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X603 VPWR VGND.t180 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X604 VPWR VGND.t285 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X605 VPWR VGND.t364 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X606 VGND VPWR.t251 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X607 VGND VPWR.t181 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X608 VPWR VGND.t257 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X609 VGND VPWR.t369 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X610 VGND VPWR.t329 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X611 VGND VPWR.t26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X612 VGND VPWR.t158 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X613 VGND VPWR.t75 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X614 VPWR VGND.t335 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X615 VGND VPWR.t293 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X616 VGND VPWR.t243 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X617 VGND VPWR.t226 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X618 VGND VPWR.t190 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X619 VGND VPWR.t205 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X620 VGND VPWR.t45 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X621 VGND VPWR.t71 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X622 VPWR VGND.t77 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X623 VGND VPWR.t249 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X624 VPWR VGND.t75 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X625 VPWR VGND.t379 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X626 VPWR VGND.t49 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X627 VPWR VGND.t243 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X628 VPWR VGND.t226 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X629 VGND VPWR.t115 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X630 VGND VPWR.t196 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X631 VPWR VGND.t190 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X632 VGND VPWR.t316 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X633 VPWR VGND.t71 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X634 VGND VPWR.t285 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X635 VGND VPWR.t23 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X636 VPWR VGND.t360 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X637 VGND VPWR.t3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X638 VGND VPWR.t52 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X639 VPWR clk.t0 clkbuf_0_clk/a_110_7# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=0 l=0
X640 input1/a_75_172# cal.t0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0 l=0
X641 VGND VPWR.t145 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X642 VGND VPWR.t191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X643 VPWR VGND.t283 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X644 VGND VPWR.t370 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X645 VPWR VGND.t316 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X646 VPWR VGND.t260 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X647 VGND VPWR.t288 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X648 VPWR VGND.t23 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X649 VPWR VGND.t137 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X650 VPWR VGND.t343 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X651 VGND VPWR.t95 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X652 VPWR VGND.t52 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X653 VPWR VGND.t351 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X654 VGND VPWR.t245 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X655 VGND VPWR.t259 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X656 VGND VPWR.t4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X657 VPWR VGND.t150 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X658 VPWR VGND.t288 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X659 VGND VPWR.t233 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X660 VPWR VGND.t79 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X661 VPWR VGND.t25 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X662 VPWR VGND.t19 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X663 VPWR VGND.t69 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X664 VGND VPWR.t78 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X665 VPWR VGND.t4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X666 VGND VPWR.t44 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X667 VPWR VGND.t47 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X668 VPWR VGND.t160 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X669 VPWR VGND.t350 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X670 VGND VPWR.t149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X671 VGND VPWR.t236 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X672 VGND VPWR.t283 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X673 VPWR VGND.t233 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X674 VPWR VGND.t381 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X675 clkbuf_0_clk/a_110_7# clk.t7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0 l=0
X676 VPWR VGND.t90 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X677 VGND VPWR.t168 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X678 VPWR VGND.t387 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X679 VGND VPWR.t265 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X680 VPWR VGND.t358 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X681 VGND VPWR.t290 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X682 VPWR VGND.t138 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X683 VGND VPWR.t374 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X684 VGND VPWR.t30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X685 VGND VPWR.t137 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X686 VGND VPWR.t315 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X687 VPWR VGND.t149 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X688 VPWR VGND.t156 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X689 VGND VPWR.t292 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X690 VPWR VGND.t135 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X691 VGND VPWR.t351 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X692 VPWR VGND.t361 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X693 VGND VPWR.t341 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X694 VGND VPWR.t286 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X695 VGND VPWR.t133 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X696 VPWR VGND.t374 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X697 VGND VPWR.t391 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X698 VGND VPWR.t320 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X699 VGND VPWR.t180 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X700 VGND VPWR.t177 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X701 VGND VPWR.t85 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X702 VPWR VGND.t345 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X703 VPWR VGND.t39 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X704 VGND VPWR.t123 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X705 VPWR VGND.t298 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X706 VGND VPWR.t291 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X707 VPWR VGND.t13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X708 VPWR VGND.t84 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X709 VGND VPWR.t258 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X710 VPWR VGND.t220 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X711 VPWR VGND.t218 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X712 VPWR VGND.t177 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X713 VGND VPWR.t48 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X714 VPWR VGND.t85 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X715 VGND VPWR.t93 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X716 VPWR VGND.t186 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X717 VGND VPWR.t135 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X718 VGND VPWR.t270 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X719 VGND VPWR.t118 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X720 VGND VPWR.t266 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X721 VPWR VGND.t258 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X722 VPWR VGND.t117 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X723 VGND VPWR.t192 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X724 VGND VPWR.t6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X725 VPWR VGND.t48 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X726 VGND VPWR.t144 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X727 VPWR VGND.t310 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X728 VGND VPWR.t37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X729 VPWR VGND.t331 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X730 VPWR VGND.t270 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X731 VPWR VGND.t109 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X732 VPWR VGND.t118 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X733 VGND VPWR.t188 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X734 VPWR VGND.t266 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X735 VPWR VGND.t64 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X736 VGND VPWR.t330 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X737 VGND VPWR.t267 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X738 VGND VPWR.t211 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X739 VGND VPWR.t389 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X740 VPWR VGND.t334 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X741 VPWR VGND.t6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X742 VGND VPWR.t84 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X743 VPWR VGND.t37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X744 VGND VPWR.t91 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X745 VGND VPWR.t376 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X746 VGND VPWR.t252 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X747 VGND VPWR.t29 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X748 VPWR VGND.t271 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X749 VGND VPWR.t343 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X750 VGND clk.t2 clkbuf_0_clk/a_110_7# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0 l=0
X751 VPWR VGND.t188 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X752 VGND VPWR.t68 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X753 VPWR VGND.t196 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X754 VPWR VGND.t211 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X755 VPWR VGND.t389 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X756 VPWR VGND.t330 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X757 VPWR VGND.t267 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X758 VPWR VGND.t355 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X759 VPWR VGND.t91 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X760 VGND VPWR.t97 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X761 VGND VPWR.t340 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X762 VGND VPWR.t277 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X763 VPWR VGND.t29 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X764 VGND VPWR.t81 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X765 VGND VPWR.t132 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X766 VPWR VGND.t131 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X767 VGND VPWR.t235 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X768 VGND VPWR.t225 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X769 VPWR VGND.t145 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X770 VGND VPWR.t25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X771 VGND VPWR.t310 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X772 VGND VPWR.t22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X773 VPWR VGND.t68 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X774 VGND VPWR.t82 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X775 VGND VPWR.t107 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X776 VPWR VGND.t114 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X777 VPWR VGND.t277 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X778 VGND VPWR.t231 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X779 VGND VPWR.t381 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X780 VGND VPWR.t248 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X781 VPWR VGND.t217 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X782 VGND VPWR.t57 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X783 VPWR VGND.t88 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X784 VGND VPWR.t108 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X785 VPWR VGND.t22 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X786 VPWR VGND.t181 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X787 VGND VPWR.t202 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X788 VPWR VGND.t369 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X789 VGND VPWR.t40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X790 VGND VPWR.t361 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X791 VPWR VGND.t248 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X792 VPWR VGND.t293 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X793 VGND VPWR.t87 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X794 VPWR VGND.t108 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X795 VGND VPWR.t74 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X796 VGND VPWR.t294 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X797 VPWR VGND.t159 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
X798 VGND VPWR.t164 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0 l=0
X799 VPWR VGND.t202 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0 l=0
R0 VPWR VPWR 5445.48
R1 VPWR VPWR 3267.29
R2 VPWR VPWR 2450.47
R3 VPWR VPWR 2317.93
R4 VPWR VPWR 2181.15
R5 VPWR VPWR 2178.19
R6 VPWR VPWR 2178.19
R7 VPWR VPWR 2175.23
R8 VPWR VPWR 2007.42
R9 VPWR VPWR 1905.92
R10 VPWR VPWR 1698.59
R11 VPWR VPWR 1698.59
R12 VPWR VPWR 1633.64
R13 VPWR VPWR 1633.64
R14 VPWR VPWR 1633.64
R15 VPWR VPWR 1633.64
R16 VPWR.n3095 VPWR 1572.7
R17 VPWR VPWR 1544.17
R18 VPWR VPWR 1314.22
R19 VPWR.n3973 VPWR 1263.87
R20 VPWR VPWR 1238.69
R21 VPWR VPWR 1238.69
R22 VPWR VPWR 1238.69
R23 VPWR VPWR 1237.01
R24 VPWR VPWR 1235.34
R25 VPWR VPWR 1235.34
R26 VPWR VPWR 1235.34
R27 VPWR VPWR 1235.34
R28 VPWR VPWR 1233.66
R29 VPWR VPWR 1233.66
R30 VPWR VPWR 1233.66
R31 VPWR VPWR 1233.66
R32 VPWR VPWR 1233.66
R33 VPWR VPWR 1233.66
R34 VPWR VPWR 1233.66
R35 VPWR VPWR 1233.66
R36 VPWR VPWR 1233.66
R37 VPWR VPWR 1159.81
R38 VPWR.n2392 VPWR 1139.41
R39 VPWR.n2347 VPWR 1139.41
R40 VPWR.n2340 VPWR 1139.41
R41 VPWR.n2339 VPWR 1139.41
R42 VPWR.n2338 VPWR 1139.41
R43 VPWR VPWR 1089.1
R44 VPWR VPWR 1089.1
R45 VPWR VPWR 1089.1
R46 VPWR VPWR 1089.1
R47 VPWR VPWR 1089.1
R48 VPWR VPWR 1089.1
R49 VPWR VPWR 1089.1
R50 VPWR VPWR 1089.1
R51 VPWR VPWR 1080.92
R52 VPWR VPWR 1080.92
R53 VPWR VPWR 1080.92
R54 VPWR VPWR 1080.92
R55 VPWR VPWR 1080.92
R56 VPWR VPWR 1080.92
R57 VPWR VPWR 1080.92
R58 VPWR VPWR 1080.92
R59 VPWR VPWR 1080.92
R60 VPWR VPWR 1080.92
R61 VPWR VPWR 1080.92
R62 VPWR VPWR 1079.24
R63 VPWR VPWR 1079.24
R64 VPWR VPWR 1079.24
R65 VPWR VPWR 1077.56
R66 VPWR VPWR 1052.39
R67 VPWR VPWR.n3438 955.035
R68 VPWR VPWR.n3972 955.035
R69 VPWR.n5270 VPWR 955.035
R70 VPWR VPWR 929.86
R71 VPWR VPWR 929.86
R72 VPWR VPWR 929.86
R73 VPWR VPWR 929.86
R74 VPWR VPWR 929.86
R75 VPWR VPWR 929.86
R76 VPWR VPWR 929.86
R77 VPWR VPWR 928.181
R78 VPWR VPWR 926.503
R79 VPWR VPWR 926.503
R80 VPWR VPWR 926.503
R81 VPWR VPWR 926.503
R82 VPWR VPWR 926.503
R83 VPWR VPWR 926.503
R84 VPWR VPWR 926.503
R85 VPWR VPWR 926.503
R86 VPWR VPWR 926.503
R87 VPWR VPWR 926.503
R88 VPWR VPWR 926.503
R89 VPWR VPWR 926.503
R90 VPWR VPWR 926.503
R91 VPWR VPWR 926.503
R92 VPWR VPWR 926.503
R93 VPWR VPWR 926.503
R94 VPWR VPWR 924.823
R95 VPWR VPWR 924.823
R96 VPWR VPWR 924.823
R97 VPWR VPWR 924.823
R98 VPWR VPWR 924.823
R99 VPWR VPWR 924.823
R100 VPWR VPWR 924.823
R101 VPWR VPWR 924.823
R102 VPWR VPWR 850.972
R103 VPWR VPWR 850.972
R104 VPWR VPWR 816.822
R105 VPWR VPWR 775.442
R106 VPWR VPWR 773.764
R107 VPWR VPWR 773.764
R108 VPWR VPWR 772.086
R109 VPWR VPWR 772.086
R110 VPWR VPWR 772.086
R111 VPWR VPWR 772.086
R112 VPWR VPWR 772.086
R113 VPWR VPWR 772.086
R114 VPWR VPWR 772.086
R115 VPWR VPWR 772.086
R116 VPWR VPWR 772.086
R117 VPWR VPWR 772.086
R118 VPWR VPWR 772.086
R119 VPWR VPWR 772.086
R120 VPWR VPWR 772.086
R121 VPWR VPWR 770.407
R122 VPWR VPWR 770.407
R123 VPWR VPWR 770.407
R124 VPWR VPWR 770.407
R125 VPWR VPWR 770.407
R126 VPWR VPWR 770.407
R127 VPWR VPWR 770.407
R128 VPWR VPWR 768.729
R129 VPWR VPWR 768.729
R130 VPWR VPWR 768.729
R131 VPWR VPWR 767.049
R132 VPWR VPWR 693.198
R133 VPWR.n6194 VPWR 646.202
R134 VPWR.n6193 VPWR 646.202
R135 VPWR.n3094 VPWR 646.202
R136 VPWR.n3092 VPWR 646.202
R137 VPWR.n3091 VPWR 646.202
R138 VPWR.n1908 VPWR 646.202
R139 VPWR VPWR.n2026 646.202
R140 VPWR VPWR.n3029 646.202
R141 VPWR VPWR.n3295 646.202
R142 VPWR VPWR.n1219 646.202
R143 VPWR VPWR.n1266 646.202
R144 VPWR.n4362 VPWR 646.202
R145 VPWR.n4361 VPWR 646.202
R146 VPWR.n4358 VPWR 646.202
R147 VPWR VPWR.n4474 646.202
R148 VPWR.n5791 VPWR 646.202
R149 VPWR.n5788 VPWR 646.202
R150 VPWR VPWR.n158 646.202
R151 VPWR.n5404 VPWR 646.202
R152 VPWR VPWR 621.025
R153 VPWR VPWR 621.025
R154 VPWR VPWR 621.025
R155 VPWR VPWR 621.025
R156 VPWR VPWR 621.025
R157 VPWR VPWR 621.025
R158 VPWR VPWR 621.025
R159 VPWR VPWR 621.025
R160 VPWR VPWR 621.025
R161 VPWR VPWR 621.025
R162 VPWR VPWR 621.025
R163 VPWR VPWR 621.025
R164 VPWR VPWR 619.346
R165 VPWR VPWR 619.346
R166 VPWR VPWR 619.346
R167 VPWR VPWR 619.346
R168 VPWR VPWR 619.346
R169 VPWR VPWR 619.346
R170 VPWR VPWR 619.346
R171 VPWR VPWR 619.346
R172 VPWR VPWR 619.346
R173 VPWR VPWR 619.346
R174 VPWR VPWR 619.346
R175 VPWR VPWR 617.668
R176 VPWR VPWR 617.668
R177 VPWR VPWR 617.668
R178 VPWR VPWR 617.668
R179 VPWR VPWR 617.668
R180 VPWR VPWR 617.668
R181 VPWR VPWR 617.668
R182 VPWR VPWR 617.668
R183 VPWR VPWR 617.668
R184 VPWR VPWR 617.668
R185 VPWR VPWR 617.668
R186 VPWR VPWR 617.668
R187 VPWR VPWR 617.668
R188 VPWR VPWR 617.668
R189 VPWR VPWR 617.668
R190 VPWR VPWR 617.668
R191 VPWR VPWR 617.668
R192 VPWR VPWR 617.668
R193 VPWR VPWR 617.668
R194 VPWR VPWR 617.668
R195 VPWR VPWR 617.668
R196 VPWR VPWR 617.668
R197 VPWR VPWR 617.668
R198 VPWR VPWR 617.668
R199 VPWR VPWR 617.668
R200 VPWR VPWR 617.668
R201 VPWR VPWR 617.668
R202 VPWR VPWR 617.668
R203 VPWR VPWR 617.668
R204 VPWR VPWR 617.668
R205 VPWR VPWR 617.668
R206 VPWR VPWR 617.668
R207 VPWR VPWR 617.668
R208 VPWR VPWR 617.668
R209 VPWR VPWR 617.668
R210 VPWR VPWR 617.668
R211 VPWR VPWR 617.668
R212 VPWR VPWR 617.668
R213 VPWR VPWR 617.668
R214 VPWR VPWR 617.668
R215 VPWR VPWR 617.668
R216 VPWR VPWR 617.668
R217 VPWR VPWR 617.668
R218 VPWR VPWR 617.668
R219 VPWR VPWR 617.668
R220 VPWR VPWR 617.668
R221 VPWR VPWR 617.668
R222 VPWR VPWR 617.668
R223 VPWR VPWR 617.668
R224 VPWR VPWR 617.668
R225 VPWR VPWR 617.668
R226 VPWR VPWR 617.668
R227 VPWR VPWR 617.668
R228 VPWR VPWR 617.668
R229 VPWR VPWR 617.668
R230 VPWR VPWR 617.668
R231 VPWR VPWR 617.668
R232 VPWR VPWR 617.668
R233 VPWR VPWR 617.668
R234 VPWR VPWR 617.668
R235 VPWR VPWR 617.668
R236 VPWR VPWR 617.668
R237 VPWR VPWR 617.668
R238 VPWR VPWR 617.668
R239 VPWR VPWR 617.668
R240 VPWR VPWR 617.668
R241 VPWR VPWR 617.668
R242 VPWR VPWR 617.668
R243 VPWR VPWR 617.668
R244 VPWR VPWR 615.99
R245 VPWR VPWR 615.99
R246 VPWR VPWR 615.99
R247 VPWR VPWR 615.99
R248 VPWR VPWR 615.99
R249 VPWR VPWR 615.99
R250 VPWR VPWR 614.312
R251 VPWR VPWR 614.312
R252 VPWR VPWR 614.312
R253 VPWR VPWR 612.634
R254 VPWR VPWR.n1267 570.672
R255 VPWR VPWR 542.139
R256 VPWR VPWR 542.139
R257 VPWR VPWR.n4084 491.784
R258 VPWR.n4829 VPWR 491.784
R259 VPWR.n4828 VPWR 491.784
R260 VPWR.n4826 VPWR 491.784
R261 VPWR VPWR 466.608
R262 VPWR VPWR 466.608
R263 VPWR VPWR 466.608
R264 VPWR VPWR 466.608
R265 VPWR VPWR 464.93
R266 VPWR VPWR 464.93
R267 VPWR VPWR 464.93
R268 VPWR VPWR 464.93
R269 VPWR VPWR 463.252
R270 VPWR VPWR 463.252
R271 VPWR VPWR 463.252
R272 VPWR VPWR 463.252
R273 VPWR VPWR 463.252
R274 VPWR VPWR 463.252
R275 VPWR VPWR 463.252
R276 VPWR VPWR 463.252
R277 VPWR VPWR 463.252
R278 VPWR VPWR 463.252
R279 VPWR VPWR 463.252
R280 VPWR VPWR 463.252
R281 VPWR VPWR 463.252
R282 VPWR VPWR 463.252
R283 VPWR VPWR 463.252
R284 VPWR VPWR 463.252
R285 VPWR VPWR 463.252
R286 VPWR VPWR 463.252
R287 VPWR VPWR 463.252
R288 VPWR VPWR 463.252
R289 VPWR VPWR 463.252
R290 VPWR VPWR 463.252
R291 VPWR VPWR 463.252
R292 VPWR VPWR 463.252
R293 VPWR VPWR 463.252
R294 VPWR VPWR 463.252
R295 VPWR VPWR 463.252
R296 VPWR VPWR 463.252
R297 VPWR VPWR 463.252
R298 VPWR VPWR 463.252
R299 VPWR VPWR 463.252
R300 VPWR VPWR 463.252
R301 VPWR VPWR 463.252
R302 VPWR VPWR 463.252
R303 VPWR VPWR 463.252
R304 VPWR VPWR 463.252
R305 VPWR VPWR 463.252
R306 VPWR VPWR 463.252
R307 VPWR VPWR 463.252
R308 VPWR VPWR 463.252
R309 VPWR VPWR 463.252
R310 VPWR VPWR 463.252
R311 VPWR VPWR 463.252
R312 VPWR VPWR 463.252
R313 VPWR VPWR 463.252
R314 VPWR VPWR 463.252
R315 VPWR VPWR 463.252
R316 VPWR VPWR 463.252
R317 VPWR VPWR 463.252
R318 VPWR VPWR 463.252
R319 VPWR VPWR 463.252
R320 VPWR VPWR 463.252
R321 VPWR VPWR 463.252
R322 VPWR VPWR 463.252
R323 VPWR VPWR 463.252
R324 VPWR VPWR 463.252
R325 VPWR VPWR 463.252
R326 VPWR VPWR 461.572
R327 VPWR VPWR 461.572
R328 VPWR VPWR 461.572
R329 VPWR VPWR 461.572
R330 VPWR VPWR 461.572
R331 VPWR VPWR 461.572
R332 VPWR VPWR 461.572
R333 VPWR VPWR 461.572
R334 VPWR VPWR 461.572
R335 VPWR VPWR 461.572
R336 VPWR VPWR 459.894
R337 VPWR VPWR 459.894
R338 VPWR VPWR 459.894
R339 VPWR VPWR 459.894
R340 VPWR VPWR 459.894
R341 VPWR VPWR 459.894
R342 VPWR VPWR 459.894
R343 VPWR VPWR 459.894
R344 VPWR VPWR 458.216
R345 VPWR VPWR 458.216
R346 VPWR VPWR 384.365
R347 VPWR VPWR 384.365
R348 VPWR.n4360 VPWR 339.046
R349 VPWR.n4359 VPWR 339.046
R350 VPWR.n1485 VPWR 337.368
R351 VPWR VPWR 312.192
R352 VPWR VPWR 312.192
R353 VPWR VPWR 312.192
R354 VPWR VPWR 312.192
R355 VPWR VPWR 312.192
R356 VPWR VPWR 312.192
R357 VPWR VPWR 312.192
R358 VPWR VPWR 312.192
R359 VPWR VPWR 312.192
R360 VPWR VPWR 312.192
R361 VPWR VPWR 312.192
R362 VPWR VPWR 312.192
R363 VPWR VPWR 310.512
R364 VPWR VPWR 310.512
R365 VPWR VPWR 310.512
R366 VPWR VPWR 310.512
R367 VPWR VPWR 310.512
R368 VPWR VPWR 310.512
R369 VPWR VPWR 310.512
R370 VPWR VPWR 308.834
R371 VPWR VPWR 308.834
R372 VPWR VPWR 308.834
R373 VPWR VPWR 308.834
R374 VPWR VPWR 308.834
R375 VPWR VPWR 308.834
R376 VPWR VPWR 308.834
R377 VPWR VPWR 308.834
R378 VPWR VPWR 308.834
R379 VPWR VPWR 308.834
R380 VPWR VPWR 308.834
R381 VPWR VPWR 308.834
R382 VPWR VPWR 308.834
R383 VPWR VPWR 308.834
R384 VPWR VPWR 308.834
R385 VPWR VPWR 308.834
R386 VPWR VPWR 308.834
R387 VPWR VPWR 308.834
R388 VPWR VPWR 308.834
R389 VPWR VPWR 308.834
R390 VPWR VPWR 308.834
R391 VPWR VPWR 308.834
R392 VPWR VPWR 308.834
R393 VPWR VPWR 308.834
R394 VPWR VPWR 308.834
R395 VPWR VPWR 308.834
R396 VPWR VPWR 308.834
R397 VPWR VPWR 308.834
R398 VPWR VPWR 308.834
R399 VPWR VPWR 308.834
R400 VPWR VPWR 308.834
R401 VPWR VPWR 308.834
R402 VPWR VPWR.n5144 308.834
R403 VPWR VPWR 308.834
R404 VPWR VPWR 308.834
R405 VPWR VPWR 308.834
R406 VPWR VPWR 308.834
R407 VPWR VPWR 308.834
R408 VPWR VPWR 308.834
R409 VPWR VPWR 308.834
R410 VPWR VPWR 308.834
R411 VPWR VPWR 308.834
R412 VPWR VPWR 308.834
R413 VPWR VPWR 307.156
R414 VPWR VPWR 307.156
R415 VPWR VPWR 307.156
R416 VPWR VPWR 307.156
R417 VPWR VPWR 307.156
R418 VPWR VPWR 305.478
R419 VPWR VPWR 272.274
R420 VPWR VPWR 272.274
R421 VPWR VPWR 272.274
R422 VPWR VPWR 272.274
R423 VPWR VPWR 272.274
R424 VPWR VPWR 272.274
R425 VPWR VPWR 229.947
R426 VPWR VPWR 228.269
R427 VPWR.n2392 VPWR 221.964
R428 VPWR VPWR.n2347 221.964
R429 VPWR VPWR.n2340 221.964
R430 VPWR VPWR.n2339 221.964
R431 VPWR VPWR.n2338 221.964
R432 VPWR VPWR.n24 182.952
R433 VPWR.n3439 VPWR 182.952
R434 VPWR.n1292 VPWR 182.952
R435 VPWR.n4997 VPWR 182.952
R436 VPWR.n5145 VPWR 182.952
R437 VPWR.n5790 VPWR 182.952
R438 VPWR.n4827 VPWR 181.273
R439 VPWR VPWR.n59 179.595
R440 VPWR VPWR.n60 179.595
R441 VPWR.n3093 VPWR 179.595
R442 VPWR.n2027 VPWR 179.595
R443 VPWR.n3296 VPWR 179.595
R444 VPWR.n3857 VPWR 179.595
R445 VPWR VPWR.n5269 179.595
R446 VPWR.n5789 VPWR 179.595
R447 VPWR.n5924 VPWR 179.595
R448 VPWR.n5403 VPWR 179.595
R449 VPWR.n5596 VPWR.t276 178.661
R450 VPWR.n0 VPWR.t260 178.661
R451 VPWR.n0 VPWR.t288 178.661
R452 VPWR.n1623 VPWR.t81 178.661
R453 VPWR.n1623 VPWR.t98 178.661
R454 VPWR.n1622 VPWR.t55 178.661
R455 VPWR.n1525 VPWR.t88 178.661
R456 VPWR.n1525 VPWR.t108 178.661
R457 VPWR.n1703 VPWR.t121 178.661
R458 VPWR.n1703 VPWR.t146 178.661
R459 VPWR.n1845 VPWR.t131 178.661
R460 VPWR.n1845 VPWR.t163 178.661
R461 VPWR.n3157 VPWR.t279 178.661
R462 VPWR.n3157 VPWR.t304 178.661
R463 VPWR.n1338 VPWR.t262 178.661
R464 VPWR.n1338 VPWR.t287 178.661
R465 VPWR.n3483 VPWR.t318 178.661
R466 VPWR.n3483 VPWR.t339 178.661
R467 VPWR.n1142 VPWR.t327 178.661
R468 VPWR.n1142 VPWR.t351 178.661
R469 VPWR.n3813 VPWR.t379 178.661
R470 VPWR.n3813 VPWR.t263 178.661
R471 VPWR.n1003 VPWR.t369 178.661
R472 VPWR.n1003 VPWR.t247 178.661
R473 VPWR.n1002 VPWR.t305 178.661
R474 VPWR.n1002 VPWR.t231 178.661
R475 VPWR.n4154 VPWR.t278 178.661
R476 VPWR.n4154 VPWR.t303 178.661
R477 VPWR.n704 VPWR.t291 178.661
R478 VPWR.n704 VPWR.t317 178.661
R479 VPWR.n4402 VPWR.t336 178.661
R480 VPWR.n4402 VPWR.t368 178.661
R481 VPWR.n4522 VPWR.t326 178.661
R482 VPWR.n4522 VPWR.t350 178.661
R483 VPWR.n4521 VPWR.t179 178.661
R484 VPWR.n267 VPWR.t234 178.661
R485 VPWR.n267 VPWR.t261 178.661
R486 VPWR.n4947 VPWR.t246 178.661
R487 VPWR.n4947 VPWR.t277 178.661
R488 VPWR.n5337 VPWR.t290 178.661
R489 VPWR.n5337 VPWR.t316 178.661
R490 VPWR.n194 VPWR.t302 178.661
R491 VPWR.n194 VPWR.t325 178.661
R492 VPWR.n5866 VPWR.t352 178.661
R493 VPWR.n5866 VPWR.t233 178.661
R494 VPWR.n5695 VPWR.t335 178.661
R495 VPWR.n5695 VPWR.t224 178.661
R496 VPWR.n5596 VPWR.t245 178.661
R497 VPWR.n203 VPWR.t202 177.762
R498 VPWR.n5865 VPWR.t212 177.762
R499 VPWR.n3626 VPWR.n1254 169.4
R500 VPWR.n2262 VPWR.t62 166.282
R501 VPWR.n2402 VPWR.t73 166.282
R502 VPWR VPWR 159.452
R503 VPWR VPWR 159.452
R504 VPWR VPWR 157.774
R505 VPWR VPWR 157.774
R506 VPWR VPWR 157.774
R507 VPWR VPWR 157.774
R508 VPWR VPWR 157.774
R509 VPWR VPWR 157.774
R510 VPWR VPWR 157.774
R511 VPWR VPWR 157.774
R512 VPWR VPWR 157.774
R513 VPWR VPWR 157.774
R514 VPWR VPWR 156.095
R515 VPWR VPWR 156.095
R516 VPWR VPWR 156.095
R517 VPWR VPWR 156.095
R518 VPWR VPWR 156.095
R519 VPWR VPWR 156.095
R520 VPWR VPWR 156.095
R521 VPWR VPWR 156.095
R522 VPWR VPWR 156.095
R523 VPWR VPWR 156.095
R524 VPWR VPWR 156.095
R525 VPWR VPWR 156.095
R526 VPWR VPWR 156.095
R527 VPWR VPWR 156.095
R528 VPWR VPWR 156.095
R529 VPWR VPWR 156.095
R530 VPWR VPWR 156.095
R531 VPWR VPWR 156.095
R532 VPWR VPWR 156.095
R533 VPWR VPWR 156.095
R534 VPWR VPWR 156.095
R535 VPWR VPWR 156.095
R536 VPWR VPWR 156.095
R537 VPWR VPWR 156.095
R538 VPWR VPWR 156.095
R539 VPWR VPWR 156.095
R540 VPWR VPWR 156.095
R541 VPWR VPWR 156.095
R542 VPWR VPWR 154.417
R543 VPWR VPWR 154.417
R544 VPWR VPWR 154.417
R545 VPWR VPWR 154.417
R546 VPWR VPWR 154.417
R547 VPWR VPWR 154.417
R548 VPWR VPWR 154.417
R549 VPWR VPWR 154.417
R550 VPWR VPWR 154.417
R551 VPWR VPWR 154.417
R552 VPWR VPWR 154.417
R553 VPWR VPWR 154.417
R554 VPWR VPWR 154.417
R555 VPWR VPWR 154.417
R556 VPWR VPWR 154.417
R557 VPWR VPWR 154.417
R558 VPWR VPWR 154.417
R559 VPWR VPWR 154.417
R560 VPWR VPWR 154.417
R561 VPWR VPWR 154.417
R562 VPWR VPWR 154.417
R563 VPWR VPWR 154.417
R564 VPWR VPWR 154.417
R565 VPWR VPWR 154.417
R566 VPWR VPWR 154.417
R567 VPWR VPWR 154.417
R568 VPWR VPWR 154.417
R569 VPWR VPWR 154.417
R570 VPWR VPWR 154.417
R571 VPWR VPWR 154.417
R572 VPWR VPWR 154.417
R573 VPWR VPWR 154.417
R574 VPWR VPWR 154.417
R575 VPWR VPWR 154.417
R576 VPWR VPWR 154.417
R577 VPWR VPWR 154.417
R578 VPWR VPWR 154.417
R579 VPWR VPWR 154.417
R580 VPWR VPWR 154.417
R581 VPWR VPWR 154.417
R582 VPWR VPWR 154.417
R583 VPWR VPWR 154.417
R584 VPWR VPWR 154.417
R585 VPWR VPWR 154.417
R586 VPWR VPWR 154.417
R587 VPWR VPWR 154.417
R588 VPWR VPWR 154.417
R589 VPWR VPWR 154.417
R590 VPWR VPWR 154.417
R591 VPWR VPWR 154.417
R592 VPWR VPWR 154.417
R593 VPWR VPWR 154.417
R594 VPWR VPWR 154.417
R595 VPWR VPWR 154.417
R596 VPWR VPWR 154.417
R597 VPWR VPWR 154.417
R598 VPWR VPWR 154.417
R599 VPWR VPWR 154.417
R600 VPWR VPWR 154.417
R601 VPWR VPWR 154.417
R602 VPWR VPWR 154.417
R603 VPWR VPWR 154.417
R604 VPWR VPWR 154.417
R605 VPWR VPWR 154.417
R606 VPWR VPWR 154.417
R607 VPWR VPWR 154.417
R608 VPWR VPWR 154.417
R609 VPWR VPWR 154.417
R610 VPWR VPWR 154.417
R611 VPWR VPWR 154.417
R612 VPWR VPWR 154.417
R613 VPWR VPWR 154.417
R614 VPWR VPWR 154.417
R615 VPWR VPWR 154.417
R616 VPWR VPWR 154.417
R617 VPWR VPWR 154.417
R618 VPWR VPWR 154.417
R619 VPWR VPWR 154.417
R620 VPWR VPWR 154.417
R621 VPWR VPWR 154.417
R622 VPWR VPWR 154.417
R623 VPWR VPWR 154.417
R624 VPWR VPWR 154.417
R625 VPWR VPWR 154.417
R626 VPWR VPWR 154.417
R627 VPWR VPWR 154.417
R628 VPWR VPWR 154.417
R629 VPWR VPWR 154.417
R630 VPWR VPWR 154.417
R631 VPWR VPWR 154.417
R632 VPWR VPWR 154.417
R633 VPWR VPWR 154.417
R634 VPWR VPWR 154.417
R635 VPWR VPWR 154.417
R636 VPWR VPWR 154.417
R637 VPWR VPWR 154.417
R638 VPWR VPWR 154.417
R639 VPWR VPWR 154.417
R640 VPWR VPWR 152.739
R641 VPWR VPWR 152.739
R642 VPWR VPWR 152.739
R643 VPWR VPWR 152.739
R644 VPWR VPWR 152.739
R645 VPWR VPWR 152.739
R646 VPWR VPWR 152.739
R647 VPWR VPWR 152.739
R648 VPWR VPWR 152.739
R649 VPWR VPWR 152.739
R650 VPWR VPWR 152.739
R651 VPWR VPWR 152.739
R652 VPWR VPWR 151.06
R653 VPWR VPWR 151.06
R654 VPWR VPWR 151.06
R655 VPWR VPWR 151.06
R656 VPWR VPWR 151.06
R657 VPWR VPWR 151.06
R658 VPWR VPWR 151.06
R659 VPWR VPWR 151.06
R660 VPWR VPWR 151.06
R661 VPWR VPWR 151.06
R662 VPWR VPWR 151.06
R663 VPWR VPWR 151.06
R664 VPWR VPWR 151.06
R665 VPWR VPWR 151.06
R666 VPWR VPWR 151.06
R667 VPWR VPWR 151.06
R668 VPWR VPWR 151.06
R669 VPWR VPWR 151.06
R670 VPWR VPWR 151.06
R671 VPWR VPWR 151.06
R672 VPWR VPWR 151.06
R673 VPWR VPWR 151.06
R674 VPWR VPWR 151.06
R675 VPWR VPWR 151.06
R676 VPWR VPWR 151.06
R677 VPWR VPWR 151.06
R678 VPWR VPWR 151.06
R679 VPWR VPWR 151.06
R680 VPWR VPWR 149.382
R681 VPWR.n3824 VPWR.t382 147.173
R682 VPWR.n708 VPWR.t192 146.809
R683 VPWR.n4406 VPWR.t356 146.809
R684 VPWR.n2856 VPWR.t52 145.663
R685 VPWR.n2773 VPWR.t16 145.663
R686 VPWR.n2777 VPWR.t85 145.663
R687 VPWR.n1812 VPWR.t84 145.663
R688 VPWR.n1813 VPWR.t194 145.663
R689 VPWR.n3404 VPWR.t59 145.663
R690 VPWR.n3377 VPWR.t259 145.663
R691 VPWR.n3324 VPWR.t199 145.663
R692 VPWR.n3303 VPWR.t114 145.663
R693 VPWR.n1290 VPWR.t323 145.663
R694 VPWR.n3898 VPWR.t320 145.663
R695 VPWR.n5110 VPWR.t112 145.663
R696 VPWR.n224 VPWR.t319 145.663
R697 VPWR.n5971 VPWR.t104 144.105
R698 VPWR.n3 VPWR.t90 143.94
R699 VPWR.n3 VPWR.t374 143.94
R700 VPWR.n6305 VPWR.t123 143.94
R701 VPWR.n6305 VPWR.t10 143.94
R702 VPWR.n6213 VPWR.t141 143.94
R703 VPWR.n6213 VPWR.t268 143.94
R704 VPWR.n1528 VPWR.t103 143.94
R705 VPWR.n1528 VPWR.t385 143.94
R706 VPWR.n3016 VPWR.t11 143.94
R707 VPWR.n3016 VPWR.t136 143.94
R708 VPWR.n1848 VPWR.t241 143.94
R709 VPWR.n1848 VPWR.t137 143.94
R710 VPWR.n1411 VPWR.t180 143.94
R711 VPWR.n1337 VPWR.t383 143.94
R712 VPWR.n1337 VPWR.t169 143.94
R713 VPWR.n3160 VPWR.t284 143.94
R714 VPWR.n3261 VPWR.t28 143.94
R715 VPWR.n3261 VPWR.t283 143.94
R716 VPWR.n1495 VPWR.t83 143.94
R717 VPWR.n1495 VPWR.t357 143.94
R718 VPWR.n1163 VPWR.t182 143.94
R719 VPWR.n1163 VPWR.t76 143.94
R720 VPWR.n1211 VPWR.t165 143.94
R721 VPWR.n3805 VPWR.t344 143.94
R722 VPWR.n3816 VPWR.t321 143.94
R723 VPWR.n3816 VPWR.t331 143.94
R724 VPWR.n1068 VPWR.t18 143.94
R725 VPWR.n1068 VPWR.t139 143.94
R726 VPWR.n820 VPWR.t164 143.94
R727 VPWR.n268 VPWR.t365 143.94
R728 VPWR.n268 VPWR.t142 143.94
R729 VPWR.n275 VPWR.t149 143.94
R730 VPWR.n503 VPWR.t370 143.94
R731 VPWR.n193 VPWR.t264 143.94
R732 VPWR.n193 VPWR.t161 143.94
R733 VPWR.n5696 VPWR.t282 143.94
R734 VPWR.n5696 VPWR.t390 143.94
R735 VPWR.n2772 VPWR.t186 143.694
R736 VPWR.n2775 VPWR.t157 143.694
R737 VPWR.n1966 VPWR.t345 143.694
R738 VPWR.n3403 VPWR.t207 143.694
R739 VPWR.n3322 VPWR.t366 143.694
R740 VPWR.n3302 VPWR.t27 143.694
R741 VPWR.n1279 VPWR.t89 143.694
R742 VPWR.n3897 VPWR.t359 143.694
R743 VPWR.n5111 VPWR.t8 143.694
R744 VPWR.n566 VPWR.t209 143.694
R745 VPWR.n1119 VPWR.t387 143.078
R746 VPWR.n4945 VPWR.t120 142.835
R747 VPWR.n1522 VPWR.t156 142.519
R748 VPWR.n1486 VPWR.t338 142.519
R749 VPWR.n5331 VPWR.t376 142.519
R750 VPWR.n191 VPWR.t306 142.519
R751 VPWR.n6197 VPWR.t130 141.607
R752 VPWR.n1764 VPWR.t185 141.607
R753 VPWR.n369 VPWR.t67 141.607
R754 VPWR.n5859 VPWR.t69 141.607
R755 VPWR.n717 VPWR.t220 141.058
R756 VPWR.n4415 VPWR.t0 141.058
R757 VPWR.n4692 VPWR.t125 141.058
R758 VPWR.n499 VPWR.t188 141.058
R759 VPWR.n4584 VPWR.t196 141.008
R760 VPWR.n5592 VPWR.t176 141.008
R761 VPWR.n4473 VPWR.t307 141.008
R762 VPWR.n501 VPWR.t162 141.008
R763 VPWR.n2646 VPWR.t78 140.714
R764 VPWR.n3397 VPWR.t58 140.714
R765 VPWR.n3171 VPWR.t35 140.714
R766 VPWR.n1144 VPWR.t166 140.714
R767 VPWR.n3703 VPWR.t214 140.714
R768 VPWR.n4031 VPWR.t105 140.714
R769 VPWR.n4510 VPWR.t173 140.714
R770 VPWR.n4594 VPWR.t77 140.714
R771 VPWR.n4941 VPWR.t22 140.714
R772 VPWR.n371 VPWR.t94 140.714
R773 VPWR.n76 VPWR.t227 140.364
R774 VPWR.n1699 VPWR.t30 140.364
R775 VPWR.n1064 VPWR.t363 140.364
R776 VPWR.n875 VPWR.t203 140.364
R777 VPWR.n4244 VPWR.t13 140.364
R778 VPWR.n4144 VPWR.t293 140.364
R779 VPWR.n5222 VPWR.t70 140.364
R780 VPWR.n5052 VPWR.t48 140.364
R781 VPWR.n4985 VPWR.t144 140.364
R782 VPWR.n5214 VPWR.t372 140.364
R783 VPWR.n494 VPWR.t367 140.364
R784 VPWR.n5525 VPWR.t175 140.364
R785 VPWR.n5482 VPWR.t80 140.364
R786 VPWR.n155 VPWR.t388 140.364
R787 VPWR.n6053 VPWR.t140 140.364
R788 VPWR.n5459 VPWR.t86 140.364
R789 VPWR.n5384 VPWR.t200 140.364
R790 VPWR.n5550 VPWR.t117 140.364
R791 VPWR.n51 VPWR.t354 135.263
R792 VPWR.n6236 VPWR.t61 134.964
R793 VPWR.n6121 VPWR.t322 134.964
R794 VPWR.n6098 VPWR.t97 134.964
R795 VPWR.n6131 VPWR.t253 134.964
R796 VPWR.n86 VPWR.t191 134.964
R797 VPWR.n6144 VPWR.t295 134.964
R798 VPWR.n6152 VPWR.t119 134.964
R799 VPWR.n6162 VPWR.t330 134.964
R800 VPWR.n2248 VPWR.t17 134.964
R801 VPWR.n2069 VPWR.t333 134.964
R802 VPWR.n2073 VPWR.t362 134.964
R803 VPWR.n2155 VPWR.t29 134.964
R804 VPWR.n2133 VPWR.t5 134.964
R805 VPWR.n2121 VPWR.t347 134.964
R806 VPWR.n2081 VPWR.t314 134.964
R807 VPWR.n2341 VPWR.t299 134.964
R808 VPWR.n2539 VPWR.t243 134.964
R809 VPWR.n2527 VPWR.t313 134.964
R810 VPWR.n2398 VPWR.t215 134.964
R811 VPWR.n2394 VPWR.t242 134.964
R812 VPWR.n2448 VPWR.t206 134.964
R813 VPWR.n1620 VPWR.t250 134.964
R814 VPWR.n1619 VPWR.t116 134.964
R815 VPWR.n1616 VPWR.t248 134.964
R816 VPWR.n1607 VPWR.t138 134.964
R817 VPWR.n1573 VPWR.t79 134.964
R818 VPWR.n2647 VPWR.t211 134.964
R819 VPWR.n2645 VPWR.t266 134.964
R820 VPWR.n2722 VPWR.t189 134.964
R821 VPWR.n2769 VPWR.t4 134.964
R822 VPWR.n1721 VPWR.t381 134.964
R823 VPWR.n1734 VPWR.t64 134.964
R824 VPWR.n1689 VPWR.t25 134.964
R825 VPWR.n1767 VPWR.t92 134.964
R826 VPWR.n2983 VPWR.t152 134.964
R827 VPWR.n2963 VPWR.t155 134.964
R828 VPWR.n1771 VPWR.t329 134.964
R829 VPWR.n1772 VPWR.t115 134.964
R830 VPWR.n2942 VPWR.t298 134.964
R831 VPWR.n1971 VPWR.t153 134.964
R832 VPWR.n1880 VPWR.t272 134.964
R833 VPWR.n1932 VPWR.t346 134.964
R834 VPWR.n3421 VPWR.t198 134.964
R835 VPWR.n1333 VPWR.t230 134.964
R836 VPWR.n1365 VPWR.t324 134.964
R837 VPWR.n1327 VPWR.t274 134.964
R838 VPWR.n1489 VPWR.t223 134.964
R839 VPWR.n3169 VPWR.t309 134.964
R840 VPWR.n3190 VPWR.t45 134.964
R841 VPWR.n3273 VPWR.t100 134.964
R842 VPWR.n1276 VPWR.t310 134.964
R843 VPWR.n3481 VPWR.t342 134.964
R844 VPWR.n3476 VPWR.t122 134.964
R845 VPWR.n3740 VPWR.t239 134.964
R846 VPWR.n1147 VPWR.t50 134.964
R847 VPWR.n1258 VPWR.t285 134.964
R848 VPWR.n3612 VPWR.t183 134.964
R849 VPWR.n1222 VPWR.t65 134.964
R850 VPWR.n1226 VPWR.t222 134.964
R851 VPWR.n1215 VPWR.t193 134.964
R852 VPWR.n1217 VPWR.t113 134.964
R853 VPWR.n3885 VPWR.t12 134.964
R854 VPWR.n999 VPWR.t378 134.964
R855 VPWR.n996 VPWR.t66 134.964
R856 VPWR.n990 VPWR.t36 134.964
R857 VPWR.n4038 VPWR.t364 134.964
R858 VPWR.n4036 VPWR.t129 134.964
R859 VPWR.n4082 VPWR.t386 134.964
R860 VPWR.n3930 VPWR.t47 134.964
R861 VPWR.n3928 VPWR.t334 134.964
R862 VPWR.n3923 VPWR.t358 134.964
R863 VPWR.n3905 VPWR.t15 134.964
R864 VPWR.n4161 VPWR.t39 134.964
R865 VPWR.n4175 VPWR.t249 134.964
R866 VPWR.n4189 VPWR.t341 134.964
R867 VPWR.n738 VPWR.t221 134.964
R868 VPWR.n943 VPWR.t235 134.964
R869 VPWR.n916 VPWR.t124 134.964
R870 VPWR.n816 VPWR.t99 134.964
R871 VPWR.n860 VPWR.t297 134.964
R872 VPWR.n4258 VPWR.t42 134.964
R873 VPWR.n4269 VPWR.t225 134.964
R874 VPWR.n4285 VPWR.t41 134.964
R875 VPWR.n761 VPWR.t328 134.964
R876 VPWR.n758 VPWR.t26 134.964
R877 VPWR.n4333 VPWR.t217 134.964
R878 VPWR.n4845 VPWR.t252 134.964
R879 VPWR.n4856 VPWR.t49 134.964
R880 VPWR.n4868 VPWR.t251 134.964
R881 VPWR.n4436 VPWR.t1 134.964
R882 VPWR.n4533 VPWR.t57 134.964
R883 VPWR.n4551 VPWR.t197 134.964
R884 VPWR.n4818 VPWR.t315 134.964
R885 VPWR.n4589 VPWR.t232 134.964
R886 VPWR.n4757 VPWR.t300 134.964
R887 VPWR.n4744 VPWR.t126 134.964
R888 VPWR.n4729 VPWR.t93 134.964
R889 VPWR.n4593 VPWR.t208 134.964
R890 VPWR.n4467 VPWR.t63 134.964
R891 VPWR.n311 VPWR.t380 134.964
R892 VPWR.n4961 VPWR.t143 134.964
R893 VPWR.n5122 VPWR.t74 134.964
R894 VPWR.n5105 VPWR.t371 134.964
R895 VPWR.n5097 VPWR.t23 134.964
R896 VPWR.n5063 VPWR.t87 134.964
R897 VPWR.n648 VPWR.t340 134.964
R898 VPWR.n5174 VPWR.t391 134.964
R899 VPWR.n5207 VPWR.t177 134.964
R900 VPWR.n5321 VPWR.t311 134.964
R901 VPWR.n498 VPWR.t265 134.964
R902 VPWR.n611 VPWR.t256 134.964
R903 VPWR.n457 VPWR.t195 134.964
R904 VPWR.n353 VPWR.t53 134.964
R905 VPWR.n354 VPWR.t257 134.964
R906 VPWR.n418 VPWR.t54 134.964
R907 VPWR.n409 VPWR.t7 134.964
R908 VPWR.n364 VPWR.t37 134.964
R909 VPWR.n374 VPWR.t229 134.964
R910 VPWR.n5864 VPWR.t38 134.964
R911 VPWR.n5508 VPWR.t389 134.964
R912 VPWR.n5993 VPWR.t267 134.964
R913 VPWR.n6005 VPWR.t213 134.964
R914 VPWR.n5621 VPWR.t296 134.964
R915 VPWR.n46 VPWR.t132 131.399
R916 VPWR.n161 VPWR.t219 128.713
R917 VPWR.n45 VPWR.t33 128.576
R918 VPWR.n184 VPWR.t216 127.45
R919 VPWR.n24 VPWR 125.883
R920 VPWR.n59 VPWR 125.883
R921 VPWR.n60 VPWR 125.883
R922 VPWR.n6196 VPWR 125.883
R923 VPWR VPWR.n6195 125.883
R924 VPWR VPWR.n6194 125.883
R925 VPWR VPWR.n6193 125.883
R926 VPWR.n3095 VPWR 125.883
R927 VPWR VPWR.n3094 125.883
R928 VPWR VPWR.n3093 125.883
R929 VPWR VPWR.n3092 125.883
R930 VPWR VPWR.n3091 125.883
R931 VPWR.n1908 VPWR 125.883
R932 VPWR.n2026 VPWR 125.883
R933 VPWR.n2027 VPWR 125.883
R934 VPWR.n3029 VPWR 125.883
R935 VPWR.n3030 VPWR 125.883
R936 VPWR.n3295 VPWR 125.883
R937 VPWR.n3296 VPWR 125.883
R938 VPWR VPWR.n1485 125.883
R939 VPWR.n3438 VPWR 125.883
R940 VPWR.n3439 VPWR 125.883
R941 VPWR.n1219 VPWR 125.883
R942 VPWR.n1220 VPWR 125.883
R943 VPWR.n1266 VPWR 125.883
R944 VPWR.n1267 VPWR 125.883
R945 VPWR.n1292 VPWR 125.883
R946 VPWR.n3857 VPWR 125.883
R947 VPWR.n3972 VPWR 125.883
R948 VPWR.n3973 VPWR 125.883
R949 VPWR.n4084 VPWR 125.883
R950 VPWR.n4085 VPWR 125.883
R951 VPWR.n4362 VPWR 125.883
R952 VPWR VPWR 125.883
R953 VPWR VPWR.n4361 125.883
R954 VPWR VPWR.n4360 125.883
R955 VPWR VPWR.n4359 125.883
R956 VPWR VPWR.n4358 125.883
R957 VPWR.n4474 VPWR 125.883
R958 VPWR.n4829 VPWR 125.883
R959 VPWR VPWR.n4828 125.883
R960 VPWR VPWR.n4827 125.883
R961 VPWR VPWR.n4826 125.883
R962 VPWR.n4997 VPWR 125.883
R963 VPWR.n5144 VPWR 125.883
R964 VPWR.n5145 VPWR 125.883
R965 VPWR.n5269 VPWR 125.883
R966 VPWR.n5270 VPWR 125.883
R967 VPWR.n5791 VPWR 125.883
R968 VPWR VPWR.n5790 125.883
R969 VPWR VPWR.n5789 125.883
R970 VPWR VPWR.n5788 125.883
R971 VPWR VPWR.n5787 125.883
R972 VPWR.n5924 VPWR 125.883
R973 VPWR VPWR.n158 125.883
R974 VPWR.n5388 VPWR 125.883
R975 VPWR.n5404 VPWR 125.883
R976 VPWR VPWR.n5403 125.883
R977 VPWR VPWR 124.206
R978 VPWR.n6229 VPWR.n60 120.481
R979 VPWR.n6194 VPWR.n74 120.481
R980 VPWR.n6195 VPWR.n73 120.481
R981 VPWR.n2338 VPWR.n2337 120.481
R982 VPWR.n2339 VPWR.n2068 120.481
R983 VPWR.n2593 VPWR.n2340 120.481
R984 VPWR.n2536 VPWR.n2347 120.481
R985 VPWR.n3091 VPWR.n3090 120.481
R986 VPWR.n3029 VPWR.n3028 120.481
R987 VPWR.n3438 VPWR.n3437 120.481
R988 VPWR.n3588 VPWR.n1267 120.481
R989 VPWR.n3974 VPWR.n3973 120.481
R990 VPWR.n3858 VPWR.n3857 120.481
R991 VPWR.n4361 VPWR.n750 120.481
R992 VPWR.n4360 VPWR.n751 120.481
R993 VPWR.n4363 VPWR.n4362 120.481
R994 VPWR.n4827 VPWR.n4476 120.481
R995 VPWR.n5144 VPWR.n5143 120.481
R996 VPWR.n5271 VPWR.n5270 120.481
R997 VPWR.n5788 VPWR.n227 120.481
R998 VPWR.n5789 VPWR.n226 120.481
R999 VPWR.n2439 VPWR.n2392 120.481
R1000 VPWR.n2026 VPWR.n2025 120.481
R1001 VPWR.n4359 VPWR.n752 120.481
R1002 VPWR.n4474 VPWR.n4447 120.481
R1003 VPWR.n5505 VPWR.n5404 120.481
R1004 VPWR.n6198 VPWR.n6196 119.094
R1005 VPWR.n3031 VPWR.n3030 119.094
R1006 VPWR.n3701 VPWR.n1220 119.094
R1007 VPWR.n5787 VPWR.n5786 119.094
R1008 VPWR.n4086 VPWR.n4085 119.094
R1009 VPWR.n4832 VPWR.n4829 118.513
R1010 VPWR.n5792 VPWR.n5791 118.484
R1011 VPWR.n1266 VPWR.n1265 118.457
R1012 VPWR.n5146 VPWR.n5145 118.457
R1013 VPWR.n3440 VPWR.n3439 118.456
R1014 VPWR.n1293 VPWR.n1292 118.456
R1015 VPWR.n2028 VPWR.n2027 117.912
R1016 VPWR.n5790 VPWR.n225 117.912
R1017 VPWR.n4998 VPWR.n4997 117.912
R1018 VPWR.n3340 VPWR.n1485 117.858
R1019 VPWR.n59 VPWR.n58 117.728
R1020 VPWR.n6290 VPWR.n24 116.73
R1021 VPWR.n3092 VPWR.n1572 116.73
R1022 VPWR.n3093 VPWR.n1571 116.73
R1023 VPWR.n3096 VPWR.n3095 116.73
R1024 VPWR.n1909 VPWR.n1908 116.73
R1025 VPWR.n3297 VPWR.n3296 116.73
R1026 VPWR.n3295 VPWR.n3294 116.73
R1027 VPWR.n1219 VPWR.n1190 116.73
R1028 VPWR.n3972 VPWR.n3971 116.73
R1029 VPWR.n4084 VPWR.n4083 116.73
R1030 VPWR.n4358 VPWR.n4357 116.73
R1031 VPWR.n4826 VPWR.n4825 116.73
R1032 VPWR.n4828 VPWR.n4475 116.73
R1033 VPWR.n5269 VPWR.n5268 116.73
R1034 VPWR.n6002 VPWR.n158 116.73
R1035 VPWR.n5403 VPWR.n5402 116.73
R1036 VPWR.n5388 VPWR.n5387 116.73
R1037 VPWR.n5933 VPWR.n5924 116.73
R1038 VPWR.n3094 VPWR.n1570 116.728
R1039 VPWR.n14 VPWR.t111 107.793
R1040 VPWR.n2489 VPWR.t273 107.793
R1041 VPWR.n2816 VPWR.t102 107.793
R1042 VPWR.n164 VPWR.t96 107.793
R1043 VPWR.n5930 VPWR.t226 107.793
R1044 VPWR.n6027 VPWR.t158 99.4427
R1045 VPWR.n5734 VPWR.t159 99.4427
R1046 VPWR.n2905 VPWR.t190 99.0895
R1047 VPWR.n4659 VPWR.t355 99.0895
R1048 VPWR.n4953 VPWR.t373 99.0895
R1049 VPWR.n490 VPWR.t348 99.0895
R1050 VPWR.n1820 VPWR.t361 97.5
R1051 VPWR.n1408 VPWR.t337 97.5
R1052 VPWR.n1817 VPWR.t205 96.1586
R1053 VPWR.n1410 VPWR.t31 96.1586
R1054 VPWR.n3161 VPWR.t3 96.1586
R1055 VPWR.n1212 VPWR.t135 96.1586
R1056 VPWR.n1270 VPWR.t109 95.5078
R1057 VPWR.n3601 VPWR.t82 95.5078
R1058 VPWR.n3808 VPWR.t294 95.5078
R1059 VPWR.n3989 VPWR.t19 95.5078
R1060 VPWR.n1128 VPWR.t40 95.5078
R1061 VPWR.n819 VPWR.t271 95.5078
R1062 VPWR.n4830 VPWR.t2 95.5078
R1063 VPWR.n4588 VPWR.t167 95.5078
R1064 VPWR.n276 VPWR.t21 95.5078
R1065 VPWR.n500 VPWR.t353 95.5078
R1066 VPWR.n89 VPWR.t270 95.5071
R1067 VPWR.n62 VPWR.t72 95.5071
R1068 VPWR.n1413 VPWR.t301 95.5071
R1069 VPWR.n709 VPWR.t150 95.5071
R1070 VPWR.n4407 VPWR.t292 95.5071
R1071 VPWR.n4583 VPWR.t286 95.5071
R1072 VPWR.n4655 VPWR.t174 95.5071
R1073 VPWR.n186 VPWR.t118 95.5071
R1074 VPWR.n5873 VPWR.t237 95.5071
R1075 VPWR.n5406 VPWR.t46 95.5071
R1076 VPWR.n5531 VPWR.t68 95.5071
R1077 VPWR.n5634 VPWR.t254 95.5071
R1078 VPWR.n2665 VPWR.t280 95.1199
R1079 VPWR.n5102 VPWR.t148 95.034
R1080 VPWR.n3807 VPWR.t360 94.8107
R1081 VPWR.n2997 VPWR.t343 94.3255
R1082 VPWR.n5100 VPWR.t171 94.1962
R1083 VPWR.n3391 VPWR.t275 93.6194
R1084 VPWR.n1254 VPWR.t134 93.6194
R1085 VPWR.n1124 VPWR.t14 93.6187
R1086 VPWR.n2652 VPWR.t168 93.2069
R1087 VPWR.n6171 VPWR.t107 91.34
R1088 VPWR.n92 VPWR.t60 91.34
R1089 VPWR.n6256 VPWR.t147 91.34
R1090 VPWR.n3253 VPWR.t44 91.34
R1091 VPWR.n1176 VPWR.t181 91.34
R1092 VPWR.n3473 VPWR.t133 91.34
R1093 VPWR.n3661 VPWR.t110 91.34
R1094 VPWR.n922 VPWR.t218 91.34
R1095 VPWR.n259 VPWR.t32 91.34
R1096 VPWR.n389 VPWR.t332 91.34
R1097 VPWR.n5327 VPWR.t312 91.34
R1098 VPWR.n595 VPWR.t228 91.34
R1099 VPWR.n5605 VPWR.t349 91.34
R1100 VPWR.n22 VPWR.t24 91.34
R1101 VPWR.n6203 VPWR.t269 91.34
R1102 VPWR.n2431 VPWR.t258 91.34
R1103 VPWR.n2274 VPWR.t255 91.34
R1104 VPWR.n1540 VPWR.t384 91.34
R1105 VPWR.n1860 VPWR.t154 91.34
R1106 VPWR.n3006 VPWR.t151 91.34
R1107 VPWR.n1709 VPWR.t187 91.34
R1108 VPWR.n3253 VPWR.t308 91.34
R1109 VPWR.n1268 VPWR.t204 91.34
R1110 VPWR.n3967 VPWR.t51 91.34
R1111 VPWR.n4021 VPWR.t170 91.34
R1112 VPWR.n4042 VPWR.t201 91.34
R1113 VPWR.n4142 VPWR.t34 91.34
R1114 VPWR.n5087 VPWR.t71 91.34
R1115 VPWR.n5216 VPWR.t91 91.34
R1116 VPWR.n5180 VPWR.t75 91.34
R1117 VPWR.n5344 VPWR.t106 91.34
R1118 VPWR.n5714 VPWR.t20 91.34
R1119 VPWR.n2765 VPWR.t95 91.2541
R1120 VPWR.n1552 VPWR.t127 91.2541
R1121 VPWR.n1974 VPWR.t375 91.2541
R1122 VPWR.n3358 VPWR.t244 91.2541
R1123 VPWR.n4241 VPWR.t236 91.2541
R1124 VPWR.n5046 VPWR.t145 91.2541
R1125 VPWR.n5894 VPWR.t56 91.2541
R1126 VPWR.n6085 VPWR.t281 91.2541
R1127 VPWR.n874 VPWR.t178 91.2541
R1128 VPWR.n4299 VPWR.t43 91.2541
R1129 VPWR.n5220 VPWR.t172 91.2541
R1130 VPWR.n4980 VPWR.t9 91.2541
R1131 VPWR.n578 VPWR.t210 91.2541
R1132 VPWR.n1251 VPWR.t184 90.7452
R1133 VPWR.n2636 VPWR.t128 88.005
R1134 VPWR.n4797 VPWR.t101 88.005
R1135 VPWR.n5887 VPWR.t238 86.1982
R1136 VPWR.n5711 VPWR.t160 86.1982
R1137 VPWR.n172 VPWR.n164 85.812
R1138 VPWR.n1858 VPWR.t240 85.8057
R1139 VPWR.n23 VPWR.n18 80.8005
R1140 VPWR.n167 VPWR.n166 80.6774
R1141 VPWR.n6299 VPWR.n17 76.0005
R1142 VPWR.n16 VPWR.n15 76.0005
R1143 VPWR.n2257 VPWR.n2256 76.0005
R1144 VPWR.n2581 VPWR.n2580 76.0005
R1145 VPWR.n2491 VPWR.n2490 76.0005
R1146 VPWR.n2502 VPWR.n2501 76.0005
R1147 VPWR.n2506 VPWR.n2505 76.0005
R1148 VPWR.n2828 VPWR.n2827 76.0005
R1149 VPWR.n2818 VPWR.n2817 76.0005
R1150 VPWR.n2824 VPWR.n2823 76.0005
R1151 VPWR.n214 VPWR.n213 76.0005
R1152 VPWR.n5932 VPWR.n5931 76.0005
R1153 VPWR.n5962 VPWR.n5961 76.0005
R1154 VPWR.n5967 VPWR.n5966 76.0005
R1155 VPWR VPWR 75.5305
R1156 VPWR VPWR 75.5305
R1157 VPWR.n6193 VPWR.n6192 60.2416
R1158 VPWR.n2255 VPWR.t6 50.5057
R1159 VPWR.n2579 VPWR.t377 50.5057
R1160 VPWR.n212 VPWR.t289 50.5057
R1161 VPWR.n45 VPWR.n41 48.8751
R1162 VPWR.n3656 VPWR.n1233 35.1785
R1163 VPWR.n3830 VPWR.n3807 35.1785
R1164 VPWR.n6219 VPWR.n66 34.6358
R1165 VPWR.n1651 VPWR.n1612 34.6358
R1166 VPWR.n1652 VPWR.n1651 34.6358
R1167 VPWR.n2971 VPWR.n2970 34.6358
R1168 VPWR.n1344 VPWR.n1343 34.6358
R1169 VPWR.n1344 VPWR.n1335 34.6358
R1170 VPWR.n3494 VPWR.n3493 34.6358
R1171 VPWR.n3494 VPWR.n3478 34.6358
R1172 VPWR.n1017 VPWR.n1016 34.6358
R1173 VPWR.n4279 VPWR.n4278 34.6358
R1174 VPWR.n4719 VPWR.n4718 34.6358
R1175 VPWR.n424 VPWR.n357 34.6358
R1176 VPWR.n420 VPWR.n357 34.6358
R1177 VPWR.n5489 VPWR.n5408 34.6358
R1178 VPWR.n5728 VPWR.n5727 34.6358
R1179 VPWR.n2558 VPWR.n2557 34.6358
R1180 VPWR.n1646 VPWR.n1645 34.6358
R1181 VPWR.n1647 VPWR.n1646 34.6358
R1182 VPWR.n1653 VPWR.n1652 34.6358
R1183 VPWR.n2892 VPWR.n2891 34.6358
R1184 VPWR.n1727 VPWR.n1695 34.6358
R1185 VPWR.n3267 VPWR.n3233 34.6358
R1186 VPWR.n3260 VPWR.n3236 34.6358
R1187 VPWR.n3729 VPWR.n3728 34.6358
R1188 VPWR.n3734 VPWR.n1209 34.6358
R1189 VPWR.n3670 VPWR.n1229 34.6358
R1190 VPWR.n3666 VPWR.n3665 34.6358
R1191 VPWR.n4050 VPWR.n4049 34.6358
R1192 VPWR.n3948 VPWR.n3926 34.6358
R1193 VPWR.n888 VPWR.n887 34.6358
R1194 VPWR.n4544 VPWR.n4519 34.6358
R1195 VPWR.n5248 VPWR.n5247 34.6358
R1196 VPWR.n203 VPWR.n202 34.6358
R1197 VPWR.n5490 VPWR.n5489 34.6358
R1198 VPWR.n5480 VPWR.n5479 34.6358
R1199 VPWR.n5989 VPWR.n5988 34.6358
R1200 VPWR.n6034 VPWR.n6033 34.6358
R1201 VPWR.n6051 VPWR.n6050 34.6358
R1202 VPWR.n5727 VPWR.n5690 34.6358
R1203 VPWR.n5546 VPWR.n5545 34.6358
R1204 VPWR.n5555 VPWR.n5554 33.1299
R1205 VPWR.n164 VPWR.n163 32.4617
R1206 VPWR.n5364 VPWR.n5363 32.0005
R1207 VPWR.n15 VPWR.n14 30.4944
R1208 VPWR.n2490 VPWR.n2489 30.4944
R1209 VPWR.n2817 VPWR.n2816 30.4944
R1210 VPWR.n5931 VPWR.n5930 30.4944
R1211 VPWR.n1030 VPWR.n1029 30.1181
R1212 VPWR.n6020 VPWR.n157 30.1181
R1213 VPWR.n6058 VPWR.n6057 30.1181
R1214 VPWR.n5464 VPWR.n5463 30.1181
R1215 VPWR.n6196 VPWR 28.5341
R1216 VPWR.n3030 VPWR 28.5341
R1217 VPWR VPWR.n1220 28.5341
R1218 VPWR.n4085 VPWR 28.5341
R1219 VPWR.n5787 VPWR 28.5341
R1220 VPWR VPWR.n5388 28.5341
R1221 VPWR.n590 VPWR.n589 28.2358
R1222 VPWR.n1653 VPWR 27.8593
R1223 VPWR.n6253 VPWR.n41 27.6743
R1224 VPWR.n6290 VPWR.n25 27.2033
R1225 VPWR.n3657 VPWR.n3656 27.2033
R1226 VPWR.n3830 VPWR.n3829 27.2033
R1227 VPWR.n4691 VPWR.n4654 27.2033
R1228 VPWR.n3164 VPWR.n3154 26.3534
R1229 VPWR.n4795 VPWR 26.3398
R1230 VPWR.n718 VPWR.n717 25.8527
R1231 VPWR.n4416 VPWR.n4415 25.8527
R1232 VPWR.n4692 VPWR.n4691 25.8527
R1233 VPWR.n549 VPWR.n499 25.8527
R1234 VPWR.n2129 VPWR.n2128 25.224
R1235 VPWR.n4015 VPWR.n4014 25.224
R1236 VPWR.n4182 VPWR.n4150 25.224
R1237 VPWR.n4959 VPWR.n4943 25.224
R1238 VPWR.n4049 VPWR.n4048 25.1912
R1239 VPWR.n3971 VPWR.n3970 25.1912
R1240 VPWR.n3906 VPWR.n3903 25.1912
R1241 VPWR.n3971 VPWR.n1123 25.1912
R1242 VPWR.n4736 VPWR.n4735 25.1912
R1243 VPWR.n6006 VPWR.n6002 25.1912
R1244 VPWR.n6122 VPWR.n6118 25.1912
R1245 VPWR.n6113 VPWR.n6112 25.1912
R1246 VPWR.n6165 VPWR.n82 25.1912
R1247 VPWR.n6205 VPWR.n6204 25.1912
R1248 VPWR.n2283 VPWR.n2282 25.1912
R1249 VPWR.n2207 VPWR.n2206 25.1912
R1250 VPWR.n2167 VPWR.n2166 25.1912
R1251 VPWR.n2122 VPWR.n2118 25.1912
R1252 VPWR.n2557 VPWR.n2344 25.1912
R1253 VPWR.n2546 VPWR.n2345 25.1912
R1254 VPWR.n2520 VPWR.n2348 25.1912
R1255 VPWR.n2417 VPWR.n2416 25.1912
R1256 VPWR.n2429 VPWR.n2428 25.1912
R1257 VPWR.n1645 VPWR.n1614 25.1912
R1258 VPWR.n1657 VPWR.n1656 25.1912
R1259 VPWR.n2688 VPWR.n1572 25.1912
R1260 VPWR.n2896 VPWR.n2895 25.1912
R1261 VPWR.n2866 VPWR.n2865 25.1912
R1262 VPWR.n1547 VPWR.n1520 25.1912
R1263 VPWR.n1715 VPWR.n1714 25.1912
R1264 VPWR.n2970 VPWR.n1770 25.1912
R1265 VPWR.n2019 VPWR.n2018 25.1912
R1266 VPWR.n1989 VPWR.n1988 25.1912
R1267 VPWR.n1953 VPWR.n1952 25.1912
R1268 VPWR.n1878 VPWR.n1877 25.1912
R1269 VPWR.n1347 VPWR.n1335 25.1912
R1270 VPWR.n1359 VPWR.n1358 25.1912
R1271 VPWR.n3329 VPWR.n1491 25.1912
R1272 VPWR.n3309 VPWR.n3308 25.1912
R1273 VPWR.n3168 VPWR.n3154 25.1912
R1274 VPWR.n3188 VPWR.n3187 25.1912
R1275 VPWR.n3571 VPWR.n1275 25.1912
R1276 VPWR.n3572 VPWR.n3571 25.1912
R1277 VPWR.n3497 VPWR.n3478 25.1912
R1278 VPWR.n3677 VPWR.n3676 25.1912
R1279 VPWR.n3671 VPWR.n3670 25.1912
R1280 VPWR.n3723 VPWR.n1216 25.1912
R1281 VPWR.n3717 VPWR.n3716 25.1912
R1282 VPWR.n3709 VPWR.n3708 25.1912
R1283 VPWR.n1010 VPWR.n1009 25.1912
R1284 VPWR.n1016 VPWR.n1015 25.1912
R1285 VPWR.n3927 VPWR.n3926 25.1912
R1286 VPWR.n3955 VPWR.n3954 25.1912
R1287 VPWR.n4169 VPWR.n4168 25.1912
R1288 VPWR.n736 VPWR.n735 25.1912
R1289 VPWR.n939 VPWR.n938 25.1912
R1290 VPWR.n915 VPWR.n914 25.1912
R1291 VPWR.n905 VPWR.n904 25.1912
R1292 VPWR.n887 VPWR.n822 25.1912
R1293 VPWR.n4295 VPWR.n4294 25.1912
R1294 VPWR.n4434 VPWR.n4433 25.1912
R1295 VPWR.n4782 VPWR.n4781 25.1912
R1296 VPWR.n4745 VPWR.n4741 25.1912
R1297 VPWR.n4730 VPWR.n4726 25.1912
R1298 VPWR.n285 VPWR.n284 25.1912
R1299 VPWR.n5234 VPWR.n5224 25.1912
R1300 VPWR.n5244 VPWR.n5243 25.1912
R1301 VPWR.n4962 VPWR.n4959 25.1912
R1302 VPWR.n5072 VPWR.n5071 25.1912
R1303 VPWR.n5048 VPWR.n5044 25.1912
R1304 VPWR.n5166 VPWR.n5165 25.1912
R1305 VPWR.n5189 VPWR.n5188 25.1912
R1306 VPWR.n5208 VPWR.n5204 25.1912
R1307 VPWR.n603 VPWR.n602 25.1912
R1308 VPWR.n452 VPWR.n451 25.1912
R1309 VPWR.n437 VPWR.n436 25.1912
R1310 VPWR.n420 VPWR.n419 25.1912
R1311 VPWR.n394 VPWR.n366 25.1912
R1312 VPWR.n380 VPWR.n379 25.1912
R1313 VPWR.n5988 VPWR.n160 25.1912
R1314 VPWR.n5538 VPWR.n5537 25.1912
R1315 VPWR.n5615 VPWR.n5614 25.1912
R1316 VPWR.n3518 VPWR.n3517 25.1799
R1317 VPWR.n6195 VPWR 25.1772
R1318 VPWR.n2495 VPWR.n2488 25.1014
R1319 VPWR.n6011 VPWR.n6010 24.9417
R1320 VPWR.n3178 VPWR.n3177 24.8476
R1321 VPWR.n5268 VPWR.n5267 24.8476
R1322 VPWR.n2297 VPWR.n2296 24.7608
R1323 VPWR.n2574 VPWR.n2573 24.7608
R1324 VPWR.n5703 VPWR.n5702 24.5079
R1325 VPWR.n4000 VPWR.n3999 24.5077
R1326 VPWR.n2860 VPWR.n1570 24.0694
R1327 VPWR.n4239 VPWR.n769 24.0618
R1328 VPWR.n4325 VPWR.n4324 24.0581
R1329 VPWR.n5268 VPWR.n315 24.0079
R1330 VPWR.n2635 VPWR.n2634 23.8912
R1331 VPWR.n4796 VPWR.n4795 23.8912
R1332 VPWR.n3297 VPWR.n1495 23.7181
R1333 VPWR.n3903 VPWR.n1129 23.7181
R1334 VPWR.n4718 VPWR.n4591 23.7181
R1335 VPWR.n6306 VPWR.n6305 23.7181
R1336 VPWR.n6213 VPWR.n6212 23.7181
R1337 VPWR.n3262 VPWR.n3261 23.7181
R1338 VPWR.n3261 VPWR.n3260 23.7181
R1339 VPWR.n3728 VPWR.n1211 23.7181
R1340 VPWR.n1155 VPWR.n1154 23.7181
R1341 VPWR.n1163 VPWR.n1140 23.7181
R1342 VPWR.n1164 VPWR.n1163 23.7181
R1343 VPWR.n3724 VPWR.n3723 23.7181
R1344 VPWR.n4195 VPWR.n4148 23.7181
R1345 VPWR.n708 VPWR.n707 23.7181
R1346 VPWR.n894 VPWR.n821 23.7181
R1347 VPWR.n4406 VPWR.n4400 23.7181
R1348 VPWR.n4684 VPWR.n4656 23.7181
R1349 VPWR.n275 VPWR.n263 23.7181
R1350 VPWR.n5257 VPWR.n5256 23.7181
R1351 VPWR.n540 VPWR.n501 23.7181
R1352 VPWR.n536 VPWR.n535 23.7181
R1353 VPWR.n207 VPWR.n188 23.7181
R1354 VPWR.n5530 VPWR.n5386 23.7181
R1355 VPWR.n5721 VPWR.n5720 23.7181
R1356 VPWR.n1711 VPWR.n1710 23.6786
R1357 VPWR.n390 VPWR.n366 23.6784
R1358 VPWR.n4324 VPWR.n764 23.6674
R1359 VPWR.n5494 VPWR.n5407 23.6011
R1360 VPWR.n2697 VPWR.n2696 23.5796
R1361 VPWR.n1023 VPWR.n1022 23.5618
R1362 VPWR.n4666 VPWR.n4665 23.458
R1363 VPWR.n1728 VPWR.n1727 23.3962
R1364 VPWR.n3961 VPWR.n3960 23.3962
R1365 VPWR.n6002 VPWR.n159 23.3962
R1366 VPWR.n2671 VPWR.n2670 22.9652
R1367 VPWR.n1009 VPWR.n1000 22.9652
R1368 VPWR.n1939 VPWR.n1938 22.9323
R1369 VPWR.n4552 VPWR.n4518 22.9323
R1370 VPWR.n5353 VPWR.n5352 22.9323
R1371 VPWR.n4850 VPWR.n4849 22.9278
R1372 VPWR.n1548 VPWR.n1547 22.9268
R1373 VPWR.n5230 VPWR.n5224 22.9268
R1374 VPWR.n3949 VPWR.n3948 22.9184
R1375 VPWR.n425 VPWR.n424 22.9139
R1376 VPWR.n6168 VPWR.n82 22.2123
R1377 VPWR.n2282 VPWR.n2260 22.2123
R1378 VPWR.n2297 VPWR.n2252 22.2123
R1379 VPWR.n2118 VPWR.n2077 22.2123
R1380 VPWR.n2521 VPWR.n2520 22.2123
R1381 VPWR.n2488 VPWR.n2349 22.2123
R1382 VPWR.n2416 VPWR.n2397 22.2123
R1383 VPWR.n2428 VPWR.n2393 22.2123
R1384 VPWR.n2843 VPWR.n2776 22.2123
R1385 VPWR.n2844 VPWR.n2843 22.2123
R1386 VPWR.n3330 VPWR.n3329 22.2123
R1387 VPWR.n3301 VPWR.n3300 22.2123
R1388 VPWR.n3955 VPWR.n3922 22.2123
R1389 VPWR.n4168 VPWR.n4152 22.2123
R1390 VPWR.n4254 VPWR.n4253 22.2123
R1391 VPWR.n4741 VPWR.n4590 22.2123
R1392 VPWR.n264 VPWR.n263 22.2123
R1393 VPWR.n5364 VPWR.n5325 22.2123
R1394 VPWR.n540 VPWR.n539 22.2123
R1395 VPWR.n202 VPWR.n192 22.2123
R1396 VPWR.n402 VPWR.n401 22.2123
R1397 VPWR.n380 VPWR.n370 22.2123
R1398 VPWR.n5702 VPWR.n5692 22.2123
R1399 VPWR.n5614 VPWR.n5594 22.2123
R1400 VPWR.n5088 VPWR.n5085 22.1794
R1401 VPWR.n930 VPWR.n929 21.7941
R1402 VPWR.n4149 VPWR.n4148 21.4593
R1403 VPWR.n868 VPWR.n867 21.4593
R1404 VPWR.n4861 VPWR.n4470 21.4593
R1405 VPWR.n6050 VPWR.n156 21.4593
R1406 VPWR VPWR.n3010 21.0829
R1407 VPWR.n1371 VPWR.n1331 20.7064
R1408 VPWR.n1741 VPWR.n1740 20.6735
R1409 VPWR.n3694 VPWR.n3693 20.6735
R1410 VPWR.n400 VPWR.n399 20.6735
R1411 VPWR.n5630 VPWR.n5629 20.6735
R1412 VPWR.n1740 VPWR.n1693 20.3299
R1413 VPWR.n6021 VPWR.n6020 20.3299
R1414 VPWR.n3414 VPWR.n3398 20.2952
R1415 VPWR.n1343 VPWR.n1342 19.9534
R1416 VPWR.n3493 VPWR.n3492 19.9534
R1417 VPWR.n402 VPWR.n362 19.9534
R1418 VPWR.n384 VPWR.n383 19.9534
R1419 VPWR.n2716 VPWR.n2715 19.5441
R1420 VPWR.n2728 VPWR.n2727 19.5441
R1421 VPWR.n4862 VPWR.n4861 19.5441
R1422 VPWR.n3268 VPWR.n3267 19.5347
R1423 VPWR.n3735 VPWR.n3734 19.5347
R1424 VPWR VPWR.n3502 19.1676
R1425 VPWR.n217 VPWR.n216 19.0196
R1426 VPWR.n171 VPWR.n170 19.0176
R1427 VPWR VPWR.n825 18.824
R1428 VPWR.n3022 VPWR.n3021 18.7912
R1429 VPWR.n3428 VPWR.n3427 18.7912
R1430 VPWR VPWR.n1352 18.7912
R1431 VPWR.n3892 VPWR.n1130 18.7912
R1432 VPWR.n872 VPWR.n825 18.7912
R1433 VPWR.n3620 VPWR.n3619 18.3906
R1434 VPWR.n3245 VPWR.n3244 18.1079
R1435 VPWR.n1940 VPWR.n1939 18.0711
R1436 VPWR.n5352 VPWR.n5329 18.0711
R1437 VPWR.n4473 VPWR.n4472 17.3181
R1438 VPWR VPWR.n4584 17.3181
R1439 VPWR.n5878 VPWR.n5877 17.3181
R1440 VPWR.n5525 VPWR.n5524 17.3181
R1441 VPWR.n5526 VPWR.n5525 17.3181
R1442 VPWR.n5483 VPWR.n5482 17.3181
R1443 VPWR.n6028 VPWR.n6027 17.3181
R1444 VPWR.n6054 VPWR.n6053 17.3181
R1445 VPWR.n6057 VPWR.n155 17.3181
R1446 VPWR.n5460 VPWR.n5459 17.3181
R1447 VPWR.n5735 VPWR.n5734 17.3181
R1448 VPWR.n5551 VPWR.n5550 17.3181
R1449 VPWR.n2128 VPWR.n2127 17.2853
R1450 VPWR.n3422 VPWR.n3396 17.2853
R1451 VPWR.n4183 VPWR.n4182 17.2853
R1452 VPWR.n4839 VPWR.n4838 17.2853
R1453 VPWR.n565 VPWR.n564 17.2853
R1454 VPWR.n4956 VPWR.n4943 17.2786
R1455 VPWR.n4278 VPWR.n767 17.1155
R1456 VPWR.n589 VPWR.n492 16.9088
R1457 VPWR.n4086 VPWR.n1066 16.6183
R1458 VPWR.n4196 VPWR.n4195 16.6183
R1459 VPWR.n4250 VPWR.n768 16.6183
R1460 VPWR.n1252 VPWR.n1251 16.295
R1461 VPWR.n6243 VPWR.n6242 15.9351
R1462 VPWR.n1867 VPWR.n1866 15.9351
R1463 VPWR.n2547 VPWR 15.8123
R1464 VPWR.n2850 VPWR.n2849 15.8123
R1465 VPWR.n3016 VPWR.n2992 15.8123
R1466 VPWR.n3164 VPWR.n3163 15.8123
R1467 VPWR.n3239 VPWR.n1495 15.8123
R1468 VPWR.n4014 VPWR.n1068 15.8123
R1469 VPWR.n5883 VPWR.n5858 15.8123
R1470 VPWR.n6099 VPWR.n6095 15.7727
R1471 VPWR.n6153 VPWR.n6150 15.7465
R1472 VPWR.n6158 VPWR.n6157 15.7465
R1473 VPWR.n2266 VPWR.n2265 15.7465
R1474 VPWR.n1639 VPWR.n1617 15.7465
R1475 VPWR.n2964 VPWR.n2960 15.7465
R1476 VPWR.n2954 VPWR.n2953 15.7465
R1477 VPWR.n2947 VPWR.n2946 15.7465
R1478 VPWR.n3595 VPWR.n3594 15.7465
R1479 VPWR.n4083 VPWR.n1067 15.7465
R1480 VPWR.n4334 VPWR.n4330 15.7465
R1481 VPWR.n5129 VPWR.n5103 15.7465
R1482 VPWR.n557 VPWR.n556 15.7465
R1483 VPWR.n4356 VPWR.n753 15.5434
R1484 VPWR.n4824 VPWR.n4479 15.5434
R1485 VPWR.n4527 VPWR.n4526 15.4029
R1486 VPWR.n4751 VPWR.n4750 15.4029
R1487 VPWR.n607 VPWR.n606 15.4029
R1488 VPWR.n6198 VPWR.n6197 15.1524
R1489 VPWR.n3031 VPWR.n1764 15.1524
R1490 VPWR.n384 VPWR.n369 15.1524
R1491 VPWR.n5877 VPWR.n5859 15.1524
R1492 VPWR.n2666 VPWR.n2665 15.1479
R1493 VPWR.n535 VPWR.n502 15.1443
R1494 VPWR.n2652 VPWR.n2651 15.1382
R1495 VPWR.n4698 VPWR.n4697 15.137
R1496 VPWR.n4949 VPWR.n4945 15.1307
R1497 VPWR.n1855 VPWR.n1854 15.1001
R1498 VPWR.n4969 VPWR.n4968 15.0593
R1499 VPWR.n5061 VPWR.n5060 15.0593
R1500 VPWR.n3565 VPWR.n3564 15.0265
R1501 VPWR.n5117 VPWR.n5116 15.0265
R1502 VPWR VPWR.n430 14.9338
R1503 VPWR.n3381 VPWR.n1412 14.6829
R1504 VPWR.n2303 VPWR.n2302 14.65
R1505 VPWR.n2113 VPWR.n2112 14.65
R1506 VPWR.n2483 VPWR.n2482 14.65
R1507 VPWR.n2411 VPWR.n2410 14.65
R1508 VPWR.n2423 VPWR.n2422 14.65
R1509 VPWR.n1036 VPWR.n1035 14.65
R1510 VPWR.n5370 VPWR.n5369 14.65
R1511 VPWR.n362 VPWR.n361 14.65
R1512 VPWR.n6095 VPWR.n91 14.3064
R1513 VPWR.n3896 VPWR.n1130 14.3064
R1514 VPWR.n567 VPWR.n565 14.3064
R1515 VPWR.n6230 VPWR.n6229 14.2735
R1516 VPWR.n6126 VPWR.n74 14.2735
R1517 VPWR.n6192 VPWR.n78 14.2735
R1518 VPWR.n2337 VPWR.n2072 14.2735
R1519 VPWR.n2161 VPWR.n2068 14.2735
R1520 VPWR.n2158 VPWR.n2068 14.2735
R1521 VPWR.n2593 VPWR.n2067 14.2735
R1522 VPWR.n2540 VPWR.n2536 14.2735
R1523 VPWR.n2536 VPWR.n2346 14.2735
R1524 VPWR.n2439 VPWR.n2391 14.2735
R1525 VPWR.n1622 VPWR.n1621 14.2735
R1526 VPWR.n3090 VPWR.n1576 14.2735
R1527 VPWR.n1704 VPWR.n1703 14.2735
R1528 VPWR.n3028 VPWR.n1768 14.2735
R1529 VPWR.n3028 VPWR.n1769 14.2735
R1530 VPWR.n2025 VPWR.n1815 14.2735
R1531 VPWR.n3369 VPWR.n1414 14.2735
R1532 VPWR.n3580 VPWR.n1271 14.2735
R1533 VPWR.n3588 VPWR.n1261 14.2735
R1534 VPWR.n3483 VPWR.n3482 14.2735
R1535 VPWR.n3589 VPWR.n3588 14.2735
R1536 VPWR.n3606 VPWR.n3605 14.2735
R1537 VPWR.n4059 VPWR.n4058 14.2735
R1538 VPWR.n3936 VPWR.n3931 14.2735
R1539 VPWR.n4155 VPWR.n4154 14.2735
R1540 VPWR.n724 VPWR.n723 14.2735
R1541 VPWR.n946 VPWR.n751 14.2735
R1542 VPWR.n899 VPWR.n750 14.2735
R1543 VPWR.n4267 VPWR.n4266 14.2735
R1544 VPWR.n4288 VPWR.n752 14.2735
R1545 VPWR.n4310 VPWR.n4309 14.2735
R1546 VPWR.n4422 VPWR.n4421 14.2735
R1547 VPWR.n4767 VPWR.n4476 14.2735
R1548 VPWR.n4764 VPWR.n4476 14.2735
R1549 VPWR.n5137 VPWR.n5136 14.2735
R1550 VPWR.n5337 VPWR.n5336 14.2735
R1551 VPWR.n614 VPWR.n226 14.2735
R1552 VPWR.n413 VPWR.n227 14.2735
R1553 VPWR.n410 VPWR.n227 14.2735
R1554 VPWR.n5509 VPWR.n5505 14.2735
R1555 VPWR.n5505 VPWR.n5504 14.2735
R1556 VPWR.n5596 VPWR.n5595 14.2735
R1557 VPWR.n6305 VPWR.n6304 14.1837
R1558 VPWR.n3492 VPWR.n3480 13.8921
R1559 VPWR.n2997 VPWR.n2995 13.6839
R1560 VPWR.n219 VPWR.n218 13.6753
R1561 VPWR.n2594 VPWR.n2593 13.664
R1562 VPWR.n2440 VPWR.n2439 13.664
R1563 VPWR.n52 VPWR.n51 13.6353
R1564 VPWR.n3016 VPWR.n3015 13.5534
R1565 VPWR.n1002 VPWR.n1001 13.5534
R1566 VPWR.n4010 VPWR.n1068 13.5534
R1567 VPWR.n4838 VPWR.n4471 13.5534
R1568 VPWR.n573 VPWR.n225 13.5534
R1569 VPWR.n4190 VPWR.n4149 13.5206
R1570 VPWR.n867 VPWR.n866 13.5206
R1571 VPWR.n4869 VPWR.n4469 13.5206
R1572 VPWR.n4874 VPWR.n4873 13.5206
R1573 VPWR.n5143 VPWR.n680 13.5156
R1574 VPWR.n5143 VPWR.n681 13.5156
R1575 VPWR.n4 VPWR.n3 13.177
R1576 VPWR.n6213 VPWR.n67 13.177
R1577 VPWR.n1529 VPWR.n1528 13.177
R1578 VPWR.n1849 VPWR.n1848 13.177
R1579 VPWR.n3386 VPWR.n1411 13.177
R1580 VPWR.n1342 VPWR.n1337 13.177
R1581 VPWR.n3817 VPWR.n3816 13.177
R1582 VPWR.n198 VPWR.n193 13.177
R1583 VPWR.n6198 VPWR.n73 12.8005
R1584 VPWR.n1623 VPWR.n1622 12.8005
R1585 VPWR.n2683 VPWR.n2650 12.8005
R1586 VPWR.n3437 VPWR.n1407 12.8005
R1587 VPWR.n3437 VPWR.n1409 12.8005
R1588 VPWR.n1338 VPWR.n1337 12.8005
R1589 VPWR.n1003 VPWR.n1002 12.8005
R1590 VPWR.n820 VPWR.n750 12.8005
R1591 VPWR.n4522 VPWR.n4521 12.8005
R1592 VPWR.n268 VPWR.n267 12.8005
R1593 VPWR.n5696 VPWR.n5695 12.8005
R1594 VPWR.n6169 VPWR.n6168 12.7676
R1595 VPWR.n2839 VPWR.n2838 12.4947
R1596 VPWR.n1980 VPWR.n1977 12.4947
R1597 VPWR.n3004 VPWR.n2995 12.4947
R1598 VPWR.n3378 VPWR.n3376 12.4947
R1599 VPWR.n219 VPWR.n211 12.4947
R1600 VPWR.n3974 VPWR.n1120 12.4348
R1601 VPWR.n4975 VPWR.n4974 12.424
R1602 VPWR.n6137 VPWR.n6136 12.386
R1603 VPWR.n2025 VPWR.n1814 12.0476
R1604 VPWR.n3409 VPWR.n3408 12.0476
R1605 VPWR.n5267 VPWR.n5217 12.0147
R1606 VPWR.n3665 VPWR.n1230 11.9991
R1607 VPWR.n5898 VPWR.n5857 11.9246
R1608 VPWR.n4075 VPWR.n4034 11.6711
R1609 VPWR.n4832 VPWR.n4831 11.4366
R1610 VPWR.n6242 VPWR.n47 11.2946
R1611 VPWR.n2666 VPWR.n2664 11.2946
R1612 VPWR.n1535 VPWR.n1524 11.2946
R1613 VPWR.n1854 VPWR.n1844 11.2946
R1614 VPWR.n3163 VPWR.n3162 11.2946
R1615 VPWR.n3824 VPWR.n3822 11.2946
R1616 VPWR.n4253 VPWR.n768 11.2946
R1617 VPWR.n3440 VPWR.n1406 11.0735
R1618 VPWR.n1293 VPWR.n1291 11.0735
R1619 VPWR.n1965 VPWR.n1816 10.9181
R1620 VPWR.n3321 VPWR.n3320 10.9181
R1621 VPWR.n5720 VPWR.n5719 10.9181
R1622 VPWR.n1174 VPWR.n1173 10.8853
R1623 VPWR.n1029 VPWR.n1028 10.8853
R1624 VPWR.n5271 VPWR.n314 10.8764
R1625 VPWR.n6132 VPWR.n74 10.8754
R1626 VPWR.n2670 VPWR.n2651 10.5417
R1627 VPWR.n1946 VPWR.n1945 10.5417
R1628 VPWR.n1868 VPWR.n1867 10.5417
R1629 VPWR.n3177 VPWR.n3152 10.5417
R1630 VPWR.n4560 VPWR.n4516 10.5417
R1631 VPWR.n573 VPWR.n496 10.5088
R1632 VPWR.n1120 VPWR.n1119 10.2607
R1633 VPWR.n3382 VPWR.n3381 10.1652
R1634 VPWR.n207 VPWR.n191 9.94141
R1635 VPWR.n1647 VPWR.n1612 9.78874
R1636 VPWR.n4682 VPWR.n4681 9.78874
R1637 VPWR.n938 VPWR.n811 9.41227
R1638 VPWR.n167 VPWR.n165 9.35435
R1639 VPWR.n2855 VPWR.n2772 9.3065
R1640 VPWR.n1967 VPWR.n1966 9.3065
R1641 VPWR.n3405 VPWR.n3403 9.3065
R1642 VPWR.n3325 VPWR.n3322 9.3065
R1643 VPWR.n3304 VPWR.n3302 9.3065
R1644 VPWR.n1280 VPWR.n1279 9.3065
R1645 VPWR.n3899 VPWR.n3897 9.3065
R1646 VPWR.n5112 VPWR.n5111 9.3065
R1647 VPWR.n2779 VPWR.n2778 9.3005
R1648 VPWR.n1587 VPWR.n1586 9.3005
R1649 VPWR.n2907 VPWR.n2906 9.3005
R1650 VPWR.n1913 VPWR.n1912 9.3005
R1651 VPWR.n1825 VPWR.n1824 9.3005
R1652 VPWR.n1827 VPWR.n1826 9.3005
R1653 VPWR.n1669 VPWR.n1668 9.3005
R1654 VPWR.n2939 VPWR.n2938 9.3005
R1655 VPWR.n3357 VPWR.n3356 9.3005
R1656 VPWR.n3291 VPWR.n3290 9.3005
R1657 VPWR.n3226 VPWR.n3225 9.3005
R1658 VPWR.n3228 VPWR.n3227 9.3005
R1659 VPWR.n3758 VPWR.n3757 9.3005
R1660 VPWR.n1202 VPWR.n1201 9.3005
R1661 VPWR.n1204 VPWR.n1203 9.3005
R1662 VPWR.n970 VPWR.n969 9.3005
R1663 VPWR.n4235 VPWR.n769 9.3005
R1664 VPWR.n830 VPWR.n829 9.3005
R1665 VPWR.n832 VPWR.n831 9.3005
R1666 VPWR.n4124 VPWR.n4123 9.3005
R1667 VPWR.n4352 VPWR.n4351 9.3005
R1668 VPWR.n4234 VPWR.n4233 9.3005
R1669 VPWR.n4459 VPWR.n4458 9.3005
R1670 VPWR.n4461 VPWR.n4460 9.3005
R1671 VPWR.n4492 VPWR.n4491 9.3005
R1672 VPWR.n4820 VPWR.n4819 9.3005
R1673 VPWR.n4699 VPWR.n4698 9.3005
R1674 VPWR.n238 VPWR.n237 9.3005
R1675 VPWR.n677 VPWR 9.3005
R1676 VPWR.n5301 VPWR.n5300 9.3005
R1677 VPWR.n462 VPWR.n461 9.3005
R1678 VPWR.n346 VPWR.n345 9.3005
R1679 VPWR.n5458 VPWR.n5457 9.3005
R1680 VPWR.n6059 VPWR.n6058 9.3005
R1681 VPWR.n5387 VPWR.n154 9.3005
R1682 VPWR.n5456 VPWR.n5455 9.3005
R1683 VPWR.n5402 VPWR.n5401 9.3005
R1684 VPWR.n5740 VPWR.n5739 9.3005
R1685 VPWR.n5412 VPWR.n5411 9.3005
R1686 VPWR.n5400 VPWR.n5399 9.3005
R1687 VPWR.n5666 VPWR.n5665 9.3005
R1688 VPWR.n5669 VPWR.n5668 9.3005
R1689 VPWR.n2595 VPWR.n2594 9.3005
R1690 VPWR.n2228 VPWR.n2227 9.3005
R1691 VPWR.n2441 VPWR.n2440 9.3005
R1692 VPWR.n1523 VPWR.n1522 9.29762
R1693 VPWR.n2856 VPWR.n2855 9.27733
R1694 VPWR.n2846 VPWR.n2773 9.27733
R1695 VPWR.n2839 VPWR.n2777 9.27733
R1696 VPWR.n1977 VPWR.n1812 9.27733
R1697 VPWR.n3405 VPWR.n3404 9.27733
R1698 VPWR.n3378 VPWR.n3377 9.27733
R1699 VPWR.n3325 VPWR.n3324 9.27733
R1700 VPWR.n3304 VPWR.n3303 9.27733
R1701 VPWR.n1290 VPWR.n1280 9.27733
R1702 VPWR.n3899 VPWR.n3898 9.27733
R1703 VPWR.n5112 VPWR.n5110 9.27733
R1704 VPWR.n5060 VPWR.n5058 9.05174
R1705 VPWR.n49 VPWR.n47 9.03579
R1706 VPWR.n4526 VPWR.n4520 9.03579
R1707 VPWR.n5116 VPWR.n5109 9.03579
R1708 VPWR.n2763 VPWR.n2762 9.0005
R1709 VPWR.n1568 VPWR.n1567 9.0005
R1710 VPWR.n2937 VPWR.n2936 9.0005
R1711 VPWR.n1823 VPWR.n1822 9.0005
R1712 VPWR.n1890 VPWR.n1889 9.0005
R1713 VPWR.n3224 VPWR.n3223 9.0005
R1714 VPWR.n3200 VPWR.n3199 9.0005
R1715 VPWR.n1200 VPWR.n1199 9.0005
R1716 VPWR.n1189 VPWR.n1188 9.0005
R1717 VPWR.n4356 VPWR.n4355 9.0005
R1718 VPWR.n4232 VPWR.n4231 9.0005
R1719 VPWR.n828 VPWR.n827 9.0005
R1720 VPWR.n748 VPWR.n747 9.0005
R1721 VPWR.n4824 VPWR.n4823 9.0005
R1722 VPWR.n4457 VPWR.n4456 9.0005
R1723 VPWR.n4446 VPWR.n4445 9.0005
R1724 VPWR.n4993 VPWR.n4992 9.0005
R1725 VPWR.n464 VPWR.n463 9.0005
R1726 VPWR.n5556 VPWR.n5555 9.0005
R1727 VPWR.n5454 VPWR.n5453 9.0005
R1728 VPWR.n5420 VPWR.n5419 9.0005
R1729 VPWR.n5671 VPWR.n5670 9.0005
R1730 VPWR.n2445 VPWR.n2444 9.0005
R1731 VPWR.n6202 VPWR.n70 8.96367
R1732 VPWR.n2904 VPWR.n2768 8.96367
R1733 VPWR.n596 VPWR.n491 8.96367
R1734 VPWR.n388 VPWR.n368 8.96367
R1735 VPWR.n5874 VPWR.n5860 8.96367
R1736 VPWR.n5972 VPWR.n5971 8.86972
R1737 VPWR.n3340 VPWR.n1486 8.74099
R1738 VPWR.n5332 VPWR.n5331 8.74099
R1739 VPWR.n6092 VPWR.n91 8.36851
R1740 VPWR.n49 VPWR.n48 8.28285
R1741 VPWR.n2727 VPWR.n2639 8.28285
R1742 VPWR.n4873 VPWR.n4469 8.28285
R1743 VPWR.n4152 VPWR.n4151 7.90638
R1744 VPWR.n401 VPWR.n400 7.90638
R1745 VPWR.n5629 VPWR.n5628 7.90638
R1746 VPWR.n215 VPWR.n214 7.87742
R1747 VPWR.n169 VPWR.n168 7.6548
R1748 VPWR.n2857 VPWR.n2856 7.59614
R1749 VPWR.n2849 VPWR.n2773 7.59614
R1750 VPWR.n2777 VPWR.n2776 7.59614
R1751 VPWR.n2028 VPWR.n1812 7.59614
R1752 VPWR.n1814 VPWR.n1813 7.59614
R1753 VPWR.n3377 VPWR.n1412 7.59614
R1754 VPWR.n3898 VPWR.n1129 7.59614
R1755 VPWR.n225 VPWR.n224 7.59614
R1756 VPWR.n1410 VPWR.n1407 7.58265
R1757 VPWR.n3162 VPWR.n3161 7.58265
R1758 VPWR.n3724 VPWR.n1212 7.58265
R1759 VPWR.n1946 VPWR.n1820 7.57422
R1760 VPWR.n1409 VPWR.n1408 7.57422
R1761 VPWR.n2852 VPWR.n2772 7.56696
R1762 VPWR.n2844 VPWR.n2775 7.56696
R1763 VPWR.n1966 VPWR.n1965 7.56696
R1764 VPWR.n3408 VPWR.n3403 7.56696
R1765 VPWR.n3322 VPWR.n3321 7.56696
R1766 VPWR.n3302 VPWR.n3301 7.56696
R1767 VPWR.n3557 VPWR.n1279 7.56696
R1768 VPWR.n3897 VPWR.n3896 7.56696
R1769 VPWR.n5111 VPWR.n5109 7.56696
R1770 VPWR.n567 VPWR.n566 7.56696
R1771 VPWR.n5884 VPWR.n5883 7.56696
R1772 VPWR.n191 VPWR.n190 7.55839
R1773 VPWR.n5720 VPWR.n5691 7.55839
R1774 VPWR.n3015 VPWR.n2993 7.52991
R1775 VPWR.n199 VPWR.n198 7.52991
R1776 VPWR.n5110 VPWR.n679 7.45536
R1777 VPWR.n277 VPWR.n262 7.15344
R1778 VPWR.n2256 VPWR.n2255 7.11866
R1779 VPWR.n2580 VPWR.n2579 7.11866
R1780 VPWR.n213 VPWR.n212 7.11866
R1781 VPWR.n1656 VPWR 6.77697
R1782 VPWR.n1001 VPWR.n1000 6.77697
R1783 VPWR.n3832 VPWR.n3806 6.48247
R1784 VPWR.n58 VPWR.n53 6.4005
R1785 VPWR VPWR.n2546 6.4005
R1786 VPWR.n3011 VPWR 6.4005
R1787 VPWR.n1353 VPWR 6.4005
R1788 VPWR.n868 VPWR 6.4005
R1789 VPWR.n4786 VPWR 6.4005
R1790 VPWR.n173 VPWR.n172 6.17645
R1791 VPWR.n3392 VPWR.n3391 6.158
R1792 VPWR.n1254 VPWR.n1253 6.158
R1793 VPWR.n1125 VPWR.n1124 6.158
R1794 VPWR.n63 VPWR.n61 6.02403
R1795 VPWR.n3503 VPWR 6.02403
R1796 VPWR.n3001 VPWR.n3000 6.01698
R1797 VPWR.n5968 VPWR.n173 5.96742
R1798 VPWR.n4952 VPWR.n4945 5.77927
R1799 VPWR.n3000 VPWR.n2999 5.76367
R1800 VPWR.n6197 VPWR.n70 5.75665
R1801 VPWR.n2905 VPWR.n2904 5.75665
R1802 VPWR.n2999 VPWR.n1764 5.75665
R1803 VPWR.n4660 VPWR.n4659 5.75665
R1804 VPWR.n4953 VPWR.n4952 5.75665
R1805 VPWR.n491 VPWR.n490 5.75665
R1806 VPWR.n369 VPWR.n368 5.75665
R1807 VPWR.n5860 VPWR.n5859 5.75665
R1808 VPWR.n2649 VPWR.n2646 5.75168
R1809 VPWR.n3419 VPWR.n3397 5.75168
R1810 VPWR.n3172 VPWR.n3171 5.75168
R1811 VPWR.n1145 VPWR.n1144 5.75168
R1812 VPWR.n3704 VPWR.n3703 5.75168
R1813 VPWR.n4032 VPWR.n4031 5.75168
R1814 VPWR.n4514 VPWR.n4510 5.75168
R1815 VPWR.n4595 VPWR.n4594 5.75168
R1816 VPWR.n4942 VPWR.n4941 5.75168
R1817 VPWR.n372 VPWR.n371 5.75168
R1818 VPWR.n820 VPWR.n819 5.70476
R1819 VPWR.n276 VPWR.n275 5.70476
R1820 VPWR.n3806 VPWR.n3805 5.70092
R1821 VPWR.n5888 VPWR.n5887 5.4882
R1822 VPWR.n5715 VPWR.n5711 5.4882
R1823 VPWR.n1250 VPWR.n1233 5.28304
R1824 VPWR.n4545 VPWR.n4544 5.2376
R1825 VPWR.n4472 VPWR 5.18145
R1826 VPWR.n4291 VPWR.n752 4.89462
R1827 VPWR.n6298 VPWR.n6297 4.73949
R1828 VPWR.n4276 VPWR.n767 4.73739
R1829 VPWR.n3239 VPWR 4.73093
R1830 VPWR.n46 VPWR.n45 4.6985
R1831 VPWR.n1710 VPWR.n1709 4.67352
R1832 VPWR.n4956 VPWR.n4955 4.67352
R1833 VPWR.n3949 VPWR.n3925 4.67352
R1834 VPWR.n6120 VPWR.n6119 4.67352
R1835 VPWR.n6097 VPWR.n6096 4.67352
R1836 VPWR.n6142 VPWR.n87 4.67352
R1837 VPWR.n6151 VPWR.n83 4.67352
R1838 VPWR.n6164 VPWR.n6163 4.67352
R1839 VPWR.n6255 VPWR.n6254 4.67352
R1840 VPWR.n6254 VPWR.n6253 4.67352
R1841 VPWR.n65 VPWR.n64 4.67352
R1842 VPWR.n6203 VPWR.n6202 4.67352
R1843 VPWR.n2071 VPWR.n2070 4.67352
R1844 VPWR.n2075 VPWR.n2074 4.67352
R1845 VPWR.n2157 VPWR.n2156 4.67352
R1846 VPWR.n2120 VPWR.n2119 4.67352
R1847 VPWR.n2066 VPWR.n2065 4.67352
R1848 VPWR.n2343 VPWR.n2342 4.67352
R1849 VPWR.n2538 VPWR.n2537 4.67352
R1850 VPWR.n2400 VPWR.n2399 4.67352
R1851 VPWR.n2396 VPWR.n2395 4.67352
R1852 VPWR.n2390 VPWR.n2389 4.67352
R1853 VPWR.n1630 VPWR.n1629 4.67352
R1854 VPWR.n1635 VPWR.n1634 4.67352
R1855 VPWR.n1641 VPWR.n1640 4.67352
R1856 VPWR.n1575 VPWR.n1574 4.67352
R1857 VPWR.n2649 VPWR.n2648 4.67352
R1858 VPWR.n2644 VPWR.n2643 4.67352
R1859 VPWR.n2733 VPWR.n2638 4.67352
R1860 VPWR.n2638 VPWR.n2637 4.67352
R1861 VPWR.n2767 VPWR.n2766 4.67352
R1862 VPWR.n2768 VPWR.n2767 4.67352
R1863 VPWR.n2771 VPWR.n2770 4.67352
R1864 VPWR.n1541 VPWR.n1540 4.67352
R1865 VPWR.n1542 VPWR.n1541 4.67352
R1866 VPWR.n1543 VPWR.n1542 4.67352
R1867 VPWR.n1709 VPWR.n1701 4.67352
R1868 VPWR.n1701 VPWR.n1700 4.67352
R1869 VPWR.n1766 VPWR.n1765 4.67352
R1870 VPWR.n2962 VPWR.n2961 4.67352
R1871 VPWR.n2959 VPWR.n2958 4.67352
R1872 VPWR.n2952 VPWR.n2951 4.67352
R1873 VPWR.n1973 VPWR.n1972 4.67352
R1874 VPWR.n1976 VPWR.n1975 4.67352
R1875 VPWR.n1981 VPWR.n1976 4.67352
R1876 VPWR.n1981 VPWR.n1980 4.67352
R1877 VPWR.n3006 VPWR.n3005 4.67352
R1878 VPWR.n3005 VPWR.n3004 4.67352
R1879 VPWR.n3420 VPWR.n3419 4.67352
R1880 VPWR.n1349 VPWR.n1348 4.67352
R1881 VPWR.n3361 VPWR.n3360 4.67352
R1882 VPWR.n3360 VPWR.n3359 4.67352
R1883 VPWR.n3339 VPWR.n1490 4.67352
R1884 VPWR.n3172 VPWR.n3170 4.67352
R1885 VPWR.n1278 VPWR.n1277 4.67352
R1886 VPWR.n1274 VPWR.n1273 4.67352
R1887 VPWR.n1269 VPWR.n1268 4.67352
R1888 VPWR.n3582 VPWR.n1269 4.67352
R1889 VPWR.n3582 VPWR.n3581 4.67352
R1890 VPWR.n3488 VPWR.n3487 4.67352
R1891 VPWR.n3499 VPWR.n3498 4.67352
R1892 VPWR.n1146 VPWR.n1145 4.67352
R1893 VPWR.n1260 VPWR.n1259 4.67352
R1894 VPWR.n3626 VPWR.n3625 4.67352
R1895 VPWR.n1224 VPWR.n1223 4.67352
R1896 VPWR.n1228 VPWR.n1227 4.67352
R1897 VPWR.n3657 VPWR.n1232 4.67352
R1898 VPWR.n1214 VPWR.n1213 4.67352
R1899 VPWR.n3705 VPWR.n3704 4.67352
R1900 VPWR.n3810 VPWR.n3809 4.67352
R1901 VPWR.n3829 VPWR.n3810 4.67352
R1902 VPWR.n998 VPWR.n997 4.67352
R1903 VPWR.n995 VPWR.n994 4.67352
R1904 VPWR.n1066 VPWR.n1065 4.67352
R1905 VPWR.n4040 VPWR.n4039 4.67352
R1906 VPWR.n4065 VPWR.n4037 4.67352
R1907 VPWR.n4081 VPWR.n4032 4.67352
R1908 VPWR.n3938 VPWR.n3937 4.67352
R1909 VPWR.n3942 VPWR.n3929 4.67352
R1910 VPWR.n3925 VPWR.n3924 4.67352
R1911 VPWR.n3904 VPWR.n1126 4.67352
R1912 VPWR.n1122 VPWR.n1121 4.67352
R1913 VPWR.n716 VPWR.n701 4.67352
R1914 VPWR.n945 VPWR.n944 4.67352
R1915 VPWR.n917 VPWR.n814 4.67352
R1916 VPWR.n818 VPWR.n817 4.67352
R1917 VPWR.n880 VPWR.n823 4.67352
R1918 VPWR.n4246 VPWR.n4242 4.67352
R1919 VPWR.n4246 VPWR.n4245 4.67352
R1920 VPWR.n4287 VPWR.n4286 4.67352
R1921 VPWR.n766 VPWR.n765 4.67352
R1922 VPWR.n763 VPWR.n762 4.67352
R1923 VPWR.n760 VPWR.n759 4.67352
R1924 VPWR.n4332 VPWR.n4331 4.67352
R1925 VPWR.n4867 VPWR.n4866 4.67352
R1926 VPWR.n4414 VPWR.n4399 4.67352
R1927 VPWR.n4550 VPWR.n4549 4.67352
R1928 VPWR.n4478 VPWR.n4477 4.67352
R1929 VPWR.n4791 VPWR.n4790 4.67352
R1930 VPWR.n4792 VPWR.n4791 4.67352
R1931 VPWR.n4772 VPWR.n4771 4.67352
R1932 VPWR.n4743 VPWR.n4742 4.67352
R1933 VPWR.n4728 VPWR.n4727 4.67352
R1934 VPWR.n4693 VPWR.n4651 4.67352
R1935 VPWR.n4653 VPWR.n4652 4.67352
R1936 VPWR.n4654 VPWR.n4653 4.67352
R1937 VPWR.n4658 VPWR.n4657 4.67352
R1938 VPWR.n5236 VPWR.n5235 4.67352
R1939 VPWR.n5237 VPWR.n5223 4.67352
R1940 VPWR.n4960 VPWR.n4942 4.67352
R1941 VPWR.n5121 VPWR.n5108 4.67352
R1942 VPWR.n5107 VPWR.n5106 4.67352
R1943 VPWR.n5131 VPWR.n5130 4.67352
R1944 VPWR.n5087 VPWR.n5086 4.67352
R1945 VPWR.n5216 VPWR.n5215 4.67352
R1946 VPWR.n5176 VPWR.n5175 4.67352
R1947 VPWR.n5183 VPWR.n5180 4.67352
R1948 VPWR.n5183 VPWR.n5182 4.67352
R1949 VPWR.n5182 VPWR.n5181 4.67352
R1950 VPWR.n5206 VPWR.n5205 4.67352
R1951 VPWR.n5344 VPWR.n5343 4.67352
R1952 VPWR.n5343 VPWR.n5334 4.67352
R1953 VPWR.n563 VPWR.n562 4.67352
R1954 VPWR.n555 VPWR.n554 4.67352
R1955 VPWR.n546 VPWR.n544 4.67352
R1956 VPWR.n546 VPWR.n545 4.67352
R1957 VPWR.n211 VPWR.n187 4.67352
R1958 VPWR.n584 VPWR.n495 4.67352
R1959 VPWR.n596 VPWR.n595 4.67352
R1960 VPWR.n489 VPWR.n488 4.67352
R1961 VPWR.n613 VPWR.n612 4.67352
R1962 VPWR.n352 VPWR.n351 4.67352
R1963 VPWR.n427 VPWR.n426 4.67352
R1964 VPWR.n417 VPWR.n359 4.67352
R1965 VPWR.n408 VPWR.n407 4.67352
R1966 VPWR.n396 VPWR.n395 4.67352
R1967 VPWR.n373 VPWR.n372 4.67352
R1968 VPWR.n5871 VPWR.n5865 4.67352
R1969 VPWR.n5507 VPWR.n5506 4.67352
R1970 VPWR.n5982 VPWR.n5979 4.67352
R1971 VPWR.n5982 VPWR.n5981 4.67352
R1972 VPWR.n5981 VPWR.n5980 4.67352
R1973 VPWR.n6004 VPWR.n6003 4.67352
R1974 VPWR.n5637 VPWR.n5636 4.67352
R1975 VPWR.n5636 VPWR.n5635 4.67352
R1976 VPWR.n5601 VPWR.n5600 4.67352
R1977 VPWR.n6130 VPWR.n6129 4.67352
R1978 VPWR.n6143 VPWR.n84 4.67352
R1979 VPWR.n6150 VPWR.n84 4.67352
R1980 VPWR.n6157 VPWR.n83 4.67352
R1981 VPWR.n6165 VPWR.n6164 4.67352
R1982 VPWR.n78 VPWR.n77 4.67352
R1983 VPWR.n6256 VPWR.n40 4.67352
R1984 VPWR.n6256 VPWR.n6255 4.67352
R1985 VPWR.n6220 VPWR.n65 4.67352
R1986 VPWR.n6204 VPWR.n6203 4.67352
R1987 VPWR.n2072 VPWR.n2071 4.67352
R1988 VPWR.n2166 VPWR.n2075 4.67352
R1989 VPWR.n2158 VPWR.n2157 4.67352
R1990 VPWR.n2067 VPWR.n2066 4.67352
R1991 VPWR.n2344 VPWR.n2343 4.67352
R1992 VPWR.n2410 VPWR.n2400 4.67352
R1993 VPWR.n2422 VPWR.n2396 4.67352
R1994 VPWR.n2391 VPWR.n2390 4.67352
R1995 VPWR.n1629 VPWR.n1621 4.67352
R1996 VPWR.n1640 VPWR.n1639 4.67352
R1997 VPWR.n1576 VPWR.n1575 4.67352
R1998 VPWR.n2684 VPWR.n2649 4.67352
R1999 VPWR.n2865 VPWR.n2771 4.67352
R2000 VPWR.n1543 VPWR.n1520 4.67352
R2001 VPWR.n2960 VPWR.n2959 4.67352
R2002 VPWR.n2953 VPWR.n2952 4.67352
R2003 VPWR.n2946 VPWR.n1773 4.67352
R2004 VPWR.n2019 VPWR.n1973 4.67352
R2005 VPWR.n1952 VPWR.n1951 4.67352
R2006 VPWR.n3419 VPWR.n3418 4.67352
R2007 VPWR.n3394 VPWR.n3393 4.67352
R2008 VPWR.n3428 VPWR.n3394 4.67352
R2009 VPWR.n1348 VPWR.n1347 4.67352
R2010 VPWR.n3369 VPWR.n3368 4.67352
R2011 VPWR.n3323 VPWR.n1491 4.67352
R2012 VPWR.n3308 VPWR.n1493 4.67352
R2013 VPWR.n3173 VPWR.n3172 4.67352
R2014 VPWR.n3565 VPWR.n1278 4.67352
R2015 VPWR.n3572 VPWR.n1274 4.67352
R2016 VPWR.n3581 VPWR.n3580 4.67352
R2017 VPWR.n3487 VPWR.n3482 4.67352
R2018 VPWR.n3498 VPWR.n3497 4.67352
R2019 VPWR.n1145 VPWR.n1141 4.67352
R2020 VPWR.n3589 VPWR.n1260 4.67352
R2021 VPWR.n1257 VPWR.n1256 4.67352
R2022 VPWR.n3595 VPWR.n1257 4.67352
R2023 VPWR.n3625 VPWR.n1255 4.67352
R2024 VPWR.n3619 VPWR.n1255 4.67352
R2025 VPWR.n3694 VPWR.n1224 4.67352
R2026 VPWR.n3671 VPWR.n1228 4.67352
R2027 VPWR.n1232 VPWR.n1231 4.67352
R2028 VPWR.n3704 VPWR.n3702 4.67352
R2029 VPWR.n4048 VPWR.n4042 4.67352
R2030 VPWR.n4059 VPWR.n4040 4.67352
R2031 VPWR.n4033 VPWR.n4032 4.67352
R2032 VPWR.n3937 VPWR.n3936 4.67352
R2033 VPWR.n3921 VPWR.n3920 4.67352
R2034 VPWR.n3961 VPWR.n3921 4.67352
R2035 VPWR.n1123 VPWR.n1122 4.67352
R2036 VPWR.n4188 VPWR.n4187 4.67352
R2037 VPWR.n723 VPWR.n701 4.67352
R2038 VPWR.n946 VPWR.n945 4.67352
R2039 VPWR.n922 VPWR.n921 4.67352
R2040 VPWR.n813 VPWR.n812 4.67352
R2041 VPWR.n929 VPWR.n813 4.67352
R2042 VPWR.n904 VPWR.n818 4.67352
R2043 VPWR.n882 VPWR.n880 4.67352
R2044 VPWR.n881 VPWR.n822 4.67352
R2045 VPWR.n873 VPWR.n872 4.67352
R2046 VPWR.n4240 VPWR.n4239 4.67352
R2047 VPWR.n4288 VPWR.n4287 4.67352
R2048 VPWR.n4309 VPWR.n766 4.67352
R2049 VPWR.n4330 VPWR.n760 4.67352
R2050 VPWR.n4331 VPWR.n753 4.67352
R2051 VPWR.n4421 VPWR.n4399 4.67352
R2052 VPWR.n4479 VPWR.n4478 4.67352
R2053 VPWR.n4697 VPWR.n4651 4.67352
R2054 VPWR.n4665 VPWR.n4657 4.67352
R2055 VPWR.n313 VPWR.n312 4.67352
R2056 VPWR.n314 VPWR.n313 4.67352
R2057 VPWR.n5237 VPWR.n5236 4.67352
R2058 VPWR.n5235 VPWR.n5234 4.67352
R2059 VPWR.n5243 VPWR.n5219 4.67352
R2060 VPWR.n4967 VPWR.n4942 4.67352
R2061 VPWR.n4955 VPWR.n4954 4.67352
R2062 VPWR.n5117 VPWR.n5108 4.67352
R2063 VPWR.n5130 VPWR.n5129 4.67352
R2064 VPWR.n5137 VPWR.n5099 4.67352
R2065 VPWR.n5088 VPWR.n5087 4.67352
R2066 VPWR.n5048 VPWR.n5047 4.67352
R2067 VPWR.n4979 VPWR.n4939 4.67352
R2068 VPWR.n5217 VPWR.n5216 4.67352
R2069 VPWR.n5180 VPWR.n316 4.67352
R2070 VPWR.n5335 VPWR.n5334 4.67352
R2071 VPWR.n5336 VPWR.n5335 4.67352
R2072 VPWR.n5328 VPWR.n5327 4.67352
R2073 VPWR.n5327 VPWR.n5326 4.67352
R2074 VPWR.n564 VPWR.n563 4.67352
R2075 VPWR.n556 VPWR.n555 4.67352
R2076 VPWR.n577 VPWR.n496 4.67352
R2077 VPWR.n585 VPWR.n584 4.67352
R2078 VPWR.n585 VPWR.n492 4.67352
R2079 VPWR.n595 VPWR.n594 4.67352
R2080 VPWR.n602 VPWR.n488 4.67352
R2081 VPWR.n614 VPWR.n613 4.67352
R2082 VPWR.n413 VPWR.n359 4.67352
R2083 VPWR.n407 VPWR.n361 4.67352
R2084 VPWR.n395 VPWR.n394 4.67352
R2085 VPWR.n372 VPWR.n228 4.67352
R2086 VPWR.n5537 VPWR.n5385 4.67352
R2087 VPWR.n5600 VPWR.n5595 4.67352
R2088 VPWR.n390 VPWR.n389 4.67351
R2089 VPWR.n426 VPWR.n425 4.67206
R2090 VPWR.n3006 VPWR.n2994 4.67166
R2091 VPWR.n4322 VPWR.n764 4.66266
R2092 VPWR.n2676 VPWR.n2675 4.65944
R2093 VPWR.n5081 VPWR.n5080 4.65624
R2094 VPWR.n425 VPWR.n356 4.65278
R2095 VPWR.n3490 VPWR.n3480 4.65151
R2096 VPWR.n5141 VPWR.n680 4.65151
R2097 VPWR.n5096 VPWR.n681 4.65151
R2098 VPWR.n3950 VPWR.n3949 4.65148
R2099 VPWR.n391 VPWR.n390 4.65148
R2100 VPWR.n6100 VPWR.n6099 4.65147
R2101 VPWR.n1710 VPWR.n1697 4.65147
R2102 VPWR.n4957 VPWR.n4956 4.65147
R2103 VPWR.n2815 VPWR.n2814 4.6505
R2104 VPWR.n2843 VPWR.n2842 4.6505
R2105 VPWR.n2851 VPWR.n2850 4.6505
R2106 VPWR.n2859 VPWR.n1570 4.6505
R2107 VPWR.n2875 VPWR.n2874 4.6505
R2108 VPWR.n2883 VPWR.n2882 4.6505
R2109 VPWR.n1530 VPWR.n1529 4.6505
R2110 VPWR.n1532 VPWR.n1531 4.6505
R2111 VPWR.n1533 VPWR.n1524 4.6505
R2112 VPWR.n1535 VPWR 4.6505
R2113 VPWR.n2820 VPWR.n2819 4.6505
R2114 VPWR.n2822 VPWR.n2821 4.6505
R2115 VPWR.n2826 VPWR.n2825 4.6505
R2116 VPWR.n2830 VPWR.n2829 4.6505
R2117 VPWR.n2832 VPWR.n2831 4.6505
R2118 VPWR.n2834 VPWR.n2833 4.6505
R2119 VPWR.n2836 VPWR.n2835 4.6505
R2120 VPWR.n2838 VPWR.n2837 4.6505
R2121 VPWR.n2849 VPWR.n2774 4.6505
R2122 VPWR.n2889 VPWR.n2888 4.6505
R2123 VPWR.n2897 VPWR.n2896 4.6505
R2124 VPWR.n2899 VPWR.n2898 4.6505
R2125 VPWR.n2902 VPWR.n2768 4.6505
R2126 VPWR.n2727 VPWR.n2726 4.6505
R2127 VPWR.n2725 VPWR.n2639 4.6505
R2128 VPWR.n2715 VPWR.n2714 4.6505
R2129 VPWR.n2707 VPWR.n2640 4.6505
R2130 VPWR.n2706 VPWR.n2641 4.6505
R2131 VPWR.n2699 VPWR.n2642 4.6505
R2132 VPWR.n2683 VPWR.n2682 4.6505
R2133 VPWR.n2681 VPWR.n2650 4.6505
R2134 VPWR.n2670 VPWR.n2669 4.6505
R2135 VPWR.n2668 VPWR.n2651 4.6505
R2136 VPWR.n2664 VPWR.n2663 4.6505
R2137 VPWR.n2662 VPWR.n2654 4.6505
R2138 VPWR.n1626 VPWR.n1622 4.6505
R2139 VPWR.n1654 VPWR.n1653 4.6505
R2140 VPWR.n1652 VPWR.n1611 4.6505
R2141 VPWR.n1651 VPWR.n1650 4.6505
R2142 VPWR.n1649 VPWR.n1612 4.6505
R2143 VPWR.n1648 VPWR.n1647 4.6505
R2144 VPWR.n1646 VPWR.n1613 4.6505
R2145 VPWR.n1645 VPWR.n1644 4.6505
R2146 VPWR.n1643 VPWR.n1614 4.6505
R2147 VPWR.n1642 VPWR.n1641 4.6505
R2148 VPWR.n1640 VPWR.n1615 4.6505
R2149 VPWR.n1639 VPWR.n1638 4.6505
R2150 VPWR.n1637 VPWR.n1617 4.6505
R2151 VPWR.n1636 VPWR.n1635 4.6505
R2152 VPWR.n1634 VPWR.n1618 4.6505
R2153 VPWR.n1633 VPWR.n1632 4.6505
R2154 VPWR.n1631 VPWR.n1630 4.6505
R2155 VPWR.n1629 VPWR.n1628 4.6505
R2156 VPWR.n1627 VPWR.n1621 4.6505
R2157 VPWR.n1660 VPWR.n1659 4.6505
R2158 VPWR.n1658 VPWR.n1657 4.6505
R2159 VPWR.n1656 VPWR.n1655 4.6505
R2160 VPWR.n2736 VPWR.n2735 4.6505
R2161 VPWR.n2733 VPWR.n2732 4.6505
R2162 VPWR.n2729 VPWR.n2728 4.6505
R2163 VPWR.n2724 VPWR.n2723 4.6505
R2164 VPWR.n2721 VPWR.n2720 4.6505
R2165 VPWR.n2719 VPWR.n2718 4.6505
R2166 VPWR.n2717 VPWR.n2716 4.6505
R2167 VPWR.n2713 VPWR.n2712 4.6505
R2168 VPWR.n2711 VPWR.n2710 4.6505
R2169 VPWR.n2709 VPWR.n2708 4.6505
R2170 VPWR.n2705 VPWR.n2704 4.6505
R2171 VPWR.n2703 VPWR.n2702 4.6505
R2172 VPWR.n2701 VPWR.n2700 4.6505
R2173 VPWR.n2698 VPWR.n2697 4.6505
R2174 VPWR.n2696 VPWR.n2695 4.6505
R2175 VPWR.n2692 VPWR.n2691 4.6505
R2176 VPWR.n2690 VPWR.n1572 4.6505
R2177 VPWR.n2689 VPWR.n2688 4.6505
R2178 VPWR.n2685 VPWR.n2684 4.6505
R2179 VPWR.n2680 VPWR.n2679 4.6505
R2180 VPWR.n2678 VPWR.n2677 4.6505
R2181 VPWR.n2672 VPWR.n2671 4.6505
R2182 VPWR VPWR.n2666 4.6505
R2183 VPWR.n2661 VPWR.n2660 4.6505
R2184 VPWR.n2659 VPWR.n2658 4.6505
R2185 VPWR.n2655 VPWR.n1576 4.6505
R2186 VPWR.n2895 VPWR.n2894 4.6505
R2187 VPWR.n2893 VPWR.n2892 4.6505
R2188 VPWR.n2891 VPWR.n2890 4.6505
R2189 VPWR.n2887 VPWR.n2886 4.6505
R2190 VPWR.n2885 VPWR.n2884 4.6505
R2191 VPWR.n2881 VPWR.n2880 4.6505
R2192 VPWR.n2879 VPWR.n2878 4.6505
R2193 VPWR.n2877 VPWR.n2876 4.6505
R2194 VPWR.n2873 VPWR.n2872 4.6505
R2195 VPWR.n2871 VPWR.n2870 4.6505
R2196 VPWR.n2869 VPWR.n2868 4.6505
R2197 VPWR.n2867 VPWR.n2866 4.6505
R2198 VPWR.n2865 VPWR.n2864 4.6505
R2199 VPWR.n2861 VPWR.n2860 4.6505
R2200 VPWR.n2849 VPWR.n2848 4.6505
R2201 VPWR.n1536 VPWR.n1535 4.6505
R2202 VPWR.n1540 VPWR.n1539 4.6505
R2203 VPWR.n1544 VPWR.n1543 4.6505
R2204 VPWR.n1545 VPWR.n1520 4.6505
R2205 VPWR.n1547 VPWR.n1546 4.6505
R2206 VPWR.n1549 VPWR.n1548 4.6505
R2207 VPWR.n1551 VPWR.n1550 4.6505
R2208 VPWR.n1554 VPWR.n1553 4.6505
R2209 VPWR.n1556 VPWR.n1555 4.6505
R2210 VPWR.n1558 VPWR.n1557 4.6505
R2211 VPWR.n1560 VPWR.n1559 4.6505
R2212 VPWR.n1563 VPWR.n1562 4.6505
R2213 VPWR.n1934 VPWR.n1933 4.6505
R2214 VPWR.n1939 VPWR.n1821 4.6505
R2215 VPWR.n1943 VPWR.n1942 4.6505
R2216 VPWR.n1945 VPWR.n1944 4.6505
R2217 VPWR.n1946 VPWR.n1819 4.6505
R2218 VPWR.n1947 VPWR.n1946 4.6505
R2219 VPWR.n1956 VPWR.n1955 4.6505
R2220 VPWR.n2025 VPWR.n2024 4.6505
R2221 VPWR.n1850 VPWR.n1849 4.6505
R2222 VPWR.n1853 VPWR.n1844 4.6505
R2223 VPWR.n1867 VPWR.n1840 4.6505
R2224 VPWR.n1869 VPWR.n1868 4.6505
R2225 VPWR.n1875 VPWR.n1874 4.6505
R2226 VPWR.n1936 VPWR.n1935 4.6505
R2227 VPWR.n1938 VPWR.n1937 4.6505
R2228 VPWR.n1970 VPWR.n1814 4.6505
R2229 VPWR.n1996 VPWR.n1995 4.6505
R2230 VPWR.n1988 VPWR.n1987 4.6505
R2231 VPWR.n1986 VPWR.n1985 4.6505
R2232 VPWR.n1982 VPWR.n1981 4.6505
R2233 VPWR.n1980 VPWR.n1979 4.6505
R2234 VPWR.n2980 VPWR.n2979 4.6505
R2235 VPWR.n3026 VPWR.n1768 4.6505
R2236 VPWR.n3021 VPWR.n3020 4.6505
R2237 VPWR.n3019 VPWR.n2991 4.6505
R2238 VPWR.n3018 VPWR.n2992 4.6505
R2239 VPWR.n3015 VPWR.n3014 4.6505
R2240 VPWR.n1737 VPWR.n1694 4.6505
R2241 VPWR.n1724 VPWR.n1696 4.6505
R2242 VPWR.n1738 VPWR.n1693 4.6505
R2243 VPWR.n1736 VPWR.n1735 4.6505
R2244 VPWR.n1733 VPWR.n1732 4.6505
R2245 VPWR.n1731 VPWR.n1730 4.6505
R2246 VPWR.n1729 VPWR.n1728 4.6505
R2247 VPWR.n1727 VPWR.n1726 4.6505
R2248 VPWR.n1725 VPWR.n1695 4.6505
R2249 VPWR.n1723 VPWR.n1722 4.6505
R2250 VPWR.n1720 VPWR.n1719 4.6505
R2251 VPWR.n1718 VPWR.n1717 4.6505
R2252 VPWR.n1716 VPWR.n1715 4.6505
R2253 VPWR.n1714 VPWR.n1713 4.6505
R2254 VPWR.n1712 VPWR.n1711 4.6505
R2255 VPWR.n1709 VPWR 4.6505
R2256 VPWR.n1708 VPWR.n1701 4.6505
R2257 VPWR.n1705 VPWR.n1704 4.6505
R2258 VPWR.n1744 VPWR.n1743 4.6505
R2259 VPWR.n1742 VPWR.n1741 4.6505
R2260 VPWR.n1740 VPWR.n1739 4.6505
R2261 VPWR.n2944 VPWR.n2943 4.6505
R2262 VPWR.n2945 VPWR.n1773 4.6505
R2263 VPWR.n2946 VPWR 4.6505
R2264 VPWR VPWR.n2947 4.6505
R2265 VPWR.n2951 VPWR.n2950 4.6505
R2266 VPWR VPWR.n2954 4.6505
R2267 VPWR.n2958 VPWR.n2957 4.6505
R2268 VPWR.n2965 VPWR.n2964 4.6505
R2269 VPWR.n2968 VPWR.n1770 4.6505
R2270 VPWR.n2970 VPWR.n2969 4.6505
R2271 VPWR.n2972 VPWR.n2971 4.6505
R2272 VPWR.n2974 VPWR.n2973 4.6505
R2273 VPWR.n2976 VPWR.n2975 4.6505
R2274 VPWR.n2978 VPWR.n2977 4.6505
R2275 VPWR.n2982 VPWR.n2981 4.6505
R2276 VPWR.n2985 VPWR.n2984 4.6505
R2277 VPWR.n2987 VPWR.n2986 4.6505
R2278 VPWR.n2989 VPWR.n2988 4.6505
R2279 VPWR.n2990 VPWR.n1769 4.6505
R2280 VPWR.n3028 VPWR.n3027 4.6505
R2281 VPWR.n3023 VPWR.n3022 4.6505
R2282 VPWR.n3012 VPWR.n3011 4.6505
R2283 VPWR.n3010 VPWR.n3009 4.6505
R2284 VPWR.n3007 VPWR.n3006 4.6505
R2285 VPWR.n3004 VPWR.n3003 4.6505
R2286 VPWR.n1990 VPWR.n1989 4.6505
R2287 VPWR.n1992 VPWR.n1991 4.6505
R2288 VPWR.n1994 VPWR.n1993 4.6505
R2289 VPWR.n1998 VPWR.n1997 4.6505
R2290 VPWR.n2000 VPWR.n1999 4.6505
R2291 VPWR.n2002 VPWR.n2001 4.6505
R2292 VPWR.n2004 VPWR.n2003 4.6505
R2293 VPWR.n2006 VPWR.n2005 4.6505
R2294 VPWR.n2008 VPWR.n2007 4.6505
R2295 VPWR.n2010 VPWR.n2009 4.6505
R2296 VPWR.n2012 VPWR.n2011 4.6505
R2297 VPWR.n2014 VPWR.n2013 4.6505
R2298 VPWR.n2016 VPWR.n2015 4.6505
R2299 VPWR.n2018 VPWR.n2017 4.6505
R2300 VPWR.n2020 VPWR.n2019 4.6505
R2301 VPWR.n2023 VPWR.n1815 4.6505
R2302 VPWR.n1969 VPWR.n1814 4.6505
R2303 VPWR.n1963 VPWR.n1816 4.6505
R2304 VPWR.n1962 VPWR.n1961 4.6505
R2305 VPWR.n1960 VPWR.n1959 4.6505
R2306 VPWR.n1958 VPWR.n1957 4.6505
R2307 VPWR.n1954 VPWR.n1953 4.6505
R2308 VPWR.n1951 VPWR.n1950 4.6505
R2309 VPWR.n1941 VPWR.n1940 4.6505
R2310 VPWR.n1852 VPWR.n1851 4.6505
R2311 VPWR.n1854 VPWR 4.6505
R2312 VPWR.n1857 VPWR.n1856 4.6505
R2313 VPWR.n1861 VPWR.n1860 4.6505
R2314 VPWR.n1866 VPWR.n1865 4.6505
R2315 VPWR.n1871 VPWR.n1870 4.6505
R2316 VPWR.n1873 VPWR.n1872 4.6505
R2317 VPWR.n1877 VPWR.n1876 4.6505
R2318 VPWR.n1879 VPWR.n1878 4.6505
R2319 VPWR.n1882 VPWR.n1881 4.6505
R2320 VPWR.n1885 VPWR.n1884 4.6505
R2321 VPWR.n3371 VPWR.n1414 4.6505
R2322 VPWR.n3381 VPWR 4.6505
R2323 VPWR.n3383 VPWR.n3382 4.6505
R2324 VPWR.n3387 VPWR.n3386 4.6505
R2325 VPWR.n3427 VPWR.n3426 4.6505
R2326 VPWR.n3425 VPWR.n3395 4.6505
R2327 VPWR.n3424 VPWR.n3396 4.6505
R2328 VPWR.n3416 VPWR.n3398 4.6505
R2329 VPWR.n3411 VPWR.n3401 4.6505
R2330 VPWR.n3264 VPWR.n3234 4.6505
R2331 VPWR.n3257 VPWR.n3237 4.6505
R2332 VPWR.n3244 VPWR.n3243 4.6505
R2333 VPWR.n3242 VPWR.n3238 4.6505
R2334 VPWR.n3241 VPWR.n3239 4.6505
R2335 VPWR.n3298 VPWR.n3297 4.6505
R2336 VPWR.n3312 VPWR.n3311 4.6505
R2337 VPWR.n3331 VPWR.n3330 4.6505
R2338 VPWR.n3335 VPWR.n3334 4.6505
R2339 VPWR.n3340 VPWR.n1487 4.6505
R2340 VPWR.n3163 VPWR.n3155 4.6505
R2341 VPWR VPWR.n3164 4.6505
R2342 VPWR.n3175 VPWR.n3152 4.6505
R2343 VPWR.n3177 VPWR.n3176 4.6505
R2344 VPWR.n3183 VPWR.n3182 4.6505
R2345 VPWR.n3275 VPWR.n3274 4.6505
R2346 VPWR.n3271 VPWR.n3270 4.6505
R2347 VPWR.n3269 VPWR.n3268 4.6505
R2348 VPWR.n3256 VPWR.n3255 4.6505
R2349 VPWR.n3254 VPWR.n3253 4.6505
R2350 VPWR.n3252 VPWR.n3251 4.6505
R2351 VPWR.n3250 VPWR.n3249 4.6505
R2352 VPWR.n3248 VPWR.n3247 4.6505
R2353 VPWR.n3246 VPWR.n3245 4.6505
R2354 VPWR.n3308 VPWR.n3307 4.6505
R2355 VPWR.n3328 VPWR.n1491 4.6505
R2356 VPWR.n3339 VPWR.n3338 4.6505
R2357 VPWR.n3362 VPWR.n3361 4.6505
R2358 VPWR.n3366 VPWR.n3365 4.6505
R2359 VPWR.n3368 VPWR.n3367 4.6505
R2360 VPWR.n3370 VPWR.n3369 4.6505
R2361 VPWR.n3389 VPWR.n1407 4.6505
R2362 VPWR.n3433 VPWR.n3432 4.6505
R2363 VPWR.n3429 VPWR.n3428 4.6505
R2364 VPWR.n3423 VPWR.n3422 4.6505
R2365 VPWR.n3418 VPWR.n3417 4.6505
R2366 VPWR.n3408 VPWR.n3402 4.6505
R2367 VPWR.n3408 VPWR.n3407 4.6505
R2368 VPWR.n1371 VPWR.n1370 4.6505
R2369 VPWR.n1368 VPWR.n1332 4.6505
R2370 VPWR.n1342 VPWR.n1341 4.6505
R2371 VPWR.n1367 VPWR.n1366 4.6505
R2372 VPWR.n1364 VPWR.n1363 4.6505
R2373 VPWR.n1362 VPWR.n1361 4.6505
R2374 VPWR.n1360 VPWR.n1359 4.6505
R2375 VPWR.n1358 VPWR.n1357 4.6505
R2376 VPWR.n1356 VPWR.n1355 4.6505
R2377 VPWR.n1354 VPWR.n1353 4.6505
R2378 VPWR.n1352 VPWR.n1351 4.6505
R2379 VPWR.n1350 VPWR.n1349 4.6505
R2380 VPWR.n1348 VPWR.n1334 4.6505
R2381 VPWR.n1347 VPWR.n1346 4.6505
R2382 VPWR VPWR.n1335 4.6505
R2383 VPWR.n1345 VPWR.n1344 4.6505
R2384 VPWR.n1343 VPWR.n1336 4.6505
R2385 VPWR.n1375 VPWR.n1374 4.6505
R2386 VPWR.n1373 VPWR.n1372 4.6505
R2387 VPWR.n1369 VPWR.n1331 4.6505
R2388 VPWR.n3413 VPWR.n3412 4.6505
R2389 VPWR.n3415 VPWR.n3414 4.6505
R2390 VPWR.n3437 VPWR.n3436 4.6505
R2391 VPWR.n3390 VPWR.n1407 4.6505
R2392 VPWR.n3385 VPWR.n3384 4.6505
R2393 VPWR.n3376 VPWR.n3375 4.6505
R2394 VPWR.n3374 VPWR.n3373 4.6505
R2395 VPWR.n3333 VPWR.n3332 4.6505
R2396 VPWR.n3329 VPWR 4.6505
R2397 VPWR.n3320 VPWR.n3319 4.6505
R2398 VPWR.n3318 VPWR.n3317 4.6505
R2399 VPWR.n3316 VPWR.n3315 4.6505
R2400 VPWR.n3314 VPWR.n3313 4.6505
R2401 VPWR.n3310 VPWR.n3309 4.6505
R2402 VPWR.n3300 VPWR.n3299 4.6505
R2403 VPWR.n3258 VPWR.n3236 4.6505
R2404 VPWR.n3260 VPWR.n3259 4.6505
R2405 VPWR.n3263 VPWR.n3262 4.6505
R2406 VPWR.n3265 VPWR.n3233 4.6505
R2407 VPWR.n3267 VPWR.n3266 4.6505
R2408 VPWR.n3165 VPWR.n3154 4.6505
R2409 VPWR.n3168 VPWR.n3167 4.6505
R2410 VPWR.n3174 VPWR.n3173 4.6505
R2411 VPWR.n3179 VPWR.n3178 4.6505
R2412 VPWR.n3181 VPWR.n3180 4.6505
R2413 VPWR.n3185 VPWR.n3184 4.6505
R2414 VPWR.n3187 VPWR.n3186 4.6505
R2415 VPWR.n3189 VPWR.n3188 4.6505
R2416 VPWR.n3192 VPWR.n3191 4.6505
R2417 VPWR.n3195 VPWR.n3194 4.6505
R2418 VPWR.n3605 VPWR.n3604 4.6505
R2419 VPWR.n3586 VPWR.n1261 4.6505
R2420 VPWR.n3564 VPWR.n3563 4.6505
R2421 VPWR.n3731 VPWR.n1210 4.6505
R2422 VPWR.n3693 VPWR.n3692 4.6505
R2423 VPWR.n3685 VPWR.n1225 4.6505
R2424 VPWR.n1154 VPWR.n1153 4.6505
R2425 VPWR.n1167 VPWR.n1166 4.6505
R2426 VPWR.n1173 VPWR.n1172 4.6505
R2427 VPWR.n3742 VPWR.n3741 4.6505
R2428 VPWR.n3738 VPWR.n3737 4.6505
R2429 VPWR.n3736 VPWR.n3735 4.6505
R2430 VPWR.n3721 VPWR.n1216 4.6505
R2431 VPWR.n3718 VPWR.n3717 4.6505
R2432 VPWR.n3706 VPWR.n3705 4.6505
R2433 VPWR.n3701 VPWR.n3700 4.6505
R2434 VPWR.n3668 VPWR.n1229 4.6505
R2435 VPWR.n3663 VPWR.n1230 4.6505
R2436 VPWR.n3662 VPWR.n3661 4.6505
R2437 VPWR.n3658 VPWR.n3657 4.6505
R2438 VPWR.n3656 VPWR.n3655 4.6505
R2439 VPWR.n3627 VPWR.n3626 4.6505
R2440 VPWR.n3625 VPWR.n3624 4.6505
R2441 VPWR.n3614 VPWR.n3613 4.6505
R2442 VPWR.n3609 VPWR.n3608 4.6505
R2443 VPWR.n3600 VPWR.n3599 4.6505
R2444 VPWR.n3596 VPWR.n3595 4.6505
R2445 VPWR.n3577 VPWR.n3576 4.6505
R2446 VPWR.n3573 VPWR.n3572 4.6505
R2447 VPWR.n3513 VPWR.n3475 4.6505
R2448 VPWR.n3492 VPWR.n3491 4.6505
R2449 VPWR.n3515 VPWR.n3514 4.6505
R2450 VPWR.n3512 VPWR.n3511 4.6505
R2451 VPWR.n3510 VPWR.n3509 4.6505
R2452 VPWR.n3508 VPWR.n3507 4.6505
R2453 VPWR.n3506 VPWR.n3505 4.6505
R2454 VPWR.n3504 VPWR.n3503 4.6505
R2455 VPWR.n3502 VPWR.n3501 4.6505
R2456 VPWR.n3500 VPWR.n3499 4.6505
R2457 VPWR.n3498 VPWR.n3477 4.6505
R2458 VPWR.n3497 VPWR.n3496 4.6505
R2459 VPWR VPWR.n3478 4.6505
R2460 VPWR.n3495 VPWR.n3494 4.6505
R2461 VPWR.n3493 VPWR.n3479 4.6505
R2462 VPWR.n3489 VPWR.n3488 4.6505
R2463 VPWR.n3487 VPWR.n3486 4.6505
R2464 VPWR.n3485 VPWR.n3482 4.6505
R2465 VPWR.n3525 VPWR.n3524 4.6505
R2466 VPWR.n3523 VPWR.n3522 4.6505
R2467 VPWR.n3521 VPWR.n3520 4.6505
R2468 VPWR.n3519 VPWR.n3518 4.6505
R2469 VPWR.n3517 VPWR.n3516 4.6505
R2470 VPWR.n3558 VPWR.n3557 4.6505
R2471 VPWR.n3560 VPWR.n3559 4.6505
R2472 VPWR.n3562 VPWR.n3561 4.6505
R2473 VPWR.n3566 VPWR.n3565 4.6505
R2474 VPWR.n3569 VPWR.n1275 4.6505
R2475 VPWR.n3571 VPWR.n3570 4.6505
R2476 VPWR.n3580 VPWR.n3579 4.6505
R2477 VPWR.n3583 VPWR.n3582 4.6505
R2478 VPWR.n3588 VPWR.n3587 4.6505
R2479 VPWR.n3590 VPWR.n3589 4.6505
R2480 VPWR.n3594 VPWR.n3593 4.6505
R2481 VPWR.n3607 VPWR.n3606 4.6505
R2482 VPWR.n3611 VPWR.n3610 4.6505
R2483 VPWR.n3616 VPWR.n3615 4.6505
R2484 VPWR.n3618 VPWR.n3617 4.6505
R2485 VPWR.n3621 VPWR.n3620 4.6505
R2486 VPWR.n3665 VPWR.n3664 4.6505
R2487 VPWR.n3667 VPWR.n3666 4.6505
R2488 VPWR.n3670 VPWR.n3669 4.6505
R2489 VPWR.n3672 VPWR.n3671 4.6505
R2490 VPWR.n3676 VPWR.n3675 4.6505
R2491 VPWR.n3678 VPWR.n3677 4.6505
R2492 VPWR.n3680 VPWR.n3679 4.6505
R2493 VPWR.n3682 VPWR.n3681 4.6505
R2494 VPWR.n3684 VPWR.n3683 4.6505
R2495 VPWR.n3687 VPWR.n3686 4.6505
R2496 VPWR.n3689 VPWR.n3688 4.6505
R2497 VPWR.n3691 VPWR.n3690 4.6505
R2498 VPWR.n3695 VPWR.n3694 4.6505
R2499 VPWR.n3699 VPWR.n3698 4.6505
R2500 VPWR.n3708 VPWR.n3707 4.6505
R2501 VPWR.n3710 VPWR.n3709 4.6505
R2502 VPWR.n3712 VPWR.n3711 4.6505
R2503 VPWR.n3714 VPWR.n3713 4.6505
R2504 VPWR.n3716 VPWR.n3715 4.6505
R2505 VPWR.n3723 VPWR.n3722 4.6505
R2506 VPWR.n3728 VPWR.n3727 4.6505
R2507 VPWR.n3730 VPWR.n3729 4.6505
R2508 VPWR.n3732 VPWR.n1209 4.6505
R2509 VPWR.n3734 VPWR.n3733 4.6505
R2510 VPWR.n1149 VPWR.n1148 4.6505
R2511 VPWR.n1152 VPWR.n1141 4.6505
R2512 VPWR.n1156 VPWR.n1155 4.6505
R2513 VPWR.n1158 VPWR.n1157 4.6505
R2514 VPWR.n1160 VPWR.n1159 4.6505
R2515 VPWR.n1161 VPWR.n1140 4.6505
R2516 VPWR.n1165 VPWR.n1164 4.6505
R2517 VPWR.n1169 VPWR.n1168 4.6505
R2518 VPWR.n1171 VPWR.n1170 4.6505
R2519 VPWR.n1175 VPWR.n1174 4.6505
R2520 VPWR.n1177 VPWR.n1176 4.6505
R2521 VPWR.n1179 VPWR.n1178 4.6505
R2522 VPWR.n1181 VPWR.n1180 4.6505
R2523 VPWR.n1184 VPWR.n1183 4.6505
R2524 VPWR.n4005 VPWR.n4004 4.6505
R2525 VPWR.n4011 VPWR.n4010 4.6505
R2526 VPWR.n4014 VPWR.n4013 4.6505
R2527 VPWR.n4018 VPWR.n4017 4.6505
R2528 VPWR.n4083 VPWR.n4030 4.6505
R2529 VPWR.n4077 VPWR.n4034 4.6505
R2530 VPWR.n4058 VPWR.n4057 4.6505
R2531 VPWR.n4054 VPWR.n4041 4.6505
R2532 VPWR.n3887 VPWR.n3886 4.6505
R2533 VPWR.n3894 VPWR.n1130 4.6505
R2534 VPWR.n3911 VPWR.n1127 4.6505
R2535 VPWR.n3971 VPWR.n3919 4.6505
R2536 VPWR.n3956 VPWR.n3922 4.6505
R2537 VPWR.n3818 VPWR.n3817 4.6505
R2538 VPWR.n3822 VPWR.n3821 4.6505
R2539 VPWR.n3824 VPWR 4.6505
R2540 VPWR.n3889 VPWR.n3888 4.6505
R2541 VPWR.n3891 VPWR.n3890 4.6505
R2542 VPWR.n3893 VPWR.n3892 4.6505
R2543 VPWR.n3911 VPWR.n3910 4.6505
R2544 VPWR.n3943 VPWR.n3942 4.6505
R2545 VPWR.n3941 VPWR.n3940 4.6505
R2546 VPWR.n3939 VPWR.n3938 4.6505
R2547 VPWR.n3993 VPWR.n3992 4.6505
R2548 VPWR.n3995 VPWR.n3994 4.6505
R2549 VPWR.n3997 VPWR.n3996 4.6505
R2550 VPWR.n3999 VPWR.n3998 4.6505
R2551 VPWR.n4001 VPWR.n4000 4.6505
R2552 VPWR.n4081 VPWR.n4080 4.6505
R2553 VPWR.n4064 VPWR.n4063 4.6505
R2554 VPWR.n4060 VPWR.n4059 4.6505
R2555 VPWR.n4049 VPWR 4.6505
R2556 VPWR.n4046 VPWR.n4042 4.6505
R2557 VPWR.n4043 VPWR.n1066 4.6505
R2558 VPWR.n1035 VPWR.n1034 4.6505
R2559 VPWR.n1029 VPWR 4.6505
R2560 VPWR.n1007 VPWR.n1000 4.6505
R2561 VPWR.n1031 VPWR.n1030 4.6505
R2562 VPWR.n1028 VPWR.n1027 4.6505
R2563 VPWR.n1024 VPWR.n1023 4.6505
R2564 VPWR.n1022 VPWR.n1021 4.6505
R2565 VPWR.n1020 VPWR.n1019 4.6505
R2566 VPWR.n1018 VPWR.n1017 4.6505
R2567 VPWR.n1016 VPWR 4.6505
R2568 VPWR.n1015 VPWR.n1014 4.6505
R2569 VPWR.n1011 VPWR.n1010 4.6505
R2570 VPWR.n1009 VPWR.n1008 4.6505
R2571 VPWR.n1039 VPWR.n1038 4.6505
R2572 VPWR.n1037 VPWR.n1036 4.6505
R2573 VPWR.n1033 VPWR.n1032 4.6505
R2574 VPWR.n4048 VPWR.n4047 4.6505
R2575 VPWR.n4051 VPWR.n4050 4.6505
R2576 VPWR.n4053 VPWR.n4052 4.6505
R2577 VPWR.n4056 VPWR.n4055 4.6505
R2578 VPWR.n4066 VPWR.n4065 4.6505
R2579 VPWR.n4072 VPWR.n4071 4.6505
R2580 VPWR.n4074 VPWR.n4073 4.6505
R2581 VPWR.n4076 VPWR.n4075 4.6505
R2582 VPWR.n4029 VPWR.n1067 4.6505
R2583 VPWR.n4028 VPWR.n4027 4.6505
R2584 VPWR.n4026 VPWR.n4025 4.6505
R2585 VPWR.n4024 VPWR.n4023 4.6505
R2586 VPWR.n4022 VPWR.n4021 4.6505
R2587 VPWR.n4020 VPWR.n4019 4.6505
R2588 VPWR.n4016 VPWR.n4015 4.6505
R2589 VPWR.n4007 VPWR.n4006 4.6505
R2590 VPWR.n4003 VPWR.n4002 4.6505
R2591 VPWR.n3936 VPWR.n3935 4.6505
R2592 VPWR.n3946 VPWR.n3926 4.6505
R2593 VPWR.n3948 VPWR.n3947 4.6505
R2594 VPWR.n3954 VPWR.n3953 4.6505
R2595 VPWR VPWR.n3955 4.6505
R2596 VPWR.n3958 VPWR.n3957 4.6505
R2597 VPWR.n3960 VPWR.n3959 4.6505
R2598 VPWR.n3962 VPWR.n3961 4.6505
R2599 VPWR.n3966 VPWR.n3965 4.6505
R2600 VPWR.n3968 VPWR.n3967 4.6505
R2601 VPWR.n3970 VPWR.n3969 4.6505
R2602 VPWR.n3918 VPWR.n1123 4.6505
R2603 VPWR.n3915 VPWR.n3914 4.6505
R2604 VPWR.n3909 VPWR.n1126 4.6505
R2605 VPWR.n3907 VPWR.n3906 4.6505
R2606 VPWR.n3903 VPWR.n3902 4.6505
R2607 VPWR.n3820 VPWR.n3819 4.6505
R2608 VPWR.n3824 VPWR.n3812 4.6505
R2609 VPWR.n3824 VPWR.n3811 4.6505
R2610 VPWR.n3825 VPWR.n3824 4.6505
R2611 VPWR.n3829 VPWR.n3828 4.6505
R2612 VPWR.n3831 VPWR.n3830 4.6505
R2613 VPWR VPWR.n768 4.6505
R2614 VPWR.n4253 VPWR.n4252 4.6505
R2615 VPWR.n4257 VPWR.n4256 4.6505
R2616 VPWR.n4268 VPWR.n4267 4.6505
R2617 VPWR.n4290 VPWR.n752 4.6505
R2618 VPWR.n4311 VPWR.n4310 4.6505
R2619 VPWR.n4313 VPWR.n4312 4.6505
R2620 VPWR.n862 VPWR.n861 4.6505
R2621 VPWR.n867 VPWR.n826 4.6505
R2622 VPWR.n870 VPWR.n825 4.6505
R2623 VPWR.n891 VPWR.n890 4.6505
R2624 VPWR.n900 VPWR.n899 4.6505
R2625 VPWR.n912 VPWR.n911 4.6505
R2626 VPWR.n725 VPWR.n724 4.6505
R2627 VPWR.n729 VPWR.n728 4.6505
R2628 VPWR.n864 VPWR.n863 4.6505
R2629 VPWR.n866 VPWR.n865 4.6505
R2630 VPWR.n873 VPWR.n824 4.6505
R2631 VPWR.n877 VPWR.n876 4.6505
R2632 VPWR.n878 VPWR.n823 4.6505
R2633 VPWR.n880 VPWR.n879 4.6505
R2634 VPWR.n883 VPWR.n882 4.6505
R2635 VPWR.n921 VPWR.n920 4.6505
R2636 VPWR.n923 VPWR.n922 4.6505
R2637 VPWR.n925 VPWR.n924 4.6505
R2638 VPWR.n929 VPWR.n928 4.6505
R2639 VPWR.n940 VPWR.n939 4.6505
R2640 VPWR.n947 VPWR.n946 4.6505
R2641 VPWR.n4239 VPWR.n4238 4.6505
R2642 VPWR.n4247 VPWR.n4246 4.6505
R2643 VPWR.n4251 VPWR.n4250 4.6505
R2644 VPWR.n4271 VPWR.n4270 4.6505
R2645 VPWR.n4273 VPWR.n4272 4.6505
R2646 VPWR.n4275 VPWR.n4274 4.6505
R2647 VPWR.n4282 VPWR.n4281 4.6505
R2648 VPWR.n4319 VPWR.n4318 4.6505
R2649 VPWR.n4326 VPWR.n4325 4.6505
R2650 VPWR.n4330 VPWR.n4329 4.6505
R2651 VPWR.n4335 VPWR.n4334 4.6505
R2652 VPWR.n4338 VPWR.n753 4.6505
R2653 VPWR.n4192 VPWR.n4149 4.6505
R2654 VPWR.n4182 VPWR.n4181 4.6505
R2655 VPWR.n4167 VPWR.n4152 4.6505
R2656 VPWR.n4191 VPWR.n4190 4.6505
R2657 VPWR.n4184 VPWR.n4183 4.6505
R2658 VPWR.n4180 VPWR.n4150 4.6505
R2659 VPWR.n4179 VPWR.n4178 4.6505
R2660 VPWR.n4177 VPWR.n4176 4.6505
R2661 VPWR.n4174 VPWR.n4173 4.6505
R2662 VPWR.n4172 VPWR.n4171 4.6505
R2663 VPWR.n4170 VPWR.n4169 4.6505
R2664 VPWR.n4168 VPWR 4.6505
R2665 VPWR.n4165 VPWR.n4164 4.6505
R2666 VPWR.n4163 VPWR.n4162 4.6505
R2667 VPWR.n4160 VPWR.n4159 4.6505
R2668 VPWR.n4158 VPWR.n4157 4.6505
R2669 VPWR.n4156 VPWR.n4155 4.6505
R2670 VPWR.n4199 VPWR.n4198 4.6505
R2671 VPWR.n4197 VPWR.n4196 4.6505
R2672 VPWR.n4195 VPWR.n4194 4.6505
R2673 VPWR.n4193 VPWR.n4148 4.6505
R2674 VPWR.n4324 VPWR.n4323 4.6505
R2675 VPWR.n4317 VPWR.n4316 4.6505
R2676 VPWR.n4315 VPWR.n4314 4.6505
R2677 VPWR.n4309 VPWR.n4308 4.6505
R2678 VPWR.n4305 VPWR.n4304 4.6505
R2679 VPWR.n4303 VPWR.n4302 4.6505
R2680 VPWR.n4301 VPWR.n4300 4.6505
R2681 VPWR.n4298 VPWR.n4297 4.6505
R2682 VPWR.n4296 VPWR.n4295 4.6505
R2683 VPWR.n4294 VPWR.n4293 4.6505
R2684 VPWR.n4292 VPWR.n4291 4.6505
R2685 VPWR.n4289 VPWR.n4288 4.6505
R2686 VPWR.n4280 VPWR.n4279 4.6505
R2687 VPWR.n4278 VPWR.n4277 4.6505
R2688 VPWR.n4266 VPWR.n4265 4.6505
R2689 VPWR.n4264 VPWR.n4263 4.6505
R2690 VPWR.n4262 VPWR.n4261 4.6505
R2691 VPWR.n4260 VPWR.n4259 4.6505
R2692 VPWR.n4255 VPWR.n4254 4.6505
R2693 VPWR.n938 VPWR.n937 4.6505
R2694 VPWR.n935 VPWR.n934 4.6505
R2695 VPWR.n933 VPWR.n932 4.6505
R2696 VPWR.n931 VPWR.n930 4.6505
R2697 VPWR.n919 VPWR.n814 4.6505
R2698 VPWR.n918 VPWR.n917 4.6505
R2699 VPWR.n914 VPWR.n913 4.6505
R2700 VPWR.n910 VPWR.n909 4.6505
R2701 VPWR.n908 VPWR.n907 4.6505
R2702 VPWR.n906 VPWR.n905 4.6505
R2703 VPWR.n904 VPWR.n903 4.6505
R2704 VPWR.n898 VPWR.n750 4.6505
R2705 VPWR.n895 VPWR.n894 4.6505
R2706 VPWR.n893 VPWR.n892 4.6505
R2707 VPWR.n889 VPWR.n888 4.6505
R2708 VPWR.n887 VPWR.n886 4.6505
R2709 VPWR.n885 VPWR.n822 4.6505
R2710 VPWR.n872 VPWR.n871 4.6505
R2711 VPWR.n869 VPWR.n868 4.6505
R2712 VPWR.n707 VPWR.n706 4.6505
R2713 VPWR.n708 VPWR.n703 4.6505
R2714 VPWR.n708 VPWR 4.6505
R2715 VPWR.n711 VPWR.n710 4.6505
R2716 VPWR.n713 VPWR.n712 4.6505
R2717 VPWR.n715 VPWR.n714 4.6505
R2718 VPWR.n719 VPWR.n718 4.6505
R2719 VPWR.n723 VPWR.n722 4.6505
R2720 VPWR.n727 VPWR.n726 4.6505
R2721 VPWR.n731 VPWR.n730 4.6505
R2722 VPWR.n735 VPWR.n734 4.6505
R2723 VPWR.n737 VPWR.n736 4.6505
R2724 VPWR.n740 VPWR.n739 4.6505
R2725 VPWR.n743 VPWR.n742 4.6505
R2726 VPWR.n4878 VPWR.n4468 4.6505
R2727 VPWR.n4873 VPWR.n4872 4.6505
R2728 VPWR.n4871 VPWR.n4469 4.6505
R2729 VPWR.n4861 VPWR.n4860 4.6505
R2730 VPWR.n4838 VPWR.n4837 4.6505
R2731 VPWR.n4836 VPWR.n4471 4.6505
R2732 VPWR.n4835 VPWR.n4472 4.6505
R2733 VPWR.n4669 VPWR.n4668 4.6505
R2734 VPWR.n4423 VPWR.n4422 4.6505
R2735 VPWR.n4427 VPWR.n4426 4.6505
R2736 VPWR.n4877 VPWR.n4876 4.6505
R2737 VPWR.n4875 VPWR.n4874 4.6505
R2738 VPWR.n4858 VPWR.n4857 4.6505
R2739 VPWR.n4855 VPWR.n4854 4.6505
R2740 VPWR.n4853 VPWR.n4852 4.6505
R2741 VPWR.n4851 VPWR.n4850 4.6505
R2742 VPWR.n4833 VPWR.n4832 4.6505
R2743 VPWR.n4691 VPWR.n4690 4.6505
R2744 VPWR.n4694 VPWR.n4693 4.6505
R2745 VPWR.n4697 VPWR.n4696 4.6505
R2746 VPWR.n4716 VPWR.n4591 4.6505
R2747 VPWR.n4740 VPWR.n4590 4.6505
R2748 VPWR.n4752 VPWR.n4751 4.6505
R2749 VPWR.n4754 VPWR.n4753 4.6505
R2750 VPWR.n4756 VPWR.n4755 4.6505
R2751 VPWR.n4766 VPWR.n4476 4.6505
R2752 VPWR.n4773 VPWR.n4586 4.6505
R2753 VPWR.n4773 VPWR.n4585 4.6505
R2754 VPWR.n4785 VPWR.n4784 4.6505
R2755 VPWR.n4560 VPWR.n4559 4.6505
R2756 VPWR.n4557 VPWR.n4517 4.6505
R2757 VPWR.n4554 VPWR.n4518 4.6505
R2758 VPWR.n4526 VPWR 4.6505
R2759 VPWR.n4525 VPWR.n4520 4.6505
R2760 VPWR.n4556 VPWR.n4555 4.6505
R2761 VPWR.n4553 VPWR.n4552 4.6505
R2762 VPWR.n4546 VPWR.n4545 4.6505
R2763 VPWR.n4544 VPWR.n4543 4.6505
R2764 VPWR.n4542 VPWR.n4519 4.6505
R2765 VPWR.n4541 VPWR.n4540 4.6505
R2766 VPWR.n4539 VPWR.n4538 4.6505
R2767 VPWR.n4537 VPWR.n4536 4.6505
R2768 VPWR.n4535 VPWR.n4534 4.6505
R2769 VPWR.n4532 VPWR.n4531 4.6505
R2770 VPWR.n4530 VPWR.n4529 4.6505
R2771 VPWR.n4528 VPWR.n4527 4.6505
R2772 VPWR.n4562 VPWR.n4561 4.6505
R2773 VPWR.n4558 VPWR.n4516 4.6505
R2774 VPWR.n4722 VPWR.n4721 4.6505
R2775 VPWR.n4724 VPWR.n4723 4.6505
R2776 VPWR.n4726 VPWR.n4725 4.6505
R2777 VPWR.n4731 VPWR.n4730 4.6505
R2778 VPWR.n4735 VPWR.n4734 4.6505
R2779 VPWR.n4737 VPWR.n4736 4.6505
R2780 VPWR.n4739 VPWR.n4738 4.6505
R2781 VPWR.n4741 VPWR 4.6505
R2782 VPWR.n4746 VPWR.n4745 4.6505
R2783 VPWR.n4750 VPWR.n4749 4.6505
R2784 VPWR.n4759 VPWR.n4758 4.6505
R2785 VPWR.n4761 VPWR.n4760 4.6505
R2786 VPWR.n4763 VPWR.n4762 4.6505
R2787 VPWR.n4765 VPWR.n4764 4.6505
R2788 VPWR.n4768 VPWR.n4767 4.6505
R2789 VPWR.n4771 VPWR.n4770 4.6505
R2790 VPWR.n4777 VPWR.n4776 4.6505
R2791 VPWR.n4779 VPWR.n4778 4.6505
R2792 VPWR.n4781 VPWR.n4780 4.6505
R2793 VPWR.n4783 VPWR.n4782 4.6505
R2794 VPWR.n4787 VPWR.n4786 4.6505
R2795 VPWR.n4790 VPWR.n4789 4.6505
R2796 VPWR.n4791 VPWR.n4582 4.6505
R2797 VPWR.n4793 VPWR.n4792 4.6505
R2798 VPWR.n4795 VPWR.n4794 4.6505
R2799 VPWR.n4800 VPWR.n4799 4.6505
R2800 VPWR.n4802 VPWR.n4801 4.6505
R2801 VPWR.n4805 VPWR.n4479 4.6505
R2802 VPWR.n4715 VPWR.n4714 4.6505
R2803 VPWR.n4718 VPWR.n4717 4.6505
R2804 VPWR.n4720 VPWR.n4719 4.6505
R2805 VPWR.n4689 VPWR.n4654 4.6505
R2806 VPWR.n4685 VPWR.n4684 4.6505
R2807 VPWR.n4683 VPWR.n4682 4.6505
R2808 VPWR.n4681 VPWR.n4680 4.6505
R2809 VPWR.n4679 VPWR.n4678 4.6505
R2810 VPWR.n4677 VPWR.n4676 4.6505
R2811 VPWR.n4675 VPWR.n4674 4.6505
R2812 VPWR.n4673 VPWR.n4672 4.6505
R2813 VPWR.n4671 VPWR.n4670 4.6505
R2814 VPWR.n4667 VPWR.n4666 4.6505
R2815 VPWR.n4665 VPWR.n4664 4.6505
R2816 VPWR.n4840 VPWR.n4839 4.6505
R2817 VPWR.n4842 VPWR.n4841 4.6505
R2818 VPWR.n4844 VPWR.n4843 4.6505
R2819 VPWR.n4847 VPWR.n4846 4.6505
R2820 VPWR.n4849 VPWR.n4848 4.6505
R2821 VPWR.n4859 VPWR.n4470 4.6505
R2822 VPWR.n4863 VPWR.n4862 4.6505
R2823 VPWR.n4870 VPWR.n4869 4.6505
R2824 VPWR.n4404 VPWR.n4400 4.6505
R2825 VPWR.n4406 VPWR.n4405 4.6505
R2826 VPWR.n4406 VPWR 4.6505
R2827 VPWR.n4409 VPWR.n4408 4.6505
R2828 VPWR.n4411 VPWR.n4410 4.6505
R2829 VPWR.n4413 VPWR.n4412 4.6505
R2830 VPWR.n4417 VPWR.n4416 4.6505
R2831 VPWR.n4421 VPWR.n4420 4.6505
R2832 VPWR.n4425 VPWR.n4424 4.6505
R2833 VPWR.n4429 VPWR.n4428 4.6505
R2834 VPWR.n4433 VPWR.n4432 4.6505
R2835 VPWR.n4435 VPWR.n4434 4.6505
R2836 VPWR.n4438 VPWR.n4437 4.6505
R2837 VPWR.n4441 VPWR.n4440 4.6505
R2838 VPWR.n5044 VPWR.n5043 4.6505
R2839 VPWR.n5062 VPWR.n5061 4.6505
R2840 VPWR.n5085 VPWR.n5084 4.6505
R2841 VPWR.n5136 VPWR.n5135 4.6505
R2842 VPWR.n5116 VPWR.n5115 4.6505
R2843 VPWR.n4950 VPWR.n4949 4.6505
R2844 VPWR VPWR.n4943 4.6505
R2845 VPWR.n4968 VPWR.n4940 4.6505
R2846 VPWR.n4970 VPWR.n4969 4.6505
R2847 VPWR.n4974 VPWR.n4973 4.6505
R2848 VPWR.n5049 VPWR.n5048 4.6505
R2849 VPWR.n5054 VPWR.n5053 4.6505
R2850 VPWR.n5056 VPWR.n5055 4.6505
R2851 VPWR.n5058 VPWR.n5057 4.6505
R2852 VPWR.n5060 VPWR.n682 4.6505
R2853 VPWR.n5060 VPWR.n5059 4.6505
R2854 VPWR.n5073 VPWR.n5072 4.6505
R2855 VPWR.n5077 VPWR.n5076 4.6505
R2856 VPWR.n5132 VPWR.n5131 4.6505
R2857 VPWR.n5127 VPWR.n5103 4.6505
R2858 VPWR.n5124 VPWR.n5123 4.6505
R2859 VPWR.n5121 VPWR.n5120 4.6505
R2860 VPWR.n5170 VPWR.n317 4.6505
R2861 VPWR.n5202 VPWR.n5201 4.6505
R2862 VPWR.n5268 VPWR.n5213 4.6505
R2863 VPWR.n5267 VPWR.n5266 4.6505
R2864 VPWR.n5256 VPWR.n5255 4.6505
R2865 VPWR.n5250 VPWR.n5218 4.6505
R2866 VPWR.n282 VPWR.n261 4.6505
R2867 VPWR.n279 VPWR.n262 4.6505
R2868 VPWR VPWR.n263 4.6505
R2869 VPWR.n273 VPWR.n264 4.6505
R2870 VPWR.n270 VPWR.n265 4.6505
R2871 VPWR.n281 VPWR.n280 4.6505
R2872 VPWR.n272 VPWR.n271 4.6505
R2873 VPWR.n292 VPWR.n291 4.6505
R2874 VPWR.n290 VPWR.n289 4.6505
R2875 VPWR.n288 VPWR.n287 4.6505
R2876 VPWR.n286 VPWR.n285 4.6505
R2877 VPWR.n284 VPWR.n283 4.6505
R2878 VPWR.n5169 VPWR.n5168 4.6505
R2879 VPWR.n5173 VPWR.n5172 4.6505
R2880 VPWR.n5177 VPWR.n5176 4.6505
R2881 VPWR.n5178 VPWR.n316 4.6505
R2882 VPWR.n5180 VPWR.n5179 4.6505
R2883 VPWR.n5184 VPWR.n5183 4.6505
R2884 VPWR.n5188 VPWR.n5187 4.6505
R2885 VPWR.n5190 VPWR.n5189 4.6505
R2886 VPWR.n5192 VPWR.n5191 4.6505
R2887 VPWR.n5194 VPWR.n5193 4.6505
R2888 VPWR.n5196 VPWR.n5195 4.6505
R2889 VPWR.n5198 VPWR.n5197 4.6505
R2890 VPWR.n5200 VPWR.n5199 4.6505
R2891 VPWR.n5204 VPWR.n5203 4.6505
R2892 VPWR.n5209 VPWR.n5208 4.6505
R2893 VPWR.n5212 VPWR.n315 4.6505
R2894 VPWR.n5265 VPWR.n5217 4.6505
R2895 VPWR.n5262 VPWR.n5261 4.6505
R2896 VPWR.n5260 VPWR.n5259 4.6505
R2897 VPWR.n5258 VPWR.n5257 4.6505
R2898 VPWR.n5254 VPWR.n5253 4.6505
R2899 VPWR.n5252 VPWR.n5251 4.6505
R2900 VPWR.n5249 VPWR.n5248 4.6505
R2901 VPWR.n5247 VPWR.n5246 4.6505
R2902 VPWR.n5245 VPWR.n5244 4.6505
R2903 VPWR.n5243 VPWR.n5242 4.6505
R2904 VPWR.n5241 VPWR.n5219 4.6505
R2905 VPWR.n5238 VPWR.n5237 4.6505
R2906 VPWR.n5234 VPWR.n5233 4.6505
R2907 VPWR.n5232 VPWR.n5224 4.6505
R2908 VPWR.n5231 VPWR.n5230 4.6505
R2909 VPWR.n5227 VPWR.n314 4.6505
R2910 VPWR.n5163 VPWR.n5162 4.6505
R2911 VPWR.n5165 VPWR.n5164 4.6505
R2912 VPWR.n5167 VPWR.n5166 4.6505
R2913 VPWR.n5118 VPWR.n5117 4.6505
R2914 VPWR.n5129 VPWR.n5128 4.6505
R2915 VPWR.n5138 VPWR.n5137 4.6505
R2916 VPWR.n5143 VPWR.n5142 4.6505
R2917 VPWR.n5095 VPWR.n5094 4.6505
R2918 VPWR.n5093 VPWR.n5092 4.6505
R2919 VPWR.n5089 VPWR.n5088 4.6505
R2920 VPWR.n5083 VPWR.n5082 4.6505
R2921 VPWR.n5079 VPWR.n5078 4.6505
R2922 VPWR.n5075 VPWR.n5074 4.6505
R2923 VPWR.n5071 VPWR.n5070 4.6505
R2924 VPWR.n5069 VPWR.n5068 4.6505
R2925 VPWR.n5067 VPWR.n5066 4.6505
R2926 VPWR.n5065 VPWR.n5064 4.6505
R2927 VPWR.n4959 VPWR.n4958 4.6505
R2928 VPWR.n4963 VPWR.n4962 4.6505
R2929 VPWR.n4967 VPWR.n4966 4.6505
R2930 VPWR.n4972 VPWR.n4971 4.6505
R2931 VPWR.n4976 VPWR.n4975 4.6505
R2932 VPWR.n4979 VPWR.n4978 4.6505
R2933 VPWR.n4982 VPWR.n4981 4.6505
R2934 VPWR.n4984 VPWR.n4983 4.6505
R2935 VPWR.n4988 VPWR.n4987 4.6505
R2936 VPWR.n537 VPWR.n536 4.6505
R2937 VPWR.n539 VPWR.n538 4.6505
R2938 VPWR.n565 VPWR.n497 4.6505
R2939 VPWR.n574 VPWR.n573 4.6505
R2940 VPWR.n589 VPWR.n588 4.6505
R2941 VPWR.n606 VPWR.n605 4.6505
R2942 VPWR.n198 VPWR.n197 4.6505
R2943 VPWR.n200 VPWR.n199 4.6505
R2944 VPWR.n201 VPWR.n192 4.6505
R2945 VPWR.n544 VPWR.n543 4.6505
R2946 VPWR.n547 VPWR.n546 4.6505
R2947 VPWR.n550 VPWR.n549 4.6505
R2948 VPWR.n558 VPWR.n557 4.6505
R2949 VPWR.n562 VPWR.n561 4.6505
R2950 VPWR.n571 VPWR.n225 4.6505
R2951 VPWR.n572 VPWR.n225 4.6505
R2952 VPWR.n580 VPWR.n579 4.6505
R2953 VPWR.n584 VPWR.n583 4.6505
R2954 VPWR.n597 VPWR.n596 4.6505
R2955 VPWR.n608 VPWR.n607 4.6505
R2956 VPWR.n615 VPWR.n614 4.6505
R2957 VPWR.n449 VPWR.n350 4.6505
R2958 VPWR.n412 VPWR.n227 4.6505
R2959 VPWR.n404 VPWR.n362 4.6505
R2960 VPWR.n401 VPWR.n363 4.6505
R2961 VPWR.n400 VPWR 4.6505
R2962 VPWR.n381 VPWR.n370 4.6505
R2963 VPWR.n5369 VPWR.n5368 4.6505
R2964 VPWR.n5365 VPWR.n5325 4.6505
R2965 VPWR.n5363 VPWR.n5362 4.6505
R2966 VPWR.n5352 VPWR.n5351 4.6505
R2967 VPWR.n5349 VPWR.n5330 4.6505
R2968 VPWR VPWR.n5364 4.6505
R2969 VPWR.n5361 VPWR.n5328 4.6505
R2970 VPWR.n5358 VPWR.n5357 4.6505
R2971 VPWR.n5356 VPWR.n5355 4.6505
R2972 VPWR.n5354 VPWR.n5353 4.6505
R2973 VPWR.n5350 VPWR.n5329 4.6505
R2974 VPWR.n5347 VPWR.n5346 4.6505
R2975 VPWR.n5343 VPWR.n5342 4.6505
R2976 VPWR.n5341 VPWR.n5334 4.6505
R2977 VPWR.n5373 VPWR.n5372 4.6505
R2978 VPWR.n5371 VPWR.n5370 4.6505
R2979 VPWR.n5367 VPWR.n5366 4.6505
R2980 VPWR.n459 VPWR.n458 4.6505
R2981 VPWR.n455 VPWR.n454 4.6505
R2982 VPWR.n453 VPWR.n452 4.6505
R2983 VPWR.n451 VPWR.n450 4.6505
R2984 VPWR.n448 VPWR.n447 4.6505
R2985 VPWR.n446 VPWR.n445 4.6505
R2986 VPWR.n444 VPWR.n443 4.6505
R2987 VPWR.n442 VPWR.n441 4.6505
R2988 VPWR.n440 VPWR.n439 4.6505
R2989 VPWR.n438 VPWR.n437 4.6505
R2990 VPWR.n436 VPWR.n435 4.6505
R2991 VPWR.n432 VPWR.n431 4.6505
R2992 VPWR.n430 VPWR.n429 4.6505
R2993 VPWR.n428 VPWR.n427 4.6505
R2994 VPWR.n426 VPWR.n355 4.6505
R2995 VPWR.n424 VPWR.n423 4.6505
R2996 VPWR.n422 VPWR.n357 4.6505
R2997 VPWR.n421 VPWR.n420 4.6505
R2998 VPWR.n419 VPWR.n358 4.6505
R2999 VPWR.n417 VPWR.n416 4.6505
R3000 VPWR.n415 VPWR.n359 4.6505
R3001 VPWR.n414 VPWR.n413 4.6505
R3002 VPWR.n411 VPWR.n410 4.6505
R3003 VPWR.n408 VPWR.n360 4.6505
R3004 VPWR.n407 VPWR.n406 4.6505
R3005 VPWR.n405 VPWR.n361 4.6505
R3006 VPWR.n403 VPWR.n402 4.6505
R3007 VPWR.n399 VPWR.n398 4.6505
R3008 VPWR.n397 VPWR.n396 4.6505
R3009 VPWR.n395 VPWR.n365 4.6505
R3010 VPWR.n394 VPWR.n393 4.6505
R3011 VPWR.n392 VPWR.n366 4.6505
R3012 VPWR.n389 VPWR.n367 4.6505
R3013 VPWR.n388 VPWR.n387 4.6505
R3014 VPWR.n385 VPWR.n384 4.6505
R3015 VPWR.n383 VPWR.n382 4.6505
R3016 VPWR VPWR.n380 4.6505
R3017 VPWR.n379 VPWR.n378 4.6505
R3018 VPWR.n375 VPWR.n228 4.6505
R3019 VPWR.n604 VPWR.n603 4.6505
R3020 VPWR.n602 VPWR.n601 4.6505
R3021 VPWR.n591 VPWR.n590 4.6505
R3022 VPWR.n587 VPWR.n492 4.6505
R3023 VPWR.n586 VPWR.n585 4.6505
R3024 VPWR.n577 VPWR.n576 4.6505
R3025 VPWR.n554 VPWR.n553 4.6505
R3026 VPWR.n541 VPWR.n540 4.6505
R3027 VPWR.n535 VPWR.n534 4.6505
R3028 VPWR.n202 VPWR 4.6505
R3029 VPWR.n204 VPWR.n203 4.6505
R3030 VPWR.n205 VPWR.n188 4.6505
R3031 VPWR.n207 VPWR.n189 4.6505
R3032 VPWR.n208 VPWR.n207 4.6505
R3033 VPWR.n211 VPWR.n210 4.6505
R3034 VPWR.n5465 VPWR.n5464 4.6505
R3035 VPWR.n5473 VPWR.n5472 4.6505
R3036 VPWR.n5493 VPWR.n5492 4.6505
R3037 VPWR.n5505 VPWR.n5405 4.6505
R3038 VPWR.n5541 VPWR.n5540 4.6505
R3039 VPWR.n5992 VPWR.n5991 4.6505
R3040 VPWR.n6015 VPWR.n6014 4.6505
R3041 VPWR.n6020 VPWR.n6019 4.6505
R3042 VPWR.n6043 VPWR.n6042 4.6505
R3043 VPWR.n6048 VPWR.n156 4.6505
R3044 VPWR.n5872 VPWR.n5862 4.6505
R3045 VPWR.n5879 VPWR.n5878 4.6505
R3046 VPWR.n5880 VPWR.n5858 4.6505
R3047 VPWR.n5965 VPWR.n5964 4.6505
R3048 VPWR.n5970 VPWR.n5969 4.6505
R3049 VPWR.n5977 VPWR.n5976 4.6505
R3050 VPWR.n5979 VPWR.n5978 4.6505
R3051 VPWR.n6017 VPWR.n6016 4.6505
R3052 VPWR.n6022 VPWR.n6021 4.6505
R3053 VPWR.n6024 VPWR.n6023 4.6505
R3054 VPWR.n6026 VPWR.n6025 4.6505
R3055 VPWR.n6029 VPWR.n6028 4.6505
R3056 VPWR.n6031 VPWR.n6030 4.6505
R3057 VPWR.n6033 VPWR.n6032 4.6505
R3058 VPWR.n6050 VPWR.n6049 4.6505
R3059 VPWR.n6052 VPWR.n6051 4.6505
R3060 VPWR.n6055 VPWR.n6054 4.6505
R3061 VPWR.n6057 VPWR.n6056 4.6505
R3062 VPWR.n5461 VPWR.n5460 4.6505
R3063 VPWR.n5463 VPWR.n5462 4.6505
R3064 VPWR.n5481 VPWR.n5480 4.6505
R3065 VPWR.n5484 VPWR.n5483 4.6505
R3066 VPWR.n5486 VPWR.n5485 4.6505
R3067 VPWR.n5487 VPWR.n5408 4.6505
R3068 VPWR.n5491 VPWR.n5490 4.6505
R3069 VPWR.n5518 VPWR.n5517 4.6505
R3070 VPWR.n5522 VPWR.n5521 4.6505
R3071 VPWR.n5524 VPWR.n5523 4.6505
R3072 VPWR.n5527 VPWR.n5526 4.6505
R3073 VPWR.n5528 VPWR.n5386 4.6505
R3074 VPWR.n5533 VPWR.n5532 4.6505
R3075 VPWR.n5537 VPWR.n5536 4.6505
R3076 VPWR.n5547 VPWR.n5546 4.6505
R3077 VPWR.n5549 VPWR.n5548 4.6505
R3078 VPWR.n5552 VPWR.n5551 4.6505
R3079 VPWR.n5554 VPWR.n5553 4.6505
R3080 VPWR.n5701 VPWR.n5692 4.6505
R3081 VPWR.n5698 VPWR.n5693 4.6505
R3082 VPWR.n5725 VPWR.n5690 4.6505
R3083 VPWR.n5724 VPWR.n5723 4.6505
R3084 VPWR.n5722 VPWR.n5721 4.6505
R3085 VPWR.n5719 VPWR.n5718 4.6505
R3086 VPWR.n5717 VPWR.n5716 4.6505
R3087 VPWR.n5706 VPWR.n5705 4.6505
R3088 VPWR.n5704 VPWR.n5703 4.6505
R3089 VPWR.n5702 VPWR 4.6505
R3090 VPWR.n5700 VPWR.n5699 4.6505
R3091 VPWR.n5738 VPWR.n5737 4.6505
R3092 VPWR.n5736 VPWR.n5735 4.6505
R3093 VPWR.n5733 VPWR.n5732 4.6505
R3094 VPWR.n5731 VPWR.n5730 4.6505
R3095 VPWR.n5729 VPWR.n5728 4.6505
R3096 VPWR.n5727 VPWR.n5726 4.6505
R3097 VPWR.n5545 VPWR.n5544 4.6505
R3098 VPWR.n5543 VPWR.n5542 4.6505
R3099 VPWR.n5539 VPWR.n5538 4.6505
R3100 VPWR.n5520 VPWR.n5519 4.6505
R3101 VPWR.n5516 VPWR.n5515 4.6505
R3102 VPWR.n5514 VPWR.n5513 4.6505
R3103 VPWR.n5510 VPWR.n5509 4.6505
R3104 VPWR.n5504 VPWR.n5503 4.6505
R3105 VPWR.n5502 VPWR.n5501 4.6505
R3106 VPWR.n5500 VPWR.n5499 4.6505
R3107 VPWR.n5498 VPWR.n5497 4.6505
R3108 VPWR.n5495 VPWR.n5494 4.6505
R3109 VPWR.n5489 VPWR.n5488 4.6505
R3110 VPWR.n5479 VPWR.n5478 4.6505
R3111 VPWR.n5477 VPWR.n5476 4.6505
R3112 VPWR.n5475 VPWR.n5474 4.6505
R3113 VPWR.n5471 VPWR.n5470 4.6505
R3114 VPWR.n5469 VPWR.n5468 4.6505
R3115 VPWR.n5467 VPWR.n5466 4.6505
R3116 VPWR.n6047 VPWR.n6046 4.6505
R3117 VPWR.n6045 VPWR.n6044 4.6505
R3118 VPWR.n6041 VPWR.n6040 4.6505
R3119 VPWR.n6039 VPWR.n6038 4.6505
R3120 VPWR.n6037 VPWR.n6036 4.6505
R3121 VPWR.n6035 VPWR.n6034 4.6505
R3122 VPWR.n6018 VPWR.n157 4.6505
R3123 VPWR.n6012 VPWR.n6011 4.6505
R3124 VPWR.n6007 VPWR.n6006 4.6505
R3125 VPWR.n6002 VPWR.n6001 4.6505
R3126 VPWR.n6000 VPWR.n159 4.6505
R3127 VPWR.n5999 VPWR.n5998 4.6505
R3128 VPWR.n5997 VPWR.n5996 4.6505
R3129 VPWR.n5995 VPWR.n5994 4.6505
R3130 VPWR.n5990 VPWR.n5989 4.6505
R3131 VPWR.n5988 VPWR.n5987 4.6505
R3132 VPWR.n5986 VPWR.n160 4.6505
R3133 VPWR.n5983 VPWR.n5982 4.6505
R3134 VPWR.n5871 VPWR.n5870 4.6505
R3135 VPWR VPWR.n5874 4.6505
R3136 VPWR.n5877 VPWR.n5876 4.6505
R3137 VPWR.n5883 VPWR.n5881 4.6505
R3138 VPWR.n5883 VPWR.n5882 4.6505
R3139 VPWR.n5886 VPWR.n5885 4.6505
R3140 VPWR.n5890 VPWR.n5889 4.6505
R3141 VPWR.n5899 VPWR.n5898 4.6505
R3142 VPWR.n2412 VPWR.n2411 4.6505
R3143 VPWR.n2415 VPWR.n2397 4.6505
R3144 VPWR.n2424 VPWR.n2423 4.6505
R3145 VPWR.n2427 VPWR.n2393 4.6505
R3146 VPWR.n2439 VPWR.n2438 4.6505
R3147 VPWR.n2484 VPWR.n2483 4.6505
R3148 VPWR.n2487 VPWR.n2349 4.6505
R3149 VPWR.n2522 VPWR.n2521 4.6505
R3150 VPWR.n2526 VPWR.n2525 4.6505
R3151 VPWR.n2541 VPWR.n2540 4.6505
R3152 VPWR.n2548 VPWR.n2547 4.6505
R3153 VPWR.n2563 VPWR.n2562 4.6505
R3154 VPWR.n2567 VPWR.n2566 4.6505
R3155 VPWR.n2114 VPWR.n2113 4.6505
R3156 VPWR.n2117 VPWR.n2077 4.6505
R3157 VPWR.n2128 VPWR.n2076 4.6505
R3158 VPWR.n2132 VPWR.n2131 4.6505
R3159 VPWR.n2143 VPWR.n2142 4.6505
R3160 VPWR.n2144 VPWR.n2143 4.6505
R3161 VPWR.n2148 VPWR.n2147 4.6505
R3162 VPWR.n2162 VPWR.n2161 4.6505
R3163 VPWR.n2170 VPWR.n2169 4.6505
R3164 VPWR.n2176 VPWR.n2175 4.6505
R3165 VPWR.n2184 VPWR.n2183 4.6505
R3166 VPWR.n2198 VPWR.n2197 4.6505
R3167 VPWR.n2204 VPWR.n2203 4.6505
R3168 VPWR.n2302 VPWR.n2301 4.6505
R3169 VPWR.n2298 VPWR.n2252 4.6505
R3170 VPWR.n2281 VPWR.n2260 4.6505
R3171 VPWR.n2278 VPWR.n2261 4.6505
R3172 VPWR.n2304 VPWR.n2303 4.6505
R3173 VPWR.n2300 VPWR.n2299 4.6505
R3174 VPWR VPWR.n2297 4.6505
R3175 VPWR.n2296 VPWR.n2295 4.6505
R3176 VPWR.n2292 VPWR.n2291 4.6505
R3177 VPWR.n2290 VPWR.n2289 4.6505
R3178 VPWR.n2288 VPWR.n2287 4.6505
R3179 VPWR.n2286 VPWR.n2285 4.6505
R3180 VPWR.n2284 VPWR.n2283 4.6505
R3181 VPWR.n2282 VPWR 4.6505
R3182 VPWR.n2280 VPWR.n2279 4.6505
R3183 VPWR.n2277 VPWR.n2276 4.6505
R3184 VPWR.n2275 VPWR.n2274 4.6505
R3185 VPWR.n2273 VPWR.n2272 4.6505
R3186 VPWR.n2271 VPWR.n2270 4.6505
R3187 VPWR.n2269 VPWR.n2268 4.6505
R3188 VPWR.n2267 VPWR.n2266 4.6505
R3189 VPWR.n2265 VPWR.n2264 4.6505
R3190 VPWR.n2306 VPWR.n2305 4.6505
R3191 VPWR.n2112 VPWR.n2111 4.6505
R3192 VPWR.n2116 VPWR.n2115 4.6505
R3193 VPWR.n2118 VPWR 4.6505
R3194 VPWR.n2123 VPWR.n2122 4.6505
R3195 VPWR.n2127 VPWR.n2126 4.6505
R3196 VPWR.n2130 VPWR.n2129 4.6505
R3197 VPWR.n2135 VPWR.n2134 4.6505
R3198 VPWR.n2137 VPWR.n2136 4.6505
R3199 VPWR.n2139 VPWR.n2138 4.6505
R3200 VPWR.n2141 VPWR.n2140 4.6505
R3201 VPWR.n2146 VPWR.n2145 4.6505
R3202 VPWR.n2150 VPWR.n2149 4.6505
R3203 VPWR.n2152 VPWR.n2151 4.6505
R3204 VPWR.n2159 VPWR.n2158 4.6505
R3205 VPWR.n2160 VPWR.n2068 4.6505
R3206 VPWR.n2166 VPWR.n2165 4.6505
R3207 VPWR.n2168 VPWR.n2167 4.6505
R3208 VPWR.n2172 VPWR.n2171 4.6505
R3209 VPWR.n2174 VPWR.n2173 4.6505
R3210 VPWR.n2178 VPWR.n2177 4.6505
R3211 VPWR.n2180 VPWR.n2179 4.6505
R3212 VPWR.n2182 VPWR.n2181 4.6505
R3213 VPWR.n2186 VPWR.n2185 4.6505
R3214 VPWR.n2188 VPWR.n2187 4.6505
R3215 VPWR.n2190 VPWR.n2189 4.6505
R3216 VPWR.n2192 VPWR.n2191 4.6505
R3217 VPWR.n2194 VPWR.n2193 4.6505
R3218 VPWR.n2196 VPWR.n2195 4.6505
R3219 VPWR.n2200 VPWR.n2199 4.6505
R3220 VPWR.n2202 VPWR.n2201 4.6505
R3221 VPWR.n2206 VPWR.n2205 4.6505
R3222 VPWR.n2208 VPWR.n2207 4.6505
R3223 VPWR.n2211 VPWR.n2072 4.6505
R3224 VPWR.n2482 VPWR.n2481 4.6505
R3225 VPWR.n2486 VPWR.n2485 4.6505
R3226 VPWR.n2488 VPWR 4.6505
R3227 VPWR.n2496 VPWR.n2495 4.6505
R3228 VPWR.n2500 VPWR.n2499 4.6505
R3229 VPWR.n2504 VPWR.n2503 4.6505
R3230 VPWR.n2508 VPWR.n2507 4.6505
R3231 VPWR.n2510 VPWR.n2509 4.6505
R3232 VPWR.n2512 VPWR.n2511 4.6505
R3233 VPWR.n2514 VPWR.n2513 4.6505
R3234 VPWR.n2516 VPWR.n2515 4.6505
R3235 VPWR.n2518 VPWR.n2517 4.6505
R3236 VPWR.n2519 VPWR.n2348 4.6505
R3237 VPWR.n2520 VPWR 4.6505
R3238 VPWR.n2524 VPWR.n2523 4.6505
R3239 VPWR.n2529 VPWR.n2528 4.6505
R3240 VPWR.n2531 VPWR.n2530 4.6505
R3241 VPWR.n2533 VPWR.n2532 4.6505
R3242 VPWR.n2534 VPWR.n2346 4.6505
R3243 VPWR.n2536 VPWR.n2535 4.6505
R3244 VPWR.n2544 VPWR.n2345 4.6505
R3245 VPWR.n2546 VPWR.n2545 4.6505
R3246 VPWR.n2550 VPWR.n2549 4.6505
R3247 VPWR.n2552 VPWR.n2551 4.6505
R3248 VPWR.n2555 VPWR.n2344 4.6505
R3249 VPWR.n2557 VPWR.n2556 4.6505
R3250 VPWR.n2559 VPWR.n2558 4.6505
R3251 VPWR.n2561 VPWR.n2560 4.6505
R3252 VPWR.n2565 VPWR.n2564 4.6505
R3253 VPWR.n2569 VPWR.n2568 4.6505
R3254 VPWR.n2571 VPWR.n2570 4.6505
R3255 VPWR.n2573 VPWR.n2572 4.6505
R3256 VPWR.n2575 VPWR.n2574 4.6505
R3257 VPWR.n2578 VPWR.n2577 4.6505
R3258 VPWR.n2583 VPWR.n2582 4.6505
R3259 VPWR.n2586 VPWR.n2585 4.6505
R3260 VPWR.n2588 VPWR.n2587 4.6505
R3261 VPWR.n2591 VPWR.n2067 4.6505
R3262 VPWR.n2593 VPWR.n2592 4.6505
R3263 VPWR.n2404 VPWR.n2403 4.6505
R3264 VPWR.n2406 VPWR.n2405 4.6505
R3265 VPWR.n2410 VPWR.n2409 4.6505
R3266 VPWR.n2414 VPWR.n2413 4.6505
R3267 VPWR.n2416 VPWR 4.6505
R3268 VPWR.n2418 VPWR.n2417 4.6505
R3269 VPWR.n2422 VPWR.n2421 4.6505
R3270 VPWR.n2426 VPWR.n2425 4.6505
R3271 VPWR.n2428 VPWR 4.6505
R3272 VPWR.n2430 VPWR.n2429 4.6505
R3273 VPWR.n2432 VPWR.n2431 4.6505
R3274 VPWR.n2434 VPWR.n2433 4.6505
R3275 VPWR.n2437 VPWR.n2391 4.6505
R3276 VPWR.n6095 VPWR 4.6505
R3277 VPWR.n6104 VPWR.n6103 4.6505
R3278 VPWR.n6104 VPWR.n90 4.6505
R3279 VPWR.n6168 VPWR.n6167 4.6505
R3280 VPWR.n6241 VPWR.n47 4.6505
R3281 VPWR.n6240 VPWR.n49 4.6505
R3282 VPWR.n6227 VPWR.n61 4.6505
R3283 VPWR.n6215 VPWR.n67 4.6505
R3284 VPWR.n6208 VPWR.n68 4.6505
R3285 VPWR.n6207 VPWR.n69 4.6505
R3286 VPWR.n5 VPWR.n4 4.6505
R3287 VPWR.n9 VPWR.n8 4.6505
R3288 VPWR.n6257 VPWR.n6256 4.6505
R3289 VPWR.n6253 VPWR 4.6505
R3290 VPWR.n6252 VPWR.n41 4.6505
R3291 VPWR.n6248 VPWR.n6247 4.6505
R3292 VPWR.n6246 VPWR.n6245 4.6505
R3293 VPWR.n6244 VPWR.n6243 4.6505
R3294 VPWR.n6242 VPWR 4.6505
R3295 VPWR.n6218 VPWR.n66 4.6505
R3296 VPWR.n6199 VPWR.n6198 4.6505
R3297 VPWR.n6087 VPWR.n6086 4.6505
R3298 VPWR.n6089 VPWR.n6088 4.6505
R3299 VPWR.n6091 VPWR.n6090 4.6505
R3300 VPWR.n6093 VPWR.n6092 4.6505
R3301 VPWR.n6138 VPWR.n6137 4.6505
R3302 VPWR.n6141 VPWR.n87 4.6505
R3303 VPWR.n6142 VPWR 4.6505
R3304 VPWR.n6146 VPWR.n6145 4.6505
R3305 VPWR VPWR.n6153 4.6505
R3306 VPWR.n6157 VPWR.n6156 4.6505
R3307 VPWR.n6170 VPWR.n6169 4.6505
R3308 VPWR.n6172 VPWR.n6171 4.6505
R3309 VPWR.n6174 VPWR.n6173 4.6505
R3310 VPWR.n6177 VPWR.n78 4.6505
R3311 VPWR VPWR.n82 4.6505
R3312 VPWR.n6166 VPWR.n6165 4.6505
R3313 VPWR.n6159 VPWR.n6158 4.6505
R3314 VPWR.n6150 VPWR.n6149 4.6505
R3315 VPWR.n6133 VPWR.n6132 4.6505
R3316 VPWR.n6128 VPWR.n74 4.6505
R3317 VPWR.n6127 VPWR.n6126 4.6505
R3318 VPWR.n6123 VPWR.n6122 4.6505
R3319 VPWR.n6118 VPWR.n6117 4.6505
R3320 VPWR.n6116 VPWR.n6115 4.6505
R3321 VPWR.n6114 VPWR.n6113 4.6505
R3322 VPWR.n6112 VPWR.n6111 4.6505
R3323 VPWR.n6110 VPWR.n6109 4.6505
R3324 VPWR.n6108 VPWR.n6107 4.6505
R3325 VPWR.n6202 VPWR.n6201 4.6505
R3326 VPWR.n6206 VPWR.n6205 4.6505
R3327 VPWR.n6210 VPWR.n6209 4.6505
R3328 VPWR.n6212 VPWR.n6211 4.6505
R3329 VPWR.n6217 VPWR.n6216 4.6505
R3330 VPWR.n6219 VPWR 4.6505
R3331 VPWR.n6221 VPWR.n6220 4.6505
R3332 VPWR.n6225 VPWR.n6224 4.6505
R3333 VPWR.n6229 VPWR.n6228 4.6505
R3334 VPWR.n6231 VPWR.n6230 4.6505
R3335 VPWR.n6233 VPWR.n6232 4.6505
R3336 VPWR.n6235 VPWR.n6234 4.6505
R3337 VPWR.n6238 VPWR.n6237 4.6505
R3338 VPWR.n7 VPWR.n6 4.6505
R3339 VPWR VPWR.n6306 4.6505
R3340 VPWR.n6304 VPWR.n6303 4.6505
R3341 VPWR VPWR.n6300 4.6505
R3342 VPWR.n6292 VPWR.n6291 4.6505
R3343 VPWR.n6290 VPWR.n6289 4.6505
R3344 VPWR.n5638 VPWR.n5637 4.6505
R3345 VPWR.n5631 VPWR.n5630 4.6505
R3346 VPWR.n5629 VPWR 4.6505
R3347 VPWR.n5628 VPWR.n5627 4.6505
R3348 VPWR.n5626 VPWR.n5625 4.6505
R3349 VPWR.n5624 VPWR.n5593 4.6505
R3350 VPWR.n5623 VPWR.n5622 4.6505
R3351 VPWR.n5620 VPWR.n5619 4.6505
R3352 VPWR.n5618 VPWR.n5617 4.6505
R3353 VPWR.n5616 VPWR.n5615 4.6505
R3354 VPWR.n5614 VPWR 4.6505
R3355 VPWR.n5613 VPWR.n5594 4.6505
R3356 VPWR.n5612 VPWR.n5611 4.6505
R3357 VPWR.n5610 VPWR.n5609 4.6505
R3358 VPWR.n5608 VPWR.n5607 4.6505
R3359 VPWR.n5606 VPWR.n5605 4.6505
R3360 VPWR.n5604 VPWR.n5603 4.6505
R3361 VPWR.n5602 VPWR.n5601 4.6505
R3362 VPWR.n5600 VPWR.n5599 4.6505
R3363 VPWR.n3090 VPWR.n3089 4.64677
R3364 VPWR.n3032 VPWR.n3031 4.64677
R3365 VPWR.n5272 VPWR.n5271 4.64677
R3366 VPWR.n5786 VPWR.n5785 4.64677
R3367 VPWR.n2337 VPWR.n2336 4.64677
R3368 VPWR.n3441 VPWR.n3440 4.64677
R3369 VPWR.n1294 VPWR.n1293 4.64677
R3370 VPWR.n4087 VPWR.n4086 4.64677
R3371 VPWR.n6192 VPWR.n6191 4.64677
R3372 VPWR.n764 VPWR.n763 4.64226
R3373 VPWR.n6145 VPWR.n6142 4.59011
R3374 VPWR.n1634 VPWR.n1633 4.59011
R3375 VPWR.n4065 VPWR.n4064 4.59011
R3376 VPWR.n3942 VPWR.n3941 4.59011
R3377 VPWR.n921 VPWR.n814 4.59011
R3378 VPWR.n5123 VPWR.n5107 4.59011
R3379 VPWR.n5176 VPWR.n316 4.59011
R3380 VPWR.n1610 VPWR.n1609 4.57427
R3381 VPWR.n2625 VPWR.n2624 4.57427
R3382 VPWR.n3097 VPWR.n3096 4.57427
R3383 VPWR.n1692 VPWR.n1691 4.57427
R3384 VPWR.n1910 VPWR.n1909 4.57427
R3385 VPWR.n1330 VPWR.n1329 4.57427
R3386 VPWR.n3294 VPWR.n3293 4.57427
R3387 VPWR.n3760 VPWR.n1190 4.57427
R3388 VPWR.n3474 VPWR.n3473 4.57427
R3389 VPWR.n993 VPWR.n992 4.57427
R3390 VPWR.n3859 VPWR.n3858 4.57427
R3391 VPWR.n4147 VPWR.n4146 4.57427
R3392 VPWR.n4364 VPWR.n4363 4.57427
R3393 VPWR.n4895 VPWR.n4447 4.57427
R3394 VPWR.n4515 VPWR.n4514 4.57427
R3395 VPWR.n4599 VPWR.n4598 4.57427
R3396 VPWR.n260 VPWR.n259 4.57427
R3397 VPWR.n5324 VPWR.n5323 4.57427
R3398 VPWR.n340 VPWR.n339 4.57427
R3399 VPWR.n5793 VPWR.n5792 4.57427
R3400 VPWR.n5410 VPWR.n5409 4.57427
R3401 VPWR.n5689 VPWR.n5688 4.57427
R3402 VPWR.n5934 VPWR.n5933 4.57427
R3403 VPWR.n2086 VPWR.n2085 4.57427
R3404 VPWR.n2454 VPWR.n2453 4.57427
R3405 VPWR.n2251 VPWR.n2250 4.57427
R3406 VPWR.n96 VPWR.n95 4.57427
R3407 VPWR.n2112 VPWR.n2078 4.52113
R3408 VPWR.n4714 VPWR.n4713 4.52113
R3409 VPWR.n5162 VPWR.n5161 4.52113
R3410 VPWR.n5430 VPWR.n5429 4.5005
R3411 VPWR.n5173 VPWR.n317 4.47674
R3412 VPWR.n1859 VPWR.n1858 4.47426
R3413 VPWR.n4146 VPWR.n4143 4.41955
R3414 VPWR.n4514 VPWR.n4512 4.41955
R3415 VPWR.n259 VPWR.n257 4.41955
R3416 VPWR.n2482 VPWR.n2350 4.21637
R3417 VPWR.n1820 VPWR.n1818 4.1826
R3418 VPWR.n503 VPWR.n502 4.17775
R3419 VPWR.n1818 VPWR.n1817 4.17318
R3420 VPWR.n1411 VPWR.n1410 4.17318
R3421 VPWR.n3161 VPWR.n3160 4.17318
R3422 VPWR.n1253 VPWR.n1252 4.17318
R3423 VPWR.n1212 VPWR.n1211 4.17318
R3424 VPWR.n6104 VPWR.n89 4.12386
R3425 VPWR.n63 VPWR.n62 4.12386
R3426 VPWR.n1414 VPWR.n1413 4.12386
R3427 VPWR.n1271 VPWR.n1270 4.12386
R3428 VPWR.n3602 VPWR.n3601 4.12386
R3429 VPWR.n3990 VPWR.n3989 4.12386
R3430 VPWR.n3911 VPWR.n1128 4.12386
R3431 VPWR.n709 VPWR.n708 4.12386
R3432 VPWR.n4407 VPWR.n4406 4.12386
R3433 VPWR.n4584 VPWR.n4583 4.12386
R3434 VPWR.n4773 VPWR.n4588 4.12386
R3435 VPWR.n4656 VPWR.n4655 4.12386
R3436 VPWR.n4830 VPWR.n4473 4.12386
R3437 VPWR.n277 VPWR.n276 4.12386
R3438 VPWR.n501 VPWR.n500 4.12386
R3439 VPWR.n5873 VPWR.n5872 4.12386
R3440 VPWR.n5407 VPWR.n5406 4.12386
R3441 VPWR.n5531 VPWR.n5530 4.12386
R3442 VPWR.n5634 VPWR.n5592 4.12386
R3443 VPWR.n1884 VPWR.n1883 4.06399
R3444 VPWR.n742 VPWR.n741 4.06399
R3445 VPWR.n4440 VPWR.n4439 4.06399
R3446 VPWR.n1562 VPWR.n1561 4.06399
R3447 VPWR.n3194 VPWR.n3193 4.06399
R3448 VPWR.n1183 VPWR.n1182 4.06399
R3449 VPWR.n4987 VPWR.n4986 4.06399
R3450 VPWR.n6291 VPWR.n6290 3.99029
R3451 VPWR.n185 VPWR.n184 3.98162
R3452 VPWR VPWR.n881 3.81002
R3453 VPWR.n5099 VPWR 3.81002
R3454 VPWR VPWR.n388 3.81002
R3455 VPWR.n3000 VPWR.n2997 3.54454
R3456 VPWR.n2756 VPWR.n2755 3.4105
R3457 VPWR.n1663 VPWR.n1662 3.4105
R3458 VPWR.n1593 VPWR.n1592 3.4105
R3459 VPWR.n3078 VPWR.n3077 3.4105
R3460 VPWR.n3085 VPWR.n3084 3.4105
R3461 VPWR.n2740 VPWR.n2739 3.4105
R3462 VPWR.n2748 VPWR.n2747 3.4105
R3463 VPWR.n2911 VPWR.n2910 3.4105
R3464 VPWR.n3114 VPWR.n3113 3.4105
R3465 VPWR.n3108 VPWR.n3107 3.4105
R3466 VPWR.n2808 VPWR.n2807 3.4105
R3467 VPWR.n1806 VPWR.n1805 3.4105
R3468 VPWR.n1747 VPWR.n1746 3.4105
R3469 VPWR.n1675 VPWR.n1674 3.4105
R3470 VPWR.n1763 VPWR.n1762 3.4105
R3471 VPWR.n3037 VPWR.n3036 3.4105
R3472 VPWR.n2935 VPWR.n2934 3.4105
R3473 VPWR.n1798 VPWR.n1797 3.4105
R3474 VPWR.n2034 VPWR.n2033 3.4105
R3475 VPWR.n1895 VPWR.n1894 3.4105
R3476 VPWR.n1906 VPWR.n1905 3.4105
R3477 VPWR.n1918 VPWR.n1917 3.4105
R3478 VPWR.n1930 VPWR.n1929 3.4105
R3479 VPWR.n1402 VPWR.n1401 3.4105
R3480 VPWR.n3345 VPWR.n3344 3.4105
R3481 VPWR.n1387 VPWR.n1386 3.4105
R3482 VPWR.n1378 VPWR.n1377 3.4105
R3483 VPWR.n1473 VPWR.n1472 3.4105
R3484 VPWR.n1465 VPWR.n1464 3.4105
R3485 VPWR.n3353 VPWR.n3352 3.4105
R3486 VPWR.n3446 VPWR.n3445 3.4105
R3487 VPWR.n3216 VPWR.n3215 3.4105
R3488 VPWR.n3210 VPWR.n3209 3.4105
R3489 VPWR.n3286 VPWR.n3285 3.4105
R3490 VPWR.n3277 VPWR.n3276 3.4105
R3491 VPWR.n3546 VPWR.n3545 3.4105
R3492 VPWR.n3654 VPWR.n3653 3.4105
R3493 VPWR.n3537 VPWR.n3536 3.4105
R3494 VPWR.n3528 VPWR.n3527 3.4105
R3495 VPWR.n3647 VPWR.n3646 3.4105
R3496 VPWR.n3639 VPWR.n3638 3.4105
R3497 VPWR.n3631 VPWR.n3630 3.4105
R3498 VPWR.n3553 VPWR.n3552 3.4105
R3499 VPWR.n3777 VPWR.n3776 3.4105
R3500 VPWR.n3771 VPWR.n3770 3.4105
R3501 VPWR.n3753 VPWR.n3752 3.4105
R3502 VPWR.n3744 VPWR.n3743 3.4105
R3503 VPWR.n1062 VPWR.n1061 3.4105
R3504 VPWR.n3979 VPWR.n3978 3.4105
R3505 VPWR.n976 VPWR.n975 3.4105
R3506 VPWR.n1042 VPWR.n1041 3.4105
R3507 VPWR.n1112 VPWR.n1111 3.4105
R3508 VPWR.n1104 VPWR.n1103 3.4105
R3509 VPWR.n3987 VPWR.n3986 3.4105
R3510 VPWR.n4092 VPWR.n4091 3.4105
R3511 VPWR.n3876 VPWR.n3875 3.4105
R3512 VPWR.n3870 VPWR.n3869 3.4105
R3513 VPWR.n3851 VPWR.n3850 3.4105
R3514 VPWR.n3884 VPWR.n3883 3.4105
R3515 VPWR.n4230 VPWR.n4229 3.4105
R3516 VPWR.n797 VPWR.n796 3.4105
R3517 VPWR.n4130 VPWR.n4129 3.4105
R3518 VPWR.n4350 VPWR.n4349 3.4105
R3519 VPWR.n953 VPWR.n952 3.4105
R3520 VPWR.n4202 VPWR.n4201 3.4105
R3521 VPWR.n805 VPWR.n804 3.4105
R3522 VPWR.n4341 VPWR.n4340 3.4105
R3523 VPWR.n4381 VPWR.n4380 3.4105
R3524 VPWR.n4375 VPWR.n4374 3.4105
R3525 VPWR.n845 VPWR.n844 3.4105
R3526 VPWR.n858 VPWR.n857 3.4105
R3527 VPWR.n4643 VPWR.n4642 3.4105
R3528 VPWR.n4565 VPWR.n4564 3.4105
R3529 VPWR.n4498 VPWR.n4497 3.4105
R3530 VPWR.n4817 VPWR.n4816 3.4105
R3531 VPWR.n4808 VPWR.n4807 3.4105
R3532 VPWR.n4635 VPWR.n4634 3.4105
R3533 VPWR.n4709 VPWR.n4708 3.4105
R3534 VPWR.n4703 VPWR.n4702 3.4105
R3535 VPWR.n4912 VPWR.n4911 3.4105
R3536 VPWR.n4906 VPWR.n4905 3.4105
R3537 VPWR.n4889 VPWR.n4888 3.4105
R3538 VPWR.n4880 VPWR.n4879 3.4105
R3539 VPWR.n657 VPWR.n656 3.4105
R3540 VPWR.n295 VPWR.n294 3.4105
R3541 VPWR.n244 VPWR.n243 3.4105
R3542 VPWR.n310 VPWR.n309 3.4105
R3543 VPWR.n5277 VPWR.n5276 3.4105
R3544 VPWR.n673 VPWR.n672 3.4105
R3545 VPWR.n5157 VPWR.n5156 3.4105
R3546 VPWR.n5151 VPWR.n5150 3.4105
R3547 VPWR.n5034 VPWR.n5033 3.4105
R3548 VPWR.n5028 VPWR.n5027 3.4105
R3549 VPWR.n5011 VPWR.n5010 3.4105
R3550 VPWR.n5042 VPWR.n5041 3.4105
R3551 VPWR.n482 VPWR.n481 3.4105
R3552 VPWR.n5376 VPWR.n5375 3.4105
R3553 VPWR.n5307 VPWR.n5306 3.4105
R3554 VPWR.n5774 VPWR.n5773 3.4105
R3555 VPWR.n5781 VPWR.n5780 3.4105
R3556 VPWR.n466 VPWR.n465 3.4105
R3557 VPWR.n474 VPWR.n473 3.4105
R3558 VPWR.n621 VPWR.n620 3.4105
R3559 VPWR.n5810 VPWR.n5809 3.4105
R3560 VPWR.n5804 VPWR.n5803 3.4105
R3561 VPWR.n518 VPWR.n517 3.4105
R3562 VPWR.n532 VPWR.n531 3.4105
R3563 VPWR.n5559 VPWR.n5558 3.4105
R3564 VPWR.n5742 VPWR.n5741 3.4105
R3565 VPWR.n5683 VPWR.n5682 3.4105
R3566 VPWR.n5398 VPWR.n5397 3.4105
R3567 VPWR.n6063 VPWR.n6062 3.4105
R3568 VPWR.n5437 VPWR.n5436 3.4105
R3569 VPWR.n5452 VPWR.n5451 3.4105
R3570 VPWR.n5951 VPWR.n5950 3.4105
R3571 VPWR.n5945 VPWR.n5944 3.4105
R3572 VPWR.n5918 VPWR.n5917 3.4105
R3573 VPWR.n5959 VPWR.n5958 3.4105
R3574 VPWR.n2107 VPWR.n2106 3.4105
R3575 VPWR.n2098 VPWR.n2097 3.4105
R3576 VPWR.n2599 VPWR.n2598 3.4105
R3577 VPWR.n2480 VPWR.n2479 3.4105
R3578 VPWR.n2462 VPWR.n2461 3.4105
R3579 VPWR.n2325 VPWR.n2324 3.4105
R3580 VPWR.n2309 VPWR.n2308 3.4105
R3581 VPWR.n2234 VPWR.n2233 3.4105
R3582 VPWR.n2332 VPWR.n2331 3.4105
R3583 VPWR.n6182 VPWR.n6181 3.4105
R3584 VPWR.n6286 VPWR.n6285 3.4105
R3585 VPWR.n6278 VPWR.n6277 3.4105
R3586 VPWR.n6269 VPWR.n6268 3.4105
R3587 VPWR.n6260 VPWR.n6259 3.4105
R3588 VPWR.n6190 VPWR.n6189 3.4105
R3589 VPWR.n5579 VPWR.n5578 3.4105
R3590 VPWR.n5641 VPWR.n5640 3.4105
R3591 VPWR.n147 VPWR.n146 3.4105
R3592 VPWR.n136 VPWR.n135 3.4105
R3593 VPWR.n128 VPWR.n127 3.4105
R3594 VPWR.n6080 VPWR.n6079 3.4105
R3595 VPWR VPWR 3.35739
R3596 VPWR VPWR 3.35739
R3597 VPWR VPWR 3.35739
R3598 VPWR VPWR 3.35739
R3599 VPWR VPWR 3.35739
R3600 VPWR VPWR 3.35739
R3601 VPWR VPWR 3.35739
R3602 VPWR.n2735 VPWR.n2635 3.31258
R3603 VPWR.n4799 VPWR.n4796 3.31258
R3604 VPWR.n13 VPWR.n12 3.30837
R3605 VPWR.n2493 VPWR.n2492 3.30837
R3606 VPWR.n1524 VPWR 3.29747
R3607 VPWR.n4469 VPWR 3.29747
R3608 VPWR.n4873 VPWR 3.29747
R3609 VPWR.n2653 VPWR.n2652 3.28365
R3610 VPWR.n5101 VPWR.n5100 3.27868
R3611 VPWR.n2665 VPWR.n2653 3.273
R3612 VPWR.n5102 VPWR.n5101 3.273
R3613 VPWR.n198 VPWR 3.24826
R3614 VPWR.n2734 VPWR.n2636 3.23
R3615 VPWR.n4798 VPWR.n4797 3.23
R3616 VPWR.n3324 VPWR.n3323 3.21792
R3617 VPWR.n3303 VPWR.n1493 3.21792
R3618 VPWR.n4659 VPWR.n4658 3.20752
R3619 VPWR.n4954 VPWR.n4953 3.20752
R3620 VPWR.n490 VPWR.n489 3.20752
R3621 VPWR.n1951 VPWR.n1817 3.20443
R3622 VPWR.n5131 VPWR.n5102 3.20311
R3623 VPWR.n2734 VPWR.n2733 3.2005
R3624 VPWR.n3340 VPWR.n3339 3.2005
R3625 VPWR.n3911 VPWR.n1126 3.2005
R3626 VPWR.n4773 VPWR.n4772 3.2005
R3627 VPWR.n5872 VPWR.n5871 3.2005
R3628 VPWR.n2254 VPWR.n2253 3.16454
R3629 VPWR.n216 VPWR.n215 3.11611
R3630 VPWR.n2084 VPWR.n2083 3.09891
R3631 VPWR.n2452 VPWR.n2451 3.09891
R3632 VPWR.n4597 VPWR.n4596 3.09891
R3633 VPWR.n5147 VPWR.n5146 3.06214
R3634 VPWR.n617 VPWR.n226 3.06214
R3635 VPWR.n1265 VPWR.n1264 3.06214
R3636 VPWR.n3975 VPWR.n3974 3.06214
R3637 VPWR.n949 VPWR.n751 3.06214
R3638 VPWR.n6288 VPWR.n25 3.06214
R3639 VPWR.n2030 VPWR.n2028 3.06213
R3640 VPWR.n3341 VPWR.n3340 3.06213
R3641 VPWR.n143 VPWR.n73 3.06213
R3642 VPWR.n2737 VPWR.n2634 3.0621
R3643 VPWR.n772 VPWR.n771 3.06205
R3644 VPWR.n89 VPWR.n88 3.00117
R3645 VPWR.n3809 VPWR.n3808 3.00117
R3646 VPWR.n710 VPWR.n709 3.00117
R3647 VPWR.n4408 VPWR.n4407 3.00117
R3648 VPWR.n4790 VPWR.n4583 3.00117
R3649 VPWR.n4588 VPWR.n4587 3.00117
R3650 VPWR.n544 VPWR.n500 3.00117
R3651 VPWR.n187 VPWR.n186 3.00117
R3652 VPWR.n5874 VPWR.n5873 3.00117
R3653 VPWR.n5532 VPWR.n5531 3.00117
R3654 VPWR.n5637 VPWR.n5634 3.00117
R3655 VPWR.n6300 VPWR.n16 2.80499
R3656 VPWR.n2258 VPWR.n2257 2.76904
R3657 VPWR.n216 VPWR.n185 2.69753
R3658 VPWR.n170 VPWR.n162 2.68875
R3659 VPWR.n169 VPWR.n167 2.68875
R3660 VPWR.n162 VPWR.n161 2.68714
R3661 VPWR.n2906 VPWR.n2905 2.598
R3662 VPWR.n1372 VPWR.n1371 2.59206
R3663 VPWR.n6304 VPWR.n11 2.51735
R3664 VPWR.n2495 VPWR.n2494 2.51735
R3665 VPWR.n44 VPWR.n43 2.50603
R3666 VPWR.n22 VPWR.n21 2.50603
R3667 VPWR.n21 VPWR.n20 2.50603
R3668 VPWR.n20 VPWR.n19 2.50603
R3669 VPWR.n1842 VPWR.n1841 2.50603
R3670 VPWR.n1843 VPWR.n1842 2.50603
R3671 VPWR.n1866 VPWR.n1843 2.50603
R3672 VPWR.n5896 VPWR.n5895 2.50603
R3673 VPWR.n5897 VPWR.n5896 2.50603
R3674 VPWR.n5898 VPWR.n5897 2.50603
R3675 VPWR.n5714 VPWR.n5713 2.50603
R3676 VPWR.n5713 VPWR.n5712 2.50603
R3677 VPWR.n4241 VPWR.n4240 2.4386
R3678 VPWR.n874 VPWR.n873 2.4386
R3679 VPWR.n5047 VPWR.n5046 2.4386
R3680 VPWR.n4980 VPWR.n4979 2.4386
R3681 VPWR.n578 VPWR.n577 2.4386
R3682 VPWR.n3807 VPWR.n3806 2.37764
R3683 VPWR.n2296 VPWR.n2259 2.37353
R3684 VPWR.n6099 VPWR.n6098 2.33701
R3685 VPWR.n6121 VPWR.n6120 2.33701
R3686 VPWR.n6098 VPWR.n6097 2.33701
R3687 VPWR.n6131 VPWR.n6130 2.33701
R3688 VPWR.n87 VPWR.n86 2.33701
R3689 VPWR.n6144 VPWR.n6143 2.33701
R3690 VPWR.n6152 VPWR.n6151 2.33701
R3691 VPWR.n6163 VPWR.n6162 2.33701
R3692 VPWR.n76 VPWR.n75 2.33701
R3693 VPWR.n77 VPWR.n76 2.33701
R3694 VPWR.n2250 VPWR.n2248 2.33701
R3695 VPWR.n2070 VPWR.n2069 2.33701
R3696 VPWR.n2074 VPWR.n2073 2.33701
R3697 VPWR.n2156 VPWR.n2155 2.33701
R3698 VPWR.n2121 VPWR.n2120 2.33701
R3699 VPWR.n2085 VPWR.n2081 2.33701
R3700 VPWR.n2342 VPWR.n2341 2.33701
R3701 VPWR.n2539 VPWR.n2538 2.33701
R3702 VPWR.n2399 VPWR.n2398 2.33701
R3703 VPWR.n2395 VPWR.n2394 2.33701
R3704 VPWR.n2453 VPWR.n2448 2.33701
R3705 VPWR.n1630 VPWR.n1620 2.33701
R3706 VPWR.n1635 VPWR.n1619 2.33701
R3707 VPWR.n1641 VPWR.n1616 2.33701
R3708 VPWR.n1609 VPWR.n1607 2.33701
R3709 VPWR.n1574 VPWR.n1573 2.33701
R3710 VPWR.n2648 VPWR.n2647 2.33701
R3711 VPWR.n2770 VPWR.n2769 2.33701
R3712 VPWR.n1540 VPWR.n1523 2.33701
R3713 VPWR.n1700 VPWR.n1699 2.33701
R3714 VPWR.n1699 VPWR.n1698 2.33701
R3715 VPWR.n1767 VPWR.n1766 2.33701
R3716 VPWR.n2984 VPWR.n2983 2.33701
R3717 VPWR.n2958 VPWR.n1771 2.33701
R3718 VPWR.n2951 VPWR.n1772 2.33701
R3719 VPWR.n2943 VPWR.n2942 2.33701
R3720 VPWR.n1881 VPWR.n1880 2.33701
R3721 VPWR.n1933 VPWR.n1932 2.33701
R3722 VPWR.n3421 VPWR.n3420 2.33701
R3723 VPWR.n1349 VPWR.n1333 2.33701
R3724 VPWR.n1329 VPWR.n1327 2.33701
R3725 VPWR.n1490 VPWR.n1489 2.33701
R3726 VPWR.n3170 VPWR.n3169 2.33701
R3727 VPWR.n3191 VPWR.n3190 2.33701
R3728 VPWR.n3274 VPWR.n3273 2.33701
R3729 VPWR.n1277 VPWR.n1276 2.33701
R3730 VPWR.n3488 VPWR.n3481 2.33701
R3731 VPWR.n3502 VPWR.n3476 2.33701
R3732 VPWR.n3499 VPWR.n3476 2.33701
R3733 VPWR.n3741 VPWR.n3740 2.33701
R3734 VPWR.n1147 VPWR.n1146 2.33701
R3735 VPWR.n1259 VPWR.n1258 2.33701
R3736 VPWR.n1227 VPWR.n1226 2.33701
R3737 VPWR.n1215 VPWR.n1214 2.33701
R3738 VPWR.n3705 VPWR.n1217 2.33701
R3739 VPWR.n999 VPWR.n998 2.33701
R3740 VPWR.n996 VPWR.n995 2.33701
R3741 VPWR.n1064 VPWR.n1063 2.33701
R3742 VPWR.n1065 VPWR.n1064 2.33701
R3743 VPWR.n4039 VPWR.n4038 2.33701
R3744 VPWR.n4037 VPWR.n4036 2.33701
R3745 VPWR.n4082 VPWR.n4081 2.33701
R3746 VPWR.n3938 VPWR.n3930 2.33701
R3747 VPWR.n3929 VPWR.n3928 2.33701
R3748 VPWR.n3924 VPWR.n3923 2.33701
R3749 VPWR.n3905 VPWR.n3904 2.33701
R3750 VPWR.n4189 VPWR.n4188 2.33701
R3751 VPWR.n944 VPWR.n943 2.33701
R3752 VPWR.n917 VPWR.n916 2.33701
R3753 VPWR.n817 VPWR.n816 2.33701
R3754 VPWR.n876 VPWR.n875 2.33701
R3755 VPWR.n875 VPWR.n823 2.33701
R3756 VPWR.n861 VPWR.n860 2.33701
R3757 VPWR.n4245 VPWR.n4244 2.33701
R3758 VPWR.n4244 VPWR.n4243 2.33701
R3759 VPWR.n4286 VPWR.n4285 2.33701
R3760 VPWR.n762 VPWR.n761 2.33701
R3761 VPWR.n759 VPWR.n758 2.33701
R3762 VPWR.n4333 VPWR.n4332 2.33701
R3763 VPWR.n4868 VPWR.n4867 2.33701
R3764 VPWR.n4551 VPWR.n4550 2.33701
R3765 VPWR.n4771 VPWR.n4589 2.33701
R3766 VPWR.n4729 VPWR.n4728 2.33701
R3767 VPWR.n4598 VPWR.n4593 2.33701
R3768 VPWR.n4468 VPWR.n4467 2.33701
R3769 VPWR.n312 VPWR.n311 2.33701
R3770 VPWR.n5222 VPWR.n5221 2.33701
R3771 VPWR.n5223 VPWR.n5222 2.33701
R3772 VPWR.n4961 VPWR.n4960 2.33701
R3773 VPWR.n5122 VPWR.n5121 2.33701
R3774 VPWR.n5106 VPWR.n5105 2.33701
R3775 VPWR.n5098 VPWR.n5097 2.33701
R3776 VPWR.n5053 VPWR.n5052 2.33701
R3777 VPWR.n4987 VPWR.n4985 2.33701
R3778 VPWR.n5215 VPWR.n5214 2.33701
R3779 VPWR.n5175 VPWR.n5174 2.33701
R3780 VPWR.n5207 VPWR.n5206 2.33701
R3781 VPWR.n5345 VPWR.n5344 2.33701
R3782 VPWR.n562 VPWR.n498 2.33701
R3783 VPWR.n494 VPWR.n493 2.33701
R3784 VPWR.n495 VPWR.n494 2.33701
R3785 VPWR.n612 VPWR.n611 2.33701
R3786 VPWR.n458 VPWR.n457 2.33701
R3787 VPWR.n353 VPWR.n352 2.33701
R3788 VPWR.n427 VPWR.n354 2.33701
R3789 VPWR.n396 VPWR.n364 2.33701
R3790 VPWR.n374 VPWR.n373 2.33701
R3791 VPWR.n5865 VPWR.n5864 2.33701
R3792 VPWR.n5508 VPWR.n5507 2.33701
R3793 VPWR.n6005 VPWR.n6004 2.33701
R3794 VPWR.n5384 VPWR.n5383 2.33701
R3795 VPWR.n5385 VPWR.n5384 2.33701
R3796 VPWR.n5622 VPWR.n5621 2.33701
R3797 VPWR.n6237 VPWR.n6236 2.33701
R3798 VPWR.n6122 VPWR.n6121 2.33701
R3799 VPWR.n6132 VPWR.n6131 2.33701
R3800 VPWR.n86 VPWR.n85 2.33701
R3801 VPWR.n6145 VPWR.n6144 2.33701
R3802 VPWR.n6153 VPWR.n6152 2.33701
R3803 VPWR.n2134 VPWR.n2133 2.33701
R3804 VPWR.n2122 VPWR.n2121 2.33701
R3805 VPWR.n2540 VPWR.n2539 2.33701
R3806 VPWR.n2528 VPWR.n2527 2.33701
R3807 VPWR.n1633 VPWR.n1620 2.33701
R3808 VPWR.n1619 VPWR.n1617 2.33701
R3809 VPWR.n1616 VPWR.n1614 2.33701
R3810 VPWR.n2696 VPWR.n2645 2.33701
R3811 VPWR.n2645 VPWR.n2644 2.33701
R3812 VPWR.n2723 VPWR.n2722 2.33701
R3813 VPWR.n1534 VPWR.n1523 2.33701
R3814 VPWR.n1722 VPWR.n1721 2.33701
R3815 VPWR.n1735 VPWR.n1734 2.33701
R3816 VPWR.n1691 VPWR.n1689 2.33701
R3817 VPWR.n1768 VPWR.n1767 2.33701
R3818 VPWR.n2964 VPWR.n2963 2.33701
R3819 VPWR.n2963 VPWR.n2962 2.33701
R3820 VPWR.n2954 VPWR.n1771 2.33701
R3821 VPWR.n2947 VPWR.n1772 2.33701
R3822 VPWR.n1972 VPWR.n1971 2.33701
R3823 VPWR.n3422 VPWR.n3421 2.33701
R3824 VPWR.n1352 VPWR.n1333 2.33701
R3825 VPWR.n1366 VPWR.n1365 2.33701
R3826 VPWR.n1489 VPWR.n1488 2.33701
R3827 VPWR.n3169 VPWR.n3168 2.33701
R3828 VPWR.n1148 VPWR.n1147 2.33701
R3829 VPWR.n3613 VPWR.n3612 2.33701
R3830 VPWR.n1223 VPWR.n1222 2.33701
R3831 VPWR.n1216 VPWR.n1215 2.33701
R3832 VPWR.n3708 VPWR.n1217 2.33701
R3833 VPWR.n3886 VPWR.n3885 2.33701
R3834 VPWR.n1015 VPWR.n999 2.33701
R3835 VPWR.n1028 VPWR.n996 2.33701
R3836 VPWR.n992 VPWR.n990 2.33701
R3837 VPWR.n4064 VPWR.n4038 2.33701
R3838 VPWR.n4036 VPWR.n4035 2.33701
R3839 VPWR.n4083 VPWR.n4082 2.33701
R3840 VPWR.n3941 VPWR.n3930 2.33701
R3841 VPWR.n3928 VPWR.n3927 2.33701
R3842 VPWR.n3906 VPWR.n3905 2.33701
R3843 VPWR.n4162 VPWR.n4161 2.33701
R3844 VPWR.n4176 VPWR.n4175 2.33701
R3845 VPWR.n4190 VPWR.n4189 2.33701
R3846 VPWR.n739 VPWR.n738 2.33701
R3847 VPWR.n916 VPWR.n915 2.33701
R3848 VPWR.n4259 VPWR.n4258 2.33701
R3849 VPWR.n4270 VPWR.n4269 2.33701
R3850 VPWR.n4334 VPWR.n4333 2.33701
R3851 VPWR.n4846 VPWR.n4845 2.33701
R3852 VPWR.n4857 VPWR.n4856 2.33701
R3853 VPWR.n4869 VPWR.n4868 2.33701
R3854 VPWR.n4437 VPWR.n4436 2.33701
R3855 VPWR.n4534 VPWR.n4533 2.33701
R3856 VPWR.n4552 VPWR.n4551 2.33701
R3857 VPWR.n4767 VPWR.n4589 2.33701
R3858 VPWR.n4758 VPWR.n4757 2.33701
R3859 VPWR.n4745 VPWR.n4744 2.33701
R3860 VPWR.n4744 VPWR.n4743 2.33701
R3861 VPWR.n4730 VPWR.n4729 2.33701
R3862 VPWR.n4962 VPWR.n4961 2.33701
R3863 VPWR.n5123 VPWR.n5122 2.33701
R3864 VPWR.n5105 VPWR.n5103 2.33701
R3865 VPWR.n5064 VPWR.n5063 2.33701
R3866 VPWR.n5174 VPWR.n5173 2.33701
R3867 VPWR.n5208 VPWR.n5207 2.33701
R3868 VPWR.n5346 VPWR.n5345 2.33701
R3869 VPWR.n5323 VPWR.n5321 2.33701
R3870 VPWR.n557 VPWR.n498 2.33701
R3871 VPWR.n436 VPWR.n353 2.33701
R3872 VPWR.n430 VPWR.n354 2.33701
R3873 VPWR.n419 VPWR.n418 2.33701
R3874 VPWR.n418 VPWR.n417 2.33701
R3875 VPWR.n410 VPWR.n409 2.33701
R3876 VPWR.n409 VPWR.n408 2.33701
R3877 VPWR.n399 VPWR.n364 2.33701
R3878 VPWR.n379 VPWR.n374 2.33701
R3879 VPWR.n5864 VPWR.n5863 2.33701
R3880 VPWR.n5509 VPWR.n5508 2.33701
R3881 VPWR.n5994 VPWR.n5993 2.33701
R3882 VPWR.n6006 VPWR.n6005 2.33701
R3883 VPWR.n3481 VPWR.n3480 2.33695
R3884 VPWR.n5097 VPWR.n680 2.33695
R3885 VPWR.n2840 VPWR.n2839 2.29662
R3886 VPWR.n2841 VPWR.n2776 2.29662
R3887 VPWR.n2845 VPWR.n2844 2.29662
R3888 VPWR.n2847 VPWR.n2846 2.29662
R3889 VPWR.n2855 VPWR.n2854 2.29662
R3890 VPWR.n2858 VPWR.n2857 2.29662
R3891 VPWR.n1965 VPWR.n1964 2.29662
R3892 VPWR.n1968 VPWR.n1967 2.29662
R3893 VPWR.n1978 VPWR.n1977 2.29662
R3894 VPWR.n3002 VPWR.n2995 2.29662
R3895 VPWR.n3301 VPWR.n1494 2.29662
R3896 VPWR.n3305 VPWR.n3304 2.29662
R3897 VPWR.n3326 VPWR.n3325 2.29662
R3898 VPWR.n3379 VPWR.n3378 2.29662
R3899 VPWR.n3380 VPWR.n1412 2.29662
R3900 VPWR.n3406 VPWR.n3405 2.29662
R3901 VPWR.n3321 VPWR.n1492 2.29662
R3902 VPWR.n3557 VPWR.n3556 2.29662
R3903 VPWR.n3555 VPWR.n1280 2.29662
R3904 VPWR.n3896 VPWR.n3895 2.29662
R3905 VPWR.n3900 VPWR.n3899 2.29662
R3906 VPWR.n3933 VPWR.n1120 2.29662
R3907 VPWR.n3824 VPWR.n3823 2.29662
R3908 VPWR.n5114 VPWR.n5109 2.29662
R3909 VPWR.n5113 VPWR.n5112 2.29662
R3910 VPWR.n570 VPWR.n569 2.29662
R3911 VPWR.n5348 VPWR.n5332 2.29662
R3912 VPWR.n568 VPWR.n567 2.29662
R3913 VPWR.n207 VPWR.n206 2.29662
R3914 VPWR.n220 VPWR.n219 2.29662
R3915 VPWR.n5973 VPWR.n5972 2.29662
R3916 VPWR.n6094 VPWR.n91 2.29662
R3917 VPWR.n2853 VPWR.n2852 2.29643
R3918 VPWR.n2674 VPWR.n2673 2.29643
R3919 VPWR.n1625 VPWR.n1622 2.29643
R3920 VPWR.n3435 VPWR.n1409 2.29643
R3921 VPWR.n3410 VPWR.n3409 2.29643
R3922 VPWR.n3162 VPWR.n3156 2.29643
R3923 VPWR.n3725 VPWR.n3724 2.29643
R3924 VPWR.n4009 VPWR.n4008 2.29643
R3925 VPWR.n4070 VPWR.n4069 2.29643
R3926 VPWR.n3901 VPWR.n1129 2.29643
R3927 VPWR.n3912 VPWR.n3911 2.29643
R3928 VPWR.n3934 VPWR.n3931 2.29643
R3929 VPWR.n733 VPWR.n732 2.29643
R3930 VPWR.n4431 VPWR.n4430 2.29643
R3931 VPWR.n4774 VPWR.n4773 2.29643
R3932 VPWR.n5136 VPWR.n5134 2.29643
R3933 VPWR.n6105 VPWR.n6104 2.29643
R3934 VPWR.n3358 VPWR.n3357 2.28621
R3935 VPWR.n3839 VPWR.n3838 2.28175
R3936 VPWR.n4999 VPWR.n4998 2.28175
R3937 VPWR.n58 VPWR.n57 2.28175
R3938 VPWR.n5933 VPWR.n5925 2.27705
R3939 VPWR.n2766 VPWR.n2765 2.23542
R3940 VPWR.n1553 VPWR.n1552 2.23542
R3941 VPWR.n1975 VPWR.n1974 2.23542
R3942 VPWR.n3361 VPWR.n3358 2.23542
R3943 VPWR.n876 VPWR.n874 2.23542
R3944 VPWR.n4242 VPWR.n4241 2.23542
R3945 VPWR.n4300 VPWR.n4299 2.23542
R3946 VPWR.n5221 VPWR.n5220 2.23542
R3947 VPWR.n5046 VPWR.n5045 2.23542
R3948 VPWR.n4981 VPWR.n4980 2.23542
R3949 VPWR.n579 VPWR.n578 2.23542
R3950 VPWR.n6220 VPWR.n6219 2.22736
R3951 VPWR.n5929 VPWR.n5928 2.19376
R3952 VPWR.n2813 VPWR.n2812 2.19376
R3953 VPWR.n2942 VPWR.n2941 2.18463
R3954 VPWR.n457 VPWR.n456 2.18463
R3955 VPWR.n1607 VPWR.n1606 2.08304
R3956 VPWR.n2248 VPWR.n2247 2.08304
R3957 VPWR.n2081 VPWR.n2080 2.08304
R3958 VPWR.n1689 VPWR.n1688 2.08304
R3959 VPWR.n990 VPWR.n989 2.08304
R3960 VPWR.n4593 VPWR.n4592 2.08304
R3961 VPWR.n5321 VPWR.n5320 2.08304
R3962 VPWR.n1932 VPWR.n1931 1.87987
R3963 VPWR.n3273 VPWR.n3272 1.87987
R3964 VPWR.n3740 VPWR.n3739 1.87987
R3965 VPWR.n860 VPWR.n859 1.87987
R3966 VPWR.n4467 VPWR.n4466 1.87987
R3967 VPWR.n5900 VPWR.n5857 1.81937
R3968 VPWR.n5639 VPWR.n5592 1.81774
R3969 VPWR.n6300 VPWR.n6299 1.79825
R3970 VPWR.n5964 VPWR.n5963 1.69039
R3971 VPWR VPWR 1.67895
R3972 VPWR VPWR 1.67895
R3973 VPWR VPWR 1.67895
R3974 VPWR VPWR 1.67895
R3975 VPWR VPWR 1.67895
R3976 VPWR VPWR 1.67895
R3977 VPWR VPWR 1.67895
R3978 VPWR VPWR 1.67895
R3979 VPWR VPWR 1.67895
R3980 VPWR VPWR 1.67895
R3981 VPWR VPWR 1.67895
R3982 VPWR VPWR 1.67895
R3983 VPWR VPWR 1.67895
R3984 VPWR.n4819 VPWR.n4818 1.67669
R3985 VPWR.n46 VPWR.n44 1.66178
R3986 VPWR.n94 VPWR.n93 1.66178
R3987 VPWR.n1482 VPWR.n1481 1.6259
R3988 VPWR.n648 VPWR.n647 1.6259
R3989 VPWR.n2503 VPWR.n2502 1.51061
R3990 VPWR.n2825 VPWR.n2824 1.51061
R3991 VPWR.n5964 VPWR.n5962 1.51061
R3992 VPWR.n1526 VPWR.n1525 1.50646
R3993 VPWR.n1846 VPWR.n1845 1.50646
R3994 VPWR.n3158 VPWR.n3157 1.50646
R3995 VPWR.n1143 VPWR.n1142 1.50646
R3996 VPWR.n3814 VPWR.n3813 1.50646
R3997 VPWR.n705 VPWR.n704 1.50646
R3998 VPWR.n4403 VPWR.n4402 1.50646
R3999 VPWR.n4948 VPWR.n4947 1.50646
R4000 VPWR.n195 VPWR.n194 1.50646
R4001 VPWR.n5867 VPWR.n5866 1.50646
R4002 VPWR.n1 VPWR.n0 1.50646
R4003 VPWR.n2904 VPWR.n2903 1.49961
R4004 VPWR.n2999 VPWR.n2998 1.49961
R4005 VPWR.n708 VPWR.n702 1.49961
R4006 VPWR.n4661 VPWR.n4660 1.49961
R4007 VPWR.n4952 VPWR.n4951 1.49961
R4008 VPWR.n598 VPWR.n491 1.49961
R4009 VPWR.n386 VPWR.n368 1.49961
R4010 VPWR.n5875 VPWR.n5860 1.49961
R4011 VPWR.n6200 VPWR.n70 1.49961
R4012 VPWR.n1624 VPWR.n1623 1.49932
R4013 VPWR.n1703 VPWR.n1702 1.49932
R4014 VPWR.n3372 VPWR.n1414 1.49932
R4015 VPWR.n1339 VPWR.n1338 1.49932
R4016 VPWR.n3484 VPWR.n3483 1.49932
R4017 VPWR.n1005 VPWR.n1002 1.49932
R4018 VPWR.n1004 VPWR.n1003 1.49932
R4019 VPWR.n4154 VPWR.n4153 1.49932
R4020 VPWR.n4406 VPWR.n4401 1.49932
R4021 VPWR.n4524 VPWR.n4521 1.49932
R4022 VPWR.n4523 VPWR.n4522 1.49932
R4023 VPWR.n267 VPWR.n266 1.49932
R4024 VPWR.n533 VPWR.n503 1.49932
R4025 VPWR.n5338 VPWR.n5337 1.49932
R4026 VPWR.n5872 VPWR.n5861 1.49932
R4027 VPWR.n5695 VPWR.n5694 1.49932
R4028 VPWR.n5597 VPWR.n5596 1.49932
R4029 VPWR.n5962 VPWR.n5960 1.47466
R4030 VPWR.n5363 VPWR.n5328 1.47445
R4031 VPWR.n58 VPWR.n40 1.47352
R4032 VPWR.n2684 VPWR.n2683 1.47352
R4033 VPWR.n2735 VPWR.n2734 1.47352
R4034 VPWR.n1535 VPWR.n1534 1.47352
R4035 VPWR.n3418 VPWR.n3398 1.47352
R4036 VPWR.n3340 VPWR.n1484 1.47352
R4037 VPWR.n1483 VPWR.n1482 1.47352
R4038 VPWR.n3173 VPWR.n3152 1.47352
R4039 VPWR.n1154 VPWR.n1141 1.47352
R4040 VPWR.n3702 VPWR.n3701 1.47352
R4041 VPWR.n4034 VPWR.n4033 1.47352
R4042 VPWR.n4145 VPWR.n4144 1.47352
R4043 VPWR.n4561 VPWR.n4560 1.47352
R4044 VPWR.n4799 VPWR.n4798 1.47352
R4045 VPWR.n4714 VPWR.n4591 1.47352
R4046 VPWR.n4968 VPWR.n4967 1.47352
R4047 VPWR.n677 VPWR.n648 1.47352
R4048 VPWR.n5346 VPWR.n5332 1.47352
R4049 VPWR.n5786 VPWR.n228 1.47352
R4050 VPWR.n4975 VPWR.n4939 1.40734
R4051 VPWR.n3010 VPWR.n2994 1.40583
R4052 VPWR.n5716 VPWR.n5715 1.30773
R4053 VPWR.n3628 VPWR.n1253 1.26921
R4054 VPWR.n3991 VPWR.n3990 1.26921
R4055 VPWR.n717 VPWR.n716 1.22883
R4056 VPWR.n4415 VPWR.n4414 1.22883
R4057 VPWR.n4693 VPWR.n4692 1.22883
R4058 VPWR.n554 VPWR.n499 1.22883
R4059 VPWR.n6085 VPWR.n6084 1.22603
R4060 VPWR.n23 VPWR.n22 1.22603
R4061 VPWR.n6086 VPWR.n6085 1.1988
R4062 VPWR.n5889 VPWR.n5888 1.1988
R4063 VPWR.n5895 VPWR.n5894 1.1988
R4064 VPWR.n5715 VPWR.n5714 1.1988
R4065 VPWR.n2265 VPWR.n2262 1.16875
R4066 VPWR.n2403 VPWR.n2402 1.16875
R4067 VPWR.n2913 VPWR.n2617 1.14176
R4068 VPWR.n3449 VPWR.n1310 1.14176
R4069 VPWR.n3467 VPWR.n3466 1.14176
R4070 VPWR.n4095 VPWR.n1043 1.14176
R4071 VPWR.n4706 VPWR.n4705 1.14176
R4072 VPWR.n5154 VPWR.n5153 1.14176
R4073 VPWR.n623 VPWR.n333 1.14176
R4074 VPWR.n2478 VPWR.n2477 1.1414
R4075 VPWR.n3117 VPWR.n3116 1.14113
R4076 VPWR.n3879 VPWR.n3878 1.14113
R4077 VPWR.n3780 VPWR.n3779 1.14113
R4078 VPWR.n3219 VPWR.n3218 1.14113
R4079 VPWR.n5813 VPWR.n5812 1.14113
R4080 VPWR.n5037 VPWR.n5036 1.14113
R4081 VPWR.n4915 VPWR.n4914 1.14113
R4082 VPWR.n5954 VPWR.n5953 1.14113
R4083 VPWR.n5842 VPWR.n5841 1.14113
R4084 VPWR.n4095 VPWR.n4094 1.14113
R4085 VPWR.n3466 VPWR.n3465 1.14113
R4086 VPWR.n3449 VPWR.n3448 1.14113
R4087 VPWR.n5744 VPWR.n5561 1.14113
R4088 VPWR.n2913 VPWR.n2912 1.14113
R4089 VPWR.n3981 VPWR.n3980 1.14113
R4090 VPWR.n1434 VPWR.n1237 1.14113
R4091 VPWR.n3347 VPWR.n3346 1.14113
R4092 VPWR.n623 VPWR.n622 1.14113
R4093 VPWR.n5153 VPWR.n5152 1.14113
R4094 VPWR.n4705 VPWR.n4704 1.14113
R4095 VPWR.n6065 VPWR.n6064 1.14113
R4096 VPWR.n149 VPWR.n148 1.14113
R4097 VPWR.n5643 VPWR.n5642 1.14002
R4098 VPWR.n5744 VPWR.n5743 1.1392
R4099 VPWR.n2311 VPWR.n2310 1.1392
R4100 VPWR.n2601 VPWR.n2047 1.1392
R4101 VPWR.n2601 VPWR.n2600 1.1392
R4102 VPWR.n3067 VPWR.n1664 1.13909
R4103 VPWR.n5763 VPWR.n5377 1.13909
R4104 VPWR.n5282 VPWR.n296 1.13909
R4105 VPWR.n4576 VPWR.n4566 1.13909
R4106 VPWR.n3125 VPWR.n3124 1.1368
R4107 VPWR.n3801 VPWR.n3800 1.1368
R4108 VPWR.n3788 VPWR.n3787 1.1368
R4109 VPWR.n3148 VPWR.n3147 1.1368
R4110 VPWR.n5821 VPWR.n5820 1.1368
R4111 VPWR.n4935 VPWR.n4934 1.1368
R4112 VPWR.n4923 VPWR.n4922 1.1368
R4113 VPWR.n5853 VPWR.n5852 1.1368
R4114 VPWR.n5661 VPWR.n5660 1.1368
R4115 VPWR.n2221 VPWR.n2220 1.1368
R4116 VPWR.n5654 VPWR.n5653 1.1368
R4117 VPWR.n2607 VPWR.n2606 1.1368
R4118 VPWR.n1089 VPWR.n1088 1.1368
R4119 VPWR.n1433 VPWR.n1432 1.1368
R4120 VPWR.n1450 VPWR.n1449 1.1368
R4121 VPWR.n6072 VPWR.n6071 1.1368
R4122 VPWR.n113 VPWR.n112 1.1368
R4123 VPWR.n2805 VPWR.n1516 1.13669
R4124 VPWR.n3881 VPWR.n3880 1.13669
R4125 VPWR.n1197 VPWR.n1136 1.13669
R4126 VPWR.n3221 VPWR.n3220 1.13669
R4127 VPWR.n529 VPWR.n180 1.13669
R4128 VPWR.n5039 VPWR.n5038 1.13669
R4129 VPWR.n4454 VPWR.n4395 1.13669
R4130 VPWR.n5956 VPWR.n5955 1.13669
R4131 VPWR.n2468 VPWR.n2467 1.13669
R4132 VPWR.n2476 VPWR.n2474 1.13669
R4133 VPWR.n3070 VPWR.n3068 1.13669
R4134 VPWR.n3066 VPWR.n3065 1.13669
R4135 VPWR.n1048 VPWR.n1047 1.13669
R4136 VPWR.n4101 VPWR.n4100 1.13669
R4137 VPWR.n3462 VPWR.n3461 1.13669
R4138 VPWR.n1307 VPWR.n1306 1.13669
R4139 VPWR.n1315 VPWR.n1314 1.13669
R4140 VPWR.n3455 VPWR.n3454 1.13669
R4141 VPWR.n5750 VPWR.n5749 1.13669
R4142 VPWR.n5766 VPWR.n5764 1.13669
R4143 VPWR.n5762 VPWR.n5761 1.13669
R4144 VPWR.n5281 VPWR.n5280 1.13669
R4145 VPWR.n5290 VPWR.n5289 1.13669
R4146 VPWR.n4579 VPWR.n4577 1.13669
R4147 VPWR.n4575 VPWR.n4574 1.13669
R4148 VPWR.n2317 VPWR.n2313 1.13669
R4149 VPWR.n2044 VPWR.n2043 1.13669
R4150 VPWR.n2614 VPWR.n2613 1.13669
R4151 VPWR.n2919 VPWR.n2918 1.13669
R4152 VPWR.n3983 VPWR.n3982 1.13669
R4153 VPWR.n1440 VPWR.n1439 1.13669
R4154 VPWR.n3349 VPWR.n3348 1.13669
R4155 VPWR.n628 VPWR.n627 1.13669
R4156 VPWR.n330 VPWR.n329 1.13669
R4157 VPWR.n641 VPWR.n640 1.13669
R4158 VPWR.n636 VPWR.n635 1.13669
R4159 VPWR.n4620 VPWR.n4619 1.13669
R4160 VPWR.n4614 VPWR.n4613 1.13669
R4161 VPWR.n5448 VPWR.n150 1.13669
R4162 VPWR.n6076 VPWR.n6075 1.13669
R4163 VPWR.n5969 VPWR.n5968 1.11511
R4164 VPWR.n6299 VPWR.n6298 1.11511
R4165 VPWR.n1948 VPWR.n1818 1.09272
R4166 VPWR.n3434 VPWR.n3392 1.09272
R4167 VPWR.n3160 VPWR.n3159 1.09272
R4168 VPWR.n3726 VPWR.n1211 1.09272
R4169 VPWR.n3913 VPWR.n1125 1.09272
R4170 VPWR.n897 VPWR.n820 1.09272
R4171 VPWR.n4834 VPWR.n4473 1.09272
R4172 VPWR.n275 VPWR.n274 1.09272
R4173 VPWR.n5974 VPWR.n173 1.09272
R4174 VPWR.n1528 VPWR.n1527 1.09216
R4175 VPWR.n1848 VPWR.n1847 1.09216
R4176 VPWR.n3017 VPWR.n3016 1.09216
R4177 VPWR.n3388 VPWR.n1411 1.09216
R4178 VPWR.n3261 VPWR.n3235 1.09216
R4179 VPWR.n3240 VPWR.n1495 1.09216
R4180 VPWR.n1340 VPWR.n1337 1.09216
R4181 VPWR.n3603 VPWR.n3602 1.09216
R4182 VPWR.n3578 VPWR.n1271 1.09216
R4183 VPWR.n1163 VPWR.n1162 1.09216
R4184 VPWR.n4012 VPWR.n1068 1.09216
R4185 VPWR.n3816 VPWR.n3815 1.09216
R4186 VPWR.n896 VPWR.n821 1.09216
R4187 VPWR.n4686 VPWR.n4656 1.09216
R4188 VPWR.n4788 VPWR.n4584 1.09216
R4189 VPWR.n278 VPWR.n277 1.09216
R4190 VPWR.n269 VPWR.n268 1.09216
R4191 VPWR.n542 VPWR.n501 1.09216
R4192 VPWR.n196 VPWR.n193 1.09216
R4193 VPWR.n5697 VPWR.n5696 1.09216
R4194 VPWR.n6214 VPWR.n6213 1.09216
R4195 VPWR.n3 VPWR.n2 1.09216
R4196 VPWR.n6305 VPWR.n10 1.09216
R4197 VPWR.n5530 VPWR.n5529 1.09203
R4198 VPWR.n5496 VPWR.n5407 1.09203
R4199 VPWR.n6226 VPWR.n63 1.09203
R4200 VPWR.n6298 VPWR.n23 1.04908
R4201 VPWR.n53 VPWR.n52 0.998665
R4202 VPWR.n679 VPWR.n678 0.990318
R4203 VPWR.n3833 VPWR.n3805 0.958125
R4204 VPWR.n2259 VPWR.n2258 0.935332
R4205 VPWR.n2577 VPWR.n2576 0.935332
R4206 VPWR.n5743 VPWR.n5742 0.872922
R4207 VPWR.n2310 VPWR.n2309 0.872922
R4208 VPWR.n2600 VPWR.n2599 0.872922
R4209 VPWR.n1664 VPWR.n1663 0.872255
R4210 VPWR.n4566 VPWR.n4565 0.872255
R4211 VPWR.n296 VPWR.n295 0.872255
R4212 VPWR.n5377 VPWR.n5376 0.872255
R4213 VPWR.n1748 VPWR.n1747 0.871602
R4214 VPWR.n2479 VPWR.n2478 0.871546
R4215 VPWR.n1378 VPWR.n1310 0.871525
R4216 VPWR.n3528 VPWR.n3467 0.871525
R4217 VPWR.n1043 VPWR.n1042 0.871525
R4218 VPWR.n5642 VPWR.n5641 0.871359
R4219 VPWR.n2912 VPWR.n2911 0.871338
R4220 VPWR.n3346 VPWR.n3345 0.871338
R4221 VPWR.n3653 VPWR.n1237 0.871338
R4222 VPWR.n3980 VPWR.n3979 0.871338
R4223 VPWR.n622 VPWR.n621 0.871338
R4224 VPWR.n5152 VPWR.n5151 0.871338
R4225 VPWR.n4704 VPWR.n4703 0.871338
R4226 VPWR.n6064 VPWR.n6063 0.871338
R4227 VPWR.n148 VPWR.n147 0.871338
R4228 VPWR.n2035 VPWR.n2034 0.871205
R4229 VPWR.n4094 VPWR.n4093 0.870036
R4230 VPWR.n3465 VPWR.n1282 0.870036
R4231 VPWR.n3448 VPWR.n3447 0.870036
R4232 VPWR.n5561 VPWR.n5560 0.870036
R4233 VPWR.n4203 VPWR.n4202 0.869838
R4234 VPWR.n954 VPWR.n953 0.86965
R4235 VPWR.n2807 VPWR.n2806 0.86965
R4236 VPWR.n1929 VPWR.n1928 0.86965
R4237 VPWR.n3277 VPWR.n3222 0.86965
R4238 VPWR.n3744 VPWR.n1198 0.86965
R4239 VPWR.n3883 VPWR.n3882 0.86965
R4240 VPWR.n857 VPWR.n856 0.86965
R4241 VPWR.n4880 VPWR.n4455 0.86965
R4242 VPWR.n5041 VPWR.n5040 0.86965
R4243 VPWR.n531 VPWR.n530 0.86965
R4244 VPWR.n5958 VPWR.n5957 0.86965
R4245 VPWR.n5644 VPWR.n81 0.869615
R4246 VPWR.n3039 VPWR.n3038 0.86907
R4247 VPWR.n5953 VPWR.n5952 0.868734
R4248 VPWR.n5812 VPWR.n5811 0.868734
R4249 VPWR.n5036 VPWR.n5035 0.868734
R4250 VPWR.n4914 VPWR.n4913 0.868734
R4251 VPWR.n3878 VPWR.n3877 0.868734
R4252 VPWR.n3779 VPWR.n3778 0.868734
R4253 VPWR.n3218 VPWR.n3217 0.868734
R4254 VPWR.n3116 VPWR.n3115 0.868734
R4255 VPWR.n5841 VPWR.n26 0.868734
R4256 VPWR.n1839 VPWR.n1838 0.868685
R4257 VPWR.n4112 VPWR.n757 0.868348
R4258 VPWR.n2319 VPWR.n2318 0.868348
R4259 VPWR.n3072 VPWR.n3071 0.868348
R4260 VPWR.n4581 VPWR.n4580 0.868348
R4261 VPWR.n5279 VPWR.n5278 0.868348
R4262 VPWR.n5768 VPWR.n5767 0.868348
R4263 VPWR.n4383 VPWR.n4382 0.867046
R4264 VPWR.n2464 VPWR.n2463 0.867046
R4265 VPWR.n2250 VPWR.n2249 0.863992
R4266 VPWR.n2085 VPWR.n2084 0.863992
R4267 VPWR.n2453 VPWR.n2452 0.863992
R4268 VPWR.n1609 VPWR.n1608 0.863992
R4269 VPWR.n2624 VPWR.n2623 0.863992
R4270 VPWR.n1691 VPWR.n1690 0.863992
R4271 VPWR.n3440 VPWR.n1405 0.863992
R4272 VPWR.n1329 VPWR.n1328 0.863992
R4273 VPWR.n1484 VPWR.n1483 0.863992
R4274 VPWR.n1293 VPWR.n1289 0.863992
R4275 VPWR.n3473 VPWR.n3472 0.863992
R4276 VPWR.n992 VPWR.n991 0.863992
R4277 VPWR.n882 VPWR 0.863992
R4278 VPWR.n4146 VPWR.n4145 0.863992
R4279 VPWR.n4514 VPWR.n4513 0.863992
R4280 VPWR.n4792 VPWR 0.863992
R4281 VPWR.n4598 VPWR.n4597 0.863992
R4282 VPWR.n259 VPWR.n258 0.863992
R4283 VPWR VPWR.n5098 0.863992
R4284 VPWR.n678 VPWR.n677 0.863992
R4285 VPWR.n5323 VPWR.n5322 0.863992
R4286 VPWR.n389 VPWR 0.863992
R4287 VPWR.n2105 VPWR.n2047 0.855994
R4288 VPWR.n2933 VPWR.n2932 0.854674
R4289 VPWR.n2629 VPWR.n2617 0.854598
R4290 VPWR.n344 VPWR.n333 0.854598
R4291 VPWR.n5155 VPWR.n5154 0.854598
R4292 VPWR.n4707 VPWR.n4706 0.854598
R4293 VPWR.n4228 VPWR.n4227 0.852723
R4294 VPWR.n6078 VPWR.n6077 0.852723
R4295 VPWR.n3351 VPWR.n3350 0.852723
R4296 VPWR.n1438 VPWR.n1244 0.852723
R4297 VPWR.n3985 VPWR.n3984 0.852723
R4298 VPWR.n5450 VPWR.n5449 0.852723
R4299 VPWR.n2667 VPWR.n2653 0.842756
R4300 VPWR.n5133 VPWR.n5101 0.842756
R4301 VPWR.n1856 VPWR.n1855 0.835507
R4302 VPWR.n431 VPWR 0.813198
R4303 VPWR.n5885 VPWR.n5884 0.802048
R4304 VPWR.n12 VPWR.n11 0.791511
R4305 VPWR.n2494 VPWR.n2493 0.791511
R4306 VPWR.n2814 VPWR.n2813 0.791511
R4307 VPWR.n5716 VPWR.n5710 0.790287
R4308 VPWR.n2083 VPWR.n2082 0.711611
R4309 VPWR.n1481 VPWR.n1480 0.711611
R4310 VPWR.n4596 VPWR.n4595 0.711611
R4311 VPWR.n647 VPWR.n646 0.711611
R4312 VPWR.n5975 VPWR.n162 0.67208
R4313 VPWR.n6251 VPWR.n46 0.67208
R4314 VPWR.n5823 VPWR.n179 0.668275
R4315 VPWR.n1405 VPWR.n1404 0.610024
R4316 VPWR.n1289 VPWR.n1288 0.610024
R4317 VPWR.n221 VPWR.n185 0.608239
R4318 VPWR.n2257 VPWR.n2254 0.539826
R4319 VPWR.n2582 VPWR.n2581 0.539826
R4320 VPWR.n16 VPWR.n13 0.503871
R4321 VPWR.n2492 VPWR.n2491 0.503871
R4322 VPWR.n2819 VPWR.n2818 0.503871
R4323 VPWR.n5933 VPWR.n5932 0.503871
R4324 VPWR.n5752 VPWR.n179 0.478275
R4325 VPWR.n1511 VPWR.n1510 0.473873
R4326 VPWR.n4213 VPWR.n690 0.473873
R4327 VPWR.n897 VPWR.n896 0.470249
R4328 VPWR.n4211 VPWR.n4210 0.469446
R4329 VPWR.n1508 VPWR.n1507 0.466417
R4330 VPWR.n95 VPWR.n94 0.463479
R4331 VPWR.n5146 VPWR.n679 0.427908
R4332 VPWR.n170 VPWR.n169 0.419768
R4333 VPWR.n5134 VPWR.n5133 0.410386
R4334 VPWR.n3159 VPWR.n3158 0.407316
R4335 VPWR.n2451 VPWR.n2450 0.406849
R4336 VPWR.n1527 VPWR.n1526 0.404857
R4337 VPWR.n1847 VPWR.n1846 0.404857
R4338 VPWR.n3815 VPWR.n3814 0.404857
R4339 VPWR.n196 VPWR.n195 0.404857
R4340 VPWR.n2 VPWR.n1 0.404857
R4341 VPWR.n221 VPWR 0.398022
R4342 VPWR.n5977 VPWR.n5975 0.397684
R4343 VPWR.n6251 VPWR.n6250 0.397684
R4344 VPWR.n93 VPWR.n92 0.381777
R4345 VPWR.n4387 VPWR.n4386 0.3805
R4346 VPWR.n4387 VPWR.n693 0.3805
R4347 VPWR.n4387 VPWR.n689 0.3805
R4348 VPWR.n4207 VPWR.n4116 0.3805
R4349 VPWR.n4207 VPWR.n4119 0.3805
R4350 VPWR.n4207 VPWR.n4206 0.3805
R4351 VPWR.n4224 VPWR.n4223 0.3805
R4352 VPWR.n4223 VPWR.n957 0.3805
R4353 VPWR.n4223 VPWR.n4222 0.3805
R4354 VPWR.n5975 VPWR 0.379742
R4355 VPWR VPWR.n6251 0.379742
R4356 VPWR.n3435 VPWR.n3434 0.356134
R4357 VPWR.n3913 VPWR.n3912 0.356134
R4358 VPWR.n699 VPWR.n698 0.342728
R4359 VPWR.n4110 VPWR.n4109 0.342728
R4360 VPWR.n784 VPWR.n783 0.342728
R4361 VPWR.n3130 VPWR.n1513 0.3424
R4362 VPWR VPWR.n2667 0.329918
R4363 VPWR.n2812 VPWR.n2811 0.324095
R4364 VPWR.n3135 VPWR.n3134 0.31175
R4365 VPWR.n3049 VPWR.n3048 0.311379
R4366 VPWR.n2927 VPWR.n2926 0.311379
R4367 VPWR.n1781 VPWR.n1780 0.311379
R4368 VPWR.n3055 VPWR.n3054 0.311321
R4369 VPWR.n3050 VPWR.n3042 0.309572
R4370 VPWR.n3050 VPWR.n1751 0.309572
R4371 VPWR.n2929 VPWR.n2928 0.309572
R4372 VPWR.n2928 VPWR.n2038 0.309572
R4373 VPWR.n3130 VPWR.n1515 0.309146
R4374 VPWR.n3130 VPWR.n1503 0.309146
R4375 VPWR.n2450 VPWR.n2449 0.305262
R4376 VPWR.n5498 VPWR.n5496 0.295115
R4377 VPWR.n6226 VPWR.n6225 0.295115
R4378 VPWR.n3603 VPWR.n3600 0.294041
R4379 VPWR.n3578 VPWR.n3577 0.294041
R4380 VPWR.n4687 VPWR.n4686 0.294041
R4381 VPWR.n270 VPWR.n269 0.294041
R4382 VPWR.n5698 VPWR.n5697 0.294041
R4383 VPWR.n3833 VPWR 0.292135
R4384 VPWR.n2810 VPWR.n2809 0.28814
R4385 VPWR.n5928 VPWR.n5927 0.28814
R4386 VPWR VPWR.n4834 0.275667
R4387 VPWR.n274 VPWR 0.274365
R4388 VPWR.n5974 VPWR 0.274365
R4389 VPWR.n5496 VPWR 0.272723
R4390 VPWR VPWR.n3017 0.271905
R4391 VPWR.n3235 VPWR 0.271905
R4392 VPWR VPWR.n3240 0.271905
R4393 VPWR.n3388 VPWR 0.271905
R4394 VPWR.n1162 VPWR 0.271905
R4395 VPWR.n4012 VPWR 0.271905
R4396 VPWR VPWR.n278 0.271905
R4397 VPWR.n10 VPWR 0.271905
R4398 VPWR.n1948 VPWR 0.26525
R4399 VPWR VPWR.n3726 0.26525
R4400 VPWR VPWR.n6226 0.263609
R4401 VPWR VPWR.n1340 0.262791
R4402 VPWR VPWR.n3603 0.262791
R4403 VPWR.n896 VPWR 0.262791
R4404 VPWR.n542 VPWR 0.262791
R4405 VPWR VPWR.n6214 0.262791
R4406 VPWR.n5529 VPWR 0.262307
R4407 VPWR VPWR.n3578 0.261489
R4408 VPWR.n4686 VPWR 0.261489
R4409 VPWR.n4788 VPWR 0.261489
R4410 VPWR.n222 VPWR.n221 0.259761
R4411 VPWR.n3993 VPWR.n3991 0.257284
R4412 VPWR.n2247 VPWR.n2246 0.254468
R4413 VPWR.n2080 VPWR.n2079 0.254468
R4414 VPWR.n2444 VPWR.n2443 0.254468
R4415 VPWR.n1606 VPWR.n1605 0.254468
R4416 VPWR.n2762 VPWR.n1571 0.254468
R4417 VPWR.n1567 VPWR.n1566 0.254468
R4418 VPWR.n1688 VPWR.n1687 0.254468
R4419 VPWR.n1889 VPWR.n1888 0.254468
R4420 VPWR.n1404 VPWR.n1403 0.254468
R4421 VPWR.n3199 VPWR.n3198 0.254468
R4422 VPWR.n1288 VPWR.n1287 0.254468
R4423 VPWR.n1188 VPWR.n1187 0.254468
R4424 VPWR.n989 VPWR.n988 0.254468
R4425 VPWR.n747 VPWR.n746 0.254468
R4426 VPWR.n4143 VPWR.n4142 0.254468
R4427 VPWR.n4445 VPWR.n4444 0.254468
R4428 VPWR.n4512 VPWR.n4511 0.254468
R4429 VPWR.n4592 VPWR.n4475 0.254468
R4430 VPWR.n257 VPWR.n256 0.254468
R4431 VPWR.n4992 VPWR.n4991 0.254468
R4432 VPWR.n5320 VPWR.n5319 0.254468
R4433 VPWR.n2667 VPWR 0.250033
R4434 VPWR.n5133 VPWR 0.250033
R4435 VPWR.n570 VPWR.n568 0.24081
R4436 VPWR.n2847 VPWR.n2845 0.240554
R4437 VPWR.n3934 VPWR.n3933 0.240185
R4438 VPWR.n5752 VPWR 0.239388
R4439 VPWR VPWR.n5861 0.23824
R4440 VPWR.n3374 VPWR.n3372 0.23824
R4441 VPWR.n4525 VPWR.n4524 0.237885
R4442 VPWR.n1505 VPWR 0.235758
R4443 VPWR.n4208 VPWR 0.233458
R4444 VPWR.n1149 VPWR.n1143 0.231108
R4445 VPWR.n706 VPWR.n705 0.231108
R4446 VPWR.n4404 VPWR.n4403 0.231108
R4447 VPWR.n4950 VPWR.n4948 0.231108
R4448 VPWR.n5868 VPWR.n5867 0.231108
R4449 VPWR VPWR.n3001 0.226156
R4450 VPWR VPWR.n6200 0.218736
R4451 VPWR.n2903 VPWR 0.217434
R4452 VPWR.n2998 VPWR 0.217434
R4453 VPWR.n3832 VPWR 0.217434
R4454 VPWR.n5875 VPWR 0.217434
R4455 VPWR.n2507 VPWR.n2506 0.21623
R4456 VPWR.n2811 VPWR.n2810 0.21623
R4457 VPWR.n2829 VPWR.n2828 0.21623
R4458 VPWR.n5927 VPWR.n5926 0.21623
R4459 VPWR.n5969 VPWR.n5967 0.21623
R4460 VPWR VPWR.n1624 0.215749
R4461 VPWR.n1702 VPWR 0.215749
R4462 VPWR.n3372 VPWR 0.215749
R4463 VPWR VPWR.n1339 0.215749
R4464 VPWR VPWR.n1005 0.215749
R4465 VPWR VPWR.n1004 0.215749
R4466 VPWR.n266 VPWR 0.215749
R4467 VPWR VPWR.n5861 0.215749
R4468 VPWR.n5694 VPWR 0.215749
R4469 VPWR.n4661 VPWR 0.208319
R4470 VPWR.n4951 VPWR 0.208319
R4471 VPWR.n598 VPWR 0.208319
R4472 VPWR VPWR.n386 0.208319
R4473 VPWR VPWR.n702 0.207017
R4474 VPWR.n4153 VPWR 0.206635
R4475 VPWR VPWR.n4523 0.206635
R4476 VPWR VPWR.n5338 0.206635
R4477 VPWR VPWR.n5597 0.205688
R4478 VPWR VPWR.n3484 0.205333
R4479 VPWR VPWR.n4401 0.205333
R4480 VPWR.n4357 VPWR.n4356 0.203675
R4481 VPWR.n4825 VPWR.n4824 0.203675
R4482 VPWR.n5529 VPWR 0.197459
R4483 VPWR VPWR.n1948 0.196835
R4484 VPWR.n3434 VPWR 0.196835
R4485 VPWR.n3159 VPWR 0.196835
R4486 VPWR.n3726 VPWR 0.196835
R4487 VPWR VPWR.n3913 0.196835
R4488 VPWR VPWR.n897 0.196835
R4489 VPWR.n4834 VPWR 0.196835
R4490 VPWR.n274 VPWR 0.196835
R4491 VPWR VPWR.n5974 0.196835
R4492 VPWR.n1527 VPWR 0.196385
R4493 VPWR.n1847 VPWR 0.196385
R4494 VPWR.n3017 VPWR 0.196385
R4495 VPWR VPWR.n3235 0.196385
R4496 VPWR.n3240 VPWR 0.196385
R4497 VPWR VPWR.n3388 0.196385
R4498 VPWR.n1340 VPWR 0.196385
R4499 VPWR.n1162 VPWR 0.196385
R4500 VPWR.n3815 VPWR 0.196385
R4501 VPWR VPWR.n4012 0.196385
R4502 VPWR VPWR.n4788 0.196385
R4503 VPWR.n278 VPWR 0.196385
R4504 VPWR.n269 VPWR 0.196385
R4505 VPWR VPWR.n196 0.196385
R4506 VPWR VPWR.n542 0.196385
R4507 VPWR.n5697 VPWR 0.196385
R4508 VPWR.n2 VPWR 0.196385
R4509 VPWR VPWR.n10 0.196385
R4510 VPWR.n6214 VPWR 0.196385
R4511 VPWR.n5753 VPWR.n5752 0.1905
R4512 VPWR.n323 VPWR.n179 0.1905
R4513 VPWR.n533 VPWR.n532 0.189708
R4514 VPWR.n5349 VPWR.n5348 0.180551
R4515 VPWR.n5973 VPWR.n5970 0.180551
R4516 VPWR.n2853 VPWR.n2851 0.179926
R4517 VPWR.n2676 VPWR.n2674 0.179926
R4518 VPWR.n2674 VPWR.n2672 0.179926
R4519 VPWR.n3411 VPWR.n3410 0.179926
R4520 VPWR.n4009 VPWR.n4007 0.179926
R4521 VPWR.n4011 VPWR.n4009 0.179926
R4522 VPWR.n4072 VPWR.n4070 0.179926
R4523 VPWR.n733 VPWR.n731 0.179926
R4524 VPWR.n734 VPWR.n733 0.179926
R4525 VPWR.n4431 VPWR.n4429 0.179926
R4526 VPWR.n4432 VPWR.n4431 0.179926
R4527 VPWR.n4775 VPWR.n4774 0.179926
R4528 VPWR.n6106 VPWR.n6105 0.179926
R4529 VPWR.n5900 VPWR 0.168958
R4530 VPWR.n3834 VPWR.n3833 0.161711
R4531 VPWR.n2264 VPWR.n2263 0.160318
R4532 VPWR.n1964 VPWR 0.159717
R4533 VPWR.n1968 VPWR 0.159717
R4534 VPWR.n3326 VPWR 0.159717
R4535 VPWR.n3556 VPWR 0.159717
R4536 VPWR VPWR.n5113 0.159717
R4537 VPWR.n3628 VPWR 0.159628
R4538 VPWR VPWR.n1492 0.159461
R4539 VPWR.n2840 VPWR 0.158415
R4540 VPWR.n2845 VPWR 0.158415
R4541 VPWR.n2854 VPWR 0.158415
R4542 VPWR.n3305 VPWR 0.158415
R4543 VPWR.n3380 VPWR 0.158415
R4544 VPWR VPWR.n3555 0.158415
R4545 VPWR.n3900 VPWR 0.158415
R4546 VPWR.n206 VPWR 0.158415
R4547 VPWR.n2841 VPWR 0.158159
R4548 VPWR.n2858 VPWR 0.158159
R4549 VPWR.n3895 VPWR 0.158159
R4550 VPWR.n568 VPWR 0.158159
R4551 VPWR.n6094 VPWR 0.158159
R4552 VPWR VPWR.n1625 0.15779
R4553 VPWR VPWR.n3156 0.15779
R4554 VPWR VPWR.n3725 0.15779
R4555 VPWR.n3901 VPWR 0.15779
R4556 VPWR VPWR.n3934 0.15779
R4557 VPWR VPWR.n5134 0.15779
R4558 VPWR.n6105 VPWR 0.15779
R4559 VPWR.n3912 VPWR 0.156488
R4560 VPWR.n4774 VPWR 0.156488
R4561 VPWR.n2404 VPWR.n2401 0.153014
R4562 VPWR.n5845 VPWR.n5844 0.151488
R4563 VPWR.n4927 VPWR.n4926 0.151488
R4564 VPWR.n4925 VPWR.n4924 0.151488
R4565 VPWR.n4394 VPWR.n4393 0.151488
R4566 VPWR.n3790 VPWR.n3789 0.151488
R4567 VPWR.n3140 VPWR.n3139 0.151488
R4568 VPWR.n2378 VPWR.n2377 0.151488
R4569 VPWR.n5656 VPWR.n5655 0.151488
R4570 VPWR.n5292 VPWR.n5291 0.151488
R4571 VPWR.n4567 VPWR.n297 0.151488
R4572 VPWR.n1301 VPWR.n1300 0.151488
R4573 VPWR.n3457 VPWR.n3456 0.151488
R4574 VPWR.n2213 VPWR.n1578 0.151488
R4575 VPWR.n6074 VPWR.n6073 0.151488
R4576 VPWR.n630 VPWR.n629 0.151488
R4577 VPWR.n4608 VPWR.n4607 0.151488
R4578 VPWR.n1425 VPWR.n1078 0.151488
R4579 VPWR.n1442 VPWR.n1441 0.151488
R4580 VPWR.n2609 VPWR.n2608 0.151488
R4581 VPWR.n3138 VPWR.n3137 0.150166
R4582 VPWR.n3044 VPWR.n3043 0.150166
R4583 VPWR.n1776 VPWR.n1424 0.150166
R4584 VPWR VPWR.n1978 0.149301
R4585 VPWR VPWR.n1494 0.149301
R4586 VPWR.n3379 VPWR 0.149301
R4587 VPWR VPWR.n3406 0.149301
R4588 VPWR.n3823 VPWR 0.149301
R4589 VPWR VPWR.n5114 0.149301
R4590 VPWR.n220 VPWR 0.149301
R4591 VPWR VPWR.n3435 0.148676
R4592 VPWR.n5640 VPWR.n5639 0.148
R4593 VPWR VPWR.n3002 0.147999
R4594 VPWR.n2585 VPWR.n2584 0.14432
R4595 VPWR.n3127 VPWR.n3126 0.142933
R4596 VPWR.n3058 VPWR.n3057 0.142933
R4597 VPWR.n2921 VPWR.n2920 0.142933
R4598 VPWR.n2903 VPWR 0.140863
R4599 VPWR.n2998 VPWR 0.140863
R4600 VPWR VPWR.n3832 0.140863
R4601 VPWR VPWR.n702 0.140863
R4602 VPWR VPWR.n4661 0.140863
R4603 VPWR.n4951 VPWR 0.140863
R4604 VPWR VPWR.n598 0.140863
R4605 VPWR.n386 VPWR 0.140863
R4606 VPWR VPWR.n5875 0.140863
R4607 VPWR.n6200 VPWR 0.140863
R4608 VPWR.n1624 VPWR 0.140584
R4609 VPWR.n1702 VPWR 0.140584
R4610 VPWR.n1339 VPWR 0.140584
R4611 VPWR.n3484 VPWR 0.140584
R4612 VPWR.n1005 VPWR 0.140584
R4613 VPWR.n1004 VPWR 0.140584
R4614 VPWR.n4153 VPWR 0.140584
R4615 VPWR VPWR.n4401 0.140584
R4616 VPWR.n4524 VPWR 0.140584
R4617 VPWR.n4523 VPWR 0.140584
R4618 VPWR.n266 VPWR 0.140584
R4619 VPWR VPWR.n533 0.140584
R4620 VPWR.n5338 VPWR 0.140584
R4621 VPWR.n5694 VPWR 0.140584
R4622 VPWR.n5597 VPWR 0.140228
R4623 VPWR.n3793 VPWR.n3792 0.137664
R4624 VPWR.n4103 VPWR.n4102 0.137664
R4625 VPWR.n1081 VPWR.n1080 0.137664
R4626 VPWR.n3001 VPWR 0.134445
R4627 VPWR.n5823 VPWR.n5822 0.131219
R4628 VPWR.n5754 VPWR.n5753 0.131219
R4629 VPWR.n324 VPWR.n323 0.131219
R4630 VPWR.n1532 VPWR.n1530 0.120292
R4631 VPWR.n1533 VPWR.n1532 0.120292
R4632 VPWR.n1539 VPWR.n1537 0.120292
R4633 VPWR.n1538 VPWR.n1521 0.120292
R4634 VPWR.n1544 VPWR.n1521 0.120292
R4635 VPWR.n1551 VPWR.n1549 0.120292
R4636 VPWR.n1554 VPWR.n1551 0.120292
R4637 VPWR.n1556 VPWR.n1554 0.120292
R4638 VPWR.n1558 VPWR.n1556 0.120292
R4639 VPWR.n1560 VPWR.n1558 0.120292
R4640 VPWR.n1563 VPWR.n1560 0.120292
R4641 VPWR.n2820 VPWR.n2815 0.120292
R4642 VPWR.n2822 VPWR.n2820 0.120292
R4643 VPWR.n2826 VPWR.n2822 0.120292
R4644 VPWR.n2830 VPWR.n2826 0.120292
R4645 VPWR.n2832 VPWR.n2830 0.120292
R4646 VPWR.n2834 VPWR.n2832 0.120292
R4647 VPWR.n2836 VPWR.n2834 0.120292
R4648 VPWR.n2837 VPWR.n2836 0.120292
R4649 VPWR.n2862 VPWR.n2861 0.120292
R4650 VPWR.n2863 VPWR.n2862 0.120292
R4651 VPWR.n2864 VPWR.n2863 0.120292
R4652 VPWR.n2869 VPWR.n2867 0.120292
R4653 VPWR.n2871 VPWR.n2869 0.120292
R4654 VPWR.n2873 VPWR.n2871 0.120292
R4655 VPWR.n2875 VPWR.n2873 0.120292
R4656 VPWR.n2877 VPWR.n2875 0.120292
R4657 VPWR.n2879 VPWR.n2877 0.120292
R4658 VPWR.n2881 VPWR.n2879 0.120292
R4659 VPWR.n2883 VPWR.n2881 0.120292
R4660 VPWR.n2885 VPWR.n2883 0.120292
R4661 VPWR.n2887 VPWR.n2885 0.120292
R4662 VPWR.n2889 VPWR.n2887 0.120292
R4663 VPWR.n2890 VPWR.n2889 0.120292
R4664 VPWR.n2894 VPWR.n2893 0.120292
R4665 VPWR.n2899 VPWR.n2897 0.120292
R4666 VPWR.n2900 VPWR.n2899 0.120292
R4667 VPWR.n2901 VPWR.n2900 0.120292
R4668 VPWR.n2902 VPWR.n2901 0.120292
R4669 VPWR.n2732 VPWR.n2731 0.120292
R4670 VPWR.n2731 VPWR.n2730 0.120292
R4671 VPWR.n2730 VPWR.n2729 0.120292
R4672 VPWR.n2725 VPWR.n2724 0.120292
R4673 VPWR.n2724 VPWR.n2721 0.120292
R4674 VPWR.n2721 VPWR.n2719 0.120292
R4675 VPWR.n2719 VPWR.n2717 0.120292
R4676 VPWR.n2714 VPWR.n2713 0.120292
R4677 VPWR.n2713 VPWR.n2711 0.120292
R4678 VPWR.n2711 VPWR.n2709 0.120292
R4679 VPWR.n2709 VPWR.n2707 0.120292
R4680 VPWR.n2707 VPWR.n2706 0.120292
R4681 VPWR.n2706 VPWR.n2705 0.120292
R4682 VPWR.n2705 VPWR.n2703 0.120292
R4683 VPWR.n2703 VPWR.n2701 0.120292
R4684 VPWR.n2701 VPWR.n2699 0.120292
R4685 VPWR.n2699 VPWR.n2698 0.120292
R4686 VPWR.n2695 VPWR.n2694 0.120292
R4687 VPWR.n2694 VPWR.n2693 0.120292
R4688 VPWR.n2693 VPWR.n2692 0.120292
R4689 VPWR.n2689 VPWR.n2687 0.120292
R4690 VPWR.n2687 VPWR.n2686 0.120292
R4691 VPWR.n2686 VPWR.n2685 0.120292
R4692 VPWR.n2681 VPWR.n2680 0.120292
R4693 VPWR.n2680 VPWR.n2678 0.120292
R4694 VPWR.n2678 VPWR.n2676 0.120292
R4695 VPWR.n2663 VPWR.n2662 0.120292
R4696 VPWR.n2662 VPWR.n2661 0.120292
R4697 VPWR.n2661 VPWR.n2659 0.120292
R4698 VPWR.n2659 VPWR.n2657 0.120292
R4699 VPWR.n2657 VPWR.n2656 0.120292
R4700 VPWR.n2656 VPWR.n2655 0.120292
R4701 VPWR.n1660 VPWR.n1658 0.120292
R4702 VPWR.n1654 VPWR.n1611 0.120292
R4703 VPWR.n1650 VPWR.n1611 0.120292
R4704 VPWR.n1650 VPWR.n1649 0.120292
R4705 VPWR.n1649 VPWR.n1648 0.120292
R4706 VPWR.n1648 VPWR.n1613 0.120292
R4707 VPWR.n1644 VPWR.n1613 0.120292
R4708 VPWR.n1643 VPWR.n1642 0.120292
R4709 VPWR.n1642 VPWR.n1615 0.120292
R4710 VPWR.n1638 VPWR.n1615 0.120292
R4711 VPWR.n1636 VPWR.n1618 0.120292
R4712 VPWR.n1632 VPWR.n1618 0.120292
R4713 VPWR.n1628 VPWR.n1627 0.120292
R4714 VPWR.n1852 VPWR.n1850 0.120292
R4715 VPWR.n1853 VPWR.n1852 0.120292
R4716 VPWR.n1861 VPWR.n1857 0.120292
R4717 VPWR.n1862 VPWR.n1861 0.120292
R4718 VPWR.n1863 VPWR.n1862 0.120292
R4719 VPWR.n1864 VPWR.n1863 0.120292
R4720 VPWR.n1865 VPWR.n1864 0.120292
R4721 VPWR.n1871 VPWR.n1869 0.120292
R4722 VPWR.n1873 VPWR.n1871 0.120292
R4723 VPWR.n1875 VPWR.n1873 0.120292
R4724 VPWR.n1876 VPWR.n1875 0.120292
R4725 VPWR.n1882 VPWR.n1879 0.120292
R4726 VPWR.n1885 VPWR.n1882 0.120292
R4727 VPWR.n1936 VPWR.n1934 0.120292
R4728 VPWR.n1937 VPWR.n1936 0.120292
R4729 VPWR.n1943 VPWR.n1941 0.120292
R4730 VPWR.n1944 VPWR.n1943 0.120292
R4731 VPWR.n1950 VPWR.n1949 0.120292
R4732 VPWR.n1956 VPWR.n1954 0.120292
R4733 VPWR.n1958 VPWR.n1956 0.120292
R4734 VPWR.n1960 VPWR.n1958 0.120292
R4735 VPWR.n1962 VPWR.n1960 0.120292
R4736 VPWR.n1963 VPWR.n1962 0.120292
R4737 VPWR.n2023 VPWR.n2022 0.120292
R4738 VPWR.n2022 VPWR.n2021 0.120292
R4739 VPWR.n2021 VPWR.n2020 0.120292
R4740 VPWR.n2017 VPWR.n2016 0.120292
R4741 VPWR.n2016 VPWR.n2014 0.120292
R4742 VPWR.n2014 VPWR.n2012 0.120292
R4743 VPWR.n2012 VPWR.n2010 0.120292
R4744 VPWR.n2010 VPWR.n2008 0.120292
R4745 VPWR.n2008 VPWR.n2006 0.120292
R4746 VPWR.n2006 VPWR.n2004 0.120292
R4747 VPWR.n2004 VPWR.n2002 0.120292
R4748 VPWR.n2002 VPWR.n2000 0.120292
R4749 VPWR.n2000 VPWR.n1998 0.120292
R4750 VPWR.n1998 VPWR.n1996 0.120292
R4751 VPWR.n1996 VPWR.n1994 0.120292
R4752 VPWR.n1994 VPWR.n1992 0.120292
R4753 VPWR.n1992 VPWR.n1990 0.120292
R4754 VPWR.n1987 VPWR.n1986 0.120292
R4755 VPWR.n1986 VPWR.n1984 0.120292
R4756 VPWR.n1984 VPWR.n1983 0.120292
R4757 VPWR.n1983 VPWR.n1982 0.120292
R4758 VPWR.n2945 VPWR.n2944 0.120292
R4759 VPWR VPWR.n2945 0.120292
R4760 VPWR.n2950 VPWR.n2949 0.120292
R4761 VPWR.n2949 VPWR.n2948 0.120292
R4762 VPWR.n2957 VPWR.n2956 0.120292
R4763 VPWR.n2956 VPWR.n2955 0.120292
R4764 VPWR.n2966 VPWR.n2965 0.120292
R4765 VPWR.n2967 VPWR.n2966 0.120292
R4766 VPWR.n2968 VPWR.n2967 0.120292
R4767 VPWR.n2974 VPWR.n2972 0.120292
R4768 VPWR.n2976 VPWR.n2974 0.120292
R4769 VPWR.n2978 VPWR.n2976 0.120292
R4770 VPWR.n2980 VPWR.n2978 0.120292
R4771 VPWR.n2982 VPWR.n2980 0.120292
R4772 VPWR.n2985 VPWR.n2982 0.120292
R4773 VPWR.n2987 VPWR.n2985 0.120292
R4774 VPWR.n2989 VPWR.n2987 0.120292
R4775 VPWR.n2990 VPWR.n2989 0.120292
R4776 VPWR.n3026 VPWR.n3025 0.120292
R4777 VPWR.n3025 VPWR.n3024 0.120292
R4778 VPWR.n3024 VPWR.n3023 0.120292
R4779 VPWR.n3020 VPWR.n3019 0.120292
R4780 VPWR.n3019 VPWR.n3018 0.120292
R4781 VPWR.n3014 VPWR.n3013 0.120292
R4782 VPWR.n3013 VPWR.n3012 0.120292
R4783 VPWR.n3008 VPWR.n3007 0.120292
R4784 VPWR.n3003 VPWR.n2996 0.120292
R4785 VPWR.n1744 VPWR.n1742 0.120292
R4786 VPWR.n1738 VPWR.n1737 0.120292
R4787 VPWR.n1737 VPWR.n1736 0.120292
R4788 VPWR.n1736 VPWR.n1733 0.120292
R4789 VPWR.n1733 VPWR.n1731 0.120292
R4790 VPWR.n1731 VPWR.n1729 0.120292
R4791 VPWR.n1725 VPWR.n1724 0.120292
R4792 VPWR.n1724 VPWR.n1723 0.120292
R4793 VPWR.n1723 VPWR.n1720 0.120292
R4794 VPWR.n1720 VPWR.n1718 0.120292
R4795 VPWR.n1718 VPWR.n1716 0.120292
R4796 VPWR.n1713 VPWR.n1712 0.120292
R4797 VPWR VPWR.n1697 0.120292
R4798 VPWR.n1708 VPWR.n1707 0.120292
R4799 VPWR.n1707 VPWR.n1706 0.120292
R4800 VPWR.n1706 VPWR.n1705 0.120292
R4801 VPWR VPWR.n3155 0.120292
R4802 VPWR.n3166 VPWR.n3153 0.120292
R4803 VPWR.n3174 VPWR.n3153 0.120292
R4804 VPWR.n3181 VPWR.n3179 0.120292
R4805 VPWR.n3183 VPWR.n3181 0.120292
R4806 VPWR.n3185 VPWR.n3183 0.120292
R4807 VPWR.n3186 VPWR.n3185 0.120292
R4808 VPWR.n3192 VPWR.n3189 0.120292
R4809 VPWR.n3195 VPWR.n3192 0.120292
R4810 VPWR.n3275 VPWR.n3271 0.120292
R4811 VPWR.n3271 VPWR.n3269 0.120292
R4812 VPWR.n3265 VPWR.n3264 0.120292
R4813 VPWR.n3264 VPWR.n3263 0.120292
R4814 VPWR.n3258 VPWR.n3257 0.120292
R4815 VPWR.n3257 VPWR.n3256 0.120292
R4816 VPWR.n3256 VPWR.n3254 0.120292
R4817 VPWR.n3254 VPWR.n3252 0.120292
R4818 VPWR.n3252 VPWR.n3250 0.120292
R4819 VPWR.n3250 VPWR.n3248 0.120292
R4820 VPWR.n3248 VPWR.n3246 0.120292
R4821 VPWR.n3243 VPWR.n3242 0.120292
R4822 VPWR.n3242 VPWR.n3241 0.120292
R4823 VPWR.n3307 VPWR.n3306 0.120292
R4824 VPWR.n3312 VPWR.n3310 0.120292
R4825 VPWR.n3314 VPWR.n3312 0.120292
R4826 VPWR.n3316 VPWR.n3314 0.120292
R4827 VPWR.n3318 VPWR.n3316 0.120292
R4828 VPWR.n3319 VPWR.n3318 0.120292
R4829 VPWR.n3328 VPWR.n3327 0.120292
R4830 VPWR.n3333 VPWR.n3331 0.120292
R4831 VPWR.n3335 VPWR.n3333 0.120292
R4832 VPWR.n3336 VPWR.n3335 0.120292
R4833 VPWR.n3337 VPWR.n3336 0.120292
R4834 VPWR.n3338 VPWR.n3337 0.120292
R4835 VPWR.n3363 VPWR.n3362 0.120292
R4836 VPWR.n3364 VPWR.n3363 0.120292
R4837 VPWR.n3366 VPWR.n3364 0.120292
R4838 VPWR.n3367 VPWR.n3366 0.120292
R4839 VPWR.n3375 VPWR.n3374 0.120292
R4840 VPWR.n3385 VPWR.n3383 0.120292
R4841 VPWR.n3387 VPWR.n3385 0.120292
R4842 VPWR.n3433 VPWR.n3431 0.120292
R4843 VPWR.n3431 VPWR.n3430 0.120292
R4844 VPWR.n3430 VPWR.n3429 0.120292
R4845 VPWR.n3426 VPWR.n3425 0.120292
R4846 VPWR.n3425 VPWR.n3424 0.120292
R4847 VPWR.n3400 VPWR.n3399 0.120292
R4848 VPWR.n3417 VPWR.n3400 0.120292
R4849 VPWR.n3415 VPWR.n3413 0.120292
R4850 VPWR.n3413 VPWR.n3411 0.120292
R4851 VPWR.n1375 VPWR.n1373 0.120292
R4852 VPWR.n1369 VPWR.n1368 0.120292
R4853 VPWR.n1368 VPWR.n1367 0.120292
R4854 VPWR.n1367 VPWR.n1364 0.120292
R4855 VPWR.n1364 VPWR.n1362 0.120292
R4856 VPWR.n1362 VPWR.n1360 0.120292
R4857 VPWR.n1357 VPWR.n1356 0.120292
R4858 VPWR.n1356 VPWR.n1354 0.120292
R4859 VPWR.n1351 VPWR.n1350 0.120292
R4860 VPWR.n1350 VPWR.n1334 0.120292
R4861 VPWR.n1346 VPWR.n1334 0.120292
R4862 VPWR.n1345 VPWR.n1336 0.120292
R4863 VPWR.n1151 VPWR.n1150 0.120292
R4864 VPWR.n1152 VPWR.n1151 0.120292
R4865 VPWR.n1158 VPWR.n1156 0.120292
R4866 VPWR.n1160 VPWR.n1158 0.120292
R4867 VPWR.n1161 VPWR.n1160 0.120292
R4868 VPWR.n1167 VPWR.n1165 0.120292
R4869 VPWR.n1169 VPWR.n1167 0.120292
R4870 VPWR.n1171 VPWR.n1169 0.120292
R4871 VPWR.n1172 VPWR.n1171 0.120292
R4872 VPWR.n1177 VPWR.n1175 0.120292
R4873 VPWR.n1179 VPWR.n1177 0.120292
R4874 VPWR.n1181 VPWR.n1179 0.120292
R4875 VPWR.n1184 VPWR.n1181 0.120292
R4876 VPWR.n3742 VPWR.n3738 0.120292
R4877 VPWR.n3738 VPWR.n3736 0.120292
R4878 VPWR.n3732 VPWR.n3731 0.120292
R4879 VPWR.n3731 VPWR.n3730 0.120292
R4880 VPWR.n3721 VPWR.n3720 0.120292
R4881 VPWR.n3720 VPWR.n3719 0.120292
R4882 VPWR.n3719 VPWR.n3718 0.120292
R4883 VPWR.n3715 VPWR.n3714 0.120292
R4884 VPWR.n3714 VPWR.n3712 0.120292
R4885 VPWR.n3712 VPWR.n3710 0.120292
R4886 VPWR.n3706 VPWR.n1218 0.120292
R4887 VPWR.n1221 VPWR.n1218 0.120292
R4888 VPWR.n3699 VPWR.n3697 0.120292
R4889 VPWR.n3697 VPWR.n3696 0.120292
R4890 VPWR.n3696 VPWR.n3695 0.120292
R4891 VPWR.n3692 VPWR.n3691 0.120292
R4892 VPWR.n3691 VPWR.n3689 0.120292
R4893 VPWR.n3689 VPWR.n3687 0.120292
R4894 VPWR.n3687 VPWR.n3685 0.120292
R4895 VPWR.n3685 VPWR.n3684 0.120292
R4896 VPWR.n3684 VPWR.n3682 0.120292
R4897 VPWR.n3682 VPWR.n3680 0.120292
R4898 VPWR.n3680 VPWR.n3678 0.120292
R4899 VPWR.n3675 VPWR.n3674 0.120292
R4900 VPWR.n3674 VPWR.n3673 0.120292
R4901 VPWR.n3673 VPWR.n3672 0.120292
R4902 VPWR.n3668 VPWR.n3667 0.120292
R4903 VPWR.n3663 VPWR.n3662 0.120292
R4904 VPWR.n3662 VPWR.n3660 0.120292
R4905 VPWR.n3660 VPWR.n3659 0.120292
R4906 VPWR.n3659 VPWR.n3658 0.120292
R4907 VPWR.n3624 VPWR.n3623 0.120292
R4908 VPWR.n3623 VPWR.n3622 0.120292
R4909 VPWR.n3621 VPWR.n3618 0.120292
R4910 VPWR.n3618 VPWR.n3616 0.120292
R4911 VPWR.n3616 VPWR.n3614 0.120292
R4912 VPWR.n3614 VPWR.n3611 0.120292
R4913 VPWR.n3611 VPWR.n3609 0.120292
R4914 VPWR.n3609 VPWR.n3607 0.120292
R4915 VPWR.n3600 VPWR.n3598 0.120292
R4916 VPWR.n3598 VPWR.n3597 0.120292
R4917 VPWR.n3597 VPWR.n3596 0.120292
R4918 VPWR.n3593 VPWR.n3592 0.120292
R4919 VPWR.n3592 VPWR.n3591 0.120292
R4920 VPWR.n3591 VPWR.n3590 0.120292
R4921 VPWR.n3586 VPWR.n3585 0.120292
R4922 VPWR.n3585 VPWR.n3584 0.120292
R4923 VPWR.n3584 VPWR.n3583 0.120292
R4924 VPWR.n3579 VPWR.n1272 0.120292
R4925 VPWR.n3577 VPWR.n3575 0.120292
R4926 VPWR.n3575 VPWR.n3574 0.120292
R4927 VPWR.n3574 VPWR.n3573 0.120292
R4928 VPWR.n3569 VPWR.n3568 0.120292
R4929 VPWR.n3568 VPWR.n3567 0.120292
R4930 VPWR.n3567 VPWR.n3566 0.120292
R4931 VPWR.n3563 VPWR.n3562 0.120292
R4932 VPWR.n3562 VPWR.n3560 0.120292
R4933 VPWR.n3560 VPWR.n3558 0.120292
R4934 VPWR.n3525 VPWR.n3523 0.120292
R4935 VPWR.n3523 VPWR.n3521 0.120292
R4936 VPWR.n3521 VPWR.n3519 0.120292
R4937 VPWR.n3516 VPWR.n3515 0.120292
R4938 VPWR.n3515 VPWR.n3513 0.120292
R4939 VPWR.n3513 VPWR.n3512 0.120292
R4940 VPWR.n3512 VPWR.n3510 0.120292
R4941 VPWR.n3510 VPWR.n3508 0.120292
R4942 VPWR.n3508 VPWR.n3506 0.120292
R4943 VPWR.n3506 VPWR.n3504 0.120292
R4944 VPWR.n3501 VPWR.n3500 0.120292
R4945 VPWR.n3500 VPWR.n3477 0.120292
R4946 VPWR.n3496 VPWR.n3477 0.120292
R4947 VPWR.n3495 VPWR.n3479 0.120292
R4948 VPWR.n3491 VPWR.n3479 0.120292
R4949 VPWR.n3491 VPWR.n3490 0.120292
R4950 VPWR.n3490 VPWR.n3489 0.120292
R4951 VPWR.n3486 VPWR.n3485 0.120292
R4952 VPWR.n3820 VPWR.n3818 0.120292
R4953 VPWR.n3821 VPWR.n3820 0.120292
R4954 VPWR.n3826 VPWR.n3825 0.120292
R4955 VPWR.n3827 VPWR.n3826 0.120292
R4956 VPWR.n3828 VPWR.n3827 0.120292
R4957 VPWR.n3889 VPWR.n3887 0.120292
R4958 VPWR.n3891 VPWR.n3889 0.120292
R4959 VPWR.n3893 VPWR.n3891 0.120292
R4960 VPWR.n3908 VPWR.n3907 0.120292
R4961 VPWR.n3916 VPWR.n3915 0.120292
R4962 VPWR.n3917 VPWR.n3916 0.120292
R4963 VPWR.n3918 VPWR.n3917 0.120292
R4964 VPWR.n3969 VPWR.n3968 0.120292
R4965 VPWR.n3968 VPWR.n3966 0.120292
R4966 VPWR.n3966 VPWR.n3964 0.120292
R4967 VPWR.n3964 VPWR.n3963 0.120292
R4968 VPWR.n3963 VPWR.n3962 0.120292
R4969 VPWR.n3959 VPWR.n3958 0.120292
R4970 VPWR.n3958 VPWR.n3956 0.120292
R4971 VPWR.n3956 VPWR 0.120292
R4972 VPWR.n3953 VPWR.n3952 0.120292
R4973 VPWR.n3952 VPWR.n3951 0.120292
R4974 VPWR.n3951 VPWR.n3950 0.120292
R4975 VPWR.n3945 VPWR.n3944 0.120292
R4976 VPWR.n3944 VPWR.n3943 0.120292
R4977 VPWR.n3935 VPWR.n3932 0.120292
R4978 VPWR.n3995 VPWR.n3993 0.120292
R4979 VPWR.n3997 VPWR.n3995 0.120292
R4980 VPWR.n3998 VPWR.n3997 0.120292
R4981 VPWR.n4003 VPWR.n4001 0.120292
R4982 VPWR.n4005 VPWR.n4003 0.120292
R4983 VPWR.n4007 VPWR.n4005 0.120292
R4984 VPWR.n4018 VPWR.n4016 0.120292
R4985 VPWR.n4020 VPWR.n4018 0.120292
R4986 VPWR.n4022 VPWR.n4020 0.120292
R4987 VPWR.n4024 VPWR.n4022 0.120292
R4988 VPWR.n4026 VPWR.n4024 0.120292
R4989 VPWR.n4028 VPWR.n4026 0.120292
R4990 VPWR.n4029 VPWR.n4028 0.120292
R4991 VPWR.n4080 VPWR.n4079 0.120292
R4992 VPWR.n4079 VPWR.n4078 0.120292
R4993 VPWR.n4076 VPWR.n4074 0.120292
R4994 VPWR.n4074 VPWR.n4072 0.120292
R4995 VPWR.n4068 VPWR.n4067 0.120292
R4996 VPWR.n4067 VPWR.n4066 0.120292
R4997 VPWR.n4062 VPWR.n4061 0.120292
R4998 VPWR.n4061 VPWR.n4060 0.120292
R4999 VPWR.n4057 VPWR.n4056 0.120292
R5000 VPWR.n4056 VPWR.n4054 0.120292
R5001 VPWR.n4054 VPWR.n4053 0.120292
R5002 VPWR.n4053 VPWR.n4051 0.120292
R5003 VPWR.n4051 VPWR 0.120292
R5004 VPWR.n4046 VPWR.n4045 0.120292
R5005 VPWR.n4045 VPWR.n4044 0.120292
R5006 VPWR.n4044 VPWR.n4043 0.120292
R5007 VPWR.n1039 VPWR.n1037 0.120292
R5008 VPWR.n1034 VPWR.n1033 0.120292
R5009 VPWR.n1033 VPWR.n1031 0.120292
R5010 VPWR.n1031 VPWR 0.120292
R5011 VPWR.n1027 VPWR.n1026 0.120292
R5012 VPWR.n1026 VPWR.n1025 0.120292
R5013 VPWR.n1025 VPWR.n1024 0.120292
R5014 VPWR.n1021 VPWR.n1020 0.120292
R5015 VPWR.n1020 VPWR.n1018 0.120292
R5016 VPWR.n1018 VPWR 0.120292
R5017 VPWR.n1014 VPWR.n1013 0.120292
R5018 VPWR.n1013 VPWR.n1012 0.120292
R5019 VPWR.n1012 VPWR.n1011 0.120292
R5020 VPWR.n1007 VPWR.n1006 0.120292
R5021 VPWR.n713 VPWR.n711 0.120292
R5022 VPWR.n715 VPWR.n713 0.120292
R5023 VPWR.n719 VPWR.n715 0.120292
R5024 VPWR.n721 VPWR.n720 0.120292
R5025 VPWR.n722 VPWR.n721 0.120292
R5026 VPWR.n727 VPWR.n725 0.120292
R5027 VPWR.n729 VPWR.n727 0.120292
R5028 VPWR.n731 VPWR.n729 0.120292
R5029 VPWR.n740 VPWR.n737 0.120292
R5030 VPWR.n743 VPWR.n740 0.120292
R5031 VPWR.n864 VPWR.n862 0.120292
R5032 VPWR.n865 VPWR.n864 0.120292
R5033 VPWR.n877 VPWR.n824 0.120292
R5034 VPWR.n878 VPWR.n877 0.120292
R5035 VPWR.n879 VPWR.n878 0.120292
R5036 VPWR.n885 VPWR.n884 0.120292
R5037 VPWR.n891 VPWR.n889 0.120292
R5038 VPWR.n893 VPWR.n891 0.120292
R5039 VPWR.n895 VPWR.n893 0.120292
R5040 VPWR.n901 VPWR.n900 0.120292
R5041 VPWR.n902 VPWR.n901 0.120292
R5042 VPWR.n903 VPWR.n902 0.120292
R5043 VPWR.n908 VPWR.n906 0.120292
R5044 VPWR.n910 VPWR.n908 0.120292
R5045 VPWR.n912 VPWR.n910 0.120292
R5046 VPWR.n913 VPWR.n912 0.120292
R5047 VPWR.n918 VPWR.n815 0.120292
R5048 VPWR.n925 VPWR.n923 0.120292
R5049 VPWR.n926 VPWR.n925 0.120292
R5050 VPWR.n927 VPWR.n926 0.120292
R5051 VPWR.n928 VPWR.n927 0.120292
R5052 VPWR.n933 VPWR.n931 0.120292
R5053 VPWR.n935 VPWR.n933 0.120292
R5054 VPWR.n936 VPWR.n935 0.120292
R5055 VPWR.n937 VPWR.n936 0.120292
R5056 VPWR.n941 VPWR.n940 0.120292
R5057 VPWR.n942 VPWR.n941 0.120292
R5058 VPWR.n947 VPWR.n942 0.120292
R5059 VPWR.n4238 VPWR.n4237 0.120292
R5060 VPWR.n4237 VPWR.n4236 0.120292
R5061 VPWR.n4248 VPWR.n4247 0.120292
R5062 VPWR.n4249 VPWR.n4248 0.120292
R5063 VPWR.n4251 VPWR.n4249 0.120292
R5064 VPWR.n4257 VPWR.n4255 0.120292
R5065 VPWR.n4260 VPWR.n4257 0.120292
R5066 VPWR.n4262 VPWR.n4260 0.120292
R5067 VPWR.n4264 VPWR.n4262 0.120292
R5068 VPWR.n4265 VPWR.n4264 0.120292
R5069 VPWR.n4271 VPWR.n4268 0.120292
R5070 VPWR.n4273 VPWR.n4271 0.120292
R5071 VPWR.n4275 VPWR.n4273 0.120292
R5072 VPWR.n4276 VPWR.n4275 0.120292
R5073 VPWR.n4283 VPWR.n4282 0.120292
R5074 VPWR.n4284 VPWR.n4283 0.120292
R5075 VPWR.n4289 VPWR.n4284 0.120292
R5076 VPWR.n4293 VPWR.n4292 0.120292
R5077 VPWR.n4298 VPWR.n4296 0.120292
R5078 VPWR.n4301 VPWR.n4298 0.120292
R5079 VPWR.n4303 VPWR.n4301 0.120292
R5080 VPWR.n4305 VPWR.n4303 0.120292
R5081 VPWR.n4306 VPWR.n4305 0.120292
R5082 VPWR.n4307 VPWR.n4306 0.120292
R5083 VPWR.n4308 VPWR.n4307 0.120292
R5084 VPWR.n4313 VPWR.n4311 0.120292
R5085 VPWR.n4315 VPWR.n4313 0.120292
R5086 VPWR.n4317 VPWR.n4315 0.120292
R5087 VPWR.n4319 VPWR.n4317 0.120292
R5088 VPWR.n4320 VPWR.n4319 0.120292
R5089 VPWR.n4321 VPWR.n4320 0.120292
R5090 VPWR.n4322 VPWR.n4321 0.120292
R5091 VPWR.n4327 VPWR.n4326 0.120292
R5092 VPWR.n4328 VPWR.n4327 0.120292
R5093 VPWR.n4329 VPWR.n4328 0.120292
R5094 VPWR.n4337 VPWR.n4336 0.120292
R5095 VPWR.n4338 VPWR.n4337 0.120292
R5096 VPWR.n4199 VPWR.n4197 0.120292
R5097 VPWR.n4191 VPWR.n4186 0.120292
R5098 VPWR.n4186 VPWR.n4185 0.120292
R5099 VPWR.n4185 VPWR.n4184 0.120292
R5100 VPWR.n4180 VPWR.n4179 0.120292
R5101 VPWR.n4179 VPWR.n4177 0.120292
R5102 VPWR.n4177 VPWR.n4174 0.120292
R5103 VPWR.n4174 VPWR.n4172 0.120292
R5104 VPWR.n4172 VPWR.n4170 0.120292
R5105 VPWR.n4167 VPWR.n4166 0.120292
R5106 VPWR.n4166 VPWR.n4165 0.120292
R5107 VPWR.n4165 VPWR.n4163 0.120292
R5108 VPWR.n4163 VPWR.n4160 0.120292
R5109 VPWR.n4160 VPWR.n4158 0.120292
R5110 VPWR.n4158 VPWR.n4156 0.120292
R5111 VPWR.n4411 VPWR.n4409 0.120292
R5112 VPWR.n4413 VPWR.n4411 0.120292
R5113 VPWR.n4417 VPWR.n4413 0.120292
R5114 VPWR.n4419 VPWR.n4418 0.120292
R5115 VPWR.n4420 VPWR.n4419 0.120292
R5116 VPWR.n4425 VPWR.n4423 0.120292
R5117 VPWR.n4427 VPWR.n4425 0.120292
R5118 VPWR.n4429 VPWR.n4427 0.120292
R5119 VPWR.n4438 VPWR.n4435 0.120292
R5120 VPWR.n4441 VPWR.n4438 0.120292
R5121 VPWR.n4878 VPWR.n4877 0.120292
R5122 VPWR.n4877 VPWR.n4875 0.120292
R5123 VPWR.n4870 VPWR.n4865 0.120292
R5124 VPWR.n4865 VPWR.n4864 0.120292
R5125 VPWR.n4864 VPWR.n4863 0.120292
R5126 VPWR.n4859 VPWR.n4858 0.120292
R5127 VPWR.n4858 VPWR.n4855 0.120292
R5128 VPWR.n4855 VPWR.n4853 0.120292
R5129 VPWR.n4853 VPWR.n4851 0.120292
R5130 VPWR.n4848 VPWR.n4847 0.120292
R5131 VPWR.n4847 VPWR.n4844 0.120292
R5132 VPWR.n4844 VPWR.n4842 0.120292
R5133 VPWR.n4842 VPWR.n4840 0.120292
R5134 VPWR.n4836 VPWR.n4835 0.120292
R5135 VPWR.n4663 VPWR.n4662 0.120292
R5136 VPWR.n4664 VPWR.n4663 0.120292
R5137 VPWR.n4669 VPWR.n4667 0.120292
R5138 VPWR.n4671 VPWR.n4669 0.120292
R5139 VPWR.n4673 VPWR.n4671 0.120292
R5140 VPWR.n4675 VPWR.n4673 0.120292
R5141 VPWR.n4677 VPWR.n4675 0.120292
R5142 VPWR.n4679 VPWR.n4677 0.120292
R5143 VPWR.n4680 VPWR.n4679 0.120292
R5144 VPWR.n4685 VPWR.n4683 0.120292
R5145 VPWR.n4688 VPWR.n4687 0.120292
R5146 VPWR.n4689 VPWR.n4688 0.120292
R5147 VPWR.n4696 VPWR.n4695 0.120292
R5148 VPWR.n4722 VPWR.n4720 0.120292
R5149 VPWR.n4724 VPWR.n4722 0.120292
R5150 VPWR.n4725 VPWR.n4724 0.120292
R5151 VPWR.n4732 VPWR.n4731 0.120292
R5152 VPWR.n4733 VPWR.n4732 0.120292
R5153 VPWR.n4734 VPWR.n4733 0.120292
R5154 VPWR.n4739 VPWR.n4737 0.120292
R5155 VPWR.n4740 VPWR.n4739 0.120292
R5156 VPWR VPWR.n4740 0.120292
R5157 VPWR.n4747 VPWR.n4746 0.120292
R5158 VPWR.n4748 VPWR.n4747 0.120292
R5159 VPWR.n4749 VPWR.n4748 0.120292
R5160 VPWR.n4754 VPWR.n4752 0.120292
R5161 VPWR.n4756 VPWR.n4754 0.120292
R5162 VPWR.n4759 VPWR.n4756 0.120292
R5163 VPWR.n4761 VPWR.n4759 0.120292
R5164 VPWR.n4763 VPWR.n4761 0.120292
R5165 VPWR.n4765 VPWR.n4763 0.120292
R5166 VPWR.n4770 VPWR.n4769 0.120292
R5167 VPWR.n4777 VPWR.n4775 0.120292
R5168 VPWR.n4779 VPWR.n4777 0.120292
R5169 VPWR.n4780 VPWR.n4779 0.120292
R5170 VPWR.n4785 VPWR.n4783 0.120292
R5171 VPWR.n4787 VPWR.n4785 0.120292
R5172 VPWR.n4789 VPWR.n4582 0.120292
R5173 VPWR.n4793 VPWR.n4582 0.120292
R5174 VPWR.n4802 VPWR.n4800 0.120292
R5175 VPWR.n4803 VPWR.n4802 0.120292
R5176 VPWR.n4804 VPWR.n4803 0.120292
R5177 VPWR.n4805 VPWR.n4804 0.120292
R5178 VPWR.n4558 VPWR.n4557 0.120292
R5179 VPWR.n4557 VPWR.n4556 0.120292
R5180 VPWR.n4556 VPWR.n4554 0.120292
R5181 VPWR.n4553 VPWR.n4548 0.120292
R5182 VPWR.n4548 VPWR.n4547 0.120292
R5183 VPWR.n4547 VPWR.n4546 0.120292
R5184 VPWR.n4542 VPWR.n4541 0.120292
R5185 VPWR.n4541 VPWR.n4539 0.120292
R5186 VPWR.n4539 VPWR.n4537 0.120292
R5187 VPWR.n4537 VPWR.n4535 0.120292
R5188 VPWR.n4535 VPWR.n4532 0.120292
R5189 VPWR.n4532 VPWR.n4530 0.120292
R5190 VPWR.n4530 VPWR.n4528 0.120292
R5191 VPWR.n4946 VPWR.n4944 0.120292
R5192 VPWR.n4957 VPWR.n4944 0.120292
R5193 VPWR.n4965 VPWR.n4964 0.120292
R5194 VPWR.n4966 VPWR.n4965 0.120292
R5195 VPWR.n4972 VPWR.n4970 0.120292
R5196 VPWR.n4973 VPWR.n4972 0.120292
R5197 VPWR.n4978 VPWR.n4977 0.120292
R5198 VPWR.n4984 VPWR.n4982 0.120292
R5199 VPWR.n4988 VPWR.n4984 0.120292
R5200 VPWR.n5050 VPWR.n5049 0.120292
R5201 VPWR.n5051 VPWR.n5050 0.120292
R5202 VPWR.n5054 VPWR.n5051 0.120292
R5203 VPWR.n5056 VPWR.n5054 0.120292
R5204 VPWR.n5057 VPWR.n5056 0.120292
R5205 VPWR.n5065 VPWR.n5062 0.120292
R5206 VPWR.n5067 VPWR.n5065 0.120292
R5207 VPWR.n5069 VPWR.n5067 0.120292
R5208 VPWR.n5070 VPWR.n5069 0.120292
R5209 VPWR.n5075 VPWR.n5073 0.120292
R5210 VPWR.n5077 VPWR.n5075 0.120292
R5211 VPWR.n5079 VPWR.n5077 0.120292
R5212 VPWR.n5081 VPWR.n5079 0.120292
R5213 VPWR.n5083 VPWR.n5081 0.120292
R5214 VPWR.n5084 VPWR.n5083 0.120292
R5215 VPWR.n5090 VPWR.n5089 0.120292
R5216 VPWR.n5091 VPWR.n5090 0.120292
R5217 VPWR.n5093 VPWR.n5091 0.120292
R5218 VPWR.n5095 VPWR.n5093 0.120292
R5219 VPWR.n5096 VPWR.n5095 0.120292
R5220 VPWR.n5141 VPWR.n5140 0.120292
R5221 VPWR.n5139 VPWR.n5138 0.120292
R5222 VPWR.n5128 VPWR.n5104 0.120292
R5223 VPWR.n5126 VPWR.n5125 0.120292
R5224 VPWR.n5125 VPWR.n5124 0.120292
R5225 VPWR.n5119 VPWR.n5118 0.120292
R5226 VPWR.n5164 VPWR.n5163 0.120292
R5227 VPWR.n5169 VPWR.n5167 0.120292
R5228 VPWR.n5170 VPWR.n5169 0.120292
R5229 VPWR.n5172 VPWR.n5171 0.120292
R5230 VPWR.n5185 VPWR.n5184 0.120292
R5231 VPWR.n5186 VPWR.n5185 0.120292
R5232 VPWR.n5187 VPWR.n5186 0.120292
R5233 VPWR.n5192 VPWR.n5190 0.120292
R5234 VPWR.n5194 VPWR.n5192 0.120292
R5235 VPWR.n5196 VPWR.n5194 0.120292
R5236 VPWR.n5198 VPWR.n5196 0.120292
R5237 VPWR.n5200 VPWR.n5198 0.120292
R5238 VPWR.n5202 VPWR.n5200 0.120292
R5239 VPWR.n5203 VPWR.n5202 0.120292
R5240 VPWR.n5210 VPWR.n5209 0.120292
R5241 VPWR.n5211 VPWR.n5210 0.120292
R5242 VPWR.n5212 VPWR.n5211 0.120292
R5243 VPWR.n5265 VPWR.n5264 0.120292
R5244 VPWR.n5264 VPWR.n5263 0.120292
R5245 VPWR.n5263 VPWR.n5262 0.120292
R5246 VPWR.n5262 VPWR.n5260 0.120292
R5247 VPWR.n5255 VPWR.n5254 0.120292
R5248 VPWR.n5254 VPWR.n5252 0.120292
R5249 VPWR.n5252 VPWR.n5250 0.120292
R5250 VPWR.n5250 VPWR.n5249 0.120292
R5251 VPWR.n5246 VPWR.n5245 0.120292
R5252 VPWR.n5241 VPWR.n5240 0.120292
R5253 VPWR.n5240 VPWR.n5239 0.120292
R5254 VPWR.n5239 VPWR.n5238 0.120292
R5255 VPWR.n5226 VPWR.n5225 0.120292
R5256 VPWR.n5233 VPWR.n5226 0.120292
R5257 VPWR.n5231 VPWR.n5229 0.120292
R5258 VPWR.n5229 VPWR.n5228 0.120292
R5259 VPWR.n5228 VPWR.n5227 0.120292
R5260 VPWR.n292 VPWR.n290 0.120292
R5261 VPWR.n290 VPWR.n288 0.120292
R5262 VPWR.n288 VPWR.n286 0.120292
R5263 VPWR.n283 VPWR.n282 0.120292
R5264 VPWR.n282 VPWR.n281 0.120292
R5265 VPWR.n281 VPWR.n279 0.120292
R5266 VPWR.n273 VPWR.n272 0.120292
R5267 VPWR.n272 VPWR.n270 0.120292
R5268 VPWR.n201 VPWR.n200 0.120292
R5269 VPWR VPWR.n201 0.120292
R5270 VPWR.n205 VPWR.n204 0.120292
R5271 VPWR.n209 VPWR.n208 0.120292
R5272 VPWR.n210 VPWR.n209 0.120292
R5273 VPWR.n538 VPWR.n537 0.120292
R5274 VPWR.n548 VPWR.n547 0.120292
R5275 VPWR.n550 VPWR.n548 0.120292
R5276 VPWR.n553 VPWR.n552 0.120292
R5277 VPWR.n552 VPWR.n551 0.120292
R5278 VPWR.n561 VPWR.n560 0.120292
R5279 VPWR.n560 VPWR.n559 0.120292
R5280 VPWR.n576 VPWR.n575 0.120292
R5281 VPWR.n581 VPWR.n580 0.120292
R5282 VPWR.n582 VPWR.n581 0.120292
R5283 VPWR.n583 VPWR.n582 0.120292
R5284 VPWR.n592 VPWR.n591 0.120292
R5285 VPWR.n593 VPWR.n592 0.120292
R5286 VPWR.n597 VPWR.n593 0.120292
R5287 VPWR.n600 VPWR.n599 0.120292
R5288 VPWR.n601 VPWR.n600 0.120292
R5289 VPWR.n605 VPWR.n604 0.120292
R5290 VPWR.n609 VPWR.n608 0.120292
R5291 VPWR.n610 VPWR.n609 0.120292
R5292 VPWR.n615 VPWR.n610 0.120292
R5293 VPWR.n459 VPWR.n455 0.120292
R5294 VPWR.n455 VPWR.n453 0.120292
R5295 VPWR.n450 VPWR.n449 0.120292
R5296 VPWR.n449 VPWR.n448 0.120292
R5297 VPWR.n448 VPWR.n446 0.120292
R5298 VPWR.n446 VPWR.n444 0.120292
R5299 VPWR.n444 VPWR.n442 0.120292
R5300 VPWR.n442 VPWR.n440 0.120292
R5301 VPWR.n440 VPWR.n438 0.120292
R5302 VPWR.n435 VPWR.n434 0.120292
R5303 VPWR.n434 VPWR.n433 0.120292
R5304 VPWR.n433 VPWR.n432 0.120292
R5305 VPWR.n428 VPWR.n355 0.120292
R5306 VPWR.n356 VPWR.n355 0.120292
R5307 VPWR.n422 VPWR.n421 0.120292
R5308 VPWR.n421 VPWR.n358 0.120292
R5309 VPWR.n416 VPWR.n358 0.120292
R5310 VPWR.n416 VPWR.n415 0.120292
R5311 VPWR.n415 VPWR.n414 0.120292
R5312 VPWR.n411 VPWR.n360 0.120292
R5313 VPWR.n406 VPWR.n360 0.120292
R5314 VPWR.n406 VPWR.n405 0.120292
R5315 VPWR.n404 VPWR.n403 0.120292
R5316 VPWR.n403 VPWR.n363 0.120292
R5317 VPWR VPWR.n363 0.120292
R5318 VPWR.n398 VPWR.n397 0.120292
R5319 VPWR.n397 VPWR.n365 0.120292
R5320 VPWR.n393 VPWR.n365 0.120292
R5321 VPWR.n391 VPWR.n367 0.120292
R5322 VPWR.n382 VPWR.n381 0.120292
R5323 VPWR.n381 VPWR 0.120292
R5324 VPWR.n377 VPWR.n376 0.120292
R5325 VPWR.n376 VPWR.n375 0.120292
R5326 VPWR.n5373 VPWR.n5371 0.120292
R5327 VPWR.n5368 VPWR.n5367 0.120292
R5328 VPWR.n5367 VPWR.n5365 0.120292
R5329 VPWR.n5365 VPWR 0.120292
R5330 VPWR.n5361 VPWR.n5360 0.120292
R5331 VPWR.n5360 VPWR.n5359 0.120292
R5332 VPWR.n5359 VPWR.n5358 0.120292
R5333 VPWR.n5358 VPWR.n5356 0.120292
R5334 VPWR.n5356 VPWR.n5354 0.120292
R5335 VPWR.n5350 VPWR.n5349 0.120292
R5336 VPWR.n5347 VPWR.n5333 0.120292
R5337 VPWR.n5341 VPWR.n5340 0.120292
R5338 VPWR.n5340 VPWR.n5339 0.120292
R5339 VPWR.n5869 VPWR.n5868 0.120292
R5340 VPWR.n5870 VPWR.n5869 0.120292
R5341 VPWR.n5880 VPWR.n5879 0.120292
R5342 VPWR.n5890 VPWR.n5886 0.120292
R5343 VPWR.n5891 VPWR.n5890 0.120292
R5344 VPWR.n5892 VPWR.n5891 0.120292
R5345 VPWR.n5893 VPWR.n5892 0.120292
R5346 VPWR.n5899 VPWR.n5893 0.120292
R5347 VPWR.n5970 VPWR.n5965 0.120292
R5348 VPWR.n5978 VPWR.n5977 0.120292
R5349 VPWR.n5984 VPWR.n5983 0.120292
R5350 VPWR.n5985 VPWR.n5984 0.120292
R5351 VPWR.n5986 VPWR.n5985 0.120292
R5352 VPWR.n5992 VPWR.n5990 0.120292
R5353 VPWR.n5995 VPWR.n5992 0.120292
R5354 VPWR.n5997 VPWR.n5995 0.120292
R5355 VPWR.n5999 VPWR.n5997 0.120292
R5356 VPWR.n6000 VPWR.n5999 0.120292
R5357 VPWR.n6008 VPWR.n6007 0.120292
R5358 VPWR.n6009 VPWR.n6008 0.120292
R5359 VPWR.n6012 VPWR.n6009 0.120292
R5360 VPWR.n6015 VPWR.n6013 0.120292
R5361 VPWR.n6017 VPWR.n6015 0.120292
R5362 VPWR.n6018 VPWR.n6017 0.120292
R5363 VPWR.n6024 VPWR.n6022 0.120292
R5364 VPWR.n6026 VPWR.n6024 0.120292
R5365 VPWR.n6029 VPWR.n6026 0.120292
R5366 VPWR.n6031 VPWR.n6029 0.120292
R5367 VPWR.n6032 VPWR.n6031 0.120292
R5368 VPWR.n6037 VPWR.n6035 0.120292
R5369 VPWR.n6039 VPWR.n6037 0.120292
R5370 VPWR.n6041 VPWR.n6039 0.120292
R5371 VPWR.n6043 VPWR.n6041 0.120292
R5372 VPWR.n6045 VPWR.n6043 0.120292
R5373 VPWR.n6047 VPWR.n6045 0.120292
R5374 VPWR.n6048 VPWR.n6047 0.120292
R5375 VPWR.n6055 VPWR.n6052 0.120292
R5376 VPWR.n6056 VPWR.n6055 0.120292
R5377 VPWR.n5462 VPWR.n5461 0.120292
R5378 VPWR.n5467 VPWR.n5465 0.120292
R5379 VPWR.n5469 VPWR.n5467 0.120292
R5380 VPWR.n5471 VPWR.n5469 0.120292
R5381 VPWR.n5473 VPWR.n5471 0.120292
R5382 VPWR.n5475 VPWR.n5473 0.120292
R5383 VPWR.n5477 VPWR.n5475 0.120292
R5384 VPWR.n5478 VPWR.n5477 0.120292
R5385 VPWR.n5484 VPWR.n5481 0.120292
R5386 VPWR.n5486 VPWR.n5484 0.120292
R5387 VPWR.n5487 VPWR.n5486 0.120292
R5388 VPWR.n5493 VPWR.n5491 0.120292
R5389 VPWR.n5495 VPWR.n5493 0.120292
R5390 VPWR.n5500 VPWR.n5498 0.120292
R5391 VPWR.n5502 VPWR.n5500 0.120292
R5392 VPWR.n5503 VPWR.n5502 0.120292
R5393 VPWR.n5511 VPWR.n5510 0.120292
R5394 VPWR.n5512 VPWR.n5511 0.120292
R5395 VPWR.n5514 VPWR.n5512 0.120292
R5396 VPWR.n5518 VPWR.n5516 0.120292
R5397 VPWR.n5520 VPWR.n5518 0.120292
R5398 VPWR.n5522 VPWR.n5520 0.120292
R5399 VPWR.n5523 VPWR.n5522 0.120292
R5400 VPWR.n5528 VPWR.n5527 0.120292
R5401 VPWR.n5534 VPWR.n5533 0.120292
R5402 VPWR.n5535 VPWR.n5534 0.120292
R5403 VPWR.n5536 VPWR.n5535 0.120292
R5404 VPWR.n5541 VPWR.n5539 0.120292
R5405 VPWR.n5543 VPWR.n5541 0.120292
R5406 VPWR.n5544 VPWR.n5543 0.120292
R5407 VPWR.n5549 VPWR.n5547 0.120292
R5408 VPWR.n5552 VPWR.n5549 0.120292
R5409 VPWR.n5553 VPWR.n5552 0.120292
R5410 VPWR.n5738 VPWR.n5736 0.120292
R5411 VPWR.n5736 VPWR.n5733 0.120292
R5412 VPWR.n5733 VPWR.n5731 0.120292
R5413 VPWR.n5731 VPWR.n5729 0.120292
R5414 VPWR.n5725 VPWR.n5724 0.120292
R5415 VPWR.n5724 VPWR.n5722 0.120292
R5416 VPWR.n5717 VPWR.n5709 0.120292
R5417 VPWR.n5709 VPWR.n5708 0.120292
R5418 VPWR.n5708 VPWR.n5707 0.120292
R5419 VPWR.n5707 VPWR.n5706 0.120292
R5420 VPWR.n5706 VPWR.n5704 0.120292
R5421 VPWR.n5701 VPWR.n5700 0.120292
R5422 VPWR.n5700 VPWR.n5698 0.120292
R5423 VPWR.n2406 VPWR.n2404 0.120292
R5424 VPWR.n2407 VPWR.n2406 0.120292
R5425 VPWR.n2408 VPWR.n2407 0.120292
R5426 VPWR.n2409 VPWR.n2408 0.120292
R5427 VPWR.n2414 VPWR.n2412 0.120292
R5428 VPWR.n2415 VPWR.n2414 0.120292
R5429 VPWR VPWR.n2415 0.120292
R5430 VPWR.n2419 VPWR.n2418 0.120292
R5431 VPWR.n2420 VPWR.n2419 0.120292
R5432 VPWR.n2421 VPWR.n2420 0.120292
R5433 VPWR.n2426 VPWR.n2424 0.120292
R5434 VPWR.n2427 VPWR.n2426 0.120292
R5435 VPWR VPWR.n2427 0.120292
R5436 VPWR.n2432 VPWR.n2430 0.120292
R5437 VPWR.n2434 VPWR.n2432 0.120292
R5438 VPWR.n2435 VPWR.n2434 0.120292
R5439 VPWR.n2436 VPWR.n2435 0.120292
R5440 VPWR.n2437 VPWR.n2436 0.120292
R5441 VPWR.n2486 VPWR.n2484 0.120292
R5442 VPWR.n2487 VPWR.n2486 0.120292
R5443 VPWR VPWR.n2487 0.120292
R5444 VPWR.n2497 VPWR.n2496 0.120292
R5445 VPWR.n2498 VPWR.n2497 0.120292
R5446 VPWR.n2500 VPWR.n2498 0.120292
R5447 VPWR.n2504 VPWR.n2500 0.120292
R5448 VPWR.n2508 VPWR.n2504 0.120292
R5449 VPWR.n2510 VPWR.n2508 0.120292
R5450 VPWR.n2512 VPWR.n2510 0.120292
R5451 VPWR.n2514 VPWR.n2512 0.120292
R5452 VPWR.n2516 VPWR.n2514 0.120292
R5453 VPWR.n2518 VPWR.n2516 0.120292
R5454 VPWR.n2519 VPWR.n2518 0.120292
R5455 VPWR.n2524 VPWR.n2522 0.120292
R5456 VPWR.n2526 VPWR.n2524 0.120292
R5457 VPWR.n2529 VPWR.n2526 0.120292
R5458 VPWR.n2531 VPWR.n2529 0.120292
R5459 VPWR.n2533 VPWR.n2531 0.120292
R5460 VPWR.n2534 VPWR.n2533 0.120292
R5461 VPWR.n2542 VPWR.n2541 0.120292
R5462 VPWR.n2543 VPWR.n2542 0.120292
R5463 VPWR.n2544 VPWR.n2543 0.120292
R5464 VPWR.n2550 VPWR.n2548 0.120292
R5465 VPWR.n2552 VPWR.n2550 0.120292
R5466 VPWR.n2553 VPWR.n2552 0.120292
R5467 VPWR.n2554 VPWR.n2553 0.120292
R5468 VPWR.n2555 VPWR.n2554 0.120292
R5469 VPWR.n2561 VPWR.n2559 0.120292
R5470 VPWR.n2563 VPWR.n2561 0.120292
R5471 VPWR.n2565 VPWR.n2563 0.120292
R5472 VPWR.n2567 VPWR.n2565 0.120292
R5473 VPWR.n2569 VPWR.n2567 0.120292
R5474 VPWR.n2571 VPWR.n2569 0.120292
R5475 VPWR.n2572 VPWR.n2571 0.120292
R5476 VPWR.n2578 VPWR.n2575 0.120292
R5477 VPWR.n2583 VPWR.n2578 0.120292
R5478 VPWR.n2586 VPWR.n2583 0.120292
R5479 VPWR.n2588 VPWR.n2586 0.120292
R5480 VPWR.n2589 VPWR.n2588 0.120292
R5481 VPWR.n2590 VPWR.n2589 0.120292
R5482 VPWR.n2591 VPWR.n2590 0.120292
R5483 VPWR.n2116 VPWR.n2114 0.120292
R5484 VPWR.n2117 VPWR.n2116 0.120292
R5485 VPWR VPWR.n2117 0.120292
R5486 VPWR.n2124 VPWR.n2123 0.120292
R5487 VPWR.n2125 VPWR.n2124 0.120292
R5488 VPWR.n2126 VPWR.n2125 0.120292
R5489 VPWR.n2132 VPWR.n2130 0.120292
R5490 VPWR.n2135 VPWR.n2132 0.120292
R5491 VPWR.n2137 VPWR.n2135 0.120292
R5492 VPWR.n2139 VPWR.n2137 0.120292
R5493 VPWR.n2141 VPWR.n2139 0.120292
R5494 VPWR.n2146 VPWR.n2144 0.120292
R5495 VPWR.n2148 VPWR.n2146 0.120292
R5496 VPWR.n2150 VPWR.n2148 0.120292
R5497 VPWR.n2152 VPWR.n2150 0.120292
R5498 VPWR.n2153 VPWR.n2152 0.120292
R5499 VPWR.n2154 VPWR.n2153 0.120292
R5500 VPWR.n2159 VPWR.n2154 0.120292
R5501 VPWR.n2163 VPWR.n2162 0.120292
R5502 VPWR.n2164 VPWR.n2163 0.120292
R5503 VPWR.n2165 VPWR.n2164 0.120292
R5504 VPWR.n2170 VPWR.n2168 0.120292
R5505 VPWR.n2172 VPWR.n2170 0.120292
R5506 VPWR.n2174 VPWR.n2172 0.120292
R5507 VPWR.n2176 VPWR.n2174 0.120292
R5508 VPWR.n2178 VPWR.n2176 0.120292
R5509 VPWR.n2180 VPWR.n2178 0.120292
R5510 VPWR.n2182 VPWR.n2180 0.120292
R5511 VPWR.n2184 VPWR.n2182 0.120292
R5512 VPWR.n2186 VPWR.n2184 0.120292
R5513 VPWR.n2188 VPWR.n2186 0.120292
R5514 VPWR.n2190 VPWR.n2188 0.120292
R5515 VPWR.n2192 VPWR.n2190 0.120292
R5516 VPWR.n2194 VPWR.n2192 0.120292
R5517 VPWR.n2196 VPWR.n2194 0.120292
R5518 VPWR.n2198 VPWR.n2196 0.120292
R5519 VPWR.n2200 VPWR.n2198 0.120292
R5520 VPWR.n2202 VPWR.n2200 0.120292
R5521 VPWR.n2204 VPWR.n2202 0.120292
R5522 VPWR.n2205 VPWR.n2204 0.120292
R5523 VPWR.n2209 VPWR.n2208 0.120292
R5524 VPWR.n2210 VPWR.n2209 0.120292
R5525 VPWR.n2211 VPWR.n2210 0.120292
R5526 VPWR.n2306 VPWR.n2304 0.120292
R5527 VPWR.n2301 VPWR.n2300 0.120292
R5528 VPWR.n2300 VPWR.n2298 0.120292
R5529 VPWR.n2298 VPWR 0.120292
R5530 VPWR.n2295 VPWR.n2294 0.120292
R5531 VPWR.n2294 VPWR.n2293 0.120292
R5532 VPWR.n2293 VPWR.n2292 0.120292
R5533 VPWR.n2292 VPWR.n2290 0.120292
R5534 VPWR.n2290 VPWR.n2288 0.120292
R5535 VPWR.n2288 VPWR.n2286 0.120292
R5536 VPWR.n2286 VPWR.n2284 0.120292
R5537 VPWR.n2281 VPWR.n2280 0.120292
R5538 VPWR.n2280 VPWR.n2278 0.120292
R5539 VPWR.n2278 VPWR.n2277 0.120292
R5540 VPWR.n2277 VPWR.n2275 0.120292
R5541 VPWR.n2275 VPWR.n2273 0.120292
R5542 VPWR.n2273 VPWR.n2271 0.120292
R5543 VPWR.n2271 VPWR.n2269 0.120292
R5544 VPWR.n2269 VPWR.n2267 0.120292
R5545 VPWR.n7 VPWR.n5 0.120292
R5546 VPWR.n9 VPWR.n7 0.120292
R5547 VPWR VPWR.n9 0.120292
R5548 VPWR.n6303 VPWR.n6302 0.120292
R5549 VPWR.n6302 VPWR.n6301 0.120292
R5550 VPWR.n6301 VPWR 0.120292
R5551 VPWR.n6297 VPWR.n6296 0.120292
R5552 VPWR.n6296 VPWR.n6295 0.120292
R5553 VPWR.n6295 VPWR.n6294 0.120292
R5554 VPWR.n6294 VPWR.n6293 0.120292
R5555 VPWR.n6293 VPWR.n6292 0.120292
R5556 VPWR.n6257 VPWR.n39 0.120292
R5557 VPWR.n42 VPWR.n39 0.120292
R5558 VPWR VPWR.n42 0.120292
R5559 VPWR.n6250 VPWR.n6249 0.120292
R5560 VPWR.n6249 VPWR.n6248 0.120292
R5561 VPWR.n6248 VPWR.n6246 0.120292
R5562 VPWR.n6246 VPWR.n6244 0.120292
R5563 VPWR.n6240 VPWR.n6239 0.120292
R5564 VPWR.n6239 VPWR.n6238 0.120292
R5565 VPWR.n6238 VPWR.n6235 0.120292
R5566 VPWR.n6235 VPWR.n6233 0.120292
R5567 VPWR.n6233 VPWR.n6231 0.120292
R5568 VPWR.n6225 VPWR.n6223 0.120292
R5569 VPWR.n6223 VPWR.n6222 0.120292
R5570 VPWR.n6222 VPWR.n6221 0.120292
R5571 VPWR.n6218 VPWR.n6217 0.120292
R5572 VPWR.n6217 VPWR.n6215 0.120292
R5573 VPWR.n6211 VPWR.n6210 0.120292
R5574 VPWR.n6210 VPWR.n6208 0.120292
R5575 VPWR.n6208 VPWR.n6207 0.120292
R5576 VPWR.n6207 VPWR.n6206 0.120292
R5577 VPWR.n72 VPWR.n71 0.120292
R5578 VPWR.n6201 VPWR.n72 0.120292
R5579 VPWR.n6089 VPWR.n6087 0.120292
R5580 VPWR.n6091 VPWR.n6089 0.120292
R5581 VPWR.n6093 VPWR.n6091 0.120292
R5582 VPWR.n6101 VPWR.n6100 0.120292
R5583 VPWR.n6102 VPWR.n6101 0.120292
R5584 VPWR.n6103 VPWR.n6102 0.120292
R5585 VPWR.n6108 VPWR.n6106 0.120292
R5586 VPWR.n6110 VPWR.n6108 0.120292
R5587 VPWR.n6111 VPWR.n6110 0.120292
R5588 VPWR.n6116 VPWR.n6114 0.120292
R5589 VPWR.n6117 VPWR.n6116 0.120292
R5590 VPWR.n6124 VPWR.n6123 0.120292
R5591 VPWR.n6125 VPWR.n6124 0.120292
R5592 VPWR.n6127 VPWR.n6125 0.120292
R5593 VPWR.n6134 VPWR.n6133 0.120292
R5594 VPWR.n6135 VPWR.n6134 0.120292
R5595 VPWR.n6138 VPWR.n6135 0.120292
R5596 VPWR.n6140 VPWR.n6139 0.120292
R5597 VPWR.n6141 VPWR.n6140 0.120292
R5598 VPWR VPWR.n6141 0.120292
R5599 VPWR.n6148 VPWR.n6147 0.120292
R5600 VPWR.n6149 VPWR.n6148 0.120292
R5601 VPWR.n6155 VPWR.n6154 0.120292
R5602 VPWR.n6156 VPWR.n6155 0.120292
R5603 VPWR.n6160 VPWR.n6159 0.120292
R5604 VPWR.n6161 VPWR.n6160 0.120292
R5605 VPWR.n6166 VPWR.n6161 0.120292
R5606 VPWR.n6172 VPWR.n6170 0.120292
R5607 VPWR.n6174 VPWR.n6172 0.120292
R5608 VPWR.n6175 VPWR.n6174 0.120292
R5609 VPWR.n6176 VPWR.n6175 0.120292
R5610 VPWR.n6177 VPWR.n6176 0.120292
R5611 VPWR.n5638 VPWR.n5633 0.120292
R5612 VPWR.n5633 VPWR.n5632 0.120292
R5613 VPWR.n5632 VPWR.n5631 0.120292
R5614 VPWR.n5627 VPWR.n5626 0.120292
R5615 VPWR.n5626 VPWR.n5624 0.120292
R5616 VPWR.n5624 VPWR.n5623 0.120292
R5617 VPWR.n5623 VPWR.n5620 0.120292
R5618 VPWR.n5620 VPWR.n5618 0.120292
R5619 VPWR.n5618 VPWR.n5616 0.120292
R5620 VPWR.n5613 VPWR.n5612 0.120292
R5621 VPWR.n5612 VPWR.n5610 0.120292
R5622 VPWR.n5610 VPWR.n5608 0.120292
R5623 VPWR.n5608 VPWR.n5606 0.120292
R5624 VPWR.n5606 VPWR.n5604 0.120292
R5625 VPWR.n5604 VPWR.n5602 0.120292
R5626 VPWR.n5599 VPWR.n5598 0.120292
R5627 VPWR.n3629 VPWR.n3628 0.118519
R5628 VPWR.n3991 VPWR.n3988 0.118519
R5629 VPWR.n2944 VPWR.n2940 0.116385
R5630 VPWR.n4715 VPWR.n4712 0.116385
R5631 VPWR.n5163 VPWR.n5160 0.116385
R5632 VPWR.n460 VPWR.n459 0.116385
R5633 VPWR.n5461 VPWR.n5458 0.116385
R5634 VPWR.n2111 VPWR.n2110 0.116385
R5635 VPWR.n6087 VPWR.n6083 0.116385
R5636 VPWR.n5639 VPWR 0.113757
R5637 VPWR.n53 VPWR.n50 0.112576
R5638 VPWR.n5932 VPWR.n5929 0.108365
R5639 VPWR.n1564 VPWR.n1563 0.104667
R5640 VPWR.n1886 VPWR.n1885 0.104667
R5641 VPWR.n3196 VPWR.n3195 0.104667
R5642 VPWR.n1185 VPWR.n1184 0.104667
R5643 VPWR.n744 VPWR.n743 0.104667
R5644 VPWR.n4442 VPWR.n4441 0.104667
R5645 VPWR.n4989 VPWR.n4988 0.104667
R5646 VPWR.n1526 VPWR 0.104136
R5647 VPWR.n1846 VPWR 0.104136
R5648 VPWR.n3158 VPWR 0.104136
R5649 VPWR.n1143 VPWR 0.104136
R5650 VPWR.n3814 VPWR 0.104136
R5651 VPWR.n705 VPWR 0.104136
R5652 VPWR.n4403 VPWR 0.104136
R5653 VPWR.n4948 VPWR 0.104136
R5654 VPWR.n195 VPWR 0.104136
R5655 VPWR.n5867 VPWR 0.104136
R5656 VPWR.n1 VPWR 0.104136
R5657 VPWR.n2263 VPWR 0.102383
R5658 VPWR.n1879 VPWR 0.0994583
R5659 VPWR VPWR.n1487 0.0994583
R5660 VPWR.n3399 VPWR 0.0994583
R5661 VPWR.n1175 VPWR 0.0994583
R5662 VPWR VPWR.n3721 0.0994583
R5663 VPWR.n3707 VPWR 0.0994583
R5664 VPWR VPWR.n3706 0.0994583
R5665 VPWR.n3675 VPWR 0.0994583
R5666 VPWR.n1272 VPWR 0.0994583
R5667 VPWR VPWR.n3569 0.0994583
R5668 VPWR.n3501 VPWR 0.0994583
R5669 VPWR VPWR 0.0994583
R5670 VPWR.n3940 VPWR 0.0994583
R5671 VPWR.n4063 VPWR 0.0994583
R5672 VPWR VPWR.n815 0.0994583
R5673 VPWR.n919 VPWR 0.0994583
R5674 VPWR.n940 VPWR 0.0994583
R5675 VPWR.n4695 VPWR 0.0994583
R5676 VPWR.n4770 VPWR 0.0994583
R5677 VPWR.n5059 VPWR 0.0994583
R5678 VPWR.n5177 VPWR 0.0994583
R5679 VPWR.n5209 VPWR 0.0994583
R5680 VPWR.n5246 VPWR 0.0994583
R5681 VPWR.n580 VPWR 0.0994583
R5682 VPWR.n608 VPWR 0.0994583
R5683 VPWR.n6049 VPWR 0.0994583
R5684 VPWR.n5481 VPWR 0.0994583
R5685 VPWR.n1530 VPWR 0.0981562
R5686 VPWR VPWR 0.0981562
R5687 VPWR.n1536 VPWR 0.0981562
R5688 VPWR VPWR.n1538 0.0981562
R5689 VPWR.n1545 VPWR 0.0981562
R5690 VPWR.n1546 VPWR 0.0981562
R5691 VPWR.n2842 VPWR 0.0981562
R5692 VPWR.n2848 VPWR 0.0981562
R5693 VPWR VPWR.n2774 0.0981562
R5694 VPWR.n2851 VPWR 0.0981562
R5695 VPWR.n2859 VPWR 0.0981562
R5696 VPWR.n2867 VPWR 0.0981562
R5697 VPWR.n2893 VPWR 0.0981562
R5698 VPWR VPWR.n2736 0.0981562
R5699 VPWR.n2732 VPWR 0.0981562
R5700 VPWR.n2726 VPWR 0.0981562
R5701 VPWR VPWR.n2725 0.0981562
R5702 VPWR.n2714 VPWR 0.0981562
R5703 VPWR.n2695 VPWR 0.0981562
R5704 VPWR VPWR.n2690 0.0981562
R5705 VPWR.n2682 VPWR 0.0981562
R5706 VPWR VPWR.n2681 0.0981562
R5707 VPWR.n2669 VPWR 0.0981562
R5708 VPWR VPWR 0.0981562
R5709 VPWR.n2663 VPWR 0.0981562
R5710 VPWR.n1661 VPWR.n1660 0.0981562
R5711 VPWR.n1655 VPWR 0.0981562
R5712 VPWR VPWR.n1643 0.0981562
R5713 VPWR VPWR.n1637 0.0981562
R5714 VPWR VPWR.n1636 0.0981562
R5715 VPWR VPWR.n1631 0.0981562
R5716 VPWR.n1628 VPWR 0.0981562
R5717 VPWR VPWR.n1626 0.0981562
R5718 VPWR.n1850 VPWR 0.0981562
R5719 VPWR VPWR 0.0981562
R5720 VPWR.n1857 VPWR 0.0981562
R5721 VPWR VPWR.n1840 0.0981562
R5722 VPWR.n1869 VPWR 0.0981562
R5723 VPWR VPWR.n1821 0.0981562
R5724 VPWR.n1947 VPWR 0.0981562
R5725 VPWR.n1950 VPWR 0.0981562
R5726 VPWR.n1954 VPWR 0.0981562
R5727 VPWR.n1969 VPWR 0.0981562
R5728 VPWR.n1970 VPWR 0.0981562
R5729 VPWR.n2024 VPWR 0.0981562
R5730 VPWR.n2017 VPWR 0.0981562
R5731 VPWR.n1979 VPWR 0.0981562
R5732 VPWR VPWR 0.0981562
R5733 VPWR.n2950 VPWR 0.0981562
R5734 VPWR VPWR 0.0981562
R5735 VPWR.n2957 VPWR 0.0981562
R5736 VPWR.n2965 VPWR 0.0981562
R5737 VPWR.n2969 VPWR 0.0981562
R5738 VPWR.n2972 VPWR 0.0981562
R5739 VPWR.n3027 VPWR 0.0981562
R5740 VPWR.n3020 VPWR 0.0981562
R5741 VPWR.n3014 VPWR 0.0981562
R5742 VPWR.n3009 VPWR 0.0981562
R5743 VPWR.n2996 VPWR 0.0981562
R5744 VPWR.n1745 VPWR.n1744 0.0981562
R5745 VPWR.n1739 VPWR 0.0981562
R5746 VPWR.n1726 VPWR 0.0981562
R5747 VPWR VPWR.n1725 0.0981562
R5748 VPWR.n1713 VPWR 0.0981562
R5749 VPWR.n1697 VPWR 0.0981562
R5750 VPWR VPWR.n1708 0.0981562
R5751 VPWR VPWR.n3155 0.0981562
R5752 VPWR.n3165 VPWR 0.0981562
R5753 VPWR VPWR.n3166 0.0981562
R5754 VPWR.n3175 VPWR 0.0981562
R5755 VPWR.n3176 VPWR 0.0981562
R5756 VPWR.n3266 VPWR 0.0981562
R5757 VPWR VPWR.n3265 0.0981562
R5758 VPWR.n3259 VPWR 0.0981562
R5759 VPWR.n3243 VPWR 0.0981562
R5760 VPWR.n3298 VPWR 0.0981562
R5761 VPWR.n3306 VPWR 0.0981562
R5762 VPWR.n3310 VPWR 0.0981562
R5763 VPWR.n3327 VPWR 0.0981562
R5764 VPWR VPWR 0.0981562
R5765 VPWR.n3331 VPWR 0.0981562
R5766 VPWR.n3362 VPWR 0.0981562
R5767 VPWR.n3370 VPWR 0.0981562
R5768 VPWR VPWR 0.0981562
R5769 VPWR.n3383 VPWR 0.0981562
R5770 VPWR.n3389 VPWR 0.0981562
R5771 VPWR.n3390 VPWR 0.0981562
R5772 VPWR.n3436 VPWR 0.0981562
R5773 VPWR VPWR.n3433 0.0981562
R5774 VPWR.n3426 VPWR 0.0981562
R5775 VPWR VPWR.n3423 0.0981562
R5776 VPWR VPWR.n3416 0.0981562
R5777 VPWR VPWR.n3415 0.0981562
R5778 VPWR.n3407 VPWR 0.0981562
R5779 VPWR.n1376 VPWR.n1375 0.0981562
R5780 VPWR.n1370 VPWR 0.0981562
R5781 VPWR VPWR.n1369 0.0981562
R5782 VPWR.n1357 VPWR 0.0981562
R5783 VPWR.n1351 VPWR 0.0981562
R5784 VPWR VPWR 0.0981562
R5785 VPWR VPWR.n1345 0.0981562
R5786 VPWR.n1341 VPWR 0.0981562
R5787 VPWR.n1153 VPWR 0.0981562
R5788 VPWR.n1156 VPWR 0.0981562
R5789 VPWR.n1165 VPWR 0.0981562
R5790 VPWR.n3733 VPWR 0.0981562
R5791 VPWR VPWR.n3732 0.0981562
R5792 VPWR.n3727 VPWR 0.0981562
R5793 VPWR.n3722 VPWR 0.0981562
R5794 VPWR.n3715 VPWR 0.0981562
R5795 VPWR.n3700 VPWR 0.0981562
R5796 VPWR.n3692 VPWR 0.0981562
R5797 VPWR.n3669 VPWR 0.0981562
R5798 VPWR VPWR.n3668 0.0981562
R5799 VPWR.n3664 VPWR 0.0981562
R5800 VPWR VPWR.n3627 0.0981562
R5801 VPWR VPWR.n3621 0.0981562
R5802 VPWR.n3604 VPWR 0.0981562
R5803 VPWR.n3593 VPWR 0.0981562
R5804 VPWR.n3587 VPWR 0.0981562
R5805 VPWR.n3570 VPWR 0.0981562
R5806 VPWR.n3563 VPWR 0.0981562
R5807 VPWR.n3526 VPWR.n3525 0.0981562
R5808 VPWR.n3516 VPWR 0.0981562
R5809 VPWR VPWR 0.0981562
R5810 VPWR VPWR.n3495 0.0981562
R5811 VPWR.n3486 VPWR 0.0981562
R5812 VPWR.n3818 VPWR 0.0981562
R5813 VPWR VPWR.n3812 0.0981562
R5814 VPWR VPWR.n3811 0.0981562
R5815 VPWR.n3825 VPWR 0.0981562
R5816 VPWR.n3894 VPWR 0.0981562
R5817 VPWR.n3902 VPWR 0.0981562
R5818 VPWR.n3907 VPWR 0.0981562
R5819 VPWR.n3909 VPWR 0.0981562
R5820 VPWR VPWR.n1127 0.0981562
R5821 VPWR.n3915 VPWR 0.0981562
R5822 VPWR.n3919 VPWR 0.0981562
R5823 VPWR.n3959 VPWR 0.0981562
R5824 VPWR.n3953 VPWR 0.0981562
R5825 VPWR.n3947 VPWR 0.0981562
R5826 VPWR VPWR.n3946 0.0981562
R5827 VPWR VPWR.n3939 0.0981562
R5828 VPWR.n3932 VPWR 0.0981562
R5829 VPWR.n4001 VPWR 0.0981562
R5830 VPWR.n4013 VPWR 0.0981562
R5831 VPWR.n4016 VPWR 0.0981562
R5832 VPWR.n4030 VPWR 0.0981562
R5833 VPWR VPWR.n4077 0.0981562
R5834 VPWR VPWR.n4076 0.0981562
R5835 VPWR VPWR.n4062 0.0981562
R5836 VPWR.n4057 VPWR 0.0981562
R5837 VPWR.n4047 VPWR 0.0981562
R5838 VPWR.n1040 VPWR.n1039 0.0981562
R5839 VPWR.n1034 VPWR 0.0981562
R5840 VPWR.n1027 VPWR 0.0981562
R5841 VPWR.n1021 VPWR 0.0981562
R5842 VPWR.n1014 VPWR 0.0981562
R5843 VPWR.n1008 VPWR 0.0981562
R5844 VPWR VPWR 0.0981562
R5845 VPWR.n711 VPWR 0.0981562
R5846 VPWR.n720 VPWR 0.0981562
R5847 VPWR.n725 VPWR 0.0981562
R5848 VPWR.n737 VPWR 0.0981562
R5849 VPWR VPWR.n826 0.0981562
R5850 VPWR.n869 VPWR 0.0981562
R5851 VPWR.n870 VPWR 0.0981562
R5852 VPWR.n883 VPWR 0.0981562
R5853 VPWR.n884 VPWR 0.0981562
R5854 VPWR.n886 VPWR 0.0981562
R5855 VPWR.n889 VPWR 0.0981562
R5856 VPWR.n898 VPWR 0.0981562
R5857 VPWR.n906 VPWR 0.0981562
R5858 VPWR.n923 VPWR 0.0981562
R5859 VPWR.n931 VPWR 0.0981562
R5860 VPWR.n4247 VPWR 0.0981562
R5861 VPWR VPWR 0.0981562
R5862 VPWR.n4252 VPWR 0.0981562
R5863 VPWR.n4268 VPWR 0.0981562
R5864 VPWR.n4277 VPWR 0.0981562
R5865 VPWR.n4282 VPWR 0.0981562
R5866 VPWR.n4290 VPWR 0.0981562
R5867 VPWR.n4311 VPWR 0.0981562
R5868 VPWR.n4323 VPWR 0.0981562
R5869 VPWR.n4326 VPWR 0.0981562
R5870 VPWR.n4335 VPWR 0.0981562
R5871 VPWR.n4336 VPWR 0.0981562
R5872 VPWR.n4200 VPWR.n4199 0.0981562
R5873 VPWR.n4194 VPWR 0.0981562
R5874 VPWR VPWR.n4193 0.0981562
R5875 VPWR VPWR.n4192 0.0981562
R5876 VPWR.n4181 VPWR 0.0981562
R5877 VPWR VPWR.n4180 0.0981562
R5878 VPWR VPWR 0.0981562
R5879 VPWR VPWR.n4167 0.0981562
R5880 VPWR VPWR 0.0981562
R5881 VPWR.n4409 VPWR 0.0981562
R5882 VPWR.n4418 VPWR 0.0981562
R5883 VPWR.n4423 VPWR 0.0981562
R5884 VPWR.n4435 VPWR 0.0981562
R5885 VPWR.n4872 VPWR 0.0981562
R5886 VPWR VPWR.n4870 0.0981562
R5887 VPWR.n4860 VPWR 0.0981562
R5888 VPWR VPWR.n4859 0.0981562
R5889 VPWR.n4848 VPWR 0.0981562
R5890 VPWR.n4837 VPWR 0.0981562
R5891 VPWR VPWR.n4836 0.0981562
R5892 VPWR VPWR.n4833 0.0981562
R5893 VPWR.n4662 VPWR 0.0981562
R5894 VPWR.n4667 VPWR 0.0981562
R5895 VPWR.n4690 VPWR 0.0981562
R5896 VPWR.n4694 VPWR 0.0981562
R5897 VPWR.n4716 VPWR 0.0981562
R5898 VPWR.n4717 VPWR 0.0981562
R5899 VPWR.n4737 VPWR 0.0981562
R5900 VPWR.n4746 VPWR 0.0981562
R5901 VPWR.n4752 VPWR 0.0981562
R5902 VPWR.n4766 VPWR 0.0981562
R5903 VPWR VPWR.n4585 0.0981562
R5904 VPWR.n4783 VPWR 0.0981562
R5905 VPWR.n4789 VPWR 0.0981562
R5906 VPWR.n4794 VPWR 0.0981562
R5907 VPWR.n4800 VPWR 0.0981562
R5908 VPWR.n4563 VPWR.n4562 0.0981562
R5909 VPWR.n4559 VPWR 0.0981562
R5910 VPWR VPWR.n4558 0.0981562
R5911 VPWR VPWR.n4553 0.0981562
R5912 VPWR.n4543 VPWR 0.0981562
R5913 VPWR VPWR 0.0981562
R5914 VPWR VPWR.n4525 0.0981562
R5915 VPWR VPWR.n4946 0.0981562
R5916 VPWR VPWR 0.0981562
R5917 VPWR.n4958 VPWR 0.0981562
R5918 VPWR.n4964 VPWR 0.0981562
R5919 VPWR VPWR.n4940 0.0981562
R5920 VPWR.n4970 VPWR 0.0981562
R5921 VPWR.n4976 VPWR 0.0981562
R5922 VPWR.n4982 VPWR 0.0981562
R5923 VPWR VPWR.n682 0.0981562
R5924 VPWR.n5062 VPWR 0.0981562
R5925 VPWR.n5073 VPWR 0.0981562
R5926 VPWR.n5089 VPWR 0.0981562
R5927 VPWR.n5142 VPWR 0.0981562
R5928 VPWR VPWR.n5139 0.0981562
R5929 VPWR VPWR.n5132 0.0981562
R5930 VPWR.n5104 VPWR 0.0981562
R5931 VPWR VPWR.n5127 0.0981562
R5932 VPWR VPWR.n5126 0.0981562
R5933 VPWR.n5120 VPWR 0.0981562
R5934 VPWR VPWR.n5119 0.0981562
R5935 VPWR.n5115 VPWR 0.0981562
R5936 VPWR.n5167 VPWR 0.0981562
R5937 VPWR.n5172 VPWR 0.0981562
R5938 VPWR.n5179 VPWR 0.0981562
R5939 VPWR.n5184 VPWR 0.0981562
R5940 VPWR.n5190 VPWR 0.0981562
R5941 VPWR.n5213 VPWR 0.0981562
R5942 VPWR VPWR.n5258 0.0981562
R5943 VPWR.n5225 VPWR 0.0981562
R5944 VPWR VPWR.n5232 0.0981562
R5945 VPWR VPWR.n5231 0.0981562
R5946 VPWR.n293 VPWR.n292 0.0981562
R5947 VPWR.n283 VPWR 0.0981562
R5948 VPWR VPWR 0.0981562
R5949 VPWR VPWR.n273 0.0981562
R5950 VPWR.n197 VPWR 0.0981562
R5951 VPWR.n200 VPWR 0.0981562
R5952 VPWR.n204 VPWR 0.0981562
R5953 VPWR VPWR.n189 0.0981562
R5954 VPWR.n208 VPWR 0.0981562
R5955 VPWR.n534 VPWR 0.0981562
R5956 VPWR.n537 VPWR 0.0981562
R5957 VPWR.n541 VPWR 0.0981562
R5958 VPWR.n543 VPWR 0.0981562
R5959 VPWR.n547 VPWR 0.0981562
R5960 VPWR.n553 VPWR 0.0981562
R5961 VPWR.n558 VPWR 0.0981562
R5962 VPWR.n561 VPWR 0.0981562
R5963 VPWR VPWR.n497 0.0981562
R5964 VPWR.n571 VPWR 0.0981562
R5965 VPWR.n574 VPWR 0.0981562
R5966 VPWR.n586 VPWR 0.0981562
R5967 VPWR.n587 VPWR 0.0981562
R5968 VPWR.n588 VPWR 0.0981562
R5969 VPWR.n591 VPWR 0.0981562
R5970 VPWR.n599 VPWR 0.0981562
R5971 VPWR.n604 VPWR 0.0981562
R5972 VPWR.n450 VPWR 0.0981562
R5973 VPWR.n435 VPWR 0.0981562
R5974 VPWR.n429 VPWR 0.0981562
R5975 VPWR VPWR.n428 0.0981562
R5976 VPWR.n423 VPWR 0.0981562
R5977 VPWR VPWR.n422 0.0981562
R5978 VPWR VPWR.n412 0.0981562
R5979 VPWR VPWR.n404 0.0981562
R5980 VPWR.n398 VPWR 0.0981562
R5981 VPWR VPWR.n392 0.0981562
R5982 VPWR.n387 VPWR 0.0981562
R5983 VPWR VPWR.n385 0.0981562
R5984 VPWR.n382 VPWR 0.0981562
R5985 VPWR.n378 VPWR 0.0981562
R5986 VPWR VPWR.n377 0.0981562
R5987 VPWR.n5374 VPWR.n5373 0.0981562
R5988 VPWR.n5368 VPWR 0.0981562
R5989 VPWR.n5362 VPWR 0.0981562
R5990 VPWR.n5351 VPWR 0.0981562
R5991 VPWR VPWR.n5347 0.0981562
R5992 VPWR.n5342 VPWR 0.0981562
R5993 VPWR VPWR.n5862 0.0981562
R5994 VPWR.n5876 VPWR 0.0981562
R5995 VPWR.n5879 VPWR 0.0981562
R5996 VPWR.n5881 VPWR 0.0981562
R5997 VPWR.n5882 VPWR 0.0981562
R5998 VPWR.n5983 VPWR 0.0981562
R5999 VPWR.n5987 VPWR 0.0981562
R6000 VPWR.n6001 VPWR 0.0981562
R6001 VPWR.n6013 VPWR 0.0981562
R6002 VPWR.n6019 VPWR 0.0981562
R6003 VPWR.n6035 VPWR 0.0981562
R6004 VPWR.n6052 VPWR 0.0981562
R6005 VPWR.n5465 VPWR 0.0981562
R6006 VPWR.n5488 VPWR 0.0981562
R6007 VPWR.n5491 VPWR 0.0981562
R6008 VPWR VPWR.n5405 0.0981562
R6009 VPWR.n5516 VPWR 0.0981562
R6010 VPWR.n5527 VPWR 0.0981562
R6011 VPWR.n5533 VPWR 0.0981562
R6012 VPWR.n5539 VPWR 0.0981562
R6013 VPWR.n5547 VPWR 0.0981562
R6014 VPWR.n5740 VPWR.n5738 0.0981562
R6015 VPWR.n5726 VPWR 0.0981562
R6016 VPWR.n5718 VPWR 0.0981562
R6017 VPWR VPWR 0.0981562
R6018 VPWR VPWR.n5701 0.0981562
R6019 VPWR.n2412 VPWR 0.0981562
R6020 VPWR.n2418 VPWR 0.0981562
R6021 VPWR.n2424 VPWR 0.0981562
R6022 VPWR.n2430 VPWR 0.0981562
R6023 VPWR.n2438 VPWR 0.0981562
R6024 VPWR.n2484 VPWR 0.0981562
R6025 VPWR.n2496 VPWR 0.0981562
R6026 VPWR VPWR 0.0981562
R6027 VPWR.n2522 VPWR 0.0981562
R6028 VPWR.n2535 VPWR 0.0981562
R6029 VPWR.n2545 VPWR 0.0981562
R6030 VPWR.n2548 VPWR 0.0981562
R6031 VPWR.n2556 VPWR 0.0981562
R6032 VPWR.n2559 VPWR 0.0981562
R6033 VPWR.n2592 VPWR 0.0981562
R6034 VPWR.n2114 VPWR 0.0981562
R6035 VPWR.n2123 VPWR 0.0981562
R6036 VPWR VPWR.n2076 0.0981562
R6037 VPWR.n2130 VPWR 0.0981562
R6038 VPWR.n2142 VPWR 0.0981562
R6039 VPWR.n2144 VPWR 0.0981562
R6040 VPWR.n2160 VPWR 0.0981562
R6041 VPWR.n2168 VPWR 0.0981562
R6042 VPWR.n2208 VPWR 0.0981562
R6043 VPWR.n2307 VPWR.n2306 0.0981562
R6044 VPWR.n2301 VPWR 0.0981562
R6045 VPWR.n2295 VPWR 0.0981562
R6046 VPWR VPWR 0.0981562
R6047 VPWR VPWR.n2281 0.0981562
R6048 VPWR.n2264 VPWR 0.0981562
R6049 VPWR.n5 VPWR 0.0981562
R6050 VPWR.n6303 VPWR 0.0981562
R6051 VPWR.n6297 VPWR 0.0981562
R6052 VPWR.n6289 VPWR 0.0981562
R6053 VPWR VPWR.n6257 0.0981562
R6054 VPWR VPWR.n6252 0.0981562
R6055 VPWR VPWR 0.0981562
R6056 VPWR VPWR.n6241 0.0981562
R6057 VPWR VPWR.n6240 0.0981562
R6058 VPWR.n6228 VPWR 0.0981562
R6059 VPWR VPWR 0.0981562
R6060 VPWR VPWR.n6218 0.0981562
R6061 VPWR.n6211 VPWR 0.0981562
R6062 VPWR.n71 VPWR 0.0981562
R6063 VPWR VPWR.n6199 0.0981562
R6064 VPWR VPWR 0.0981562
R6065 VPWR.n6100 VPWR 0.0981562
R6066 VPWR VPWR.n90 0.0981562
R6067 VPWR.n6114 VPWR 0.0981562
R6068 VPWR.n6123 VPWR 0.0981562
R6069 VPWR.n6128 VPWR 0.0981562
R6070 VPWR.n6139 VPWR 0.0981562
R6071 VPWR.n6146 VPWR 0.0981562
R6072 VPWR.n6147 VPWR 0.0981562
R6073 VPWR VPWR 0.0981562
R6074 VPWR.n6154 VPWR 0.0981562
R6075 VPWR.n6159 VPWR 0.0981562
R6076 VPWR VPWR 0.0981562
R6077 VPWR.n6167 VPWR 0.0981562
R6078 VPWR VPWR.n5638 0.0981562
R6079 VPWR VPWR 0.0981562
R6080 VPWR.n5627 VPWR 0.0981562
R6081 VPWR VPWR 0.0981562
R6082 VPWR VPWR.n5613 0.0981562
R6083 VPWR.n5599 VPWR 0.0981562
R6084 VPWR VPWR.n1654 0.0968542
R6085 VPWR.n1941 VPWR 0.0968542
R6086 VPWR VPWR.n1738 0.0968542
R6087 VPWR.n3179 VPWR 0.0968542
R6088 VPWR VPWR.n3258 0.0968542
R6089 VPWR.n3624 VPWR 0.0968542
R6090 VPWR VPWR.n4068 0.0968542
R6091 VPWR VPWR.n1007 0.0968542
R6092 VPWR.n4255 VPWR 0.0968542
R6093 VPWR.n4280 VPWR 0.0968542
R6094 VPWR VPWR.n4191 0.0968542
R6095 VPWR VPWR.n4871 0.0968542
R6096 VPWR.n4683 VPWR 0.0968542
R6097 VPWR.n4720 VPWR 0.0968542
R6098 VPWR VPWR.n4542 0.0968542
R6099 VPWR.n5255 VPWR 0.0968542
R6100 VPWR VPWR.n5350 0.0968542
R6101 VPWR VPWR.n5341 0.0968542
R6102 VPWR.n5990 VPWR 0.0968542
R6103 VPWR VPWR.n5725 0.0968542
R6104 VPWR.n4210 VPWR.n4207 0.0942472
R6105 VPWR.n4223 VPWR.n4213 0.0942472
R6106 VPWR.n3410 VPWR 0.0913841
R6107 VPWR.n1537 VPWR 0.0890417
R6108 VPWR.n2861 VPWR 0.0890417
R6109 VPWR VPWR.n2689 0.0890417
R6110 VPWR VPWR.n2668 0.0890417
R6111 VPWR VPWR.n1819 0.0890417
R6112 VPWR VPWR.n2023 0.0890417
R6113 VPWR VPWR.n3026 0.0890417
R6114 VPWR VPWR.n3008 0.0890417
R6115 VPWR.n3167 VPWR 0.0890417
R6116 VPWR.n3189 VPWR 0.0890417
R6117 VPWR.n3299 VPWR 0.0890417
R6118 VPWR.n3371 VPWR 0.0890417
R6119 VPWR.n3402 VPWR 0.0890417
R6120 VPWR.n1150 VPWR 0.0890417
R6121 VPWR VPWR.n3699 0.0890417
R6122 VPWR VPWR.n3663 0.0890417
R6123 VPWR.n3655 VPWR 0.0890417
R6124 VPWR VPWR.n3586 0.0890417
R6125 VPWR.n3910 VPWR 0.0890417
R6126 VPWR.n3969 VPWR 0.0890417
R6127 VPWR VPWR.n3945 0.0890417
R6128 VPWR.n4080 VPWR 0.0890417
R6129 VPWR VPWR.n4046 0.0890417
R6130 VPWR VPWR.n703 0.0890417
R6131 VPWR.n871 VPWR 0.0890417
R6132 VPWR VPWR.n824 0.0890417
R6133 VPWR.n900 VPWR 0.0890417
R6134 VPWR.n920 VPWR 0.0890417
R6135 VPWR.n4292 VPWR 0.0890417
R6136 VPWR.n4405 VPWR 0.0890417
R6137 VPWR.n4731 VPWR 0.0890417
R6138 VPWR.n4768 VPWR 0.0890417
R6139 VPWR.n4963 VPWR 0.0890417
R6140 VPWR.n4977 VPWR 0.0890417
R6141 VPWR VPWR.n5141 0.0890417
R6142 VPWR.n5178 VPWR 0.0890417
R6143 VPWR.n5266 VPWR 0.0890417
R6144 VPWR VPWR.n5265 0.0890417
R6145 VPWR VPWR.n5241 0.0890417
R6146 VPWR.n572 VPWR 0.0890417
R6147 VPWR VPWR.n411 0.0890417
R6148 VPWR VPWR.n391 0.0890417
R6149 VPWR VPWR.n5361 0.0890417
R6150 VPWR.n5886 VPWR 0.0890417
R6151 VPWR.n6007 VPWR 0.0890417
R6152 VPWR.n6022 VPWR 0.0890417
R6153 VPWR.n5510 VPWR 0.0890417
R6154 VPWR VPWR.n5717 0.0890417
R6155 VPWR.n2541 VPWR 0.0890417
R6156 VPWR.n2162 VPWR 0.0890417
R6157 VPWR VPWR.n6227 0.0890417
R6158 VPWR.n6133 VPWR 0.0890417
R6159 VPWR.n6170 VPWR 0.0890417
R6160 VPWR.n1549 VPWR 0.0877396
R6161 VPWR.n2897 VPWR 0.0877396
R6162 VPWR.n1987 VPWR 0.0877396
R6163 VPWR.n3831 VPWR 0.0877396
R6164 VPWR.n4238 VPWR 0.0877396
R6165 VPWR.n4296 VPWR 0.0877396
R6166 VPWR VPWR.n4586 0.0877396
R6167 VPWR.n5049 VPWR 0.0877396
R6168 VPWR.n5135 VPWR 0.0877396
R6169 VPWR.n5242 VPWR 0.0877396
R6170 VPWR.n575 VPWR 0.0877396
R6171 VPWR.n2575 VPWR 0.0877396
R6172 VPWR VPWR.n6288 0.0869256
R6173 VPWR.n4070 VPWR 0.0835716
R6174 VPWR VPWR.n2841 0.0828946
R6175 VPWR VPWR.n2858 0.0828946
R6176 VPWR.n3895 VPWR 0.0828946
R6177 VPWR VPWR.n6094 0.0828946
R6178 VPWR VPWR.n2840 0.0826382
R6179 VPWR VPWR.n2847 0.0826382
R6180 VPWR.n2854 VPWR 0.0826382
R6181 VPWR VPWR.n1968 0.0826382
R6182 VPWR.n1978 VPWR 0.0826382
R6183 VPWR.n3002 VPWR 0.0826382
R6184 VPWR VPWR.n3379 0.0826382
R6185 VPWR VPWR.n3380 0.0826382
R6186 VPWR.n3406 VPWR 0.0826382
R6187 VPWR VPWR.n3305 0.0826382
R6188 VPWR VPWR.n3326 0.0826382
R6189 VPWR.n3556 VPWR 0.0826382
R6190 VPWR.n3555 VPWR 0.0826382
R6191 VPWR VPWR.n3900 0.0826382
R6192 VPWR.n3933 VPWR 0.0826382
R6193 VPWR.n3823 VPWR 0.0826382
R6194 VPWR.n5113 VPWR 0.0826382
R6195 VPWR VPWR.n570 0.0826382
R6196 VPWR.n206 VPWR 0.0826382
R6197 VPWR VPWR.n220 0.0826382
R6198 VPWR.n5348 VPWR 0.0826382
R6199 VPWR VPWR.n5973 0.0826382
R6200 VPWR VPWR.n2853 0.0822696
R6201 VPWR.n1625 VPWR 0.0822696
R6202 VPWR.n3156 VPWR 0.0822696
R6203 VPWR.n3725 VPWR 0.0822696
R6204 VPWR VPWR.n3901 0.0822696
R6205 VPWR.n1492 VPWR 0.0815925
R6206 VPWR.n1964 VPWR 0.0813361
R6207 VPWR.n5114 VPWR 0.0813361
R6208 VPWR.n2441 VPWR 0.0734167
R6209 VPWR.n2815 VPWR.n2808 0.0721146
R6210 VPWR.n1934 VPWR.n1930 0.0721146
R6211 VPWR.n3276 VPWR.n3275 0.0721146
R6212 VPWR.n3743 VPWR.n3742 0.0721146
R6213 VPWR.n3887 VPWR.n3884 0.0721146
R6214 VPWR.n862 VPWR.n858 0.0721146
R6215 VPWR.n4879 VPWR.n4878 0.0721146
R6216 VPWR.n5043 VPWR.n5042 0.0721146
R6217 VPWR.n5965 VPWR.n5959 0.0721146
R6218 VPWR.n2481 VPWR.n2480 0.0721146
R6219 VPWR.n6259 VPWR.n6258 0.0721146
R6220 VPWR.n2401 VPWR 0.0657573
R6221 VPWR.n1494 VPWR 0.0605028
R6222 VPWR VPWR.n1577 0.0590938
R6223 VPWR VPWR.n1753 0.0590938
R6224 VPWR VPWR.n1319 0.0590938
R6225 VPWR VPWR.n3554 0.0590938
R6226 VPWR VPWR.n1052 0.0590938
R6227 VPWR.n4806 VPWR 0.0590938
R6228 VPWR VPWR.n300 0.0590938
R6229 VPWR VPWR.n229 0.0590938
R6230 VPWR VPWR.n5381 0.0590938
R6231 VPWR.n2212 VPWR 0.0590938
R6232 VPWR.n6178 VPWR 0.0590938
R6233 VPWR.n5901 VPWR.n5900 0.0572053
R6234 VPWR.n1860 VPWR.n1859 0.0549681
R6235 VPWR.n3130 VPWR.n1511 0.0545016
R6236 VPWR.n4387 VPWR.n690 0.0545016
R6237 VPWR.n4339 VPWR 0.0499792
R6238 VPWR.n1602 VPWR.n1601 0.0460729
R6239 VPWR.n1684 VPWR.n1683 0.0460729
R6240 VPWR.n1324 VPWR.n1323 0.0460729
R6241 VPWR.n3469 VPWR.n3468 0.0460729
R6242 VPWR.n985 VPWR.n984 0.0460729
R6243 VPWR.n4139 VPWR.n4138 0.0460729
R6244 VPWR.n4507 VPWR.n4506 0.0460729
R6245 VPWR.n253 VPWR.n252 0.0460729
R6246 VPWR.n5316 VPWR.n5315 0.0460729
R6247 VPWR.n5685 VPWR.n5684 0.0460729
R6248 VPWR.n2243 VPWR.n2242 0.0460729
R6249 VPWR.n5588 VPWR.n5587 0.0460729
R6250 VPWR.n1247 VPWR.n1246 0.0444602
R6251 VPWR.n1071 VPWR.n1070 0.0444602
R6252 VPWR.n773 VPWR.n772 0.0444602
R6253 VPWR.n3110 VPWR.n3109 0.0434688
R6254 VPWR.n1891 VPWR.n1835 0.0434688
R6255 VPWR.n3212 VPWR.n3211 0.0434688
R6256 VPWR.n3773 VPWR.n3772 0.0434688
R6257 VPWR.n3872 VPWR.n3871 0.0434688
R6258 VPWR.n4377 VPWR.n4376 0.0434688
R6259 VPWR.n4908 VPWR.n4907 0.0434688
R6260 VPWR.n5030 VPWR.n5029 0.0434688
R6261 VPWR.n5806 VPWR.n5805 0.0434688
R6262 VPWR.n5947 VPWR.n5946 0.0434688
R6263 VPWR.n2458 VPWR.n2457 0.0434688
R6264 VPWR.n31 VPWR.n30 0.0434688
R6265 VPWR.n2031 VPWR.n2030 0.039085
R6266 VPWR.n3342 VPWR.n3341 0.0390849
R6267 VPWR.n144 VPWR.n143 0.0390849
R6268 VPWR.n1264 VPWR.n1263 0.0387485
R6269 VPWR.n3976 VPWR.n3975 0.0387485
R6270 VPWR.n950 VPWR.n949 0.0387485
R6271 VPWR.n5148 VPWR.n5147 0.0387485
R6272 VPWR.n618 VPWR.n617 0.0387485
R6273 VPWR.n1546 VPWR 0.0330521
R6274 VPWR.n2894 VPWR 0.0330521
R6275 VPWR.n1990 VPWR 0.0330521
R6276 VPWR.n3003 VPWR 0.0330521
R6277 VPWR.n3828 VPWR 0.0330521
R6278 VPWR.n703 VPWR 0.0330521
R6279 VPWR.n4293 VPWR 0.0330521
R6280 VPWR.n4405 VPWR 0.0330521
R6281 VPWR VPWR.n4685 0.0330521
R6282 VPWR.n4769 VPWR 0.0330521
R6283 VPWR.n5245 VPWR 0.0330521
R6284 VPWR VPWR.n574 0.0330521
R6285 VPWR.n2572 VPWR 0.0330521
R6286 VPWR VPWR.n1536 0.03175
R6287 VPWR VPWR.n2859 0.03175
R6288 VPWR.n2690 VPWR 0.03175
R6289 VPWR.n2669 VPWR 0.03175
R6290 VPWR.n1944 VPWR 0.03175
R6291 VPWR VPWR.n1947 0.03175
R6292 VPWR.n2024 VPWR 0.03175
R6293 VPWR.n1979 VPWR 0.03175
R6294 VPWR.n3027 VPWR 0.03175
R6295 VPWR.n3009 VPWR 0.03175
R6296 VPWR VPWR.n3165 0.03175
R6297 VPWR.n3186 VPWR 0.03175
R6298 VPWR VPWR.n3298 0.03175
R6299 VPWR.n3299 VPWR 0.03175
R6300 VPWR.n3375 VPWR 0.03175
R6301 VPWR.n3436 VPWR 0.03175
R6302 VPWR.n3407 VPWR 0.03175
R6303 VPWR.n1341 VPWR 0.03175
R6304 VPWR VPWR.n1149 0.03175
R6305 VPWR.n3727 VPWR 0.03175
R6306 VPWR.n3664 VPWR 0.03175
R6307 VPWR.n3658 VPWR 0.03175
R6308 VPWR.n3604 VPWR 0.03175
R6309 VPWR.n3587 VPWR 0.03175
R6310 VPWR VPWR.n3812 0.03175
R6311 VPWR VPWR.n3909 0.03175
R6312 VPWR VPWR.n3919 0.03175
R6313 VPWR.n3946 VPWR 0.03175
R6314 VPWR VPWR.n4030 0.03175
R6315 VPWR.n4047 VPWR 0.03175
R6316 VPWR.n706 VPWR 0.03175
R6317 VPWR VPWR.n870 0.03175
R6318 VPWR.n871 VPWR 0.03175
R6319 VPWR VPWR.n895 0.03175
R6320 VPWR VPWR.n898 0.03175
R6321 VPWR VPWR.n919 0.03175
R6322 VPWR VPWR.n4290 0.03175
R6323 VPWR VPWR.n4404 0.03175
R6324 VPWR.n4833 VPWR 0.03175
R6325 VPWR.n4725 VPWR 0.03175
R6326 VPWR VPWR.n4766 0.03175
R6327 VPWR VPWR.n4950 0.03175
R6328 VPWR.n4958 VPWR 0.03175
R6329 VPWR VPWR.n4976 0.03175
R6330 VPWR.n5142 VPWR 0.03175
R6331 VPWR.n5115 VPWR 0.03175
R6332 VPWR VPWR.n5177 0.03175
R6333 VPWR VPWR.n5213 0.03175
R6334 VPWR.n5266 VPWR 0.03175
R6335 VPWR.n5242 VPWR 0.03175
R6336 VPWR.n210 VPWR 0.03175
R6337 VPWR VPWR.n571 0.03175
R6338 VPWR VPWR.n597 0.03175
R6339 VPWR.n412 VPWR 0.03175
R6340 VPWR.n392 VPWR 0.03175
R6341 VPWR.n387 VPWR 0.03175
R6342 VPWR.n5362 VPWR 0.03175
R6343 VPWR.n5882 VPWR 0.03175
R6344 VPWR.n6001 VPWR 0.03175
R6345 VPWR.n6019 VPWR 0.03175
R6346 VPWR.n5405 VPWR 0.03175
R6347 VPWR.n5718 VPWR 0.03175
R6348 VPWR.n2438 VPWR 0.03175
R6349 VPWR.n2535 VPWR 0.03175
R6350 VPWR.n2592 VPWR 0.03175
R6351 VPWR VPWR.n2160 0.03175
R6352 VPWR.n6289 VPWR 0.03175
R6353 VPWR.n6228 VPWR 0.03175
R6354 VPWR.n6227 VPWR 0.03175
R6355 VPWR.n6215 VPWR 0.03175
R6356 VPWR VPWR.n6128 0.03175
R6357 VPWR.n6167 VPWR 0.03175
R6358 VPWR.n3080 VPWR.n3079 0.0304479
R6359 VPWR.n3074 VPWR.n3073 0.0304479
R6360 VPWR.n3076 VPWR.n3075 0.0304479
R6361 VPWR.n1759 VPWR.n1758 0.0304479
R6362 VPWR.n1761 VPWR.n1760 0.0304479
R6363 VPWR.n1755 VPWR.n1754 0.0304479
R6364 VPWR.n1398 VPWR.n1397 0.0304479
R6365 VPWR.n1400 VPWR.n1399 0.0304479
R6366 VPWR.n1394 VPWR.n1393 0.0304479
R6367 VPWR.n3548 VPWR.n3547 0.0304479
R6368 VPWR.n1284 VPWR.n1283 0.0304479
R6369 VPWR.n3544 VPWR.n3543 0.0304479
R6370 VPWR.n1058 VPWR.n1057 0.0304479
R6371 VPWR.n1060 VPWR.n1059 0.0304479
R6372 VPWR.n1054 VPWR.n1053 0.0304479
R6373 VPWR.n4346 VPWR.n4345 0.0304479
R6374 VPWR.n4348 VPWR.n4347 0.0304479
R6375 VPWR.n756 VPWR.n755 0.0304479
R6376 VPWR.n4813 VPWR.n4812 0.0304479
R6377 VPWR.n4815 VPWR.n4814 0.0304479
R6378 VPWR.n4482 VPWR.n4481 0.0304479
R6379 VPWR.n306 VPWR.n305 0.0304479
R6380 VPWR.n308 VPWR.n307 0.0304479
R6381 VPWR.n302 VPWR.n301 0.0304479
R6382 VPWR.n5776 VPWR.n5775 0.0304479
R6383 VPWR.n5770 VPWR.n5769 0.0304479
R6384 VPWR.n5772 VPWR.n5771 0.0304479
R6385 VPWR.n5394 VPWR.n5393 0.0304479
R6386 VPWR.n5396 VPWR.n5395 0.0304479
R6387 VPWR.n5390 VPWR.n5389 0.0304479
R6388 VPWR.n2323 VPWR.n2322 0.0304479
R6389 VPWR.n2327 VPWR.n2326 0.0304479
R6390 VPWR.n2321 VPWR.n2320 0.0304479
R6391 VPWR.n6187 VPWR.n6186 0.0304479
R6392 VPWR.n1417 VPWR.n1416 0.0291458
R6393 VPWR VPWR.n4235 0.0291458
R6394 VPWR.n4601 VPWR.n4600 0.0291458
R6395 VPWR VPWR.n676 0.0291458
R6396 VPWR.n5413 VPWR.n5412 0.0291458
R6397 VPWR.n2088 VPWR.n2087 0.0291458
R6398 VPWR.n98 VPWR.n97 0.0291458
R6399 VPWR.n2737 VPWR 0.0283802
R6400 VPWR.n2101 VPWR.n2100 0.0278438
R6401 VPWR.n2363 VPWR.n2362 0.0278438
R6402 VPWR.n2745 VPWR.n2744 0.0278438
R6403 VPWR.n2781 VPWR.n2780 0.0278438
R6404 VPWR.n2784 VPWR.n2783 0.0278438
R6405 VPWR.n2792 VPWR.n2791 0.0278438
R6406 VPWR.n1795 VPWR.n1794 0.0278438
R6407 VPWR.n1915 VPWR.n1914 0.0278438
R6408 VPWR.n1833 VPWR.n1832 0.0278438
R6409 VPWR.n1462 VPWR.n1461 0.0278438
R6410 VPWR.n3289 VPWR.n3288 0.0278438
R6411 VPWR.n1498 VPWR.n1497 0.0278438
R6412 VPWR.n3636 VPWR.n3635 0.0278438
R6413 VPWR.n3756 VPWR.n3755 0.0278438
R6414 VPWR.n1192 VPWR.n1191 0.0278438
R6415 VPWR.n1101 VPWR.n1100 0.0278438
R6416 VPWR.n3854 VPWR.n3853 0.0278438
R6417 VPWR.n3851 VPWR.n3840 0.0278438
R6418 VPWR.n3842 VPWR.n3841 0.0278438
R6419 VPWR.n794 VPWR.n793 0.0278438
R6420 VPWR.n842 VPWR.n841 0.0278438
R6421 VPWR.n838 VPWR.n837 0.0278438
R6422 VPWR.n4632 VPWR.n4631 0.0278438
R6423 VPWR.n4892 VPWR.n4891 0.0278438
R6424 VPWR.n4449 VPWR.n4448 0.0278438
R6425 VPWR.n670 VPWR.n669 0.0278438
R6426 VPWR.n5014 VPWR.n5013 0.0278438
R6427 VPWR.n5011 VPWR.n5000 0.0278438
R6428 VPWR.n5002 VPWR.n5001 0.0278438
R6429 VPWR.n471 VPWR.n470 0.0278438
R6430 VPWR.n515 VPWR.n514 0.0278438
R6431 VPWR.n511 VPWR.n510 0.0278438
R6432 VPWR.n5440 VPWR.n5439 0.0278438
R6433 VPWR.n5921 VPWR.n5920 0.0278438
R6434 VPWR.n5918 VPWR.n5907 0.0278438
R6435 VPWR.n5909 VPWR.n5908 0.0278438
R6436 VPWR.n36 VPWR.n35 0.0278438
R6437 VPWR.n2352 VPWR.n2351 0.0278438
R6438 VPWR.n2355 VPWR.n2354 0.0278438
R6439 VPWR.n6272 VPWR.n6271 0.0278438
R6440 VPWR.n6269 VPWR.n32 0.0278438
R6441 VPWR.n125 VPWR.n124 0.0278438
R6442 VPWR.n1515 VPWR.n1514 0.0272664
R6443 VPWR.n2603 VPWR.n2602 0.0259094
R6444 VPWR.n3064 VPWR.n3063 0.0259094
R6445 VPWR.n3063 VPWR.n3062 0.0259094
R6446 VPWR.n2917 VPWR.n2916 0.0259094
R6447 VPWR.n3123 VPWR.n3122 0.0259094
R6448 VPWR.n3122 VPWR.n3121 0.0259094
R6449 VPWR.n3052 VPWR.n3051 0.0259094
R6450 VPWR.n2924 VPWR.n2923 0.0259094
R6451 VPWR.n3133 VPWR.n3132 0.0259094
R6452 VPWR.n1448 VPWR.n1447 0.0259094
R6453 VPWR.n1447 VPWR.n1446 0.0259094
R6454 VPWR.n3453 VPWR.n3452 0.0259094
R6455 VPWR.n3146 VPWR.n3145 0.0259094
R6456 VPWR.n3145 VPWR.n3144 0.0259094
R6457 VPWR.n1431 VPWR.n1430 0.0259094
R6458 VPWR.n1430 VPWR.n1429 0.0259094
R6459 VPWR.n1305 VPWR.n1304 0.0259094
R6460 VPWR.n3786 VPWR.n3785 0.0259094
R6461 VPWR.n3785 VPWR.n3784 0.0259094
R6462 VPWR.n1087 VPWR.n1086 0.0259094
R6463 VPWR.n1086 VPWR.n1085 0.0259094
R6464 VPWR.n4099 VPWR.n4098 0.0259094
R6465 VPWR.n3799 VPWR.n3798 0.0259094
R6466 VPWR.n3798 VPWR.n3797 0.0259094
R6467 VPWR.n4106 VPWR.n4105 0.0259094
R6468 VPWR.n782 VPWR.n781 0.0259094
R6469 VPWR.n697 VPWR.n696 0.0259094
R6470 VPWR.n4573 VPWR.n4572 0.0259094
R6471 VPWR.n4572 VPWR.n4571 0.0259094
R6472 VPWR.n4612 VPWR.n4611 0.0259094
R6473 VPWR.n4921 VPWR.n4920 0.0259094
R6474 VPWR.n4920 VPWR.n4919 0.0259094
R6475 VPWR.n5288 VPWR.n5287 0.0259094
R6476 VPWR.n5287 VPWR.n5286 0.0259094
R6477 VPWR.n634 VPWR.n633 0.0259094
R6478 VPWR.n4933 VPWR.n4932 0.0259094
R6479 VPWR.n4932 VPWR.n4931 0.0259094
R6480 VPWR.n5760 VPWR.n5759 0.0259094
R6481 VPWR.n5759 VPWR.n5758 0.0259094
R6482 VPWR.n328 VPWR.n327 0.0259094
R6483 VPWR.n5819 VPWR.n5818 0.0259094
R6484 VPWR.n5818 VPWR.n5817 0.0259094
R6485 VPWR.n6070 VPWR.n6069 0.0259094
R6486 VPWR.n6069 VPWR.n6068 0.0259094
R6487 VPWR.n5746 VPWR.n5745 0.0259094
R6488 VPWR.n5851 VPWR.n5850 0.0259094
R6489 VPWR.n5850 VPWR.n5849 0.0259094
R6490 VPWR.n5835 VPWR.n5834 0.0259094
R6491 VPWR.n5834 VPWR.n5833 0.0259094
R6492 VPWR.n2473 VPWR.n2472 0.0259094
R6493 VPWR.n2472 VPWR.n2471 0.0259094
R6494 VPWR.n2216 VPWR.n2215 0.0259094
R6495 VPWR.n2217 VPWR.n2216 0.0259094
R6496 VPWR.n5652 VPWR.n5651 0.0259094
R6497 VPWR.n5651 VPWR.n5650 0.0259094
R6498 VPWR.n111 VPWR.n110 0.0259094
R6499 VPWR.n110 VPWR.n109 0.0259094
R6500 VPWR.n2908 VPWR.n2907 0.0252396
R6501 VPWR.n3077 VPWR 0.0252396
R6502 VPWR VPWR.n1763 0.0252396
R6503 VPWR VPWR.n1402 0.0252396
R6504 VPWR.n3545 VPWR 0.0252396
R6505 VPWR VPWR.n1062 0.0252396
R6506 VPWR VPWR.n4350 0.0252396
R6507 VPWR.n4700 VPWR.n4699 0.0252396
R6508 VPWR VPWR.n4817 0.0252396
R6509 VPWR VPWR.n310 0.0252396
R6510 VPWR.n5773 VPWR 0.0252396
R6511 VPWR.n6060 VPWR.n6059 0.0252396
R6512 VPWR VPWR.n5398 0.0252396
R6513 VPWR.n2596 VPWR.n2595 0.0252396
R6514 VPWR.n2324 VPWR 0.0252396
R6515 VPWR VPWR.n6190 0.0252396
R6516 VPWR.n2057 VPWR.n2056 0.0239375
R6517 VPWR.n2056 VPWR.n2055 0.0239375
R6518 VPWR.n2102 VPWR.n2101 0.0239375
R6519 VPWR.n2386 VPWR.n2385 0.0239375
R6520 VPWR.n3081 VPWR.n3080 0.0239375
R6521 VPWR.n1596 VPWR.n1595 0.0239375
R6522 VPWR.n2760 VPWR.n2759 0.0239375
R6523 VPWR.n2759 VPWR.n2758 0.0239375
R6524 VPWR.n2744 VPWR.n2743 0.0239375
R6525 VPWR.n2910 VPWR 0.0239375
R6526 VPWR.n2752 VPWR.n2751 0.0239375
R6527 VPWR.n1655 VPWR 0.0239375
R6528 VPWR.n3101 VPWR.n3100 0.0239375
R6529 VPWR.n1758 VPWR.n1757 0.0239375
R6530 VPWR.n1678 VPWR.n1677 0.0239375
R6531 VPWR.n1810 VPWR.n1809 0.0239375
R6532 VPWR.n1809 VPWR.n1808 0.0239375
R6533 VPWR.n1794 VPWR.n1793 0.0239375
R6534 VPWR.n1821 VPWR 0.0239375
R6535 VPWR.n2033 VPWR 0.0239375
R6536 VPWR.n1802 VPWR.n1801 0.0239375
R6537 VPWR.n1739 VPWR 0.0239375
R6538 VPWR.n1899 VPWR.n1898 0.0239375
R6539 VPWR.n1477 VPWR.n1476 0.0239375
R6540 VPWR.n1476 VPWR.n1475 0.0239375
R6541 VPWR.n1461 VPWR.n1460 0.0239375
R6542 VPWR.n1397 VPWR.n1396 0.0239375
R6543 VPWR.n1384 VPWR.n1383 0.0239375
R6544 VPWR.n3176 VPWR 0.0239375
R6545 VPWR.n3259 VPWR 0.0239375
R6546 VPWR.n3344 VPWR 0.0239375
R6547 VPWR.n1469 VPWR.n1468 0.0239375
R6548 VPWR.n3203 VPWR.n3202 0.0239375
R6549 VPWR.n3651 VPWR.n3650 0.0239375
R6550 VPWR.n3650 VPWR.n3649 0.0239375
R6551 VPWR.n3635 VPWR.n3634 0.0239375
R6552 VPWR.n3549 VPWR.n3548 0.0239375
R6553 VPWR.n3534 VPWR.n3533 0.0239375
R6554 VPWR VPWR.n3654 0.0239375
R6555 VPWR.n3643 VPWR.n3642 0.0239375
R6556 VPWR.n3627 VPWR 0.0239375
R6557 VPWR.n3764 VPWR.n3763 0.0239375
R6558 VPWR.n1116 VPWR.n1115 0.0239375
R6559 VPWR.n1115 VPWR.n1114 0.0239375
R6560 VPWR.n1100 VPWR.n1099 0.0239375
R6561 VPWR.n1057 VPWR.n1056 0.0239375
R6562 VPWR.n979 VPWR.n978 0.0239375
R6563 VPWR.n1127 VPWR 0.0239375
R6564 VPWR.n3978 VPWR 0.0239375
R6565 VPWR.n1108 VPWR.n1107 0.0239375
R6566 VPWR.n1008 VPWR 0.0239375
R6567 VPWR.n3863 VPWR.n3862 0.0239375
R6568 VPWR.n4345 VPWR.n4344 0.0239375
R6569 VPWR.n4133 VPWR.n4132 0.0239375
R6570 VPWR.n809 VPWR.n808 0.0239375
R6571 VPWR.n808 VPWR.n807 0.0239375
R6572 VPWR.n793 VPWR.n792 0.0239375
R6573 VPWR.n952 VPWR 0.0239375
R6574 VPWR.n801 VPWR.n800 0.0239375
R6575 VPWR.n4252 VPWR 0.0239375
R6576 VPWR.n4277 VPWR 0.0239375
R6577 VPWR.n4192 VPWR 0.0239375
R6578 VPWR.n4368 VPWR.n4367 0.0239375
R6579 VPWR.n4812 VPWR.n4811 0.0239375
R6580 VPWR.n4501 VPWR.n4500 0.0239375
R6581 VPWR.n4647 VPWR.n4646 0.0239375
R6582 VPWR.n4646 VPWR.n4645 0.0239375
R6583 VPWR.n4631 VPWR.n4630 0.0239375
R6584 VPWR.n4872 VPWR 0.0239375
R6585 VPWR.n4680 VPWR 0.0239375
R6586 VPWR.n4702 VPWR 0.0239375
R6587 VPWR.n4639 VPWR.n4638 0.0239375
R6588 VPWR.n4717 VPWR 0.0239375
R6589 VPWR.n4585 VPWR 0.0239375
R6590 VPWR.n4543 VPWR 0.0239375
R6591 VPWR.n4899 VPWR.n4898 0.0239375
R6592 VPWR.n305 VPWR.n304 0.0239375
R6593 VPWR.n247 VPWR.n246 0.0239375
R6594 VPWR.n650 VPWR.n649 0.0239375
R6595 VPWR.n651 VPWR.n650 0.0239375
R6596 VPWR.n669 VPWR.n668 0.0239375
R6597 VPWR.n5043 VPWR 0.0239375
R6598 VPWR.n5150 VPWR 0.0239375
R6599 VPWR.n661 VPWR.n660 0.0239375
R6600 VPWR.n5021 VPWR.n5020 0.0239375
R6601 VPWR.n5777 VPWR.n5776 0.0239375
R6602 VPWR.n5310 VPWR.n5309 0.0239375
R6603 VPWR.n486 VPWR.n485 0.0239375
R6604 VPWR.n485 VPWR.n484 0.0239375
R6605 VPWR.n470 VPWR.n469 0.0239375
R6606 VPWR.n620 VPWR 0.0239375
R6607 VPWR.n478 VPWR.n477 0.0239375
R6608 VPWR.n5351 VPWR 0.0239375
R6609 VPWR.n5342 VPWR 0.0239375
R6610 VPWR.n5797 VPWR.n5796 0.0239375
R6611 VPWR.n5423 VPWR.n5422 0.0239375
R6612 VPWR.n5424 VPWR.n5423 0.0239375
R6613 VPWR.n5441 VPWR.n5440 0.0239375
R6614 VPWR.n5393 VPWR.n5392 0.0239375
R6615 VPWR.n5680 VPWR.n5679 0.0239375
R6616 VPWR.n5987 VPWR 0.0239375
R6617 VPWR.n6062 VPWR 0.0239375
R6618 VPWR.n5433 VPWR.n5432 0.0239375
R6619 VPWR.n5726 VPWR 0.0239375
R6620 VPWR.n5938 VPWR.n5937 0.0239375
R6621 VPWR.n6282 VPWR.n6281 0.0239375
R6622 VPWR.n35 VPWR.n34 0.0239375
R6623 VPWR.n2328 VPWR.n2327 0.0239375
R6624 VPWR.n2237 VPWR.n2236 0.0239375
R6625 VPWR.n6186 VPWR.n6185 0.0239375
R6626 VPWR.n5569 VPWR.n5568 0.0239375
R6627 VPWR.n5582 VPWR.n5581 0.0239375
R6628 VPWR.n132 VPWR.n131 0.0239375
R6629 VPWR.n140 VPWR.n139 0.0239375
R6630 VPWR.n139 VPWR.n138 0.0239375
R6631 VPWR.n124 VPWR.n123 0.0239375
R6632 VPWR.n3089 VPWR 0.0237788
R6633 VPWR.n3441 VPWR 0.0237788
R6634 VPWR VPWR.n1294 0.0237788
R6635 VPWR.n5272 VPWR 0.0237788
R6636 VPWR.n2336 VPWR 0.0237788
R6637 VPWR.n6191 VPWR 0.0237788
R6638 VPWR.n1597 VPWR.n1596 0.0226354
R6639 VPWR VPWR.n1533 0.0226354
R6640 VPWR.n1539 VPWR 0.0226354
R6641 VPWR VPWR.n1544 0.0226354
R6642 VPWR VPWR.n1545 0.0226354
R6643 VPWR.n2837 VPWR 0.0226354
R6644 VPWR.n2842 VPWR 0.0226354
R6645 VPWR.n2848 VPWR 0.0226354
R6646 VPWR.n2774 VPWR 0.0226354
R6647 VPWR.n2864 VPWR 0.0226354
R6648 VPWR.n2890 VPWR 0.0226354
R6649 VPWR VPWR.n2902 0.0226354
R6650 VPWR.n2630 VPWR.n2625 0.0226354
R6651 VPWR.n2736 VPWR 0.0226354
R6652 VPWR.n2729 VPWR 0.0226354
R6653 VPWR.n2726 VPWR 0.0226354
R6654 VPWR.n2717 VPWR 0.0226354
R6655 VPWR.n2698 VPWR 0.0226354
R6656 VPWR.n2692 VPWR 0.0226354
R6657 VPWR.n2685 VPWR 0.0226354
R6658 VPWR.n2682 VPWR 0.0226354
R6659 VPWR.n2672 VPWR 0.0226354
R6660 VPWR VPWR 0.0226354
R6661 VPWR.n2655 VPWR 0.0226354
R6662 VPWR.n1658 VPWR 0.0226354
R6663 VPWR.n1644 VPWR 0.0226354
R6664 VPWR.n1638 VPWR 0.0226354
R6665 VPWR.n1637 VPWR 0.0226354
R6666 VPWR.n1632 VPWR 0.0226354
R6667 VPWR.n1631 VPWR 0.0226354
R6668 VPWR.n1627 VPWR 0.0226354
R6669 VPWR.n1626 VPWR 0.0226354
R6670 VPWR.n1679 VPWR.n1678 0.0226354
R6671 VPWR VPWR.n1853 0.0226354
R6672 VPWR.n1865 VPWR 0.0226354
R6673 VPWR.n1840 VPWR 0.0226354
R6674 VPWR.n1937 VPWR 0.0226354
R6675 VPWR.n1819 VPWR 0.0226354
R6676 VPWR.n1949 VPWR 0.0226354
R6677 VPWR VPWR.n1969 0.0226354
R6678 VPWR VPWR.n1970 0.0226354
R6679 VPWR.n2020 VPWR 0.0226354
R6680 VPWR.n1982 VPWR 0.0226354
R6681 VPWR.n2948 VPWR 0.0226354
R6682 VPWR.n2955 VPWR 0.0226354
R6683 VPWR VPWR.n2968 0.0226354
R6684 VPWR.n2969 VPWR 0.0226354
R6685 VPWR VPWR.n2990 0.0226354
R6686 VPWR.n3023 VPWR 0.0226354
R6687 VPWR.n3018 VPWR 0.0226354
R6688 VPWR.n3012 VPWR 0.0226354
R6689 VPWR.n3007 VPWR 0.0226354
R6690 VPWR.n1742 VPWR 0.0226354
R6691 VPWR.n1729 VPWR 0.0226354
R6692 VPWR.n1726 VPWR 0.0226354
R6693 VPWR.n1716 VPWR 0.0226354
R6694 VPWR.n1712 VPWR 0.0226354
R6695 VPWR.n1705 VPWR 0.0226354
R6696 VPWR.n1383 VPWR.n1382 0.0226354
R6697 VPWR.n3167 VPWR 0.0226354
R6698 VPWR VPWR.n3174 0.0226354
R6699 VPWR VPWR.n3175 0.0226354
R6700 VPWR.n3269 VPWR 0.0226354
R6701 VPWR.n3266 VPWR 0.0226354
R6702 VPWR.n3263 VPWR 0.0226354
R6703 VPWR.n3246 VPWR 0.0226354
R6704 VPWR.n3241 VPWR 0.0226354
R6705 VPWR.n3307 VPWR 0.0226354
R6706 VPWR VPWR.n3328 0.0226354
R6707 VPWR.n1487 VPWR 0.0226354
R6708 VPWR.n1416 VPWR.n1415 0.0226354
R6709 VPWR.n3367 VPWR 0.0226354
R6710 VPWR VPWR.n3370 0.0226354
R6711 VPWR VPWR.n3371 0.0226354
R6712 VPWR VPWR.n3387 0.0226354
R6713 VPWR VPWR.n3389 0.0226354
R6714 VPWR VPWR.n3390 0.0226354
R6715 VPWR.n3429 VPWR 0.0226354
R6716 VPWR.n3424 VPWR 0.0226354
R6717 VPWR.n3417 VPWR 0.0226354
R6718 VPWR.n3416 VPWR 0.0226354
R6719 VPWR VPWR.n3402 0.0226354
R6720 VPWR.n1373 VPWR 0.0226354
R6721 VPWR.n1370 VPWR 0.0226354
R6722 VPWR.n1360 VPWR 0.0226354
R6723 VPWR.n1354 VPWR 0.0226354
R6724 VPWR.n1346 VPWR 0.0226354
R6725 VPWR VPWR.n1336 0.0226354
R6726 VPWR.n3533 VPWR.n3532 0.0226354
R6727 VPWR VPWR.n1152 0.0226354
R6728 VPWR.n1153 VPWR 0.0226354
R6729 VPWR.n3736 VPWR 0.0226354
R6730 VPWR.n3733 VPWR 0.0226354
R6731 VPWR.n3730 VPWR 0.0226354
R6732 VPWR.n3718 VPWR 0.0226354
R6733 VPWR VPWR.n1221 0.0226354
R6734 VPWR.n3700 VPWR 0.0226354
R6735 VPWR.n3695 VPWR 0.0226354
R6736 VPWR.n3672 VPWR 0.0226354
R6737 VPWR.n3669 VPWR 0.0226354
R6738 VPWR.n3667 VPWR 0.0226354
R6739 VPWR.n3655 VPWR 0.0226354
R6740 VPWR.n3622 VPWR 0.0226354
R6741 VPWR.n3596 VPWR 0.0226354
R6742 VPWR.n3590 VPWR 0.0226354
R6743 VPWR.n3579 VPWR 0.0226354
R6744 VPWR.n3573 VPWR 0.0226354
R6745 VPWR.n3566 VPWR 0.0226354
R6746 VPWR.n3519 VPWR 0.0226354
R6747 VPWR.n3496 VPWR 0.0226354
R6748 VPWR.n3489 VPWR 0.0226354
R6749 VPWR.n3485 VPWR 0.0226354
R6750 VPWR.n980 VPWR.n979 0.0226354
R6751 VPWR.n3811 VPWR 0.0226354
R6752 VPWR VPWR.n3831 0.0226354
R6753 VPWR VPWR.n3893 0.0226354
R6754 VPWR VPWR.n3894 0.0226354
R6755 VPWR.n3902 VPWR 0.0226354
R6756 VPWR VPWR.n3908 0.0226354
R6757 VPWR.n3910 VPWR 0.0226354
R6758 VPWR VPWR.n3918 0.0226354
R6759 VPWR.n3962 VPWR 0.0226354
R6760 VPWR.n3950 VPWR 0.0226354
R6761 VPWR.n3947 VPWR 0.0226354
R6762 VPWR.n3940 VPWR 0.0226354
R6763 VPWR.n3939 VPWR 0.0226354
R6764 VPWR.n3935 VPWR 0.0226354
R6765 VPWR.n3998 VPWR 0.0226354
R6766 VPWR VPWR.n4011 0.0226354
R6767 VPWR.n4013 VPWR 0.0226354
R6768 VPWR.n4078 VPWR 0.0226354
R6769 VPWR.n4077 VPWR 0.0226354
R6770 VPWR.n4063 VPWR 0.0226354
R6771 VPWR.n4060 VPWR 0.0226354
R6772 VPWR.n4043 VPWR 0.0226354
R6773 VPWR.n1037 VPWR 0.0226354
R6774 VPWR.n1024 VPWR 0.0226354
R6775 VPWR.n1011 VPWR 0.0226354
R6776 VPWR.n1006 VPWR 0.0226354
R6777 VPWR.n4134 VPWR.n4133 0.0226354
R6778 VPWR VPWR.n719 0.0226354
R6779 VPWR.n722 VPWR 0.0226354
R6780 VPWR.n734 VPWR 0.0226354
R6781 VPWR.n865 VPWR 0.0226354
R6782 VPWR.n826 VPWR 0.0226354
R6783 VPWR VPWR.n869 0.0226354
R6784 VPWR.n879 VPWR 0.0226354
R6785 VPWR VPWR.n883 0.0226354
R6786 VPWR VPWR.n885 0.0226354
R6787 VPWR.n886 VPWR 0.0226354
R6788 VPWR.n903 VPWR 0.0226354
R6789 VPWR.n920 VPWR 0.0226354
R6790 VPWR.n928 VPWR 0.0226354
R6791 VPWR VPWR.n947 0.0226354
R6792 VPWR.n4236 VPWR 0.0226354
R6793 VPWR VPWR.n4251 0.0226354
R6794 VPWR.n4265 VPWR 0.0226354
R6795 VPWR VPWR.n4276 0.0226354
R6796 VPWR VPWR.n4280 0.0226354
R6797 VPWR VPWR.n4289 0.0226354
R6798 VPWR.n4308 VPWR 0.0226354
R6799 VPWR VPWR.n4322 0.0226354
R6800 VPWR.n4323 VPWR 0.0226354
R6801 VPWR.n4329 VPWR 0.0226354
R6802 VPWR VPWR.n4335 0.0226354
R6803 VPWR VPWR.n4338 0.0226354
R6804 VPWR.n4197 VPWR 0.0226354
R6805 VPWR.n4194 VPWR 0.0226354
R6806 VPWR.n4193 VPWR 0.0226354
R6807 VPWR.n4184 VPWR 0.0226354
R6808 VPWR.n4181 VPWR 0.0226354
R6809 VPWR.n4170 VPWR 0.0226354
R6810 VPWR.n4156 VPWR 0.0226354
R6811 VPWR.n4502 VPWR.n4501 0.0226354
R6812 VPWR VPWR.n4417 0.0226354
R6813 VPWR.n4420 VPWR 0.0226354
R6814 VPWR.n4432 VPWR 0.0226354
R6815 VPWR.n4875 VPWR 0.0226354
R6816 VPWR.n4871 VPWR 0.0226354
R6817 VPWR.n4863 VPWR 0.0226354
R6818 VPWR.n4860 VPWR 0.0226354
R6819 VPWR.n4851 VPWR 0.0226354
R6820 VPWR.n4840 VPWR 0.0226354
R6821 VPWR.n4837 VPWR 0.0226354
R6822 VPWR.n4664 VPWR 0.0226354
R6823 VPWR VPWR.n4689 0.0226354
R6824 VPWR.n4690 VPWR 0.0226354
R6825 VPWR.n4696 VPWR 0.0226354
R6826 VPWR.n4600 VPWR.n4599 0.0226354
R6827 VPWR VPWR.n4715 0.0226354
R6828 VPWR VPWR.n4716 0.0226354
R6829 VPWR.n4734 VPWR 0.0226354
R6830 VPWR.n4749 VPWR 0.0226354
R6831 VPWR VPWR.n4765 0.0226354
R6832 VPWR.n4586 VPWR 0.0226354
R6833 VPWR.n4780 VPWR 0.0226354
R6834 VPWR VPWR.n4787 0.0226354
R6835 VPWR VPWR.n4793 0.0226354
R6836 VPWR.n4794 VPWR 0.0226354
R6837 VPWR.n4562 VPWR 0.0226354
R6838 VPWR.n4559 VPWR 0.0226354
R6839 VPWR.n4554 VPWR 0.0226354
R6840 VPWR.n4546 VPWR 0.0226354
R6841 VPWR.n4528 VPWR 0.0226354
R6842 VPWR.n248 VPWR.n247 0.0226354
R6843 VPWR VPWR.n4957 0.0226354
R6844 VPWR VPWR.n4963 0.0226354
R6845 VPWR.n4966 VPWR 0.0226354
R6846 VPWR.n4940 VPWR 0.0226354
R6847 VPWR.n4973 VPWR 0.0226354
R6848 VPWR.n4978 VPWR 0.0226354
R6849 VPWR.n5057 VPWR 0.0226354
R6850 VPWR.n5059 VPWR 0.0226354
R6851 VPWR.n5070 VPWR 0.0226354
R6852 VPWR.n5084 VPWR 0.0226354
R6853 VPWR VPWR.n5096 0.0226354
R6854 VPWR.n5140 VPWR 0.0226354
R6855 VPWR.n5138 VPWR 0.0226354
R6856 VPWR.n5135 VPWR 0.0226354
R6857 VPWR.n5132 VPWR 0.0226354
R6858 VPWR.n5128 VPWR 0.0226354
R6859 VPWR.n5127 VPWR 0.0226354
R6860 VPWR.n5124 VPWR 0.0226354
R6861 VPWR.n5120 VPWR 0.0226354
R6862 VPWR.n5118 VPWR 0.0226354
R6863 VPWR VPWR.n674 0.0226354
R6864 VPWR.n5164 VPWR 0.0226354
R6865 VPWR VPWR.n5170 0.0226354
R6866 VPWR VPWR.n5178 0.0226354
R6867 VPWR.n5179 VPWR 0.0226354
R6868 VPWR.n5187 VPWR 0.0226354
R6869 VPWR VPWR.n5212 0.0226354
R6870 VPWR.n5260 VPWR 0.0226354
R6871 VPWR.n5258 VPWR 0.0226354
R6872 VPWR.n5238 VPWR 0.0226354
R6873 VPWR.n5233 VPWR 0.0226354
R6874 VPWR.n5232 VPWR 0.0226354
R6875 VPWR.n5227 VPWR 0.0226354
R6876 VPWR.n286 VPWR 0.0226354
R6877 VPWR.n279 VPWR 0.0226354
R6878 VPWR.n5311 VPWR.n5310 0.0226354
R6879 VPWR.n197 VPWR 0.0226354
R6880 VPWR VPWR.n205 0.0226354
R6881 VPWR.n189 VPWR 0.0226354
R6882 VPWR.n534 VPWR 0.0226354
R6883 VPWR.n538 VPWR 0.0226354
R6884 VPWR VPWR.n541 0.0226354
R6885 VPWR.n543 VPWR 0.0226354
R6886 VPWR VPWR.n550 0.0226354
R6887 VPWR.n551 VPWR 0.0226354
R6888 VPWR VPWR.n558 0.0226354
R6889 VPWR.n559 VPWR 0.0226354
R6890 VPWR.n497 VPWR 0.0226354
R6891 VPWR VPWR.n572 0.0226354
R6892 VPWR.n583 VPWR 0.0226354
R6893 VPWR VPWR.n586 0.0226354
R6894 VPWR VPWR.n587 0.0226354
R6895 VPWR.n588 VPWR 0.0226354
R6896 VPWR.n601 VPWR 0.0226354
R6897 VPWR VPWR.n615 0.0226354
R6898 VPWR.n346 VPWR.n340 0.0226354
R6899 VPWR.n453 VPWR 0.0226354
R6900 VPWR.n438 VPWR 0.0226354
R6901 VPWR.n429 VPWR 0.0226354
R6902 VPWR VPWR.n356 0.0226354
R6903 VPWR.n423 VPWR 0.0226354
R6904 VPWR.n414 VPWR 0.0226354
R6905 VPWR.n405 VPWR 0.0226354
R6906 VPWR.n393 VPWR 0.0226354
R6907 VPWR VPWR.n367 0.0226354
R6908 VPWR.n385 VPWR 0.0226354
R6909 VPWR.n378 VPWR 0.0226354
R6910 VPWR.n375 VPWR 0.0226354
R6911 VPWR.n5371 VPWR 0.0226354
R6912 VPWR.n5354 VPWR 0.0226354
R6913 VPWR VPWR.n5333 0.0226354
R6914 VPWR.n5339 VPWR 0.0226354
R6915 VPWR.n5679 VPWR.n5678 0.0226354
R6916 VPWR.n5870 VPWR 0.0226354
R6917 VPWR.n5862 VPWR 0.0226354
R6918 VPWR.n5876 VPWR 0.0226354
R6919 VPWR VPWR.n5880 0.0226354
R6920 VPWR VPWR.n5881 0.0226354
R6921 VPWR VPWR.n5899 0.0226354
R6922 VPWR.n5978 VPWR 0.0226354
R6923 VPWR VPWR.n5986 0.0226354
R6924 VPWR VPWR.n6000 0.0226354
R6925 VPWR VPWR.n6012 0.0226354
R6926 VPWR VPWR.n6018 0.0226354
R6927 VPWR.n6032 VPWR 0.0226354
R6928 VPWR.n6049 VPWR 0.0226354
R6929 VPWR.n6056 VPWR 0.0226354
R6930 VPWR.n5412 VPWR.n5410 0.0226354
R6931 VPWR.n5462 VPWR 0.0226354
R6932 VPWR VPWR.n5487 0.0226354
R6933 VPWR.n5488 VPWR 0.0226354
R6934 VPWR VPWR.n5495 0.0226354
R6935 VPWR.n5503 VPWR 0.0226354
R6936 VPWR VPWR.n5514 0.0226354
R6937 VPWR.n5523 VPWR 0.0226354
R6938 VPWR VPWR.n5528 0.0226354
R6939 VPWR.n5536 VPWR 0.0226354
R6940 VPWR.n5544 VPWR 0.0226354
R6941 VPWR.n5553 VPWR 0.0226354
R6942 VPWR.n5729 VPWR 0.0226354
R6943 VPWR.n5722 VPWR 0.0226354
R6944 VPWR.n5704 VPWR 0.0226354
R6945 VPWR.n2409 VPWR 0.0226354
R6946 VPWR.n2421 VPWR 0.0226354
R6947 VPWR VPWR.n2437 0.0226354
R6948 VPWR.n2481 VPWR 0.0226354
R6949 VPWR VPWR.n2519 0.0226354
R6950 VPWR VPWR.n2534 0.0226354
R6951 VPWR VPWR.n2544 0.0226354
R6952 VPWR.n2545 VPWR 0.0226354
R6953 VPWR VPWR.n2555 0.0226354
R6954 VPWR.n2556 VPWR 0.0226354
R6955 VPWR VPWR.n2591 0.0226354
R6956 VPWR.n2087 VPWR.n2086 0.0226354
R6957 VPWR.n2111 VPWR 0.0226354
R6958 VPWR.n2126 VPWR 0.0226354
R6959 VPWR.n2076 VPWR 0.0226354
R6960 VPWR VPWR.n2141 0.0226354
R6961 VPWR.n2142 VPWR 0.0226354
R6962 VPWR VPWR.n2159 0.0226354
R6963 VPWR.n2165 VPWR 0.0226354
R6964 VPWR.n2205 VPWR 0.0226354
R6965 VPWR VPWR.n2211 0.0226354
R6966 VPWR.n2304 VPWR 0.0226354
R6967 VPWR.n2284 VPWR 0.0226354
R6968 VPWR.n2267 VPWR 0.0226354
R6969 VPWR.n2238 VPWR.n2237 0.0226354
R6970 VPWR.n5583 VPWR.n5582 0.0226354
R6971 VPWR.n6292 VPWR 0.0226354
R6972 VPWR.n6258 VPWR 0.0226354
R6973 VPWR.n6252 VPWR 0.0226354
R6974 VPWR.n6244 VPWR 0.0226354
R6975 VPWR.n6241 VPWR 0.0226354
R6976 VPWR.n6231 VPWR 0.0226354
R6977 VPWR.n6221 VPWR 0.0226354
R6978 VPWR.n6206 VPWR 0.0226354
R6979 VPWR.n6199 VPWR 0.0226354
R6980 VPWR.n97 VPWR.n96 0.0226354
R6981 VPWR VPWR.n6093 0.0226354
R6982 VPWR.n6103 VPWR 0.0226354
R6983 VPWR.n90 VPWR 0.0226354
R6984 VPWR.n6111 VPWR 0.0226354
R6985 VPWR.n6117 VPWR 0.0226354
R6986 VPWR VPWR.n6127 0.0226354
R6987 VPWR VPWR.n6138 0.0226354
R6988 VPWR VPWR.n6146 0.0226354
R6989 VPWR.n6156 VPWR 0.0226354
R6990 VPWR VPWR.n6166 0.0226354
R6991 VPWR VPWR.n6177 0.0226354
R6992 VPWR.n5631 VPWR 0.0226354
R6993 VPWR.n5616 VPWR 0.0226354
R6994 VPWR.n5602 VPWR 0.0226354
R6995 VPWR.n5598 VPWR 0.0226354
R6996 VPWR.n2093 VPWR.n2092 0.0213333
R6997 VPWR.n2367 VPWR.n2366 0.0213333
R6998 VPWR.n2369 VPWR.n2368 0.0213333
R6999 VPWR.n2628 VPWR.n2627 0.0213333
R7000 VPWR.n2750 VPWR.n2749 0.0213333
R7001 VPWR.n2668 VPWR 0.0213333
R7002 VPWR.n1662 VPWR.n1661 0.0213333
R7003 VPWR.n2796 VPWR.n2795 0.0213333
R7004 VPWR.n2798 VPWR.n2797 0.0213333
R7005 VPWR.n1791 VPWR.n1790 0.0213333
R7006 VPWR.n1876 VPWR 0.0213333
R7007 VPWR VPWR.n1963 0.0213333
R7008 VPWR.n1800 VPWR.n1799 0.0213333
R7009 VPWR.n1746 VPWR.n1745 0.0213333
R7010 VPWR.n1920 VPWR.n1919 0.0213333
R7011 VPWR.n1922 VPWR.n1921 0.0213333
R7012 VPWR.n1458 VPWR.n1457 0.0213333
R7013 VPWR.n3319 VPWR 0.0213333
R7014 VPWR.n3338 VPWR 0.0213333
R7015 VPWR.n1467 VPWR.n1466 0.0213333
R7016 VPWR.n3423 VPWR 0.0213333
R7017 VPWR.n1377 VPWR.n1376 0.0213333
R7018 VPWR.n3284 VPWR.n3283 0.0213333
R7019 VPWR.n3282 VPWR.n3281 0.0213333
R7020 VPWR.n1243 VPWR.n1242 0.0213333
R7021 VPWR VPWR.n1161 0.0213333
R7022 VPWR.n1172 VPWR 0.0213333
R7023 VPWR.n3722 VPWR 0.0213333
R7024 VPWR.n3710 VPWR 0.0213333
R7025 VPWR.n3707 VPWR 0.0213333
R7026 VPWR.n3678 VPWR 0.0213333
R7027 VPWR.n3641 VPWR.n3640 0.0213333
R7028 VPWR.n3607 VPWR 0.0213333
R7029 VPWR.n3583 VPWR 0.0213333
R7030 VPWR.n3570 VPWR 0.0213333
R7031 VPWR.n3558 VPWR 0.0213333
R7032 VPWR.n3527 VPWR.n3526 0.0213333
R7033 VPWR.n3504 VPWR 0.0213333
R7034 VPWR.n3751 VPWR.n3750 0.0213333
R7035 VPWR.n3749 VPWR.n3748 0.0213333
R7036 VPWR.n1097 VPWR.n1096 0.0213333
R7037 VPWR.n3821 VPWR 0.0213333
R7038 VPWR.n3943 VPWR 0.0213333
R7039 VPWR.n1106 VPWR.n1105 0.0213333
R7040 VPWR VPWR.n4029 0.0213333
R7041 VPWR.n4066 VPWR 0.0213333
R7042 VPWR VPWR 0.0213333
R7043 VPWR.n1041 VPWR.n1040 0.0213333
R7044 VPWR.n3849 VPWR.n3848 0.0213333
R7045 VPWR.n3847 VPWR.n3846 0.0213333
R7046 VPWR.n790 VPWR.n789 0.0213333
R7047 VPWR.n913 VPWR 0.0213333
R7048 VPWR VPWR.n918 0.0213333
R7049 VPWR.n937 VPWR 0.0213333
R7050 VPWR.n799 VPWR.n798 0.0213333
R7051 VPWR.n4201 VPWR.n4200 0.0213333
R7052 VPWR.n847 VPWR.n846 0.0213333
R7053 VPWR.n849 VPWR.n848 0.0213333
R7054 VPWR.n4628 VPWR.n4627 0.0213333
R7055 VPWR.n4835 VPWR 0.0213333
R7056 VPWR VPWR.n4694 0.0213333
R7057 VPWR.n4637 VPWR.n4636 0.0213333
R7058 VPWR VPWR.n4768 0.0213333
R7059 VPWR VPWR.n4805 0.0213333
R7060 VPWR.n4564 VPWR.n4563 0.0213333
R7061 VPWR.n4887 VPWR.n4886 0.0213333
R7062 VPWR.n4885 VPWR.n4884 0.0213333
R7063 VPWR.n666 VPWR.n665 0.0213333
R7064 VPWR VPWR.n682 0.0213333
R7065 VPWR.n663 VPWR.n662 0.0213333
R7066 VPWR.n5171 VPWR 0.0213333
R7067 VPWR.n5203 VPWR 0.0213333
R7068 VPWR.n5249 VPWR 0.0213333
R7069 VPWR.n294 VPWR.n293 0.0213333
R7070 VPWR.n5009 VPWR.n5008 0.0213333
R7071 VPWR.n5007 VPWR.n5006 0.0213333
R7072 VPWR.n343 VPWR.n342 0.0213333
R7073 VPWR.n576 VPWR 0.0213333
R7074 VPWR.n605 VPWR 0.0213333
R7075 VPWR.n476 VPWR.n475 0.0213333
R7076 VPWR.n432 VPWR 0.0213333
R7077 VPWR.n5375 VPWR.n5374 0.0213333
R7078 VPWR.n520 VPWR.n519 0.0213333
R7079 VPWR.n522 VPWR.n521 0.0213333
R7080 VPWR.n5418 VPWR.n5417 0.0213333
R7081 VPWR VPWR.n6048 0.0213333
R7082 VPWR.n5435 VPWR.n5434 0.0213333
R7083 VPWR.n5478 VPWR 0.0213333
R7084 VPWR.n5741 VPWR.n5740 0.0213333
R7085 VPWR.n5916 VPWR.n5915 0.0213333
R7086 VPWR.n5914 VPWR.n5913 0.0213333
R7087 VPWR.n6267 VPWR.n6266 0.0213333
R7088 VPWR.n6265 VPWR.n6264 0.0213333
R7089 VPWR.n2096 VPWR.n2095 0.0213333
R7090 VPWR.n2308 VPWR.n2307 0.0213333
R7091 VPWR.n6201 VPWR 0.0213333
R7092 VPWR.n130 VPWR.n129 0.0213333
R7093 VPWR.n6149 VPWR 0.0213333
R7094 VPWR VPWR 0.0213333
R7095 VPWR.n121 VPWR.n120 0.0213333
R7096 VPWR.n5824 VPWR.n5823 0.0207687
R7097 VPWR.n5753 VPWR.n5751 0.0207687
R7098 VPWR.n323 VPWR.n322 0.0207687
R7099 VPWR.n1581 VPWR.n1580 0.0202124
R7100 VPWR.n2804 VPWR.n2803 0.0202124
R7101 VPWR.n1423 VPWR.n1422 0.0202124
R7102 VPWR.n1502 VPWR.n1501 0.0202124
R7103 VPWR.n1437 VPWR.n1436 0.0202124
R7104 VPWR.n1196 VPWR.n1195 0.0202124
R7105 VPWR.n1077 VPWR.n1076 0.0202124
R7106 VPWR.n1135 VPWR.n1134 0.0202124
R7107 VPWR.n4486 VPWR.n4485 0.0202124
R7108 VPWR.n4453 VPWR.n4452 0.0202124
R7109 VPWR.n232 VPWR.n231 0.0202124
R7110 VPWR.n687 VPWR.n686 0.0202124
R7111 VPWR.n5295 VPWR.n5294 0.0202124
R7112 VPWR.n528 VPWR.n527 0.0202124
R7113 VPWR.n5447 VPWR.n5446 0.0202124
R7114 VPWR.n178 VPWR.n177 0.0202124
R7115 VPWR.n5839 VPWR.n5838 0.0202124
R7116 VPWR.n5830 VPWR.n5829 0.0202124
R7117 VPWR.n2466 VPWR.n2465 0.0202124
R7118 VPWR.n2375 VPWR.n2374 0.0202124
R7119 VPWR.n2316 VPWR.n2315 0.0202124
R7120 VPWR.n5647 VPWR.n5646 0.0202124
R7121 VPWR.n5566 VPWR.n5565 0.0202124
R7122 VPWR.n105 VPWR.n104 0.0202124
R7123 VPWR.n2058 VPWR.n2057 0.0200312
R7124 VPWR.n2385 VPWR.n2384 0.0200312
R7125 VPWR.n2371 VPWR.n2370 0.0200312
R7126 VPWR.n1599 VPWR.n1598 0.0200312
R7127 VPWR.n2761 VPWR.n2760 0.0200312
R7128 VPWR.n2789 VPWR.n2788 0.0200312
R7129 VPWR.n2909 VPWR.n2908 0.0200312
R7130 VPWR.n2631 VPWR 0.0200312
R7131 VPWR.n1604 VPWR.n1603 0.0200312
R7132 VPWR.n3102 VPWR.n3101 0.0200312
R7133 VPWR.n2800 VPWR.n2799 0.0200312
R7134 VPWR.n1681 VPWR.n1680 0.0200312
R7135 VPWR.n1811 VPWR.n1810 0.0200312
R7136 VPWR.n1830 VPWR.n1829 0.0200312
R7137 VPWR.n2032 VPWR.n2031 0.0200312
R7138 VPWR VPWR.n1786 0.0200312
R7139 VPWR.n1686 VPWR.n1685 0.0200312
R7140 VPWR.n1900 VPWR.n1899 0.0200312
R7141 VPWR.n1924 VPWR.n1923 0.0200312
R7142 VPWR.n1478 VPWR.n1477 0.0200312
R7143 VPWR.n1381 VPWR.n1380 0.0200312
R7144 VPWR.n3231 VPWR.n3230 0.0200312
R7145 VPWR.n3343 VPWR.n3342 0.0200312
R7146 VPWR.n1326 VPWR.n1325 0.0200312
R7147 VPWR.n3204 VPWR.n3203 0.0200312
R7148 VPWR.n3280 VPWR.n3279 0.0200312
R7149 VPWR.n3652 VPWR.n3651 0.0200312
R7150 VPWR.n3531 VPWR.n3530 0.0200312
R7151 VPWR.n1207 VPWR.n1206 0.0200312
R7152 VPWR.n1263 VPWR.n1234 0.0200312
R7153 VPWR.n3471 VPWR.n3470 0.0200312
R7154 VPWR.n3765 VPWR.n3764 0.0200312
R7155 VPWR.n3747 VPWR.n3746 0.0200312
R7156 VPWR.n1117 VPWR.n1116 0.0200312
R7157 VPWR.n982 VPWR.n981 0.0200312
R7158 VPWR.n3977 VPWR.n3976 0.0200312
R7159 VPWR.n987 VPWR.n986 0.0200312
R7160 VPWR.n3864 VPWR.n3863 0.0200312
R7161 VPWR.n3845 VPWR.n3844 0.0200312
R7162 VPWR.n4136 VPWR.n4135 0.0200312
R7163 VPWR.n810 VPWR.n809 0.0200312
R7164 VPWR.n835 VPWR.n834 0.0200312
R7165 VPWR.n951 VPWR.n950 0.0200312
R7166 VPWR.n4141 VPWR.n4140 0.0200312
R7167 VPWR.n4369 VPWR.n4368 0.0200312
R7168 VPWR.n851 VPWR.n850 0.0200312
R7169 VPWR.n4504 VPWR.n4503 0.0200312
R7170 VPWR.n4648 VPWR.n4647 0.0200312
R7171 VPWR.n4464 VPWR.n4463 0.0200312
R7172 VPWR.n4701 VPWR.n4700 0.0200312
R7173 VPWR.n4509 VPWR.n4508 0.0200312
R7174 VPWR.n4900 VPWR.n4899 0.0200312
R7175 VPWR.n4883 VPWR.n4882 0.0200312
R7176 VPWR.n250 VPWR.n249 0.0200312
R7177 VPWR.n649 VPWR.n644 0.0200312
R7178 VPWR.n5149 VPWR.n5148 0.0200312
R7179 VPWR.n255 VPWR.n254 0.0200312
R7180 VPWR.n5022 VPWR.n5021 0.0200312
R7181 VPWR.n5005 VPWR.n5004 0.0200312
R7182 VPWR.n5313 VPWR.n5312 0.0200312
R7183 VPWR.n487 VPWR.n486 0.0200312
R7184 VPWR.n508 VPWR.n507 0.0200312
R7185 VPWR.n619 VPWR.n618 0.0200312
R7186 VPWR.n347 VPWR 0.0200312
R7187 VPWR.n5318 VPWR.n5317 0.0200312
R7188 VPWR.n5798 VPWR.n5797 0.0200312
R7189 VPWR.n524 VPWR.n523 0.0200312
R7190 VPWR.n5422 VPWR.n153 0.0200312
R7191 VPWR.n5677 VPWR.n5676 0.0200312
R7192 VPWR.n6061 VPWR.n6060 0.0200312
R7193 VPWR.n5687 VPWR.n5686 0.0200312
R7194 VPWR.n5939 VPWR.n5938 0.0200312
R7195 VPWR.n5912 VPWR.n5911 0.0200312
R7196 VPWR.n6281 VPWR.n6280 0.0200312
R7197 VPWR.n6263 VPWR.n6262 0.0200312
R7198 VPWR.n2360 VPWR.n2359 0.0200312
R7199 VPWR.n2597 VPWR.n2596 0.0200312
R7200 VPWR.n2245 VPWR.n2244 0.0200312
R7201 VPWR.n2240 VPWR.n2239 0.0200312
R7202 VPWR.n5585 VPWR.n5584 0.0200312
R7203 VPWR.n145 VPWR.n144 0.0200312
R7204 VPWR.n5590 VPWR.n5589 0.0200312
R7205 VPWR.n141 VPWR.n140 0.0200312
R7206 VPWR.n3083 VPWR.n3082 0.0187292
R7207 VPWR.n3087 VPWR.n3086 0.0187292
R7208 VPWR.n1756 VPWR.n1752 0.0187292
R7209 VPWR.n2939 VPWR.n2937 0.0187292
R7210 VPWR.n3035 VPWR.n3034 0.0187292
R7211 VPWR.n1395 VPWR.n1318 0.0187292
R7212 VPWR.n3355 VPWR.n3354 0.0187292
R7213 VPWR.n3356 VPWR 0.0187292
R7214 VPWR.n3444 VPWR.n3443 0.0187292
R7215 VPWR.n3551 VPWR.n3550 0.0187292
R7216 VPWR.n1285 VPWR.n1281 0.0187292
R7217 VPWR.n1055 VPWR.n1051 0.0187292
R7218 VPWR.n4090 VPWR.n4089 0.0187292
R7219 VPWR.n4343 VPWR.n4342 0.0187292
R7220 VPWR.n4234 VPWR.n4232 0.0187292
R7221 VPWR.n4355 VPWR.n754 0.0187292
R7222 VPWR.n4810 VPWR.n4809 0.0187292
R7223 VPWR.n4711 VPWR.n4710 0.0187292
R7224 VPWR.n4823 VPWR.n4480 0.0187292
R7225 VPWR.n303 VPWR.n299 0.0187292
R7226 VPWR.n5159 VPWR.n5158 0.0187292
R7227 VPWR.n5275 VPWR.n5274 0.0187292
R7228 VPWR.n5779 VPWR.n5778 0.0187292
R7229 VPWR.n464 VPWR.n462 0.0187292
R7230 VPWR.n5783 VPWR.n5782 0.0187292
R7231 VPWR.n5391 VPWR.n5380 0.0187292
R7232 VPWR.n5456 VPWR.n5454 0.0187292
R7233 VPWR.n5557 VPWR.n5556 0.0187292
R7234 VPWR.n2109 VPWR.n2108 0.0187292
R7235 VPWR.n2334 VPWR.n2333 0.0187292
R7236 VPWR.n2330 VPWR.n2329 0.0187292
R7237 VPWR.n6184 VPWR.n6183 0.0187292
R7238 VPWR.n6082 VPWR.n6081 0.0187292
R7239 VPWR.n6180 VPWR.n6179 0.0187292
R7240 VPWR.n3404 VPWR.n1406 0.0179168
R7241 VPWR.n1291 VPWR.n1290 0.0179168
R7242 VPWR.n2052 VPWR.n2051 0.0174271
R7243 VPWR.n2103 VPWR.n2102 0.0174271
R7244 VPWR.n2106 VPWR.n2105 0.0174271
R7245 VPWR.n2388 VPWR.n2387 0.0174271
R7246 VPWR.n2380 VPWR.n2379 0.0174271
R7247 VPWR.n1585 VPWR.n1584 0.0174271
R7248 VPWR.n2622 VPWR.n2621 0.0174271
R7249 VPWR.n2743 VPWR.n2742 0.0174271
R7250 VPWR.n2740 VPWR.n2629 0.0174271
R7251 VPWR.n3112 VPWR.n3111 0.0174271
R7252 VPWR.n3109 VPWR.n3108 0.0174271
R7253 VPWR.n3097 VPWR.n1569 0.0174271
R7254 VPWR.n2632 VPWR.n2631 0.0174271
R7255 VPWR.n2739 VPWR.n2738 0.0174271
R7256 VPWR.n1591 VPWR.n1590 0.0174271
R7257 VPWR.n3099 VPWR.n1519 0.0174271
R7258 VPWR.n3105 VPWR.n3104 0.0174271
R7259 VPWR.n1667 VPWR.n1666 0.0174271
R7260 VPWR.n1784 VPWR.n1783 0.0174271
R7261 VPWR.n1793 VPWR.n1792 0.0174271
R7262 VPWR.n2934 VPWR.n2933 0.0174271
R7263 VPWR.n1893 VPWR.n1892 0.0174271
R7264 VPWR.n1906 VPWR.n1835 0.0174271
R7265 VPWR.n1911 VPWR.n1910 0.0174271
R7266 VPWR.n1786 VPWR.n1785 0.0174271
R7267 VPWR.n2937 VPWR.n2935 0.0174271
R7268 VPWR.n1673 VPWR.n1672 0.0174271
R7269 VPWR.n1897 VPWR.n1896 0.0174271
R7270 VPWR.n1903 VPWR.n1902 0.0174271
R7271 VPWR.n1455 VPWR.n1454 0.0174271
R7272 VPWR.n1460 VPWR.n1459 0.0174271
R7273 VPWR.n3352 VPWR.n3351 0.0174271
R7274 VPWR.n1322 VPWR.n1321 0.0174271
R7275 VPWR.n3214 VPWR.n3213 0.0174271
R7276 VPWR.n3211 VPWR.n3210 0.0174271
R7277 VPWR.n3293 VPWR.n3292 0.0174271
R7278 VPWR.n1418 VPWR.n1417 0.0174271
R7279 VPWR.n3354 VPWR.n3353 0.0174271
R7280 VPWR.n3201 VPWR.n3151 0.0174271
R7281 VPWR.n3207 VPWR.n3206 0.0174271
R7282 VPWR.n1240 VPWR.n1239 0.0174271
R7283 VPWR.n3634 VPWR.n3633 0.0174271
R7284 VPWR.n3631 VPWR.n1244 0.0174271
R7285 VPWR.n1297 VPWR.n1296 0.0174271
R7286 VPWR.n3775 VPWR.n3774 0.0174271
R7287 VPWR.n3772 VPWR.n3771 0.0174271
R7288 VPWR.n3760 VPWR.n3759 0.0174271
R7289 VPWR.n1248 VPWR.n1247 0.0174271
R7290 VPWR.n3630 VPWR.n3629 0.0174271
R7291 VPWR.n3762 VPWR.n1139 0.0174271
R7292 VPWR.n3768 VPWR.n3767 0.0174271
R7293 VPWR.n1094 VPWR.n1093 0.0174271
R7294 VPWR.n1099 VPWR.n1098 0.0174271
R7295 VPWR.n3986 VPWR.n3985 0.0174271
R7296 VPWR.n968 VPWR.n967 0.0174271
R7297 VPWR.n3874 VPWR.n3873 0.0174271
R7298 VPWR.n3871 VPWR.n3870 0.0174271
R7299 VPWR.n3859 VPWR.n3856 0.0174271
R7300 VPWR.n3836 VPWR 0.0174271
R7301 VPWR.n1072 VPWR.n1071 0.0174271
R7302 VPWR.n3988 VPWR.n3987 0.0174271
R7303 VPWR.n974 VPWR.n973 0.0174271
R7304 VPWR.n3861 VPWR.n3804 0.0174271
R7305 VPWR.n3867 VPWR.n3866 0.0174271
R7306 VPWR.n4122 VPWR.n4121 0.0174271
R7307 VPWR.n787 VPWR.n786 0.0174271
R7308 VPWR.n792 VPWR.n791 0.0174271
R7309 VPWR.n4229 VPWR.n4228 0.0174271
R7310 VPWR.n4379 VPWR.n4378 0.0174271
R7311 VPWR.n4376 VPWR.n4375 0.0174271
R7312 VPWR.n4364 VPWR.n749 0.0174271
R7313 VPWR.n774 VPWR.n773 0.0174271
R7314 VPWR.n4232 VPWR.n4230 0.0174271
R7315 VPWR.n4353 VPWR.n4352 0.0174271
R7316 VPWR.n4128 VPWR.n4127 0.0174271
R7317 VPWR.n4366 VPWR.n700 0.0174271
R7318 VPWR.n4372 VPWR.n4371 0.0174271
R7319 VPWR.n4490 VPWR.n4489 0.0174271
R7320 VPWR.n4625 VPWR.n4624 0.0174271
R7321 VPWR.n4630 VPWR.n4629 0.0174271
R7322 VPWR.n4708 VPWR.n4707 0.0174271
R7323 VPWR.n4910 VPWR.n4909 0.0174271
R7324 VPWR.n4907 VPWR.n4906 0.0174271
R7325 VPWR.n4895 VPWR.n4894 0.0174271
R7326 VPWR.n4602 VPWR.n4601 0.0174271
R7327 VPWR.n4710 VPWR.n4709 0.0174271
R7328 VPWR.n4821 VPWR.n4820 0.0174271
R7329 VPWR.n4496 VPWR.n4495 0.0174271
R7330 VPWR.n4897 VPWR.n4398 0.0174271
R7331 VPWR.n4903 VPWR.n4902 0.0174271
R7332 VPWR.n236 VPWR.n235 0.0174271
R7333 VPWR.n655 VPWR.n654 0.0174271
R7334 VPWR.n668 VPWR.n667 0.0174271
R7335 VPWR.n5156 VPWR.n5155 0.0174271
R7336 VPWR.n5032 VPWR.n5031 0.0174271
R7337 VPWR.n5029 VPWR.n5028 0.0174271
R7338 VPWR.n5017 VPWR.n5016 0.0174271
R7339 VPWR.n676 VPWR.n675 0.0174271
R7340 VPWR.n5158 VPWR.n5157 0.0174271
R7341 VPWR.n242 VPWR.n241 0.0174271
R7342 VPWR.n5019 VPWR.n4938 0.0174271
R7343 VPWR.n5025 VPWR.n5024 0.0174271
R7344 VPWR.n5299 VPWR.n5298 0.0174271
R7345 VPWR.n338 VPWR.n337 0.0174271
R7346 VPWR.n469 VPWR.n468 0.0174271
R7347 VPWR.n466 VPWR.n344 0.0174271
R7348 VPWR.n5808 VPWR.n5807 0.0174271
R7349 VPWR.n5805 VPWR.n5804 0.0174271
R7350 VPWR.n5793 VPWR.n223 0.0174271
R7351 VPWR.n348 VPWR.n347 0.0174271
R7352 VPWR.n465 VPWR.n464 0.0174271
R7353 VPWR.n5305 VPWR.n5304 0.0174271
R7354 VPWR.n5795 VPWR.n183 0.0174271
R7355 VPWR.n5801 VPWR.n5800 0.0174271
R7356 VPWR.n5429 VPWR.n5428 0.0174271
R7357 VPWR.n5442 VPWR.n5441 0.0174271
R7358 VPWR.n5451 VPWR.n5450 0.0174271
R7359 VPWR.n5675 VPWR.n5674 0.0174271
R7360 VPWR.n5949 VPWR.n5948 0.0174271
R7361 VPWR.n5946 VPWR.n5945 0.0174271
R7362 VPWR.n5934 VPWR.n5923 0.0174271
R7363 VPWR.n5903 VPWR 0.0174271
R7364 VPWR.n5414 VPWR.n5413 0.0174271
R7365 VPWR.n5454 VPWR.n5452 0.0174271
R7366 VPWR.n5401 VPWR.n5400 0.0174271
R7367 VPWR.n5672 VPWR.n5671 0.0174271
R7368 VPWR.n5936 VPWR.n5856 0.0174271
R7369 VPWR.n5942 VPWR.n5941 0.0174271
R7370 VPWR.n6284 VPWR.n6283 0.0174271
R7371 VPWR.n34 VPWR.n33 0.0174271
R7372 VPWR.n2460 VPWR.n2459 0.0174271
R7373 VPWR.n2457 VPWR.n2456 0.0174271
R7374 VPWR.n2454 VPWR.n2447 0.0174271
R7375 VPWR.n2061 VPWR.n2060 0.0174271
R7376 VPWR.n2089 VPWR.n2088 0.0174271
R7377 VPWR.n2108 VPWR.n2107 0.0174271
R7378 VPWR.n2232 VPWR.n2231 0.0174271
R7379 VPWR.n2226 VPWR.n2225 0.0174271
R7380 VPWR.n5571 VPWR.n5570 0.0174271
R7381 VPWR.n29 VPWR.n28 0.0174271
R7382 VPWR.n6277 VPWR.n31 0.0174271
R7383 VPWR.n6275 VPWR.n6274 0.0174271
R7384 VPWR.n55 VPWR 0.0174271
R7385 VPWR.n99 VPWR.n98 0.0174271
R7386 VPWR.n6081 VPWR.n6080 0.0174271
R7387 VPWR.n5577 VPWR.n5576 0.0174271
R7388 VPWR.n118 VPWR.n117 0.0174271
R7389 VPWR.n123 VPWR.n122 0.0174271
R7390 VPWR.n6079 VPWR.n6078 0.0174271
R7391 VPWR.n4116 VPWR.n4115 0.0173639
R7392 VPWR.n4224 VPWR.n778 0.0173639
R7393 VPWR.n689 VPWR.n688 0.0173639
R7394 VPWR.n3839 VPWR.n3837 0.0172647
R7395 VPWR.n4999 VPWR.n4996 0.0172647
R7396 VPWR.n506 VPWR.n505 0.0172647
R7397 VPWR.n57 VPWR.n56 0.0172647
R7398 VPWR.n2043 VPWR.n2041 0.0168788
R7399 VPWR.n2606 VPWR.n2605 0.0168788
R7400 VPWR.n3065 VPWR.n3060 0.0168788
R7401 VPWR.n2918 VPWR.n2915 0.0168788
R7402 VPWR.n2613 VPWR.n2612 0.0168788
R7403 VPWR.n3124 VPWR.n3119 0.0168788
R7404 VPWR.n3048 VPWR.n3046 0.0168788
R7405 VPWR.n3054 VPWR.n3053 0.0168788
R7406 VPWR.n1780 VPWR.n1778 0.0168788
R7407 VPWR.n2926 VPWR.n2925 0.0168788
R7408 VPWR.n3134 VPWR.n3131 0.0168788
R7409 VPWR.n1449 VPWR.n1444 0.0168788
R7410 VPWR.n3454 VPWR.n3451 0.0168788
R7411 VPWR.n1314 VPWR.n1313 0.0168788
R7412 VPWR.n3147 VPWR.n3142 0.0168788
R7413 VPWR.n1432 VPWR.n1427 0.0168788
R7414 VPWR.n1306 VPWR.n1303 0.0168788
R7415 VPWR.n3461 VPWR.n3460 0.0168788
R7416 VPWR.n3787 VPWR.n3782 0.0168788
R7417 VPWR.n1088 VPWR.n1083 0.0168788
R7418 VPWR.n4100 VPWR.n4097 0.0168788
R7419 VPWR.n1047 VPWR.n1046 0.0168788
R7420 VPWR.n3800 VPWR.n3795 0.0168788
R7421 VPWR.n4119 VPWR.n4117 0.0168788
R7422 VPWR.n4109 VPWR.n4108 0.0168788
R7423 VPWR.n783 VPWR.n780 0.0168788
R7424 VPWR.n4222 VPWR.n4221 0.0168788
R7425 VPWR.n698 VPWR.n695 0.0168788
R7426 VPWR.n693 VPWR.n692 0.0168788
R7427 VPWR.n4574 VPWR.n4569 0.0168788
R7428 VPWR.n4613 VPWR.n4610 0.0168788
R7429 VPWR.n4619 VPWR.n4618 0.0168788
R7430 VPWR.n4922 VPWR.n4917 0.0168788
R7431 VPWR.n5289 VPWR.n5284 0.0168788
R7432 VPWR.n635 VPWR.n632 0.0168788
R7433 VPWR.n640 VPWR.n639 0.0168788
R7434 VPWR.n4934 VPWR.n4929 0.0168788
R7435 VPWR.n5761 VPWR.n5756 0.0168788
R7436 VPWR.n329 VPWR.n326 0.0168788
R7437 VPWR.n627 VPWR.n626 0.0168788
R7438 VPWR.n5820 VPWR.n5815 0.0168788
R7439 VPWR.n6071 VPWR.n6067 0.0168788
R7440 VPWR.n5445 VPWR.n5444 0.0168788
R7441 VPWR.n5660 VPWR.n5658 0.0168788
R7442 VPWR.n5749 VPWR.n5748 0.0168788
R7443 VPWR.n5852 VPWR.n5847 0.0168788
R7444 VPWR.n5837 VPWR.n5836 0.0168788
R7445 VPWR.n5832 VPWR.n5831 0.0168788
R7446 VPWR.n2474 VPWR.n2469 0.0168788
R7447 VPWR.n2220 VPWR.n2219 0.0168788
R7448 VPWR.n5653 VPWR.n5648 0.0168788
R7449 VPWR.n112 VPWR.n108 0.0168788
R7450 VPWR.n103 VPWR.n102 0.0168788
R7451 VPWR.n3840 VPWR.n3839 0.0166259
R7452 VPWR.n5000 VPWR.n4999 0.0166259
R7453 VPWR.n505 VPWR.n504 0.0166259
R7454 VPWR.n57 VPWR.n32 0.0166259
R7455 VPWR.n1565 VPWR.n1564 0.016125
R7456 VPWR.n2907 VPWR.n2764 0.016125
R7457 VPWR.n1887 VPWR.n1886 0.016125
R7458 VPWR.n3197 VPWR.n3196 0.016125
R7459 VPWR.n1389 VPWR 0.016125
R7460 VPWR.n1186 VPWR.n1185 0.016125
R7461 VPWR.n3539 VPWR 0.016125
R7462 VPWR.n745 VPWR.n744 0.016125
R7463 VPWR.n4443 VPWR.n4442 0.016125
R7464 VPWR.n4699 VPWR.n4650 0.016125
R7465 VPWR.n4990 VPWR.n4989 0.016125
R7466 VPWR.n6059 VPWR.n154 0.016125
R7467 VPWR.n2442 VPWR.n2441 0.016125
R7468 VPWR.n2595 VPWR.n2064 0.016125
R7469 VPWR.n1787 VPWR 0.0158144
R7470 VPWR.n3792 VPWR.n3791 0.0153171
R7471 VPWR.n4104 VPWR.n4103 0.0153171
R7472 VPWR.n1080 VPWR.n1079 0.0153171
R7473 VPWR.n2738 VPWR.n2737 0.0149528
R7474 VPWR.n2599 VPWR.n2058 0.0148229
R7475 VPWR.n2106 VPWR.n2104 0.0148229
R7476 VPWR.n2462 VPWR.n2388 0.0148229
R7477 VPWR.n3084 VPWR.n3083 0.0148229
R7478 VPWR.n2911 VPWR.n2761 0.0148229
R7479 VPWR.n2741 VPWR.n2740 0.0148229
R7480 VPWR.n2910 VPWR.n2909 0.0148229
R7481 VPWR.n2739 VPWR.n2633 0.0148229
R7482 VPWR.n3086 VPWR.n3085 0.0148229
R7483 VPWR.n3114 VPWR.n1519 0.0148229
R7484 VPWR.n3037 VPWR.n1752 0.0148229
R7485 VPWR.n2034 VPWR.n1811 0.0148229
R7486 VPWR.n2934 VPWR.n1775 0.0148229
R7487 VPWR.n2033 VPWR.n2032 0.0148229
R7488 VPWR.n2935 VPWR.n1774 0.0148229
R7489 VPWR.n3036 VPWR.n3035 0.0148229
R7490 VPWR.n1896 VPWR.n1895 0.0148229
R7491 VPWR.n3345 VPWR.n1478 0.0148229
R7492 VPWR.n3352 VPWR.n1420 0.0148229
R7493 VPWR.n3446 VPWR.n1318 0.0148229
R7494 VPWR.n3344 VPWR.n3343 0.0148229
R7495 VPWR.n3353 VPWR.n1419 0.0148229
R7496 VPWR.n3445 VPWR.n3444 0.0148229
R7497 VPWR.n1393 VPWR.n1392 0.0148229
R7498 VPWR.n3216 VPWR.n3151 0.0148229
R7499 VPWR.n3653 VPWR.n3652 0.0148229
R7500 VPWR.n3632 VPWR.n3631 0.0148229
R7501 VPWR.n3552 VPWR.n3551 0.0148229
R7502 VPWR.n3654 VPWR.n1234 0.0148229
R7503 VPWR.n3630 VPWR.n1249 0.0148229
R7504 VPWR.n3553 VPWR.n1281 0.0148229
R7505 VPWR.n3543 VPWR.n3542 0.0148229
R7506 VPWR.n3777 VPWR.n1139 0.0148229
R7507 VPWR.n3979 VPWR.n1117 0.0148229
R7508 VPWR.n3986 VPWR.n1074 0.0148229
R7509 VPWR.n4092 VPWR.n1051 0.0148229
R7510 VPWR.n3978 VPWR.n3977 0.0148229
R7511 VPWR.n3987 VPWR.n1073 0.0148229
R7512 VPWR.n4091 VPWR.n4090 0.0148229
R7513 VPWR.n3876 VPWR.n3804 0.0148229
R7514 VPWR.n4342 VPWR.n4341 0.0148229
R7515 VPWR.n953 VPWR.n810 0.0148229
R7516 VPWR.n4229 VPWR.n776 0.0148229
R7517 VPWR.n952 VPWR.n951 0.0148229
R7518 VPWR.n4230 VPWR.n775 0.0148229
R7519 VPWR.n4340 VPWR.n754 0.0148229
R7520 VPWR.n4352 VPWR 0.0148229
R7521 VPWR.n4381 VPWR.n700 0.0148229
R7522 VPWR.n4809 VPWR.n4808 0.0148229
R7523 VPWR.n4703 VPWR.n4648 0.0148229
R7524 VPWR.n4708 VPWR.n4604 0.0148229
R7525 VPWR.n4702 VPWR.n4701 0.0148229
R7526 VPWR.n4709 VPWR.n4603 0.0148229
R7527 VPWR.n4807 VPWR.n4480 0.0148229
R7528 VPWR.n4820 VPWR 0.0148229
R7529 VPWR.n4912 VPWR.n4398 0.0148229
R7530 VPWR.n5277 VPWR.n299 0.0148229
R7531 VPWR.n5151 VPWR.n644 0.0148229
R7532 VPWR.n5156 VPWR.n319 0.0148229
R7533 VPWR.n5150 VPWR.n5149 0.0148229
R7534 VPWR.n5157 VPWR.n318 0.0148229
R7535 VPWR.n5276 VPWR.n5275 0.0148229
R7536 VPWR.n5034 VPWR.n4938 0.0148229
R7537 VPWR.n5780 VPWR.n5779 0.0148229
R7538 VPWR.n621 VPWR.n487 0.0148229
R7539 VPWR.n467 VPWR.n466 0.0148229
R7540 VPWR.n620 VPWR.n619 0.0148229
R7541 VPWR.n465 VPWR.n349 0.0148229
R7542 VPWR.n5782 VPWR.n5781 0.0148229
R7543 VPWR.n5810 VPWR.n183 0.0148229
R7544 VPWR.n6063 VPWR.n153 0.0148229
R7545 VPWR.n5451 VPWR.n5443 0.0148229
R7546 VPWR.n5559 VPWR.n5380 0.0148229
R7547 VPWR.n6062 VPWR.n6061 0.0148229
R7548 VPWR.n5452 VPWR.n5415 0.0148229
R7549 VPWR.n5558 VPWR.n5557 0.0148229
R7550 VPWR.n5400 VPWR 0.0148229
R7551 VPWR.n5951 VPWR.n5856 0.0148229
R7552 VPWR.n6285 VPWR.n6284 0.0148229
R7553 VPWR.n2461 VPWR.n2460 0.0148229
R7554 VPWR.n2598 VPWR 0.0148229
R7555 VPWR.n2598 VPWR.n2597 0.0148229
R7556 VPWR.n2107 VPWR.n2090 0.0148229
R7557 VPWR.n2333 VPWR.n2332 0.0148229
R7558 VPWR.n2331 VPWR.n2330 0.0148229
R7559 VPWR.n6183 VPWR.n6182 0.0148229
R7560 VPWR.n146 VPWR 0.0148229
R7561 VPWR.n146 VPWR.n145 0.0148229
R7562 VPWR.n6080 VPWR.n100 0.0148229
R7563 VPWR.n6181 VPWR.n6180 0.0148229
R7564 VPWR.n5573 VPWR.n5572 0.0148229
R7565 VPWR.n147 VPWR.n141 0.0148229
R7566 VPWR.n6079 VPWR.n101 0.0148229
R7567 VPWR.n3032 VPWR 0.0146642
R7568 VPWR.n5785 VPWR 0.0146642
R7569 VPWR.n4087 VPWR 0.0146642
R7570 VPWR.n5710 VPWR.n5691 0.0138584
R7571 VPWR.n2051 VPWR.n2050 0.0135208
R7572 VPWR.n2381 VPWR.n2380 0.0135208
R7573 VPWR.n1584 VPWR.n1583 0.0135208
R7574 VPWR.n1600 VPWR.n1599 0.0135208
R7575 VPWR.n2621 VPWR.n2620 0.0135208
R7576 VPWR.n3113 VPWR 0.0135208
R7577 VPWR.n3098 VPWR.n3097 0.0135208
R7578 VPWR.n2753 VPWR.n2752 0.0135208
R7579 VPWR.n1610 VPWR.n1604 0.0135208
R7580 VPWR.n3106 VPWR.n3105 0.0135208
R7581 VPWR.n1666 VPWR.n1665 0.0135208
R7582 VPWR.n1682 VPWR.n1681 0.0135208
R7583 VPWR.n1783 VPWR.n1782 0.0135208
R7584 VPWR.n1894 VPWR 0.0135208
R7585 VPWR.n1910 VPWR.n1907 0.0135208
R7586 VPWR.n1803 VPWR.n1802 0.0135208
R7587 VPWR.n1692 VPWR.n1686 0.0135208
R7588 VPWR.n1904 VPWR.n1903 0.0135208
R7589 VPWR.n1454 VPWR.n1453 0.0135208
R7590 VPWR.n1321 VPWR.n1320 0.0135208
R7591 VPWR.n1380 VPWR.n1379 0.0135208
R7592 VPWR.n3215 VPWR 0.0135208
R7593 VPWR.n3293 VPWR.n1496 0.0135208
R7594 VPWR.n1470 VPWR.n1469 0.0135208
R7595 VPWR.n1330 VPWR.n1326 0.0135208
R7596 VPWR.n3208 VPWR.n3207 0.0135208
R7597 VPWR.n1239 VPWR.n1238 0.0135208
R7598 VPWR.n1296 VPWR.n1295 0.0135208
R7599 VPWR.n3530 VPWR.n3529 0.0135208
R7600 VPWR.n3776 VPWR 0.0135208
R7601 VPWR.n3761 VPWR.n3760 0.0135208
R7602 VPWR.n3644 VPWR.n3643 0.0135208
R7603 VPWR.n3474 VPWR.n3471 0.0135208
R7604 VPWR.n3769 VPWR.n3768 0.0135208
R7605 VPWR.n1093 VPWR.n1092 0.0135208
R7606 VPWR.n967 VPWR.n966 0.0135208
R7607 VPWR.n983 VPWR.n982 0.0135208
R7608 VPWR.n3875 VPWR 0.0135208
R7609 VPWR.n3860 VPWR.n3859 0.0135208
R7610 VPWR.n1109 VPWR.n1108 0.0135208
R7611 VPWR.n993 VPWR.n987 0.0135208
R7612 VPWR.n3868 VPWR.n3867 0.0135208
R7613 VPWR.n4121 VPWR.n4120 0.0135208
R7614 VPWR.n4137 VPWR.n4136 0.0135208
R7615 VPWR.n786 VPWR.n785 0.0135208
R7616 VPWR.n4380 VPWR 0.0135208
R7617 VPWR.n4365 VPWR.n4364 0.0135208
R7618 VPWR.n802 VPWR.n801 0.0135208
R7619 VPWR.n4147 VPWR.n4141 0.0135208
R7620 VPWR.n4373 VPWR.n4372 0.0135208
R7621 VPWR.n4489 VPWR.n4488 0.0135208
R7622 VPWR.n4505 VPWR.n4504 0.0135208
R7623 VPWR.n4624 VPWR.n4623 0.0135208
R7624 VPWR.n4911 VPWR 0.0135208
R7625 VPWR.n4896 VPWR.n4895 0.0135208
R7626 VPWR.n4640 VPWR.n4639 0.0135208
R7627 VPWR.n4515 VPWR.n4509 0.0135208
R7628 VPWR.n4904 VPWR.n4903 0.0135208
R7629 VPWR.n235 VPWR.n234 0.0135208
R7630 VPWR.n251 VPWR.n250 0.0135208
R7631 VPWR.n654 VPWR.n653 0.0135208
R7632 VPWR.n5033 VPWR 0.0135208
R7633 VPWR.n5018 VPWR.n5017 0.0135208
R7634 VPWR.n660 VPWR.n659 0.0135208
R7635 VPWR.n260 VPWR.n255 0.0135208
R7636 VPWR.n5026 VPWR.n5025 0.0135208
R7637 VPWR.n5298 VPWR.n5297 0.0135208
R7638 VPWR.n5314 VPWR.n5313 0.0135208
R7639 VPWR.n337 VPWR.n336 0.0135208
R7640 VPWR.n5809 VPWR 0.0135208
R7641 VPWR.n5794 VPWR.n5793 0.0135208
R7642 VPWR.n479 VPWR.n478 0.0135208
R7643 VPWR.n5324 VPWR.n5318 0.0135208
R7644 VPWR.n5802 VPWR.n5801 0.0135208
R7645 VPWR.n5428 VPWR.n5427 0.0135208
R7646 VPWR.n5674 VPWR.n5673 0.0135208
R7647 VPWR.n5676 VPWR.n5664 0.0135208
R7648 VPWR.n5950 VPWR 0.0135208
R7649 VPWR.n5935 VPWR.n5934 0.0135208
R7650 VPWR.n5421 VPWR.n5420 0.0135208
R7651 VPWR.n5432 VPWR.n5431 0.0135208
R7652 VPWR.n5689 VPWR.n5687 0.0135208
R7653 VPWR.n5943 VPWR.n5942 0.0135208
R7654 VPWR.n33 VPWR.n27 0.0135208
R7655 VPWR.n2455 VPWR.n2454 0.0135208
R7656 VPWR.n2063 VPWR.n2062 0.0135208
R7657 VPWR.n2060 VPWR.n2059 0.0135208
R7658 VPWR.n2251 VPWR.n2245 0.0135208
R7659 VPWR.n2225 VPWR.n2224 0.0135208
R7660 VPWR.n2241 VPWR.n2240 0.0135208
R7661 VPWR.n5570 VPWR.n5569 0.0135208
R7662 VPWR.n5586 VPWR.n5585 0.0135208
R7663 VPWR.n6286 VPWR 0.0135208
R7664 VPWR.n6276 VPWR.n6275 0.0135208
R7665 VPWR.n133 VPWR.n132 0.0135208
R7666 VPWR.n5591 VPWR.n5590 0.0135208
R7667 VPWR.n117 VPWR.n116 0.0135208
R7668 VPWR.n3089 VPWR.n3088 0.0133621
R7669 VPWR.n3033 VPWR.n3032 0.0133621
R7670 VPWR.n5273 VPWR.n5272 0.0133621
R7671 VPWR.n5785 VPWR.n5784 0.0133621
R7672 VPWR.n2336 VPWR.n2335 0.0133621
R7673 VPWR.n3442 VPWR.n3441 0.0133621
R7674 VPWR.n1294 VPWR.n1286 0.0133621
R7675 VPWR.n4088 VPWR.n4087 0.0133621
R7676 VPWR.n6191 VPWR.n79 0.0133621
R7677 VPWR.n2041 VPWR.n2040 0.0130912
R7678 VPWR.n2605 VPWR.n2604 0.0130912
R7679 VPWR.n3060 VPWR.n3059 0.0130912
R7680 VPWR.n1580 VPWR.n1579 0.0130912
R7681 VPWR.n2915 VPWR.n2914 0.0130912
R7682 VPWR.n2612 VPWR.n2611 0.0130912
R7683 VPWR.n3119 VPWR.n3118 0.0130912
R7684 VPWR.n2803 VPWR.n2802 0.0130912
R7685 VPWR.n1444 VPWR.n1443 0.0130912
R7686 VPWR.n1422 VPWR.n1421 0.0130912
R7687 VPWR.n3451 VPWR.n3450 0.0130912
R7688 VPWR.n1313 VPWR.n1312 0.0130912
R7689 VPWR.n3142 VPWR.n3141 0.0130912
R7690 VPWR.n1501 VPWR.n1500 0.0130912
R7691 VPWR.n1427 VPWR.n1426 0.0130912
R7692 VPWR.n1436 VPWR.n1435 0.0130912
R7693 VPWR.n1303 VPWR.n1302 0.0130912
R7694 VPWR.n3460 VPWR.n3459 0.0130912
R7695 VPWR.n3782 VPWR.n3781 0.0130912
R7696 VPWR.n1195 VPWR.n1194 0.0130912
R7697 VPWR.n1083 VPWR.n1082 0.0130912
R7698 VPWR.n1076 VPWR.n1075 0.0130912
R7699 VPWR.n4097 VPWR.n4096 0.0130912
R7700 VPWR.n1046 VPWR.n1045 0.0130912
R7701 VPWR.n3795 VPWR.n3794 0.0130912
R7702 VPWR.n1134 VPWR.n1133 0.0130912
R7703 VPWR.n4108 VPWR.n4107 0.0130912
R7704 VPWR.n780 VPWR.n779 0.0130912
R7705 VPWR.n695 VPWR.n694 0.0130912
R7706 VPWR.n4569 VPWR.n4568 0.0130912
R7707 VPWR.n4485 VPWR.n4484 0.0130912
R7708 VPWR.n4610 VPWR.n4609 0.0130912
R7709 VPWR.n4618 VPWR.n4617 0.0130912
R7710 VPWR.n4917 VPWR.n4916 0.0130912
R7711 VPWR.n4452 VPWR.n4451 0.0130912
R7712 VPWR.n5284 VPWR.n5283 0.0130912
R7713 VPWR.n231 VPWR.n230 0.0130912
R7714 VPWR.n632 VPWR.n631 0.0130912
R7715 VPWR.n639 VPWR.n638 0.0130912
R7716 VPWR.n4929 VPWR.n4928 0.0130912
R7717 VPWR.n686 VPWR.n685 0.0130912
R7718 VPWR.n5756 VPWR.n5755 0.0130912
R7719 VPWR.n5294 VPWR.n5293 0.0130912
R7720 VPWR.n326 VPWR.n325 0.0130912
R7721 VPWR.n626 VPWR.n625 0.0130912
R7722 VPWR.n5815 VPWR.n5814 0.0130912
R7723 VPWR.n527 VPWR.n526 0.0130912
R7724 VPWR.n6067 VPWR.n6066 0.0130912
R7725 VPWR.n5446 VPWR.n5445 0.0130912
R7726 VPWR.n5658 VPWR.n5657 0.0130912
R7727 VPWR.n5748 VPWR.n5747 0.0130912
R7728 VPWR.n5847 VPWR.n5846 0.0130912
R7729 VPWR.n177 VPWR.n176 0.0130912
R7730 VPWR.n5838 VPWR.n5837 0.0130912
R7731 VPWR.n5831 VPWR.n5830 0.0130912
R7732 VPWR.n2374 VPWR.n2373 0.0130912
R7733 VPWR.n2315 VPWR.n2314 0.0130912
R7734 VPWR.n2219 VPWR.n2218 0.0130912
R7735 VPWR.n5648 VPWR.n5647 0.0130912
R7736 VPWR.n5565 VPWR.n5564 0.0130912
R7737 VPWR.n108 VPWR.n107 0.0130912
R7738 VPWR.n104 VPWR.n103 0.0130912
R7739 VPWR.n2372 VPWR.n2371 0.0122188
R7740 VPWR.n2787 VPWR.n2786 0.0122188
R7741 VPWR.n2790 VPWR.n2789 0.0122188
R7742 VPWR.n2801 VPWR.n2800 0.0122188
R7743 VPWR.n1828 VPWR.n1827 0.0122188
R7744 VPWR.n1831 VPWR.n1830 0.0122188
R7745 VPWR.n1925 VPWR.n1924 0.0122188
R7746 VPWR.n3229 VPWR.n3228 0.0122188
R7747 VPWR.n3232 VPWR.n3231 0.0122188
R7748 VPWR.n3279 VPWR.n3278 0.0122188
R7749 VPWR.n1205 VPWR.n1204 0.0122188
R7750 VPWR.n1208 VPWR.n1207 0.0122188
R7751 VPWR.n3746 VPWR.n3745 0.0122188
R7752 VPWR.n3835 VPWR.n1131 0.0122188
R7753 VPWR.n3844 VPWR.n1132 0.0122188
R7754 VPWR.n833 VPWR.n832 0.0122188
R7755 VPWR.n836 VPWR.n835 0.0122188
R7756 VPWR.n852 VPWR.n851 0.0122188
R7757 VPWR.n4462 VPWR.n4461 0.0122188
R7758 VPWR.n4465 VPWR.n4464 0.0122188
R7759 VPWR.n4882 VPWR.n4881 0.0122188
R7760 VPWR VPWR.n4994 0.0122188
R7761 VPWR.n4994 VPWR.n683 0.0122188
R7762 VPWR.n5004 VPWR.n684 0.0122188
R7763 VPWR.n509 VPWR.n508 0.0122188
R7764 VPWR.n525 VPWR.n524 0.0122188
R7765 VPWR.n5905 VPWR.n5904 0.0122188
R7766 VPWR.n5902 VPWR.n174 0.0122188
R7767 VPWR.n5911 VPWR.n175 0.0122188
R7768 VPWR.n6262 VPWR.n6261 0.0122188
R7769 VPWR.n2358 VPWR.n2357 0.0122188
R7770 VPWR.n2361 VPWR.n2360 0.0122188
R7771 VPWR.n54 VPWR.n38 0.0122188
R7772 VPWR.n218 VPWR.n217 0.0117355
R7773 VPWR.n5147 VPWR.n645 0.011097
R7774 VPWR.n617 VPWR.n616 0.011097
R7775 VPWR.n1264 VPWR.n1262 0.011097
R7776 VPWR.n3975 VPWR.n1118 0.011097
R7777 VPWR.n949 VPWR.n948 0.011097
R7778 VPWR.n6288 VPWR.n6287 0.011097
R7779 VPWR.n2384 VPWR.n2383 0.0109167
R7780 VPWR.n2785 VPWR.n2784 0.0109167
R7781 VPWR.n3103 VPWR.n3102 0.0109167
R7782 VPWR.n1825 VPWR.n1823 0.0109167
R7783 VPWR.n1901 VPWR.n1900 0.0109167
R7784 VPWR.n3226 VPWR.n3224 0.0109167
R7785 VPWR.n3205 VPWR.n3204 0.0109167
R7786 VPWR.n1202 VPWR.n1200 0.0109167
R7787 VPWR VPWR 0.0109167
R7788 VPWR VPWR 0.0109167
R7789 VPWR.n3766 VPWR.n3765 0.0109167
R7790 VPWR.n3865 VPWR.n3864 0.0109167
R7791 VPWR.n830 VPWR.n828 0.0109167
R7792 VPWR.n4370 VPWR.n4369 0.0109167
R7793 VPWR.n4459 VPWR.n4457 0.0109167
R7794 VPWR VPWR 0.0109167
R7795 VPWR.n4901 VPWR.n4900 0.0109167
R7796 VPWR VPWR 0.0109167
R7797 VPWR.n5023 VPWR.n5022 0.0109167
R7798 VPWR.n5799 VPWR.n5798 0.0109167
R7799 VPWR.n5907 VPWR.n5906 0.0109167
R7800 VPWR VPWR 0.0109167
R7801 VPWR.n5940 VPWR.n5939 0.0109167
R7802 VPWR.n6280 VPWR.n6279 0.0109167
R7803 VPWR.n2356 VPWR.n2355 0.0109167
R7804 VPWR VPWR 0.0109167
R7805 VPWR.n5575 VPWR.n5574 0.0108178
R7806 VPWR.n2030 VPWR.n2029 0.0107609
R7807 VPWR.n3341 VPWR.n1479 0.0107609
R7808 VPWR.n143 VPWR.n142 0.0107609
R7809 VPWR.n3128 VPWR.n3127 0.0100114
R7810 VPWR.n3057 VPWR.n3056 0.0100114
R7811 VPWR.n2922 VPWR.n2921 0.0100114
R7812 VPWR.n2049 VPWR.n2048 0.00975758
R7813 VPWR.n2046 VPWR.n2045 0.00975758
R7814 VPWR.n3070 VPWR.n3069 0.00975758
R7815 VPWR.n1582 VPWR.n1581 0.00975758
R7816 VPWR.n2619 VPWR.n2618 0.00975758
R7817 VPWR.n2616 VPWR.n2615 0.00975758
R7818 VPWR.n1518 VPWR.n1517 0.00975758
R7819 VPWR.n2805 VPWR.n2804 0.00975758
R7820 VPWR.n3041 VPWR.n3040 0.00975758
R7821 VPWR.n1750 VPWR.n1749 0.00975758
R7822 VPWR.n2037 VPWR.n2036 0.00975758
R7823 VPWR.n2931 VPWR.n2930 0.00975758
R7824 VPWR.n1837 VPWR.n1836 0.00975758
R7825 VPWR.n1927 VPWR.n1926 0.00975758
R7826 VPWR.n1452 VPWR.n1451 0.00975758
R7827 VPWR.n3349 VPWR.n1423 0.00975758
R7828 VPWR.n1317 VPWR.n1316 0.00975758
R7829 VPWR.n1309 VPWR.n1308 0.00975758
R7830 VPWR.n3150 VPWR.n3149 0.00975758
R7831 VPWR.n3221 VPWR.n1502 0.00975758
R7832 VPWR.n1236 VPWR.n1235 0.00975758
R7833 VPWR.n1439 VPWR.n1437 0.00975758
R7834 VPWR.n3464 VPWR.n3463 0.00975758
R7835 VPWR.n1299 VPWR.n1298 0.00975758
R7836 VPWR.n1138 VPWR.n1137 0.00975758
R7837 VPWR.n1197 VPWR.n1196 0.00975758
R7838 VPWR.n1091 VPWR.n1090 0.00975758
R7839 VPWR.n3983 VPWR.n1077 0.00975758
R7840 VPWR.n1050 VPWR.n1049 0.00975758
R7841 VPWR.n965 VPWR.n964 0.00975758
R7842 VPWR.n3803 VPWR.n3802 0.00975758
R7843 VPWR.n3881 VPWR.n1135 0.00975758
R7844 VPWR.n4114 VPWR.n4113 0.00975758
R7845 VPWR.n4205 VPWR.n4204 0.00975758
R7846 VPWR.n956 VPWR.n955 0.00975758
R7847 VPWR.n4226 VPWR.n4225 0.00975758
R7848 VPWR.n4385 VPWR.n4384 0.00975758
R7849 VPWR.n855 VPWR.n854 0.00975758
R7850 VPWR.n4579 VPWR.n4578 0.00975758
R7851 VPWR.n4487 VPWR.n4486 0.00975758
R7852 VPWR.n4622 VPWR.n4621 0.00975758
R7853 VPWR.n4606 VPWR.n4605 0.00975758
R7854 VPWR.n4397 VPWR.n4396 0.00975758
R7855 VPWR.n4454 VPWR.n4453 0.00975758
R7856 VPWR.n5280 VPWR.n298 0.00975758
R7857 VPWR.n233 VPWR.n232 0.00975758
R7858 VPWR.n643 VPWR.n642 0.00975758
R7859 VPWR.n321 VPWR.n320 0.00975758
R7860 VPWR.n4937 VPWR.n4936 0.00975758
R7861 VPWR.n5039 VPWR.n687 0.00975758
R7862 VPWR.n5766 VPWR.n5765 0.00975758
R7863 VPWR.n5296 VPWR.n5295 0.00975758
R7864 VPWR.n335 VPWR.n334 0.00975758
R7865 VPWR.n332 VPWR.n331 0.00975758
R7866 VPWR.n182 VPWR.n181 0.00975758
R7867 VPWR.n529 VPWR.n528 0.00975758
R7868 VPWR.n152 VPWR.n151 0.00975758
R7869 VPWR.n5448 VPWR.n5447 0.00975758
R7870 VPWR.n5379 VPWR.n5378 0.00975758
R7871 VPWR.n5663 VPWR.n5662 0.00975758
R7872 VPWR.n5855 VPWR.n5854 0.00975758
R7873 VPWR.n5956 VPWR.n178 0.00975758
R7874 VPWR.n5840 VPWR.n5839 0.00975758
R7875 VPWR.n5829 VPWR.n5828 0.00975758
R7876 VPWR.n2467 VPWR.n2466 0.00975758
R7877 VPWR.n2376 VPWR.n2375 0.00975758
R7878 VPWR.n2317 VPWR.n2316 0.00975758
R7879 VPWR.n2223 VPWR.n2222 0.00975758
R7880 VPWR.n5646 VPWR.n5645 0.00975758
R7881 VPWR.n5567 VPWR.n5566 0.00975758
R7882 VPWR.n115 VPWR.n114 0.00975758
R7883 VPWR.n6076 VPWR.n105 0.00975758
R7884 VPWR.n4227 VPWR.n777 0.00975384
R7885 VPWR.n2092 VPWR.n2091 0.00961458
R7886 VPWR.n2368 VPWR.n2367 0.00961458
R7887 VPWR.n2627 VPWR.n2626 0.00961458
R7888 VPWR VPWR.n2779 0.00961458
R7889 VPWR.n2780 VPWR 0.00961458
R7890 VPWR VPWR.n2753 0.00961458
R7891 VPWR.n2751 VPWR.n2750 0.00961458
R7892 VPWR.n2748 VPWR.n2625 0.00961458
R7893 VPWR VPWR.n2630 0.00961458
R7894 VPWR.n1588 VPWR.n1587 0.00961458
R7895 VPWR.n2797 VPWR.n2796 0.00961458
R7896 VPWR.n1790 VPWR.n1789 0.00961458
R7897 VPWR VPWR.n1913 0.00961458
R7898 VPWR.n1914 VPWR 0.00961458
R7899 VPWR VPWR.n1803 0.00961458
R7900 VPWR.n1801 VPWR.n1800 0.00961458
R7901 VPWR.n1798 VPWR.n1788 0.00961458
R7902 VPWR VPWR 0.00961458
R7903 VPWR VPWR 0.00961458
R7904 VPWR.n1670 VPWR.n1669 0.00961458
R7905 VPWR.n1921 VPWR.n1920 0.00961458
R7906 VPWR.n1457 VPWR.n1456 0.00961458
R7907 VPWR.n3291 VPWR 0.00961458
R7908 VPWR VPWR.n3289 0.00961458
R7909 VPWR VPWR.n1470 0.00961458
R7910 VPWR.n1468 VPWR.n1467 0.00961458
R7911 VPWR VPWR 0.00961458
R7912 VPWR.n1392 VPWR.n1391 0.00961458
R7913 VPWR.n3283 VPWR.n3282 0.00961458
R7914 VPWR.n1242 VPWR.n1241 0.00961458
R7915 VPWR.n3758 VPWR 0.00961458
R7916 VPWR VPWR.n3756 0.00961458
R7917 VPWR VPWR 0.00961458
R7918 VPWR VPWR.n3644 0.00961458
R7919 VPWR.n3642 VPWR.n3641 0.00961458
R7920 VPWR.n3542 VPWR.n3541 0.00961458
R7921 VPWR.n3750 VPWR.n3749 0.00961458
R7922 VPWR.n1096 VPWR.n1095 0.00961458
R7923 VPWR.n3855 VPWR 0.00961458
R7924 VPWR VPWR.n3854 0.00961458
R7925 VPWR VPWR.n1109 0.00961458
R7926 VPWR.n1107 VPWR.n1106 0.00961458
R7927 VPWR VPWR 0.00961458
R7928 VPWR.n971 VPWR.n970 0.00961458
R7929 VPWR.n3848 VPWR.n3847 0.00961458
R7930 VPWR.n789 VPWR.n788 0.00961458
R7931 VPWR VPWR.n840 0.00961458
R7932 VPWR.n841 VPWR 0.00961458
R7933 VPWR VPWR.n802 0.00961458
R7934 VPWR.n800 VPWR.n799 0.00961458
R7935 VPWR VPWR 0.00961458
R7936 VPWR.n4125 VPWR.n4124 0.00961458
R7937 VPWR VPWR 0.00961458
R7938 VPWR.n848 VPWR.n847 0.00961458
R7939 VPWR.n4627 VPWR.n4626 0.00961458
R7940 VPWR.n4893 VPWR 0.00961458
R7941 VPWR VPWR.n4892 0.00961458
R7942 VPWR VPWR.n4640 0.00961458
R7943 VPWR.n4638 VPWR.n4637 0.00961458
R7944 VPWR.n4493 VPWR.n4492 0.00961458
R7945 VPWR VPWR 0.00961458
R7946 VPWR.n4886 VPWR.n4885 0.00961458
R7947 VPWR.n665 VPWR.n664 0.00961458
R7948 VPWR.n5015 VPWR 0.00961458
R7949 VPWR VPWR.n5014 0.00961458
R7950 VPWR VPWR 0.00961458
R7951 VPWR.n659 VPWR 0.00961458
R7952 VPWR.n662 VPWR.n661 0.00961458
R7953 VPWR.n674 VPWR.n673 0.00961458
R7954 VPWR.n239 VPWR.n238 0.00961458
R7955 VPWR.n5008 VPWR.n5007 0.00961458
R7956 VPWR.n342 VPWR.n341 0.00961458
R7957 VPWR VPWR.n513 0.00961458
R7958 VPWR.n514 VPWR 0.00961458
R7959 VPWR VPWR 0.00961458
R7960 VPWR VPWR.n479 0.00961458
R7961 VPWR.n477 VPWR.n476 0.00961458
R7962 VPWR.n474 VPWR.n340 0.00961458
R7963 VPWR VPWR.n346 0.00961458
R7964 VPWR VPWR 0.00961458
R7965 VPWR.n5302 VPWR.n5301 0.00961458
R7966 VPWR VPWR 0.00961458
R7967 VPWR.n521 VPWR.n520 0.00961458
R7968 VPWR.n5417 VPWR.n5416 0.00961458
R7969 VPWR.n5922 VPWR 0.00961458
R7970 VPWR VPWR.n5921 0.00961458
R7971 VPWR.n5431 VPWR 0.00961458
R7972 VPWR.n5434 VPWR.n5433 0.00961458
R7973 VPWR.n5667 VPWR.n5666 0.00961458
R7974 VPWR.n5684 VPWR 0.00961458
R7975 VPWR.n5915 VPWR.n5914 0.00961458
R7976 VPWR.n6266 VPWR.n6265 0.00961458
R7977 VPWR.n2095 VPWR.n2094 0.00961458
R7978 VPWR.n2229 VPWR.n2228 0.00961458
R7979 VPWR.n6273 VPWR 0.00961458
R7980 VPWR VPWR.n6272 0.00961458
R7981 VPWR VPWR 0.00961458
R7982 VPWR VPWR.n133 0.00961458
R7983 VPWR.n131 VPWR.n130 0.00961458
R7984 VPWR.n5574 VPWR.n5573 0.00961458
R7985 VPWR.n120 VPWR.n119 0.00961458
R7986 VPWR.n4112 VPWR.n4111 0.00900406
R7987 VPWR.n856 VPWR.n853 0.00900406
R7988 VPWR.n1507 VPWR.n1506 0.00837842
R7989 VPWR.n4209 VPWR.n4208 0.00837842
R7990 VPWR.n1509 VPWR.n1508 0.00837842
R7991 VPWR.n2786 VPWR.n2785 0.0083125
R7992 VPWR.n2754 VPWR 0.0083125
R7993 VPWR.n1827 VPWR.n1825 0.0083125
R7994 VPWR.n1804 VPWR 0.0083125
R7995 VPWR.n3228 VPWR.n3226 0.0083125
R7996 VPWR.n1471 VPWR 0.0083125
R7997 VPWR.n1204 VPWR.n1202 0.0083125
R7998 VPWR.n3645 VPWR 0.0083125
R7999 VPWR.n1110 VPWR 0.0083125
R8000 VPWR.n832 VPWR.n830 0.0083125
R8001 VPWR.n803 VPWR 0.0083125
R8002 VPWR.n4461 VPWR.n4459 0.0083125
R8003 VPWR.n4641 VPWR 0.0083125
R8004 VPWR.n4995 VPWR 0.0083125
R8005 VPWR VPWR.n658 0.0083125
R8006 VPWR.n480 VPWR 0.0083125
R8007 VPWR.n5906 VPWR.n5905 0.0083125
R8008 VPWR VPWR.n5430 0.0083125
R8009 VPWR.n2357 VPWR.n2356 0.0083125
R8010 VPWR.n134 VPWR 0.0083125
R8011 VPWR.n1788 VPWR.n1787 0.00828576
R8012 VPWR.n1246 VPWR.n1245 0.00828576
R8013 VPWR.n1070 VPWR.n1069 0.00828576
R8014 VPWR.n772 VPWR.n770 0.00828576
R8015 VPWR.n4212 VPWR.n4211 0.00803709
R8016 VPWR.n1751 VPWR.n1750 0.00736036
R8017 VPWR.n3042 VPWR.n3041 0.00736036
R8018 VPWR.n2038 VPWR.n2037 0.00736036
R8019 VPWR.n2930 VPWR.n2929 0.00736036
R8020 VPWR.n2055 VPWR.n2054 0.00701042
R8021 VPWR.n2054 VPWR.n2053 0.00701042
R8022 VPWR.n2099 VPWR.n2098 0.00701042
R8023 VPWR.n2383 VPWR.n2382 0.00701042
R8024 VPWR.n2366 VPWR.n2365 0.00701042
R8025 VPWR.n3079 VPWR.n3078 0.00701042
R8026 VPWR.n1594 VPWR.n1593 0.00701042
R8027 VPWR.n1595 VPWR.n1594 0.00701042
R8028 VPWR.n2758 VPWR.n2757 0.00701042
R8029 VPWR.n2757 VPWR.n2756 0.00701042
R8030 VPWR.n2747 VPWR.n2746 0.00701042
R8031 VPWR.n1568 VPWR.n1565 0.00701042
R8032 VPWR.n2764 VPWR.n2763 0.00701042
R8033 VPWR.n1589 VPWR.n1588 0.00701042
R8034 VPWR.n1590 VPWR.n1589 0.00701042
R8035 VPWR.n3107 VPWR.n3103 0.00701042
R8036 VPWR.n2795 VPWR.n2794 0.00701042
R8037 VPWR.n1762 VPWR.n1759 0.00701042
R8038 VPWR.n1676 VPWR.n1675 0.00701042
R8039 VPWR.n1677 VPWR.n1676 0.00701042
R8040 VPWR.n1808 VPWR.n1807 0.00701042
R8041 VPWR.n1807 VPWR.n1806 0.00701042
R8042 VPWR.n1797 VPWR.n1796 0.00701042
R8043 VPWR.n1890 VPWR.n1887 0.00701042
R8044 VPWR.n1671 VPWR.n1670 0.00701042
R8045 VPWR.n1672 VPWR.n1671 0.00701042
R8046 VPWR.n1905 VPWR.n1901 0.00701042
R8047 VPWR.n1919 VPWR.n1918 0.00701042
R8048 VPWR.n1475 VPWR.n1474 0.00701042
R8049 VPWR.n1474 VPWR.n1473 0.00701042
R8050 VPWR.n1464 VPWR.n1463 0.00701042
R8051 VPWR.n1401 VPWR.n1398 0.00701042
R8052 VPWR.n1386 VPWR.n1385 0.00701042
R8053 VPWR.n1385 VPWR.n1384 0.00701042
R8054 VPWR.n3200 VPWR.n3197 0.00701042
R8055 VPWR.n1391 VPWR.n1390 0.00701042
R8056 VPWR.n1390 VPWR.n1389 0.00701042
R8057 VPWR.n3209 VPWR.n3205 0.00701042
R8058 VPWR.n3285 VPWR.n3284 0.00701042
R8059 VPWR.n3649 VPWR.n3648 0.00701042
R8060 VPWR.n3648 VPWR.n3647 0.00701042
R8061 VPWR.n3638 VPWR.n3637 0.00701042
R8062 VPWR.n3547 VPWR.n3546 0.00701042
R8063 VPWR.n3536 VPWR.n3535 0.00701042
R8064 VPWR.n3535 VPWR.n3534 0.00701042
R8065 VPWR.n1189 VPWR.n1186 0.00701042
R8066 VPWR.n3541 VPWR.n3540 0.00701042
R8067 VPWR.n3540 VPWR.n3539 0.00701042
R8068 VPWR.n3770 VPWR.n3766 0.00701042
R8069 VPWR.n3752 VPWR.n3751 0.00701042
R8070 VPWR.n1114 VPWR.n1113 0.00701042
R8071 VPWR.n1113 VPWR.n1112 0.00701042
R8072 VPWR.n1103 VPWR.n1102 0.00701042
R8073 VPWR.n1061 VPWR.n1058 0.00701042
R8074 VPWR.n977 VPWR.n976 0.00701042
R8075 VPWR.n978 VPWR.n977 0.00701042
R8076 VPWR.n972 VPWR.n971 0.00701042
R8077 VPWR.n973 VPWR.n972 0.00701042
R8078 VPWR.n3869 VPWR.n3865 0.00701042
R8079 VPWR.n3850 VPWR.n3849 0.00701042
R8080 VPWR.n4349 VPWR.n4346 0.00701042
R8081 VPWR.n4131 VPWR.n4130 0.00701042
R8082 VPWR.n4132 VPWR.n4131 0.00701042
R8083 VPWR.n807 VPWR.n806 0.00701042
R8084 VPWR.n806 VPWR.n805 0.00701042
R8085 VPWR.n796 VPWR.n795 0.00701042
R8086 VPWR.n748 VPWR.n745 0.00701042
R8087 VPWR.n4126 VPWR.n4125 0.00701042
R8088 VPWR.n4127 VPWR.n4126 0.00701042
R8089 VPWR.n4374 VPWR.n4370 0.00701042
R8090 VPWR.n846 VPWR.n845 0.00701042
R8091 VPWR.n4816 VPWR.n4813 0.00701042
R8092 VPWR.n4499 VPWR.n4498 0.00701042
R8093 VPWR.n4500 VPWR.n4499 0.00701042
R8094 VPWR.n4645 VPWR.n4644 0.00701042
R8095 VPWR.n4644 VPWR.n4643 0.00701042
R8096 VPWR.n4634 VPWR.n4633 0.00701042
R8097 VPWR.n4446 VPWR.n4443 0.00701042
R8098 VPWR.n4650 VPWR.n4649 0.00701042
R8099 VPWR.n4494 VPWR.n4493 0.00701042
R8100 VPWR.n4495 VPWR.n4494 0.00701042
R8101 VPWR.n4905 VPWR.n4901 0.00701042
R8102 VPWR.n4888 VPWR.n4887 0.00701042
R8103 VPWR.n309 VPWR.n306 0.00701042
R8104 VPWR.n245 VPWR.n244 0.00701042
R8105 VPWR.n246 VPWR.n245 0.00701042
R8106 VPWR.n652 VPWR.n651 0.00701042
R8107 VPWR.n656 VPWR.n652 0.00701042
R8108 VPWR.n672 VPWR.n671 0.00701042
R8109 VPWR.n4993 VPWR.n4990 0.00701042
R8110 VPWR.n240 VPWR.n239 0.00701042
R8111 VPWR.n241 VPWR.n240 0.00701042
R8112 VPWR.n5027 VPWR.n5023 0.00701042
R8113 VPWR.n5010 VPWR.n5009 0.00701042
R8114 VPWR.n5775 VPWR.n5774 0.00701042
R8115 VPWR.n5308 VPWR.n5307 0.00701042
R8116 VPWR.n5309 VPWR.n5308 0.00701042
R8117 VPWR.n484 VPWR.n483 0.00701042
R8118 VPWR.n483 VPWR.n482 0.00701042
R8119 VPWR.n473 VPWR.n472 0.00701042
R8120 VPWR.n5303 VPWR.n5302 0.00701042
R8121 VPWR.n5304 VPWR.n5303 0.00701042
R8122 VPWR.n5803 VPWR.n5799 0.00701042
R8123 VPWR.n519 VPWR.n518 0.00701042
R8124 VPWR.n5425 VPWR.n5424 0.00701042
R8125 VPWR.n5426 VPWR.n5425 0.00701042
R8126 VPWR.n5438 VPWR.n5437 0.00701042
R8127 VPWR.n5397 VPWR.n5394 0.00701042
R8128 VPWR.n5682 VPWR.n5681 0.00701042
R8129 VPWR.n5681 VPWR.n5680 0.00701042
R8130 VPWR.n5420 VPWR.n154 0.00701042
R8131 VPWR.n5669 VPWR.n5667 0.00701042
R8132 VPWR.n5671 VPWR.n5669 0.00701042
R8133 VPWR.n5944 VPWR.n5940 0.00701042
R8134 VPWR.n5917 VPWR.n5916 0.00701042
R8135 VPWR.n6279 VPWR.n6278 0.00701042
R8136 VPWR.n6268 VPWR.n6267 0.00701042
R8137 VPWR.n2445 VPWR.n2442 0.00701042
R8138 VPWR.n2064 VPWR.n2063 0.00701042
R8139 VPWR.n2230 VPWR.n2229 0.00701042
R8140 VPWR.n2231 VPWR.n2230 0.00701042
R8141 VPWR.n2326 VPWR.n2325 0.00701042
R8142 VPWR.n2235 VPWR.n2234 0.00701042
R8143 VPWR.n2236 VPWR.n2235 0.00701042
R8144 VPWR.n6189 VPWR.n6187 0.00701042
R8145 VPWR.n5580 VPWR.n5579 0.00701042
R8146 VPWR.n5581 VPWR.n5580 0.00701042
R8147 VPWR.n138 VPWR.n137 0.00701042
R8148 VPWR.n137 VPWR.n136 0.00701042
R8149 VPWR.n127 VPWR.n126 0.00701042
R8150 VPWR.n1506 VPWR.n1505 0.00696227
R8151 VPWR.n1926 VPWR.n1515 0.00690179
R8152 VPWR.n1836 VPWR.n1503 0.00690178
R8153 VPWR.n1510 VPWR.n1509 0.00657697
R8154 VPWR.n4213 VPWR.n4212 0.00657697
R8155 VPWR.n4210 VPWR.n4209 0.00657697
R8156 VPWR.n3056 VPWR.n3055 0.00590801
R8157 VPWR.n2779 VPWR.n1569 0.00570833
R8158 VPWR.n1913 VPWR.n1911 0.00570833
R8159 VPWR.n3292 VPWR.n3291 0.00570833
R8160 VPWR.n3759 VPWR.n3758 0.00570833
R8161 VPWR.n3856 VPWR.n3855 0.00570833
R8162 VPWR.n840 VPWR.n749 0.00570833
R8163 VPWR.n4894 VPWR.n4893 0.00570833
R8164 VPWR.n5016 VPWR.n5015 0.00570833
R8165 VPWR.n513 VPWR.n223 0.00570833
R8166 VPWR.n5923 VPWR.n5922 0.00570833
R8167 VPWR.n2447 VPWR.n2446 0.00570833
R8168 VPWR.n6274 VPWR.n6273 0.00570833
R8169 VPWR.n3136 VPWR.n3135 0.00554564
R8170 VPWR.n3049 VPWR.n3045 0.00500002
R8171 VPWR.n2927 VPWR.n2922 0.00500002
R8172 VPWR.n1781 VPWR.n1777 0.00500002
R8173 VPWR.n5826 VPWR.n5825 0.00460158
R8174 VPWR.n5853 VPWR.n5845 0.00460158
R8175 VPWR.n5822 VPWR.n5821 0.00460158
R8176 VPWR.n4935 VPWR.n4927 0.00460158
R8177 VPWR.n4924 VPWR.n4923 0.00460158
R8178 VPWR.n3801 VPWR.n3793 0.00460158
R8179 VPWR.n3789 VPWR.n3788 0.00460158
R8180 VPWR.n3148 VPWR.n3140 0.00460158
R8181 VPWR.n3126 VPWR.n3125 0.00460158
R8182 VPWR.n5661 VPWR.n5656 0.00460158
R8183 VPWR.n2221 VPWR.n2213 0.00460158
R8184 VPWR.n5655 VPWR.n5654 0.00460158
R8185 VPWR.n113 VPWR.n106 0.00460158
R8186 VPWR.n6073 VPWR.n6072 0.00460158
R8187 VPWR.n1089 VPWR.n1081 0.00460158
R8188 VPWR.n1433 VPWR.n1425 0.00460158
R8189 VPWR.n1450 VPWR.n1442 0.00460158
R8190 VPWR.n2608 VPWR.n2607 0.00460158
R8191 VPWR.n1252 VPWR.n1250 0.00442876
R8192 VPWR.n2053 VPWR.n2052 0.00440625
R8193 VPWR.n2098 VPWR.n2093 0.00440625
R8194 VPWR.n2382 VPWR.n2381 0.00440625
R8195 VPWR.n2365 VPWR.n2364 0.00440625
R8196 VPWR.n3078 VPWR.n3074 0.00440625
R8197 VPWR.n1593 VPWR.n1585 0.00440625
R8198 VPWR.n2756 VPWR.n2622 0.00440625
R8199 VPWR.n2747 VPWR.n2628 0.00440625
R8200 VPWR.n3108 VPWR.n3098 0.00440625
R8201 VPWR.n2783 VPWR.n2782 0.00440625
R8202 VPWR.n2755 VPWR.n2754 0.00440625
R8203 VPWR.n2749 VPWR.n2748 0.00440625
R8204 VPWR.n3077 VPWR.n3076 0.00440625
R8205 VPWR.n1592 VPWR.n1591 0.00440625
R8206 VPWR.n3107 VPWR.n3106 0.00440625
R8207 VPWR.n2794 VPWR.n2793 0.00440625
R8208 VPWR.n1762 VPWR.n1761 0.00440625
R8209 VPWR.n1675 VPWR.n1667 0.00440625
R8210 VPWR.n1806 VPWR.n1784 0.00440625
R8211 VPWR.n1797 VPWR.n1791 0.00440625
R8212 VPWR.n1907 VPWR.n1906 0.00440625
R8213 VPWR.n1917 VPWR.n1916 0.00440625
R8214 VPWR.n1805 VPWR.n1804 0.00440625
R8215 VPWR.n1799 VPWR.n1798 0.00440625
R8216 VPWR.n2940 VPWR.n2939 0.00440625
R8217 VPWR.n1763 VPWR.n1755 0.00440625
R8218 VPWR.n1674 VPWR.n1673 0.00440625
R8219 VPWR.n1905 VPWR.n1904 0.00440625
R8220 VPWR.n1918 VPWR.n1834 0.00440625
R8221 VPWR.n1473 VPWR.n1455 0.00440625
R8222 VPWR.n1464 VPWR.n1458 0.00440625
R8223 VPWR.n1401 VPWR.n1400 0.00440625
R8224 VPWR.n1386 VPWR.n1322 0.00440625
R8225 VPWR.n3210 VPWR.n1496 0.00440625
R8226 VPWR.n3287 VPWR.n3286 0.00440625
R8227 VPWR.n1472 VPWR.n1471 0.00440625
R8228 VPWR.n1466 VPWR.n1465 0.00440625
R8229 VPWR.n3356 VPWR.n3355 0.00440625
R8230 VPWR.n1402 VPWR.n1394 0.00440625
R8231 VPWR.n1388 VPWR.n1387 0.00440625
R8232 VPWR.n3209 VPWR.n3208 0.00440625
R8233 VPWR.n3285 VPWR.n1499 0.00440625
R8234 VPWR.n3647 VPWR.n1240 0.00440625
R8235 VPWR.n3638 VPWR.n1243 0.00440625
R8236 VPWR.n3546 VPWR.n1284 0.00440625
R8237 VPWR.n3536 VPWR.n1297 0.00440625
R8238 VPWR.n3771 VPWR.n3761 0.00440625
R8239 VPWR.n3754 VPWR.n3753 0.00440625
R8240 VPWR.n3646 VPWR.n3645 0.00440625
R8241 VPWR.n3640 VPWR.n3639 0.00440625
R8242 VPWR.n3545 VPWR.n3544 0.00440625
R8243 VPWR.n3538 VPWR.n3537 0.00440625
R8244 VPWR.n3770 VPWR.n3769 0.00440625
R8245 VPWR.n3752 VPWR.n1193 0.00440625
R8246 VPWR.n1112 VPWR.n1094 0.00440625
R8247 VPWR.n1103 VPWR.n1097 0.00440625
R8248 VPWR.n1061 VPWR.n1060 0.00440625
R8249 VPWR.n976 VPWR.n968 0.00440625
R8250 VPWR.n3870 VPWR.n3860 0.00440625
R8251 VPWR.n3852 VPWR.n3851 0.00440625
R8252 VPWR.n1111 VPWR.n1110 0.00440625
R8253 VPWR.n1105 VPWR.n1104 0.00440625
R8254 VPWR.n1062 VPWR.n1054 0.00440625
R8255 VPWR.n975 VPWR.n974 0.00440625
R8256 VPWR.n3869 VPWR.n3868 0.00440625
R8257 VPWR.n3850 VPWR.n3843 0.00440625
R8258 VPWR.n4349 VPWR.n4348 0.00440625
R8259 VPWR.n4130 VPWR.n4122 0.00440625
R8260 VPWR.n805 VPWR.n787 0.00440625
R8261 VPWR.n796 VPWR.n790 0.00440625
R8262 VPWR.n4375 VPWR.n4365 0.00440625
R8263 VPWR.n844 VPWR.n843 0.00440625
R8264 VPWR.n804 VPWR.n803 0.00440625
R8265 VPWR.n798 VPWR.n797 0.00440625
R8266 VPWR.n4235 VPWR.n4234 0.00440625
R8267 VPWR.n4354 VPWR.n4353 0.00440625
R8268 VPWR.n4350 VPWR.n756 0.00440625
R8269 VPWR.n4129 VPWR.n4128 0.00440625
R8270 VPWR.n4374 VPWR.n4373 0.00440625
R8271 VPWR.n845 VPWR.n839 0.00440625
R8272 VPWR.n4816 VPWR.n4815 0.00440625
R8273 VPWR.n4498 VPWR.n4490 0.00440625
R8274 VPWR.n4643 VPWR.n4625 0.00440625
R8275 VPWR.n4634 VPWR.n4628 0.00440625
R8276 VPWR.n4906 VPWR.n4896 0.00440625
R8277 VPWR.n4890 VPWR.n4889 0.00440625
R8278 VPWR.n4642 VPWR.n4641 0.00440625
R8279 VPWR.n4636 VPWR.n4635 0.00440625
R8280 VPWR.n4712 VPWR.n4711 0.00440625
R8281 VPWR.n4822 VPWR.n4821 0.00440625
R8282 VPWR.n4817 VPWR.n4482 0.00440625
R8283 VPWR.n4497 VPWR.n4496 0.00440625
R8284 VPWR.n4905 VPWR.n4904 0.00440625
R8285 VPWR.n4888 VPWR.n4450 0.00440625
R8286 VPWR.n309 VPWR.n308 0.00440625
R8287 VPWR.n244 VPWR.n236 0.00440625
R8288 VPWR.n656 VPWR.n655 0.00440625
R8289 VPWR.n672 VPWR.n666 0.00440625
R8290 VPWR.n5028 VPWR.n5018 0.00440625
R8291 VPWR.n5012 VPWR.n5011 0.00440625
R8292 VPWR.n658 VPWR.n657 0.00440625
R8293 VPWR.n673 VPWR.n663 0.00440625
R8294 VPWR.n5160 VPWR.n5159 0.00440625
R8295 VPWR.n310 VPWR.n302 0.00440625
R8296 VPWR.n243 VPWR.n242 0.00440625
R8297 VPWR.n5027 VPWR.n5026 0.00440625
R8298 VPWR.n5010 VPWR.n5003 0.00440625
R8299 VPWR.n5774 VPWR.n5770 0.00440625
R8300 VPWR.n5307 VPWR.n5299 0.00440625
R8301 VPWR.n482 VPWR.n338 0.00440625
R8302 VPWR.n473 VPWR.n343 0.00440625
R8303 VPWR.n5804 VPWR.n5794 0.00440625
R8304 VPWR.n517 VPWR.n516 0.00440625
R8305 VPWR.n481 VPWR.n480 0.00440625
R8306 VPWR.n475 VPWR.n474 0.00440625
R8307 VPWR.n462 VPWR.n460 0.00440625
R8308 VPWR.n5773 VPWR.n5772 0.00440625
R8309 VPWR.n5306 VPWR.n5305 0.00440625
R8310 VPWR.n5803 VPWR.n5802 0.00440625
R8311 VPWR.n518 VPWR.n512 0.00440625
R8312 VPWR.n5429 VPWR.n5426 0.00440625
R8313 VPWR.n5437 VPWR.n5418 0.00440625
R8314 VPWR.n5397 VPWR.n5396 0.00440625
R8315 VPWR.n5682 VPWR.n5675 0.00440625
R8316 VPWR.n5945 VPWR.n5935 0.00440625
R8317 VPWR.n5919 VPWR.n5918 0.00440625
R8318 VPWR.n5436 VPWR.n5435 0.00440625
R8319 VPWR.n5458 VPWR.n5456 0.00440625
R8320 VPWR.n5401 VPWR.n5382 0.00440625
R8321 VPWR.n5398 VPWR.n5390 0.00440625
R8322 VPWR.n5683 VPWR.n5672 0.00440625
R8323 VPWR VPWR.n5683 0.00440625
R8324 VPWR.n5944 VPWR.n5943 0.00440625
R8325 VPWR.n5917 VPWR.n5910 0.00440625
R8326 VPWR.n6278 VPWR.n27 0.00440625
R8327 VPWR.n6268 VPWR.n37 0.00440625
R8328 VPWR.n2456 VPWR.n2455 0.00440625
R8329 VPWR.n2354 VPWR.n2353 0.00440625
R8330 VPWR.n2062 VPWR.n2061 0.00440625
R8331 VPWR.n2097 VPWR.n2096 0.00440625
R8332 VPWR.n2110 VPWR.n2109 0.00440625
R8333 VPWR.n2324 VPWR.n2323 0.00440625
R8334 VPWR.n2233 VPWR.n2232 0.00440625
R8335 VPWR.n2325 VPWR.n2321 0.00440625
R8336 VPWR.n2234 VPWR.n2226 0.00440625
R8337 VPWR.n6189 VPWR.n6188 0.00440625
R8338 VPWR.n5579 VPWR.n5571 0.00440625
R8339 VPWR.n6277 VPWR.n6276 0.00440625
R8340 VPWR.n6270 VPWR.n6269 0.00440625
R8341 VPWR.n135 VPWR.n134 0.00440625
R8342 VPWR.n129 VPWR.n128 0.00440625
R8343 VPWR.n6083 VPWR.n6082 0.00440625
R8344 VPWR.n6190 VPWR.n80 0.00440625
R8345 VPWR.n5578 VPWR.n5577 0.00440625
R8346 VPWR.n136 VPWR.n118 0.00440625
R8347 VPWR.n127 VPWR.n121 0.00440625
R8348 VPWR.n4831 VPWR.n4830 0.00434825
R8349 VPWR.n1511 VPWR.n1504 0.00434475
R8350 VPWR.n4204 VPWR.n4203 0.0042754
R8351 VPWR.n5576 VPWR.n5575 0.00420071
R8352 VPWR.n2043 VPWR.n2042 0.00406061
R8353 VPWR.n2606 VPWR.n2603 0.00406061
R8354 VPWR.n3065 VPWR.n3064 0.00406061
R8355 VPWR.n3062 VPWR.n3061 0.00406061
R8356 VPWR.n2918 VPWR.n2917 0.00406061
R8357 VPWR.n2613 VPWR.n2610 0.00406061
R8358 VPWR.n3124 VPWR.n3123 0.00406061
R8359 VPWR.n3121 VPWR.n3120 0.00406061
R8360 VPWR.n3048 VPWR.n3047 0.00406061
R8361 VPWR.n3054 VPWR.n3052 0.00406061
R8362 VPWR.n1780 VPWR.n1779 0.00406061
R8363 VPWR.n2926 VPWR.n2924 0.00406061
R8364 VPWR.n3134 VPWR.n3133 0.00406061
R8365 VPWR.n1513 VPWR.n1512 0.00406061
R8366 VPWR.n1449 VPWR.n1448 0.00406061
R8367 VPWR.n1446 VPWR.n1445 0.00406061
R8368 VPWR.n3454 VPWR.n3453 0.00406061
R8369 VPWR.n1314 VPWR.n1311 0.00406061
R8370 VPWR.n3147 VPWR.n3146 0.00406061
R8371 VPWR.n3144 VPWR.n3143 0.00406061
R8372 VPWR.n1432 VPWR.n1431 0.00406061
R8373 VPWR.n1429 VPWR.n1428 0.00406061
R8374 VPWR.n1306 VPWR.n1305 0.00406061
R8375 VPWR.n3461 VPWR.n3458 0.00406061
R8376 VPWR.n3787 VPWR.n3786 0.00406061
R8377 VPWR.n3784 VPWR.n3783 0.00406061
R8378 VPWR.n1088 VPWR.n1087 0.00406061
R8379 VPWR.n1085 VPWR.n1084 0.00406061
R8380 VPWR.n4100 VPWR.n4099 0.00406061
R8381 VPWR.n1047 VPWR.n1044 0.00406061
R8382 VPWR.n3800 VPWR.n3799 0.00406061
R8383 VPWR.n3797 VPWR.n3796 0.00406061
R8384 VPWR.n4119 VPWR.n4118 0.00406061
R8385 VPWR.n4109 VPWR.n4106 0.00406061
R8386 VPWR.n783 VPWR.n782 0.00406061
R8387 VPWR.n4222 VPWR.n4220 0.00406061
R8388 VPWR.n698 VPWR.n697 0.00406061
R8389 VPWR.n693 VPWR.n691 0.00406061
R8390 VPWR.n4574 VPWR.n4573 0.00406061
R8391 VPWR.n4571 VPWR.n4570 0.00406061
R8392 VPWR.n4613 VPWR.n4612 0.00406061
R8393 VPWR.n4619 VPWR.n4616 0.00406061
R8394 VPWR.n4922 VPWR.n4921 0.00406061
R8395 VPWR.n4919 VPWR.n4918 0.00406061
R8396 VPWR.n5289 VPWR.n5288 0.00406061
R8397 VPWR.n5286 VPWR.n5285 0.00406061
R8398 VPWR.n635 VPWR.n634 0.00406061
R8399 VPWR.n640 VPWR.n637 0.00406061
R8400 VPWR.n4934 VPWR.n4933 0.00406061
R8401 VPWR.n4931 VPWR.n4930 0.00406061
R8402 VPWR.n5761 VPWR.n5760 0.00406061
R8403 VPWR.n5758 VPWR.n5757 0.00406061
R8404 VPWR.n329 VPWR.n328 0.00406061
R8405 VPWR.n627 VPWR.n624 0.00406061
R8406 VPWR.n5820 VPWR.n5819 0.00406061
R8407 VPWR.n5817 VPWR.n5816 0.00406061
R8408 VPWR.n6071 VPWR.n6070 0.00406061
R8409 VPWR.n5660 VPWR.n5659 0.00406061
R8410 VPWR.n5749 VPWR.n5746 0.00406061
R8411 VPWR.n5852 VPWR.n5851 0.00406061
R8412 VPWR.n5849 VPWR.n5848 0.00406061
R8413 VPWR.n5836 VPWR.n5835 0.00406061
R8414 VPWR.n5833 VPWR.n5832 0.00406061
R8415 VPWR.n2474 VPWR.n2473 0.00406061
R8416 VPWR.n2471 VPWR.n2470 0.00406061
R8417 VPWR.n2215 VPWR.n2214 0.00406061
R8418 VPWR.n2220 VPWR.n2217 0.00406061
R8419 VPWR.n5653 VPWR.n5652 0.00406061
R8420 VPWR.n5650 VPWR.n5649 0.00406061
R8421 VPWR.n112 VPWR.n111 0.00406061
R8422 VPWR.n5955 VPWR.n5824 0.00393497
R8423 VPWR.n4926 VPWR.n180 0.00393497
R8424 VPWR.n5038 VPWR.n4925 0.00393497
R8425 VPWR.n4395 VPWR.n4394 0.00393497
R8426 VPWR.n3880 VPWR.n3790 0.00393497
R8427 VPWR.n3139 VPWR.n1136 0.00393497
R8428 VPWR.n3220 VPWR.n3138 0.00393497
R8429 VPWR.n2377 VPWR.n1516 0.00393497
R8430 VPWR.n2476 VPWR.n2475 0.00393497
R8431 VPWR.n5844 VPWR.n5843 0.00393497
R8432 VPWR.n2468 VPWR.n2378 0.00393497
R8433 VPWR.n5762 VPWR.n5754 0.00393497
R8434 VPWR.n5764 VPWR.n5292 0.00393497
R8435 VPWR.n5291 VPWR.n5290 0.00393497
R8436 VPWR.n5281 VPWR.n297 0.00393497
R8437 VPWR.n4575 VPWR.n4567 0.00393497
R8438 VPWR.n4577 VPWR.n4483 0.00393497
R8439 VPWR.n1300 VPWR.n1048 0.00393497
R8440 VPWR.n3462 VPWR.n3457 0.00393497
R8441 VPWR.n3043 VPWR.n1315 0.00393497
R8442 VPWR.n3066 VPWR.n3058 0.00393497
R8443 VPWR.n3068 VPWR.n1578 0.00393497
R8444 VPWR.n2313 VPWR.n2312 0.00393497
R8445 VPWR.n4102 VPWR.n4101 0.00393497
R8446 VPWR.n1307 VPWR.n1301 0.00393497
R8447 VPWR.n3456 VPWR.n3455 0.00393497
R8448 VPWR.n5751 VPWR.n5750 0.00393497
R8449 VPWR.n629 VPWR.n628 0.00393497
R8450 VPWR.n4607 VPWR.n641 0.00393497
R8451 VPWR.n4620 VPWR.n4615 0.00393497
R8452 VPWR.n3982 VPWR.n1078 0.00393497
R8453 VPWR.n1441 VPWR.n1440 0.00393497
R8454 VPWR.n3348 VPWR.n1424 0.00393497
R8455 VPWR.n2614 VPWR.n2609 0.00393497
R8456 VPWR.n6075 VPWR.n6074 0.00393497
R8457 VPWR.n2920 VPWR.n2919 0.00393497
R8458 VPWR.n322 VPWR.n150 0.00393497
R8459 VPWR.n330 VPWR.n324 0.00393497
R8460 VPWR.n636 VPWR.n630 0.00393497
R8461 VPWR.n4614 VPWR.n4608 0.00393497
R8462 VPWR.n2044 VPWR.n2039 0.00393497
R8463 VPWR.n4227 VPWR.n4226 0.00390143
R8464 VPWR.n4384 VPWR.n4383 0.00390143
R8465 VPWR.n955 VPWR.n954 0.00390143
R8466 VPWR.n2806 VPWR.n2805 0.00365283
R8467 VPWR.n1928 VPWR.n1927 0.00365283
R8468 VPWR.n3222 VPWR.n3221 0.00365283
R8469 VPWR.n1198 VPWR.n1197 0.00365283
R8470 VPWR.n3882 VPWR.n3881 0.00365283
R8471 VPWR.n856 VPWR.n855 0.00365283
R8472 VPWR.n4455 VPWR.n4454 0.00365283
R8473 VPWR.n5040 VPWR.n5039 0.00365283
R8474 VPWR.n530 VPWR.n529 0.00365283
R8475 VPWR.n5957 VPWR.n5956 0.00365283
R8476 VPWR.n5828 VPWR.n5827 0.00365283
R8477 VPWR.n2467 VPWR.n2464 0.00365283
R8478 VPWR.n2318 VPWR.n2317 0.00365283
R8479 VPWR.n4113 VPWR.n4112 0.00365283
R8480 VPWR.n6077 VPWR.n6076 0.00365283
R8481 VPWR.n3071 VPWR.n3070 0.00365283
R8482 VPWR.n3350 VPWR.n3349 0.00365283
R8483 VPWR.n1439 VPWR.n1438 0.00365283
R8484 VPWR.n3984 VPWR.n3983 0.00365283
R8485 VPWR.n4580 VPWR.n4579 0.00365283
R8486 VPWR.n5280 VPWR.n5279 0.00365283
R8487 VPWR.n5767 VPWR.n5766 0.00365283
R8488 VPWR.n5449 VPWR.n5448 0.00365283
R8489 VPWR.n2932 VPWR.n2931 0.00350892
R8490 VPWR.n1749 VPWR.n1748 0.00350844
R8491 VPWR.n4116 VPWR.n4114 0.00334848
R8492 VPWR.n4206 VPWR.n4205 0.00334848
R8493 VPWR.n957 VPWR.n956 0.00334848
R8494 VPWR.n4225 VPWR.n4224 0.00334848
R8495 VPWR.n4386 VPWR.n4385 0.00334848
R8496 VPWR.n854 VPWR.n689 0.00334848
R8497 VPWR.n1838 VPWR.n1837 0.00326041
R8498 VPWR.n3129 VPWR.n3128 0.0032017
R8499 VPWR.n3130 VPWR.n3129 0.0032017
R8500 VPWR.n5643 VPWR.n5563 0.0032017
R8501 VPWR.n5563 VPWR.n5562 0.0032017
R8502 VPWR.n172 VPWR.n171 0.00318898
R8503 VPWR.n2475 VPWR 0.00314375
R8504 VPWR.n2312 VPWR 0.00314375
R8505 VPWR.n2039 VPWR 0.00314375
R8506 VPWR.n2100 VPWR.n2099 0.00310417
R8507 VPWR.n2104 VPWR.n2103 0.00310417
R8508 VPWR.n2463 VPWR.n2462 0.00310417
R8509 VPWR.n2387 VPWR.n2386 0.00310417
R8510 VPWR.n2364 VPWR.n2363 0.00310417
R8511 VPWR.n2370 VPWR.n2369 0.00310417
R8512 VPWR.n2479 VPWR.n2372 0.00310417
R8513 VPWR.n2746 VPWR.n2745 0.00310417
R8514 VPWR.n2742 VPWR.n2741 0.00310417
R8515 VPWR.n3113 VPWR.n1568 0.00310417
R8516 VPWR.n3111 VPWR.n3110 0.00310417
R8517 VPWR.n2782 VPWR.n2781 0.00310417
R8518 VPWR.n2788 VPWR.n2787 0.00310417
R8519 VPWR.n2808 VPWR.n2790 0.00310417
R8520 VPWR.n2633 VPWR.n2632 0.00310417
R8521 VPWR.n3115 VPWR.n3114 0.00310417
R8522 VPWR.n3100 VPWR.n3099 0.00310417
R8523 VPWR.n2793 VPWR.n2792 0.00310417
R8524 VPWR.n2799 VPWR.n2798 0.00310417
R8525 VPWR.n2807 VPWR.n2801 0.00310417
R8526 VPWR.n1796 VPWR.n1795 0.00310417
R8527 VPWR.n1792 VPWR.n1775 0.00310417
R8528 VPWR.n1894 VPWR.n1890 0.00310417
R8529 VPWR.n1892 VPWR.n1891 0.00310417
R8530 VPWR.n1916 VPWR.n1915 0.00310417
R8531 VPWR.n1829 VPWR.n1828 0.00310417
R8532 VPWR.n1930 VPWR.n1831 0.00310417
R8533 VPWR.n1785 VPWR.n1774 0.00310417
R8534 VPWR.n1895 VPWR.n1839 0.00310417
R8535 VPWR.n1898 VPWR.n1897 0.00310417
R8536 VPWR.n1834 VPWR.n1833 0.00310417
R8537 VPWR.n1923 VPWR.n1922 0.00310417
R8538 VPWR.n1929 VPWR.n1925 0.00310417
R8539 VPWR.n1463 VPWR.n1462 0.00310417
R8540 VPWR.n1459 VPWR.n1420 0.00310417
R8541 VPWR.n3215 VPWR.n3200 0.00310417
R8542 VPWR.n3213 VPWR.n3212 0.00310417
R8543 VPWR.n3288 VPWR.n3287 0.00310417
R8544 VPWR.n3230 VPWR.n3229 0.00310417
R8545 VPWR.n3276 VPWR.n3232 0.00310417
R8546 VPWR.n1419 VPWR.n1418 0.00310417
R8547 VPWR.n3217 VPWR.n3216 0.00310417
R8548 VPWR.n3202 VPWR.n3201 0.00310417
R8549 VPWR.n1499 VPWR.n1498 0.00310417
R8550 VPWR.n3281 VPWR.n3280 0.00310417
R8551 VPWR.n3278 VPWR.n3277 0.00310417
R8552 VPWR.n3637 VPWR.n3636 0.00310417
R8553 VPWR.n3633 VPWR.n3632 0.00310417
R8554 VPWR.n3776 VPWR.n1189 0.00310417
R8555 VPWR.n3774 VPWR.n3773 0.00310417
R8556 VPWR.n3755 VPWR.n3754 0.00310417
R8557 VPWR.n1206 VPWR.n1205 0.00310417
R8558 VPWR.n3743 VPWR.n1208 0.00310417
R8559 VPWR.n1249 VPWR.n1248 0.00310417
R8560 VPWR.n3778 VPWR.n3777 0.00310417
R8561 VPWR.n3763 VPWR.n3762 0.00310417
R8562 VPWR.n1193 VPWR.n1192 0.00310417
R8563 VPWR.n3748 VPWR.n3747 0.00310417
R8564 VPWR.n3745 VPWR.n3744 0.00310417
R8565 VPWR.n1102 VPWR.n1101 0.00310417
R8566 VPWR.n1098 VPWR.n1074 0.00310417
R8567 VPWR.n3875 VPWR.n3834 0.00310417
R8568 VPWR.n3873 VPWR.n3872 0.00310417
R8569 VPWR.n3853 VPWR.n3852 0.00310417
R8570 VPWR.n3837 VPWR.n3836 0.00310417
R8571 VPWR VPWR.n3835 0.00310417
R8572 VPWR.n3884 VPWR.n1131 0.00310417
R8573 VPWR.n1073 VPWR.n1072 0.00310417
R8574 VPWR.n3877 VPWR.n3876 0.00310417
R8575 VPWR.n3862 VPWR.n3861 0.00310417
R8576 VPWR.n3843 VPWR.n3842 0.00310417
R8577 VPWR.n3846 VPWR.n3845 0.00310417
R8578 VPWR.n3883 VPWR.n1132 0.00310417
R8579 VPWR.n795 VPWR.n794 0.00310417
R8580 VPWR.n791 VPWR.n776 0.00310417
R8581 VPWR.n4380 VPWR.n748 0.00310417
R8582 VPWR.n4378 VPWR.n4377 0.00310417
R8583 VPWR.n843 VPWR.n842 0.00310417
R8584 VPWR.n834 VPWR.n833 0.00310417
R8585 VPWR.n858 VPWR.n836 0.00310417
R8586 VPWR.n775 VPWR.n774 0.00310417
R8587 VPWR.n4382 VPWR.n4381 0.00310417
R8588 VPWR.n4367 VPWR.n4366 0.00310417
R8589 VPWR.n839 VPWR.n838 0.00310417
R8590 VPWR.n850 VPWR.n849 0.00310417
R8591 VPWR.n857 VPWR.n852 0.00310417
R8592 VPWR.n4633 VPWR.n4632 0.00310417
R8593 VPWR.n4629 VPWR.n4604 0.00310417
R8594 VPWR.n4911 VPWR.n4446 0.00310417
R8595 VPWR.n4909 VPWR.n4908 0.00310417
R8596 VPWR.n4891 VPWR.n4890 0.00310417
R8597 VPWR.n4463 VPWR.n4462 0.00310417
R8598 VPWR.n4879 VPWR.n4465 0.00310417
R8599 VPWR.n4603 VPWR.n4602 0.00310417
R8600 VPWR.n4913 VPWR.n4912 0.00310417
R8601 VPWR.n4898 VPWR.n4897 0.00310417
R8602 VPWR.n4450 VPWR.n4449 0.00310417
R8603 VPWR.n4884 VPWR.n4883 0.00310417
R8604 VPWR.n4881 VPWR.n4880 0.00310417
R8605 VPWR.n671 VPWR.n670 0.00310417
R8606 VPWR.n667 VPWR.n319 0.00310417
R8607 VPWR.n5033 VPWR.n4993 0.00310417
R8608 VPWR.n5031 VPWR.n5030 0.00310417
R8609 VPWR.n5013 VPWR.n5012 0.00310417
R8610 VPWR.n4996 VPWR.n4995 0.00310417
R8611 VPWR.n5042 VPWR.n683 0.00310417
R8612 VPWR.n675 VPWR.n318 0.00310417
R8613 VPWR.n5035 VPWR.n5034 0.00310417
R8614 VPWR.n5020 VPWR.n5019 0.00310417
R8615 VPWR.n5003 VPWR.n5002 0.00310417
R8616 VPWR.n5006 VPWR.n5005 0.00310417
R8617 VPWR.n5041 VPWR.n684 0.00310417
R8618 VPWR.n472 VPWR.n471 0.00310417
R8619 VPWR.n468 VPWR.n467 0.00310417
R8620 VPWR.n5809 VPWR.n222 0.00310417
R8621 VPWR.n5807 VPWR.n5806 0.00310417
R8622 VPWR.n516 VPWR.n515 0.00310417
R8623 VPWR.n507 VPWR.n506 0.00310417
R8624 VPWR.n532 VPWR.n509 0.00310417
R8625 VPWR.n349 VPWR.n348 0.00310417
R8626 VPWR.n5811 VPWR.n5810 0.00310417
R8627 VPWR.n5796 VPWR.n5795 0.00310417
R8628 VPWR.n512 VPWR.n511 0.00310417
R8629 VPWR.n523 VPWR.n522 0.00310417
R8630 VPWR.n531 VPWR.n525 0.00310417
R8631 VPWR.n5439 VPWR.n5438 0.00310417
R8632 VPWR.n5443 VPWR.n5442 0.00310417
R8633 VPWR.n5950 VPWR.n5901 0.00310417
R8634 VPWR.n5948 VPWR.n5947 0.00310417
R8635 VPWR.n5920 VPWR.n5919 0.00310417
R8636 VPWR.n5904 VPWR.n5903 0.00310417
R8637 VPWR VPWR.n5902 0.00310417
R8638 VPWR.n5959 VPWR.n174 0.00310417
R8639 VPWR VPWR.n5421 0.00310417
R8640 VPWR.n5415 VPWR.n5414 0.00310417
R8641 VPWR.n5952 VPWR.n5951 0.00310417
R8642 VPWR.n5937 VPWR.n5936 0.00310417
R8643 VPWR.n5910 VPWR.n5909 0.00310417
R8644 VPWR.n5913 VPWR.n5912 0.00310417
R8645 VPWR.n5958 VPWR.n175 0.00310417
R8646 VPWR.n6285 VPWR.n26 0.00310417
R8647 VPWR.n6283 VPWR.n6282 0.00310417
R8648 VPWR.n37 VPWR.n36 0.00310417
R8649 VPWR.n6264 VPWR.n6263 0.00310417
R8650 VPWR.n6261 VPWR.n6260 0.00310417
R8651 VPWR.n2461 VPWR.n2445 0.00310417
R8652 VPWR.n2459 VPWR.n2458 0.00310417
R8653 VPWR.n2353 VPWR.n2352 0.00310417
R8654 VPWR.n2359 VPWR.n2358 0.00310417
R8655 VPWR.n2480 VPWR.n2361 0.00310417
R8656 VPWR.n2090 VPWR.n2089 0.00310417
R8657 VPWR.n6287 VPWR.n6286 0.00310417
R8658 VPWR.n30 VPWR.n29 0.00310417
R8659 VPWR.n6271 VPWR.n6270 0.00310417
R8660 VPWR.n56 VPWR.n55 0.00310417
R8661 VPWR VPWR.n54 0.00310417
R8662 VPWR.n6259 VPWR.n38 0.00310417
R8663 VPWR.n100 VPWR.n99 0.00310417
R8664 VPWR.n126 VPWR.n125 0.00310417
R8665 VPWR.n122 VPWR.n101 0.00310417
R8666 VPWR.n2036 VPWR.n2035 0.00309601
R8667 VPWR.n3040 VPWR.n3039 0.00305268
R8668 VPWR.n5954 VPWR.n5853 0.0028004
R8669 VPWR.n5821 VPWR.n5813 0.0028004
R8670 VPWR.n5037 VPWR.n4935 0.0028004
R8671 VPWR.n4923 VPWR.n4915 0.0028004
R8672 VPWR.n3879 VPWR.n3801 0.0028004
R8673 VPWR.n3788 VPWR.n3780 0.0028004
R8674 VPWR.n3219 VPWR.n3148 0.0028004
R8675 VPWR.n3125 VPWR.n3117 0.0028004
R8676 VPWR.n5842 VPWR.n5826 0.0028004
R8677 VPWR.n5744 VPWR.n5661 0.0028004
R8678 VPWR.n2311 VPWR.n2221 0.0028004
R8679 VPWR.n5654 VPWR.n5643 0.0028004
R8680 VPWR.n149 VPWR.n113 0.0028004
R8681 VPWR.n2607 VPWR.n2601 0.0028004
R8682 VPWR.n3347 VPWR.n1450 0.0028004
R8683 VPWR.n1434 VPWR.n1433 0.0028004
R8684 VPWR.n3981 VPWR.n1089 0.0028004
R8685 VPWR.n6072 VPWR.n6065 0.0028004
R8686 VPWR.n3791 VPWR.n699 0.00271707
R8687 VPWR.n4110 VPWR.n4104 0.00271707
R8688 VPWR.n1079 VPWR.n784 0.00271707
R8689 VPWR.n1043 VPWR.n965 0.00271013
R8690 VPWR.n3467 VPWR.n1299 0.00271013
R8691 VPWR.n1310 VPWR.n1309 0.00271013
R8692 VPWR.n2617 VPWR.n2616 0.00271013
R8693 VPWR.n333 VPWR.n332 0.00271013
R8694 VPWR.n5154 VPWR.n321 0.00271013
R8695 VPWR.n4706 VPWR.n4606 0.00271013
R8696 VPWR.n2478 VPWR.n2376 0.00262794
R8697 VPWR.n5843 VPWR.n5842 0.00246749
R8698 VPWR.n2477 VPWR.n2468 0.00246749
R8699 VPWR.n5955 VPWR.n5954 0.00246749
R8700 VPWR.n5813 VPWR.n180 0.00246749
R8701 VPWR.n5038 VPWR.n5037 0.00246749
R8702 VPWR.n4915 VPWR.n4395 0.00246749
R8703 VPWR.n3880 VPWR.n3879 0.00246749
R8704 VPWR.n3780 VPWR.n1136 0.00246749
R8705 VPWR.n3220 VPWR.n3219 0.00246749
R8706 VPWR.n3117 VPWR.n1516 0.00246749
R8707 VPWR.n2477 VPWR.n2476 0.00246749
R8708 VPWR.n5750 VPWR.n5744 0.00246749
R8709 VPWR.n4101 VPWR.n4095 0.00246749
R8710 VPWR.n3466 VPWR.n1307 0.00246749
R8711 VPWR.n3455 VPWR.n3449 0.00246749
R8712 VPWR.n2313 VPWR.n2311 0.00246749
R8713 VPWR.n3068 VPWR.n3067 0.00246749
R8714 VPWR.n3067 VPWR.n3066 0.00246749
R8715 VPWR.n4095 VPWR.n1048 0.00246749
R8716 VPWR.n3466 VPWR.n3462 0.00246749
R8717 VPWR.n3449 VPWR.n1315 0.00246749
R8718 VPWR.n4577 VPWR.n4576 0.00246749
R8719 VPWR.n5282 VPWR.n5281 0.00246749
R8720 VPWR.n5764 VPWR.n5763 0.00246749
R8721 VPWR.n5763 VPWR.n5762 0.00246749
R8722 VPWR.n5290 VPWR.n5282 0.00246749
R8723 VPWR.n4576 VPWR.n4575 0.00246749
R8724 VPWR.n6075 VPWR.n149 0.00246749
R8725 VPWR.n6065 VPWR.n150 0.00246749
R8726 VPWR.n623 VPWR.n330 0.00246749
R8727 VPWR.n5153 VPWR.n636 0.00246749
R8728 VPWR.n4705 VPWR.n4614 0.00246749
R8729 VPWR.n2919 VPWR.n2913 0.00246749
R8730 VPWR.n2601 VPWR.n2044 0.00246749
R8731 VPWR.n2913 VPWR.n2614 0.00246749
R8732 VPWR.n3348 VPWR.n3347 0.00246749
R8733 VPWR.n1440 VPWR.n1434 0.00246749
R8734 VPWR.n3982 VPWR.n3981 0.00246749
R8735 VPWR.n628 VPWR.n623 0.00246749
R8736 VPWR.n5153 VPWR.n641 0.00246749
R8737 VPWR.n4705 VPWR.n4620 0.00246749
R8738 VPWR.n5645 VPWR.n5644 0.00244614
R8739 VPWR.n2600 VPWR.n2049 0.00237907
R8740 VPWR.n5743 VPWR.n5663 0.00237907
R8741 VPWR.n2310 VPWR.n2223 0.00237907
R8742 VPWR.n2047 VPWR.n2046 0.00237907
R8743 VPWR.n2912 VPWR.n2619 0.00233584
R8744 VPWR.n3116 VPWR.n1518 0.00233584
R8745 VPWR.n3346 VPWR.n1452 0.00233584
R8746 VPWR.n3448 VPWR.n1317 0.00233584
R8747 VPWR.n3218 VPWR.n3150 0.00233584
R8748 VPWR.n1237 VPWR.n1236 0.00233584
R8749 VPWR.n3465 VPWR.n3464 0.00233584
R8750 VPWR.n3779 VPWR.n1138 0.00233584
R8751 VPWR.n3980 VPWR.n1091 0.00233584
R8752 VPWR.n4094 VPWR.n1050 0.00233584
R8753 VPWR.n3878 VPWR.n3803 0.00233584
R8754 VPWR.n4704 VPWR.n4622 0.00233584
R8755 VPWR.n4914 VPWR.n4397 0.00233584
R8756 VPWR.n5152 VPWR.n643 0.00233584
R8757 VPWR.n5036 VPWR.n4937 0.00233584
R8758 VPWR.n622 VPWR.n335 0.00233584
R8759 VPWR.n5812 VPWR.n182 0.00233584
R8760 VPWR.n6064 VPWR.n152 0.00233584
R8761 VPWR.n5561 VPWR.n5379 0.00233584
R8762 VPWR.n5953 VPWR.n5855 0.00233584
R8763 VPWR.n5841 VPWR.n5840 0.00233584
R8764 VPWR.n148 VPWR.n115 0.00233584
R8765 VPWR.n4389 VPWR.n4388 0.00224993
R8766 VPWR.n963 VPWR.n962 0.00224993
R8767 VPWR.n4219 VPWR.n4218 0.00224993
R8768 VPWR.n4388 VPWR.n4387 0.00224603
R8769 VPWR.n4207 VPWR.n963 0.00224603
R8770 VPWR.n4223 VPWR.n4219 0.00224603
R8771 VPWR.n4392 VPWR.n4391 0.00210121
R8772 VPWR.n4390 VPWR.n4389 0.00210121
R8773 VPWR.n4391 VPWR.n4390 0.00210121
R8774 VPWR.n4393 VPWR.n4392 0.00210121
R8775 VPWR.n960 VPWR.n959 0.00210121
R8776 VPWR.n962 VPWR.n961 0.00210121
R8777 VPWR.n959 VPWR.n958 0.00210121
R8778 VPWR.n961 VPWR.n960 0.00210121
R8779 VPWR.n4216 VPWR.n4215 0.00210121
R8780 VPWR.n4217 VPWR.n4216 0.00210121
R8781 VPWR.n4215 VPWR.n4214 0.00210121
R8782 VPWR.n4218 VPWR.n4217 0.00210121
R8783 VPWR.n1664 VPWR.n1582 0.00204637
R8784 VPWR.n4566 VPWR.n4487 0.00204637
R8785 VPWR.n296 VPWR.n233 0.00204637
R8786 VPWR.n5377 VPWR.n5296 0.00204637
R8787 VPWR.n5642 VPWR.n5567 0.00200456
R8788 VPWR.n3135 VPWR.n3130 0.00185526
R8789 VPWR.n3137 VPWR.n3136 0.00182188
R8790 VPWR.n3045 VPWR.n3044 0.00182188
R8791 VPWR.n1777 VPWR.n1776 0.00182188
R8792 VPWR.n3084 VPWR.n3072 0.00180208
R8793 VPWR.n3082 VPWR.n3081 0.00180208
R8794 VPWR.n1598 VPWR.n1597 0.00180208
R8795 VPWR.n1663 VPWR.n1600 0.00180208
R8796 VPWR VPWR.n3112 0.00180208
R8797 VPWR.n3085 VPWR.n1577 0.00180208
R8798 VPWR.n3088 VPWR.n3087 0.00180208
R8799 VPWR.n1603 VPWR.n1602 0.00180208
R8800 VPWR.n1662 VPWR.n1610 0.00180208
R8801 VPWR.n3038 VPWR.n3037 0.00180208
R8802 VPWR.n1757 VPWR.n1756 0.00180208
R8803 VPWR.n1680 VPWR.n1679 0.00180208
R8804 VPWR.n1747 VPWR.n1682 0.00180208
R8805 VPWR VPWR.n1893 0.00180208
R8806 VPWR.n3036 VPWR.n1753 0.00180208
R8807 VPWR.n3034 VPWR.n3033 0.00180208
R8808 VPWR.n1685 VPWR.n1684 0.00180208
R8809 VPWR.n1746 VPWR.n1692 0.00180208
R8810 VPWR.n3447 VPWR.n3446 0.00180208
R8811 VPWR.n1396 VPWR.n1395 0.00180208
R8812 VPWR.n1382 VPWR.n1381 0.00180208
R8813 VPWR.n1379 VPWR.n1378 0.00180208
R8814 VPWR VPWR.n3214 0.00180208
R8815 VPWR.n3445 VPWR.n1319 0.00180208
R8816 VPWR.n3443 VPWR.n3442 0.00180208
R8817 VPWR VPWR.n1388 0.00180208
R8818 VPWR.n1325 VPWR.n1324 0.00180208
R8819 VPWR.n1377 VPWR.n1330 0.00180208
R8820 VPWR.n3552 VPWR.n1282 0.00180208
R8821 VPWR.n3550 VPWR.n3549 0.00180208
R8822 VPWR.n3532 VPWR.n3531 0.00180208
R8823 VPWR.n3529 VPWR.n3528 0.00180208
R8824 VPWR VPWR 0.00180208
R8825 VPWR VPWR.n3775 0.00180208
R8826 VPWR VPWR 0.00180208
R8827 VPWR.n3554 VPWR.n3553 0.00180208
R8828 VPWR.n1286 VPWR.n1285 0.00180208
R8829 VPWR VPWR.n3538 0.00180208
R8830 VPWR.n3470 VPWR.n3469 0.00180208
R8831 VPWR.n3527 VPWR.n3474 0.00180208
R8832 VPWR.n4093 VPWR.n4092 0.00180208
R8833 VPWR.n1056 VPWR.n1055 0.00180208
R8834 VPWR.n981 VPWR.n980 0.00180208
R8835 VPWR.n1042 VPWR.n983 0.00180208
R8836 VPWR VPWR.n3874 0.00180208
R8837 VPWR VPWR 0.00180208
R8838 VPWR VPWR 0.00180208
R8839 VPWR.n4091 VPWR.n1052 0.00180208
R8840 VPWR.n4089 VPWR.n4088 0.00180208
R8841 VPWR.n986 VPWR.n985 0.00180208
R8842 VPWR.n1041 VPWR.n993 0.00180208
R8843 VPWR.n4341 VPWR.n757 0.00180208
R8844 VPWR.n4344 VPWR.n4343 0.00180208
R8845 VPWR.n4135 VPWR.n4134 0.00180208
R8846 VPWR.n4202 VPWR.n4137 0.00180208
R8847 VPWR VPWR.n4379 0.00180208
R8848 VPWR.n4340 VPWR.n4339 0.00180208
R8849 VPWR.n4355 VPWR.n4354 0.00180208
R8850 VPWR.n4140 VPWR.n4139 0.00180208
R8851 VPWR.n4201 VPWR.n4147 0.00180208
R8852 VPWR.n4808 VPWR.n4581 0.00180208
R8853 VPWR.n4811 VPWR.n4810 0.00180208
R8854 VPWR.n4503 VPWR.n4502 0.00180208
R8855 VPWR.n4565 VPWR.n4505 0.00180208
R8856 VPWR VPWR.n4910 0.00180208
R8857 VPWR VPWR 0.00180208
R8858 VPWR.n4807 VPWR.n4806 0.00180208
R8859 VPWR.n4823 VPWR.n4822 0.00180208
R8860 VPWR.n4508 VPWR.n4507 0.00180208
R8861 VPWR.n4564 VPWR.n4515 0.00180208
R8862 VPWR.n5278 VPWR.n5277 0.00180208
R8863 VPWR.n304 VPWR.n303 0.00180208
R8864 VPWR.n249 VPWR.n248 0.00180208
R8865 VPWR.n295 VPWR.n251 0.00180208
R8866 VPWR VPWR.n5032 0.00180208
R8867 VPWR VPWR 0.00180208
R8868 VPWR.n5276 VPWR.n300 0.00180208
R8869 VPWR.n5274 VPWR.n5273 0.00180208
R8870 VPWR.n254 VPWR.n253 0.00180208
R8871 VPWR.n294 VPWR.n260 0.00180208
R8872 VPWR.n5780 VPWR.n5768 0.00180208
R8873 VPWR.n5778 VPWR.n5777 0.00180208
R8874 VPWR.n5312 VPWR.n5311 0.00180208
R8875 VPWR.n5376 VPWR.n5314 0.00180208
R8876 VPWR VPWR.n5808 0.00180208
R8877 VPWR VPWR 0.00180208
R8878 VPWR.n5781 VPWR.n229 0.00180208
R8879 VPWR.n5784 VPWR.n5783 0.00180208
R8880 VPWR.n5317 VPWR.n5316 0.00180208
R8881 VPWR.n5375 VPWR.n5324 0.00180208
R8882 VPWR.n5560 VPWR.n5559 0.00180208
R8883 VPWR.n5392 VPWR.n5391 0.00180208
R8884 VPWR.n5678 VPWR.n5677 0.00180208
R8885 VPWR.n5742 VPWR.n5664 0.00180208
R8886 VPWR VPWR.n5949 0.00180208
R8887 VPWR.n5430 VPWR 0.00180208
R8888 VPWR.n5558 VPWR.n5381 0.00180208
R8889 VPWR.n5556 VPWR.n5382 0.00180208
R8890 VPWR.n5686 VPWR.n5685 0.00180208
R8891 VPWR.n5741 VPWR.n5689 0.00180208
R8892 VPWR.n2332 VPWR.n2212 0.00180208
R8893 VPWR.n2335 VPWR.n2334 0.00180208
R8894 VPWR.n2244 VPWR.n2243 0.00180208
R8895 VPWR.n2308 VPWR.n2251 0.00180208
R8896 VPWR.n2331 VPWR.n2319 0.00180208
R8897 VPWR.n2329 VPWR.n2328 0.00180208
R8898 VPWR.n2239 VPWR.n2238 0.00180208
R8899 VPWR.n2309 VPWR.n2241 0.00180208
R8900 VPWR.n6182 VPWR.n81 0.00180208
R8901 VPWR.n6185 VPWR.n6184 0.00180208
R8902 VPWR.n5584 VPWR.n5583 0.00180208
R8903 VPWR.n5641 VPWR.n5586 0.00180208
R8904 VPWR.n28 VPWR 0.00180208
R8905 VPWR VPWR 0.00180208
R8906 VPWR VPWR 0.00180208
R8907 VPWR.n6181 VPWR.n6178 0.00180208
R8908 VPWR.n6179 VPWR.n79 0.00180208
R8909 VPWR.n5589 VPWR.n5588 0.00180208
R8910 VPWR.n5640 VPWR.n5591 0.00180208
R8911 VPWR.n3055 VPWR.n3050 0.0014919
R8912 VPWR.n3050 VPWR.n3049 0.00140106
R8913 VPWR.n2928 VPWR.n1781 0.00140106
R8914 VPWR.n2928 VPWR.n2927 0.00140106
R8915 VPWR.n4387 VPWR.n699 0.00119134
R8916 VPWR.n4207 VPWR.n4110 0.00119134
R8917 VPWR.n4223 VPWR.n784 0.00119134
R8918 VGND.n225 VGND.n224 6.95552e+06
R8919 VGND.n226 VGND.n127 6.95552e+06
R8920 VGND.n5013 VGND.n231 6.95552e+06
R8921 VGND.n5014 VGND.n230 6.95552e+06
R8922 VGND.n5010 VGND.n233 6.95552e+06
R8923 VGND.n5011 VGND.n232 6.95552e+06
R8924 VGND.n5007 VGND.n235 6.95552e+06
R8925 VGND.n5008 VGND.n234 6.95552e+06
R8926 VGND.n5004 VGND.n237 6.95552e+06
R8927 VGND.n5005 VGND.n236 6.95552e+06
R8928 VGND.n5001 VGND.n239 6.95552e+06
R8929 VGND.n5002 VGND.n238 6.95552e+06
R8930 VGND.n4998 VGND.n241 6.95552e+06
R8931 VGND.n4999 VGND.n240 6.95552e+06
R8932 VGND.n4995 VGND.n243 6.95552e+06
R8933 VGND.n4996 VGND.n242 6.95552e+06
R8934 VGND.n4992 VGND.n245 6.95552e+06
R8935 VGND.n4993 VGND.n244 6.95552e+06
R8936 VGND.n4989 VGND.n247 6.95552e+06
R8937 VGND.n4990 VGND.n246 6.95552e+06
R8938 VGND.n5016 VGND.n229 6.95552e+06
R8939 VGND.n5017 VGND.n228 6.95552e+06
R8940 VGND.n4975 VGND.n4974 131565
R8941 VGND.n4988 VGND.n4987 68558.8
R8942 VGND.n5018 VGND.n127 40822.2
R8943 VGND.n5018 VGND.n5017 40822.2
R8944 VGND.n5016 VGND.n5015 40822.2
R8945 VGND.n5015 VGND.n5014 40822.2
R8946 VGND.n5013 VGND.n5012 40822.2
R8947 VGND.n5012 VGND.n5011 40822.2
R8948 VGND.n5010 VGND.n5009 40822.2
R8949 VGND.n5009 VGND.n5008 40822.2
R8950 VGND.n5007 VGND.n5006 40822.2
R8951 VGND.n5006 VGND.n5005 40822.2
R8952 VGND.n5004 VGND.n5003 40822.2
R8953 VGND.n5003 VGND.n5002 40822.2
R8954 VGND.n5001 VGND.n5000 40822.2
R8955 VGND.n5000 VGND.n4999 40822.2
R8956 VGND.n4998 VGND.n4997 40822.2
R8957 VGND.n4997 VGND.n4996 40822.2
R8958 VGND.n4995 VGND.n4994 40822.2
R8959 VGND.n4994 VGND.n4993 40822.2
R8960 VGND.n4992 VGND.n4991 40822.2
R8961 VGND.n4991 VGND.n4990 40822.2
R8962 VGND.n4989 VGND.n4988 40822.2
R8963 VGND.n224 VGND 19898.8
R8964 VGND VGND 12407.7
R8965 VGND VGND 11615.3
R8966 VGND VGND 8530.27
R8967 VGND.n225 VGND 8272.92
R8968 VGND VGND 7754.79
R8969 VGND VGND 7754.79
R8970 VGND VGND 7754.79
R8971 VGND VGND 7754.79
R8972 VGND VGND 7746.36
R8973 VGND.n307 VGND.n246 7652.17
R8974 VGND.n4974 VGND.n247 7652.17
R8975 VGND.n397 VGND.n244 7652.17
R8976 VGND.n307 VGND.n245 7652.17
R8977 VGND.n701 VGND.n242 7652.17
R8978 VGND.n397 VGND.n243 7652.17
R8979 VGND.n769 VGND.n240 7652.17
R8980 VGND.n701 VGND.n241 7652.17
R8981 VGND.n1050 VGND.n238 7652.17
R8982 VGND.n769 VGND.n239 7652.17
R8983 VGND.n1139 VGND.n236 7652.17
R8984 VGND.n1050 VGND.n237 7652.17
R8985 VGND.n1352 VGND.n234 7652.17
R8986 VGND.n1139 VGND.n235 7652.17
R8987 VGND.n2123 VGND.n232 7652.17
R8988 VGND.n1352 VGND.n233 7652.17
R8989 VGND.n228 VGND.n227 7652.17
R8990 VGND.n1533 VGND.n229 7652.17
R8991 VGND.n1533 VGND.n230 7652.17
R8992 VGND.n2123 VGND.n231 7652.17
R8993 VGND.n227 VGND.n226 7652.17
R8994 VGND.n224 VGND.n127 7007.41
R8995 VGND.n5017 VGND.n5016 7007.41
R8996 VGND.n5014 VGND.n5013 7007.41
R8997 VGND.n5011 VGND.n5010 7007.41
R8998 VGND.n5008 VGND.n5007 7007.41
R8999 VGND.n5005 VGND.n5004 7007.41
R9000 VGND.n5002 VGND.n5001 7007.41
R9001 VGND.n4999 VGND.n4998 7007.41
R9002 VGND.n4996 VGND.n4995 7007.41
R9003 VGND.n4993 VGND.n4992 7007.41
R9004 VGND.n4990 VGND.n4989 7007.41
R9005 VGND VGND 6515.71
R9006 VGND VGND 6220.69
R9007 VGND VGND 6203.83
R9008 VGND VGND 6203.83
R9009 VGND VGND 6203.83
R9010 VGND VGND 6203.83
R9011 VGND VGND 6203.83
R9012 VGND VGND 6203.83
R9013 VGND VGND 6195.4
R9014 VGND VGND 6195.4
R9015 VGND VGND 6195.4
R9016 VGND VGND 6195.4
R9017 VGND VGND 6195.4
R9018 VGND VGND 6195.4
R9019 VGND VGND 6195.4
R9020 VGND VGND 6195.4
R9021 VGND VGND 6195.4
R9022 VGND VGND 6195.4
R9023 VGND VGND 5731.8
R9024 VGND VGND 5445.21
R9025 VGND VGND 5445.21
R9026 VGND VGND 5436.78
R9027 VGND VGND 5428.35
R9028 VGND VGND 5428.35
R9029 VGND VGND 5428.35
R9030 VGND VGND 5428.35
R9031 VGND VGND 5428.35
R9032 VGND VGND 5428.35
R9033 VGND VGND 5428.35
R9034 VGND VGND 5428.35
R9035 VGND VGND 5428.35
R9036 VGND VGND 5428.35
R9037 VGND VGND 5411.49
R9038 VGND VGND 5403.07
R9039 VGND.n3200 VGND 4796.17
R9040 VGND VGND 4669.73
R9041 VGND VGND 4661.3
R9042 VGND VGND 4661.3
R9043 VGND VGND 4652.87
R9044 VGND VGND 4652.87
R9045 VGND VGND 4652.87
R9046 VGND VGND 4652.87
R9047 VGND VGND 4652.87
R9048 VGND VGND 4652.87
R9049 VGND VGND 4652.87
R9050 VGND VGND 4652.87
R9051 VGND VGND 4652.87
R9052 VGND VGND 4652.87
R9053 VGND VGND 4652.87
R9054 VGND VGND 4652.87
R9055 VGND VGND 4652.87
R9056 VGND VGND 4652.87
R9057 VGND VGND 4652.87
R9058 VGND VGND 4652.87
R9059 VGND VGND 4652.87
R9060 VGND VGND 4652.87
R9061 VGND VGND 4652.87
R9062 VGND VGND 4652.87
R9063 VGND VGND 4644.44
R9064 VGND VGND 4644.44
R9065 VGND VGND 4644.44
R9066 VGND VGND 4644.44
R9067 VGND VGND 4644.44
R9068 VGND VGND 4644.44
R9069 VGND VGND 4644.44
R9070 VGND VGND 4644.44
R9071 VGND VGND 4644.44
R9072 VGND VGND 4644.44
R9073 VGND VGND 4644.44
R9074 VGND VGND 4644.44
R9075 VGND VGND 4644.44
R9076 VGND VGND 4644.44
R9077 VGND VGND 4636.02
R9078 VGND VGND 4031.2
R9079 VGND VGND 3894.25
R9080 VGND VGND 3894.25
R9081 VGND VGND 3885.82
R9082 VGND VGND 3885.82
R9083 VGND VGND 3877.39
R9084 VGND VGND 3877.39
R9085 VGND VGND 3877.39
R9086 VGND VGND 3877.39
R9087 VGND VGND 3877.39
R9088 VGND VGND 3877.39
R9089 VGND VGND 3877.39
R9090 VGND VGND 3877.39
R9091 VGND VGND 3877.39
R9092 VGND VGND 3868.97
R9093 VGND VGND 3868.97
R9094 VGND VGND 3868.97
R9095 VGND VGND 3868.97
R9096 VGND VGND 3868.97
R9097 VGND VGND 3868.97
R9098 VGND VGND 3695.27
R9099 VGND VGND 3413.79
R9100 VGND VGND 3405.36
R9101 VGND VGND.n4588 3245.21
R9102 VGND.n4589 VGND 3245.21
R9103 VGND VGND.n4747 3245.21
R9104 VGND.n4748 VGND 3245.21
R9105 VGND VGND.n484 3245.21
R9106 VGND.n4092 VGND 3245.21
R9107 VGND.n702 VGND 3245.21
R9108 VGND VGND.n884 3245.21
R9109 VGND.n3575 VGND 3245.21
R9110 VGND VGND.n3199 3245.21
R9111 VGND VGND.n3348 3245.21
R9112 VGND VGND.n1241 3245.21
R9113 VGND VGND.n1249 3245.21
R9114 VGND.n2946 VGND 3245.21
R9115 VGND VGND.n2734 3245.21
R9116 VGND.n2408 VGND 3245.21
R9117 VGND.n2018 VGND 3245.21
R9118 VGND.n2017 VGND 3245.21
R9119 VGND.n4971 VGND 3245.21
R9120 VGND.n4968 VGND 3245.21
R9121 VGND.n4967 VGND 3245.21
R9122 VGND.n222 VGND 3245.21
R9123 VGND.n5020 VGND 3245.21
R9124 VGND.n5019 VGND 3245.21
R9125 VGND VGND 3118.77
R9126 VGND VGND 3118.77
R9127 VGND VGND 3118.77
R9128 VGND VGND 3110.34
R9129 VGND VGND 3110.34
R9130 VGND VGND 3110.34
R9131 VGND VGND 3110.34
R9132 VGND VGND 3110.34
R9133 VGND VGND 3110.34
R9134 VGND VGND 3110.34
R9135 VGND VGND 3110.34
R9136 VGND VGND 3110.34
R9137 VGND VGND 3110.34
R9138 VGND VGND 3110.34
R9139 VGND VGND 3110.34
R9140 VGND VGND 3110.34
R9141 VGND VGND 3110.34
R9142 VGND VGND 3101.92
R9143 VGND VGND 3101.92
R9144 VGND VGND 3101.92
R9145 VGND VGND 3101.92
R9146 VGND VGND 3101.92
R9147 VGND VGND 3101.92
R9148 VGND VGND 3101.92
R9149 VGND VGND 3101.92
R9150 VGND VGND 3101.92
R9151 VGND VGND 3101.92
R9152 VGND VGND 3101.92
R9153 VGND VGND 3101.92
R9154 VGND VGND 3101.92
R9155 VGND VGND 3101.92
R9156 VGND VGND 3101.92
R9157 VGND VGND 3101.92
R9158 VGND VGND 3101.92
R9159 VGND VGND 3101.92
R9160 VGND VGND 3101.92
R9161 VGND VGND 3101.92
R9162 VGND VGND 3101.92
R9163 VGND VGND 3101.92
R9164 VGND VGND 3101.92
R9165 VGND VGND 3101.92
R9166 VGND VGND 3101.92
R9167 VGND VGND 3101.92
R9168 VGND VGND 3101.92
R9169 VGND VGND 3101.92
R9170 VGND VGND 3101.92
R9171 VGND VGND 3101.92
R9172 VGND VGND 3101.92
R9173 VGND VGND 3101.92
R9174 VGND VGND 3101.92
R9175 VGND VGND 3101.92
R9176 VGND VGND 3101.92
R9177 VGND VGND 3101.92
R9178 VGND VGND 3101.92
R9179 VGND VGND 3101.92
R9180 VGND VGND 3101.92
R9181 VGND VGND 3101.92
R9182 VGND VGND 3101.92
R9183 VGND VGND 3101.92
R9184 VGND VGND 3101.92
R9185 VGND VGND 3101.92
R9186 VGND VGND 3101.92
R9187 VGND VGND 3101.92
R9188 VGND VGND 3101.92
R9189 VGND VGND 3101.92
R9190 VGND VGND 3101.92
R9191 VGND VGND 3101.92
R9192 VGND VGND 3101.92
R9193 VGND VGND 3101.92
R9194 VGND VGND 3101.92
R9195 VGND VGND 3101.92
R9196 VGND VGND 3101.92
R9197 VGND VGND 3101.92
R9198 VGND VGND 3101.92
R9199 VGND VGND 3101.92
R9200 VGND VGND 3101.92
R9201 VGND VGND 3093.49
R9202 VGND VGND 3093.49
R9203 VGND VGND 3093.49
R9204 VGND VGND 3093.49
R9205 VGND VGND 3093.49
R9206 VGND VGND 3093.49
R9207 VGND VGND 3093.49
R9208 VGND VGND 3093.49
R9209 VGND VGND 3093.49
R9210 VGND VGND 3093.49
R9211 VGND VGND 3093.49
R9212 VGND VGND 3093.49
R9213 VGND VGND 3093.49
R9214 VGND VGND 3093.49
R9215 VGND VGND 3093.49
R9216 VGND VGND 3085.06
R9217 VGND VGND 3023.4
R9218 VGND VGND 2975.48
R9219 VGND VGND 2950.19
R9220 VGND VGND.n3885 2781.61
R9221 VGND.n5568 VGND 2749.54
R9222 VGND.n247 VGND.n246 2742.03
R9223 VGND.n245 VGND.n244 2742.03
R9224 VGND.n243 VGND.n242 2742.03
R9225 VGND.n241 VGND.n240 2742.03
R9226 VGND.n239 VGND.n238 2742.03
R9227 VGND.n237 VGND.n236 2742.03
R9228 VGND.n235 VGND.n234 2742.03
R9229 VGND.n233 VGND.n232 2742.03
R9230 VGND.n229 VGND.n228 2742.03
R9231 VGND.n231 VGND.n230 2742.03
R9232 VGND.n226 VGND.n225 2742.03
R9233 VGND VGND 2683.82
R9234 VGND VGND 2683.82
R9235 VGND VGND 2638.31
R9236 VGND VGND 2638.31
R9237 VGND VGND.n494 2469.73
R9238 VGND.n3574 VGND 2469.73
R9239 VGND VGND.n1248 2469.73
R9240 VGND.n2646 VGND 2469.73
R9241 VGND.n2735 VGND 2469.73
R9242 VGND VGND 2351.54
R9243 VGND VGND 2351.54
R9244 VGND VGND 2351.54
R9245 VGND VGND 2351.54
R9246 VGND VGND 2351.54
R9247 VGND VGND 2343.29
R9248 VGND VGND 2343.29
R9249 VGND VGND 2334.87
R9250 VGND VGND 2334.87
R9251 VGND VGND 2334.87
R9252 VGND VGND 2334.87
R9253 VGND VGND 2334.87
R9254 VGND VGND 2334.87
R9255 VGND VGND 2334.87
R9256 VGND VGND 2334.87
R9257 VGND VGND 2326.44
R9258 VGND VGND 2326.44
R9259 VGND VGND 2326.44
R9260 VGND VGND 2326.44
R9261 VGND VGND 2326.44
R9262 VGND VGND 2326.44
R9263 VGND VGND 2326.44
R9264 VGND VGND 2326.44
R9265 VGND VGND 2326.44
R9266 VGND VGND 2326.44
R9267 VGND VGND 2326.44
R9268 VGND VGND 2326.44
R9269 VGND VGND 2326.44
R9270 VGND VGND 2326.44
R9271 VGND VGND 2326.44
R9272 VGND VGND 2326.44
R9273 VGND VGND 2326.44
R9274 VGND VGND 2326.44
R9275 VGND VGND 2326.44
R9276 VGND VGND 2326.44
R9277 VGND VGND 2326.44
R9278 VGND VGND 2326.44
R9279 VGND VGND 2326.44
R9280 VGND VGND 2326.44
R9281 VGND VGND 2326.44
R9282 VGND VGND 2326.44
R9283 VGND VGND 2326.44
R9284 VGND VGND 2326.44
R9285 VGND VGND 2326.44
R9286 VGND VGND 2326.44
R9287 VGND VGND 2326.44
R9288 VGND VGND 2326.44
R9289 VGND VGND 2326.44
R9290 VGND VGND 2326.44
R9291 VGND VGND 2326.44
R9292 VGND VGND 2326.44
R9293 VGND VGND 2326.44
R9294 VGND VGND 2326.44
R9295 VGND VGND 2326.44
R9296 VGND VGND 2326.44
R9297 VGND VGND 2326.44
R9298 VGND VGND 2326.44
R9299 VGND VGND 2326.44
R9300 VGND VGND 2326.44
R9301 VGND VGND 2326.44
R9302 VGND VGND 2326.44
R9303 VGND VGND 2326.44
R9304 VGND VGND 2326.44
R9305 VGND VGND 2326.44
R9306 VGND VGND 2326.44
R9307 VGND VGND 2326.44
R9308 VGND VGND 2326.44
R9309 VGND VGND 2326.44
R9310 VGND VGND 2326.44
R9311 VGND VGND 2326.44
R9312 VGND VGND 2326.44
R9313 VGND VGND 2326.44
R9314 VGND VGND 2326.44
R9315 VGND VGND 2326.44
R9316 VGND VGND 2326.44
R9317 VGND VGND 2318.01
R9318 VGND VGND 2318.01
R9319 VGND VGND 2318.01
R9320 VGND VGND 2318.01
R9321 VGND VGND 2318.01
R9322 VGND VGND 2318.01
R9323 VGND VGND 2318.01
R9324 VGND VGND 2318.01
R9325 VGND VGND 2318.01
R9326 VGND VGND 2318.01
R9327 VGND VGND 2318.01
R9328 VGND VGND 2318.01
R9329 VGND VGND 2318.01
R9330 VGND VGND 2318.01
R9331 VGND VGND 2318.01
R9332 VGND VGND 2318.01
R9333 VGND VGND 2318.01
R9334 VGND VGND 2309.58
R9335 VGND VGND 2309.58
R9336 VGND VGND 2309.58
R9337 VGND VGND 2309.58
R9338 VGND VGND 2309.58
R9339 VGND VGND 2309.58
R9340 VGND VGND 2309.58
R9341 VGND VGND 2309.58
R9342 VGND VGND 2015.6
R9343 VGND VGND 2015.6
R9344 VGND VGND 2015.6
R9345 VGND VGND 2014.56
R9346 VGND VGND 1997.7
R9347 VGND.n3800 VGND 1694.25
R9348 VGND.n4972 VGND 1694.25
R9349 VGND VGND 1679.67
R9350 VGND.n1041 VGND 1677.39
R9351 VGND.n1353 VGND 1677.39
R9352 VGND VGND.n1641 1677.39
R9353 VGND VGND 1567.82
R9354 VGND VGND 1567.82
R9355 VGND VGND 1567.82
R9356 VGND VGND 1559.39
R9357 VGND VGND 1559.39
R9358 VGND VGND 1559.39
R9359 VGND VGND 1559.39
R9360 VGND VGND 1559.39
R9361 VGND VGND 1559.39
R9362 VGND VGND 1550.96
R9363 VGND VGND 1550.96
R9364 VGND VGND 1550.96
R9365 VGND VGND 1550.96
R9366 VGND VGND 1550.96
R9367 VGND VGND 1550.96
R9368 VGND VGND 1550.96
R9369 VGND VGND 1550.96
R9370 VGND VGND 1550.96
R9371 VGND VGND 1550.96
R9372 VGND VGND 1550.96
R9373 VGND VGND 1550.96
R9374 VGND VGND 1550.96
R9375 VGND VGND 1550.96
R9376 VGND VGND 1550.96
R9377 VGND VGND.n2645 1550.96
R9378 VGND VGND 1550.96
R9379 VGND VGND 1550.96
R9380 VGND VGND 1550.96
R9381 VGND VGND 1550.96
R9382 VGND VGND 1550.96
R9383 VGND VGND 1550.96
R9384 VGND VGND 1550.96
R9385 VGND VGND 1550.96
R9386 VGND VGND 1550.96
R9387 VGND VGND 1550.96
R9388 VGND VGND 1550.96
R9389 VGND VGND 1550.96
R9390 VGND VGND 1550.96
R9391 VGND VGND 1542.53
R9392 VGND VGND 1542.53
R9393 VGND VGND 1542.53
R9394 VGND VGND 1542.53
R9395 VGND VGND 1542.53
R9396 VGND VGND 1542.53
R9397 VGND VGND 1542.53
R9398 VGND VGND 1542.53
R9399 VGND VGND 1542.53
R9400 VGND VGND 1542.53
R9401 VGND VGND 1542.53
R9402 VGND VGND 1542.53
R9403 VGND VGND 1542.53
R9404 VGND VGND 1542.53
R9405 VGND VGND 1534.1
R9406 VGND VGND 1534.1
R9407 VGND VGND 1534.1
R9408 VGND VGND 1534.1
R9409 VGND VGND 1534.1
R9410 VGND VGND 1534.1
R9411 VGND VGND 1534.1
R9412 VGND VGND 1525.67
R9413 VGND VGND.n307 1432.95
R9414 VGND VGND.n397 1432.95
R9415 VGND VGND.n701 1432.95
R9416 VGND VGND.n769 1432.95
R9417 VGND VGND.n1050 1432.95
R9418 VGND VGND.n1139 1432.95
R9419 VGND VGND.n1352 1432.95
R9420 VGND VGND.n2123 1432.95
R9421 VGND VGND.n1533 1432.95
R9422 VGND.n4974 VGND 1432.95
R9423 VGND.n227 VGND 1432.95
R9424 VGND.n5572 VGND 1405.81
R9425 VGND.n5569 VGND 1405.81
R9426 VGND VGND 1343.73
R9427 VGND VGND 1343.73
R9428 VGND VGND 1343.73
R9429 VGND VGND 1343.73
R9430 VGND VGND 1343.73
R9431 VGND VGND 1343.73
R9432 VGND VGND 1343.73
R9433 VGND VGND 1239.08
R9434 VGND VGND 1239.08
R9435 VGND VGND 1239.08
R9436 VGND VGND 1007.8
R9437 VGND VGND 1007.8
R9438 VGND.n4269 VGND.n4266 990.732
R9439 VGND.n302 VGND 927.203
R9440 VGND VGND.n877 927.203
R9441 VGND VGND.n2407 927.203
R9442 VGND VGND.n1634 927.203
R9443 VGND.n4969 VGND 927.203
R9444 VGND.n223 VGND 927.203
R9445 VGND.n4093 VGND 918.774
R9446 VGND.n3886 VGND 918.774
R9447 VGND.n3573 VGND 918.774
R9448 VGND VGND.n2224 918.774
R9449 VGND.n2225 VGND 918.774
R9450 VGND.n1486 VGND 918.774
R9451 VGND.n4973 VGND 918.774
R9452 VGND.n2947 VGND 910.346
R9453 VGND VGND 800.766
R9454 VGND VGND 800.766
R9455 VGND VGND 792.337
R9456 VGND VGND 792.337
R9457 VGND VGND 792.337
R9458 VGND VGND 792.337
R9459 VGND VGND 792.337
R9460 VGND VGND 792.337
R9461 VGND VGND 792.337
R9462 VGND VGND 792.337
R9463 VGND VGND 783.909
R9464 VGND VGND 783.909
R9465 VGND VGND 783.909
R9466 VGND VGND 783.909
R9467 VGND VGND 783.909
R9468 VGND VGND 783.909
R9469 VGND VGND 783.909
R9470 VGND VGND 783.909
R9471 VGND VGND 783.909
R9472 VGND VGND 783.909
R9473 VGND VGND 783.909
R9474 VGND VGND 783.909
R9475 VGND VGND 783.909
R9476 VGND VGND 783.909
R9477 VGND VGND 783.909
R9478 VGND VGND 783.909
R9479 VGND VGND 783.909
R9480 VGND VGND 783.909
R9481 VGND VGND 783.909
R9482 VGND VGND 783.909
R9483 VGND VGND 783.909
R9484 VGND VGND 783.909
R9485 VGND VGND 783.909
R9486 VGND VGND 783.909
R9487 VGND VGND 783.909
R9488 VGND VGND 783.909
R9489 VGND VGND 783.909
R9490 VGND VGND 783.909
R9491 VGND VGND 783.909
R9492 VGND VGND 783.909
R9493 VGND VGND 783.909
R9494 VGND VGND 783.909
R9495 VGND VGND 783.909
R9496 VGND VGND 783.909
R9497 VGND VGND 783.909
R9498 VGND VGND 783.909
R9499 VGND VGND 783.909
R9500 VGND VGND 783.909
R9501 VGND VGND 783.909
R9502 VGND VGND 783.909
R9503 VGND VGND 783.909
R9504 VGND VGND 783.909
R9505 VGND VGND 783.909
R9506 VGND VGND 783.909
R9507 VGND VGND 783.909
R9508 VGND VGND 783.909
R9509 VGND VGND 783.909
R9510 VGND.n4979 VGND.n4978 782.61
R9511 VGND VGND 775.48
R9512 VGND VGND 775.48
R9513 VGND VGND 775.48
R9514 VGND VGND 775.48
R9515 VGND VGND 775.48
R9516 VGND VGND 775.48
R9517 VGND VGND 775.48
R9518 VGND VGND 775.48
R9519 VGND VGND 775.48
R9520 VGND VGND 775.48
R9521 VGND VGND 775.48
R9522 VGND VGND 775.48
R9523 VGND VGND 775.48
R9524 VGND VGND 775.48
R9525 VGND VGND 775.48
R9526 VGND VGND 775.48
R9527 VGND VGND 775.48
R9528 VGND VGND 775.48
R9529 VGND VGND 775.48
R9530 VGND VGND 775.48
R9531 VGND VGND 775.48
R9532 VGND VGND 775.48
R9533 VGND VGND 775.48
R9534 VGND VGND 775.48
R9535 VGND VGND 775.48
R9536 VGND VGND 775.48
R9537 VGND VGND 775.48
R9538 VGND VGND 775.48
R9539 VGND VGND 775.48
R9540 VGND VGND 775.48
R9541 VGND VGND 775.48
R9542 VGND VGND 775.48
R9543 VGND VGND 775.48
R9544 VGND VGND 775.48
R9545 VGND VGND 775.48
R9546 VGND VGND 775.48
R9547 VGND VGND 775.48
R9548 VGND VGND 775.48
R9549 VGND VGND 775.48
R9550 VGND VGND 775.48
R9551 VGND VGND 775.48
R9552 VGND VGND 775.48
R9553 VGND VGND 775.48
R9554 VGND VGND 775.48
R9555 VGND VGND 775.48
R9556 VGND VGND 775.48
R9557 VGND VGND 775.48
R9558 VGND VGND 775.48
R9559 VGND VGND 775.48
R9560 VGND VGND 775.48
R9561 VGND VGND 775.48
R9562 VGND VGND 775.48
R9563 VGND VGND 775.48
R9564 VGND VGND 775.48
R9565 VGND VGND 775.48
R9566 VGND VGND 775.48
R9567 VGND VGND 775.48
R9568 VGND VGND 775.48
R9569 VGND VGND 775.48
R9570 VGND VGND 775.48
R9571 VGND VGND 775.48
R9572 VGND VGND 775.48
R9573 VGND VGND 775.48
R9574 VGND VGND 775.48
R9575 VGND VGND 775.48
R9576 VGND VGND 775.48
R9577 VGND VGND 775.48
R9578 VGND VGND 775.48
R9579 VGND VGND 775.48
R9580 VGND VGND 775.48
R9581 VGND VGND 775.48
R9582 VGND VGND 775.48
R9583 VGND VGND 775.48
R9584 VGND VGND 775.48
R9585 VGND VGND 775.48
R9586 VGND VGND 775.48
R9587 VGND VGND 775.48
R9588 VGND VGND 775.48
R9589 VGND VGND 775.48
R9590 VGND VGND 775.48
R9591 VGND VGND 775.48
R9592 VGND VGND 775.48
R9593 VGND VGND 775.48
R9594 VGND VGND 775.48
R9595 VGND VGND 775.48
R9596 VGND VGND 775.48
R9597 VGND VGND 775.48
R9598 VGND VGND 775.48
R9599 VGND VGND 775.48
R9600 VGND VGND 775.48
R9601 VGND VGND 775.48
R9602 VGND VGND 775.48
R9603 VGND VGND 775.48
R9604 VGND VGND 775.48
R9605 VGND VGND 775.48
R9606 VGND VGND 775.48
R9607 VGND VGND 775.48
R9608 VGND VGND 775.48
R9609 VGND VGND 775.48
R9610 VGND VGND 775.48
R9611 VGND VGND 775.48
R9612 VGND VGND 775.48
R9613 VGND VGND 775.48
R9614 VGND VGND 775.48
R9615 VGND VGND 775.48
R9616 VGND VGND 775.48
R9617 VGND VGND 767.051
R9618 VGND VGND 767.051
R9619 VGND VGND 767.051
R9620 VGND VGND 767.051
R9621 VGND VGND 767.051
R9622 VGND VGND 767.051
R9623 VGND VGND 767.051
R9624 VGND VGND 767.051
R9625 VGND VGND 767.051
R9626 VGND VGND 767.051
R9627 VGND VGND 767.051
R9628 VGND VGND 767.051
R9629 VGND VGND 767.051
R9630 VGND VGND 767.051
R9631 VGND VGND 767.051
R9632 VGND VGND 767.051
R9633 VGND VGND 767.051
R9634 VGND VGND 767.051
R9635 VGND VGND 767.051
R9636 VGND VGND 767.051
R9637 VGND.n4985 VGND.n4984 765.217
R9638 VGND VGND 758.621
R9639 VGND VGND 758.621
R9640 VGND VGND 758.621
R9641 VGND VGND 750.192
R9642 VGND VGND 750.192
R9643 VGND.n4976 VGND.n4975 730.436
R9644 VGND.n4980 VGND.n4979 730.436
R9645 VGND.n4978 VGND.n4977 652.174
R9646 VGND.n4977 VGND.n4976 643.479
R9647 VGND.n4588 VGND 632.184
R9648 VGND.n4589 VGND 632.184
R9649 VGND VGND.n302 632.184
R9650 VGND.n4747 VGND 632.184
R9651 VGND.n4748 VGND 632.184
R9652 VGND.n484 VGND 632.184
R9653 VGND.n494 VGND 632.184
R9654 VGND.n4093 VGND 632.184
R9655 VGND VGND.n4092 632.184
R9656 VGND VGND.n4091 632.184
R9657 VGND.n702 VGND 632.184
R9658 VGND.n3799 VGND 632.184
R9659 VGND.n3800 VGND 632.184
R9660 VGND.n3885 VGND 632.184
R9661 VGND.n3886 VGND 632.184
R9662 VGND.n877 VGND 632.184
R9663 VGND.n884 VGND 632.184
R9664 VGND.n3575 VGND 632.184
R9665 VGND VGND.n3574 632.184
R9666 VGND VGND.n3573 632.184
R9667 VGND.n3199 VGND 632.184
R9668 VGND.n3200 VGND 632.184
R9669 VGND VGND.n1041 632.184
R9670 VGND.n3348 VGND 632.184
R9671 VGND.n3349 VGND 632.184
R9672 VGND.n1241 VGND 632.184
R9673 VGND.n1248 VGND 632.184
R9674 VGND.n1249 VGND 632.184
R9675 VGND.n2947 VGND 632.184
R9676 VGND.n1353 VGND 632.184
R9677 VGND.n2645 VGND 632.184
R9678 VGND.n2646 VGND 632.184
R9679 VGND.n2734 VGND 632.184
R9680 VGND.n2735 VGND 632.184
R9681 VGND.n2224 VGND 632.184
R9682 VGND.n2225 VGND 632.184
R9683 VGND VGND.n1486 632.184
R9684 VGND.n2407 VGND 632.184
R9685 VGND.n2408 VGND 632.184
R9686 VGND.n1634 VGND 632.184
R9687 VGND.n1641 VGND 632.184
R9688 VGND.n2018 VGND 632.184
R9689 VGND VGND.n2017 632.184
R9690 VGND.n1705 VGND 632.184
R9691 VGND VGND.n4973 632.184
R9692 VGND VGND.n4972 632.184
R9693 VGND VGND.n4971 632.184
R9694 VGND VGND.n4970 632.184
R9695 VGND VGND.n4969 632.184
R9696 VGND VGND.n4968 632.184
R9697 VGND VGND.n4967 632.184
R9698 VGND VGND.n223 632.184
R9699 VGND VGND.n222 632.184
R9700 VGND VGND.n221 632.184
R9701 VGND.n5020 VGND 632.184
R9702 VGND VGND.n5019 632.184
R9703 VGND VGND 623.755
R9704 VGND VGND.n2946 623.755
R9705 VGND.n4981 VGND.n4980 617.391
R9706 VGND.n5573 VGND.n5572 613.249
R9707 VGND.n5571 VGND.n27 613.249
R9708 VGND.n5570 VGND.n28 613.249
R9709 VGND.n5569 VGND.n29 613.249
R9710 VGND.n4971 VGND.n250 613.249
R9711 VGND.n1641 VGND.n1640 613.249
R9712 VGND.n2019 VGND.n2018 613.249
R9713 VGND.n4590 VGND.n4589 613.249
R9714 VGND.n4747 VGND.n4746 613.249
R9715 VGND.n4804 VGND.n4748 613.249
R9716 VGND.n4092 VGND.n495 613.249
R9717 VGND.n3885 VGND.n3884 613.249
R9718 VGND.n703 VGND.n702 613.249
R9719 VGND.n884 VGND.n883 613.249
R9720 VGND.n877 VGND.n876 613.249
R9721 VGND.n3348 VGND.n3347 613.249
R9722 VGND.n3268 VGND.n1041 613.249
R9723 VGND.n3199 VGND.n3198 613.249
R9724 VGND.n2948 VGND.n2947 613.249
R9725 VGND.n3014 VGND.n1249 613.249
R9726 VGND.n1241 VGND.n1240 613.249
R9727 VGND.n2645 VGND.n2644 613.249
R9728 VGND.n2734 VGND.n2733 613.249
R9729 VGND.n1404 VGND.n1353 613.249
R9730 VGND.n2407 VGND.n2406 613.249
R9731 VGND.n2017 VGND.n2016 613.249
R9732 VGND.n5021 VGND.n5020 613.249
R9733 VGND.n5019 VGND.n126 613.249
R9734 VGND.n5568 VGND.n5567 613.249
R9735 VGND.n4970 VGND.n251 611.862
R9736 VGND.n1706 VGND.n1705 611.862
R9737 VGND.n4091 VGND.n4090 611.862
R9738 VGND.n3799 VGND.n3798 611.862
R9739 VGND.n3574 VGND.n885 611.862
R9740 VGND.n3350 VGND.n3349 611.862
R9741 VGND.n2946 VGND.n2945 611.862
R9742 VGND.n2648 VGND.n2646 611.862
R9743 VGND.n2787 VGND.n2735 611.862
R9744 VGND.n221 VGND.n107 611.862
R9745 VGND.n4973 VGND.n248 611.225
R9746 VGND.n4095 VGND.n4093 611.225
R9747 VGND.n3933 VGND.n3886 611.225
R9748 VGND.n3573 VGND.n3572 611.225
R9749 VGND.n1248 VGND.n1247 611.225
R9750 VGND.n2226 VGND.n2225 611.225
R9751 VGND.n2224 VGND.n2223 611.225
R9752 VGND.n4972 VGND.n249 611.211
R9753 VGND.n1634 VGND.n1633 610.78
R9754 VGND.n4662 VGND.n302 610.679
R9755 VGND.n2317 VGND.n1486 610.679
R9756 VGND.n4968 VGND.n253 609.497
R9757 VGND.n4588 VGND.n4587 609.497
R9758 VGND.n494 VGND.n493 609.497
R9759 VGND.n484 VGND.n483 609.497
R9760 VGND.n3801 VGND.n3800 609.497
R9761 VGND.n3576 VGND.n3575 609.497
R9762 VGND.n3201 VGND.n3200 609.497
R9763 VGND.n2469 VGND.n2408 609.497
R9764 VGND.n222 VGND.n220 609.497
R9765 VGND.n4969 VGND.n252 609.497
R9766 VGND.n223 VGND.n211 609.497
R9767 VGND.n4982 VGND.n4981 608.697
R9768 VGND.n4984 VGND.n4983 600
R9769 VGND.n4986 VGND.n4985 582.61
R9770 VGND.n4983 VGND.n4982 565.217
R9771 VGND.n4991 VGND 564.751
R9772 VGND.n4994 VGND 564.751
R9773 VGND.n4997 VGND 564.751
R9774 VGND.n5000 VGND 564.751
R9775 VGND.n5003 VGND 564.751
R9776 VGND.n5006 VGND 564.751
R9777 VGND.n5009 VGND 564.751
R9778 VGND.n5012 VGND 564.751
R9779 VGND.n5015 VGND 564.751
R9780 VGND.n4988 VGND 564.751
R9781 VGND VGND.n5018 564.751
R9782 VGND VGND 463.603
R9783 VGND VGND 463.603
R9784 VGND.n5571 VGND 401.661
R9785 VGND.n5570 VGND 401.661
R9786 VGND VGND 335.935
R9787 VGND VGND 335.935
R9788 VGND VGND 335.935
R9789 VGND VGND 335.935
R9790 VGND VGND 335.935
R9791 VGND VGND 335.935
R9792 VGND VGND 335.935
R9793 VGND.n4967 VGND.n4966 306.625
R9794 VGND.n5572 VGND 273.86
R9795 VGND VGND.n5571 273.86
R9796 VGND VGND.n5570 273.86
R9797 VGND VGND.n5569 273.86
R9798 VGND VGND.n5568 273.86
R9799 VGND.n4987 VGND.n4986 208.696
R9800 VGND.n4928 VGND.t81 191.915
R9801 VGND.n4928 VGND.t62 191.915
R9802 VGND.n4927 VGND.t55 191.915
R9803 VGND.n4223 VGND.t88 191.915
R9804 VGND.n4223 VGND.t73 191.915
R9805 VGND.n1663 VGND.t335 191.915
R9806 VGND.n1663 VGND.t316 191.915
R9807 VGND.n1594 VGND.t352 191.915
R9808 VGND.n1594 VGND.t325 191.915
R9809 VGND.n4760 VGND.t121 191.915
R9810 VGND.n4760 VGND.t98 191.915
R9811 VGND.n316 VGND.t131 191.915
R9812 VGND.n316 VGND.t108 191.915
R9813 VGND.n4049 VGND.t262 191.915
R9814 VGND.n4049 VGND.t146 191.915
R9815 VGND.n405 VGND.t279 191.915
R9816 VGND.n405 VGND.t163 191.915
R9817 VGND.n3897 VGND.t318 191.915
R9818 VGND.n3897 VGND.t287 191.915
R9819 VGND.n676 VGND.t327 191.915
R9820 VGND.n676 VGND.t304 191.915
R9821 VGND.n839 VGND.t379 191.915
R9822 VGND.n839 VGND.t351 191.915
R9823 VGND.n3524 VGND.t369 191.915
R9824 VGND.n3524 VGND.t339 191.915
R9825 VGND.n3359 VGND.t278 191.915
R9826 VGND.n3359 VGND.t247 191.915
R9827 VGND.n3358 VGND.t231 191.915
R9828 VGND.n1056 VGND.t291 191.915
R9829 VGND.n1056 VGND.t263 191.915
R9830 VGND.n2909 VGND.t326 191.915
R9831 VGND.n2909 VGND.t303 191.915
R9832 VGND.n1151 VGND.t336 191.915
R9833 VGND.n1151 VGND.t317 191.915
R9834 VGND.n2744 VGND.t234 191.915
R9835 VGND.n2744 VGND.t350 191.915
R9836 VGND.n2743 VGND.t179 191.915
R9837 VGND.n1367 VGND.t246 191.915
R9838 VGND.n1367 VGND.t368 191.915
R9839 VGND.n2425 VGND.t290 191.915
R9840 VGND.n2425 VGND.t261 191.915
R9841 VGND.n2133 VGND.t302 191.915
R9842 VGND.n2133 VGND.t277 191.915
R9843 VGND.n1888 VGND.t245 191.915
R9844 VGND.n1888 VGND.t224 191.915
R9845 VGND.n137 VGND.t260 191.915
R9846 VGND.n137 VGND.t233 191.915
R9847 VGND.n1592 VGND.t202 190.931
R9848 VGND.n142 VGND.t212 188.97
R9849 VGND.n2 VGND.t288 183.082
R9850 VGND.n3522 VGND.t305 183.082
R9851 VGND.n5517 VGND.t276 183.082
R9852 VGND.n4094 VGND.t84 153.644
R9853 VGND.n3932 VGND.t59 153.644
R9854 VGND.n886 VGND.t323 153.644
R9855 VGND.n2257 VGND.t319 153.644
R9856 VGND.n4882 VGND.t362 150.329
R9857 VGND.n4409 VGND.t314 150.329
R9858 VGND.n1606 VGND.t69 150.329
R9859 VGND.n363 VGND.t345 150.329
R9860 VGND.n4751 VGND.t248 150.329
R9861 VGND.n502 VGND.t198 150.329
R9862 VGND.n440 VGND.t28 150.329
R9863 VGND.n395 VGND.t223 150.329
R9864 VGND.n4005 VGND.t92 150.329
R9865 VGND.n518 VGND.t180 150.329
R9866 VGND.n634 VGND.t89 150.329
R9867 VGND.n644 VGND.t338 150.329
R9868 VGND.n3512 VGND.t363 150.329
R9869 VGND.n1043 VGND.t358 150.329
R9870 VGND.n1071 VGND.t382 150.329
R9871 VGND.n1097 VGND.t359 150.329
R9872 VGND.n1271 VGND.t26 150.329
R9873 VGND.n1364 VGND.t120 150.329
R9874 VGND.n2823 VGND.t232 150.329
R9875 VGND.n1488 VGND.t256 150.329
R9876 VGND.n2128 VGND.t306 150.329
R9877 VGND.n4215 VGND.t206 150.204
R9878 VGND.n1582 VGND.t162 148.918
R9879 VGND.n254 VGND.t138 148.862
R9880 VGND.n254 VGND.t17 148.862
R9881 VGND.n255 VGND.t79 148.862
R9882 VGND.n255 VGND.t333 148.862
R9883 VGND.n4226 VGND.t103 148.862
R9884 VGND.n4226 VGND.t215 148.862
R9885 VGND.n4207 VGND.t186 148.862
R9886 VGND.n4207 VGND.t313 148.862
R9887 VGND.n1662 VGND.t282 148.862
R9888 VGND.n1597 VGND.t38 148.862
R9889 VGND.n1597 VGND.t161 148.862
R9890 VGND.n1630 VGND.t104 148.862
R9891 VGND.n319 VGND.t241 148.862
R9892 VGND.n319 VGND.t385 148.862
R9893 VGND.n4568 VGND.t85 148.862
R9894 VGND.n4681 VGND.t329 148.862
R9895 VGND.n4681 VGND.t189 148.862
R9896 VGND.n4052 VGND.t383 148.862
R9897 VGND.n408 VGND.t137 148.862
R9898 VGND.n402 VGND.t35 148.862
R9899 VGND.n447 VGND.t83 148.862
R9900 VGND.n447 VGND.t194 148.862
R9901 VGND.n3896 VGND.t342 148.862
R9902 VGND.n3896 VGND.t169 148.862
R9903 VGND.n651 VGND.t193 148.862
R9904 VGND.n687 VGND.t182 148.862
R9905 VGND.n687 VGND.t309 148.862
R9906 VGND.n842 VGND.t321 148.862
R9907 VGND.n842 VGND.t50 148.862
R9908 VGND.n1051 VGND.t221 148.862
R9909 VGND.n3406 VGND.t217 148.862
R9910 VGND.n2895 VGND.t173 148.862
R9911 VGND.n1328 VGND.t70 148.862
R9912 VGND.n1347 VGND.t251 148.862
R9913 VGND.n2173 VGND.t87 148.862
R9914 VGND.n259 VGND.t78 148.846
R9915 VGND.n1547 VGND.t188 148.846
R9916 VGND.n366 VGND.t52 148.846
R9917 VGND.n4756 VGND.t381 148.846
R9918 VGND.n1052 VGND.t220 148.846
R9919 VGND.n1100 VGND.t203 148.846
R9920 VGND.n1323 VGND.t372 148.846
R9921 VGND.n2146 VGND.t22 148.846
R9922 VGND.n2315 VGND.t112 148.846
R9923 VGND.n4209 VGND.t157 148.843
R9924 VGND.n4236 VGND.t242 148.843
R9925 VGND.n1718 VGND.t67 148.843
R9926 VGND.n1727 VGND.t37 148.843
R9927 VGND.n1654 VGND.t94 148.843
R9928 VGND.n497 VGND.t185 148.843
R9929 VGND.n504 VGND.t136 148.843
R9930 VGND.n521 VGND.t259 148.843
R9931 VGND.n524 VGND.t115 148.843
R9932 VGND.n655 VGND.t165 148.843
R9933 VGND.n672 VGND.t166 148.843
R9934 VGND.n648 VGND.t214 148.843
R9935 VGND.n1062 VGND.t192 148.843
R9936 VGND.n1195 VGND.t49 148.843
R9937 VGND.n3059 VGND.t99 148.843
R9938 VGND.n1338 VGND.t340 148.843
R9939 VGND.n1754 VGND.t53 148.843
R9940 VGND.n156 VGND.t123 148.843
R9941 VGND.n106 VGND.t388 148.843
R9942 VGND.n4768 VGND.t250 148.083
R9943 VGND.n4138 VGND.t153 148.083
R9944 VGND.n3579 VGND.t387 148.083
R9945 VGND.n761 VGND.t222 148.083
R9946 VGND.n888 VGND.t364 148.083
R9947 VGND.n3301 VGND.t139 148.083
R9948 VGND.n2282 VGND.t367 148.083
R9949 VGND.n2188 VGND.t265 148.083
R9950 VGND.n136 VGND.t90 148.083
R9951 VGND.n4222 VGND.t156 147.28
R9952 VGND.n1651 VGND.t200 147.28
R9953 VGND.n1646 VGND.t175 147.28
R9954 VGND.n1710 VGND.t117 147.28
R9955 VGND.n499 VGND.t207 147.28
R9956 VGND.n545 VGND.t155 147.28
R9957 VGND.n657 VGND.t283 147.28
R9958 VGND.n675 VGND.t284 147.28
R9959 VGND.n735 VGND.t357 147.28
R9960 VGND.n810 VGND.t320 147.28
R9961 VGND.n967 VGND.t386 147.28
R9962 VGND.n3357 VGND.t39 147.28
R9963 VGND.n1055 VGND.t331 147.28
R9964 VGND.n1150 VGND.t356 147.28
R9965 VGND.n2742 VGND.t365 147.28
R9966 VGND.n2786 VGND.t315 147.28
R9967 VGND.n2590 VGND.t371 147.28
R9968 VGND.n2647 VGND.t208 147.28
R9969 VGND.n2135 VGND.t264 147.28
R9970 VGND.n1780 VGND.t80 147.28
R9971 VGND.n5091 VGND.t130 147.28
R9972 VGND.n4091 VGND 143.296
R9973 VGND VGND.n3799 143.296
R9974 VGND.n3349 VGND 143.296
R9975 VGND.n1705 VGND 143.296
R9976 VGND.n4970 VGND 143.296
R9977 VGND.n221 VGND 143.296
R9978 VGND.n5257 VGND.t61 142.308
R9979 VGND.n5204 VGND.t354 142.308
R9980 VGND.n5589 VGND.t10 142.308
R9981 VGND.n1 VGND.t374 142.308
R9982 VGND.n5418 VGND.t322 142.308
R9983 VGND.n5345 VGND.t268 142.308
R9984 VGND.n5458 VGND.t253 142.308
R9985 VGND.n5473 VGND.t295 142.308
R9986 VGND.n5488 VGND.t330 142.308
R9987 VGND.n5503 VGND.t227 142.308
R9988 VGND.n4921 VGND.t116 142.308
R9989 VGND.n4328 VGND.t29 142.308
R9990 VGND.n4325 VGND.t5 142.308
R9991 VGND.n4321 VGND.t347 142.308
R9992 VGND.n4310 VGND.t299 142.308
R9993 VGND.n4464 VGND.t243 142.308
R9994 VGND.n1550 VGND.t209 142.308
R9995 VGND.n1757 VGND.t86 142.308
R9996 VGND.n2023 VGND.t140 142.308
R9997 VGND.n1737 VGND.t7 142.308
R9998 VGND.n4762 VGND.t30 142.308
R9999 VGND.n355 VGND.t346 142.308
R10000 VGND.n309 VGND.t272 142.308
R10001 VGND.n361 VGND.t16 142.308
R10002 VGND.n4613 VGND.t4 142.308
R10003 VGND.n4785 VGND.t64 142.308
R10004 VGND.n4798 VGND.t25 142.308
R10005 VGND.n4838 VGND.t11 142.308
R10006 VGND.n4852 VGND.t211 142.308
R10007 VGND.n4667 VGND.t298 142.308
R10008 VGND.n4708 VGND.t266 142.308
R10009 VGND.n4060 VGND.t230 142.308
R10010 VGND.n4072 VGND.t324 142.308
R10011 VGND.n4084 VGND.t274 142.308
R10012 VGND.n399 VGND.t45 142.308
R10013 VGND.n438 VGND.t100 142.308
R10014 VGND.n4110 VGND.t199 142.308
R10015 VGND.n390 VGND.t114 142.308
R10016 VGND.n564 VGND.t152 142.308
R10017 VGND.n3907 VGND.t122 142.308
R10018 VGND.n3950 VGND.t58 142.308
R10019 VGND.n709 VGND.t239 142.308
R10020 VGND.n3776 VGND.t27 142.308
R10021 VGND.n3752 VGND.t366 142.308
R10022 VGND.n772 VGND.t12 142.308
R10023 VGND.n827 VGND.t344 142.308
R10024 VGND.n836 VGND.t76 142.308
R10025 VGND.n764 VGND.t334 142.308
R10026 VGND.n783 VGND.t113 142.308
R10027 VGND.n3621 VGND.t65 142.308
R10028 VGND.n3515 VGND.t36 142.308
R10029 VGND.n3537 VGND.t378 142.308
R10030 VGND.n3552 VGND.t66 142.308
R10031 VGND.n3495 VGND.t310 142.308
R10032 VGND.n905 VGND.t183 142.308
R10033 VGND.n903 VGND.t18 142.308
R10034 VGND.n960 VGND.t285 142.308
R10035 VGND.n3371 VGND.t249 142.308
R10036 VGND.n3385 VGND.t341 142.308
R10037 VGND.n3399 VGND.t293 142.308
R10038 VGND.n3262 VGND.t235 142.308
R10039 VGND.n3253 VGND.t47 142.308
R10040 VGND.n1094 VGND.t297 142.308
R10041 VGND.n1103 VGND.t15 142.308
R10042 VGND.n3417 VGND.t328 142.308
R10043 VGND.n3428 VGND.t129 142.308
R10044 VGND.n3444 VGND.t105 142.308
R10045 VGND.n3306 VGND.t225 142.308
R10046 VGND.n2917 VGND.t57 142.308
R10047 VGND.n2899 VGND.t197 142.308
R10048 VGND.n2880 VGND.t196 142.308
R10049 VGND.n3017 VGND.t125 142.308
R10050 VGND.n3042 VGND.t124 142.308
R10051 VGND.n1146 VGND.t0 142.308
R10052 VGND.n1181 VGND.t1 142.308
R10053 VGND.n1234 VGND.t63 142.308
R10054 VGND.n1201 VGND.t164 142.308
R10055 VGND.n3008 VGND.t77 142.308
R10056 VGND.n1251 VGND.t13 142.308
R10057 VGND.n1254 VGND.t93 142.308
R10058 VGND.n2986 VGND.t42 142.308
R10059 VGND.n1257 VGND.t126 142.308
R10060 VGND.n2966 VGND.t41 142.308
R10061 VGND.n2790 VGND.t380 142.308
R10062 VGND.n2593 VGND.t8 142.308
R10063 VGND.n1359 VGND.t143 142.308
R10064 VGND.n1399 VGND.t144 142.308
R10065 VGND.n1345 VGND.t252 142.308
R10066 VGND.n1446 VGND.t307 142.308
R10067 VGND.n1336 VGND.t391 142.308
R10068 VGND.n2695 VGND.t300 142.308
R10069 VGND.n2463 VGND.t311 142.308
R10070 VGND.n2421 VGND.t142 142.308
R10071 VGND.n2418 VGND.t376 142.308
R10072 VGND.n2438 VGND.t149 142.308
R10073 VGND.n2472 VGND.t229 142.308
R10074 VGND.n2303 VGND.t74 142.308
R10075 VGND.n2170 VGND.t370 142.308
R10076 VGND.n2207 VGND.t48 142.308
R10077 VGND.n2276 VGND.t23 142.308
R10078 VGND.n2322 VGND.t195 142.308
R10079 VGND.n1480 VGND.t257 142.308
R10080 VGND.n2360 VGND.t177 142.308
R10081 VGND.n1803 VGND.t54 142.308
R10082 VGND.n1886 VGND.t390 142.308
R10083 VGND.n5109 VGND.t141 142.308
R10084 VGND.n179 VGND.t267 142.308
R10085 VGND.n5129 VGND.t213 142.308
R10086 VGND.n1921 VGND.t176 142.308
R10087 VGND.n1954 VGND.t119 142.308
R10088 VGND.n1965 VGND.t191 142.308
R10089 VGND.n1973 VGND.t389 142.308
R10090 VGND.n113 VGND.t97 142.308
R10091 VGND.n5535 VGND.t296 142.308
R10092 VGND.n1542 VGND.n1541 105.487
R10093 VGND.n173 VGND.t132 101.097
R10094 VGND.n175 VGND.t219 98.9756
R10095 VGND.n1631 VGND.t216 98.9623
R10096 VGND.n130 VGND.t111 98.822
R10097 VGND.n202 VGND.t226 98.8213
R10098 VGND.n4211 VGND.t273 98.4768
R10099 VGND.n205 VGND.t147 85.3257
R10100 VGND.n256 VGND.t168 84.847
R10101 VGND.n4317 VGND.t128 84.847
R10102 VGND.n1657 VGND.t159 84.847
R10103 VGND.n1523 VGND.t158 84.847
R10104 VGND.n442 VGND.t44 84.847
R10105 VGND.n3887 VGND.t133 84.847
R10106 VGND.n663 VGND.t181 84.847
R10107 VGND.n3243 VGND.t218 84.847
R10108 VGND.n2891 VGND.t101 84.847
R10109 VGND.n2737 VGND.t32 84.847
R10110 VGND.n1490 VGND.t228 84.847
R10111 VGND.n108 VGND.t60 84.847
R10112 VGND.n23 VGND.t24 84.847
R10113 VGND.n75 VGND.t269 84.847
R10114 VGND.n4924 VGND.t255 84.847
R10115 VGND.n1528 VGND.t348 84.847
R10116 VGND.n4029 VGND.t151 84.847
R10117 VGND.n630 VGND.t337 84.847
R10118 VGND.n639 VGND.t31 84.847
R10119 VGND.n775 VGND.t135 84.847
R10120 VGND.n889 VGND.t204 84.847
R10121 VGND.n1045 VGND.t51 84.847
R10122 VGND.n1031 VGND.t170 84.847
R10123 VGND.n2131 VGND.t373 84.847
R10124 VGND.n1462 VGND.t91 84.847
R10125 VGND.n1482 VGND.t75 84.847
R10126 VGND.n1880 VGND.t20 84.847
R10127 VGND.n5513 VGND.t349 84.847
R10128 VGND.n4824 VGND.t280 84.2473
R10129 VGND.n4664 VGND.t190 84.2473
R10130 VGND.n460 VGND.t205 84.2473
R10131 VGND.n409 VGND.t3 83.9505
R10132 VGND.n2258 VGND.t71 82.587
R10133 VGND.n2623 VGND.t355 82.587
R10134 VGND.n357 VGND.t361 82.3353
R10135 VGND.n1661 VGND.t106 82.3353
R10136 VGND.n4053 VGND.t187 82.3353
R10137 VGND.n415 VGND.t154 82.3353
R10138 VGND.n133 VGND.t238 80.3196
R10139 VGND.n653 VGND.t308 80.3195
R10140 VGND.n3407 VGND.t201 80.3195
R10141 VGND.n1270 VGND.t34 80.3195
R10142 VGND.n2486 VGND.t332 78.7329
R10143 VGND.n1931 VGND.t107 78.7329
R10144 VGND.n4218 VGND.t258 78.7329
R10145 VGND.n314 VGND.t384 78.7329
R10146 VGND.n908 VGND.t184 78.7329
R10147 VGND.n1412 VGND.t145 77.3299
R10148 VGND.n1088 VGND.t360 77.3292
R10149 VGND.n1130 VGND.t2 76.7791
R10150 VGND.n2042 VGND.t210 76.1558
R10151 VGND.n1148 VGND.t150 76.1558
R10152 VGND.n2601 VGND.t174 76.1558
R10153 VGND.n1361 VGND.t292 76.1558
R10154 VGND.n5232 VGND.n5231 76.0005
R10155 VGND.n5239 VGND.n5238 76.0005
R10156 VGND.n5228 VGND.n5227 76.0005
R10157 VGND.n65 VGND.n64 76.0005
R10158 VGND.n71 VGND.n70 76.0005
R10159 VGND.n5327 VGND.n5326 76.0005
R10160 VGND.n4947 VGND.n4946 76.0005
R10161 VGND.n4268 VGND.n4267 76.0005
R10162 VGND.n4277 VGND.n4276 76.0005
R10163 VGND.n4281 VGND.n4280 76.0005
R10164 VGND.n1679 VGND.n1678 76.0005
R10165 VGND.n1577 VGND.n1576 76.0005
R10166 VGND.n1570 VGND.n1569 76.0005
R10167 VGND.n4812 VGND.n4811 76.0005
R10168 VGND.n3963 VGND.n3962 76.0005
R10169 VGND.n3816 VGND.n3815 76.0005
R10170 VGND.n3836 VGND.n3835 76.0005
R10171 VGND.n831 VGND.n830 76.0005
R10172 VGND.n780 VGND.n779 76.0005
R10173 VGND.n917 VGND.n916 76.0005
R10174 VGND.n1037 VGND.n1036 76.0005
R10175 VGND.n2761 VGND.n2760 76.0005
R10176 VGND.n2802 VGND.n2801 76.0005
R10177 VGND.n2584 VGND.n2583 76.0005
R10178 VGND.n1473 VGND.n1472 76.0005
R10179 VGND.n1872 VGND.n1871 76.0005
R10180 VGND.n5044 VGND.n5043 76.0005
R10181 VGND.n5554 VGND.n5553 76.0005
R10182 VGND.n641 VGND.t82 75.7712
R10183 VGND.n1590 VGND.t118 75.7704
R10184 VGND.n3729 VGND.t110 75.3998
R10185 VGND.n2414 VGND.t312 75.3998
R10186 VGND.n4654 VGND.t375 75.1361
R10187 VGND.n532 VGND.t244 75.1361
R10188 VGND.n4010 VGND.t275 75.1361
R10189 VGND.n1193 VGND.t178 75.1361
R10190 VGND.n135 VGND.t237 75.1353
R10191 VGND.n2175 VGND.t353 74.7175
R10192 VGND.n1492 VGND.t148 74.6516
R10193 VGND.n1536 VGND.t56 73.7275
R10194 VGND.n313 VGND.t240 73.7275
R10195 VGND.n3153 VGND.t271 73.7275
R10196 VGND.n2164 VGND.t289 73.7275
R10197 VGND.n4416 VGND.t377 73.7268
R10198 VGND.n3153 VGND.t14 73.7268
R10199 VGND.n2862 VGND.t43 73.7268
R10200 VGND.n4216 VGND.t127 68.948
R10201 VGND.n2218 VGND.t9 68.948
R10202 VGND.n5237 VGND.t33 68.6994
R10203 VGND.n4279 VGND.t102 68.6994
R10204 VGND.n1568 VGND.t96 68.6994
R10205 VGND.n4414 VGND.t95 68.3876
R10206 VGND.n2863 VGND.t167 68.3876
R10207 VGND.n731 VGND.n730 34.6358
R10208 VGND.n3744 VGND.n3743 34.6358
R10209 VGND.n1211 VGND.n1210 34.6358
R10210 VGND.n1210 VGND.n1209 34.6358
R10211 VGND.n2667 VGND.n2666 34.6358
R10212 VGND.n1787 VGND.n1786 34.6358
R10213 VGND.n4901 VGND.n258 34.6358
R10214 VGND.n4387 VGND.n4326 34.6358
R10215 VGND.n4435 VGND.n4434 34.6358
R10216 VGND.n539 VGND.n538 34.6358
R10217 VGND.n413 VGND.n404 34.6358
R10218 VGND.n475 VGND.n439 34.6358
R10219 VGND.n4107 VGND.n394 34.6358
R10220 VGND.n730 VGND.n729 34.6358
R10221 VGND.n714 VGND.n660 34.6358
R10222 VGND.n848 VGND.n838 34.6358
R10223 VGND.n3534 VGND.n3520 34.6358
R10224 VGND.n3544 VGND.n3543 34.6358
R10225 VGND.n3506 VGND.n3505 34.6358
R10226 VGND.n3506 VGND.n887 34.6358
R10227 VGND.n3368 VGND.n3355 34.6358
R10228 VGND.n2925 VGND.n2924 34.6358
R10229 VGND.n2925 VGND.n2900 34.6358
R10230 VGND.n1169 VGND.n1168 34.6358
R10231 VGND.n1174 VGND.n1173 34.6358
R10232 VGND.n1175 VGND.n1174 34.6358
R10233 VGND.n1175 VGND.n1142 34.6358
R10234 VGND.n1217 VGND.n1216 34.6358
R10235 VGND.n2610 VGND.n2587 34.6358
R10236 VGND.n1387 VGND.n1386 34.6358
R10237 VGND.n1392 VGND.n1391 34.6358
R10238 VGND.n1393 VGND.n1392 34.6358
R10239 VGND.n1393 VGND.n1355 34.6358
R10240 VGND.n1406 VGND.n1405 34.6358
R10241 VGND.n2455 VGND.n2454 34.6358
R10242 VGND.n2352 VGND.n2351 34.6358
R10243 VGND.n1907 VGND.n1906 34.6358
R10244 VGND.n1962 VGND.n1866 34.6358
R10245 VGND.n69 VGND.t281 34.2973
R10246 VGND.n63 VGND.t270 34.2973
R10247 VGND.n5325 VGND.t72 34.2973
R10248 VGND.n5552 VGND.t254 34.2973
R10249 VGND.n4945 VGND.t6 34.2973
R10250 VGND.n1677 VGND.t160 34.2973
R10251 VGND.n4810 VGND.t343 34.2973
R10252 VGND.n3961 VGND.t109 34.2973
R10253 VGND.n3834 VGND.t301 34.2973
R10254 VGND.n3814 VGND.t134 34.2973
R10255 VGND.n829 VGND.t294 34.2973
R10256 VGND.n778 VGND.t40 34.2973
R10257 VGND.n915 VGND.t19 34.2973
R10258 VGND.n1035 VGND.t236 34.2973
R10259 VGND.n2759 VGND.t21 34.2973
R10260 VGND.n2800 VGND.t286 34.2973
R10261 VGND.n2582 VGND.t171 34.2973
R10262 VGND.n1471 VGND.t172 34.2973
R10263 VGND.n5042 VGND.t46 34.2973
R10264 VGND.n1870 VGND.t68 34.2973
R10265 VGND.n2334 VGND.n1485 32.0005
R10266 VGND.n5238 VGND.n5237 31.4781
R10267 VGND.n4280 VGND.n4279 31.4781
R10268 VGND.n1569 VGND.n1568 31.4781
R10269 VGND.n1211 VGND.n1199 29.8804
R10270 VGND.n1581 VGND.n1542 29.4862
R10271 VGND.n4257 VGND.n4256 28.4695
R10272 VGND.n2043 VGND.n2042 28.4695
R10273 VGND.n4824 VGND.n4823 28.4695
R10274 VGND.n4665 VGND.n4664 28.4695
R10275 VGND.n1162 VGND.n1148 28.4695
R10276 VGND.n2601 VGND.n2600 28.4695
R10277 VGND.n1380 VGND.n1361 28.4695
R10278 VGND.n2220 VGND.n2219 28.4695
R10279 VGND.n1324 VGND.n1322 27.4829
R10280 VGND.n5216 VGND.n5214 26.001
R10281 VGND.n1695 VGND.n1659 25.977
R10282 VGND.n4579 VGND.n4578 25.977
R10283 VGND.n4795 VGND.n4749 25.977
R10284 VGND.n691 VGND.n690 25.977
R10285 VGND.n691 VGND.n665 25.977
R10286 VGND.n849 VGND.n848 25.977
R10287 VGND.n2929 VGND.n2900 25.977
R10288 VGND.n4587 VGND.n310 25.6926
R10289 VGND.n3048 VGND.n3047 25.6926
R10290 VGND.n2469 VGND.n2410 25.6926
R10291 VGND.n5581 VGND.n5580 25.6926
R10292 VGND.n5595 VGND.n5594 25.6926
R10293 VGND.n5412 VGND.n5411 25.6926
R10294 VGND.n5361 VGND.n5359 25.6926
R10295 VGND.n5350 VGND.n5349 25.6926
R10296 VGND.n5470 VGND.n5468 25.6926
R10297 VGND.n5477 VGND.n32 25.6926
R10298 VGND.n5492 VGND.n31 25.6926
R10299 VGND.n4388 VGND.n4387 25.6926
R10300 VGND.n2053 VGND.n1521 25.6926
R10301 VGND.n4618 VGND.n4617 25.6926
R10302 VGND.n4831 VGND.n4830 25.6926
R10303 VGND.n4836 VGND.n4835 25.6926
R10304 VGND.n4844 VGND.n4843 25.6926
R10305 VGND.n4850 VGND.n4849 25.6926
R10306 VGND.n4673 VGND.n300 25.6926
R10307 VGND.n4649 VGND.n4647 25.6926
R10308 VGND.n4071 VGND.n4070 25.6926
R10309 VGND.n414 VGND.n413 25.6926
R10310 VGND.n431 VGND.n430 25.6926
R10311 VGND.n483 VGND.n401 25.6926
R10312 VGND.n476 VGND.n475 25.6926
R10313 VGND.n4108 VGND.n4107 25.6926
R10314 VGND.n4116 VGND.n4115 25.6926
R10315 VGND.n3906 VGND.n3905 25.6926
R10316 VGND.n3939 VGND.n3938 25.6926
R10317 VGND.n3948 VGND.n3947 25.6926
R10318 VGND.n710 VGND.n660 25.6926
R10319 VGND.n3774 VGND.n3773 25.6926
R10320 VGND.n3758 VGND.n3757 25.6926
R10321 VGND.n3750 VGND.n3749 25.6926
R10322 VGND.n822 VGND.n770 25.6926
R10323 VGND.n3619 VGND.n3618 25.6926
R10324 VGND.n805 VGND.n804 25.6926
R10325 VGND.n3535 VGND.n3534 25.6926
R10326 VGND.n3543 VGND.n3542 25.6926
R10327 VGND.n3558 VGND.n3557 25.6926
R10328 VGND.n3510 VGND.n887 25.6926
R10329 VGND.n3502 VGND.n3501 25.6926
R10330 VGND.n946 VGND.n945 25.6926
R10331 VGND.n956 VGND.n955 25.6926
R10332 VGND.n3369 VGND.n3368 25.6926
R10333 VGND.n3397 VGND.n3396 25.6926
R10334 VGND.n3250 VGND.n3248 25.6926
R10335 VGND.n3238 VGND.n1044 25.6926
R10336 VGND.n1082 VGND.n1081 25.6926
R10337 VGND.n3415 VGND.n3414 25.6926
R10338 VGND.n3426 VGND.n3425 25.6926
R10339 VGND.n3434 VGND.n3433 25.6926
R10340 VGND.n3442 VGND.n3441 25.6926
R10341 VGND.n2916 VGND.n2904 25.6926
R10342 VGND.n1168 VGND.n1167 25.6926
R10343 VGND.n1230 VGND.n1190 25.6926
R10344 VGND.n2978 VGND.n2977 25.6926
R10345 VGND.n2973 VGND.n2972 25.6926
R10346 VGND.n2796 VGND.n1332 25.6926
R10347 VGND.n1386 VGND.n1385 25.6926
R10348 VGND.n2659 VGND.n2658 25.6926
R10349 VGND.n2666 VGND.n1337 25.6926
R10350 VGND.n2454 VGND.n2413 25.6926
R10351 VGND.n2470 VGND.n2469 25.6926
R10352 VGND.n2150 VGND.n2125 25.6926
R10353 VGND.n2194 VGND.n2193 25.6926
R10354 VGND.n2351 VGND.n1481 25.6926
R10355 VGND.n2356 VGND.n2355 25.6926
R10356 VGND.n5115 VGND.n5114 25.6926
R10357 VGND.n5127 VGND.n5126 25.6926
R10358 VGND.n1906 VGND.n1879 25.6926
R10359 VGND.n1919 VGND.n1918 25.6926
R10360 VGND.n1963 VGND.n1962 25.6926
R10361 VGND.n5070 VGND.n5069 25.6926
R10362 VGND.n5058 VGND.n5057 25.6926
R10363 VGND.n5533 VGND.n5532 25.6926
R10364 VGND.n1216 VGND.n1215 25.6506
R10365 VGND.n4398 VGND.n4322 25.224
R10366 VGND.n4079 VGND.n4078 25.224
R10367 VGND.n4035 VGND.n500 25.224
R10368 VGND.n3588 VGND.n766 25.224
R10369 VGND.n3382 VGND.n3354 25.224
R10370 VGND.n2588 VGND.n2587 25.224
R10371 VGND.n2493 VGND.n1467 25.224
R10372 VGND.n5246 VGND.n5200 24.9894
R10373 VGND.n5406 VGND.n5405 24.9894
R10374 VGND.n5384 VGND.n74 24.9894
R10375 VGND.n5334 VGND.n77 24.9894
R10376 VGND.n926 VGND.n925 24.9894
R10377 VGND.n2797 VGND.n2796 24.9894
R10378 VGND.n2611 VGND.n2610 24.9894
R10379 VGND.n2478 VGND.n1476 24.9894
R10380 VGND.n5547 VGND.n5546 24.9894
R10381 VGND.n2885 VGND.n1273 24.9308
R10382 VGND.n4573 VGND.n4572 24.9283
R10383 VGND.n3601 VGND.n3600 24.9283
R10384 VGND.n4244 VGND.n4243 24.8035
R10385 VGND.n5247 VGND.n5246 24.4711
R10386 VGND.n5214 VGND.n5201 24.4711
R10387 VGND.n5581 VGND.n21 24.4711
R10388 VGND.n5385 VGND.n5384 24.4711
R10389 VGND.n5335 VGND.n5334 24.4711
R10390 VGND.n5468 VGND.n33 24.4711
R10391 VGND.n5478 VGND.n5477 24.4711
R10392 VGND.n5493 VGND.n5492 24.4711
R10393 VGND.n4243 VGND.n4220 24.4711
R10394 VGND.n4674 VGND.n4673 24.4711
R10395 VGND.n551 VGND.n550 24.4711
R10396 VGND.n685 VGND.n671 24.4711
R10397 VGND.n3558 VGND.n3517 24.4711
R10398 VGND.n3233 VGND.n1044 24.4711
R10399 VGND.n1066 VGND.n1054 24.4711
R10400 VGND.n2905 VGND.n2904 24.4711
R10401 VGND.n2753 VGND.n2740 24.4711
R10402 VGND.n2455 VGND.n2411 24.4711
R10403 VGND.n1884 VGND.n1882 24.4711
R10404 VGND.n5546 VGND.n5509 24.4711
R10405 VGND.n5532 VGND.n5511 24.4711
R10406 VGND.n4587 VGND.n311 24.3747
R10407 VGND.n2886 VGND.n2885 24.1648
R10408 VGND.n2910 VGND.n2907 24.0946
R10409 VGND.n483 VGND.n400 24.0841
R10410 VGND.n2461 VGND.n2460 24.0841
R10411 VGND.n410 VGND.n404 23.7181
R10412 VGND.n843 VGND.n842 23.7181
R10413 VGND.n3248 VGND.n1042 23.7181
R10414 VGND.n3058 VGND.n1131 23.7181
R10415 VGND.n2782 VGND.n2738 23.7181
R10416 VGND.n2148 VGND.n2147 23.7181
R10417 VGND.n1786 VGND.n1753 23.7181
R10418 VGND.n5368 VGND.n28 23.7181
R10419 VGND.n4887 VGND.n4886 23.7181
R10420 VGND.n4434 VGND.n4315 23.7181
R10421 VGND.n1706 VGND.n1704 23.7181
R10422 VGND.n1549 VGND.n1548 23.7181
R10423 VGND.n4682 VGND.n4681 23.7181
R10424 VGND.n4036 VGND.n4035 23.7181
R10425 VGND.n4020 VGND.n4019 23.7181
R10426 VGND.n538 VGND.n523 23.7181
R10427 VGND.n3891 VGND.n3890 23.7181
R10428 VGND.n876 VGND.n770 23.7181
R10429 VGND.n805 VGND.n776 23.7181
R10430 VGND.n1063 VGND.n1054 23.7181
R10431 VGND.n3409 VGND.n3408 23.7181
R10432 VGND.n3269 VGND.n3268 23.7181
R10433 VGND.n2910 VGND.n2909 23.7181
R10434 VGND.n1154 VGND.n1151 23.7181
R10435 VGND.n1155 VGND.n1154 23.7181
R10436 VGND.n2851 VGND.n2850 23.7181
R10437 VGND.n1405 VGND.n1404 23.7181
R10438 VGND.n2493 VGND.n2492 23.7181
R10439 VGND.n2197 VGND.n2176 23.7181
R10440 VGND.n1882 VGND.n1881 23.7181
R10441 VGND.n3475 VGND.n3474 23.6966
R10442 VGND.n1704 VGND.n1656 23.4101
R10443 VGND.n3726 VGND.n3724 23.4101
R10444 VGND.n2478 VGND.n2477 23.4101
R10445 VGND.n3006 VGND.n3005 23.4027
R10446 VGND.n1406 VGND.n1349 23.4027
R10447 VGND.n5269 VGND.n27 22.9652
R10448 VGND.n3905 VGND.n3895 22.9652
R10449 VGND.n715 VGND.n714 22.9652
R10450 VGND.n1169 VGND.n1144 22.4034
R10451 VGND.n1387 VGND.n1357 22.4034
R10452 VGND.n1728 VGND.n1726 22.2123
R10453 VGND.n4066 VGND.n4044 22.2123
R10454 VGND.n4070 VGND.n4044 22.2123
R10455 VGND.n2941 VGND.n2940 22.2123
R10456 VGND.n3288 VGND.n1040 21.9776
R10457 VGND.n3902 VGND.n3895 21.4593
R10458 VGND.n2940 VGND.n2896 21.4593
R10459 VGND.n5069 VGND.n114 21.4593
R10460 VGND.n2043 VGND.n2040 21.283
R10461 VGND.n4767 VGND.n4757 21.283
R10462 VGND.n4823 VGND.n296 21.283
R10463 VGND.n457 VGND.n456 21.283
R10464 VGND.n4137 VGND.n392 21.283
R10465 VGND.n528 VGND.n527 21.283
R10466 VGND.n3931 VGND.n3889 21.283
R10467 VGND.n3801 VGND.n645 21.283
R10468 VGND.n3595 VGND.n3594 21.283
R10469 VGND.n3569 VGND.n3568 21.283
R10470 VGND.n3497 VGND.n3494 21.283
R10471 VGND.n3577 VGND.n3576 21.283
R10472 VGND.n3308 VGND.n3305 21.283
R10473 VGND.n1163 VGND.n1162 21.283
R10474 VGND.n2600 VGND.n2595 21.283
R10475 VGND.n1381 VGND.n1380 21.283
R10476 VGND.n2443 VGND.n2416 21.283
R10477 VGND.n2289 VGND.n1494 21.283
R10478 VGND.n2220 VGND.n2217 21.283
R10479 VGND.n2187 VGND.n2179 21.283
R10480 VGND.n147 VGND.n146 21.283
R10481 VGND.n177 VGND.n176 21.0829
R10482 VGND.n3273 VGND.n3272 20.7985
R10483 VGND.n4372 VGND.n4371 20.422
R10484 VGND.n4959 VGND.n4920 20.0456
R10485 VGND VGND.n4065 20.0456
R10486 VGND.n2878 VGND 20.0456
R10487 VGND.n3902 VGND.n3901 19.9534
R10488 VGND VGND.n3912 19.6691
R10489 VGND.n4910 VGND.n4909 19.577
R10490 VGND.n4768 VGND.n4767 19.3636
R10491 VGND.n4138 VGND.n4137 19.3636
R10492 VGND.n3595 VGND.n761 19.3636
R10493 VGND.n3494 VGND.n888 19.3636
R10494 VGND.n2188 VGND.n2187 19.3636
R10495 VGND.n146 VGND.n136 19.3636
R10496 VGND.n4556 VGND.n4555 19.2926
R10497 VGND.n4078 VGND.n4077 19.2926
R10498 VGND.n817 VGND.n816 19.2926
R10499 VGND.n1438 VGND.n1437 19.2499
R10500 VGND.n2754 VGND.n2753 18.9637
R10501 VGND.n729 VGND.n650 18.824
R10502 VGND.n686 VGND.n685 18.824
R10503 VGND.n2924 VGND.n2923 18.824
R10504 VGND.n1206 VGND 18.78
R10505 VGND.n863 VGND.n862 18.5894
R10506 VGND.n734 VGND 18.0711
R10507 VGND.n4083 VGND.n4040 17.7867
R10508 VGND.n869 VGND.n868 17.7867
R10509 VGND.n766 VGND.n765 17.7867
R10510 VGND.n3383 VGND.n3382 17.7867
R10511 VGND.n3191 VGND.n3190 17.7867
R10512 VGND.n1437 VGND.n1346 17.7867
R10513 VGND.n5075 VGND.n111 17.7867
R10514 VGND.n1179 VGND.n1142 17.7459
R10515 VGND.n1397 VGND.n1355 17.7459
R10516 VGND.n444 VGND.n443 17.3181
R10517 VGND.n2140 VGND.n2130 17.3181
R10518 VGND.n110 VGND.n109 17.3181
R10519 VGND.n4257 VGND.n4215 16.9936
R10520 VGND.n3932 VGND.n3931 16.9936
R10521 VGND.n3732 VGND.n645 16.9936
R10522 VGND.n3569 VGND.n886 16.9936
R10523 VGND.n2444 VGND.n2443 16.9936
R10524 VGND.n2820 VGND.n1322 16.9417
R10525 VGND VGND 16.8587
R10526 VGND VGND 16.8587
R10527 VGND VGND 16.8587
R10528 VGND VGND 16.8587
R10529 VGND VGND 16.8587
R10530 VGND VGND 16.8587
R10531 VGND.n2432 VGND.n2431 16.7494
R10532 VGND.n4935 VGND.n4934 16.7494
R10533 VGND.n939 VGND.n938 16.7494
R10534 VGND.n3259 VGND.n3257 16.7494
R10535 VGND.n3313 VGND.n1033 16.7494
R10536 VGND.n2997 VGND.n2996 16.7494
R10537 VGND.n2992 VGND.n2991 16.7494
R10538 VGND.n2985 VGND.n2984 16.7494
R10539 VGND.n2437 VGND.n2436 16.7494
R10540 VGND.n2281 VGND.n1495 16.7494
R10541 VGND.n2213 VGND.n2212 16.7494
R10542 VGND.n2206 VGND.n2172 16.7494
R10543 VGND.n1971 VGND.n1970 16.7494
R10544 VGND.n2923 VGND.n2902 16.6573
R10545 VGND.n2935 VGND.n2897 16.6573
R10546 VGND.n2773 VGND.n2739 16.6573
R10547 VGND.n1563 VGND.n1549 16.5652
R10548 VGND.n1944 VGND.n1943 16.3306
R10549 VGND.n4580 VGND.n4579 16.2808
R10550 VGND.n4555 VGND.n4554 16.2808
R10551 VGND.n4782 VGND.n4753 16.2808
R10552 VGND.n4796 VGND.n4795 16.2808
R10553 VGND.n3175 VGND.n3174 16.2808
R10554 VGND.n2930 VGND.n2929 16.2808
R10555 VGND.n2141 VGND.n2140 16.2808
R10556 VGND.n4240 VGND.n4220 16.1887
R10557 VGND.n3821 VGND.n3820 16.0462
R10558 VGND.n3841 VGND.n3840 16.0462
R10559 VGND.n790 VGND.n789 16.0462
R10560 VGND.n4940 VGND.n4939 16.0462
R10561 VGND.n3956 VGND.n3955 16.0462
R10562 VGND.n3488 VGND.n3486 15.9516
R10563 VGND.n2028 VGND.n1531 15.9044
R10564 VGND.n1939 VGND.n1875 15.9044
R10565 VGND VGND.n535 15.8505
R10566 VGND VGND.n153 15.8505
R10567 VGND.n447 VGND.n446 15.8123
R10568 VGND.n811 VGND.n774 15.8123
R10569 VGND.n1197 VGND.n1196 15.8123
R10570 VGND.n338 VGND.n337 15.7682
R10571 VGND.n1764 VGND.n1763 15.5279
R10572 VGND.n324 VGND.n315 15.5279
R10573 VGND.n4132 VGND.n4131 15.5279
R10574 VGND.n2308 VGND.n1489 15.5279
R10575 VGND.n2310 VGND.n2308 15.5279
R10576 VGND.n5107 VGND.n5106 15.5279
R10577 VGND.n4783 VGND.n4782 15.4968
R10578 VGND.n1231 VGND.n1230 15.4358
R10579 VGND.n850 VGND.n849 15.3918
R10580 VGND.n1957 VGND.n1867 15.3918
R10581 VGND.n5209 VGND.n5208 15.1514
R10582 VGND.n5587 VGND.n5586 15.1514
R10583 VGND.n14 VGND.n13 15.1514
R10584 VGND.n5463 VGND.n5462 15.1514
R10585 VGND.n4447 VGND.n4446 15.1514
R10586 VGND.n1668 VGND.n1660 15.1514
R10587 VGND.n1735 VGND.n1734 15.1514
R10588 VGND.n4055 VGND.n4047 15.1514
R10589 VGND.n3550 VGND.n3549 15.1514
R10590 VGND.n1067 VGND.n1066 15.1514
R10591 VGND.n3189 VGND.n3188 15.1514
R10592 VGND.n1630 VGND.n1539 15.0834
R10593 VGND.n157 VGND.n134 15.0834
R10594 VGND.n4308 VGND 15.0593
R10595 VGND.n501 VGND.n500 15.0593
R10596 VGND.n3564 VGND.n3563 14.9001
R10597 VGND.n3524 VGND.n3523 14.8179
R10598 VGND.n5516 VGND.n5514 14.8179
R10599 VGND.n5260 VGND.n27 14.775
R10600 VGND.n5573 VGND.n26 14.775
R10601 VGND.n5419 VGND.n29 14.775
R10602 VGND.n5567 VGND.n30 14.775
R10603 VGND.n4319 VGND.n4318 14.775
R10604 VGND.n252 VGND.n251 14.775
R10605 VGND.n2019 VGND.n1532 14.775
R10606 VGND.n1527 VGND.n1525 14.775
R10607 VGND.n4761 VGND.n4760 14.775
R10608 VGND.n4804 VGND.n298 14.775
R10609 VGND.n4704 VGND.n4703 14.775
R10610 VGND.n4090 VGND.n496 14.775
R10611 VGND.n3976 VGND.n629 14.775
R10612 VGND.n703 VGND.n662 14.775
R10613 VGND.n876 VGND.n875 14.775
R10614 VGND.n3390 VGND.n3353 14.775
R10615 VGND.n3352 VGND.n3350 14.775
R10616 VGND.n3297 VGND.n3296 14.775
R10617 VGND.n3015 VGND.n3014 14.775
R10618 VGND.n1240 VGND.n1140 14.775
R10619 VGND.n1240 VGND.n1239 14.775
R10620 VGND.n3014 VGND.n1138 14.775
R10621 VGND.n2788 VGND.n2787 14.775
R10622 VGND.n2648 VGND.n1340 14.775
R10623 VGND.n1368 VGND.n1367 14.775
R10624 VGND.n1404 VGND.n1351 14.775
R10625 VGND.n2426 VGND.n2425 14.775
R10626 VGND.n2300 VGND.n2298 14.775
R10627 VGND.n2319 VGND.n2317 14.775
R10628 VGND.n1888 VGND.n1887 14.775
R10629 VGND.n1926 VGND.n126 14.775
R10630 VGND.n1929 VGND.n126 14.775
R10631 VGND.n5567 VGND.n5566 14.775
R10632 VGND.n1650 VGND.n1649 14.6829
R10633 VGND.n688 VGND.n687 14.6829
R10634 VGND.n687 VGND.n686 14.6829
R10635 VGND.n3169 VGND.n1105 14.6388
R10636 VGND.n1659 VGND.n1658 14.3064
R10637 VGND.n420 VGND.n402 14.3064
R10638 VGND.n723 VGND.n722 14.3064
R10639 VGND.n1076 VGND.n1075 14.3064
R10640 VGND.n2906 VGND.n2905 14.3064
R10641 VGND.n4805 VGND.n4804 14.0717
R10642 VGND.n4059 VGND.n4058 14.022
R10643 VGND.n1233 VGND.n1232 14.022
R10644 VGND.n4233 VGND.n4232 13.5534
R10645 VGND.n4290 VGND.n4208 13.5534
R10646 VGND.n1603 VGND.n1602 13.5534
R10647 VGND.n1645 VGND.n1644 13.5534
R10648 VGND.n4568 VGND.n4567 13.5534
R10649 VGND.n724 VGND.n723 13.5534
R10650 VGND.n722 VGND.n654 13.5534
R10651 VGND.n717 VGND.n716 13.5534
R10652 VGND.n3183 VGND.n3182 13.5534
R10653 VGND.n1327 VGND.n1326 13.5534
R10654 VGND.n190 VGND.n176 13.5534
R10655 VGND.n1672 VGND.n1671 13.3188
R10656 VGND.n4024 VGND.n503 13.2691
R10657 VGND.n4917 VGND.n254 13.177
R10658 VGND.n4914 VGND.n255 13.177
R10659 VGND.n4227 VGND.n4226 13.177
R10660 VGND.n4238 VGND.n4237 13.177
R10661 VGND.n1598 VGND.n1597 13.177
R10662 VGND.n4776 VGND.n4755 13.177
R10663 VGND.n320 VGND.n319 13.177
R10664 VGND.n3901 VGND.n3896 13.177
R10665 VGND.n3227 VGND.n3226 13.177
R10666 VGND.n1417 VGND.n1347 13.177
R10667 VGND.n1222 VGND.n1192 12.9808
R10668 VGND.n5573 VGND.n24 12.8005
R10669 VGND.n76 VGND.n28 12.8005
R10670 VGND.n4928 VGND.n4927 12.8005
R10671 VGND.n4966 VGND.n254 12.8005
R10672 VGND.n4966 VGND.n255 12.8005
R10673 VGND.n4207 VGND.n250 12.8005
R10674 VGND.n1663 VGND.n1662 12.8005
R10675 VGND.n4052 VGND.n4049 12.8005
R10676 VGND.n421 VGND.n420 12.8005
R10677 VGND.n3897 VGND.n3896 12.8005
R10678 VGND.n703 VGND.n700 12.8005
R10679 VGND.n677 VGND.n676 12.8005
R10680 VGND.n3359 VGND.n3358 12.8005
R10681 VGND.n3198 VGND.n1051 12.8005
R10682 VGND.n2945 VGND.n1269 12.8005
R10683 VGND.n2744 VGND.n2743 12.8005
R10684 VGND.n4256 VGND.n4216 12.7128
R10685 VGND.n2219 VGND.n2218 12.7128
R10686 VGND.n3198 VGND.n3197 12.4838
R10687 VGND.n1217 VGND.n1197 12.424
R10688 VGND.n4301 VGND.n250 12.3566
R10689 VGND.n202 VGND.n201 12.3437
R10690 VGND.n130 VGND.n128 12.3437
R10691 VGND.n1719 VGND.n1717 12.0476
R10692 VGND.n1943 VGND.n1875 12.0476
R10693 VGND.n4430 VGND.n4315 11.7989
R10694 VGND.n2854 VGND.n2851 11.7989
R10695 VGND.n2492 VGND.n1470 11.7989
R10696 VGND.n4291 VGND.n4290 11.6711
R10697 VGND.n682 VGND.n671 11.6711
R10698 VGND.n1671 VGND.n1660 11.2946
R10699 VGND.n4058 VGND.n4047 11.2946
R10700 VGND.n3174 VGND.n3173 11.2946
R10701 VGND.n2343 VGND.n1483 11.2946
R10702 VGND.n3182 VGND.n3181 11.0103
R10703 VGND.n2344 VGND.n2343 11.0103
R10704 VGND.n1617 VGND.n1590 11.0085
R10705 VGND.n3852 VGND.n641 11.0085
R10706 VGND.n2623 VGND.n2622 11.0085
R10707 VGND.n2259 VGND.n2258 11.0085
R10708 VGND.n4446 VGND.n4311 10.9181
R10709 VGND.n550 VGND.n520 10.9181
R10710 VGND.n3289 VGND.n3288 10.9181
R10711 VGND.n2871 VGND.n2870 10.9181
R10712 VGND.n1418 VGND.n1417 10.9181
R10713 VGND.n4079 VGND.n4040 10.9181
R10714 VGND.n4262 VGND.n4261 10.9046
R10715 VGND.n211 VGND.n128 10.9046
R10716 VGND.n4408 VGND.n4316 10.8605
R10717 VGND.n1607 VGND.n1591 10.8605
R10718 VGND.n4030 VGND.n4028 10.8605
R10719 VGND.n4013 VGND.n4009 10.8605
R10720 VGND.n563 VGND.n519 10.8605
R10721 VGND.n3805 VGND.n3804 10.8605
R10722 VGND.n3853 VGND.n3852 10.8605
R10723 VGND.n3244 VGND.n3242 10.8605
R10724 VGND.n2892 VGND.n2890 10.8605
R10725 VGND.n2622 VGND.n2580 10.8605
R10726 VGND.n1373 VGND.n1372 10.8605
R10727 VGND.n462 VGND.n441 10.8605
R10728 VGND.n4419 VGND.n251 10.7135
R10729 VGND.n4233 VGND.n4222 10.7135
R10730 VGND.n4237 VGND.n4236 10.7135
R10731 VGND.n4209 VGND.n4208 10.7135
R10732 VGND.n1719 VGND.n1718 10.7135
R10733 VGND.n1651 VGND.n1650 10.7135
R10734 VGND.n1728 VGND.n1727 10.7135
R10735 VGND.n1646 VGND.n1645 10.7135
R10736 VGND.n1711 VGND.n1710 10.7135
R10737 VGND.n1706 VGND.n1654 10.7135
R10738 VGND.n4090 VGND.n497 10.7135
R10739 VGND.n4036 VGND.n499 10.7135
R10740 VGND.n4019 VGND.n504 10.7135
R10741 VGND.n546 VGND.n545 10.7135
R10742 VGND.n521 VGND.n520 10.7135
R10743 VGND.n524 VGND.n523 10.7135
R10744 VGND.n653 VGND.n650 10.7135
R10745 VGND.n724 VGND.n653 10.7135
R10746 VGND.n655 VGND.n654 10.7135
R10747 VGND.n717 VGND.n657 10.7135
R10748 VGND.n681 VGND.n672 10.7135
R10749 VGND.n677 VGND.n675 10.7135
R10750 VGND.n735 VGND.n734 10.7135
R10751 VGND.n811 VGND.n810 10.7135
R10752 VGND.n3357 VGND.n3356 10.7135
R10753 VGND.n1058 VGND.n1055 10.7135
R10754 VGND.n1063 VGND.n1062 10.7135
R10755 VGND.n3407 VGND.n3350 10.7135
R10756 VGND.n3408 VGND.n3407 10.7135
R10757 VGND.n2941 VGND.n1270 10.7135
R10758 VGND.n2945 VGND.n1270 10.7135
R10759 VGND.n1155 VGND.n1150 10.7135
R10760 VGND.n1196 VGND.n1195 10.7135
R10761 VGND.n3059 VGND.n3058 10.7135
R10762 VGND.n2870 VGND.n1275 10.7135
R10763 VGND.n2787 VGND.n2786 10.7135
R10764 VGND.n1330 VGND.n1327 10.7135
R10765 VGND.n2590 VGND.n2589 10.7135
R10766 VGND.n2652 VGND.n1338 10.7135
R10767 VGND.n2648 VGND.n2647 10.7135
R10768 VGND.n2136 VGND.n2135 10.7135
R10769 VGND.n2176 VGND.n2175 10.7135
R10770 VGND.n1781 VGND.n1780 10.7135
R10771 VGND.n1754 VGND.n1753 10.7135
R10772 VGND.n157 VGND.n156 10.7135
R10773 VGND.n5092 VGND.n5091 10.7135
R10774 VGND.n107 VGND.n106 10.7135
R10775 VGND.n1781 VGND.n1779 10.5417
R10776 VGND.n2653 VGND.n2652 10.5417
R10777 VGND.n5092 VGND.n105 10.5417
R10778 VGND.n1603 VGND.n1592 10.4353
R10779 VGND.n348 VGND.n347 10.2509
R10780 VGND.n695 VGND.n665 10.2509
R10781 VGND.n1173 VGND.n1144 10.171
R10782 VGND.n1391 VGND.n1357 10.171
R10783 VGND.n1215 VGND.n1199 10.0827
R10784 VGND.n201 VGND.n170 10.0462
R10785 VGND.n1618 VGND.n1617 10.0021
R10786 VGND.n3040 VGND.n3039 9.86687
R10787 VGND.n1711 VGND.n1653 9.78874
R10788 VGND.n690 VGND.n689 9.78874
R10789 VGND.n682 VGND.n681 9.78874
R10790 VGND.n4712 VGND.n4711 9.3005
R10791 VGND.n4735 VGND.n4734 9.3005
R10792 VGND.n4737 VGND.n4736 9.3005
R10793 VGND.n566 VGND.n565 9.3005
R10794 VGND.n488 VGND.n487 9.3005
R10795 VGND.n493 VGND.n492 9.3005
R10796 VGND.n571 VGND.n570 9.3005
R10797 VGND.n573 VGND.n572 9.3005
R10798 VGND.n3873 VGND.n3872 9.3005
R10799 VGND.n3875 VGND.n3874 9.3005
R10800 VGND.n964 VGND.n963 9.3005
R10801 VGND.n3650 VGND.n3649 9.3005
R10802 VGND.n3138 VGND.n3137 9.3005
R10803 VGND.n3202 VGND.n3201 9.3005
R10804 VGND.n3336 VGND.n3335 9.3005
R10805 VGND.n3338 VGND.n3337 9.3005
R10806 VGND.n2965 VGND.n2964 9.3005
R10807 VGND.n2699 VGND.n2698 9.3005
R10808 VGND.n2722 VGND.n2721 9.3005
R10809 VGND.n2724 VGND.n2723 9.3005
R10810 VGND.n2563 VGND.n2562 9.3005
R10811 VGND.n2364 VGND.n2363 9.3005
R10812 VGND.n2390 VGND.n2389 9.3005
R10813 VGND.n2388 VGND.n2387 9.3005
R10814 VGND.n1807 VGND.n1806 9.3005
R10815 VGND.n2005 VGND.n2004 9.3005
R10816 VGND.n2007 VGND.n2006 9.3005
R10817 VGND.n2081 VGND.n2080 9.3005
R10818 VGND.n215 VGND.n214 9.3005
R10819 VGND.n220 VGND.n219 9.3005
R10820 VGND.n1861 VGND.n1860 9.3005
R10821 VGND.n1859 VGND.n1858 9.3005
R10822 VGND.n5158 VGND.n5157 9.3005
R10823 VGND.n4476 VGND.n4475 9.3005
R10824 VGND.n4371 VGND.n4370 9.3005
R10825 VGND.n4357 VGND.n4356 9.3005
R10826 VGND.n4350 VGND.n4349 9.3005
R10827 VGND.n4369 VGND.n253 9.3005
R10828 VGND.n4348 VGND.n4347 9.3005
R10829 VGND.n4479 VGND.n4478 9.3005
R10830 VGND.n4306 VGND.n4305 9.3005
R10831 VGND.n5427 VGND.n5426 9.3005
R10832 VGND.n5302 VGND.n5301 9.3005
R10833 VGND.n5305 VGND.n5304 9.3005
R10834 VGND.n5434 VGND.n5433 9.3005
R10835 VGND.n5425 VGND.n5424 9.3005
R10836 VGND.n716 VGND.n715 9.03579
R10837 VGND.n4302 VGND.n4301 9.00185
R10838 VGND.n4718 VGND.n4717 9.0005
R10839 VGND.n4739 VGND.n4738 9.0005
R10840 VGND.n4733 VGND.n4732 9.0005
R10841 VGND.n598 VGND.n597 9.0005
R10842 VGND.n491 VGND.n490 9.0005
R10843 VGND.n486 VGND.n485 9.0005
R10844 VGND.n575 VGND.n574 9.0005
R10845 VGND.n569 VGND.n568 9.0005
R10846 VGND.n3877 VGND.n3876 9.0005
R10847 VGND.n3871 VGND.n3870 9.0005
R10848 VGND.n993 VGND.n992 9.0005
R10849 VGND.n3655 VGND.n3654 9.0005
R10850 VGND.n3204 VGND.n3203 9.0005
R10851 VGND.n3140 VGND.n3139 9.0005
R10852 VGND.n3340 VGND.n3339 9.0005
R10853 VGND.n3334 VGND.n3333 9.0005
R10854 VGND.n2962 VGND.n2961 9.0005
R10855 VGND.n2705 VGND.n2704 9.0005
R10856 VGND.n2558 VGND.n2557 9.0005
R10857 VGND.n2726 VGND.n2725 9.0005
R10858 VGND.n2720 VGND.n2719 9.0005
R10859 VGND.n2370 VGND.n2369 9.0005
R10860 VGND.n2273 VGND.n2272 9.0005
R10861 VGND.n2392 VGND.n2391 9.0005
R10862 VGND.n2386 VGND.n2385 9.0005
R10863 VGND.n1824 VGND.n1823 9.0005
R10864 VGND.n2009 VGND.n2008 9.0005
R10865 VGND.n2003 VGND.n2002 9.0005
R10866 VGND.n2086 VGND.n2085 9.0005
R10867 VGND.n1857 VGND.n1856 9.0005
R10868 VGND.n1863 VGND.n1862 9.0005
R10869 VGND.n218 VGND.n217 9.0005
R10870 VGND.n213 VGND.n212 9.0005
R10871 VGND.n5163 VGND.n5162 9.0005
R10872 VGND.n4368 VGND.n4329 9.0005
R10873 VGND.n4362 VGND.n4361 9.0005
R10874 VGND.n4352 VGND.n4351 9.0005
R10875 VGND.n4346 VGND.n4345 9.0005
R10876 VGND.n4474 VGND.n4473 9.0005
R10877 VGND.n4481 VGND.n4480 9.0005
R10878 VGND.n5307 VGND.n5306 9.0005
R10879 VGND.n5300 VGND.n5299 9.0005
R10880 VGND.n5270 VGND.n5269 9.0005
R10881 VGND.n5429 VGND.n5428 9.0005
R10882 VGND.n5439 VGND.n5438 9.0005
R10883 VGND.n5423 VGND.n5422 9.0005
R10884 VGND.n190 VGND.n175 8.97441
R10885 VGND.n1606 VGND.n1605 8.88606
R10886 VGND.n4460 VGND.n4459 8.75144
R10887 VGND.n4399 VGND.n4398 8.70217
R10888 VGND.n1464 VGND.n1463 8.65932
R10889 VGND VGND 8.42962
R10890 VGND VGND 8.42962
R10891 VGND VGND 8.42962
R10892 VGND VGND 8.42962
R10893 VGND VGND 8.42962
R10894 VGND VGND 8.42962
R10895 VGND VGND 8.42962
R10896 VGND VGND 8.42962
R10897 VGND VGND 8.42962
R10898 VGND VGND 8.42962
R10899 VGND VGND 8.42962
R10900 VGND VGND 8.42962
R10901 VGND VGND 8.42962
R10902 VGND VGND 8.42962
R10903 VGND VGND 8.42962
R10904 VGND VGND 8.42962
R10905 VGND VGND 8.42962
R10906 VGND.n2335 VGND.n2334 8.3666
R10907 VGND.n1159 VGND.n1158 8.36259
R10908 VGND.n2603 VGND.n2591 8.36259
R10909 VGND.n1232 VGND.n1231 8.28285
R10910 VGND.n1193 VGND.n1192 7.83347
R10911 VGND.n4255 VGND.n248 7.82272
R10912 VGND.n4095 VGND.n4094 7.82272
R10913 VGND.n3933 VGND.n3932 7.82272
R10914 VGND.n3572 VGND.n886 7.82272
R10915 VGND.n2223 VGND.n2124 7.82272
R10916 VGND.n4215 VGND.n249 7.76113
R10917 VGND.n4825 VGND.n294 7.65314
R10918 VGND.n461 VGND.n459 7.65314
R10919 VGND.n4655 VGND.n4654 7.56414
R10920 VGND.n4011 VGND.n4010 7.56414
R10921 VGND.n535 VGND.n532 7.56414
R10922 VGND.n153 VGND.n135 7.56414
R10923 VGND.n1599 VGND.n1598 7.52991
R10924 VGND.n4567 VGND.n4566 7.52991
R10925 VGND.n3850 VGND.n3849 7.34052
R10926 VGND.n2624 VGND.n2623 7.23528
R10927 VGND.n4458 VGND 7.15344
R10928 VGND.n2897 VGND.n2896 7.15344
R10929 VGND.n5126 VGND.n100 7.15344
R10930 VGND.n4211 VGND.n4210 6.82364
R10931 VGND.n4654 VGND.n301 6.82364
R10932 VGND.n4010 VGND.n505 6.82364
R10933 VGND.n532 VGND.n525 6.82364
R10934 VGND.n1194 VGND.n1193 6.82364
R10935 VGND.n155 VGND.n135 6.82364
R10936 VGND.n4918 VGND.n4917 6.77697
R10937 VGND.n2907 VGND.n2906 6.77697
R10938 VGND.n4261 VGND.n4215 6.61527
R10939 VGND.n4883 VGND.n259 6.57117
R10940 VGND.n4883 VGND.n4882 6.57117
R10941 VGND.n4409 VGND.n4408 6.57117
R10942 VGND.n1547 VGND.n1546 6.57117
R10943 VGND.n1607 VGND.n1606 6.57117
R10944 VGND.n365 VGND.n363 6.57117
R10945 VGND.n366 VGND.n365 6.57117
R10946 VGND.n4756 VGND.n4754 6.57117
R10947 VGND.n4028 VGND.n502 6.57117
R10948 VGND.n441 VGND.n440 6.57117
R10949 VGND.n396 VGND.n395 6.57117
R10950 VGND.n4094 VGND.n396 6.57117
R10951 VGND.n519 VGND.n518 6.57117
R10952 VGND.n635 VGND.n634 6.57117
R10953 VGND.n3932 VGND.n635 6.57117
R10954 VGND.n3804 VGND.n644 6.57117
R10955 VGND.n3513 VGND.n3512 6.57117
R10956 VGND.n3513 VGND.n886 6.57117
R10957 VGND.n3242 VGND.n1043 6.57117
R10958 VGND.n1072 VGND.n1052 6.57117
R10959 VGND.n1072 VGND.n1071 6.57117
R10960 VGND.n1100 VGND.n1099 6.57117
R10961 VGND.n1099 VGND.n1097 6.57117
R10962 VGND.n2890 VGND.n1271 6.57117
R10963 VGND.n1372 VGND.n1364 6.57117
R10964 VGND.n1323 VGND.n1321 6.57117
R10965 VGND.n2145 VGND.n2128 6.57117
R10966 VGND.n2146 VGND.n2145 6.57117
R10967 VGND.n2259 VGND.n2257 6.57117
R10968 VGND.n2314 VGND.n1488 6.57117
R10969 VGND.n2315 VGND.n2314 6.57117
R10970 VGND.n1605 VGND.n1592 6.4005
R10971 VGND.n3529 VGND.n3528 6.4005
R10972 VGND.n5516 VGND.n5515 6.4005
R10973 VGND.n4663 VGND.n301 6.38812
R10974 VGND.n809 VGND.n775 6.38812
R10975 VGND.n968 VGND.n889 6.38812
R10976 VGND.n2785 VGND.n2737 6.38812
R10977 VGND.n1493 VGND.n1490 6.38812
R10978 VGND.n2132 VGND.n2131 6.38812
R10979 VGND.n2 VGND 6.27264
R10980 VGND.n5216 VGND.n5215 6.26433
R10981 VGND.n26 VGND.n25 6.26433
R10982 VGND.n5580 VGND.n22 6.26433
R10983 VGND.n5594 VGND.n20 6.26433
R10984 VGND.n5361 VGND.n5360 6.26433
R10985 VGND.n5470 VGND.n5469 6.26433
R10986 VGND.n4934 VGND.n4926 6.26433
R10987 VGND.n4939 VGND.n4923 6.26433
R10988 VGND.n4959 VGND.n4958 6.26433
R10989 VGND.n4903 VGND.n4902 6.26433
R10990 VGND.n4402 VGND.n4319 6.26433
R10991 VGND.n4410 VGND.n252 6.26433
R10992 VGND.n1668 VGND.n1667 6.26433
R10993 VGND.n1656 VGND.n1655 6.26433
R10994 VGND.n2028 VGND.n2027 6.26433
R10995 VGND.n1527 VGND.n1526 6.26433
R10996 VGND.n2040 VGND.n1524 6.26433
R10997 VGND.n2053 VGND.n2052 6.26433
R10998 VGND.n4763 VGND.n4757 6.26433
R10999 VGND.n327 VGND.n315 6.26433
R11000 VGND.n4554 VGND.n4553 6.26433
R11001 VGND.n298 VGND.n297 6.26433
R11002 VGND.n4830 VGND.n293 6.26433
R11003 VGND.n4843 VGND.n291 6.26433
R11004 VGND.n4649 VGND.n4648 6.26433
R11005 VGND.n4055 VGND.n4054 6.26433
R11006 VGND.n4065 VGND.n4045 6.26433
R11007 VGND.n4077 VGND.n4042 6.26433
R11008 VGND.n416 VGND.n414 6.26433
R11009 VGND.n467 VGND.n466 6.26433
R11010 VGND.n4100 VGND.n4099 6.26433
R11011 VGND.n4115 VGND.n393 6.26433
R11012 VGND.n3912 VGND.n3893 6.26433
R11013 VGND.n3938 VGND.n633 6.26433
R11014 VGND.n3955 VGND.n631 6.26433
R11015 VGND.n629 VGND.n628 6.26433
R11016 VGND.n707 VGND.n662 6.26433
R11017 VGND.n696 VGND.n695 6.26433
R11018 VGND.n3726 VGND.n3725 6.26433
R11019 VGND.n3757 VGND.n3727 6.26433
R11020 VGND.n3542 VGND.n3519 6.26433
R11021 VGND.n3557 VGND.n3518 6.26433
R11022 VGND.n3568 VGND.n3516 6.26433
R11023 VGND.n3511 VGND.n3510 6.26433
R11024 VGND.n3488 VGND.n3487 6.26433
R11025 VGND.n3390 VGND.n3389 6.26433
R11026 VGND.n3352 VGND.n3351 6.26433
R11027 VGND.n3259 VGND.n3258 6.26433
R11028 VGND.n3239 VGND.n3238 6.26433
R11029 VGND.n1089 VGND.n1087 6.26433
R11030 VGND.n3188 VGND.n3187 6.26433
R11031 VGND.n3433 VGND.n1024 6.26433
R11032 VGND.n3308 VGND.n3307 6.26433
R11033 VGND.n3314 VGND.n3313 6.26433
R11034 VGND.n2919 VGND.n2902 6.26433
R11035 VGND.n2879 VGND.n2878 6.26433
R11036 VGND.n3022 VGND.n1136 6.26433
R11037 VGND.n3047 VGND.n1132 6.26433
R11038 VGND.n1180 VGND.n1179 6.26433
R11039 VGND.n1239 VGND.n1186 6.26433
R11040 VGND.n1235 VGND.n1186 6.26433
R11041 VGND.n1226 VGND.n1190 6.26433
R11042 VGND.n1138 VGND.n1137 6.26433
R11043 VGND.n2996 VGND.n1252 6.26433
R11044 VGND.n2773 VGND.n2772 6.26433
R11045 VGND.n2595 VGND.n2594 6.26433
R11046 VGND.n1369 VGND.n1368 6.26433
R11047 VGND.n1374 VGND.n1373 6.26433
R11048 VGND.n1398 VGND.n1397 6.26433
R11049 VGND.n1413 VGND.n1411 6.26433
R11050 VGND.n2431 VGND.n2423 6.26433
R11051 VGND.n2436 VGND.n2420 6.26433
R11052 VGND.n2413 VGND.n2412 6.26433
R11053 VGND.n2410 VGND.n2409 6.26433
R11054 VGND.n2477 VGND.n1477 6.26433
R11055 VGND.n2300 VGND.n2299 6.26433
R11056 VGND.n2291 VGND.n2289 6.26433
R11057 VGND.n2284 VGND.n2281 6.26433
R11058 VGND.n2142 VGND.n2141 6.26433
R11059 VGND.n2154 VGND.n2125 6.26433
R11060 VGND.n2208 VGND.n2171 6.26433
R11061 VGND.n2202 VGND.n2172 6.26433
R11062 VGND.n2189 VGND.n2178 6.26433
R11063 VGND.n2183 VGND.n2179 6.26433
R11064 VGND.n2319 VGND.n2318 6.26433
R11065 VGND.n2310 VGND.n2309 6.26433
R11066 VGND.n161 VGND.n134 6.26433
R11067 VGND.n5114 VGND.n102 6.26433
R11068 VGND.n1879 VGND.n1878 6.26433
R11069 VGND.n1926 VGND.n1925 6.26433
R11070 VGND.n1939 VGND.n1938 6.26433
R11071 VGND.n1970 VGND.n1865 6.26433
R11072 VGND.n5566 VGND.n5508 6.26433
R11073 VGND.n4926 VGND.n4925 6.26433
R11074 VGND.n4923 VGND.n4922 6.26433
R11075 VGND.n4214 VGND.n4213 6.26433
R11076 VGND.n4266 VGND.n4214 6.26433
R11077 VGND.n1586 VGND.n1540 6.26433
R11078 VGND.n1612 VGND.n1591 6.26433
R11079 VGND.n4770 VGND.n4769 6.26433
R11080 VGND.n4753 VGND.n4752 6.26433
R11081 VGND.n296 VGND.n295 6.26433
R11082 VGND.n4669 VGND.n4668 6.26433
R11083 VGND.n4061 VGND.n4045 6.26433
R11084 VGND.n4073 VGND.n4042 6.26433
R11085 VGND.n4086 VGND.n496 6.26433
R11086 VGND.n4086 VGND.n4085 6.26433
R11087 VGND.n392 VGND.n391 6.26433
R11088 VGND.n4139 VGND.n389 6.26433
R11089 VGND.n4013 VGND.n4012 6.26433
R11090 VGND.n534 VGND.n533 6.26433
R11091 VGND.n3908 VGND.n3893 6.26433
R11092 VGND.n3889 VGND.n3888 6.26433
R11093 VGND.n708 VGND.n707 6.26433
R11094 VGND.n697 VGND.n696 6.26433
R11095 VGND.n3848 VGND.n3847 6.26433
R11096 VGND.n3594 VGND.n763 6.26433
R11097 VGND.n3599 VGND.n3598 6.26433
R11098 VGND.n3497 VGND.n3496 6.26433
R11099 VGND.n3250 VGND.n3249 6.26433
R11100 VGND.n2919 VGND.n2918 6.26433
R11101 VGND.n2935 VGND.n2934 6.26433
R11102 VGND.n2934 VGND.n2933 6.26433
R11103 VGND.n2881 VGND.n2879 6.26433
R11104 VGND.n1164 VGND.n1163 6.26433
R11105 VGND.n1182 VGND.n1180 6.26433
R11106 VGND.n1226 VGND.n1225 6.26433
R11107 VGND.n1225 VGND.n1224 6.26433
R11108 VGND.n2987 VGND.n1255 6.26433
R11109 VGND.n1332 VGND.n1331 6.26433
R11110 VGND.n1382 VGND.n1381 6.26433
R11111 VGND.n1400 VGND.n1398 6.26433
R11112 VGND.n1411 VGND.n1410 6.26433
R11113 VGND.n2423 VGND.n2422 6.26433
R11114 VGND.n2420 VGND.n2419 6.26433
R11115 VGND.n2439 VGND.n2416 6.26433
R11116 VGND.n2291 VGND.n2290 6.26433
R11117 VGND.n2284 VGND.n2283 6.26433
R11118 VGND.n2217 VGND.n2169 6.26433
R11119 VGND.n1893 VGND.n1892 6.26433
R11120 VGND.n211 VGND.n129 6.26433
R11121 VGND.n152 VGND.n151 6.26433
R11122 VGND.n143 VGND.n142 6.26433
R11123 VGND.n1410 VGND.n1349 6.26374
R11124 VGND.n4572 VGND.n4571 6.2636
R11125 VGND.n3600 VGND.n3599 6.2636
R11126 VGND.n2887 VGND.n2886 6.26328
R11127 VGND.n5518 VGND.n5517 6.2505
R11128 VGND.n1530 VGND.n1529 6.02403
R11129 VGND.n3913 VGND 6.02403
R11130 VGND.n1209 VGND 6.02403
R11131 VGND.n4459 VGND 5.72682
R11132 VGND.n5268 VGND.n5267 5.64756
R11133 VGND.n4066 VGND 5.64756
R11134 VGND.n731 VGND 5.64756
R11135 VGND.n689 VGND.n688 5.64756
R11136 VGND.n2875 VGND 5.64756
R11137 VGND.n1614 VGND.n1613 5.47606
R11138 VGND.n1586 VGND.n1585 5.37524
R11139 VGND.n328 VGND.n327 5.37524
R11140 VGND.n3576 VGND.n768 5.37524
R11141 VGND.n2155 VGND.n2154 5.37524
R11142 VGND.n203 VGND.n129 5.37524
R11143 VGND.n162 VGND.n161 5.37524
R11144 VGND.n4886 VGND.n259 5.35702
R11145 VGND.n1548 VGND.n1547 5.35702
R11146 VGND.n4549 VGND.n366 5.35702
R11147 VGND.n4776 VGND.n4756 5.35702
R11148 VGND.n4663 VGND.n4662 5.35702
R11149 VGND.n410 VGND.n409 5.35702
R11150 VGND.n1075 VGND.n1052 5.35702
R11151 VGND.n3183 VGND.n1100 5.35702
R11152 VGND.n2820 VGND.n1323 5.35702
R11153 VGND.n2147 VGND.n2146 5.35702
R11154 VGND.n2317 VGND.n2315 5.35702
R11155 VGND.n1493 VGND.n1492 5.33915
R11156 VGND.n4256 VGND.n4255 5.28304
R11157 VGND.n2219 VGND.n2124 5.28304
R11158 VGND.n4920 VGND.n4919 5.27109
R11159 VGND.n1485 VGND.n1484 5.27109
R11160 VGND.n4025 VGND 5.24305
R11161 VGND.n133 VGND.n130 5.23624
R11162 VGND.n205 VGND.n202 5.23624
R11163 VGND.n1633 VGND.n1632 5.17489
R11164 VGND.n2602 VGND.n2592 5.12314
R11165 VGND.n2625 VGND 5.10688
R11166 VGND.n4287 VGND.n4212 5.09669
R11167 VGND.n1160 VGND.n1149 5.08226
R11168 VGND.n175 VGND.n174 4.97399
R11169 VGND.n1631 VGND.n1630 4.94421
R11170 VGND.n70 VGND.n69 4.85762
R11171 VGND.n64 VGND.n63 4.85762
R11172 VGND.n5326 VGND.n5325 4.85762
R11173 VGND.n5553 VGND.n5552 4.85762
R11174 VGND.n4946 VGND.n4945 4.85762
R11175 VGND.n1678 VGND.n1677 4.85762
R11176 VGND.n4811 VGND.n4810 4.85762
R11177 VGND.n3962 VGND.n3961 4.85762
R11178 VGND.n3835 VGND.n3834 4.85762
R11179 VGND.n3815 VGND.n3814 4.85762
R11180 VGND.n830 VGND.n829 4.85762
R11181 VGND.n779 VGND.n778 4.85762
R11182 VGND.n916 VGND.n915 4.85762
R11183 VGND.n1036 VGND.n1035 4.85762
R11184 VGND.n2760 VGND.n2759 4.85762
R11185 VGND.n2801 VGND.n2800 4.85762
R11186 VGND.n2583 VGND.n2582 4.85762
R11187 VGND.n1472 VGND.n1471 4.85762
R11188 VGND.n5043 VGND.n5042 4.85762
R11189 VGND.n1871 VGND.n1870 4.85762
R11190 VGND.n3 VGND.n2 4.8005
R11191 VGND.n3528 VGND.n3522 4.8005
R11192 VGND.n857 VGND.n855 4.76901
R11193 VGND.n920 VGND.n913 4.76901
R11194 VGND.n1950 VGND.n1949 4.76901
R11195 VGND.n3486 VGND.n3485 4.70498
R11196 VGND.n3480 VGND.n3479 4.70498
R11197 VGND.n3614 VGND.n3613 4.67844
R11198 VGND.n951 VGND.n950 4.67844
R11199 VGND.n3921 VGND.n3920 4.65418
R11200 VGND.n1215 VGND.n1214 4.65418
R11201 VGND.n3484 VGND.n3483 4.65256
R11202 VGND.n2886 VGND.n1272 4.65245
R11203 VGND.n558 VGND.n557 4.65216
R11204 VGND.n3600 VGND.n760 4.65211
R11205 VGND.n1896 VGND.n1895 4.65211
R11206 VGND.n3197 VGND.n3196 4.65209
R11207 VGND.n4784 VGND.n4783 4.65205
R11208 VGND.n3007 VGND.n3006 4.65205
R11209 VGND.n1408 VGND.n1349 4.65205
R11210 VGND.n2883 VGND.n1273 4.65131
R11211 VGND.n4612 VGND.n4611 4.6505
R11212 VGND.n4621 VGND.n4620 4.6505
R11213 VGND.n4675 VGND.n4674 4.6505
R11214 VGND.n4677 VGND.n4676 4.6505
R11215 VGND.n4679 VGND.n4678 4.6505
R11216 VGND.n4695 VGND.n4694 4.6505
R11217 VGND.n4703 VGND.n4702 4.6505
R11218 VGND.n321 VGND.n320 4.6505
R11219 VGND.n325 VGND.n324 4.6505
R11220 VGND.n339 VGND.n338 4.6505
R11221 VGND.n341 VGND.n340 4.6505
R11222 VGND.n343 VGND.n342 4.6505
R11223 VGND.n347 VGND.n346 4.6505
R11224 VGND.n4579 VGND.n356 4.6505
R11225 VGND.n4567 VGND.n359 4.6505
R11226 VGND.n4566 VGND.n4565 4.6505
R11227 VGND.n4555 VGND.n362 4.6505
R11228 VGND.n4615 VGND.n4614 4.6505
R11229 VGND.n4617 VGND.n4616 4.6505
R11230 VGND.n4666 VGND.n4665 4.6505
R11231 VGND.n4670 VGND.n4669 4.6505
R11232 VGND.n4691 VGND.n4690 4.6505
R11233 VGND.n4699 VGND.n4698 4.6505
R11234 VGND.n4705 VGND.n4704 4.6505
R11235 VGND.n4707 VGND.n4706 4.6505
R11236 VGND.n4710 VGND.n4709 4.6505
R11237 VGND.n4833 VGND.n292 4.6505
R11238 VGND.n4804 VGND.n4803 4.6505
R11239 VGND.n4795 VGND.n4794 4.6505
R11240 VGND.n4792 VGND.n4750 4.6505
R11241 VGND.n4782 VGND.n4781 4.6505
R11242 VGND.n4774 VGND.n4755 4.6505
R11243 VGND.n4847 VGND.n4846 4.6505
R11244 VGND.n4845 VGND.n4844 4.6505
R11245 VGND.n4843 VGND.n4842 4.6505
R11246 VGND.n4840 VGND.n4839 4.6505
R11247 VGND.n4837 VGND.n4836 4.6505
R11248 VGND.n4835 VGND.n4834 4.6505
R11249 VGND.n4832 VGND.n4831 4.6505
R11250 VGND.n4830 VGND.n4829 4.6505
R11251 VGND.n4827 VGND.n4826 4.6505
R11252 VGND.n4823 VGND.n4822 4.6505
R11253 VGND.n4821 VGND.n296 4.6505
R11254 VGND.n4819 VGND.n4818 4.6505
R11255 VGND.n4817 VGND.n4816 4.6505
R11256 VGND.n4814 VGND.n4813 4.6505
R11257 VGND.n4809 VGND.n4808 4.6505
R11258 VGND.n4806 VGND.n4805 4.6505
R11259 VGND.n4802 VGND.n298 4.6505
R11260 VGND.n4800 VGND.n4799 4.6505
R11261 VGND.n4797 VGND.n4796 4.6505
R11262 VGND.n4793 VGND.n4749 4.6505
R11263 VGND.n4791 VGND.n4790 4.6505
R11264 VGND.n4789 VGND.n4788 4.6505
R11265 VGND.n4787 VGND.n4786 4.6505
R11266 VGND.n4780 VGND.n4753 4.6505
R11267 VGND.n4777 VGND.n4776 4.6505
R11268 VGND.n4776 VGND.n4775 4.6505
R11269 VGND.n4773 VGND.n4772 4.6505
R11270 VGND.n4771 VGND.n4770 4.6505
R11271 VGND.n4769 VGND 4.6505
R11272 VGND.n4767 VGND.n4766 4.6505
R11273 VGND.n4765 VGND.n4757 4.6505
R11274 VGND.n4764 VGND.n4763 4.6505
R11275 VGND.n4856 VGND.n4855 4.6505
R11276 VGND.n4854 VGND.n4853 4.6505
R11277 VGND.n4851 VGND.n4850 4.6505
R11278 VGND.n4849 VGND.n4848 4.6505
R11279 VGND.n4701 VGND.n4700 4.6505
R11280 VGND.n4697 VGND.n4696 4.6505
R11281 VGND.n4693 VGND.n4692 4.6505
R11282 VGND.n4689 VGND.n4688 4.6505
R11283 VGND.n4687 VGND.n4686 4.6505
R11284 VGND.n4685 VGND.n4684 4.6505
R11285 VGND.n4683 VGND.n4682 4.6505
R11286 VGND.n4673 VGND 4.6505
R11287 VGND.n4672 VGND.n300 4.6505
R11288 VGND.n4639 VGND.n4638 4.6505
R11289 VGND.n4637 VGND.n4636 4.6505
R11290 VGND.n4635 VGND.n4634 4.6505
R11291 VGND.n4633 VGND.n4632 4.6505
R11292 VGND.n4631 VGND.n4630 4.6505
R11293 VGND.n4629 VGND.n4628 4.6505
R11294 VGND.n4627 VGND.n4626 4.6505
R11295 VGND.n4625 VGND.n4624 4.6505
R11296 VGND.n4623 VGND.n4622 4.6505
R11297 VGND.n4619 VGND.n4618 4.6505
R11298 VGND.n323 VGND.n322 4.6505
R11299 VGND VGND.n315 4.6505
R11300 VGND.n327 VGND.n326 4.6505
R11301 VGND.n329 VGND.n328 4.6505
R11302 VGND.n331 VGND.n330 4.6505
R11303 VGND.n333 VGND.n332 4.6505
R11304 VGND.n337 VGND.n336 4.6505
R11305 VGND.n345 VGND.n344 4.6505
R11306 VGND.n349 VGND.n348 4.6505
R11307 VGND.n351 VGND.n350 4.6505
R11308 VGND.n353 VGND.n310 4.6505
R11309 VGND.n4587 VGND.n4586 4.6505
R11310 VGND.n4585 VGND.n311 4.6505
R11311 VGND.n4584 VGND.n4583 4.6505
R11312 VGND.n4581 VGND.n4580 4.6505
R11313 VGND.n4578 VGND.n4577 4.6505
R11314 VGND.n4576 VGND.n4575 4.6505
R11315 VGND.n4574 VGND.n4573 4.6505
R11316 VGND.n4571 VGND.n4570 4.6505
R11317 VGND.n4564 VGND.n4563 4.6505
R11318 VGND.n4562 VGND.n4561 4.6505
R11319 VGND.n4560 VGND.n4559 4.6505
R11320 VGND.n4557 VGND.n4556 4.6505
R11321 VGND.n4553 VGND.n4552 4.6505
R11322 VGND.n4550 VGND.n4549 4.6505
R11323 VGND.n4641 VGND.n4640 4.6505
R11324 VGND.n4647 VGND.n4646 4.6505
R11325 VGND.n4645 VGND.n4644 4.6505
R11326 VGND.n4643 VGND.n4642 4.6505
R11327 VGND.n4657 VGND.n4656 4.6505
R11328 VGND.n4653 VGND.n4652 4.6505
R11329 VGND.n4650 VGND.n4649 4.6505
R11330 VGND.n4662 VGND.n4660 4.6505
R11331 VGND.n4662 VGND.n4661 4.6505
R11332 VGND.n4140 VGND.n389 4.6505
R11333 VGND.n4131 VGND.n4130 4.6505
R11334 VGND.n538 VGND 4.6505
R11335 VGND.n544 VGND.n543 4.6505
R11336 VGND.n552 VGND.n551 4.6505
R11337 VGND.n556 VGND.n555 4.6505
R11338 VGND.n420 VGND.n419 4.6505
R11339 VGND.n422 VGND.n421 4.6505
R11340 VGND.n424 VGND.n423 4.6505
R11341 VGND.n428 VGND.n427 4.6505
R11342 VGND.n451 VGND.n444 4.6505
R11343 VGND.n450 VGND.n445 4.6505
R11344 VGND.n449 VGND.n446 4.6505
R11345 VGND VGND.n4139 4.6505
R11346 VGND.n4137 VGND.n4136 4.6505
R11347 VGND.n4103 VGND.n4102 4.6505
R11348 VGND.n540 VGND.n539 4.6505
R11349 VGND.n547 VGND.n546 4.6505
R11350 VGND.n549 VGND.n520 4.6505
R11351 VGND.n563 VGND.n562 4.6505
R11352 VGND.n4021 VGND.n4020 4.6505
R11353 VGND.n4022 VGND.n503 4.6505
R11354 VGND.n4033 VGND.n500 4.6505
R11355 VGND.n4037 VGND.n4036 4.6505
R11356 VGND.n4088 VGND.n496 4.6505
R11357 VGND.n4081 VGND.n4040 4.6505
R11358 VGND.n4078 VGND.n4041 4.6505
R11359 VGND.n4068 VGND.n4044 4.6505
R11360 VGND.n4058 VGND 4.6505
R11361 VGND.n4057 VGND.n4047 4.6505
R11362 VGND.n4019 VGND.n4018 4.6505
R11363 VGND.n4024 VGND.n4023 4.6505
R11364 VGND.n4026 VGND.n4025 4.6505
R11365 VGND.n4031 VGND.n4030 4.6505
R11366 VGND.n4035 VGND.n4034 4.6505
R11367 VGND.n4090 VGND.n4089 4.6505
R11368 VGND.n4087 VGND.n4086 4.6505
R11369 VGND.n4085 VGND.n4039 4.6505
R11370 VGND.n4083 VGND.n4082 4.6505
R11371 VGND.n4080 VGND.n4079 4.6505
R11372 VGND.n4077 VGND.n4076 4.6505
R11373 VGND.n4075 VGND.n4042 4.6505
R11374 VGND.n4074 VGND.n4073 4.6505
R11375 VGND.n4071 VGND.n4043 4.6505
R11376 VGND.n4070 VGND.n4069 4.6505
R11377 VGND.n4067 VGND.n4066 4.6505
R11378 VGND.n4065 VGND.n4064 4.6505
R11379 VGND.n4063 VGND.n4045 4.6505
R11380 VGND.n4062 VGND.n4061 4.6505
R11381 VGND.n4059 VGND.n4046 4.6505
R11382 VGND.n4056 VGND.n4055 4.6505
R11383 VGND.n4054 VGND.n4048 4.6505
R11384 VGND.n4007 VGND.n4006 4.6505
R11385 VGND.n4014 VGND.n4013 4.6505
R11386 VGND.n560 VGND.n559 4.6505
R11387 VGND.n554 VGND.n553 4.6505
R11388 VGND.n550 VGND 4.6505
R11389 VGND.n542 VGND.n541 4.6505
R11390 VGND.n4099 VGND.n4098 4.6505
R11391 VGND.n4101 VGND.n4100 4.6505
R11392 VGND.n4105 VGND.n4104 4.6505
R11393 VGND.n4106 VGND.n394 4.6505
R11394 VGND.n4107 VGND 4.6505
R11395 VGND.n4109 VGND.n4108 4.6505
R11396 VGND.n4112 VGND.n4111 4.6505
R11397 VGND.n4115 VGND.n4114 4.6505
R11398 VGND.n4117 VGND.n4116 4.6505
R11399 VGND.n4119 VGND.n4118 4.6505
R11400 VGND.n4121 VGND.n4120 4.6505
R11401 VGND.n4123 VGND.n4122 4.6505
R11402 VGND.n4125 VGND.n4124 4.6505
R11403 VGND.n4127 VGND.n4126 4.6505
R11404 VGND.n4129 VGND.n4128 4.6505
R11405 VGND.n4133 VGND.n4132 4.6505
R11406 VGND.n4135 VGND.n392 4.6505
R11407 VGND.n412 VGND.n404 4.6505
R11408 VGND.n413 VGND 4.6505
R11409 VGND.n417 VGND.n416 4.6505
R11410 VGND.n426 VGND.n425 4.6505
R11411 VGND.n430 VGND.n429 4.6505
R11412 VGND.n432 VGND.n431 4.6505
R11413 VGND.n434 VGND.n433 4.6505
R11414 VGND.n436 VGND.n400 4.6505
R11415 VGND.n483 VGND.n482 4.6505
R11416 VGND.n481 VGND.n401 4.6505
R11417 VGND.n480 VGND.n479 4.6505
R11418 VGND.n477 VGND.n476 4.6505
R11419 VGND.n475 VGND.n474 4.6505
R11420 VGND.n473 VGND.n439 4.6505
R11421 VGND.n472 VGND.n471 4.6505
R11422 VGND.n470 VGND.n469 4.6505
R11423 VGND.n468 VGND.n467 4.6505
R11424 VGND.n466 VGND.n465 4.6505
R11425 VGND.n463 VGND.n462 4.6505
R11426 VGND.n458 VGND.n457 4.6505
R11427 VGND.n456 VGND.n455 4.6505
R11428 VGND.n454 VGND.n453 4.6505
R11429 VGND.n537 VGND.n523 4.6505
R11430 VGND.n529 VGND.n528 4.6505
R11431 VGND.n534 VGND.n531 4.6505
R11432 VGND.n527 VGND.n526 4.6505
R11433 VGND.n4096 VGND.n4095 4.6505
R11434 VGND.n3780 VGND.n3726 4.6505
R11435 VGND.n678 VGND.n677 4.6505
R11436 VGND.n683 VGND.n682 4.6505
R11437 VGND.n684 VGND.n671 4.6505
R11438 VGND.n686 VGND.n670 4.6505
R11439 VGND.n688 VGND.n668 4.6505
R11440 VGND.n689 VGND.n667 4.6505
R11441 VGND.n690 VGND.n666 4.6505
R11442 VGND.n693 VGND.n665 4.6505
R11443 VGND.n704 VGND.n703 4.6505
R11444 VGND.n715 VGND.n659 4.6505
R11445 VGND.n716 VGND.n658 4.6505
R11446 VGND.n718 VGND.n717 4.6505
R11447 VGND.n722 VGND.n721 4.6505
R11448 VGND.n723 VGND.n652 4.6505
R11449 VGND.n725 VGND.n724 4.6505
R11450 VGND.n729 VGND.n728 4.6505
R11451 VGND.n3778 VGND.n3777 4.6505
R11452 VGND.n3775 VGND.n3774 4.6505
R11453 VGND.n3773 VGND.n3772 4.6505
R11454 VGND.n3822 VGND.n3821 4.6505
R11455 VGND.n3824 VGND.n3823 4.6505
R11456 VGND.n3826 VGND.n3825 4.6505
R11457 VGND.n3828 VGND.n3827 4.6505
R11458 VGND.n3838 VGND.n3837 4.6505
R11459 VGND.n3840 VGND.n3839 4.6505
R11460 VGND.n3842 VGND.n3841 4.6505
R11461 VGND.n3854 VGND.n3853 4.6505
R11462 VGND.n3941 VGND.n632 4.6505
R11463 VGND.n3926 VGND.n3891 4.6505
R11464 VGND.n3915 VGND.n3892 4.6505
R11465 VGND.n3904 VGND.n3895 4.6505
R11466 VGND.n3901 VGND.n3900 4.6505
R11467 VGND.n3972 VGND.n3971 4.6505
R11468 VGND.n3970 VGND.n3969 4.6505
R11469 VGND.n3968 VGND.n3967 4.6505
R11470 VGND.n3965 VGND.n3964 4.6505
R11471 VGND.n3960 VGND.n3959 4.6505
R11472 VGND.n3957 VGND.n3956 4.6505
R11473 VGND.n3955 VGND.n3954 4.6505
R11474 VGND.n3952 VGND.n3951 4.6505
R11475 VGND.n3949 VGND.n3948 4.6505
R11476 VGND.n3947 VGND.n3946 4.6505
R11477 VGND.n3945 VGND.n3944 4.6505
R11478 VGND.n3943 VGND.n3942 4.6505
R11479 VGND.n3940 VGND.n3939 4.6505
R11480 VGND.n3938 VGND.n3937 4.6505
R11481 VGND.n3936 VGND.n633 4.6505
R11482 VGND.n3934 VGND.n3933 4.6505
R11483 VGND.n3931 VGND.n3930 4.6505
R11484 VGND.n3929 VGND.n3889 4.6505
R11485 VGND.n3925 VGND.n3924 4.6505
R11486 VGND.n3923 VGND.n3922 4.6505
R11487 VGND.n3919 VGND.n3918 4.6505
R11488 VGND.n3917 VGND.n3916 4.6505
R11489 VGND.n3914 VGND.n3913 4.6505
R11490 VGND.n3912 VGND.n3911 4.6505
R11491 VGND.n3910 VGND.n3893 4.6505
R11492 VGND.n3909 VGND.n3908 4.6505
R11493 VGND.n3906 VGND.n3894 4.6505
R11494 VGND.n3905 VGND 4.6505
R11495 VGND.n3903 VGND.n3902 4.6505
R11496 VGND.n3981 VGND.n3980 4.6505
R11497 VGND.n3979 VGND.n3978 4.6505
R11498 VGND.n3977 VGND.n3976 4.6505
R11499 VGND.n3974 VGND.n629 4.6505
R11500 VGND.n3844 VGND.n3843 4.6505
R11501 VGND.n3820 VGND.n3819 4.6505
R11502 VGND.n3818 VGND.n3817 4.6505
R11503 VGND.n3808 VGND.n3807 4.6505
R11504 VGND.n3806 VGND.n3805 4.6505
R11505 VGND.n3763 VGND.n3762 4.6505
R11506 VGND.n3765 VGND.n3764 4.6505
R11507 VGND.n3767 VGND.n3766 4.6505
R11508 VGND.n3769 VGND.n3768 4.6505
R11509 VGND.n3771 VGND.n3770 4.6505
R11510 VGND.n681 VGND.n680 4.6505
R11511 VGND.n685 VGND 4.6505
R11512 VGND.n692 VGND.n691 4.6505
R11513 VGND.n695 VGND.n694 4.6505
R11514 VGND.n696 VGND.n664 4.6505
R11515 VGND.n698 VGND.n697 4.6505
R11516 VGND.n705 VGND.n662 4.6505
R11517 VGND.n707 VGND.n706 4.6505
R11518 VGND.n708 VGND.n661 4.6505
R11519 VGND.n711 VGND.n710 4.6505
R11520 VGND.n712 VGND.n660 4.6505
R11521 VGND.n714 VGND.n713 4.6505
R11522 VGND.n720 VGND.n654 4.6505
R11523 VGND.n727 VGND.n650 4.6505
R11524 VGND.n730 VGND.n649 4.6505
R11525 VGND.n732 VGND.n731 4.6505
R11526 VGND.n734 VGND.n733 4.6505
R11527 VGND.n3761 VGND.n3760 4.6505
R11528 VGND.n3759 VGND.n3758 4.6505
R11529 VGND.n3757 VGND.n3756 4.6505
R11530 VGND.n3754 VGND.n3753 4.6505
R11531 VGND.n3751 VGND.n3750 4.6505
R11532 VGND.n3749 VGND.n3748 4.6505
R11533 VGND.n3745 VGND.n3744 4.6505
R11534 VGND.n3747 VGND.n3746 4.6505
R11535 VGND.n3743 VGND.n3742 4.6505
R11536 VGND.n3734 VGND.n3733 4.6505
R11537 VGND.n3737 VGND.n3736 4.6505
R11538 VGND.n3739 VGND.n3738 4.6505
R11539 VGND.n3741 VGND.n3740 4.6505
R11540 VGND.n3728 VGND.n645 4.6505
R11541 VGND.n3802 VGND.n3801 4.6505
R11542 VGND.n3624 VGND.n759 4.6505
R11543 VGND.n3590 VGND.n766 4.6505
R11544 VGND.n953 VGND.n952 4.6505
R11545 VGND.n849 VGND.n837 4.6505
R11546 VGND.n864 VGND.n863 4.6505
R11547 VGND.n868 VGND.n867 4.6505
R11548 VGND.n876 VGND.n825 4.6505
R11549 VGND.n816 VGND.n815 4.6505
R11550 VGND.n814 VGND.n773 4.6505
R11551 VGND.n813 VGND.n774 4.6505
R11552 VGND.n3623 VGND.n3622 4.6505
R11553 VGND.n3620 VGND.n3619 4.6505
R11554 VGND.n3604 VGND.n3603 4.6505
R11555 VGND.n3598 VGND.n3597 4.6505
R11556 VGND.n3596 VGND.n3595 4.6505
R11557 VGND.n909 VGND.n768 4.6505
R11558 VGND.n913 VGND.n912 4.6505
R11559 VGND.n933 VGND.n932 4.6505
R11560 VGND.n935 VGND.n934 4.6505
R11561 VGND.n938 VGND.n937 4.6505
R11562 VGND.n942 VGND.n941 4.6505
R11563 VGND.n957 VGND.n956 4.6505
R11564 VGND.n959 VGND.n958 4.6505
R11565 VGND.n962 VGND.n961 4.6505
R11566 VGND.n3563 VGND.n3562 4.6505
R11567 VGND.n3559 VGND.n3517 4.6505
R11568 VGND.n3549 VGND.n3548 4.6505
R11569 VGND.n3531 VGND.n3521 4.6505
R11570 VGND.n3478 VGND.n3477 4.6505
R11571 VGND.n3482 VGND.n3481 4.6505
R11572 VGND.n3489 VGND.n3488 4.6505
R11573 VGND.n3492 VGND.n3491 4.6505
R11574 VGND.n3494 VGND.n3493 4.6505
R11575 VGND.n3498 VGND.n3497 4.6505
R11576 VGND.n3501 VGND.n3500 4.6505
R11577 VGND.n3503 VGND.n3502 4.6505
R11578 VGND.n3505 VGND.n3504 4.6505
R11579 VGND VGND.n3506 4.6505
R11580 VGND.n3507 VGND.n887 4.6505
R11581 VGND.n3510 VGND.n3509 4.6505
R11582 VGND.n3572 VGND.n3571 4.6505
R11583 VGND.n3570 VGND.n3569 4.6505
R11584 VGND.n3568 VGND.n3567 4.6505
R11585 VGND.n3565 VGND.n3564 4.6505
R11586 VGND.n3561 VGND.n3560 4.6505
R11587 VGND VGND.n3558 4.6505
R11588 VGND.n3557 VGND.n3556 4.6505
R11589 VGND.n3554 VGND.n3553 4.6505
R11590 VGND.n3551 VGND.n3550 4.6505
R11591 VGND.n3547 VGND.n3546 4.6505
R11592 VGND.n3545 VGND.n3544 4.6505
R11593 VGND.n3543 VGND 4.6505
R11594 VGND.n3542 VGND.n3541 4.6505
R11595 VGND.n3539 VGND.n3538 4.6505
R11596 VGND.n3536 VGND.n3535 4.6505
R11597 VGND.n3534 VGND.n3533 4.6505
R11598 VGND.n3532 VGND.n3520 4.6505
R11599 VGND.n3530 VGND.n3529 4.6505
R11600 VGND.n3528 VGND.n3527 4.6505
R11601 VGND.n3476 VGND.n3475 4.6505
R11602 VGND.n955 VGND.n954 4.6505
R11603 VGND.n949 VGND.n948 4.6505
R11604 VGND.n947 VGND.n946 4.6505
R11605 VGND.n945 VGND.n944 4.6505
R11606 VGND.n940 VGND.n939 4.6505
R11607 VGND.n931 VGND.n930 4.6505
R11608 VGND.n929 VGND.n928 4.6505
R11609 VGND.n927 VGND.n926 4.6505
R11610 VGND.n925 VGND.n924 4.6505
R11611 VGND.n921 VGND.n920 4.6505
R11612 VGND.n3589 VGND.n3588 4.6505
R11613 VGND.n3592 VGND.n763 4.6505
R11614 VGND.n3594 VGND.n3593 4.6505
R11615 VGND.n3602 VGND.n3601 4.6505
R11616 VGND.n3606 VGND.n3605 4.6505
R11617 VGND.n3608 VGND.n3607 4.6505
R11618 VGND.n3610 VGND.n3609 4.6505
R11619 VGND.n3612 VGND.n3611 4.6505
R11620 VGND.n3616 VGND.n3615 4.6505
R11621 VGND.n3618 VGND.n3617 4.6505
R11622 VGND.n844 VGND.n843 4.6505
R11623 VGND.n846 VGND.n845 4.6505
R11624 VGND.n847 VGND.n838 4.6505
R11625 VGND.n848 VGND 4.6505
R11626 VGND.n851 VGND.n850 4.6505
R11627 VGND.n855 VGND.n854 4.6505
R11628 VGND.n858 VGND.n857 4.6505
R11629 VGND.n862 VGND.n861 4.6505
R11630 VGND.n866 VGND.n865 4.6505
R11631 VGND.n870 VGND.n869 4.6505
R11632 VGND.n872 VGND.n871 4.6505
R11633 VGND.n875 VGND.n874 4.6505
R11634 VGND.n824 VGND.n770 4.6505
R11635 VGND.n823 VGND.n822 4.6505
R11636 VGND.n821 VGND.n820 4.6505
R11637 VGND.n818 VGND.n817 4.6505
R11638 VGND.n812 VGND.n811 4.6505
R11639 VGND.n806 VGND.n805 4.6505
R11640 VGND.n804 VGND.n803 4.6505
R11641 VGND.n802 VGND.n801 4.6505
R11642 VGND.n800 VGND.n799 4.6505
R11643 VGND.n798 VGND.n797 4.6505
R11644 VGND.n796 VGND.n795 4.6505
R11645 VGND.n791 VGND.n790 4.6505
R11646 VGND.n789 VGND.n788 4.6505
R11647 VGND.n787 VGND.n786 4.6505
R11648 VGND.n785 VGND.n784 4.6505
R11649 VGND.n3587 VGND.n3586 4.6505
R11650 VGND.n3581 VGND.n3580 4.6505
R11651 VGND.n3583 VGND.n3582 4.6505
R11652 VGND.n3585 VGND.n3584 4.6505
R11653 VGND.n3578 VGND.n3577 4.6505
R11654 VGND.n3576 VGND.n767 4.6505
R11655 VGND.n3222 VGND.n3221 4.6505
R11656 VGND.n3228 VGND.n3227 4.6505
R11657 VGND.n3248 VGND.n3247 4.6505
R11658 VGND.n3272 VGND.n3271 4.6505
R11659 VGND.n3288 VGND.n3287 4.6505
R11660 VGND.n3290 VGND.n3289 4.6505
R11661 VGND.n3292 VGND.n3291 4.6505
R11662 VGND.n3294 VGND.n3293 4.6505
R11663 VGND.n3296 VGND.n3295 4.6505
R11664 VGND.n1064 VGND.n1063 4.6505
R11665 VGND.n1066 VGND.n1065 4.6505
R11666 VGND.n1075 VGND.n1074 4.6505
R11667 VGND.n1075 VGND.n1053 4.6505
R11668 VGND.n1077 VGND.n1076 4.6505
R11669 VGND.n3198 VGND.n1092 4.6505
R11670 VGND.n3190 VGND.n1095 4.6505
R11671 VGND.n3189 VGND.n1096 4.6505
R11672 VGND.n3182 VGND.n1101 4.6505
R11673 VGND.n3174 VGND.n1104 4.6505
R11674 VGND.n3173 VGND.n3172 4.6505
R11675 VGND.n3171 VGND.n1105 4.6505
R11676 VGND.n3224 VGND.n3223 4.6505
R11677 VGND.n3236 VGND.n3235 4.6505
R11678 VGND.n3238 VGND.n3237 4.6505
R11679 VGND.n3240 VGND.n3239 4.6505
R11680 VGND.n3245 VGND.n3244 4.6505
R11681 VGND.n3251 VGND.n3250 4.6505
R11682 VGND.n3255 VGND.n3254 4.6505
R11683 VGND.n3257 VGND.n3256 4.6505
R11684 VGND.n3298 VGND.n3297 4.6505
R11685 VGND.n3300 VGND.n3299 4.6505
R11686 VGND.n3303 VGND.n3302 4.6505
R11687 VGND.n3305 VGND.n3304 4.6505
R11688 VGND.n3309 VGND.n3308 4.6505
R11689 VGND.n3313 VGND.n3312 4.6505
R11690 VGND.n3315 VGND.n3314 4.6505
R11691 VGND.n3317 VGND.n3316 4.6505
R11692 VGND.n3439 VGND.n1022 4.6505
R11693 VGND.n3436 VGND.n1023 4.6505
R11694 VGND.n3412 VGND.n1025 4.6505
R11695 VGND.n3411 VGND.n1026 4.6505
R11696 VGND.n3408 VGND.n1027 4.6505
R11697 VGND.n3403 VGND.n3352 4.6505
R11698 VGND.n3392 VGND.n3353 4.6505
R11699 VGND.n3382 VGND.n3381 4.6505
R11700 VGND.n3362 VGND.n3356 4.6505
R11701 VGND.n3438 VGND.n3437 4.6505
R11702 VGND.n3435 VGND.n3434 4.6505
R11703 VGND.n3433 VGND.n3432 4.6505
R11704 VGND.n3430 VGND.n3429 4.6505
R11705 VGND.n3427 VGND.n3426 4.6505
R11706 VGND.n3425 VGND.n3424 4.6505
R11707 VGND.n3423 VGND.n3422 4.6505
R11708 VGND.n3421 VGND.n3420 4.6505
R11709 VGND.n3419 VGND.n3418 4.6505
R11710 VGND.n3416 VGND.n3415 4.6505
R11711 VGND.n3414 VGND.n3413 4.6505
R11712 VGND.n3410 VGND.n3409 4.6505
R11713 VGND.n3404 VGND.n3350 4.6505
R11714 VGND.n3401 VGND.n3400 4.6505
R11715 VGND.n3398 VGND.n3397 4.6505
R11716 VGND.n3396 VGND.n3395 4.6505
R11717 VGND.n3394 VGND.n3393 4.6505
R11718 VGND.n3391 VGND.n3390 4.6505
R11719 VGND.n3387 VGND.n3386 4.6505
R11720 VGND.n3384 VGND.n3383 4.6505
R11721 VGND.n3380 VGND.n3354 4.6505
R11722 VGND.n3379 VGND.n3378 4.6505
R11723 VGND.n3377 VGND.n3376 4.6505
R11724 VGND.n3375 VGND.n3374 4.6505
R11725 VGND.n3373 VGND.n3372 4.6505
R11726 VGND.n3370 VGND.n3369 4.6505
R11727 VGND.n3368 VGND 4.6505
R11728 VGND.n3367 VGND.n3355 4.6505
R11729 VGND.n3366 VGND.n3365 4.6505
R11730 VGND.n3364 VGND.n3363 4.6505
R11731 VGND.n3448 VGND.n3447 4.6505
R11732 VGND.n3446 VGND.n3445 4.6505
R11733 VGND.n3443 VGND.n3442 4.6505
R11734 VGND.n3441 VGND.n3440 4.6505
R11735 VGND.n3311 VGND.n1033 4.6505
R11736 VGND.n3286 VGND.n1040 4.6505
R11737 VGND.n3283 VGND.n3282 4.6505
R11738 VGND.n3280 VGND.n3279 4.6505
R11739 VGND.n3278 VGND.n3277 4.6505
R11740 VGND.n3276 VGND.n3275 4.6505
R11741 VGND.n3274 VGND.n3273 4.6505
R11742 VGND.n3270 VGND.n3269 4.6505
R11743 VGND.n3266 VGND.n3265 4.6505
R11744 VGND.n3264 VGND.n3263 4.6505
R11745 VGND.n3260 VGND.n3259 4.6505
R11746 VGND VGND.n1044 4.6505
R11747 VGND.n3231 VGND.n3230 4.6505
R11748 VGND.n1059 VGND.n1058 4.6505
R11749 VGND VGND.n1054 4.6505
R11750 VGND.n1068 VGND.n1067 4.6505
R11751 VGND.n1070 VGND.n1069 4.6505
R11752 VGND.n1079 VGND.n1078 4.6505
R11753 VGND.n1081 VGND.n1080 4.6505
R11754 VGND.n1083 VGND.n1082 4.6505
R11755 VGND.n1085 VGND.n1084 4.6505
R11756 VGND.n1090 VGND.n1089 4.6505
R11757 VGND.n3195 VGND.n3194 4.6505
R11758 VGND.n3192 VGND.n3191 4.6505
R11759 VGND.n3187 VGND.n3186 4.6505
R11760 VGND.n3181 VGND.n3180 4.6505
R11761 VGND.n3179 VGND.n3178 4.6505
R11762 VGND.n3176 VGND.n3175 4.6505
R11763 VGND.n3170 VGND.n3169 4.6505
R11764 VGND.n3168 VGND.n3167 4.6505
R11765 VGND.n3166 VGND.n3165 4.6505
R11766 VGND.n3164 VGND.n3163 4.6505
R11767 VGND.n3162 VGND.n3161 4.6505
R11768 VGND.n3160 VGND.n3159 4.6505
R11769 VGND.n3158 VGND.n3157 4.6505
R11770 VGND.n3268 VGND.n3267 4.6505
R11771 VGND.n3056 VGND.n1131 4.6505
R11772 VGND.n3037 VGND.n1133 4.6505
R11773 VGND.n3028 VGND.n1134 4.6505
R11774 VGND.n3025 VGND.n1135 4.6505
R11775 VGND.n2975 VGND.n1258 4.6505
R11776 VGND.n1240 VGND.n1185 4.6505
R11777 VGND.n1232 VGND.n1188 4.6505
R11778 VGND.n1231 VGND.n1189 4.6505
R11779 VGND.n1220 VGND.n1196 4.6505
R11780 VGND.n1219 VGND.n1197 4.6505
R11781 VGND.n3058 VGND.n3057 4.6505
R11782 VGND.n3049 VGND.n3048 4.6505
R11783 VGND.n3047 VGND.n3046 4.6505
R11784 VGND.n3044 VGND.n3043 4.6505
R11785 VGND.n3041 VGND.n3040 4.6505
R11786 VGND.n3003 VGND.n3002 4.6505
R11787 VGND.n3001 VGND.n3000 4.6505
R11788 VGND.n2998 VGND.n2997 4.6505
R11789 VGND.n2995 VGND.n1252 4.6505
R11790 VGND.n2993 VGND.n2992 4.6505
R11791 VGND.n2991 VGND.n2990 4.6505
R11792 VGND.n2988 VGND.n2987 4.6505
R11793 VGND.n2985 VGND 4.6505
R11794 VGND.n2972 VGND.n2971 4.6505
R11795 VGND.n2970 VGND.n2969 4.6505
R11796 VGND.n2968 VGND.n2967 4.6505
R11797 VGND.n2851 VGND.n1276 4.6505
R11798 VGND.n2872 VGND.n2871 4.6505
R11799 VGND.n2874 VGND.n2873 4.6505
R11800 VGND.n2945 VGND.n2944 4.6505
R11801 VGND.n2940 VGND.n2939 4.6505
R11802 VGND.n2938 VGND.n2896 4.6505
R11803 VGND.n2937 VGND.n2897 4.6505
R11804 VGND.n2929 VGND.n2928 4.6505
R11805 VGND.n2923 VGND.n2922 4.6505
R11806 VGND.n2914 VGND.n2905 4.6505
R11807 VGND.n2913 VGND.n2906 4.6505
R11808 VGND.n2912 VGND.n2907 4.6505
R11809 VGND.n2850 VGND.n2849 4.6505
R11810 VGND.n2855 VGND.n2854 4.6505
R11811 VGND.n2859 VGND.n2858 4.6505
R11812 VGND.n2861 VGND.n2860 4.6505
R11813 VGND.n2866 VGND.n2865 4.6505
R11814 VGND.n2868 VGND.n2867 4.6505
R11815 VGND.n2870 VGND.n2869 4.6505
R11816 VGND.n2876 VGND.n2875 4.6505
R11817 VGND.n2878 VGND.n2877 4.6505
R11818 VGND.n2879 VGND.n1274 4.6505
R11819 VGND.n2882 VGND.n2881 4.6505
R11820 VGND.n2885 VGND.n2884 4.6505
R11821 VGND.n2888 VGND.n2887 4.6505
R11822 VGND.n2893 VGND.n2892 4.6505
R11823 VGND.n2942 VGND.n2941 4.6505
R11824 VGND.n2936 VGND.n2935 4.6505
R11825 VGND.n2934 VGND.n2898 4.6505
R11826 VGND.n2933 VGND.n2932 4.6505
R11827 VGND.n2931 VGND.n2930 4.6505
R11828 VGND.n2927 VGND.n2900 4.6505
R11829 VGND.n2926 VGND.n2925 4.6505
R11830 VGND.n2924 VGND.n2901 4.6505
R11831 VGND.n2921 VGND.n2902 4.6505
R11832 VGND.n2920 VGND.n2919 4.6505
R11833 VGND.n2918 VGND.n2903 4.6505
R11834 VGND.n2916 VGND.n2915 4.6505
R11835 VGND VGND.n2904 4.6505
R11836 VGND.n2911 VGND.n2910 4.6505
R11837 VGND.n2974 VGND.n2973 4.6505
R11838 VGND.n2977 VGND.n2976 4.6505
R11839 VGND.n2979 VGND.n2978 4.6505
R11840 VGND.n2982 VGND.n2981 4.6505
R11841 VGND.n2984 VGND.n2983 4.6505
R11842 VGND.n2996 VGND 4.6505
R11843 VGND.n3005 VGND.n3004 4.6505
R11844 VGND.n3010 VGND.n3009 4.6505
R11845 VGND.n3012 VGND.n1138 4.6505
R11846 VGND.n3016 VGND.n3015 4.6505
R11847 VGND.n3019 VGND.n3018 4.6505
R11848 VGND.n3022 VGND.n3021 4.6505
R11849 VGND.n3024 VGND.n3023 4.6505
R11850 VGND.n3027 VGND.n3026 4.6505
R11851 VGND.n3030 VGND.n3029 4.6505
R11852 VGND.n3032 VGND.n3031 4.6505
R11853 VGND.n3034 VGND.n3033 4.6505
R11854 VGND.n3036 VGND.n3035 4.6505
R11855 VGND.n3039 VGND.n3038 4.6505
R11856 VGND.n3051 VGND.n3050 4.6505
R11857 VGND.n3053 VGND.n3052 4.6505
R11858 VGND.n3055 VGND.n3054 4.6505
R11859 VGND.n1154 VGND.n1153 4.6505
R11860 VGND.n1156 VGND.n1155 4.6505
R11861 VGND VGND.n1159 4.6505
R11862 VGND.n1162 VGND.n1161 4.6505
R11863 VGND.n1163 VGND.n1147 4.6505
R11864 VGND.n1165 VGND.n1164 4.6505
R11865 VGND.n1167 VGND.n1166 4.6505
R11866 VGND.n1168 VGND.n1145 4.6505
R11867 VGND.n1170 VGND.n1169 4.6505
R11868 VGND.n1171 VGND.n1144 4.6505
R11869 VGND.n1173 VGND.n1172 4.6505
R11870 VGND.n1174 VGND.n1143 4.6505
R11871 VGND.n1176 VGND.n1175 4.6505
R11872 VGND.n1177 VGND.n1142 4.6505
R11873 VGND.n1179 VGND.n1178 4.6505
R11874 VGND.n1180 VGND.n1141 4.6505
R11875 VGND.n1183 VGND.n1182 4.6505
R11876 VGND.n1184 VGND.n1140 4.6505
R11877 VGND.n1239 VGND.n1238 4.6505
R11878 VGND.n1237 VGND.n1186 4.6505
R11879 VGND.n1236 VGND.n1235 4.6505
R11880 VGND.n1233 VGND.n1187 4.6505
R11881 VGND.n1230 VGND.n1229 4.6505
R11882 VGND.n1228 VGND.n1190 4.6505
R11883 VGND.n1227 VGND.n1226 4.6505
R11884 VGND.n1225 VGND.n1191 4.6505
R11885 VGND.n1224 VGND.n1223 4.6505
R11886 VGND.n1218 VGND.n1217 4.6505
R11887 VGND.n1216 VGND.n1198 4.6505
R11888 VGND.n1213 VGND.n1199 4.6505
R11889 VGND.n1212 VGND.n1211 4.6505
R11890 VGND.n1210 VGND.n1200 4.6505
R11891 VGND.n1209 VGND.n1208 4.6505
R11892 VGND.n1207 VGND.n1206 4.6505
R11893 VGND.n1205 VGND.n1204 4.6505
R11894 VGND.n1203 VGND.n1202 4.6505
R11895 VGND.n3014 VGND.n3013 4.6505
R11896 VGND.n2627 VGND.n2578 4.6505
R11897 VGND.n2607 VGND.n2588 4.6505
R11898 VGND.n2606 VGND.n2589 4.6505
R11899 VGND.n2654 VGND.n2653 4.6505
R11900 VGND.n2672 VGND.n2671 4.6505
R11901 VGND.n2690 VGND.n2689 4.6505
R11902 VGND.n1404 VGND.n1403 4.6505
R11903 VGND.n1417 VGND.n1416 4.6505
R11904 VGND.n1421 VGND.n1420 4.6505
R11905 VGND.n1437 VGND.n1436 4.6505
R11906 VGND.n1441 VGND.n1440 4.6505
R11907 VGND.n2626 VGND.n2625 4.6505
R11908 VGND.n2604 VGND.n2603 4.6505
R11909 VGND.n2600 VGND.n2599 4.6505
R11910 VGND.n2598 VGND.n2595 4.6505
R11911 VGND.n2686 VGND.n2685 4.6505
R11912 VGND.n2692 VGND.n2691 4.6505
R11913 VGND.n2694 VGND.n2693 4.6505
R11914 VGND.n2697 VGND.n2696 4.6505
R11915 VGND.n2818 VGND.n1322 4.6505
R11916 VGND.n2817 VGND.n1324 4.6505
R11917 VGND.n2810 VGND.n1325 4.6505
R11918 VGND.n2807 VGND.n1326 4.6505
R11919 VGND.n2806 VGND.n1327 4.6505
R11920 VGND.n2787 VGND.n2736 4.6505
R11921 VGND.n2780 VGND.n2738 4.6505
R11922 VGND.n2775 VGND.n2739 4.6505
R11923 VGND.n2752 VGND.n2740 4.6505
R11924 VGND.n2747 VGND.n2741 4.6505
R11925 VGND.n2820 VGND.n2819 4.6505
R11926 VGND.n2816 VGND.n2815 4.6505
R11927 VGND.n2814 VGND.n2813 4.6505
R11928 VGND.n2812 VGND.n2811 4.6505
R11929 VGND.n2809 VGND.n2808 4.6505
R11930 VGND.n2804 VGND.n2803 4.6505
R11931 VGND.n2796 VGND.n2795 4.6505
R11932 VGND.n2794 VGND.n1332 4.6505
R11933 VGND.n2792 VGND.n2791 4.6505
R11934 VGND.n2789 VGND.n2788 4.6505
R11935 VGND.n2783 VGND.n2782 4.6505
R11936 VGND.n2779 VGND.n2778 4.6505
R11937 VGND.n2777 VGND.n2776 4.6505
R11938 VGND.n2774 VGND.n2773 4.6505
R11939 VGND.n2770 VGND.n2769 4.6505
R11940 VGND.n2768 VGND.n2767 4.6505
R11941 VGND.n2766 VGND.n2765 4.6505
R11942 VGND.n2763 VGND.n2762 4.6505
R11943 VGND.n2758 VGND.n2757 4.6505
R11944 VGND.n2755 VGND.n2754 4.6505
R11945 VGND.n2753 VGND 4.6505
R11946 VGND.n2751 VGND.n2750 4.6505
R11947 VGND.n2749 VGND.n2748 4.6505
R11948 VGND.n2825 VGND.n2824 4.6505
R11949 VGND.n2821 VGND.n2820 4.6505
R11950 VGND.n2688 VGND.n2687 4.6505
R11951 VGND.n2684 VGND.n2683 4.6505
R11952 VGND.n2682 VGND.n2681 4.6505
R11953 VGND.n2680 VGND.n2679 4.6505
R11954 VGND.n2678 VGND.n2677 4.6505
R11955 VGND.n2676 VGND.n2675 4.6505
R11956 VGND.n2674 VGND.n2673 4.6505
R11957 VGND.n2670 VGND.n2669 4.6505
R11958 VGND.n2668 VGND.n2667 4.6505
R11959 VGND.n2666 VGND.n2665 4.6505
R11960 VGND.n2664 VGND.n1337 4.6505
R11961 VGND.n2662 VGND.n2661 4.6505
R11962 VGND.n2660 VGND.n2659 4.6505
R11963 VGND.n2658 VGND.n2657 4.6505
R11964 VGND.n2656 VGND.n2655 4.6505
R11965 VGND.n2596 VGND.n1340 4.6505
R11966 VGND.n2608 VGND.n2587 4.6505
R11967 VGND.n2610 VGND.n2609 4.6505
R11968 VGND.n2612 VGND.n2611 4.6505
R11969 VGND.n2617 VGND.n2616 4.6505
R11970 VGND.n2619 VGND.n2618 4.6505
R11971 VGND.n2620 VGND.n2580 4.6505
R11972 VGND.n1368 VGND.n1365 4.6505
R11973 VGND.n1370 VGND.n1369 4.6505
R11974 VGND.n1373 VGND.n1363 4.6505
R11975 VGND.n1375 VGND.n1374 4.6505
R11976 VGND.n1378 VGND.n1377 4.6505
R11977 VGND.n1380 VGND.n1379 4.6505
R11978 VGND.n1381 VGND.n1360 4.6505
R11979 VGND.n1383 VGND.n1382 4.6505
R11980 VGND.n1385 VGND.n1384 4.6505
R11981 VGND.n1386 VGND.n1358 4.6505
R11982 VGND.n1388 VGND.n1387 4.6505
R11983 VGND.n1389 VGND.n1357 4.6505
R11984 VGND.n1391 VGND.n1390 4.6505
R11985 VGND.n1392 VGND.n1356 4.6505
R11986 VGND.n1394 VGND.n1393 4.6505
R11987 VGND.n1395 VGND.n1355 4.6505
R11988 VGND.n1397 VGND.n1396 4.6505
R11989 VGND.n1398 VGND.n1354 4.6505
R11990 VGND.n1401 VGND.n1400 4.6505
R11991 VGND.n1402 VGND.n1351 4.6505
R11992 VGND.n1405 VGND.n1350 4.6505
R11993 VGND.n1407 VGND.n1406 4.6505
R11994 VGND.n1410 VGND.n1409 4.6505
R11995 VGND.n1411 VGND.n1348 4.6505
R11996 VGND.n1414 VGND.n1413 4.6505
R11997 VGND.n1419 VGND.n1418 4.6505
R11998 VGND.n1423 VGND.n1422 4.6505
R11999 VGND.n1425 VGND.n1424 4.6505
R12000 VGND.n1427 VGND.n1426 4.6505
R12001 VGND.n1429 VGND.n1428 4.6505
R12002 VGND.n1431 VGND.n1430 4.6505
R12003 VGND.n1433 VGND.n1432 4.6505
R12004 VGND.n1435 VGND.n1346 4.6505
R12005 VGND.n1439 VGND.n1438 4.6505
R12006 VGND.n1443 VGND.n1442 4.6505
R12007 VGND.n1445 VGND.n1444 4.6505
R12008 VGND.n1448 VGND.n1447 4.6505
R12009 VGND.n2652 VGND.n2651 4.6505
R12010 VGND.n2649 VGND.n2648 4.6505
R12011 VGND.n2275 VGND.n2274 4.6505
R12012 VGND.n2301 VGND.n2300 4.6505
R12013 VGND.n2330 VGND.n2329 4.6505
R12014 VGND.n2332 VGND.n1485 4.6505
R12015 VGND.n2343 VGND.n2342 4.6505
R12016 VGND.n2140 VGND 4.6505
R12017 VGND.n2147 VGND.n2127 4.6505
R12018 VGND.n2147 VGND.n2126 4.6505
R12019 VGND.n2199 VGND.n2176 4.6505
R12020 VGND.n2196 VGND.n2177 4.6505
R12021 VGND.n2278 VGND.n2277 4.6505
R12022 VGND.n2279 VGND.n1495 4.6505
R12023 VGND.n2281 VGND.n2280 4.6505
R12024 VGND.n2287 VGND.n1494 4.6505
R12025 VGND.n2289 VGND.n2288 4.6505
R12026 VGND.n2292 VGND.n2291 4.6505
R12027 VGND.n2295 VGND.n2294 4.6505
R12028 VGND.n2298 VGND.n2297 4.6505
R12029 VGND.n2305 VGND.n2304 4.6505
R12030 VGND.n2306 VGND.n1489 4.6505
R12031 VGND.n2320 VGND.n2319 4.6505
R12032 VGND.n2336 VGND.n2335 4.6505
R12033 VGND.n2338 VGND.n2337 4.6505
R12034 VGND.n2340 VGND.n2339 4.6505
R12035 VGND.n2353 VGND.n2352 4.6505
R12036 VGND.n2357 VGND.n2356 4.6505
R12037 VGND.n2359 VGND.n2358 4.6505
R12038 VGND.n2362 VGND.n2361 4.6505
R12039 VGND.n2500 VGND.n1464 4.6505
R12040 VGND.n2497 VGND.n1465 4.6505
R12041 VGND.n2496 VGND.n1466 4.6505
R12042 VGND.n2495 VGND.n1467 4.6505
R12043 VGND.n2492 VGND.n2491 4.6505
R12044 VGND.n2456 VGND.n2411 4.6505
R12045 VGND.n2507 VGND.n2506 4.6505
R12046 VGND.n2505 VGND.n2504 4.6505
R12047 VGND.n2503 VGND.n2502 4.6505
R12048 VGND.n2499 VGND.n2498 4.6505
R12049 VGND.n2494 VGND.n2493 4.6505
R12050 VGND.n2490 VGND.n1470 4.6505
R12051 VGND.n2487 VGND.n2486 4.6505
R12052 VGND.n2485 VGND.n2484 4.6505
R12053 VGND.n2482 VGND.n2481 4.6505
R12054 VGND VGND.n2478 4.6505
R12055 VGND.n2477 VGND.n2476 4.6505
R12056 VGND.n2474 VGND.n2473 4.6505
R12057 VGND.n2471 VGND.n2470 4.6505
R12058 VGND.n2469 VGND.n2468 4.6505
R12059 VGND.n2467 VGND.n2410 4.6505
R12060 VGND.n2465 VGND.n2464 4.6505
R12061 VGND.n2462 VGND.n2461 4.6505
R12062 VGND.n2460 VGND.n2459 4.6505
R12063 VGND.n2458 VGND.n2457 4.6505
R12064 VGND VGND.n2455 4.6505
R12065 VGND.n2454 VGND.n2453 4.6505
R12066 VGND.n2452 VGND.n2413 4.6505
R12067 VGND.n2450 VGND.n2449 4.6505
R12068 VGND.n2448 VGND.n2447 4.6505
R12069 VGND.n2446 VGND.n2445 4.6505
R12070 VGND.n2443 VGND.n2442 4.6505
R12071 VGND.n2441 VGND.n2416 4.6505
R12072 VGND.n2440 VGND.n2439 4.6505
R12073 VGND.n2436 VGND 4.6505
R12074 VGND.n2435 VGND.n2420 4.6505
R12075 VGND.n2433 VGND.n2432 4.6505
R12076 VGND.n2431 VGND.n2430 4.6505
R12077 VGND.n2429 VGND.n2423 4.6505
R12078 VGND.n2427 VGND.n2426 4.6505
R12079 VGND.n2355 VGND.n2354 4.6505
R12080 VGND.n2351 VGND.n2350 4.6505
R12081 VGND.n2349 VGND.n1481 4.6505
R12082 VGND.n2347 VGND.n2346 4.6505
R12083 VGND.n2345 VGND.n2344 4.6505
R12084 VGND.n2334 VGND.n2333 4.6505
R12085 VGND.n2328 VGND.n2327 4.6505
R12086 VGND.n2326 VGND.n2325 4.6505
R12087 VGND.n2324 VGND.n2323 4.6505
R12088 VGND.n2285 VGND.n2284 4.6505
R12089 VGND.n2137 VGND.n2136 4.6505
R12090 VGND.n2143 VGND.n2142 4.6505
R12091 VGND.n2149 VGND.n2148 4.6505
R12092 VGND.n2151 VGND.n2150 4.6505
R12093 VGND.n2152 VGND.n2125 4.6505
R12094 VGND.n2154 VGND.n2153 4.6505
R12095 VGND.n2156 VGND.n2155 4.6505
R12096 VGND.n2158 VGND.n2157 4.6505
R12097 VGND.n2160 VGND.n2159 4.6505
R12098 VGND.n2168 VGND.n2167 4.6505
R12099 VGND.n2223 VGND.n2222 4.6505
R12100 VGND.n2221 VGND.n2220 4.6505
R12101 VGND.n2217 VGND.n2216 4.6505
R12102 VGND.n2214 VGND.n2213 4.6505
R12103 VGND.n2212 VGND.n2211 4.6505
R12104 VGND.n2209 VGND.n2208 4.6505
R12105 VGND.n2206 VGND.n2205 4.6505
R12106 VGND.n2204 VGND.n2172 4.6505
R12107 VGND.n2203 VGND.n2202 4.6505
R12108 VGND.n2198 VGND.n2197 4.6505
R12109 VGND.n2195 VGND.n2194 4.6505
R12110 VGND.n2193 VGND.n2192 4.6505
R12111 VGND.n2190 VGND.n2189 4.6505
R12112 VGND.n2187 VGND.n2186 4.6505
R12113 VGND.n2185 VGND.n2179 4.6505
R12114 VGND.n2184 VGND.n2183 4.6505
R12115 VGND.n2308 VGND.n2307 4.6505
R12116 VGND.n2311 VGND.n2310 4.6505
R12117 VGND.n2317 VGND.n1487 4.6505
R12118 VGND.n2317 VGND.n2316 4.6505
R12119 VGND.n2055 VGND.n1521 4.6505
R12120 VGND.n2036 VGND.n1527 4.6505
R12121 VGND.n2031 VGND.n1530 4.6505
R12122 VGND.n2030 VGND.n1531 4.6505
R12123 VGND.n1758 VGND.n1532 4.6505
R12124 VGND.n1765 VGND.n1764 4.6505
R12125 VGND.n1775 VGND.n1774 4.6505
R12126 VGND.n1777 VGND.n1776 4.6505
R12127 VGND.n1779 VGND.n1778 4.6505
R12128 VGND.n1784 VGND.n1753 4.6505
R12129 VGND.n1790 VGND.n1789 4.6505
R12130 VGND.n1796 VGND.n1795 4.6505
R12131 VGND.n1598 VGND.n1593 4.6505
R12132 VGND.n1600 VGND.n1599 4.6505
R12133 VGND.n1602 VGND.n1601 4.6505
R12134 VGND.n1589 VGND.n1539 4.6505
R12135 VGND.n1565 VGND.n1549 4.6505
R12136 VGND.n2054 VGND.n2053 4.6505
R12137 VGND.n2050 VGND.n2049 4.6505
R12138 VGND.n2048 VGND.n2047 4.6505
R12139 VGND.n2045 VGND.n1522 4.6505
R12140 VGND.n2044 VGND.n2043 4.6505
R12141 VGND.n2040 VGND.n2039 4.6505
R12142 VGND.n2034 VGND.n2033 4.6505
R12143 VGND.n1786 VGND.n1785 4.6505
R12144 VGND.n1800 VGND.n1799 4.6505
R12145 VGND.n1802 VGND.n1801 4.6505
R12146 VGND.n1805 VGND.n1804 4.6505
R12147 VGND.n1734 VGND.n1733 4.6505
R12148 VGND.n1731 VGND.n1644 4.6505
R12149 VGND VGND.n1645 4.6505
R12150 VGND.n1726 VGND.n1725 4.6505
R12151 VGND.n1724 VGND.n1648 4.6505
R12152 VGND.n1723 VGND.n1649 4.6505
R12153 VGND.n1722 VGND.n1650 4.6505
R12154 VGND.n1717 VGND.n1716 4.6505
R12155 VGND.n1713 VGND.n1653 4.6505
R12156 VGND.n1704 VGND.n1703 4.6505
R12157 VGND.n1697 VGND.n1659 4.6505
R12158 VGND.n1671 VGND 4.6505
R12159 VGND.n1670 VGND.n1660 4.6505
R12160 VGND.n1729 VGND.n1728 4.6505
R12161 VGND.n1720 VGND.n1719 4.6505
R12162 VGND.n1715 VGND.n1714 4.6505
R12163 VGND.n1712 VGND.n1711 4.6505
R12164 VGND.n1707 VGND.n1706 4.6505
R12165 VGND.n1702 VGND.n1656 4.6505
R12166 VGND.n1700 VGND.n1699 4.6505
R12167 VGND.n1696 VGND.n1695 4.6505
R12168 VGND.n1694 VGND.n1693 4.6505
R12169 VGND.n1692 VGND.n1691 4.6505
R12170 VGND.n1690 VGND.n1689 4.6505
R12171 VGND.n1688 VGND.n1687 4.6505
R12172 VGND.n1686 VGND.n1685 4.6505
R12173 VGND.n1684 VGND.n1683 4.6505
R12174 VGND.n1681 VGND.n1680 4.6505
R12175 VGND.n1676 VGND.n1675 4.6505
R12176 VGND.n1673 VGND.n1672 4.6505
R12177 VGND.n1669 VGND.n1668 4.6505
R12178 VGND.n1741 VGND.n1740 4.6505
R12179 VGND.n1739 VGND.n1738 4.6505
R12180 VGND.n1736 VGND.n1735 4.6505
R12181 VGND.n1732 VGND.n1643 4.6505
R12182 VGND.n1798 VGND.n1797 4.6505
R12183 VGND.n1794 VGND.n1793 4.6505
R12184 VGND.n1792 VGND.n1791 4.6505
R12185 VGND.n1788 VGND.n1787 4.6505
R12186 VGND.n1782 VGND.n1781 4.6505
R12187 VGND.n1773 VGND.n1772 4.6505
R12188 VGND.n1771 VGND.n1770 4.6505
R12189 VGND.n1769 VGND.n1768 4.6505
R12190 VGND.n1767 VGND.n1766 4.6505
R12191 VGND.n1763 VGND.n1762 4.6505
R12192 VGND.n1760 VGND.n1759 4.6505
R12193 VGND.n2020 VGND.n2019 4.6505
R12194 VGND.n2022 VGND.n2021 4.6505
R12195 VGND.n2025 VGND.n2024 4.6505
R12196 VGND.n2029 VGND.n2028 4.6505
R12197 VGND.n2038 VGND.n1524 4.6505
R12198 VGND VGND.n1603 4.6505
R12199 VGND.n1612 VGND.n1611 4.6505
R12200 VGND.n1615 VGND.n1614 4.6505
R12201 VGND.n1619 VGND.n1618 4.6505
R12202 VGND.n1621 VGND.n1620 4.6505
R12203 VGND.n1623 VGND.n1622 4.6505
R12204 VGND.n1626 VGND.n1538 4.6505
R12205 VGND.n1627 VGND.n1534 4.6505
R12206 VGND.n1628 VGND.n1534 4.6505
R12207 VGND.n1587 VGND.n1586 4.6505
R12208 VGND.n1581 VGND.n1580 4.6505
R12209 VGND.n1579 VGND.n1578 4.6505
R12210 VGND.n1575 VGND.n1574 4.6505
R12211 VGND.n1573 VGND.n1572 4.6505
R12212 VGND.n1564 VGND.n1563 4.6505
R12213 VGND.n1562 VGND.n1561 4.6505
R12214 VGND.n1560 VGND.n1559 4.6505
R12215 VGND.n1558 VGND.n1557 4.6505
R12216 VGND.n1556 VGND.n1555 4.6505
R12217 VGND.n1554 VGND.n1553 4.6505
R12218 VGND.n1552 VGND.n1551 4.6505
R12219 VGND.n5132 VGND.n99 4.6505
R12220 VGND.n5119 VGND.n101 4.6505
R12221 VGND.n5106 VGND.n5105 4.6505
R12222 VGND.n5096 VGND.n103 4.6505
R12223 VGND.n5095 VGND.n104 4.6505
R12224 VGND.n5094 VGND.n105 4.6505
R12225 VGND.n5088 VGND.n107 4.6505
R12226 VGND.n5080 VGND.n110 4.6505
R12227 VGND.n5077 VGND.n111 4.6505
R12228 VGND.n5067 VGND.n114 4.6505
R12229 VGND.n5060 VGND.n115 4.6505
R12230 VGND.n188 VGND.n176 4.6505
R12231 VGND.n187 VGND.n177 4.6505
R12232 VGND.n186 VGND.n178 4.6505
R12233 VGND.n5131 VGND.n5130 4.6505
R12234 VGND.n5128 VGND.n5127 4.6505
R12235 VGND.n5085 VGND.n5084 4.6505
R12236 VGND.n5057 VGND.n5056 4.6505
R12237 VGND.n5055 VGND.n5054 4.6505
R12238 VGND.n5053 VGND.n5052 4.6505
R12239 VGND.n5051 VGND.n5050 4.6505
R12240 VGND.n5049 VGND.n5048 4.6505
R12241 VGND.n5046 VGND.n5045 4.6505
R12242 VGND.n5041 VGND.n5040 4.6505
R12243 VGND.n1959 VGND.n1867 4.6505
R12244 VGND.n1943 VGND.n1942 4.6505
R12245 VGND.n1941 VGND.n1875 4.6505
R12246 VGND.n1928 VGND.n126 4.6505
R12247 VGND.n1916 VGND.n1876 4.6505
R12248 VGND.n1913 VGND.n1877 4.6505
R12249 VGND VGND.n1882 4.6505
R12250 VGND.n1899 VGND.n1884 4.6505
R12251 VGND.n1897 VGND.n1885 4.6505
R12252 VGND.n1967 VGND.n1966 4.6505
R12253 VGND.n1964 VGND.n1963 4.6505
R12254 VGND.n1962 VGND.n1961 4.6505
R12255 VGND.n1960 VGND.n1866 4.6505
R12256 VGND.n1958 VGND.n1957 4.6505
R12257 VGND.n1951 VGND.n1950 4.6505
R12258 VGND.n1949 VGND.n1948 4.6505
R12259 VGND.n1945 VGND.n1944 4.6505
R12260 VGND.n1940 VGND.n1939 4.6505
R12261 VGND.n1936 VGND.n1935 4.6505
R12262 VGND.n1934 VGND.n1933 4.6505
R12263 VGND.n1932 VGND.n1931 4.6505
R12264 VGND.n1930 VGND.n1929 4.6505
R12265 VGND.n1927 VGND.n1926 4.6505
R12266 VGND.n1923 VGND.n1922 4.6505
R12267 VGND.n1920 VGND.n1919 4.6505
R12268 VGND.n1918 VGND.n1917 4.6505
R12269 VGND.n1915 VGND.n1914 4.6505
R12270 VGND.n1912 VGND.n1911 4.6505
R12271 VGND.n1910 VGND.n1909 4.6505
R12272 VGND.n1908 VGND.n1907 4.6505
R12273 VGND.n1906 VGND.n1905 4.6505
R12274 VGND.n1904 VGND.n1879 4.6505
R12275 VGND.n1902 VGND.n1901 4.6505
R12276 VGND.n1894 VGND.n1893 4.6505
R12277 VGND.n1892 VGND.n1891 4.6505
R12278 VGND.n1977 VGND.n1976 4.6505
R12279 VGND.n1975 VGND.n1974 4.6505
R12280 VGND.n1972 VGND.n1971 4.6505
R12281 VGND.n1970 VGND.n1969 4.6505
R12282 VGND.n5059 VGND.n5058 4.6505
R12283 VGND.n5062 VGND.n5061 4.6505
R12284 VGND.n5064 VGND.n5063 4.6505
R12285 VGND.n5066 VGND.n5065 4.6505
R12286 VGND.n5069 VGND.n5068 4.6505
R12287 VGND.n5071 VGND.n5070 4.6505
R12288 VGND.n5074 VGND.n5073 4.6505
R12289 VGND.n5076 VGND.n5075 4.6505
R12290 VGND.n5079 VGND.n5078 4.6505
R12291 VGND.n5083 VGND.n5082 4.6505
R12292 VGND.n5087 VGND.n5086 4.6505
R12293 VGND.n5093 VGND.n5092 4.6505
R12294 VGND.n5098 VGND.n5097 4.6505
R12295 VGND.n5100 VGND.n5099 4.6505
R12296 VGND.n5102 VGND.n5101 4.6505
R12297 VGND.n5104 VGND.n5103 4.6505
R12298 VGND.n5108 VGND.n5107 4.6505
R12299 VGND.n5111 VGND.n5110 4.6505
R12300 VGND.n5114 VGND.n5113 4.6505
R12301 VGND.n5116 VGND.n5115 4.6505
R12302 VGND.n5118 VGND.n5117 4.6505
R12303 VGND.n5121 VGND.n5120 4.6505
R12304 VGND.n5123 VGND.n5122 4.6505
R12305 VGND.n5126 VGND.n5125 4.6505
R12306 VGND.n140 VGND.n139 4.6505
R12307 VGND.n144 VGND.n143 4.6505
R12308 VGND.n146 VGND.n145 4.6505
R12309 VGND.n148 VGND.n147 4.6505
R12310 VGND.n152 VGND.n150 4.6505
R12311 VGND.n158 VGND.n157 4.6505
R12312 VGND.n161 VGND.n160 4.6505
R12313 VGND.n163 VGND.n162 4.6505
R12314 VGND.n165 VGND.n164 4.6505
R12315 VGND.n211 VGND.n210 4.6505
R12316 VGND.n209 VGND.n129 4.6505
R12317 VGND.n199 VGND.n170 4.6505
R12318 VGND.n198 VGND.n197 4.6505
R12319 VGND.n196 VGND.n195 4.6505
R12320 VGND.n191 VGND.n190 4.6505
R12321 VGND.n190 VGND.n189 4.6505
R12322 VGND.n185 VGND.n184 4.6505
R12323 VGND.n183 VGND.n182 4.6505
R12324 VGND.n181 VGND.n180 4.6505
R12325 VGND.n4228 VGND.n4227 4.6505
R12326 VGND.n4230 VGND.n4229 4.6505
R12327 VGND.n4232 VGND.n4231 4.6505
R12328 VGND.n4237 VGND.n4221 4.6505
R12329 VGND.n4239 VGND.n4238 4.6505
R12330 VGND.n4241 VGND.n4240 4.6505
R12331 VGND.n4242 VGND.n4220 4.6505
R12332 VGND VGND.n4208 4.6505
R12333 VGND.n4290 VGND.n4289 4.6505
R12334 VGND.n4292 VGND.n4291 4.6505
R12335 VGND.n4294 VGND.n4293 4.6505
R12336 VGND.n4296 VGND.n250 4.6505
R12337 VGND.n4456 VGND.n4308 4.6505
R12338 VGND.n4446 VGND.n4445 4.6505
R12339 VGND.n4439 VGND.n4312 4.6505
R12340 VGND.n4438 VGND.n4313 4.6505
R12341 VGND.n4437 VGND.n4314 4.6505
R12342 VGND.n4432 VGND.n4315 4.6505
R12343 VGND.n4412 VGND.n252 4.6505
R12344 VGND.n4404 VGND.n4319 4.6505
R12345 VGND.n4398 VGND.n4397 4.6505
R12346 VGND.n4395 VGND.n4323 4.6505
R12347 VGND.n4888 VGND.n4887 4.6505
R12348 VGND.n4909 VGND 4.6505
R12349 VGND.n4911 VGND.n4910 4.6505
R12350 VGND.n4913 VGND.n4912 4.6505
R12351 VGND.n4915 VGND.n4914 4.6505
R12352 VGND.n4963 VGND.n4917 4.6505
R12353 VGND.n4962 VGND.n4918 4.6505
R12354 VGND.n4961 VGND.n4919 4.6505
R12355 VGND VGND.n4920 4.6505
R12356 VGND.n4455 VGND.n4454 4.6505
R12357 VGND.n4453 VGND.n4452 4.6505
R12358 VGND.n4451 VGND.n4450 4.6505
R12359 VGND.n4448 VGND.n4447 4.6505
R12360 VGND.n4444 VGND.n4311 4.6505
R12361 VGND.n4443 VGND.n4442 4.6505
R12362 VGND.n4441 VGND.n4440 4.6505
R12363 VGND.n4436 VGND.n4435 4.6505
R12364 VGND.n4434 VGND.n4433 4.6505
R12365 VGND.n4431 VGND.n4430 4.6505
R12366 VGND.n4429 VGND.n4428 4.6505
R12367 VGND.n4427 VGND.n4426 4.6505
R12368 VGND.n4425 VGND.n4424 4.6505
R12369 VGND.n4421 VGND.n4420 4.6505
R12370 VGND.n4413 VGND.n251 4.6505
R12371 VGND.n4411 VGND.n4410 4.6505
R12372 VGND.n4406 VGND.n4316 4.6505
R12373 VGND.n4403 VGND.n4402 4.6505
R12374 VGND.n4400 VGND.n4399 4.6505
R12375 VGND.n4396 VGND.n4322 4.6505
R12376 VGND.n4394 VGND.n4393 4.6505
R12377 VGND.n4392 VGND.n4391 4.6505
R12378 VGND.n4389 VGND.n4388 4.6505
R12379 VGND.n4387 VGND.n4386 4.6505
R12380 VGND.n4385 VGND.n4326 4.6505
R12381 VGND.n4384 VGND.n4383 4.6505
R12382 VGND.n4382 VGND.n4381 4.6505
R12383 VGND.n4380 VGND.n4379 4.6505
R12384 VGND.n4378 VGND.n4377 4.6505
R12385 VGND.n4376 VGND.n4375 4.6505
R12386 VGND.n4373 VGND.n4372 4.6505
R12387 VGND.n4890 VGND.n4889 4.6505
R12388 VGND.n4892 VGND.n4891 4.6505
R12389 VGND.n4894 VGND.n4893 4.6505
R12390 VGND.n4896 VGND.n4895 4.6505
R12391 VGND.n4898 VGND.n4897 4.6505
R12392 VGND.n4899 VGND.n258 4.6505
R12393 VGND.n4901 VGND.n4900 4.6505
R12394 VGND.n4904 VGND.n4903 4.6505
R12395 VGND.n4907 VGND.n4906 4.6505
R12396 VGND.n4960 VGND.n4959 4.6505
R12397 VGND.n4956 VGND.n4955 4.6505
R12398 VGND.n4954 VGND.n4953 4.6505
R12399 VGND.n4952 VGND.n4951 4.6505
R12400 VGND.n4949 VGND.n4948 4.6505
R12401 VGND.n4944 VGND.n4943 4.6505
R12402 VGND.n4941 VGND.n4940 4.6505
R12403 VGND.n4939 VGND 4.6505
R12404 VGND.n4938 VGND.n4923 4.6505
R12405 VGND.n4936 VGND.n4935 4.6505
R12406 VGND.n4934 VGND.n4933 4.6505
R12407 VGND.n4932 VGND.n4926 4.6505
R12408 VGND.n4461 VGND.n4460 4.6505
R12409 VGND.n4458 VGND.n4457 4.6505
R12410 VGND VGND.n4233 4.6505
R12411 VGND.n4243 VGND 4.6505
R12412 VGND.n4245 VGND.n4244 4.6505
R12413 VGND.n4247 VGND.n4246 4.6505
R12414 VGND.n4249 VGND.n4248 4.6505
R12415 VGND.n4254 VGND.n4253 4.6505
R12416 VGND.n4252 VGND.n248 4.6505
R12417 VGND.n4258 VGND.n4257 4.6505
R12418 VGND.n4259 VGND.n249 4.6505
R12419 VGND.n4263 VGND.n4262 4.6505
R12420 VGND.n4265 VGND.n4214 4.6505
R12421 VGND.n4266 VGND 4.6505
R12422 VGND.n4270 VGND.n4269 4.6505
R12423 VGND.n4272 VGND.n4271 4.6505
R12424 VGND.n4286 VGND.n4285 4.6505
R12425 VGND.n4966 VGND.n4965 4.6505
R12426 VGND.n5520 VGND.n5516 4.6505
R12427 VGND.n5319 VGND.n5318 4.6505
R12428 VGND.n5336 VGND.n5335 4.6505
R12429 VGND.n5340 VGND.n5339 4.6505
R12430 VGND.n5369 VGND.n5368 4.6505
R12431 VGND.n5386 VGND.n5385 4.6505
R12432 VGND.n5390 VGND.n5389 4.6505
R12433 VGND.n5409 VGND.n5408 4.6505
R12434 VGND.n15 VGND.n14 4.6505
R12435 VGND.n19 VGND.n18 4.6505
R12436 VGND.n5586 VGND.n5585 4.6505
R12437 VGND.n5582 VGND.n21 4.6505
R12438 VGND.n5202 VGND.n26 4.6505
R12439 VGND.n5210 VGND.n5209 4.6505
R12440 VGND.n5213 VGND.n5201 4.6505
R12441 VGND.n5248 VGND.n5247 4.6505
R12442 VGND.n5252 VGND.n5251 4.6505
R12443 VGND.n5321 VGND.n5320 4.6505
R12444 VGND.n5324 VGND.n5323 4.6505
R12445 VGND.n5329 VGND.n5328 4.6505
R12446 VGND.n5332 VGND.n5331 4.6505
R12447 VGND.n5333 VGND.n77 4.6505
R12448 VGND.n5342 VGND.n5341 4.6505
R12449 VGND.n5344 VGND.n5343 4.6505
R12450 VGND.n5347 VGND.n5346 4.6505
R12451 VGND.n5349 VGND.n5348 4.6505
R12452 VGND.n5362 VGND.n5361 4.6505
R12453 VGND.n5365 VGND.n5364 4.6505
R12454 VGND.n5367 VGND.n28 4.6505
R12455 VGND.n5371 VGND.n5370 4.6505
R12456 VGND.n5373 VGND.n5372 4.6505
R12457 VGND.n5375 VGND.n5374 4.6505
R12458 VGND.n5377 VGND.n5376 4.6505
R12459 VGND.n5380 VGND.n5379 4.6505
R12460 VGND.n5383 VGND.n74 4.6505
R12461 VGND.n5392 VGND.n5391 4.6505
R12462 VGND.n5394 VGND.n5393 4.6505
R12463 VGND.n5396 VGND.n5395 4.6505
R12464 VGND.n5398 VGND.n5397 4.6505
R12465 VGND.n5401 VGND.n5400 4.6505
R12466 VGND.n5405 VGND.n5404 4.6505
R12467 VGND.n5413 VGND.n5412 4.6505
R12468 VGND.n5415 VGND.n5414 4.6505
R12469 VGND.n5420 VGND.n5419 4.6505
R12470 VGND.n5411 VGND.n5410 4.6505
R12471 VGND.n5407 VGND.n5406 4.6505
R12472 VGND.n5388 VGND.n5387 4.6505
R12473 VGND.n5384 VGND 4.6505
R12474 VGND.n5359 VGND.n5358 4.6505
R12475 VGND.n5357 VGND.n5356 4.6505
R12476 VGND.n5355 VGND.n5354 4.6505
R12477 VGND.n5353 VGND.n5352 4.6505
R12478 VGND.n5351 VGND.n5350 4.6505
R12479 VGND.n5338 VGND.n5337 4.6505
R12480 VGND.n5334 VGND 4.6505
R12481 VGND.n4 VGND.n3 4.6505
R12482 VGND.n6 VGND.n5 4.6505
R12483 VGND.n8 VGND.n7 4.6505
R12484 VGND.n10 VGND.n9 4.6505
R12485 VGND.n13 VGND.n12 4.6505
R12486 VGND.n17 VGND.n16 4.6505
R12487 VGND VGND.n5595 4.6505
R12488 VGND.n5594 VGND.n5593 4.6505
R12489 VGND.n5591 VGND.n5590 4.6505
R12490 VGND.n5588 VGND.n5587 4.6505
R12491 VGND.n5584 VGND.n5583 4.6505
R12492 VGND VGND.n5581 4.6505
R12493 VGND.n5580 VGND.n5579 4.6505
R12494 VGND.n5577 VGND.n5576 4.6505
R12495 VGND.n5574 VGND.n5573 4.6505
R12496 VGND.n5206 VGND.n5205 4.6505
R12497 VGND.n5208 VGND.n5207 4.6505
R12498 VGND.n5212 VGND.n5211 4.6505
R12499 VGND.n5214 VGND 4.6505
R12500 VGND.n5217 VGND.n5216 4.6505
R12501 VGND.n5220 VGND.n5219 4.6505
R12502 VGND.n5222 VGND.n5221 4.6505
R12503 VGND.n5224 VGND.n5223 4.6505
R12504 VGND.n5226 VGND.n5225 4.6505
R12505 VGND.n5230 VGND.n5229 4.6505
R12506 VGND.n5234 VGND.n5233 4.6505
R12507 VGND.n5236 VGND.n5235 4.6505
R12508 VGND.n5241 VGND.n5240 4.6505
R12509 VGND.n5244 VGND.n5243 4.6505
R12510 VGND.n5245 VGND.n5200 4.6505
R12511 VGND.n5246 VGND 4.6505
R12512 VGND.n5250 VGND.n5249 4.6505
R12513 VGND.n5254 VGND.n5253 4.6505
R12514 VGND.n5256 VGND.n5255 4.6505
R12515 VGND.n5259 VGND.n5258 4.6505
R12516 VGND.n5261 VGND.n5260 4.6505
R12517 VGND.n5262 VGND.n27 4.6505
R12518 VGND.n5460 VGND.n5459 4.6505
R12519 VGND.n5462 VGND.n5461 4.6505
R12520 VGND.n5464 VGND.n5463 4.6505
R12521 VGND.n5466 VGND.n5465 4.6505
R12522 VGND.n5467 VGND.n33 4.6505
R12523 VGND.n5468 VGND 4.6505
R12524 VGND.n5471 VGND.n5470 4.6505
R12525 VGND.n5475 VGND.n5474 4.6505
R12526 VGND.n5476 VGND.n32 4.6505
R12527 VGND.n5477 VGND 4.6505
R12528 VGND.n5479 VGND.n5478 4.6505
R12529 VGND.n5481 VGND.n5480 4.6505
R12530 VGND.n5483 VGND.n5482 4.6505
R12531 VGND.n5485 VGND.n5484 4.6505
R12532 VGND.n5487 VGND.n5486 4.6505
R12533 VGND.n5490 VGND.n5489 4.6505
R12534 VGND.n5491 VGND.n31 4.6505
R12535 VGND.n5492 VGND 4.6505
R12536 VGND.n5494 VGND.n5493 4.6505
R12537 VGND.n5496 VGND.n5495 4.6505
R12538 VGND.n5498 VGND.n5497 4.6505
R12539 VGND.n5500 VGND.n5499 4.6505
R12540 VGND.n5502 VGND.n5501 4.6505
R12541 VGND.n5505 VGND.n5504 4.6505
R12542 VGND.n5506 VGND.n30 4.6505
R12543 VGND.n5567 VGND.n5507 4.6505
R12544 VGND.n5566 VGND.n5565 4.6505
R12545 VGND.n5563 VGND.n5562 4.6505
R12546 VGND.n5561 VGND.n5560 4.6505
R12547 VGND.n5559 VGND.n5558 4.6505
R12548 VGND.n5556 VGND.n5555 4.6505
R12549 VGND.n5551 VGND.n5550 4.6505
R12550 VGND.n5548 VGND.n5547 4.6505
R12551 VGND.n5546 VGND 4.6505
R12552 VGND.n5545 VGND.n5509 4.6505
R12553 VGND.n5544 VGND.n5543 4.6505
R12554 VGND.n5542 VGND.n5510 4.6505
R12555 VGND.n5541 VGND.n5540 4.6505
R12556 VGND.n5539 VGND.n5538 4.6505
R12557 VGND.n5537 VGND.n5536 4.6505
R12558 VGND.n5534 VGND.n5533 4.6505
R12559 VGND.n5532 VGND 4.6505
R12560 VGND.n5531 VGND.n5511 4.6505
R12561 VGND.n5530 VGND.n5529 4.6505
R12562 VGND.n5528 VGND.n5512 4.6505
R12563 VGND.n5527 VGND.n5526 4.6505
R12564 VGND.n5525 VGND.n5524 4.6505
R12565 VGND.n5523 VGND.n5522 4.6505
R12566 VGND.n2577 VGND.n2576 4.57589
R12567 VGND.n304 VGND.n303 4.57427
R12568 VGND.n4151 VGND.n4150 4.57427
R12569 VGND.n3724 VGND.n3723 4.57427
R12570 VGND.n3635 VGND.n3634 4.57427
R12571 VGND.n1047 VGND.n1046 4.57427
R12572 VGND.n2241 VGND.n2240 4.57427
R12573 VGND.n2066 VGND.n2065 4.57427
R12574 VGND.n5143 VGND.n5142 4.57427
R12575 VGND.n4466 VGND.n4465 4.57427
R12576 VGND.n5315 VGND.n5314 4.57427
R12577 VGND.n4746 VGND.n4745 4.57412
R12578 VGND.n581 VGND.n495 4.57412
R12579 VGND.n3884 VGND.n3883 4.57412
R12580 VGND.n976 VGND.n885 4.57412
R12581 VGND.n3347 VGND.n3346 4.57412
R12582 VGND.n2949 VGND.n2948 4.57412
R12583 VGND.n2733 VGND.n2732 4.57412
R12584 VGND.n2406 VGND.n2405 4.57412
R12585 VGND.n2016 VGND.n2015 4.57412
R12586 VGND.n5022 VGND.n5021 4.57412
R12587 VGND.n4549 VGND.n4548 4.57412
R12588 VGND.n2260 VGND.n2259 4.57412
R12589 VGND.n4591 VGND.n4590 4.57282
R12590 VGND.n3798 VGND.n3797 4.57282
R12591 VGND.n883 VGND.n882 4.57282
R12592 VGND.n1247 VGND.n1246 4.57282
R12593 VGND.n2644 VGND.n2643 4.57282
R12594 VGND.n2227 VGND.n2226 4.57282
R12595 VGND.n1640 VGND.n1639 4.57282
R12596 VGND.n1613 VGND.n1612 4.5622
R12597 VGND.n4656 VGND.n4655 4.5622
R12598 VGND.n4012 VGND.n4011 4.5622
R12599 VGND.n535 VGND.n534 4.5622
R12600 VGND.n2603 VGND.n2602 4.5622
R12601 VGND.n153 VGND.n152 4.5622
R12602 VGND.n1159 VGND.n1149 4.56192
R12603 VGND.n1374 VGND.n1362 4.56157
R12604 VGND.n3849 VGND.n3848 4.54121
R12605 VGND.n3793 VGND.n3792 4.5005
R12606 VGND.n4418 VGND.n4414 4.44939
R12607 VGND.n2864 VGND.n2863 4.44939
R12608 VGND.n4925 VGND.n4924 4.28986
R12609 VGND.n4410 VGND.n4409 4.28986
R12610 VGND.n1524 VGND.n1523 4.28986
R12611 VGND.n4571 VGND.n357 4.28986
R12612 VGND.n4553 VGND.n363 4.28986
R12613 VGND.n4752 VGND.n4751 4.28986
R12614 VGND.n4826 VGND.n4825 4.28986
R12615 VGND.n4054 VGND.n4053 4.28986
R12616 VGND.n4030 VGND.n4029 4.28986
R12617 VGND.n4025 VGND.n502 4.28986
R12618 VGND.n416 VGND.n415 4.28986
R12619 VGND.n466 VGND.n440 4.28986
R12620 VGND.n462 VGND.n461 4.28986
R12621 VGND.n4099 VGND.n395 4.28986
R12622 VGND.n4006 VGND.n4005 4.28986
R12623 VGND.n3888 VGND.n3887 4.28986
R12624 VGND.n634 VGND.n633 4.28986
R12625 VGND.n697 VGND.n663 4.28986
R12626 VGND.n3731 VGND.n3730 4.28986
R12627 VGND.n3733 VGND.n3732 4.28986
R12628 VGND.n3801 VGND.n644 4.28986
R12629 VGND.n3512 VGND.n3511 4.28986
R12630 VGND.n3244 VGND.n3243 4.28986
R12631 VGND.n3239 VGND.n1043 4.28986
R12632 VGND.n1089 VGND.n1088 4.28986
R12633 VGND.n3187 VGND.n1097 4.28986
R12634 VGND.n2892 VGND.n2891 4.28986
R12635 VGND.n1369 VGND.n1364 4.28986
R12636 VGND.n2625 VGND.n2624 4.28986
R12637 VGND.n2824 VGND.n2823 4.28986
R12638 VGND.n2445 VGND.n2444 4.28986
R12639 VGND.n2142 VGND.n2128 4.28986
R12640 VGND.n2175 VGND.n2174 4.28986
R12641 VGND.n2183 VGND.n2182 4.28986
R12642 VGND.n2309 VGND.n1488 4.28986
R12643 VGND.n1224 VGND.n1192 4.26609
R12644 VGND.n1884 VGND.n1883 4.14168
R12645 VGND.n24 VGND.n23 4.07323
R12646 VGND.n76 VGND.n75 4.07323
R12647 VGND.n257 VGND.n256 4.07323
R12648 VGND.n4318 VGND.n4317 4.07323
R12649 VGND.n4235 VGND.n4222 4.07323
R12650 VGND.n4236 VGND.n4235 4.07323
R12651 VGND.n4210 VGND.n4209 4.07323
R12652 VGND.n1658 VGND.n1657 4.07323
R12653 VGND.n1652 VGND.n1651 4.07323
R12654 VGND.n1718 VGND.n1652 4.07323
R12655 VGND.n1529 VGND.n1528 4.07323
R12656 VGND.n1647 VGND.n1646 4.07323
R12657 VGND.n1727 VGND.n1647 4.07323
R12658 VGND.n1710 VGND.n1709 4.07323
R12659 VGND.n1709 VGND.n1654 4.07323
R12660 VGND.n499 VGND.n498 4.07323
R12661 VGND.n498 VGND.n497 4.07323
R12662 VGND.n4029 VGND.n501 4.07323
R12663 VGND.n443 VGND.n442 4.07323
R12664 VGND.n505 VGND.n504 4.07323
R12665 VGND.n522 VGND.n521 4.07323
R12666 VGND.n545 VGND.n522 4.07323
R12667 VGND.n525 VGND.n524 4.07323
R12668 VGND.n656 VGND.n655 4.07323
R12669 VGND.n657 VGND.n656 4.07323
R12670 VGND.n700 VGND.n663 4.07323
R12671 VGND.n673 VGND.n672 4.07323
R12672 VGND.n675 VGND.n673 4.07323
R12673 VGND.n736 VGND.n648 4.07323
R12674 VGND.n736 VGND.n735 4.07323
R12675 VGND.n3976 VGND.n630 4.07323
R12676 VGND.n640 VGND.n639 4.07323
R12677 VGND.n810 VGND.n809 4.07323
R12678 VGND.n776 VGND.n775 4.07323
R12679 VGND.n3474 VGND.n889 4.07323
R12680 VGND.n968 VGND.n967 4.07323
R12681 VGND.n3358 VGND.n3357 4.07323
R12682 VGND.n3226 VGND.n1045 4.07323
R12683 VGND.n1062 VGND.n1061 4.07323
R12684 VGND.n1061 VGND.n1055 4.07323
R12685 VGND.n1032 VGND.n1031 4.07323
R12686 VGND.n2891 VGND.n1269 4.07323
R12687 VGND.n1158 VGND.n1150 4.07323
R12688 VGND.n1195 VGND.n1194 4.07323
R12689 VGND.n3060 VGND.n1130 4.07323
R12690 VGND.n3060 VGND.n3059 4.07323
R12691 VGND.n2743 VGND.n2742 4.07323
R12692 VGND.n2782 VGND.n2737 4.07323
R12693 VGND.n2786 VGND.n2785 4.07323
R12694 VGND.n2591 VGND.n2590 4.07323
R12695 VGND.n1339 VGND.n1338 4.07323
R12696 VGND.n2647 VGND.n1339 4.07323
R12697 VGND.n2298 VGND.n1490 4.07323
R12698 VGND.n2135 VGND.n2132 4.07323
R12699 VGND.n2131 VGND.n2130 4.07323
R12700 VGND.n1463 VGND.n1462 4.07323
R12701 VGND.n1483 VGND.n1482 4.07323
R12702 VGND.n1780 VGND.n1755 4.07323
R12703 VGND.n1755 VGND.n1754 4.07323
R12704 VGND.n156 VGND.n155 4.07323
R12705 VGND.n1881 VGND.n1880 4.07323
R12706 VGND.n5091 VGND.n5090 4.07323
R12707 VGND.n5090 VGND.n106 4.07323
R12708 VGND.n109 VGND.n108 4.07323
R12709 VGND.n5514 VGND.n5513 4.07323
R12710 VGND.n4232 VGND 3.95686
R12711 VGND.n4903 VGND.n4901 3.85748
R12712 VGND.n3023 VGND.n3022 3.85748
R12713 VGND.n4909 VGND.n257 3.76521
R12714 VGND.n3849 VGND.n641 3.71925
R12715 VGND.n1613 VGND.n1590 3.69828
R12716 VGND.n1632 VGND.n1631 3.65764
R12717 VGND.n4825 VGND.n4824 3.61789
R12718 VGND.n4664 VGND.n4663 3.61789
R12719 VGND.n461 VGND.n460 3.61789
R12720 VGND.n1377 VGND.n1362 3.56403
R12721 VGND.n3813 VGND.n3812 3.50735
R12722 VGND.n919 VGND.n918 3.50735
R12723 VGND.n1874 VGND.n1873 3.50735
R12724 VGND.n3833 VGND.n3832 3.50735
R12725 VGND.n2041 VGND.n1522 3.47666
R12726 VGND.n4218 VGND.n4217 3.44377
R12727 VGND.n1585 VGND.n1584 3.44377
R12728 VGND.n1584 VGND.n1583 3.44377
R12729 VGND.n1538 VGND.n1537 3.44377
R12730 VGND.n337 VGND.n314 3.44377
R12731 VGND.n835 VGND.n834 3.44377
R12732 VGND.n908 VGND.n907 3.44377
R12733 VGND.n913 VGND.n908 3.44377
R12734 VGND.n2854 VGND.n2853 3.44377
R12735 VGND.n2853 VGND.n2852 3.44377
R12736 VGND.n1470 VGND.n1469 3.44377
R12737 VGND.n1469 VGND.n1468 3.44377
R12738 VGND.n204 VGND.n203 3.44377
R12739 VGND.n132 VGND.n131 3.44377
R12740 VGND.n1957 VGND.n1956 3.44377
R12741 VGND.n1956 VGND.n1955 3.44377
R12742 VGND.n4729 VGND.n4728 3.4105
R12743 VGND.n4545 VGND.n4544 3.4105
R12744 VGND.n4600 VGND 3.4105
R12745 VGND.n4609 VGND.n4608 3.4105
R12746 VGND.n592 VGND.n591 3.4105
R12747 VGND.n4171 VGND.n4170 3.4105
R12748 VGND.n4156 VGND 3.4105
R12749 VGND.n4149 VGND.n4148 3.4105
R12750 VGND.n3867 VGND.n3866 3.4105
R12751 VGND.n3705 VGND.n3704 3.4105
R12752 VGND.n3791 VGND 3.4105
R12753 VGND.n3783 VGND.n3782 3.4105
R12754 VGND.n987 VGND.n986 3.4105
R12755 VGND.n3658 VGND.n3657 3.4105
R12756 VGND.n3640 VGND 3.4105
R12757 VGND.n3633 VGND.n3632 3.4105
R12758 VGND.n3330 VGND.n3329 3.4105
R12759 VGND.n3151 VGND.n3150 3.4105
R12760 VGND.n3210 VGND 3.4105
R12761 VGND.n3219 VGND.n3218 3.4105
R12762 VGND.n2953 VGND.n2952 3.4105
R12763 VGND.n3091 VGND.n3090 3.4105
R12764 VGND.n3076 VGND 3.4105
R12765 VGND.n3070 VGND.n3069 3.4105
R12766 VGND.n2716 VGND.n2715 3.4105
R12767 VGND.n2553 VGND.n2552 3.4105
R12768 VGND VGND.n2638 3.4105
R12769 VGND.n2630 VGND.n2629 3.4105
R12770 VGND.n2381 VGND.n2380 3.4105
R12771 VGND.n2264 VGND.n2263 3.4105
R12772 VGND.n2246 VGND 3.4105
R12773 VGND.n2239 VGND.n2238 3.4105
R12774 VGND.n1818 VGND.n1817 3.4105
R12775 VGND.n2089 VGND.n2088 3.4105
R12776 VGND.n2071 VGND 3.4105
R12777 VGND.n2064 VGND.n2063 3.4105
R12778 VGND.n5026 VGND.n5025 3.4105
R12779 VGND.n5166 VGND.n5165 3.4105
R12780 VGND.n5148 VGND 3.4105
R12781 VGND.n5141 VGND.n5140 3.4105
R12782 VGND.n5273 VGND.n5272 3.4105
R12783 VGND.n4420 VGND.n4418 3.36892
R12784 VGND.n3157 VGND.n3156 3.36892
R12785 VGND.n1649 VGND 3.29747
R12786 VGND.n3182 VGND 3.29747
R12787 VGND.n1232 VGND 3.29747
R12788 VGND.n2343 VGND 3.29747
R12789 VGND.n4285 VGND.n4212 3.28385
R12790 VGND VGND.n1271 3.26859
R12791 VGND.n3731 VGND.n3729 3.26272
R12792 VGND.n2415 VGND.n2414 3.26272
R12793 VGND.n4917 VGND 3.24826
R12794 VGND.n1598 VGND 3.24826
R12795 VGND.n66 VGND.n65 3.2005
R12796 VGND.n72 VGND.n71 3.2005
R12797 VGND.n3817 VGND.n3816 3.2005
R12798 VGND.n3837 VGND.n3836 3.2005
R12799 VGND.n832 VGND.n831 3.2005
R12800 VGND.n781 VGND.n780 3.2005
R12801 VGND.n917 VGND.n914 3.2005
R12802 VGND.n1038 VGND.n1037 3.2005
R12803 VGND.n2802 VGND.n2799 3.2005
R12804 VGND.n2585 VGND.n2584 3.2005
R12805 VGND.n1474 VGND.n1473 3.2005
R12806 VGND.n1872 VGND.n1869 3.2005
R12807 VGND.n2880 VGND.n1273 3.13259
R12808 VGND.n13 VGND.n1 3.13242
R12809 VGND.n5419 VGND.n5418 3.13242
R12810 VGND.n4372 VGND.n4328 3.13242
R12811 VGND.n4388 VGND.n4325 3.13242
R12812 VGND.n4399 VGND.n4321 3.13242
R12813 VGND.n4447 VGND.n4310 3.13242
R12814 VGND.n1551 VGND.n1550 3.13242
R12815 VGND.n1757 VGND.n1756 3.13242
R12816 VGND.n1763 VGND.n1757 3.13242
R12817 VGND.n4762 VGND.n4761 3.13242
R12818 VGND.n310 VGND.n309 3.13242
R12819 VGND.n4580 VGND.n355 3.13242
R12820 VGND.n4556 VGND.n361 3.13242
R12821 VGND.n4667 VGND.n300 3.13242
R12822 VGND.n4060 VGND.n4059 3.13242
R12823 VGND.n4073 VGND.n4072 3.13242
R12824 VGND.n4072 VGND.n4071 3.13242
R12825 VGND.n4084 VGND.n4083 3.13242
R12826 VGND.n400 VGND.n399 3.13242
R12827 VGND.n476 VGND.n438 3.13242
R12828 VGND.n3907 VGND.n3906 3.13242
R12829 VGND.n710 VGND.n709 3.13242
R12830 VGND.n817 VGND.n772 3.13242
R12831 VGND.n827 VGND.n826 3.13242
R12832 VGND.n875 VGND.n827 3.13242
R12833 VGND.n764 VGND.n763 3.13242
R12834 VGND.n765 VGND.n764 3.13242
R12835 VGND.n938 VGND.n905 3.13242
R12836 VGND.n945 VGND.n903 3.13242
R12837 VGND.n3263 VGND.n3262 3.13242
R12838 VGND.n3191 VGND.n1094 3.13242
R12839 VGND.n3175 VGND.n1103 3.13242
R12840 VGND.n3306 VGND.n1033 3.13242
R12841 VGND.n2918 VGND.n2917 3.13242
R12842 VGND.n2917 VGND.n2916 3.13242
R12843 VGND.n2930 VGND.n2899 3.13242
R12844 VGND.n1167 VGND.n1146 3.13242
R12845 VGND.n1182 VGND.n1181 3.13242
R12846 VGND.n1181 VGND.n1140 3.13242
R12847 VGND.n1234 VGND.n1233 3.13242
R12848 VGND.n2997 VGND.n1251 3.13242
R12849 VGND.n2992 VGND.n1254 3.13242
R12850 VGND.n2986 VGND.n2985 3.13242
R12851 VGND.n2978 VGND.n1257 3.13242
R12852 VGND.n2593 VGND.n1340 3.13242
R12853 VGND.n1385 VGND.n1359 3.13242
R12854 VGND.n1400 VGND.n1399 3.13242
R12855 VGND.n1399 VGND.n1351 3.13242
R12856 VGND.n1346 VGND.n1345 3.13242
R12857 VGND.n1337 VGND.n1336 3.13242
R12858 VGND.n2438 VGND.n2437 3.13242
R12859 VGND.n2213 VGND.n2170 3.13242
R12860 VGND.n2207 VGND.n2206 3.13242
R12861 VGND.n1481 VGND.n1480 3.13242
R12862 VGND.n1887 VGND.n1886 3.13242
R12863 VGND.n5110 VGND.n5109 3.13242
R12864 VGND.n5070 VGND.n113 3.13242
R12865 VGND.n5258 VGND.n5257 3.13241
R12866 VGND.n5205 VGND.n5204 3.13241
R12867 VGND.n5590 VGND.n5589 3.13241
R12868 VGND.n1 VGND.n0 3.13241
R12869 VGND.n5418 VGND.n5417 3.13241
R12870 VGND.n5346 VGND.n5345 3.13241
R12871 VGND.n5459 VGND.n5458 3.13241
R12872 VGND.n5474 VGND.n5473 3.13241
R12873 VGND.n5489 VGND.n5488 3.13241
R12874 VGND.n5504 VGND.n5503 3.13241
R12875 VGND.n4922 VGND.n4921 3.13241
R12876 VGND.n4328 VGND.n4327 3.13241
R12877 VGND.n4325 VGND.n4324 3.13241
R12878 VGND.n4321 VGND.n4320 3.13241
R12879 VGND.n4310 VGND.n4309 3.13241
R12880 VGND.n4465 VGND.n4464 3.13241
R12881 VGND.n2024 VGND.n2023 3.13241
R12882 VGND.n1738 VGND.n1737 3.13241
R12883 VGND.n4763 VGND.n4762 3.13241
R12884 VGND.n309 VGND.n308 3.13241
R12885 VGND.n355 VGND.n354 3.13241
R12886 VGND.n361 VGND.n360 3.13241
R12887 VGND.n4614 VGND.n4613 3.13241
R12888 VGND.n4786 VGND.n4785 3.13241
R12889 VGND.n4799 VGND.n4798 3.13241
R12890 VGND.n4839 VGND.n4838 3.13241
R12891 VGND.n4853 VGND.n4852 3.13241
R12892 VGND.n4668 VGND.n4667 3.13241
R12893 VGND.n4709 VGND.n4708 3.13241
R12894 VGND.n4061 VGND.n4060 3.13241
R12895 VGND.n4085 VGND.n4084 3.13241
R12896 VGND.n399 VGND.n398 3.13241
R12897 VGND.n438 VGND.n437 3.13241
R12898 VGND.n4111 VGND.n4110 3.13241
R12899 VGND.n391 VGND.n390 3.13241
R12900 VGND.n564 VGND.n563 3.13241
R12901 VGND.n3908 VGND.n3907 3.13241
R12902 VGND.n3951 VGND.n3950 3.13241
R12903 VGND.n709 VGND.n708 3.13241
R12904 VGND.n3777 VGND.n3776 3.13241
R12905 VGND.n3753 VGND.n3752 3.13241
R12906 VGND.n772 VGND.n771 3.13241
R12907 VGND.n784 VGND.n783 3.13241
R12908 VGND.n3622 VGND.n3621 3.13241
R12909 VGND.n3538 VGND.n3537 3.13241
R12910 VGND.n3553 VGND.n3552 3.13241
R12911 VGND.n3516 VGND.n3515 3.13241
R12912 VGND.n3496 VGND.n3495 3.13241
R12913 VGND.n905 VGND.n904 3.13241
R12914 VGND.n903 VGND.n902 3.13241
R12915 VGND.n961 VGND.n960 3.13241
R12916 VGND.n3372 VGND.n3371 3.13241
R12917 VGND.n3386 VGND.n3385 3.13241
R12918 VGND.n3400 VGND.n3399 3.13241
R12919 VGND.n3254 VGND.n3253 3.13241
R12920 VGND.n1094 VGND.n1093 3.13241
R12921 VGND.n1103 VGND.n1102 3.13241
R12922 VGND.n3418 VGND.n3417 3.13241
R12923 VGND.n3429 VGND.n3428 3.13241
R12924 VGND.n3445 VGND.n3444 3.13241
R12925 VGND.n3307 VGND.n3306 3.13241
R12926 VGND.n2933 VGND.n2899 3.13241
R12927 VGND.n2881 VGND.n2880 3.13241
R12928 VGND.n3018 VGND.n3017 3.13241
R12929 VGND.n3043 VGND.n3042 3.13241
R12930 VGND.n1164 VGND.n1146 3.13241
R12931 VGND.n1235 VGND.n1234 3.13241
R12932 VGND.n3009 VGND.n3008 3.13241
R12933 VGND.n1251 VGND.n1250 3.13241
R12934 VGND.n1254 VGND.n1253 3.13241
R12935 VGND.n2987 VGND.n2986 3.13241
R12936 VGND.n1257 VGND.n1256 3.13241
R12937 VGND.n2967 VGND.n2966 3.13241
R12938 VGND.n2791 VGND.n2790 3.13241
R12939 VGND.n2594 VGND.n2593 3.13241
R12940 VGND.n1382 VGND.n1359 3.13241
R12941 VGND VGND.n1412 3.13241
R12942 VGND.n1345 VGND.n1344 3.13241
R12943 VGND.n1447 VGND.n1446 3.13241
R12944 VGND.n1336 VGND.n1335 3.13241
R12945 VGND.n2696 VGND.n2695 3.13241
R12946 VGND.n2422 VGND.n2421 3.13241
R12947 VGND.n2419 VGND.n2418 3.13241
R12948 VGND.n2439 VGND.n2438 3.13241
R12949 VGND.n2464 VGND.n2463 3.13241
R12950 VGND.n2473 VGND.n2472 3.13241
R12951 VGND.n2304 VGND.n2303 3.13241
R12952 VGND.n2170 VGND.n2169 3.13241
R12953 VGND.n2208 VGND.n2207 3.13241
R12954 VGND.n2277 VGND.n2276 3.13241
R12955 VGND.n2323 VGND.n2322 3.13241
R12956 VGND.n1480 VGND.n1479 3.13241
R12957 VGND.n2361 VGND.n2360 3.13241
R12958 VGND.n1804 VGND.n1803 3.13241
R12959 VGND.n1892 VGND.n1886 3.13241
R12960 VGND.n180 VGND.n179 3.13241
R12961 VGND.n5130 VGND.n5129 3.13241
R12962 VGND.n1922 VGND.n1921 3.13241
R12963 VGND.n1966 VGND.n1965 3.13241
R12964 VGND.n1974 VGND.n1973 3.13241
R12965 VGND.n113 VGND.n112 3.13241
R12966 VGND.n5536 VGND.n5535 3.13241
R12967 VGND.n5421 VGND.n29 3.06214
R12968 VGND.n4537 VGND.n4536 3.0005
R12969 VGND.n4163 VGND.n4162 3.0005
R12970 VGND.n3714 VGND.n3713 3.0005
R12971 VGND.n3647 VGND.n3646 3.0005
R12972 VGND.n3143 VGND.n3142 3.0005
R12973 VGND.n1287 VGND.n1286 3.0005
R12974 VGND.n3083 VGND.n3082 3.0005
R12975 VGND.n2567 VGND.n2566 3.0005
R12976 VGND.n2401 VGND.n2400 3.0005
R12977 VGND.n2253 VGND.n2252 3.0005
R12978 VGND.n2078 VGND.n2077 3.0005
R12979 VGND.n5155 VGND.n5154 3.0005
R12980 VGND.n4484 VGND.n4483 3.0005
R12981 VGND.n5297 VGND.n5296 3.0005
R12982 VGND.n1662 VGND.n1661 2.9514
R12983 VGND.n4568 VGND.n357 2.9514
R12984 VGND.n4053 VGND.n4052 2.9514
R12985 VGND.n409 VGND.n408 2.9514
R12986 VGND.n415 VGND.n402 2.9514
R12987 VGND.n653 VGND.n651 2.9514
R12988 VGND.n1088 VGND.n1051 2.9514
R12989 VGND.n3407 VGND.n3406 2.9514
R12990 VGND.n2895 VGND.n1270 2.9514
R12991 VGND.n1330 VGND.n1328 2.9514
R12992 VGND.n1412 VGND.n1347 2.9514
R12993 VGND.n2175 VGND.n2173 2.9514
R12994 VGND.n5405 VGND.n67 2.89365
R12995 VGND.n74 VGND.n73 2.89365
R12996 VGND.n3820 VGND.n643 2.89365
R12997 VGND.n3840 VGND.n642 2.89365
R12998 VGND.n862 VGND.n833 2.89365
R12999 VGND.n790 VGND.n782 2.89365
R13000 VGND.n925 VGND.n906 2.89365
R13001 VGND.n1040 VGND.n1039 2.89365
R13002 VGND.n2798 VGND.n2797 2.89365
R13003 VGND.n2611 VGND.n2586 2.89365
R13004 VGND.n1476 VGND.n1475 2.89365
R13005 VGND.n1578 VGND.n1542 2.76214
R13006 VGND.n1572 VGND.n1571 2.76214
R13007 VGND.n2803 VGND.n1330 2.76214
R13008 VGND.n2483 VGND.n2482 2.76214
R13009 VGND.n4283 VGND.n4282 2.64086
R13010 VGND.n4459 VGND.n4458 2.63579
R13011 VGND.n1231 VGND 2.53073
R13012 VGND.n4719 VGND.n4718 2.47351
R13013 VGND.n4858 VGND.n4857 2.47351
R13014 VGND.n599 VGND.n598 2.47351
R13015 VGND.n4004 VGND.n4003 2.47351
R13016 VGND.n3857 VGND.n3856 2.47351
R13017 VGND.n3983 VGND.n3982 2.47351
R13018 VGND.n994 VGND.n993 2.47351
R13019 VGND.n3471 VGND.n3470 2.47351
R13020 VGND.n3320 VGND.n3319 2.47351
R13021 VGND.n3450 VGND.n3449 2.47351
R13022 VGND.n2962 VGND.n2959 2.47351
R13023 VGND.n2848 VGND.n2847 2.47351
R13024 VGND.n2706 VGND.n2705 2.47351
R13025 VGND.n2827 VGND.n2826 2.47351
R13026 VGND.n2371 VGND.n2370 2.47351
R13027 VGND.n2509 VGND.n2508 2.47351
R13028 VGND.n1825 VGND.n1824 2.47351
R13029 VGND.n2000 VGND.n1999 2.47351
R13030 VGND.n5033 VGND.n5032 2.47351
R13031 VGND.n1979 VGND.n1978 2.47351
R13032 VGND.n4368 VGND.n4344 2.47351
R13033 VGND.n4881 VGND.n4880 2.47351
R13034 VGND.n5457 VGND.n5456 2.47351
R13035 VGND.n5446 VGND.n5445 2.47351
R13036 VGND.n2042 VGND.n2041 2.45595
R13037 VGND.n1362 VGND.n1361 2.44917
R13038 VGND.n1149 VGND.n1148 2.44882
R13039 VGND.n2602 VGND.n2601 2.44756
R13040 VGND.n172 VGND.n171 2.43325
R13041 VGND.n205 VGND.n204 2.43325
R13042 VGND.n133 VGND.n132 2.43325
R13043 VGND.n4212 VGND.n4211 2.4297
R13044 VGND.n4281 VGND.n4278 2.35386
R13045 VGND.n4778 VGND.n4754 2.29662
R13046 VGND.n4551 VGND.n365 2.29662
R13047 VGND.n4097 VGND.n396 2.29662
R13048 VGND.n561 VGND.n519 2.29662
R13049 VGND.n4028 VGND.n4027 2.29662
R13050 VGND.n4009 VGND.n4008 2.29662
R13051 VGND.n464 VGND.n441 2.29662
R13052 VGND.n3804 VGND.n3803 2.29662
R13053 VGND.n3852 VGND.n3851 2.29662
R13054 VGND.n3935 VGND.n635 2.29662
R13055 VGND.n3976 VGND.n3975 2.29662
R13056 VGND.n737 VGND.n736 2.29662
R13057 VGND.n3514 VGND.n3513 2.29662
R13058 VGND.n3242 VGND.n3241 2.29662
R13059 VGND.n1073 VGND.n1072 2.29662
R13060 VGND.n3185 VGND.n1099 2.29662
R13061 VGND.n2890 VGND.n2889 2.29662
R13062 VGND.n2622 VGND.n2621 2.29662
R13063 VGND.n2782 VGND.n2781 2.29662
R13064 VGND.n2822 VGND.n1321 2.29662
R13065 VGND.n1372 VGND.n1371 2.29662
R13066 VGND.n1377 VGND.n1376 2.29662
R13067 VGND.n2298 VGND.n1491 2.29662
R13068 VGND.n2145 VGND.n2144 2.29662
R13069 VGND.n2314 VGND.n2313 2.29662
R13070 VGND.n2046 VGND.n1522 2.29662
R13071 VGND.n1605 VGND.n1604 2.29662
R13072 VGND.n1608 VGND.n1607 2.29662
R13073 VGND.n1617 VGND.n1616 2.29662
R13074 VGND.n1567 VGND.n1546 2.29662
R13075 VGND.n1566 VGND.n1548 2.29662
R13076 VGND.n169 VGND.n128 2.29662
R13077 VGND.n201 VGND.n200 2.29662
R13078 VGND.n193 VGND.n172 2.29662
R13079 VGND.n4408 VGND.n4407 2.29662
R13080 VGND.n4884 VGND.n4883 2.29662
R13081 VGND.n4886 VGND.n4885 2.29662
R13082 VGND.n4261 VGND.n4260 2.29662
R13083 VGND.n411 VGND.n410 2.29643
R13084 VGND.n3184 VGND.n3183 2.29643
R13085 VGND.n3061 VGND.n3060 2.29643
R13086 VGND.n969 VGND.n968 2.28155
R13087 VGND.n1283 VGND.n1282 2.28144
R13088 VGND.n5039 VGND.n5038 2.27995
R13089 VGND.n565 VGND.n564 2.17922
R13090 VGND.n5233 VGND.n5232 2.01694
R13091 VGND.n1578 VGND.n1577 2.01694
R13092 VGND.n1577 VGND.n1575 2.01694
R13093 VGND.n174 VGND.n173 2.00532
R13094 VGND.n3733 VGND.n3731 1.97497
R13095 VGND.n2445 VGND.n2415 1.97497
R13096 VGND.n4285 VGND.n4284 1.89467
R13097 VGND.n4416 VGND.n4415 1.79699
R13098 VGND.n4219 VGND.n4218 1.79699
R13099 VGND.n1536 VGND.n1535 1.79699
R13100 VGND.n313 VGND.n312 1.79699
R13101 VGND.n2164 VGND.n2163 1.79699
R13102 VGND.n2166 VGND.n2165 1.79699
R13103 VGND.n836 VGND.n835 1.72214
R13104 VGND.n855 VGND.n836 1.72214
R13105 VGND.n1202 VGND.n1201 1.72214
R13106 VGND.n1955 VGND.n1954 1.72214
R13107 VGND.n3234 VGND.n3233 1.7005
R13108 VGND.n4769 VGND.n4768 1.6905
R13109 VGND.n4139 VGND.n4138 1.6905
R13110 VGND.n3598 VGND.n761 1.6905
R13111 VGND.n3491 VGND.n888 1.6905
R13112 VGND.n3580 VGND.n3579 1.6905
R13113 VGND.n3302 VGND.n3301 1.6905
R13114 VGND.n2283 VGND.n2282 1.6905
R13115 VGND.n2189 VGND.n2188 1.6905
R13116 VGND.n143 VGND.n136 1.6905
R13117 VGND.n4417 VGND.n4416 1.64728
R13118 VGND.n4254 VGND.n4219 1.64728
R13119 VGND.n1537 VGND.n1536 1.64728
R13120 VGND.n314 VGND.n313 1.64728
R13121 VGND.n3157 VGND.n3153 1.64728
R13122 VGND.n2865 VGND.n2862 1.64728
R13123 VGND.n2165 VGND.n2164 1.64728
R13124 VGND.n2167 VGND.n2166 1.64728
R13125 VGND.n3523 VGND.n3522 1.6005
R13126 VGND.n317 VGND.n316 1.50646
R13127 VGND.n406 VGND.n405 1.50646
R13128 VGND.n676 VGND.n674 1.50646
R13129 VGND.n840 VGND.n839 1.50646
R13130 VGND.n1057 VGND.n1056 1.50646
R13131 VGND.n1152 VGND.n1151 1.50646
R13132 VGND.n1367 VGND.n1366 1.50646
R13133 VGND.n2134 VGND.n2133 1.50646
R13134 VGND.n1595 VGND.n1594 1.50646
R13135 VGND.n138 VGND.n137 1.50646
R13136 VGND.n4224 VGND.n4223 1.50646
R13137 VGND.n3190 VGND.n3189 1.50638
R13138 VGND.n1582 VGND.n1581 1.50008
R13139 VGND.n4659 VGND.n301 1.49961
R13140 VGND.n548 VGND.n522 1.49961
R13141 VGND.n4017 VGND.n505 1.49961
R13142 VGND.n4032 VGND.n501 1.49961
R13143 VGND.n4038 VGND.n498 1.49961
R13144 VGND.n536 VGND.n525 1.49961
R13145 VGND.n3927 VGND.n3890 1.49961
R13146 VGND.n679 VGND.n673 1.49961
R13147 VGND.n700 VGND.n699 1.49961
R13148 VGND.n719 VGND.n656 1.49961
R13149 VGND.n3474 VGND.n3473 1.49961
R13150 VGND.n809 VGND.n808 1.49961
R13151 VGND.n3226 VGND.n3225 1.49961
R13152 VGND.n3361 VGND.n3358 1.49961
R13153 VGND.n1061 VGND.n1060 1.49961
R13154 VGND.n2894 VGND.n1269 1.49961
R13155 VGND.n1158 VGND.n1157 1.49961
R13156 VGND.n1221 VGND.n1194 1.49961
R13157 VGND.n2605 VGND.n2591 1.49961
R13158 VGND.n2785 VGND.n2784 1.49961
R13159 VGND.n2746 VGND.n2743 1.49961
R13160 VGND.n2650 VGND.n1339 1.49961
R13161 VGND.n2296 VGND.n1493 1.49961
R13162 VGND.n2341 VGND.n1483 1.49961
R13163 VGND.n2501 VGND.n1463 1.49961
R13164 VGND.n2138 VGND.n2132 1.49961
R13165 VGND.n2032 VGND.n1529 1.49961
R13166 VGND.n1783 VGND.n1755 1.49961
R13167 VGND.n1730 VGND.n1647 1.49961
R13168 VGND.n1721 VGND.n1652 1.49961
R13169 VGND.n1709 VGND.n1708 1.49961
R13170 VGND.n1698 VGND.n1658 1.49961
R13171 VGND.n5090 VGND.n5089 1.49961
R13172 VGND.n1900 VGND.n1881 1.49961
R13173 VGND.n155 VGND.n154 1.49961
R13174 VGND.n4405 VGND.n4318 1.49961
R13175 VGND.n4908 VGND.n257 1.49961
R13176 VGND.n4930 VGND.n4927 1.49961
R13177 VGND.n4235 VGND.n4234 1.49961
R13178 VGND.n4288 VGND.n4210 1.49961
R13179 VGND.n5366 VGND.n76 1.49961
R13180 VGND.n5575 VGND.n24 1.49961
R13181 VGND.n2037 VGND.n1525 1.49956
R13182 VGND.n3246 VGND.n1042 1.49933
R13183 VGND.n4760 VGND.n4759 1.49932
R13184 VGND.n452 VGND.n443 1.49932
R13185 VGND.n448 VGND.n447 1.49932
R13186 VGND.n4050 VGND.n4049 1.49932
R13187 VGND.n3898 VGND.n3897 1.49932
R13188 VGND.n807 VGND.n776 1.49932
R13189 VGND.n3525 VGND.n3524 1.49932
R13190 VGND.n3360 VGND.n3359 1.49932
R13191 VGND.n2909 VGND.n2908 1.49932
R13192 VGND.n2745 VGND.n2744 1.49932
R13193 VGND.n2139 VGND.n2130 1.49932
R13194 VGND.n2425 VGND.n2424 1.49932
R13195 VGND.n1664 VGND.n1663 1.49932
R13196 VGND.n5081 VGND.n109 1.49932
R13197 VGND.n1889 VGND.n1888 1.49932
R13198 VGND.n4929 VGND.n4928 1.49932
R13199 VGND.n5521 VGND.n5514 1.49932
R13200 VGND.n4278 VGND.n4277 1.32068
R13201 VGND.n3855 VGND.n640 1.27165
R13202 VGND.n3318 VGND.n1032 1.27165
R13203 VGND.n1413 VGND 1.15795
R13204 VGND VGND.n2578 1.15795
R13205 VGND.n5455 VGND.n5454 1.14176
R13206 VGND.n4527 VGND.n4524 1.14113
R13207 VGND.n4174 VGND.n4173 1.14113
R13208 VGND.n3697 VGND.n3694 1.14113
R13209 VGND.n3661 VGND.n3660 1.14113
R13210 VGND.n3126 VGND.n3123 1.14113
R13211 VGND.n3094 VGND.n3093 1.14113
R13212 VGND.n2545 VGND.n2542 1.14113
R13213 VGND.n2267 VGND.n2266 1.14113
R13214 VGND.n2092 VGND.n2091 1.14113
R13215 VGND.n5169 VGND.n5168 1.14113
R13216 VGND.n5198 VGND.n5183 1.14113
R13217 VGND.n5454 VGND.n5447 1.14113
R13218 VGND.n4860 VGND.n273 1.14113
R13219 VGND.n3999 VGND.n600 1.14113
R13220 VGND.n3985 VGND.n610 1.14113
R13221 VGND.n3466 VGND.n995 1.14113
R13222 VGND.n3452 VGND.n1004 1.14113
R13223 VGND.n2843 VGND.n1262 1.14113
R13224 VGND.n2829 VGND.n1303 1.14113
R13225 VGND.n2511 VGND.n1453 1.14113
R13226 VGND.n1995 VGND.n1826 1.14113
R13227 VGND.n1981 VGND.n119 1.14113
R13228 VGND.n5243 VGND.n5242 1.14023
R13229 VGND.n67 VGND.n66 1.14023
R13230 VGND.n73 VGND.n72 1.14023
R13231 VGND.n5331 VGND.n5330 1.14023
R13232 VGND.n4943 VGND.n4942 1.14023
R13233 VGND.n1675 VGND.n1674 1.14023
R13234 VGND.n4808 VGND.n4807 1.14023
R13235 VGND.n3959 VGND.n3958 1.14023
R13236 VGND.n3817 VGND.n643 1.14023
R13237 VGND.n3837 VGND.n642 1.14023
R13238 VGND.n833 VGND.n832 1.14023
R13239 VGND.n782 VGND.n781 1.14023
R13240 VGND.n914 VGND.n906 1.14023
R13241 VGND.n1039 VGND.n1038 1.14023
R13242 VGND.n2757 VGND.n2756 1.14023
R13243 VGND.n2799 VGND.n2798 1.14023
R13244 VGND.n2586 VGND.n2585 1.14023
R13245 VGND.n1475 VGND.n1474 1.14023
R13246 VGND.n1869 VGND.n1868 1.14023
R13247 VGND.n5040 VGND.n5039 1.14023
R13248 VGND.n5550 VGND.n5549 1.14023
R13249 VGND.n4860 VGND.n4859 1.1392
R13250 VGND.n4002 VGND.n3999 1.1392
R13251 VGND.n3985 VGND.n3984 1.1392
R13252 VGND.n3469 VGND.n3466 1.1392
R13253 VGND.n3452 VGND.n3451 1.1392
R13254 VGND.n2846 VGND.n2843 1.1392
R13255 VGND.n2829 VGND.n2828 1.1392
R13256 VGND.n2511 VGND.n2510 1.1392
R13257 VGND.n1998 VGND.n1995 1.1392
R13258 VGND.n1981 VGND.n1980 1.1392
R13259 VGND.n4879 VGND.n4876 1.1392
R13260 VGND.n4522 VGND.n4521 1.13717
R13261 VGND.n4181 VGND.n4180 1.13717
R13262 VGND.n3692 VGND.n3691 1.13717
R13263 VGND.n3668 VGND.n3667 1.13717
R13264 VGND.n3121 VGND.n3120 1.13717
R13265 VGND.n3101 VGND.n3100 1.13717
R13266 VGND.n2540 VGND.n2539 1.13717
R13267 VGND.n2271 VGND.n2270 1.13717
R13268 VGND.n2099 VGND.n2098 1.13717
R13269 VGND.n85 VGND.n84 1.13717
R13270 VGND.n4502 VGND.n4501 1.13717
R13271 VGND.n4192 VGND.n4191 1.1368
R13272 VGND.n376 VGND.n375 1.1368
R13273 VGND.n3683 VGND.n3682 1.1368
R13274 VGND.n746 VGND.n745 1.1368
R13275 VGND.n3112 VGND.n3111 1.1368
R13276 VGND.n1114 VGND.n1113 1.1368
R13277 VGND.n2531 VGND.n2530 1.1368
R13278 VGND.n2110 VGND.n2109 1.1368
R13279 VGND.n1508 VGND.n1507 1.1368
R13280 VGND.n5177 VGND.n5176 1.1368
R13281 VGND.n5453 VGND.n5452 1.1368
R13282 VGND.n279 VGND.n278 1.1368
R13283 VGND.n3998 VGND.n3997 1.1368
R13284 VGND.n616 VGND.n615 1.1368
R13285 VGND.n3465 VGND.n3464 1.1368
R13286 VGND.n1010 VGND.n1009 1.1368
R13287 VGND.n2842 VGND.n2841 1.1368
R13288 VGND.n1309 VGND.n1308 1.1368
R13289 VGND.n1458 VGND.n1457 1.1368
R13290 VGND.n1994 VGND.n1993 1.1368
R13291 VGND.n1841 VGND.n1840 1.1368
R13292 VGND.n4875 VGND.n4874 1.1368
R13293 VGND.n4523 VGND.n4522 1.13669
R13294 VGND.n4182 VGND.n4181 1.13669
R13295 VGND.n3693 VGND.n3692 1.13669
R13296 VGND.n3669 VGND.n3668 1.13669
R13297 VGND.n3122 VGND.n3121 1.13669
R13298 VGND.n3102 VGND.n3101 1.13669
R13299 VGND.n2541 VGND.n2540 1.13669
R13300 VGND.n2270 VGND.n2268 1.13669
R13301 VGND.n2100 VGND.n2099 1.13669
R13302 VGND.n86 VGND.n85 1.13669
R13303 VGND.n4513 VGND.n4496 1.13669
R13304 VGND.n4511 VGND.n4509 1.13669
R13305 VGND.n4865 VGND.n4864 1.13669
R13306 VGND.n607 VGND.n606 1.13669
R13307 VGND.n3990 VGND.n3989 1.13669
R13308 VGND.n1001 VGND.n1000 1.13669
R13309 VGND.n3457 VGND.n3456 1.13669
R13310 VGND.n1300 VGND.n1299 1.13669
R13311 VGND.n2834 VGND.n2833 1.13669
R13312 VGND.n2517 VGND.n2516 1.13669
R13313 VGND.n1834 VGND.n1833 1.13669
R13314 VGND.n1987 VGND.n1986 1.13669
R13315 VGND.n4333 VGND.n270 1.13669
R13316 VGND.n50 VGND.n49 1.13669
R13317 VGND.n4512 VGND.n4503 1.13648
R13318 VGND.n4052 VGND.n4051 1.09272
R13319 VGND.n408 VGND.n407 1.09272
R13320 VGND.n726 VGND.n651 1.09272
R13321 VGND.n3406 VGND.n3405 1.09272
R13322 VGND.n2943 VGND.n2895 1.09272
R13323 VGND.n2805 VGND.n1328 1.09272
R13324 VGND.n2200 VGND.n2173 1.09272
R13325 VGND.n1665 VGND.n1662 1.09272
R13326 VGND.n1630 VGND.n1629 1.09272
R13327 VGND.n192 VGND.n174 1.09272
R13328 VGND.n4681 VGND.n4680 1.09216
R13329 VGND.n319 VGND.n318 1.09216
R13330 VGND.n4569 VGND.n4568 1.09216
R13331 VGND.n418 VGND.n402 1.09216
R13332 VGND.n687 VGND.n669 1.09216
R13333 VGND.n3899 VGND.n3896 1.09216
R13334 VGND.n842 VGND.n841 1.09216
R13335 VGND.n1091 VGND.n1051 1.09216
R13336 VGND.n1415 VGND.n1347 1.09216
R13337 VGND.n1597 VGND.n1596 1.09216
R13338 VGND.n168 VGND.n133 1.09216
R13339 VGND.n206 VGND.n205 1.09216
R13340 VGND.n4226 VGND.n4225 1.09216
R13341 VGND.n4295 VGND.n4207 1.09216
R13342 VGND.n4916 VGND.n255 1.09216
R13343 VGND.n4964 VGND.n254 1.09216
R13344 VGND.n4420 VGND.n4419 1.08588
R13345 VGND.n4255 VGND.n4254 1.08588
R13346 VGND.n1632 VGND.n1538 1.08588
R13347 VGND.n2867 VGND.n1275 1.08588
R13348 VGND.n2167 VGND.n2124 1.08588
R13349 VGND VGND.n4024 1.02178
R13350 VGND.n2887 VGND 1.02178
R13351 VGND.n2484 VGND.n2483 1.00931
R13352 VGND.n2562 VGND.n2561 0.953691
R13353 VGND.n1583 VGND.n1582 0.882934
R13354 VGND.n4859 VGND.n4858 0.872922
R13355 VGND.n4003 VGND.n4002 0.872922
R13356 VGND.n3984 VGND.n3983 0.872922
R13357 VGND.n3470 VGND.n3469 0.872922
R13358 VGND.n3451 VGND.n3450 0.872922
R13359 VGND.n2847 VGND.n2846 0.872922
R13360 VGND.n2828 VGND.n2827 0.872922
R13361 VGND.n2510 VGND.n2509 0.872922
R13362 VGND.n1999 VGND.n1998 0.872922
R13363 VGND.n1980 VGND.n1979 0.872922
R13364 VGND.n4880 VGND.n4879 0.872922
R13365 VGND.n5456 VGND.n5455 0.871525
R13366 VGND.n4719 VGND.n273 0.871338
R13367 VGND.n600 VGND.n599 0.871338
R13368 VGND.n3857 VGND.n610 0.871338
R13369 VGND.n995 VGND.n994 0.871338
R13370 VGND.n3320 VGND.n1004 0.871338
R13371 VGND.n2959 VGND.n1262 0.871338
R13372 VGND.n2706 VGND.n1303 0.871338
R13373 VGND.n2371 VGND.n1453 0.871338
R13374 VGND.n1826 VGND.n1825 0.871338
R13375 VGND.n5032 VGND.n119 0.871338
R13376 VGND.n5447 VGND.n5446 0.871338
R13377 VGND.n4344 VGND.n4334 0.86965
R13378 VGND.n5168 VGND.n5167 0.867431
R13379 VGND.n2091 VGND.n2090 0.867431
R13380 VGND.n2266 VGND.n2265 0.867431
R13381 VGND.n2546 VGND.n2545 0.867431
R13382 VGND.n3093 VGND.n3092 0.867431
R13383 VGND.n3127 VGND.n3126 0.867431
R13384 VGND.n3660 VGND.n3659 0.867431
R13385 VGND.n3698 VGND.n3697 0.867431
R13386 VGND.n4173 VGND.n4172 0.867431
R13387 VGND.n4528 VGND.n4527 0.867431
R13388 VGND.n5199 VGND.n5198 0.867431
R13389 VGND.n4493 VGND.n4492 0.865744
R13390 VGND.n65 VGND.n62 0.833377
R13391 VGND.n71 VGND.n68 0.833377
R13392 VGND.n5328 VGND.n5327 0.833377
R13393 VGND.n4948 VGND.n4947 0.833377
R13394 VGND.n1680 VGND.n1679 0.833377
R13395 VGND.n4813 VGND.n4812 0.833377
R13396 VGND.n3964 VGND.n3963 0.833377
R13397 VGND.n3816 VGND.n3813 0.833377
R13398 VGND.n3836 VGND.n3833 0.833377
R13399 VGND.n831 VGND.n828 0.833377
R13400 VGND.n780 VGND.n777 0.833377
R13401 VGND.n918 VGND.n917 0.833377
R13402 VGND.n1037 VGND.n1034 0.833377
R13403 VGND.n2762 VGND.n2761 0.833377
R13404 VGND.n2803 VGND.n2802 0.833377
R13405 VGND.n2584 VGND.n2581 0.833377
R13406 VGND.n2482 VGND.n1473 0.833377
R13407 VGND.n1873 VGND.n1872 0.833377
R13408 VGND.n5045 VGND.n5044 0.833377
R13409 VGND.n5555 VGND.n5554 0.833377
R13410 VGND.n3235 VGND.n3234 0.8005
R13411 VGND.n5269 VGND.n5268 0.753441
R13412 VGND.n4284 VGND.n4283 0.746688
R13413 VGND.n3674 VGND.n3673 0.668275
R13414 VGND.n2522 VGND.n2521 0.668275
R13415 VGND.n5038 VGND.n5037 0.614199
R13416 VGND.n3155 VGND.n3154 0.561904
R13417 VGND.n1129 VGND.n1128 0.561904
R13418 VGND.n5400 VGND.n5399 0.526527
R13419 VGND.n5379 VGND.n5378 0.526527
R13420 VGND.n5323 VGND.n5322 0.526527
R13421 VGND.n4951 VGND.n4950 0.526527
R13422 VGND.n1683 VGND.n1682 0.526527
R13423 VGND.n4816 VGND.n4815 0.526527
R13424 VGND.n3967 VGND.n3966 0.526527
R13425 VGND.n3812 VGND.n3811 0.526527
R13426 VGND.n3832 VGND.n3831 0.526527
R13427 VGND.n857 VGND.n856 0.526527
R13428 VGND.n795 VGND.n794 0.526527
R13429 VGND.n920 VGND.n919 0.526527
R13430 VGND.n3282 VGND.n3281 0.526527
R13431 VGND.n2765 VGND.n2764 0.526527
R13432 VGND.n2616 VGND.n2615 0.526527
R13433 VGND.n1949 VGND.n1874 0.526527
R13434 VGND.n5048 VGND.n5047 0.526527
R13435 VGND.n5558 VGND.n5557 0.526527
R13436 VGND.n1130 VGND.n1129 0.524477
R13437 VGND.n3673 VGND 0.478275
R13438 VGND.n2521 VGND 0.478275
R13439 VGND.n5229 VGND.n5228 0.438856
R13440 VGND.n5240 VGND.n5239 0.438856
R13441 VGND.n1572 VGND.n1570 0.438856
R13442 VGND.n407 VGND.n406 0.407316
R13443 VGND.n318 VGND.n317 0.404857
R13444 VGND.n841 VGND.n840 0.404857
R13445 VGND.n1596 VGND.n1595 0.404857
R13446 VGND.n4225 VGND.n4224 0.404857
R13447 VGND.n3230 VGND.n3229 0.4005
R13448 VGND.n193 VGND.n192 0.356503
R13449 VGND.n4051 VGND.n4048 0.2965
R13450 VGND.n2201 VGND.n2200 0.2965
R13451 VGND.n1666 VGND.n1665 0.2965
R13452 VGND.n4680 VGND.n4679 0.294041
R13453 VGND.n168 VGND.n167 0.294041
R13454 VGND.n207 VGND.n206 0.294041
R13455 VGND.n4295 VGND.n4294 0.294041
R13456 VGND.n4269 VGND.n4268 0.287496
R13457 VGND.n4282 VGND.n4281 0.287496
R13458 VGND.n726 VGND 0.275667
R13459 VGND.n3405 VGND 0.274365
R13460 VGND VGND.n4569 0.271905
R13461 VGND.n418 VGND 0.271905
R13462 VGND.n1091 VGND 0.271905
R13463 VGND.n1415 VGND 0.271905
R13464 VGND.n4916 VGND 0.271905
R13465 VGND VGND.n2805 0.26525
R13466 VGND.n1629 VGND 0.26525
R13467 VGND VGND.n2943 0.263948
R13468 VGND VGND.n669 0.262791
R13469 VGND VGND.n3899 0.262791
R13470 VGND VGND.n4964 0.261489
R13471 VGND.n3855 VGND.n3854 0.253789
R13472 VGND.n3318 VGND.n3317 0.253789
R13473 VGND.n699 VGND.n698 0.239569
R13474 VGND.n3928 VGND.n3927 0.239569
R13475 VGND.n3225 VGND.n3224 0.239569
R13476 VGND.n1222 VGND.n1221 0.239569
R13477 VGND.n2747 VGND.n2746 0.239569
R13478 VGND.n2296 VGND.n2295 0.239569
R13479 VGND.n2341 VGND.n2340 0.239569
R13480 VGND.n2503 VGND.n2501 0.239569
R13481 VGND.n2034 VGND.n2032 0.239569
R13482 VGND.n1700 VGND.n1698 0.239569
R13483 VGND.n1902 VGND.n1900 0.239569
R13484 VGND.n4406 VGND.n4405 0.239569
R13485 VGND.n4908 VGND.n4907 0.239569
R13486 VGND.n4931 VGND.n4930 0.239569
R13487 VGND.n5366 VGND.n5365 0.239569
R13488 VGND.n5577 VGND.n5575 0.239569
R13489 VGND.n2038 VGND.n2037 0.239393
R13490 VGND.n1161 VGND.n1160 0.238519
R13491 VGND.n3246 VGND.n3245 0.238116
R13492 VGND.n454 VGND.n452 0.237885
R13493 VGND.n5083 VGND.n5081 0.237885
R13494 VGND.n5523 VGND.n5521 0.237885
R13495 VGND.n678 VGND.n674 0.231108
R13496 VGND.n1059 VGND.n1057 0.231108
R13497 VGND.n1153 VGND.n1152 0.231108
R13498 VGND.n1366 VGND.n1365 0.231108
R13499 VGND.n2137 VGND.n2134 0.231108
R13500 VGND.n140 VGND.n138 0.231108
R13501 VGND.n4659 VGND 0.217434
R13502 VGND.n4017 VGND 0.217434
R13503 VGND.n4032 VGND 0.217434
R13504 VGND.n4038 VGND 0.217434
R13505 VGND.n536 VGND 0.217434
R13506 VGND.n3473 VGND 0.217434
R13507 VGND VGND.n3361 0.217434
R13508 VGND.n1160 VGND 0.217434
R13509 VGND.n2894 VGND 0.217434
R13510 VGND.n2592 VGND 0.217434
R13511 VGND.n1783 VGND 0.217434
R13512 VGND VGND.n1730 0.217434
R13513 VGND.n1708 VGND 0.217434
R13514 VGND.n5089 VGND 0.217434
R13515 VGND.n154 VGND 0.217434
R13516 VGND.n4234 VGND 0.217434
R13517 VGND.n4287 VGND 0.217434
R13518 VGND.n4288 VGND 0.217434
R13519 VGND.n4759 VGND 0.215749
R13520 VGND VGND.n448 0.215749
R13521 VGND VGND.n4050 0.215749
R13522 VGND VGND.n3898 0.215749
R13523 VGND VGND.n807 0.215749
R13524 VGND VGND.n3360 0.215749
R13525 VGND VGND.n2745 0.215749
R13526 VGND.n2139 VGND 0.215749
R13527 VGND VGND.n1664 0.215749
R13528 VGND VGND.n4929 0.215749
R13529 VGND.n548 VGND 0.208319
R13530 VGND.n679 VGND 0.208319
R13531 VGND.n719 VGND 0.208319
R13532 VGND.n808 VGND 0.208319
R13533 VGND.n1060 VGND 0.208319
R13534 VGND.n2138 VGND 0.208319
R13535 VGND VGND.n1721 0.208319
R13536 VGND.n2784 VGND 0.207017
R13537 VGND.n2650 VGND 0.207017
R13538 VGND.n2908 VGND 0.206635
R13539 VGND.n2424 VGND 0.206635
R13540 VGND.n1157 VGND 0.205715
R13541 VGND VGND.n2605 0.205715
R13542 VGND.n4717 VGND.n4716 0.204755
R13543 VGND.n597 VGND.n596 0.204755
R13544 VGND.n992 VGND.n991 0.204755
R13545 VGND.n2961 VGND.n2960 0.204755
R13546 VGND.n2704 VGND.n2703 0.204755
R13547 VGND.n2369 VGND.n2368 0.204755
R13548 VGND.n1823 VGND.n1822 0.204755
R13549 VGND VGND.n3525 0.204031
R13550 VGND VGND.n1889 0.204031
R13551 VGND.n448 VGND.n380 0.201782
R13552 VGND.n407 VGND 0.196835
R13553 VGND.n4051 VGND 0.196835
R13554 VGND VGND.n726 0.196835
R13555 VGND.n3405 VGND 0.196835
R13556 VGND.n2943 VGND 0.196835
R13557 VGND.n2805 VGND 0.196835
R13558 VGND.n2200 VGND 0.196835
R13559 VGND.n1629 VGND 0.196835
R13560 VGND.n1665 VGND 0.196835
R13561 VGND.n192 VGND 0.196835
R13562 VGND.n318 VGND 0.196385
R13563 VGND.n4569 VGND 0.196385
R13564 VGND.n4680 VGND 0.196385
R13565 VGND VGND.n418 0.196385
R13566 VGND.n669 VGND 0.196385
R13567 VGND.n3899 VGND 0.196385
R13568 VGND.n841 VGND 0.196385
R13569 VGND VGND.n1091 0.196385
R13570 VGND VGND.n1415 0.196385
R13571 VGND.n1596 VGND 0.196385
R13572 VGND VGND.n168 0.196385
R13573 VGND.n206 VGND 0.196385
R13574 VGND.n4225 VGND 0.196385
R13575 VGND VGND.n4295 0.196385
R13576 VGND VGND.n4916 0.196385
R13577 VGND.n4964 VGND 0.196385
R13578 VGND.n3673 VGND.n3672 0.1905
R13579 VGND.n2521 VGND.n2520 0.1905
R13580 VGND.n1633 VGND.n1534 0.185802
R13581 VGND.n4779 VGND.n4778 0.180551
R13582 VGND.n561 VGND.n560 0.180551
R13583 VGND.n4008 VGND.n4007 0.180551
R13584 VGND.n3850 VGND.n3846 0.180551
R13585 VGND.n1073 VGND.n1070 0.180551
R13586 VGND.n2825 VGND.n2822 0.180551
R13587 VGND.n1376 VGND.n1375 0.180551
R13588 VGND.n2048 VGND.n2046 0.180551
R13589 VGND.n1573 VGND.n1567 0.180551
R13590 VGND.n194 VGND.n193 0.180551
R13591 VGND.n459 VGND.n458 0.180294
R13592 VGND.n2889 VGND 0.16102
R13593 VGND.n3975 VGND 0.159717
R13594 VGND.n737 VGND 0.159717
R13595 VGND.n2313 VGND 0.159717
R13596 VGND.n294 VGND 0.158415
R13597 VGND VGND.n4551 0.158415
R13598 VGND.n3851 VGND 0.158415
R13599 VGND.n3514 VGND 0.158415
R13600 VGND.n2781 VGND 0.158415
R13601 VGND.n2144 VGND 0.158415
R13602 VGND.n1604 VGND 0.158415
R13603 VGND.n1608 VGND 0.158415
R13604 VGND VGND.n1566 0.158415
R13605 VGND.n169 VGND 0.158415
R13606 VGND.n200 VGND 0.158415
R13607 VGND.n4885 VGND 0.158415
R13608 VGND VGND.n1491 0.158159
R13609 VGND.n411 VGND 0.15779
R13610 VGND VGND.n3184 0.15779
R13611 VGND.n459 VGND 0.157113
R13612 VGND.n3062 VGND.n3061 0.155186
R13613 VGND.n5179 VGND.n5178 0.151488
R13614 VGND.n1500 VGND.n1499 0.151488
R13615 VGND.n2102 VGND.n2101 0.151488
R13616 VGND.n2533 VGND.n2532 0.151488
R13617 VGND.n3104 VGND.n3103 0.151488
R13618 VGND.n3114 VGND.n3113 0.151488
R13619 VGND.n3685 VGND.n3684 0.151488
R13620 VGND.n4184 VGND.n4183 0.151488
R13621 VGND.n4515 VGND.n4514 0.151488
R13622 VGND.n1836 VGND.n1835 0.151488
R13623 VGND.n1989 VGND.n1988 0.151488
R13624 VGND.n1828 VGND.n1827 0.151488
R13625 VGND.n2836 VGND.n2835 0.151488
R13626 VGND.n1295 VGND.n1294 0.151488
R13627 VGND.n3459 VGND.n3458 0.151488
R13628 VGND.n3992 VGND.n3991 0.151488
R13629 VGND.n602 VGND.n601 0.151488
R13630 VGND.n4867 VGND.n4866 0.151488
R13631 VGND VGND.n2592 0.149977
R13632 VGND VGND.n4097 0.149301
R13633 VGND.n4027 VGND 0.149301
R13634 VGND VGND.n464 0.149301
R13635 VGND VGND.n3935 0.149301
R13636 VGND.n3241 VGND 0.149301
R13637 VGND VGND.n3185 0.149301
R13638 VGND.n1616 VGND 0.149301
R13639 VGND.n4407 VGND 0.149301
R13640 VGND.n3803 VGND 0.147999
R13641 VGND.n4260 VGND 0.147999
R13642 VGND.n2621 VGND 0.146697
R13643 VGND.n1371 VGND 0.146697
R13644 VGND.n738 VGND.n737 0.143836
R13645 VGND VGND.n3246 0.141328
R13646 VGND.n2037 VGND 0.141026
R13647 VGND VGND.n4659 0.140863
R13648 VGND VGND.n548 0.140863
R13649 VGND VGND.n4017 0.140863
R13650 VGND VGND.n4032 0.140863
R13651 VGND VGND.n4038 0.140863
R13652 VGND VGND.n536 0.140863
R13653 VGND VGND.n679 0.140863
R13654 VGND.n699 VGND 0.140863
R13655 VGND VGND.n719 0.140863
R13656 VGND.n3927 VGND 0.140863
R13657 VGND.n808 VGND 0.140863
R13658 VGND.n3473 VGND 0.140863
R13659 VGND.n3225 VGND 0.140863
R13660 VGND.n1060 VGND 0.140863
R13661 VGND.n3361 VGND 0.140863
R13662 VGND.n1157 VGND 0.140863
R13663 VGND.n1221 VGND 0.140863
R13664 VGND VGND.n2894 0.140863
R13665 VGND.n2605 VGND 0.140863
R13666 VGND.n2784 VGND 0.140863
R13667 VGND.n2746 VGND 0.140863
R13668 VGND VGND.n2650 0.140863
R13669 VGND VGND.n2296 0.140863
R13670 VGND VGND.n2341 0.140863
R13671 VGND VGND.n2138 0.140863
R13672 VGND.n2501 VGND 0.140863
R13673 VGND.n2032 VGND 0.140863
R13674 VGND VGND.n1783 0.140863
R13675 VGND.n1730 VGND 0.140863
R13676 VGND.n1721 VGND 0.140863
R13677 VGND.n1708 VGND 0.140863
R13678 VGND.n1698 VGND 0.140863
R13679 VGND.n5089 VGND 0.140863
R13680 VGND.n154 VGND 0.140863
R13681 VGND.n1900 VGND 0.140863
R13682 VGND.n4234 VGND 0.140863
R13683 VGND VGND.n4287 0.140863
R13684 VGND VGND.n4288 0.140863
R13685 VGND VGND.n4908 0.140863
R13686 VGND.n4930 VGND 0.140863
R13687 VGND VGND.n5366 0.140863
R13688 VGND.n5575 VGND 0.140863
R13689 VGND.n4759 VGND 0.140584
R13690 VGND.n452 VGND 0.140584
R13691 VGND.n4050 VGND 0.140584
R13692 VGND.n3898 VGND 0.140584
R13693 VGND.n807 VGND 0.140584
R13694 VGND.n3525 VGND 0.140584
R13695 VGND.n3360 VGND 0.140584
R13696 VGND.n2908 VGND 0.140584
R13697 VGND.n2745 VGND 0.140584
R13698 VGND VGND.n2139 0.140584
R13699 VGND.n2424 VGND 0.140584
R13700 VGND.n1664 VGND 0.140584
R13701 VGND.n5081 VGND 0.140584
R13702 VGND.n1889 VGND 0.140584
R13703 VGND.n4929 VGND 0.140584
R13704 VGND.n5521 VGND 0.140584
R13705 VGND.n3472 VGND.n3471 0.137582
R13706 VGND.n4884 VGND.n4881 0.137582
R13707 VGND.n5438 VGND.n5437 0.13667
R13708 VGND.n4361 VGND.n4360 0.13667
R13709 VGND.n2085 VGND.n2084 0.13667
R13710 VGND.n3654 VGND.n3653 0.13667
R13711 VGND.n2557 VGND.n2556 0.13667
R13712 VGND.n5162 VGND.n5161 0.13667
R13713 VGND.n4301 VGND.n4300 0.136287
R13714 VGND.n5037 VGND.n5036 0.132007
R13715 VGND.n323 VGND.n321 0.120292
R13716 VGND.n325 VGND.n323 0.120292
R13717 VGND.n331 VGND.n329 0.120292
R13718 VGND.n333 VGND.n331 0.120292
R13719 VGND.n334 VGND.n333 0.120292
R13720 VGND.n335 VGND.n334 0.120292
R13721 VGND.n336 VGND.n335 0.120292
R13722 VGND.n341 VGND.n339 0.120292
R13723 VGND.n343 VGND.n341 0.120292
R13724 VGND.n345 VGND.n343 0.120292
R13725 VGND.n346 VGND.n345 0.120292
R13726 VGND.n351 VGND.n349 0.120292
R13727 VGND.n352 VGND.n351 0.120292
R13728 VGND.n353 VGND.n352 0.120292
R13729 VGND.n4585 VGND.n4584 0.120292
R13730 VGND.n4584 VGND.n4582 0.120292
R13731 VGND.n4582 VGND.n4581 0.120292
R13732 VGND.n4577 VGND.n4576 0.120292
R13733 VGND.n4576 VGND.n4574 0.120292
R13734 VGND.n4570 VGND.n358 0.120292
R13735 VGND.n4565 VGND.n4564 0.120292
R13736 VGND.n4564 VGND.n4562 0.120292
R13737 VGND.n4562 VGND.n4560 0.120292
R13738 VGND.n4560 VGND.n4558 0.120292
R13739 VGND.n4558 VGND.n4557 0.120292
R13740 VGND.n4552 VGND.n364 0.120292
R13741 VGND.n4615 VGND.n4612 0.120292
R13742 VGND.n4616 VGND.n4615 0.120292
R13743 VGND.n4621 VGND.n4619 0.120292
R13744 VGND.n4623 VGND.n4621 0.120292
R13745 VGND.n4625 VGND.n4623 0.120292
R13746 VGND.n4627 VGND.n4625 0.120292
R13747 VGND.n4629 VGND.n4627 0.120292
R13748 VGND.n4631 VGND.n4629 0.120292
R13749 VGND.n4633 VGND.n4631 0.120292
R13750 VGND.n4635 VGND.n4633 0.120292
R13751 VGND.n4637 VGND.n4635 0.120292
R13752 VGND.n4639 VGND.n4637 0.120292
R13753 VGND.n4641 VGND.n4639 0.120292
R13754 VGND.n4643 VGND.n4641 0.120292
R13755 VGND.n4645 VGND.n4643 0.120292
R13756 VGND.n4646 VGND.n4645 0.120292
R13757 VGND.n4651 VGND.n4650 0.120292
R13758 VGND.n4653 VGND.n4651 0.120292
R13759 VGND.n4657 VGND.n4653 0.120292
R13760 VGND.n4658 VGND.n4657 0.120292
R13761 VGND.n4672 VGND.n4671 0.120292
R13762 VGND.n4677 VGND.n4675 0.120292
R13763 VGND.n4679 VGND.n4677 0.120292
R13764 VGND.n4685 VGND.n4683 0.120292
R13765 VGND.n4687 VGND.n4685 0.120292
R13766 VGND.n4689 VGND.n4687 0.120292
R13767 VGND.n4691 VGND.n4689 0.120292
R13768 VGND.n4693 VGND.n4691 0.120292
R13769 VGND.n4695 VGND.n4693 0.120292
R13770 VGND.n4697 VGND.n4695 0.120292
R13771 VGND.n4699 VGND.n4697 0.120292
R13772 VGND.n4701 VGND.n4699 0.120292
R13773 VGND.n4702 VGND.n4701 0.120292
R13774 VGND.n4707 VGND.n4705 0.120292
R13775 VGND.n4710 VGND.n4707 0.120292
R13776 VGND.n4856 VGND.n4854 0.120292
R13777 VGND.n4854 VGND.n4851 0.120292
R13778 VGND.n4848 VGND.n4847 0.120292
R13779 VGND.n4847 VGND.n4845 0.120292
R13780 VGND.n4842 VGND.n4841 0.120292
R13781 VGND.n4841 VGND.n4840 0.120292
R13782 VGND.n4840 VGND.n4837 0.120292
R13783 VGND.n4834 VGND.n4833 0.120292
R13784 VGND.n4833 VGND.n4832 0.120292
R13785 VGND.n4829 VGND.n4828 0.120292
R13786 VGND.n4828 VGND.n4827 0.120292
R13787 VGND.n4821 VGND.n4820 0.120292
R13788 VGND.n4820 VGND.n4819 0.120292
R13789 VGND.n4819 VGND.n4817 0.120292
R13790 VGND.n4817 VGND.n4814 0.120292
R13791 VGND.n4814 VGND.n4809 0.120292
R13792 VGND.n4809 VGND.n4806 0.120292
R13793 VGND.n4802 VGND.n4801 0.120292
R13794 VGND.n4801 VGND.n4800 0.120292
R13795 VGND.n4800 VGND.n4797 0.120292
R13796 VGND.n4793 VGND.n4792 0.120292
R13797 VGND.n4792 VGND.n4791 0.120292
R13798 VGND.n4791 VGND.n4789 0.120292
R13799 VGND.n4789 VGND.n4787 0.120292
R13800 VGND.n4787 VGND.n4784 0.120292
R13801 VGND.n4780 VGND.n4779 0.120292
R13802 VGND.n4774 VGND.n4773 0.120292
R13803 VGND.n4773 VGND.n4771 0.120292
R13804 VGND.n4771 VGND 0.120292
R13805 VGND.n4764 VGND.n4758 0.120292
R13806 VGND VGND.n412 0.120292
R13807 VGND.n417 VGND.n403 0.120292
R13808 VGND.n424 VGND.n422 0.120292
R13809 VGND.n426 VGND.n424 0.120292
R13810 VGND.n428 VGND.n426 0.120292
R13811 VGND.n429 VGND.n428 0.120292
R13812 VGND.n434 VGND.n432 0.120292
R13813 VGND.n435 VGND.n434 0.120292
R13814 VGND.n436 VGND.n435 0.120292
R13815 VGND.n481 VGND.n480 0.120292
R13816 VGND.n480 VGND.n478 0.120292
R13817 VGND.n478 VGND.n477 0.120292
R13818 VGND.n473 VGND.n472 0.120292
R13819 VGND.n472 VGND.n470 0.120292
R13820 VGND.n470 VGND.n468 0.120292
R13821 VGND.n455 VGND.n454 0.120292
R13822 VGND.n451 VGND.n450 0.120292
R13823 VGND.n450 VGND.n449 0.120292
R13824 VGND.n4140 VGND 0.120292
R13825 VGND.n4135 VGND.n4134 0.120292
R13826 VGND.n4134 VGND.n4133 0.120292
R13827 VGND.n4130 VGND.n4129 0.120292
R13828 VGND.n4129 VGND.n4127 0.120292
R13829 VGND.n4127 VGND.n4125 0.120292
R13830 VGND.n4125 VGND.n4123 0.120292
R13831 VGND.n4123 VGND.n4121 0.120292
R13832 VGND.n4121 VGND.n4119 0.120292
R13833 VGND.n4119 VGND.n4117 0.120292
R13834 VGND.n4114 VGND.n4113 0.120292
R13835 VGND.n4113 VGND.n4112 0.120292
R13836 VGND.n4112 VGND.n4109 0.120292
R13837 VGND.n4106 VGND.n4105 0.120292
R13838 VGND.n4105 VGND.n4103 0.120292
R13839 VGND.n4103 VGND.n4101 0.120292
R13840 VGND.n530 VGND.n529 0.120292
R13841 VGND.n531 VGND.n530 0.120292
R13842 VGND VGND.n531 0.120292
R13843 VGND.n542 VGND.n540 0.120292
R13844 VGND.n544 VGND.n542 0.120292
R13845 VGND.n547 VGND.n544 0.120292
R13846 VGND.n554 VGND.n552 0.120292
R13847 VGND.n556 VGND.n554 0.120292
R13848 VGND.n558 VGND.n556 0.120292
R13849 VGND.n560 VGND.n558 0.120292
R13850 VGND.n4015 VGND.n4014 0.120292
R13851 VGND.n4016 VGND.n4015 0.120292
R13852 VGND.n4022 VGND.n4021 0.120292
R13853 VGND.n4034 VGND.n4033 0.120292
R13854 VGND.n4088 VGND.n4087 0.120292
R13855 VGND.n4087 VGND.n4039 0.120292
R13856 VGND.n4082 VGND.n4039 0.120292
R13857 VGND.n4080 VGND.n4041 0.120292
R13858 VGND.n4076 VGND.n4041 0.120292
R13859 VGND.n4076 VGND.n4075 0.120292
R13860 VGND.n4075 VGND.n4074 0.120292
R13861 VGND.n4074 VGND.n4043 0.120292
R13862 VGND.n4069 VGND.n4068 0.120292
R13863 VGND.n4068 VGND.n4067 0.120292
R13864 VGND.n4064 VGND.n4063 0.120292
R13865 VGND.n4063 VGND.n4062 0.120292
R13866 VGND.n4062 VGND.n4046 0.120292
R13867 VGND.n4056 VGND.n4048 0.120292
R13868 VGND.n684 VGND.n683 0.120292
R13869 VGND VGND.n684 0.120292
R13870 VGND.n668 VGND.n667 0.120292
R13871 VGND.n667 VGND.n666 0.120292
R13872 VGND.n692 VGND.n666 0.120292
R13873 VGND.n693 VGND.n692 0.120292
R13874 VGND.n694 VGND.n664 0.120292
R13875 VGND.n698 VGND.n664 0.120292
R13876 VGND.n706 VGND.n705 0.120292
R13877 VGND.n706 VGND.n661 0.120292
R13878 VGND.n711 VGND.n661 0.120292
R13879 VGND.n713 VGND.n659 0.120292
R13880 VGND.n659 VGND.n658 0.120292
R13881 VGND.n721 VGND.n652 0.120292
R13882 VGND.n725 VGND.n652 0.120292
R13883 VGND.n728 VGND.n649 0.120292
R13884 VGND.n732 VGND.n649 0.120292
R13885 VGND.n3780 VGND.n3779 0.120292
R13886 VGND.n3779 VGND.n3778 0.120292
R13887 VGND.n3778 VGND.n3775 0.120292
R13888 VGND.n3772 VGND.n3771 0.120292
R13889 VGND.n3771 VGND.n3769 0.120292
R13890 VGND.n3769 VGND.n3767 0.120292
R13891 VGND.n3767 VGND.n3765 0.120292
R13892 VGND.n3765 VGND.n3763 0.120292
R13893 VGND.n3763 VGND.n3761 0.120292
R13894 VGND.n3761 VGND.n3759 0.120292
R13895 VGND.n3756 VGND.n3755 0.120292
R13896 VGND.n3755 VGND.n3754 0.120292
R13897 VGND.n3754 VGND.n3751 0.120292
R13898 VGND.n3748 VGND.n3747 0.120292
R13899 VGND.n3747 VGND.n3745 0.120292
R13900 VGND.n3741 VGND.n3739 0.120292
R13901 VGND.n3739 VGND.n3737 0.120292
R13902 VGND.n3737 VGND.n3735 0.120292
R13903 VGND.n3735 VGND.n3734 0.120292
R13904 VGND.n3808 VGND.n3806 0.120292
R13905 VGND.n3809 VGND.n3808 0.120292
R13906 VGND.n3810 VGND.n3809 0.120292
R13907 VGND.n3818 VGND.n3810 0.120292
R13908 VGND.n3824 VGND.n3822 0.120292
R13909 VGND.n3826 VGND.n3824 0.120292
R13910 VGND.n3828 VGND.n3826 0.120292
R13911 VGND.n3829 VGND.n3828 0.120292
R13912 VGND.n3830 VGND.n3829 0.120292
R13913 VGND.n3838 VGND.n3830 0.120292
R13914 VGND.n3844 VGND.n3842 0.120292
R13915 VGND.n3845 VGND.n3844 0.120292
R13916 VGND.n3846 VGND.n3845 0.120292
R13917 VGND.n3981 VGND.n3979 0.120292
R13918 VGND.n3979 VGND.n3977 0.120292
R13919 VGND.n3974 VGND.n3973 0.120292
R13920 VGND.n3973 VGND.n3972 0.120292
R13921 VGND.n3972 VGND.n3970 0.120292
R13922 VGND.n3970 VGND.n3968 0.120292
R13923 VGND.n3968 VGND.n3965 0.120292
R13924 VGND.n3965 VGND.n3960 0.120292
R13925 VGND.n3960 VGND.n3957 0.120292
R13926 VGND.n3954 VGND.n3953 0.120292
R13927 VGND.n3953 VGND.n3952 0.120292
R13928 VGND.n3952 VGND.n3949 0.120292
R13929 VGND.n3946 VGND.n3945 0.120292
R13930 VGND.n3945 VGND.n3943 0.120292
R13931 VGND.n3943 VGND.n3941 0.120292
R13932 VGND.n3941 VGND.n3940 0.120292
R13933 VGND.n3929 VGND.n3928 0.120292
R13934 VGND.n3926 VGND.n3925 0.120292
R13935 VGND.n3925 VGND.n3923 0.120292
R13936 VGND.n3923 VGND.n3921 0.120292
R13937 VGND.n3921 VGND.n3919 0.120292
R13938 VGND.n3919 VGND.n3917 0.120292
R13939 VGND.n3917 VGND.n3915 0.120292
R13940 VGND.n3915 VGND.n3914 0.120292
R13941 VGND.n3911 VGND.n3910 0.120292
R13942 VGND.n3910 VGND.n3909 0.120292
R13943 VGND.n3909 VGND.n3894 0.120292
R13944 VGND.n3904 VGND.n3903 0.120292
R13945 VGND.n846 VGND.n844 0.120292
R13946 VGND.n847 VGND.n846 0.120292
R13947 VGND VGND.n847 0.120292
R13948 VGND.n852 VGND.n851 0.120292
R13949 VGND.n853 VGND.n852 0.120292
R13950 VGND.n854 VGND.n853 0.120292
R13951 VGND.n859 VGND.n858 0.120292
R13952 VGND.n860 VGND.n859 0.120292
R13953 VGND.n861 VGND.n860 0.120292
R13954 VGND.n866 VGND.n864 0.120292
R13955 VGND.n867 VGND.n866 0.120292
R13956 VGND.n872 VGND.n870 0.120292
R13957 VGND.n873 VGND.n872 0.120292
R13958 VGND.n874 VGND.n873 0.120292
R13959 VGND.n823 VGND.n821 0.120292
R13960 VGND.n821 VGND.n819 0.120292
R13961 VGND.n819 VGND.n818 0.120292
R13962 VGND.n815 VGND.n814 0.120292
R13963 VGND.n814 VGND.n813 0.120292
R13964 VGND.n803 VGND.n802 0.120292
R13965 VGND.n802 VGND.n800 0.120292
R13966 VGND.n800 VGND.n798 0.120292
R13967 VGND.n798 VGND.n796 0.120292
R13968 VGND.n796 VGND.n793 0.120292
R13969 VGND.n793 VGND.n792 0.120292
R13970 VGND.n792 VGND.n791 0.120292
R13971 VGND.n788 VGND.n787 0.120292
R13972 VGND.n787 VGND.n785 0.120292
R13973 VGND.n3624 VGND.n3623 0.120292
R13974 VGND.n3623 VGND.n3620 0.120292
R13975 VGND.n3617 VGND.n3616 0.120292
R13976 VGND.n3616 VGND.n3614 0.120292
R13977 VGND.n3614 VGND.n3612 0.120292
R13978 VGND.n3612 VGND.n3610 0.120292
R13979 VGND.n3610 VGND.n3608 0.120292
R13980 VGND.n3608 VGND.n3606 0.120292
R13981 VGND.n3606 VGND.n3604 0.120292
R13982 VGND.n3604 VGND.n3602 0.120292
R13983 VGND.n762 VGND.n760 0.120292
R13984 VGND.n3592 VGND.n3591 0.120292
R13985 VGND.n3589 VGND.n3587 0.120292
R13986 VGND.n3587 VGND.n3585 0.120292
R13987 VGND.n3585 VGND.n3583 0.120292
R13988 VGND.n3583 VGND.n3581 0.120292
R13989 VGND.n910 VGND.n909 0.120292
R13990 VGND.n911 VGND.n910 0.120292
R13991 VGND.n912 VGND.n911 0.120292
R13992 VGND.n923 VGND.n922 0.120292
R13993 VGND.n924 VGND.n923 0.120292
R13994 VGND.n929 VGND.n927 0.120292
R13995 VGND.n931 VGND.n929 0.120292
R13996 VGND.n933 VGND.n931 0.120292
R13997 VGND.n935 VGND.n933 0.120292
R13998 VGND.n936 VGND.n935 0.120292
R13999 VGND.n937 VGND.n936 0.120292
R14000 VGND.n942 VGND.n940 0.120292
R14001 VGND.n943 VGND.n942 0.120292
R14002 VGND.n944 VGND.n943 0.120292
R14003 VGND.n949 VGND.n947 0.120292
R14004 VGND.n951 VGND.n949 0.120292
R14005 VGND.n953 VGND.n951 0.120292
R14006 VGND.n954 VGND.n953 0.120292
R14007 VGND.n959 VGND.n957 0.120292
R14008 VGND.n962 VGND.n959 0.120292
R14009 VGND.n3478 VGND.n3476 0.120292
R14010 VGND.n3480 VGND.n3478 0.120292
R14011 VGND.n3482 VGND.n3480 0.120292
R14012 VGND.n3484 VGND.n3482 0.120292
R14013 VGND.n3485 VGND.n3484 0.120292
R14014 VGND.n3490 VGND.n3489 0.120292
R14015 VGND.n3492 VGND.n3490 0.120292
R14016 VGND.n3499 VGND.n3498 0.120292
R14017 VGND.n3500 VGND.n3499 0.120292
R14018 VGND.n3504 VGND.n3503 0.120292
R14019 VGND VGND.n3504 0.120292
R14020 VGND.n3509 VGND.n3508 0.120292
R14021 VGND.n3567 VGND.n3566 0.120292
R14022 VGND.n3566 VGND.n3565 0.120292
R14023 VGND.n3562 VGND.n3561 0.120292
R14024 VGND.n3561 VGND.n3559 0.120292
R14025 VGND.n3559 VGND 0.120292
R14026 VGND.n3556 VGND.n3555 0.120292
R14027 VGND.n3555 VGND.n3554 0.120292
R14028 VGND.n3554 VGND.n3551 0.120292
R14029 VGND.n3548 VGND.n3547 0.120292
R14030 VGND.n3547 VGND.n3545 0.120292
R14031 VGND.n3545 VGND 0.120292
R14032 VGND.n3541 VGND.n3540 0.120292
R14033 VGND.n3540 VGND.n3539 0.120292
R14034 VGND.n3539 VGND.n3536 0.120292
R14035 VGND.n3532 VGND.n3531 0.120292
R14036 VGND.n3531 VGND.n3530 0.120292
R14037 VGND.n3527 VGND.n3526 0.120292
R14038 VGND.n1070 VGND.n1068 0.120292
R14039 VGND.n1079 VGND.n1077 0.120292
R14040 VGND.n1080 VGND.n1079 0.120292
R14041 VGND.n1085 VGND.n1083 0.120292
R14042 VGND.n1086 VGND.n1085 0.120292
R14043 VGND.n1090 VGND.n1086 0.120292
R14044 VGND.n3196 VGND.n3195 0.120292
R14045 VGND.n3195 VGND.n3193 0.120292
R14046 VGND.n3193 VGND.n3192 0.120292
R14047 VGND.n3186 VGND.n1098 0.120292
R14048 VGND.n3180 VGND.n3179 0.120292
R14049 VGND.n3179 VGND.n3177 0.120292
R14050 VGND.n3177 VGND.n3176 0.120292
R14051 VGND.n3172 VGND.n3171 0.120292
R14052 VGND.n3170 VGND.n3168 0.120292
R14053 VGND.n3168 VGND.n3166 0.120292
R14054 VGND.n3166 VGND.n3164 0.120292
R14055 VGND.n3164 VGND.n3162 0.120292
R14056 VGND.n3162 VGND.n3160 0.120292
R14057 VGND.n3160 VGND.n3158 0.120292
R14058 VGND.n3224 VGND.n3222 0.120292
R14059 VGND.n3231 VGND.n3228 0.120292
R14060 VGND.n3236 VGND.n3231 0.120292
R14061 VGND VGND.n3236 0.120292
R14062 VGND.n3252 VGND.n3251 0.120292
R14063 VGND.n3255 VGND.n3252 0.120292
R14064 VGND.n3256 VGND.n3255 0.120292
R14065 VGND.n3261 VGND.n3260 0.120292
R14066 VGND.n3264 VGND.n3261 0.120292
R14067 VGND.n3266 VGND.n3264 0.120292
R14068 VGND.n3271 VGND.n3270 0.120292
R14069 VGND.n3276 VGND.n3274 0.120292
R14070 VGND.n3278 VGND.n3276 0.120292
R14071 VGND.n3280 VGND.n3278 0.120292
R14072 VGND.n3283 VGND.n3280 0.120292
R14073 VGND.n3284 VGND.n3283 0.120292
R14074 VGND.n3285 VGND.n3284 0.120292
R14075 VGND.n3286 VGND.n3285 0.120292
R14076 VGND.n3292 VGND.n3290 0.120292
R14077 VGND.n3294 VGND.n3292 0.120292
R14078 VGND.n3295 VGND.n3294 0.120292
R14079 VGND.n3300 VGND.n3298 0.120292
R14080 VGND.n3303 VGND.n3300 0.120292
R14081 VGND.n3304 VGND.n3303 0.120292
R14082 VGND.n3311 VGND.n3310 0.120292
R14083 VGND.n3317 VGND.n3315 0.120292
R14084 VGND.n3448 VGND.n3446 0.120292
R14085 VGND.n3446 VGND.n3443 0.120292
R14086 VGND.n3440 VGND.n3439 0.120292
R14087 VGND.n3439 VGND.n3438 0.120292
R14088 VGND.n3438 VGND.n3436 0.120292
R14089 VGND.n3436 VGND.n3435 0.120292
R14090 VGND.n3432 VGND.n3431 0.120292
R14091 VGND.n3431 VGND.n3430 0.120292
R14092 VGND.n3430 VGND.n3427 0.120292
R14093 VGND.n3424 VGND.n3423 0.120292
R14094 VGND.n3423 VGND.n3421 0.120292
R14095 VGND.n3421 VGND.n3419 0.120292
R14096 VGND.n3419 VGND.n3416 0.120292
R14097 VGND.n3413 VGND.n3412 0.120292
R14098 VGND.n3412 VGND.n3411 0.120292
R14099 VGND.n3411 VGND.n3410 0.120292
R14100 VGND.n3403 VGND.n3402 0.120292
R14101 VGND.n3402 VGND.n3401 0.120292
R14102 VGND.n3401 VGND.n3398 0.120292
R14103 VGND.n3395 VGND.n3394 0.120292
R14104 VGND.n3394 VGND.n3392 0.120292
R14105 VGND.n3391 VGND.n3388 0.120292
R14106 VGND.n3388 VGND.n3387 0.120292
R14107 VGND.n3387 VGND.n3384 0.120292
R14108 VGND.n3380 VGND.n3379 0.120292
R14109 VGND.n3379 VGND.n3377 0.120292
R14110 VGND.n3377 VGND.n3375 0.120292
R14111 VGND.n3375 VGND.n3373 0.120292
R14112 VGND.n3373 VGND.n3370 0.120292
R14113 VGND.n3367 VGND.n3366 0.120292
R14114 VGND.n3366 VGND.n3364 0.120292
R14115 VGND.n3364 VGND.n3362 0.120292
R14116 VGND.n1165 VGND.n1147 0.120292
R14117 VGND.n1166 VGND.n1165 0.120292
R14118 VGND.n1170 VGND.n1145 0.120292
R14119 VGND.n1171 VGND.n1170 0.120292
R14120 VGND.n1172 VGND.n1171 0.120292
R14121 VGND.n1172 VGND.n1143 0.120292
R14122 VGND.n1176 VGND.n1143 0.120292
R14123 VGND.n1177 VGND.n1176 0.120292
R14124 VGND.n1178 VGND.n1141 0.120292
R14125 VGND.n1183 VGND.n1141 0.120292
R14126 VGND.n1184 VGND.n1183 0.120292
R14127 VGND.n1238 VGND.n1237 0.120292
R14128 VGND.n1237 VGND.n1236 0.120292
R14129 VGND.n1236 VGND.n1187 0.120292
R14130 VGND.n1228 VGND.n1227 0.120292
R14131 VGND.n1227 VGND.n1191 0.120292
R14132 VGND.n1223 VGND.n1191 0.120292
R14133 VGND.n1223 VGND.n1222 0.120292
R14134 VGND.n1219 VGND.n1218 0.120292
R14135 VGND.n1218 VGND.n1198 0.120292
R14136 VGND.n1214 VGND.n1198 0.120292
R14137 VGND.n1214 VGND.n1213 0.120292
R14138 VGND.n1213 VGND.n1212 0.120292
R14139 VGND.n1212 VGND.n1200 0.120292
R14140 VGND.n1208 VGND.n1200 0.120292
R14141 VGND.n1207 VGND.n1205 0.120292
R14142 VGND.n1205 VGND.n1203 0.120292
R14143 VGND.n3056 VGND.n3055 0.120292
R14144 VGND.n3055 VGND.n3053 0.120292
R14145 VGND.n3053 VGND.n3051 0.120292
R14146 VGND.n3051 VGND.n3049 0.120292
R14147 VGND.n3046 VGND.n3045 0.120292
R14148 VGND.n3045 VGND.n3044 0.120292
R14149 VGND.n3044 VGND.n3041 0.120292
R14150 VGND.n3038 VGND.n3037 0.120292
R14151 VGND.n3037 VGND.n3036 0.120292
R14152 VGND.n3036 VGND.n3034 0.120292
R14153 VGND.n3034 VGND.n3032 0.120292
R14154 VGND.n3032 VGND.n3030 0.120292
R14155 VGND.n3030 VGND.n3028 0.120292
R14156 VGND.n3028 VGND.n3027 0.120292
R14157 VGND.n3027 VGND.n3025 0.120292
R14158 VGND.n3025 VGND.n3024 0.120292
R14159 VGND.n3021 VGND.n3020 0.120292
R14160 VGND.n3020 VGND.n3019 0.120292
R14161 VGND.n3019 VGND.n3016 0.120292
R14162 VGND.n3012 VGND.n3011 0.120292
R14163 VGND.n3011 VGND.n3010 0.120292
R14164 VGND.n3010 VGND.n3007 0.120292
R14165 VGND.n3003 VGND.n3001 0.120292
R14166 VGND.n3001 VGND.n2999 0.120292
R14167 VGND.n2999 VGND.n2998 0.120292
R14168 VGND.n2995 VGND.n2994 0.120292
R14169 VGND.n2994 VGND.n2993 0.120292
R14170 VGND.n2990 VGND.n2989 0.120292
R14171 VGND.n2989 VGND.n2988 0.120292
R14172 VGND.n2988 VGND 0.120292
R14173 VGND.n2983 VGND.n2982 0.120292
R14174 VGND.n2982 VGND.n2980 0.120292
R14175 VGND.n2980 VGND.n2979 0.120292
R14176 VGND.n2976 VGND.n2975 0.120292
R14177 VGND.n2975 VGND.n2974 0.120292
R14178 VGND.n2971 VGND.n2970 0.120292
R14179 VGND.n2970 VGND.n2968 0.120292
R14180 VGND.n2856 VGND.n2855 0.120292
R14181 VGND.n2857 VGND.n2856 0.120292
R14182 VGND.n2859 VGND.n2857 0.120292
R14183 VGND.n2861 VGND.n2859 0.120292
R14184 VGND.n2866 VGND.n2861 0.120292
R14185 VGND.n2868 VGND.n2866 0.120292
R14186 VGND.n2874 VGND.n2872 0.120292
R14187 VGND.n2876 VGND.n2874 0.120292
R14188 VGND.n2877 VGND.n1274 0.120292
R14189 VGND.n2882 VGND.n1274 0.120292
R14190 VGND.n2883 VGND.n2882 0.120292
R14191 VGND.n2888 VGND.n1272 0.120292
R14192 VGND.n2938 VGND.n2937 0.120292
R14193 VGND.n2936 VGND.n2898 0.120292
R14194 VGND.n2932 VGND.n2898 0.120292
R14195 VGND.n2932 VGND.n2931 0.120292
R14196 VGND.n2927 VGND.n2926 0.120292
R14197 VGND.n2926 VGND.n2901 0.120292
R14198 VGND.n2922 VGND.n2901 0.120292
R14199 VGND.n2922 VGND.n2921 0.120292
R14200 VGND.n2921 VGND.n2920 0.120292
R14201 VGND.n2920 VGND.n2903 0.120292
R14202 VGND.n2915 VGND.n2903 0.120292
R14203 VGND.n2914 VGND.n2913 0.120292
R14204 VGND.n2913 VGND.n2912 0.120292
R14205 VGND.n2912 VGND.n2911 0.120292
R14206 VGND.n1370 VGND.n1365 0.120292
R14207 VGND.n1375 VGND.n1363 0.120292
R14208 VGND.n1383 VGND.n1360 0.120292
R14209 VGND.n1384 VGND.n1383 0.120292
R14210 VGND.n1388 VGND.n1358 0.120292
R14211 VGND.n1389 VGND.n1388 0.120292
R14212 VGND.n1390 VGND.n1389 0.120292
R14213 VGND.n1390 VGND.n1356 0.120292
R14214 VGND.n1394 VGND.n1356 0.120292
R14215 VGND.n1395 VGND.n1394 0.120292
R14216 VGND.n1396 VGND.n1354 0.120292
R14217 VGND.n1401 VGND.n1354 0.120292
R14218 VGND.n1402 VGND.n1401 0.120292
R14219 VGND.n1407 VGND.n1350 0.120292
R14220 VGND.n1409 VGND.n1408 0.120292
R14221 VGND.n1409 VGND.n1348 0.120292
R14222 VGND.n1414 VGND.n1348 0.120292
R14223 VGND.n1421 VGND.n1419 0.120292
R14224 VGND.n1423 VGND.n1421 0.120292
R14225 VGND.n1425 VGND.n1423 0.120292
R14226 VGND.n1427 VGND.n1425 0.120292
R14227 VGND.n1429 VGND.n1427 0.120292
R14228 VGND.n1431 VGND.n1429 0.120292
R14229 VGND.n1433 VGND.n1431 0.120292
R14230 VGND.n1434 VGND.n1433 0.120292
R14231 VGND.n1435 VGND.n1434 0.120292
R14232 VGND.n1441 VGND.n1439 0.120292
R14233 VGND.n1443 VGND.n1441 0.120292
R14234 VGND.n1445 VGND.n1443 0.120292
R14235 VGND.n1448 VGND.n1445 0.120292
R14236 VGND.n2626 VGND.n2579 0.120292
R14237 VGND.n2620 VGND.n2619 0.120292
R14238 VGND.n2619 VGND.n2617 0.120292
R14239 VGND.n2617 VGND.n2614 0.120292
R14240 VGND.n2614 VGND.n2613 0.120292
R14241 VGND.n2613 VGND.n2612 0.120292
R14242 VGND.n2607 VGND.n2606 0.120292
R14243 VGND.n2597 VGND.n2596 0.120292
R14244 VGND.n2656 VGND.n2654 0.120292
R14245 VGND.n2657 VGND.n2656 0.120292
R14246 VGND.n2662 VGND.n2660 0.120292
R14247 VGND.n2663 VGND.n2662 0.120292
R14248 VGND.n2664 VGND.n2663 0.120292
R14249 VGND.n2670 VGND.n2668 0.120292
R14250 VGND.n2672 VGND.n2670 0.120292
R14251 VGND.n2674 VGND.n2672 0.120292
R14252 VGND.n2676 VGND.n2674 0.120292
R14253 VGND.n2678 VGND.n2676 0.120292
R14254 VGND.n2680 VGND.n2678 0.120292
R14255 VGND.n2682 VGND.n2680 0.120292
R14256 VGND.n2684 VGND.n2682 0.120292
R14257 VGND.n2686 VGND.n2684 0.120292
R14258 VGND.n2688 VGND.n2686 0.120292
R14259 VGND.n2690 VGND.n2688 0.120292
R14260 VGND.n2692 VGND.n2690 0.120292
R14261 VGND.n2694 VGND.n2692 0.120292
R14262 VGND.n2697 VGND.n2694 0.120292
R14263 VGND.n2817 VGND.n2816 0.120292
R14264 VGND.n2816 VGND.n2814 0.120292
R14265 VGND.n2814 VGND.n2812 0.120292
R14266 VGND.n2812 VGND.n2810 0.120292
R14267 VGND.n2810 VGND.n2809 0.120292
R14268 VGND.n2809 VGND.n2807 0.120292
R14269 VGND.n2804 VGND.n1329 0.120292
R14270 VGND.n1333 VGND.n1329 0.120292
R14271 VGND.n2794 VGND.n2793 0.120292
R14272 VGND.n2793 VGND.n2792 0.120292
R14273 VGND.n2792 VGND.n2789 0.120292
R14274 VGND.n2780 VGND.n2779 0.120292
R14275 VGND.n2779 VGND.n2777 0.120292
R14276 VGND.n2777 VGND.n2775 0.120292
R14277 VGND.n2774 VGND.n2771 0.120292
R14278 VGND.n2771 VGND.n2770 0.120292
R14279 VGND.n2770 VGND.n2768 0.120292
R14280 VGND.n2768 VGND.n2766 0.120292
R14281 VGND.n2766 VGND.n2763 0.120292
R14282 VGND.n2763 VGND.n2758 0.120292
R14283 VGND.n2758 VGND.n2755 0.120292
R14284 VGND.n2752 VGND.n2751 0.120292
R14285 VGND.n2751 VGND.n2749 0.120292
R14286 VGND.n2749 VGND.n2747 0.120292
R14287 VGND.n2143 VGND.n2129 0.120292
R14288 VGND.n2151 VGND.n2149 0.120292
R14289 VGND.n2158 VGND.n2156 0.120292
R14290 VGND.n2160 VGND.n2158 0.120292
R14291 VGND.n2161 VGND.n2160 0.120292
R14292 VGND.n2162 VGND.n2161 0.120292
R14293 VGND.n2168 VGND.n2162 0.120292
R14294 VGND.n2215 VGND.n2214 0.120292
R14295 VGND.n2211 VGND.n2210 0.120292
R14296 VGND.n2210 VGND.n2209 0.120292
R14297 VGND.n2203 VGND.n2201 0.120292
R14298 VGND.n2198 VGND.n2196 0.120292
R14299 VGND.n2196 VGND.n2195 0.120292
R14300 VGND.n2192 VGND.n2191 0.120292
R14301 VGND.n2191 VGND.n2190 0.120292
R14302 VGND.n2184 VGND.n2181 0.120292
R14303 VGND.n2181 VGND.n2180 0.120292
R14304 VGND.n2278 VGND.n2275 0.120292
R14305 VGND.n2279 VGND.n2278 0.120292
R14306 VGND.n2286 VGND.n2285 0.120292
R14307 VGND.n2287 VGND.n2286 0.120292
R14308 VGND.n2293 VGND.n2292 0.120292
R14309 VGND.n2295 VGND.n2293 0.120292
R14310 VGND.n2302 VGND.n2301 0.120292
R14311 VGND.n2305 VGND.n2302 0.120292
R14312 VGND.n2306 VGND.n2305 0.120292
R14313 VGND.n2312 VGND.n2311 0.120292
R14314 VGND.n2321 VGND.n2320 0.120292
R14315 VGND.n2324 VGND.n2321 0.120292
R14316 VGND.n2326 VGND.n2324 0.120292
R14317 VGND.n2330 VGND.n2328 0.120292
R14318 VGND.n2331 VGND.n2330 0.120292
R14319 VGND.n2332 VGND.n2331 0.120292
R14320 VGND.n2338 VGND.n2336 0.120292
R14321 VGND.n2340 VGND.n2338 0.120292
R14322 VGND.n2347 VGND.n2345 0.120292
R14323 VGND.n2348 VGND.n2347 0.120292
R14324 VGND.n2349 VGND.n2348 0.120292
R14325 VGND.n2354 VGND.n2353 0.120292
R14326 VGND.n2359 VGND.n2357 0.120292
R14327 VGND.n2362 VGND.n2359 0.120292
R14328 VGND.n2507 VGND.n2505 0.120292
R14329 VGND.n2505 VGND.n2503 0.120292
R14330 VGND.n2500 VGND.n2499 0.120292
R14331 VGND.n2499 VGND.n2497 0.120292
R14332 VGND.n2497 VGND.n2496 0.120292
R14333 VGND.n2496 VGND.n2495 0.120292
R14334 VGND.n2490 VGND.n2489 0.120292
R14335 VGND.n2489 VGND.n2488 0.120292
R14336 VGND.n2488 VGND.n2487 0.120292
R14337 VGND.n2487 VGND.n2485 0.120292
R14338 VGND.n2481 VGND.n2480 0.120292
R14339 VGND.n2480 VGND.n2479 0.120292
R14340 VGND.n2476 VGND.n2475 0.120292
R14341 VGND.n2475 VGND.n2474 0.120292
R14342 VGND.n2474 VGND.n2471 0.120292
R14343 VGND.n2467 VGND.n2466 0.120292
R14344 VGND.n2466 VGND.n2465 0.120292
R14345 VGND.n2465 VGND.n2462 0.120292
R14346 VGND.n2459 VGND.n2458 0.120292
R14347 VGND.n2458 VGND.n2456 0.120292
R14348 VGND.n2456 VGND 0.120292
R14349 VGND.n2452 VGND.n2451 0.120292
R14350 VGND.n2451 VGND.n2450 0.120292
R14351 VGND.n2450 VGND.n2448 0.120292
R14352 VGND.n2448 VGND.n2446 0.120292
R14353 VGND.n2440 VGND.n2417 0.120292
R14354 VGND.n2435 VGND.n2434 0.120292
R14355 VGND.n2434 VGND.n2433 0.120292
R14356 VGND.n2429 VGND.n2428 0.120292
R14357 VGND.n2428 VGND.n2427 0.120292
R14358 VGND.n1601 VGND.n1600 0.120292
R14359 VGND VGND.n1601 0.120292
R14360 VGND.n1611 VGND.n1609 0.120292
R14361 VGND.n1611 VGND.n1610 0.120292
R14362 VGND.n1621 VGND.n1619 0.120292
R14363 VGND.n1623 VGND.n1621 0.120292
R14364 VGND.n1624 VGND.n1623 0.120292
R14365 VGND.n1625 VGND.n1624 0.120292
R14366 VGND.n1626 VGND.n1625 0.120292
R14367 VGND.n1589 VGND.n1588 0.120292
R14368 VGND.n1588 VGND.n1587 0.120292
R14369 VGND.n1544 VGND.n1543 0.120292
R14370 VGND.n1545 VGND.n1544 0.120292
R14371 VGND.n1580 VGND.n1545 0.120292
R14372 VGND.n1574 VGND.n1573 0.120292
R14373 VGND.n1564 VGND.n1562 0.120292
R14374 VGND.n1562 VGND.n1560 0.120292
R14375 VGND.n1560 VGND.n1558 0.120292
R14376 VGND.n1558 VGND.n1556 0.120292
R14377 VGND.n1556 VGND.n1554 0.120292
R14378 VGND.n1554 VGND.n1552 0.120292
R14379 VGND.n2054 VGND.n2051 0.120292
R14380 VGND.n2051 VGND.n2050 0.120292
R14381 VGND.n2050 VGND.n2048 0.120292
R14382 VGND.n2036 VGND.n2035 0.120292
R14383 VGND.n2035 VGND.n2034 0.120292
R14384 VGND.n2031 VGND.n2030 0.120292
R14385 VGND.n2029 VGND.n2026 0.120292
R14386 VGND.n2026 VGND.n2025 0.120292
R14387 VGND.n2025 VGND.n2022 0.120292
R14388 VGND.n1760 VGND.n1758 0.120292
R14389 VGND.n1761 VGND.n1760 0.120292
R14390 VGND.n1762 VGND.n1761 0.120292
R14391 VGND.n1767 VGND.n1765 0.120292
R14392 VGND.n1769 VGND.n1767 0.120292
R14393 VGND.n1771 VGND.n1769 0.120292
R14394 VGND.n1773 VGND.n1771 0.120292
R14395 VGND.n1775 VGND.n1773 0.120292
R14396 VGND.n1777 VGND.n1775 0.120292
R14397 VGND.n1778 VGND.n1777 0.120292
R14398 VGND.n1790 VGND.n1788 0.120292
R14399 VGND.n1792 VGND.n1790 0.120292
R14400 VGND.n1794 VGND.n1792 0.120292
R14401 VGND.n1796 VGND.n1794 0.120292
R14402 VGND.n1798 VGND.n1796 0.120292
R14403 VGND.n1800 VGND.n1798 0.120292
R14404 VGND.n1802 VGND.n1800 0.120292
R14405 VGND.n1805 VGND.n1802 0.120292
R14406 VGND.n1741 VGND.n1739 0.120292
R14407 VGND.n1739 VGND.n1736 0.120292
R14408 VGND.n1733 VGND.n1732 0.120292
R14409 VGND.n1732 VGND.n1731 0.120292
R14410 VGND.n1731 VGND 0.120292
R14411 VGND.n1725 VGND.n1724 0.120292
R14412 VGND.n1724 VGND.n1723 0.120292
R14413 VGND.n1716 VGND.n1715 0.120292
R14414 VGND.n1715 VGND.n1713 0.120292
R14415 VGND.n1702 VGND.n1701 0.120292
R14416 VGND.n1701 VGND.n1700 0.120292
R14417 VGND.n1696 VGND.n1694 0.120292
R14418 VGND.n1694 VGND.n1692 0.120292
R14419 VGND.n1692 VGND.n1690 0.120292
R14420 VGND.n1690 VGND.n1688 0.120292
R14421 VGND.n1688 VGND.n1686 0.120292
R14422 VGND.n1686 VGND.n1684 0.120292
R14423 VGND.n1684 VGND.n1681 0.120292
R14424 VGND.n1681 VGND.n1676 0.120292
R14425 VGND.n1676 VGND.n1673 0.120292
R14426 VGND.n1669 VGND.n1666 0.120292
R14427 VGND.n141 VGND.n140 0.120292
R14428 VGND.n144 VGND.n141 0.120292
R14429 VGND.n149 VGND.n148 0.120292
R14430 VGND.n150 VGND.n149 0.120292
R14431 VGND VGND.n150 0.120292
R14432 VGND.n160 VGND.n159 0.120292
R14433 VGND.n165 VGND.n163 0.120292
R14434 VGND.n166 VGND.n165 0.120292
R14435 VGND.n167 VGND.n166 0.120292
R14436 VGND.n208 VGND.n207 0.120292
R14437 VGND.n199 VGND.n198 0.120292
R14438 VGND.n198 VGND.n196 0.120292
R14439 VGND.n196 VGND.n194 0.120292
R14440 VGND.n187 VGND.n186 0.120292
R14441 VGND.n186 VGND.n185 0.120292
R14442 VGND.n185 VGND.n183 0.120292
R14443 VGND.n183 VGND.n181 0.120292
R14444 VGND.n5132 VGND.n5131 0.120292
R14445 VGND.n5131 VGND.n5128 0.120292
R14446 VGND.n5125 VGND.n5124 0.120292
R14447 VGND.n5124 VGND.n5123 0.120292
R14448 VGND.n5123 VGND.n5121 0.120292
R14449 VGND.n5121 VGND.n5119 0.120292
R14450 VGND.n5119 VGND.n5118 0.120292
R14451 VGND.n5118 VGND.n5116 0.120292
R14452 VGND.n5113 VGND.n5112 0.120292
R14453 VGND.n5112 VGND.n5111 0.120292
R14454 VGND.n5111 VGND.n5108 0.120292
R14455 VGND.n5105 VGND.n5104 0.120292
R14456 VGND.n5104 VGND.n5102 0.120292
R14457 VGND.n5102 VGND.n5100 0.120292
R14458 VGND.n5100 VGND.n5098 0.120292
R14459 VGND.n5098 VGND.n5096 0.120292
R14460 VGND.n5096 VGND.n5095 0.120292
R14461 VGND.n5095 VGND.n5094 0.120292
R14462 VGND.n5087 VGND.n5085 0.120292
R14463 VGND.n5085 VGND.n5083 0.120292
R14464 VGND.n5080 VGND.n5079 0.120292
R14465 VGND.n5079 VGND.n5077 0.120292
R14466 VGND.n5076 VGND.n5074 0.120292
R14467 VGND.n5074 VGND.n5072 0.120292
R14468 VGND.n5072 VGND.n5071 0.120292
R14469 VGND.n5067 VGND.n5066 0.120292
R14470 VGND.n5066 VGND.n5064 0.120292
R14471 VGND.n5064 VGND.n5062 0.120292
R14472 VGND.n5062 VGND.n5060 0.120292
R14473 VGND.n5060 VGND.n5059 0.120292
R14474 VGND.n5056 VGND.n5055 0.120292
R14475 VGND.n5055 VGND.n5053 0.120292
R14476 VGND.n5053 VGND.n5051 0.120292
R14477 VGND.n5051 VGND.n5049 0.120292
R14478 VGND.n5049 VGND.n5046 0.120292
R14479 VGND.n5046 VGND.n5041 0.120292
R14480 VGND.n1977 VGND.n1975 0.120292
R14481 VGND.n1975 VGND.n1972 0.120292
R14482 VGND.n1969 VGND.n1968 0.120292
R14483 VGND.n1968 VGND.n1967 0.120292
R14484 VGND.n1967 VGND.n1964 0.120292
R14485 VGND.n1960 VGND.n1959 0.120292
R14486 VGND.n1958 VGND.n1953 0.120292
R14487 VGND.n1953 VGND.n1952 0.120292
R14488 VGND.n1952 VGND.n1951 0.120292
R14489 VGND.n1948 VGND.n1947 0.120292
R14490 VGND.n1947 VGND.n1946 0.120292
R14491 VGND.n1946 VGND.n1945 0.120292
R14492 VGND.n1940 VGND.n1937 0.120292
R14493 VGND.n1937 VGND.n1936 0.120292
R14494 VGND.n1936 VGND.n1934 0.120292
R14495 VGND.n1934 VGND.n1932 0.120292
R14496 VGND.n1932 VGND.n1930 0.120292
R14497 VGND.n1927 VGND.n1924 0.120292
R14498 VGND.n1924 VGND.n1923 0.120292
R14499 VGND.n1923 VGND.n1920 0.120292
R14500 VGND.n1917 VGND.n1916 0.120292
R14501 VGND.n1916 VGND.n1915 0.120292
R14502 VGND.n1915 VGND.n1913 0.120292
R14503 VGND.n1913 VGND.n1912 0.120292
R14504 VGND.n1912 VGND.n1910 0.120292
R14505 VGND.n1910 VGND.n1908 0.120292
R14506 VGND.n1904 VGND.n1903 0.120292
R14507 VGND.n1903 VGND.n1902 0.120292
R14508 VGND.n1899 VGND.n1898 0.120292
R14509 VGND.n1898 VGND.n1897 0.120292
R14510 VGND.n1897 VGND.n1896 0.120292
R14511 VGND.n1896 VGND.n1894 0.120292
R14512 VGND.n1891 VGND.n1890 0.120292
R14513 VGND.n4230 VGND.n4228 0.120292
R14514 VGND.n4231 VGND.n4230 0.120292
R14515 VGND.n4241 VGND.n4239 0.120292
R14516 VGND VGND.n4242 0.120292
R14517 VGND.n4247 VGND.n4245 0.120292
R14518 VGND.n4249 VGND.n4247 0.120292
R14519 VGND.n4250 VGND.n4249 0.120292
R14520 VGND.n4251 VGND.n4250 0.120292
R14521 VGND.n4253 VGND.n4251 0.120292
R14522 VGND.n4264 VGND.n4263 0.120292
R14523 VGND.n4265 VGND.n4264 0.120292
R14524 VGND VGND.n4265 0.120292
R14525 VGND.n4272 VGND.n4270 0.120292
R14526 VGND.n4273 VGND.n4272 0.120292
R14527 VGND.n4274 VGND.n4273 0.120292
R14528 VGND.n4275 VGND.n4274 0.120292
R14529 VGND.n4286 VGND.n4275 0.120292
R14530 VGND.n4294 VGND.n4292 0.120292
R14531 VGND.n4456 VGND.n4455 0.120292
R14532 VGND.n4455 VGND.n4453 0.120292
R14533 VGND.n4453 VGND.n4451 0.120292
R14534 VGND.n4451 VGND.n4449 0.120292
R14535 VGND.n4449 VGND.n4448 0.120292
R14536 VGND.n4444 VGND.n4443 0.120292
R14537 VGND.n4443 VGND.n4441 0.120292
R14538 VGND.n4441 VGND.n4439 0.120292
R14539 VGND.n4439 VGND.n4438 0.120292
R14540 VGND.n4438 VGND.n4437 0.120292
R14541 VGND.n4437 VGND.n4436 0.120292
R14542 VGND.n4431 VGND.n4429 0.120292
R14543 VGND.n4429 VGND.n4427 0.120292
R14544 VGND.n4427 VGND.n4425 0.120292
R14545 VGND.n4425 VGND.n4423 0.120292
R14546 VGND.n4423 VGND.n4422 0.120292
R14547 VGND.n4422 VGND.n4421 0.120292
R14548 VGND.n4403 VGND.n4401 0.120292
R14549 VGND.n4401 VGND.n4400 0.120292
R14550 VGND.n4396 VGND.n4395 0.120292
R14551 VGND.n4395 VGND.n4394 0.120292
R14552 VGND.n4394 VGND.n4392 0.120292
R14553 VGND.n4392 VGND.n4390 0.120292
R14554 VGND.n4390 VGND.n4389 0.120292
R14555 VGND.n4385 VGND.n4384 0.120292
R14556 VGND.n4384 VGND.n4382 0.120292
R14557 VGND.n4382 VGND.n4380 0.120292
R14558 VGND.n4380 VGND.n4378 0.120292
R14559 VGND.n4378 VGND.n4376 0.120292
R14560 VGND.n4376 VGND.n4374 0.120292
R14561 VGND.n4374 VGND.n4373 0.120292
R14562 VGND.n4890 VGND.n4888 0.120292
R14563 VGND.n4892 VGND.n4890 0.120292
R14564 VGND.n4894 VGND.n4892 0.120292
R14565 VGND.n4896 VGND.n4894 0.120292
R14566 VGND.n4898 VGND.n4896 0.120292
R14567 VGND.n4899 VGND.n4898 0.120292
R14568 VGND.n4905 VGND.n4904 0.120292
R14569 VGND.n4907 VGND.n4905 0.120292
R14570 VGND.n4913 VGND.n4911 0.120292
R14571 VGND.n4915 VGND.n4913 0.120292
R14572 VGND.n4962 VGND.n4961 0.120292
R14573 VGND.n4961 VGND 0.120292
R14574 VGND.n4960 VGND.n4957 0.120292
R14575 VGND.n4957 VGND.n4956 0.120292
R14576 VGND.n4956 VGND.n4954 0.120292
R14577 VGND.n4954 VGND.n4952 0.120292
R14578 VGND.n4952 VGND.n4949 0.120292
R14579 VGND.n4949 VGND.n4944 0.120292
R14580 VGND.n4944 VGND.n4941 0.120292
R14581 VGND.n4938 VGND.n4937 0.120292
R14582 VGND.n4937 VGND.n4936 0.120292
R14583 VGND.n4932 VGND.n4931 0.120292
R14584 VGND.n6 VGND.n4 0.120292
R14585 VGND.n8 VGND.n6 0.120292
R14586 VGND.n10 VGND.n8 0.120292
R14587 VGND.n11 VGND.n10 0.120292
R14588 VGND.n12 VGND.n11 0.120292
R14589 VGND.n17 VGND.n15 0.120292
R14590 VGND.n19 VGND.n17 0.120292
R14591 VGND VGND.n19 0.120292
R14592 VGND.n5593 VGND.n5592 0.120292
R14593 VGND.n5592 VGND.n5591 0.120292
R14594 VGND.n5591 VGND.n5588 0.120292
R14595 VGND.n5585 VGND.n5584 0.120292
R14596 VGND.n5584 VGND.n5582 0.120292
R14597 VGND.n5582 VGND 0.120292
R14598 VGND.n5579 VGND.n5578 0.120292
R14599 VGND.n5578 VGND.n5577 0.120292
R14600 VGND.n5203 VGND.n5202 0.120292
R14601 VGND.n5206 VGND.n5203 0.120292
R14602 VGND.n5207 VGND.n5206 0.120292
R14603 VGND.n5212 VGND.n5210 0.120292
R14604 VGND.n5213 VGND.n5212 0.120292
R14605 VGND VGND.n5213 0.120292
R14606 VGND.n5218 VGND.n5217 0.120292
R14607 VGND.n5220 VGND.n5218 0.120292
R14608 VGND.n5222 VGND.n5220 0.120292
R14609 VGND.n5224 VGND.n5222 0.120292
R14610 VGND.n5226 VGND.n5224 0.120292
R14611 VGND.n5230 VGND.n5226 0.120292
R14612 VGND.n5234 VGND.n5230 0.120292
R14613 VGND.n5236 VGND.n5234 0.120292
R14614 VGND.n5241 VGND.n5236 0.120292
R14615 VGND.n5244 VGND.n5241 0.120292
R14616 VGND.n5245 VGND.n5244 0.120292
R14617 VGND.n5250 VGND.n5248 0.120292
R14618 VGND.n5252 VGND.n5250 0.120292
R14619 VGND.n5254 VGND.n5252 0.120292
R14620 VGND.n5256 VGND.n5254 0.120292
R14621 VGND.n5259 VGND.n5256 0.120292
R14622 VGND.n5261 VGND.n5259 0.120292
R14623 VGND.n5321 VGND.n5319 0.120292
R14624 VGND.n5324 VGND.n5321 0.120292
R14625 VGND.n5329 VGND.n5324 0.120292
R14626 VGND.n5332 VGND.n5329 0.120292
R14627 VGND.n5333 VGND.n5332 0.120292
R14628 VGND.n5338 VGND.n5336 0.120292
R14629 VGND.n5340 VGND.n5338 0.120292
R14630 VGND.n5342 VGND.n5340 0.120292
R14631 VGND.n5344 VGND.n5342 0.120292
R14632 VGND.n5347 VGND.n5344 0.120292
R14633 VGND.n5348 VGND.n5347 0.120292
R14634 VGND.n5353 VGND.n5351 0.120292
R14635 VGND.n5355 VGND.n5353 0.120292
R14636 VGND.n5357 VGND.n5355 0.120292
R14637 VGND.n5358 VGND.n5357 0.120292
R14638 VGND.n5363 VGND.n5362 0.120292
R14639 VGND.n5365 VGND.n5363 0.120292
R14640 VGND.n5373 VGND.n5371 0.120292
R14641 VGND.n5375 VGND.n5373 0.120292
R14642 VGND.n5377 VGND.n5375 0.120292
R14643 VGND.n5380 VGND.n5377 0.120292
R14644 VGND.n5381 VGND.n5380 0.120292
R14645 VGND.n5382 VGND.n5381 0.120292
R14646 VGND.n5383 VGND.n5382 0.120292
R14647 VGND.n5388 VGND.n5386 0.120292
R14648 VGND.n5390 VGND.n5388 0.120292
R14649 VGND.n5392 VGND.n5390 0.120292
R14650 VGND.n5394 VGND.n5392 0.120292
R14651 VGND.n5396 VGND.n5394 0.120292
R14652 VGND.n5398 VGND.n5396 0.120292
R14653 VGND.n5401 VGND.n5398 0.120292
R14654 VGND.n5402 VGND.n5401 0.120292
R14655 VGND.n5403 VGND.n5402 0.120292
R14656 VGND.n5404 VGND.n5403 0.120292
R14657 VGND.n5409 VGND.n5407 0.120292
R14658 VGND.n5410 VGND.n5409 0.120292
R14659 VGND.n5415 VGND.n5413 0.120292
R14660 VGND.n5416 VGND.n5415 0.120292
R14661 VGND.n5420 VGND.n5416 0.120292
R14662 VGND.n5461 VGND.n5460 0.120292
R14663 VGND.n5466 VGND.n5464 0.120292
R14664 VGND.n5467 VGND.n5466 0.120292
R14665 VGND VGND.n5467 0.120292
R14666 VGND.n5472 VGND.n5471 0.120292
R14667 VGND.n5475 VGND.n5472 0.120292
R14668 VGND.n5476 VGND.n5475 0.120292
R14669 VGND.n5481 VGND.n5479 0.120292
R14670 VGND.n5483 VGND.n5481 0.120292
R14671 VGND.n5485 VGND.n5483 0.120292
R14672 VGND.n5487 VGND.n5485 0.120292
R14673 VGND.n5490 VGND.n5487 0.120292
R14674 VGND.n5491 VGND.n5490 0.120292
R14675 VGND.n5496 VGND.n5494 0.120292
R14676 VGND.n5498 VGND.n5496 0.120292
R14677 VGND.n5500 VGND.n5498 0.120292
R14678 VGND.n5502 VGND.n5500 0.120292
R14679 VGND.n5505 VGND.n5502 0.120292
R14680 VGND.n5506 VGND.n5505 0.120292
R14681 VGND.n5565 VGND.n5564 0.120292
R14682 VGND.n5564 VGND.n5563 0.120292
R14683 VGND.n5563 VGND.n5561 0.120292
R14684 VGND.n5561 VGND.n5559 0.120292
R14685 VGND.n5559 VGND.n5556 0.120292
R14686 VGND.n5556 VGND.n5551 0.120292
R14687 VGND.n5551 VGND.n5548 0.120292
R14688 VGND.n5545 VGND.n5544 0.120292
R14689 VGND.n5544 VGND.n5542 0.120292
R14690 VGND.n5542 VGND.n5541 0.120292
R14691 VGND.n5541 VGND.n5539 0.120292
R14692 VGND.n5539 VGND.n5537 0.120292
R14693 VGND.n5537 VGND.n5534 0.120292
R14694 VGND.n5531 VGND.n5530 0.120292
R14695 VGND.n5530 VGND.n5528 0.120292
R14696 VGND.n5528 VGND.n5527 0.120292
R14697 VGND.n5527 VGND.n5525 0.120292
R14698 VGND.n5525 VGND.n5523 0.120292
R14699 VGND.n5520 VGND.n5519 0.120292
R14700 VGND.n5519 VGND.n5518 0.120292
R14701 VGND.n4405 VGND 0.118727
R14702 VGND.n3856 VGND.n3855 0.107365
R14703 VGND.n3319 VGND.n3318 0.107365
R14704 VGND.n317 VGND 0.104136
R14705 VGND.n406 VGND 0.104136
R14706 VGND.n674 VGND 0.104136
R14707 VGND.n840 VGND 0.104136
R14708 VGND.n1057 VGND 0.104136
R14709 VGND.n1152 VGND 0.104136
R14710 VGND.n1366 VGND 0.104136
R14711 VGND.n2134 VGND 0.104136
R14712 VGND.n1595 VGND 0.104136
R14713 VGND.n138 VGND 0.104136
R14714 VGND.n4224 VGND 0.104136
R14715 VGND.n4712 VGND.n4710 0.102062
R14716 VGND.n964 VGND.n962 0.102062
R14717 VGND.n2968 VGND.n2965 0.102062
R14718 VGND.n2699 VGND.n2697 0.102062
R14719 VGND.n2364 VGND.n2362 0.102062
R14720 VGND.n1807 VGND.n1805 0.102062
R14721 VGND.n5041 VGND.n5035 0.102062
R14722 VGND.n4026 VGND 0.10076
R14723 VGND.n4064 VGND 0.10076
R14724 VGND.n733 VGND 0.10076
R14725 VGND.n2877 VGND 0.10076
R14726 VGND VGND 0.10076
R14727 VGND.n3235 VGND.n3232 0.1005
R14728 VGND.n349 VGND 0.0994583
R14729 VGND.n364 VGND 0.0994583
R14730 VGND.n4829 VGND 0.0994583
R14731 VGND.n4114 VGND 0.0994583
R14732 VGND.n694 VGND 0.0994583
R14733 VGND.n3756 VGND 0.0994583
R14734 VGND VGND.n3728 0.0994583
R14735 VGND.n3839 VGND 0.0994583
R14736 VGND.n3937 VGND 0.0994583
R14737 VGND.n3911 VGND 0.0994583
R14738 VGND.n760 VGND 0.0994583
R14739 VGND.n3489 VGND 0.0994583
R14740 VGND.n3493 VGND 0.0994583
R14741 VGND.n1068 VGND 0.0994583
R14742 VGND.n3240 VGND 0.0994583
R14743 VGND.n3251 VGND 0.0994583
R14744 VGND.n1027 VGND 0.0994583
R14745 VGND VGND.n1207 0.0994583
R14746 VGND.n3046 VGND 0.0994583
R14747 VGND VGND.n2597 0.0994583
R14748 VGND VGND.n2203 0.0994583
R14749 VGND.n2311 VGND 0.0994583
R14750 VGND.n2333 VGND 0.0994583
R14751 VGND.n2345 VGND 0.0994583
R14752 VGND.n2357 VGND 0.0994583
R14753 VGND VGND.n2494 0.0994583
R14754 VGND VGND.n2029 0.0994583
R14755 VGND.n1782 VGND 0.0994583
R14756 VGND VGND.n5093 0.0994583
R14757 VGND VGND.n1941 0.0994583
R14758 VGND.n321 VGND 0.0981562
R14759 VGND VGND 0.0981562
R14760 VGND.n326 VGND 0.0981562
R14761 VGND.n339 VGND 0.0981562
R14762 VGND.n4586 VGND 0.0981562
R14763 VGND.n356 VGND 0.0981562
R14764 VGND.n359 VGND 0.0981562
R14765 VGND.n4565 VGND 0.0981562
R14766 VGND.n362 VGND 0.0981562
R14767 VGND VGND.n4550 0.0981562
R14768 VGND.n4619 VGND 0.0981562
R14769 VGND.n4660 VGND 0.0981562
R14770 VGND.n4670 VGND 0.0981562
R14771 VGND.n4671 VGND 0.0981562
R14772 VGND VGND 0.0981562
R14773 VGND.n4675 VGND 0.0981562
R14774 VGND.n4683 VGND 0.0981562
R14775 VGND.n4705 VGND 0.0981562
R14776 VGND.n4848 VGND 0.0981562
R14777 VGND.n4842 VGND 0.0981562
R14778 VGND.n4834 VGND 0.0981562
R14779 VGND VGND.n4821 0.0981562
R14780 VGND.n4803 VGND 0.0981562
R14781 VGND.n4794 VGND 0.0981562
R14782 VGND.n4781 VGND 0.0981562
R14783 VGND VGND.n4780 0.0981562
R14784 VGND VGND.n4777 0.0981562
R14785 VGND.n4775 VGND 0.0981562
R14786 VGND VGND.n4774 0.0981562
R14787 VGND.n4766 VGND 0.0981562
R14788 VGND VGND.n4765 0.0981562
R14789 VGND VGND.n4764 0.0981562
R14790 VGND.n412 VGND 0.0981562
R14791 VGND VGND.n403 0.0981562
R14792 VGND.n419 VGND 0.0981562
R14793 VGND.n482 VGND 0.0981562
R14794 VGND.n474 VGND 0.0981562
R14795 VGND VGND.n473 0.0981562
R14796 VGND.n465 VGND 0.0981562
R14797 VGND VGND.n463 0.0981562
R14798 VGND.n455 VGND 0.0981562
R14799 VGND VGND.n451 0.0981562
R14800 VGND.n4136 VGND 0.0981562
R14801 VGND VGND.n4135 0.0981562
R14802 VGND.n4130 VGND 0.0981562
R14803 VGND VGND 0.0981562
R14804 VGND VGND.n4106 0.0981562
R14805 VGND.n4098 VGND 0.0981562
R14806 VGND VGND.n4096 0.0981562
R14807 VGND.n529 VGND 0.0981562
R14808 VGND.n537 VGND 0.0981562
R14809 VGND VGND 0.0981562
R14810 VGND.n540 VGND 0.0981562
R14811 VGND.n549 VGND 0.0981562
R14812 VGND VGND 0.0981562
R14813 VGND.n552 VGND 0.0981562
R14814 VGND.n562 VGND 0.0981562
R14815 VGND.n4014 VGND 0.0981562
R14816 VGND.n4018 VGND 0.0981562
R14817 VGND.n4021 VGND 0.0981562
R14818 VGND.n4023 VGND 0.0981562
R14819 VGND.n4031 VGND 0.0981562
R14820 VGND.n4033 VGND 0.0981562
R14821 VGND.n4089 VGND 0.0981562
R14822 VGND VGND.n4081 0.0981562
R14823 VGND VGND.n4080 0.0981562
R14824 VGND.n4069 VGND 0.0981562
R14825 VGND VGND 0.0981562
R14826 VGND VGND.n4057 0.0981562
R14827 VGND VGND.n4056 0.0981562
R14828 VGND.n680 VGND 0.0981562
R14829 VGND.n683 VGND 0.0981562
R14830 VGND VGND.n670 0.0981562
R14831 VGND VGND.n668 0.0981562
R14832 VGND.n704 VGND 0.0981562
R14833 VGND.n712 VGND 0.0981562
R14834 VGND.n713 VGND 0.0981562
R14835 VGND.n718 VGND 0.0981562
R14836 VGND.n720 VGND 0.0981562
R14837 VGND.n727 VGND 0.0981562
R14838 VGND.n728 VGND 0.0981562
R14839 VGND.n3772 VGND 0.0981562
R14840 VGND.n3748 VGND 0.0981562
R14841 VGND.n3742 VGND 0.0981562
R14842 VGND.n3802 VGND 0.0981562
R14843 VGND.n3806 VGND 0.0981562
R14844 VGND.n3819 VGND 0.0981562
R14845 VGND.n3854 VGND 0.0981562
R14846 VGND.n3954 VGND 0.0981562
R14847 VGND.n3946 VGND 0.0981562
R14848 VGND VGND.n3936 0.0981562
R14849 VGND VGND.n3934 0.0981562
R14850 VGND VGND.n3929 0.0981562
R14851 VGND VGND.n3926 0.0981562
R14852 VGND VGND 0.0981562
R14853 VGND VGND.n3904 0.0981562
R14854 VGND.n3900 VGND 0.0981562
R14855 VGND.n844 VGND 0.0981562
R14856 VGND VGND.n837 0.0981562
R14857 VGND.n858 VGND 0.0981562
R14858 VGND.n864 VGND 0.0981562
R14859 VGND.n870 VGND 0.0981562
R14860 VGND VGND.n825 0.0981562
R14861 VGND.n815 VGND 0.0981562
R14862 VGND VGND.n812 0.0981562
R14863 VGND VGND.n806 0.0981562
R14864 VGND.n788 VGND 0.0981562
R14865 VGND.n3617 VGND 0.0981562
R14866 VGND.n3597 VGND 0.0981562
R14867 VGND.n3593 VGND 0.0981562
R14868 VGND VGND.n3592 0.0981562
R14869 VGND VGND.n3590 0.0981562
R14870 VGND VGND.n3589 0.0981562
R14871 VGND.n767 VGND 0.0981562
R14872 VGND.n921 VGND 0.0981562
R14873 VGND.n927 VGND 0.0981562
R14874 VGND.n940 VGND 0.0981562
R14875 VGND.n947 VGND 0.0981562
R14876 VGND.n957 VGND 0.0981562
R14877 VGND.n3476 VGND 0.0981562
R14878 VGND.n3498 VGND 0.0981562
R14879 VGND.n3503 VGND 0.0981562
R14880 VGND.n3507 VGND 0.0981562
R14881 VGND.n3571 VGND 0.0981562
R14882 VGND.n3567 VGND 0.0981562
R14883 VGND.n3562 VGND 0.0981562
R14884 VGND.n3556 VGND 0.0981562
R14885 VGND.n3548 VGND 0.0981562
R14886 VGND.n3541 VGND 0.0981562
R14887 VGND.n3533 VGND 0.0981562
R14888 VGND.n3527 VGND 0.0981562
R14889 VGND.n1064 VGND 0.0981562
R14890 VGND VGND 0.0981562
R14891 VGND.n1065 VGND 0.0981562
R14892 VGND.n1074 VGND 0.0981562
R14893 VGND VGND.n1053 0.0981562
R14894 VGND.n1077 VGND 0.0981562
R14895 VGND.n1092 VGND 0.0981562
R14896 VGND.n1095 VGND 0.0981562
R14897 VGND.n1096 VGND 0.0981562
R14898 VGND.n1098 VGND 0.0981562
R14899 VGND.n1101 VGND 0.0981562
R14900 VGND.n3180 VGND 0.0981562
R14901 VGND.n1104 VGND 0.0981562
R14902 VGND.n3228 VGND 0.0981562
R14903 VGND.n3237 VGND 0.0981562
R14904 VGND.n3245 VGND 0.0981562
R14905 VGND.n3247 VGND 0.0981562
R14906 VGND.n3260 VGND 0.0981562
R14907 VGND.n3267 VGND 0.0981562
R14908 VGND.n3287 VGND 0.0981562
R14909 VGND.n3298 VGND 0.0981562
R14910 VGND.n3309 VGND 0.0981562
R14911 VGND.n3310 VGND 0.0981562
R14912 VGND.n3312 VGND 0.0981562
R14913 VGND.n3440 VGND 0.0981562
R14914 VGND.n3424 VGND 0.0981562
R14915 VGND.n3413 VGND 0.0981562
R14916 VGND VGND.n3404 0.0981562
R14917 VGND.n3395 VGND 0.0981562
R14918 VGND.n3381 VGND 0.0981562
R14919 VGND VGND.n3380 0.0981562
R14920 VGND VGND 0.0981562
R14921 VGND VGND.n3367 0.0981562
R14922 VGND VGND 0.0981562
R14923 VGND VGND.n1147 0.0981562
R14924 VGND VGND.n1145 0.0981562
R14925 VGND.n1178 VGND 0.0981562
R14926 VGND.n1185 VGND 0.0981562
R14927 VGND.n1188 VGND 0.0981562
R14928 VGND.n1229 VGND 0.0981562
R14929 VGND VGND.n1220 0.0981562
R14930 VGND VGND.n1219 0.0981562
R14931 VGND.n3057 VGND 0.0981562
R14932 VGND VGND.n3056 0.0981562
R14933 VGND.n3038 VGND 0.0981562
R14934 VGND.n3021 VGND 0.0981562
R14935 VGND.n3013 VGND 0.0981562
R14936 VGND.n3004 VGND 0.0981562
R14937 VGND VGND.n2995 0.0981562
R14938 VGND.n2990 VGND 0.0981562
R14939 VGND.n2983 VGND 0.0981562
R14940 VGND.n2976 VGND 0.0981562
R14941 VGND.n2971 VGND 0.0981562
R14942 VGND.n2869 VGND 0.0981562
R14943 VGND.n2872 VGND 0.0981562
R14944 VGND.n2884 VGND 0.0981562
R14945 VGND VGND.n1272 0.0981562
R14946 VGND.n2893 VGND 0.0981562
R14947 VGND VGND.n2942 0.0981562
R14948 VGND.n2939 VGND 0.0981562
R14949 VGND VGND.n2938 0.0981562
R14950 VGND VGND.n2936 0.0981562
R14951 VGND.n2928 VGND 0.0981562
R14952 VGND VGND 0.0981562
R14953 VGND VGND.n2914 0.0981562
R14954 VGND VGND.n1363 0.0981562
R14955 VGND.n1378 VGND 0.0981562
R14956 VGND VGND.n1360 0.0981562
R14957 VGND VGND.n1358 0.0981562
R14958 VGND.n1396 VGND 0.0981562
R14959 VGND.n1403 VGND 0.0981562
R14960 VGND.n1416 VGND 0.0981562
R14961 VGND.n1419 VGND 0.0981562
R14962 VGND.n1436 VGND 0.0981562
R14963 VGND.n1439 VGND 0.0981562
R14964 VGND VGND.n2626 0.0981562
R14965 VGND VGND.n2620 0.0981562
R14966 VGND.n2609 VGND 0.0981562
R14967 VGND VGND.n2608 0.0981562
R14968 VGND VGND.n2604 0.0981562
R14969 VGND VGND.n2598 0.0981562
R14970 VGND.n2649 VGND 0.0981562
R14971 VGND.n2651 VGND 0.0981562
R14972 VGND.n2654 VGND 0.0981562
R14973 VGND.n2660 VGND 0.0981562
R14974 VGND.n2665 VGND 0.0981562
R14975 VGND.n2668 VGND 0.0981562
R14976 VGND VGND.n2821 0.0981562
R14977 VGND VGND.n2818 0.0981562
R14978 VGND VGND.n2804 0.0981562
R14979 VGND.n2795 VGND 0.0981562
R14980 VGND VGND.n2794 0.0981562
R14981 VGND.n2736 VGND 0.0981562
R14982 VGND VGND.n2783 0.0981562
R14983 VGND VGND.n2780 0.0981562
R14984 VGND VGND.n2774 0.0981562
R14985 VGND VGND 0.0981562
R14986 VGND VGND.n2752 0.0981562
R14987 VGND VGND 0.0981562
R14988 VGND VGND.n2129 0.0981562
R14989 VGND VGND.n2127 0.0981562
R14990 VGND VGND.n2126 0.0981562
R14991 VGND.n2149 VGND 0.0981562
R14992 VGND.n2153 VGND 0.0981562
R14993 VGND.n2222 VGND 0.0981562
R14994 VGND.n2216 VGND 0.0981562
R14995 VGND.n2211 VGND 0.0981562
R14996 VGND.n2205 VGND 0.0981562
R14997 VGND VGND.n2199 0.0981562
R14998 VGND VGND.n2198 0.0981562
R14999 VGND.n2192 VGND 0.0981562
R15000 VGND.n2186 VGND 0.0981562
R15001 VGND VGND.n2185 0.0981562
R15002 VGND VGND.n2184 0.0981562
R15003 VGND.n2280 VGND 0.0981562
R15004 VGND.n2285 VGND 0.0981562
R15005 VGND.n2288 VGND 0.0981562
R15006 VGND.n2292 VGND 0.0981562
R15007 VGND.n2297 VGND 0.0981562
R15008 VGND.n2301 VGND 0.0981562
R15009 VGND.n2307 VGND 0.0981562
R15010 VGND VGND.n1487 0.0981562
R15011 VGND.n2328 VGND 0.0981562
R15012 VGND.n2342 VGND 0.0981562
R15013 VGND.n2350 VGND 0.0981562
R15014 VGND.n2353 VGND 0.0981562
R15015 VGND VGND.n2500 0.0981562
R15016 VGND.n2481 VGND 0.0981562
R15017 VGND VGND 0.0981562
R15018 VGND.n2476 VGND 0.0981562
R15019 VGND.n2468 VGND 0.0981562
R15020 VGND.n2459 VGND 0.0981562
R15021 VGND.n2453 VGND 0.0981562
R15022 VGND.n2442 VGND 0.0981562
R15023 VGND VGND.n2441 0.0981562
R15024 VGND VGND 0.0981562
R15025 VGND VGND.n2435 0.0981562
R15026 VGND.n2430 VGND 0.0981562
R15027 VGND VGND.n1593 0.0981562
R15028 VGND.n1609 VGND 0.0981562
R15029 VGND.n1615 VGND 0.0981562
R15030 VGND.n1619 VGND 0.0981562
R15031 VGND.n1627 VGND 0.0981562
R15032 VGND VGND.n1589 0.0981562
R15033 VGND.n1543 VGND 0.0981562
R15034 VGND VGND.n1579 0.0981562
R15035 VGND.n1574 VGND 0.0981562
R15036 VGND VGND.n1565 0.0981562
R15037 VGND VGND.n1564 0.0981562
R15038 VGND VGND.n2045 0.0981562
R15039 VGND.n2039 VGND 0.0981562
R15040 VGND VGND.n2038 0.0981562
R15041 VGND VGND.n2031 0.0981562
R15042 VGND VGND.n2020 0.0981562
R15043 VGND.n1765 VGND 0.0981562
R15044 VGND.n1784 VGND 0.0981562
R15045 VGND.n1785 VGND 0.0981562
R15046 VGND.n1788 VGND 0.0981562
R15047 VGND.n1733 VGND 0.0981562
R15048 VGND VGND.n1729 0.0981562
R15049 VGND.n1725 VGND 0.0981562
R15050 VGND VGND.n1722 0.0981562
R15051 VGND VGND.n1720 0.0981562
R15052 VGND.n1716 VGND 0.0981562
R15053 VGND VGND.n1712 0.0981562
R15054 VGND VGND.n1707 0.0981562
R15055 VGND VGND.n1697 0.0981562
R15056 VGND VGND 0.0981562
R15057 VGND VGND.n1670 0.0981562
R15058 VGND VGND.n1669 0.0981562
R15059 VGND.n145 VGND 0.0981562
R15060 VGND.n148 VGND 0.0981562
R15061 VGND.n158 VGND 0.0981562
R15062 VGND.n159 VGND 0.0981562
R15063 VGND.n163 VGND 0.0981562
R15064 VGND.n210 VGND 0.0981562
R15065 VGND VGND.n199 0.0981562
R15066 VGND VGND.n191 0.0981562
R15067 VGND.n189 VGND 0.0981562
R15068 VGND VGND.n188 0.0981562
R15069 VGND.n5125 VGND 0.0981562
R15070 VGND.n5105 VGND 0.0981562
R15071 VGND VGND.n5088 0.0981562
R15072 VGND VGND.n5080 0.0981562
R15073 VGND VGND.n5076 0.0981562
R15074 VGND.n5068 VGND 0.0981562
R15075 VGND VGND.n5067 0.0981562
R15076 VGND.n5056 VGND 0.0981562
R15077 VGND.n1969 VGND 0.0981562
R15078 VGND.n1961 VGND 0.0981562
R15079 VGND VGND.n1960 0.0981562
R15080 VGND.n1948 VGND 0.0981562
R15081 VGND.n1942 VGND 0.0981562
R15082 VGND VGND.n1928 0.0981562
R15083 VGND.n1917 VGND 0.0981562
R15084 VGND.n1905 VGND 0.0981562
R15085 VGND VGND 0.0981562
R15086 VGND VGND.n1899 0.0981562
R15087 VGND.n1891 VGND 0.0981562
R15088 VGND.n4228 VGND 0.0981562
R15089 VGND VGND.n4221 0.0981562
R15090 VGND.n4239 VGND 0.0981562
R15091 VGND.n4242 VGND 0.0981562
R15092 VGND VGND.n4252 0.0981562
R15093 VGND.n4259 VGND 0.0981562
R15094 VGND.n4263 VGND 0.0981562
R15095 VGND.n4270 VGND 0.0981562
R15096 VGND VGND 0.0981562
R15097 VGND.n4289 VGND 0.0981562
R15098 VGND.n4292 VGND 0.0981562
R15099 VGND.n4296 VGND 0.0981562
R15100 VGND.n4457 VGND 0.0981562
R15101 VGND.n4445 VGND 0.0981562
R15102 VGND VGND.n4444 0.0981562
R15103 VGND.n4433 VGND 0.0981562
R15104 VGND VGND.n4413 0.0981562
R15105 VGND VGND.n4406 0.0981562
R15106 VGND VGND.n4404 0.0981562
R15107 VGND VGND.n4403 0.0981562
R15108 VGND.n4397 VGND 0.0981562
R15109 VGND VGND.n4396 0.0981562
R15110 VGND.n4386 VGND 0.0981562
R15111 VGND VGND.n4385 0.0981562
R15112 VGND.n4888 VGND 0.0981562
R15113 VGND.n4900 VGND 0.0981562
R15114 VGND VGND 0.0981562
R15115 VGND.n4911 VGND 0.0981562
R15116 VGND.n4965 VGND 0.0981562
R15117 VGND VGND.n4963 0.0981562
R15118 VGND VGND.n4960 0.0981562
R15119 VGND VGND 0.0981562
R15120 VGND VGND.n4938 0.0981562
R15121 VGND.n4933 VGND 0.0981562
R15122 VGND VGND.n4932 0.0981562
R15123 VGND.n4 VGND 0.0981562
R15124 VGND.n15 VGND 0.0981562
R15125 VGND.n5593 VGND 0.0981562
R15126 VGND.n5585 VGND 0.0981562
R15127 VGND.n5579 VGND 0.0981562
R15128 VGND VGND.n5574 0.0981562
R15129 VGND.n5210 VGND 0.0981562
R15130 VGND.n5217 VGND 0.0981562
R15131 VGND VGND 0.0981562
R15132 VGND.n5248 VGND 0.0981562
R15133 VGND.n5262 VGND 0.0981562
R15134 VGND VGND 0.0981562
R15135 VGND.n5336 VGND 0.0981562
R15136 VGND.n5351 VGND 0.0981562
R15137 VGND.n5362 VGND 0.0981562
R15138 VGND.n5367 VGND 0.0981562
R15139 VGND VGND 0.0981562
R15140 VGND.n5386 VGND 0.0981562
R15141 VGND.n5407 VGND 0.0981562
R15142 VGND.n5413 VGND 0.0981562
R15143 VGND.n5464 VGND 0.0981562
R15144 VGND.n5471 VGND 0.0981562
R15145 VGND VGND 0.0981562
R15146 VGND.n5479 VGND 0.0981562
R15147 VGND VGND 0.0981562
R15148 VGND.n5494 VGND 0.0981562
R15149 VGND.n5507 VGND 0.0981562
R15150 VGND VGND 0.0981562
R15151 VGND VGND.n5545 0.0981562
R15152 VGND VGND 0.0981562
R15153 VGND VGND.n5531 0.0981562
R15154 VGND VGND.n5520 0.0981562
R15155 VGND.n2522 VGND.n1450 0.0971438
R15156 VGND.n2520 VGND.n2518 0.0971438
R15157 VGND.n4577 VGND 0.0968542
R15158 VGND VGND.n4793 0.0968542
R15159 VGND.n422 VGND 0.0968542
R15160 VGND.n721 VGND 0.0968542
R15161 VGND.n922 VGND 0.0968542
R15162 VGND VGND.n3532 0.0968542
R15163 VGND.n3172 VGND 0.0968542
R15164 VGND.n3290 VGND 0.0968542
R15165 VGND.n3315 VGND 0.0968542
R15166 VGND.n3432 VGND 0.0968542
R15167 VGND VGND.n3391 0.0968542
R15168 VGND.n1189 VGND 0.0968542
R15169 VGND VGND.n3003 0.0968542
R15170 VGND VGND.n2927 0.0968542
R15171 VGND VGND.n2607 0.0968542
R15172 VGND.n2819 VGND 0.0968542
R15173 VGND VGND.n2817 0.0968542
R15174 VGND VGND.n2215 0.0968542
R15175 VGND VGND.n2440 0.0968542
R15176 VGND VGND.n2429 0.0968542
R15177 VGND VGND.n1696 0.0968542
R15178 VGND VGND.n187 0.0968542
R15179 VGND VGND.n4962 0.0968542
R15180 VGND.n4612 VGND.n4610 0.0955521
R15181 VGND.n4141 VGND.n4140 0.0955521
R15182 VGND.n3625 VGND.n3624 0.0955521
R15183 VGND.n3222 VGND.n3220 0.0955521
R15184 VGND.n2628 VGND.n2627 0.0955521
R15185 VGND.n2275 VGND.n2273 0.0955521
R15186 VGND.n1600 VGND 0.0955521
R15187 VGND.n2056 VGND.n2055 0.0955521
R15188 VGND.n5133 VGND.n5132 0.0955521
R15189 VGND.n4462 VGND.n4461 0.0955521
R15190 VGND VGND.n4456 0.0955521
R15191 VGND.n5319 VGND.n5317 0.0955521
R15192 VGND.n5421 VGND 0.0946285
R15193 VGND VGND.n294 0.0943569
R15194 VGND.n3674 VGND.n3670 0.0900938
R15195 VGND.n329 VGND 0.0890417
R15196 VGND.n358 VGND 0.0890417
R15197 VGND.n4666 VGND 0.0890417
R15198 VGND.n432 VGND 0.0890417
R15199 VGND.n4037 VGND 0.0890417
R15200 VGND VGND.n3780 0.0890417
R15201 VGND VGND.n3741 0.0890417
R15202 VGND.n3822 VGND 0.0890417
R15203 VGND.n3842 VGND 0.0890417
R15204 VGND.n851 VGND 0.0890417
R15205 VGND VGND.n823 0.0890417
R15206 VGND.n803 VGND 0.0890417
R15207 VGND VGND.n3596 0.0890417
R15208 VGND VGND.n3578 0.0890417
R15209 VGND.n3509 VGND 0.0890417
R15210 VGND VGND.n3170 0.0890417
R15211 VGND.n1156 VGND 0.0890417
R15212 VGND VGND.n1228 0.0890417
R15213 VGND VGND 0.0890417
R15214 VGND.n2944 VGND 0.0890417
R15215 VGND.n1379 VGND 0.0890417
R15216 VGND.n2599 VGND 0.0890417
R15217 VGND.n2152 VGND 0.0890417
R15218 VGND.n2156 VGND 0.0890417
R15219 VGND VGND.n2204 0.0890417
R15220 VGND.n2320 VGND 0.0890417
R15221 VGND.n2336 VGND 0.0890417
R15222 VGND.n2491 VGND 0.0890417
R15223 VGND VGND.n2452 0.0890417
R15224 VGND VGND.n2044 0.0890417
R15225 VGND VGND.n2036 0.0890417
R15226 VGND VGND.n1702 0.0890417
R15227 VGND VGND.n208 0.0890417
R15228 VGND.n5113 VGND 0.0890417
R15229 VGND VGND.n1940 0.0890417
R15230 VGND VGND.n1904 0.0890417
R15231 VGND.n4904 VGND 0.0890417
R15232 VGND.n5371 VGND 0.0890417
R15233 VGND VGND.n4585 0.0877396
R15234 VGND.n4661 VGND 0.0877396
R15235 VGND VGND.n4802 0.0877396
R15236 VGND VGND.n481 0.0877396
R15237 VGND.n526 VGND 0.0877396
R15238 VGND VGND.n4088 0.0877396
R15239 VGND.n705 VGND 0.0877396
R15240 VGND.n3930 VGND 0.0877396
R15241 VGND VGND.n824 0.0877396
R15242 VGND.n909 VGND 0.0877396
R15243 VGND VGND.n3570 0.0877396
R15244 VGND.n3196 VGND 0.0877396
R15245 VGND.n3270 VGND 0.0877396
R15246 VGND VGND.n3403 0.0877396
R15247 VGND.n1238 VGND 0.0877396
R15248 VGND VGND.n3012 0.0877396
R15249 VGND VGND.n1350 0.0877396
R15250 VGND VGND.n2221 0.0877396
R15251 VGND.n2316 VGND 0.0877396
R15252 VGND VGND.n2467 0.0877396
R15253 VGND.n1628 VGND 0.0877396
R15254 VGND.n1758 VGND 0.0877396
R15255 VGND.n1703 VGND 0.0877396
R15256 VGND VGND.n209 0.0877396
R15257 VGND VGND.n5087 0.0877396
R15258 VGND VGND.n1927 0.0877396
R15259 VGND.n4258 VGND 0.0877396
R15260 VGND VGND.n4412 0.0877396
R15261 VGND VGND.n4411 0.0877396
R15262 VGND.n5202 VGND 0.0877396
R15263 VGND.n5369 VGND 0.0877396
R15264 VGND.n5565 VGND 0.0877396
R15265 VGND.n4650 VGND 0.0864375
R15266 VGND.n4822 VGND 0.0864375
R15267 VGND VGND.n3974 0.0864375
R15268 VGND.n1083 VGND 0.0864375
R15269 VGND.n3274 VGND 0.0864375
R15270 VGND VGND.n1276 0.0864375
R15271 VGND.n2855 VGND 0.0864375
R15272 VGND.n1408 VGND 0.0864375
R15273 VGND VGND.n2806 0.0864375
R15274 VGND VGND.n2490 0.0864375
R15275 VGND VGND.n2054 0.0864375
R15276 VGND VGND.n1958 0.0864375
R15277 VGND.n4245 VGND 0.0864375
R15278 VGND VGND.n4432 0.0864375
R15279 VGND VGND.n4431 0.0864375
R15280 VGND.n785 VGND.n750 0.0838333
R15281 VGND.n3158 VGND.n3152 0.0838333
R15282 VGND.n1203 VGND.n1118 0.0838333
R15283 VGND.n1449 VGND.n1448 0.0838333
R15284 VGND.n2180 VGND.n2114 0.0838333
R15285 VGND.n1552 VGND.n1512 0.0838333
R15286 VGND.n181 VGND.n90 0.0838333
R15287 VGND.n4510 VGND 0.0830437
R15288 VGND.n269 VGND 0.0830437
R15289 VGND.n1491 VGND 0.0828946
R15290 VGND.n4551 VGND 0.0826382
R15291 VGND.n4778 VGND 0.0826382
R15292 VGND.n4097 VGND 0.0826382
R15293 VGND VGND.n561 0.0826382
R15294 VGND.n464 VGND 0.0826382
R15295 VGND.n4008 VGND 0.0826382
R15296 VGND.n4027 VGND 0.0826382
R15297 VGND.n3803 VGND 0.0826382
R15298 VGND VGND.n3850 0.0826382
R15299 VGND.n3851 VGND 0.0826382
R15300 VGND.n3975 VGND 0.0826382
R15301 VGND.n3935 VGND 0.0826382
R15302 VGND VGND.n3472 0.0826382
R15303 VGND VGND.n3514 0.0826382
R15304 VGND.n3241 VGND 0.0826382
R15305 VGND VGND.n1073 0.0826382
R15306 VGND.n3185 VGND 0.0826382
R15307 VGND.n2889 VGND 0.0826382
R15308 VGND.n2621 VGND 0.0826382
R15309 VGND.n1371 VGND 0.0826382
R15310 VGND.n2822 VGND 0.0826382
R15311 VGND.n2781 VGND 0.0826382
R15312 VGND.n2144 VGND 0.0826382
R15313 VGND.n2313 VGND 0.0826382
R15314 VGND.n2046 VGND 0.0826382
R15315 VGND.n1604 VGND 0.0826382
R15316 VGND VGND.n1608 0.0826382
R15317 VGND.n1616 VGND 0.0826382
R15318 VGND.n1567 VGND 0.0826382
R15319 VGND.n1566 VGND 0.0826382
R15320 VGND VGND.n169 0.0826382
R15321 VGND.n200 VGND 0.0826382
R15322 VGND.n4260 VGND 0.0826382
R15323 VGND.n4407 VGND 0.0826382
R15324 VGND VGND.n4884 0.0826382
R15325 VGND.n4885 VGND 0.0826382
R15326 VGND VGND.n411 0.0822696
R15327 VGND.n3184 VGND 0.0822696
R15328 VGND.n3061 VGND 0.0822696
R15329 VGND.n566 VGND 0.0799271
R15330 VGND.n4370 VGND 0.0799271
R15331 VGND.n4857 VGND.n4856 0.0773229
R15332 VGND.n4007 VGND.n4004 0.0773229
R15333 VGND.n3982 VGND.n3981 0.0773229
R15334 VGND.n3449 VGND.n3448 0.0773229
R15335 VGND.n2849 VGND.n2848 0.0773229
R15336 VGND.n2826 VGND.n2825 0.0773229
R15337 VGND.n2508 VGND.n2507 0.0773229
R15338 VGND.n2000 VGND.n1741 0.0773229
R15339 VGND.n1978 VGND.n1977 0.0773229
R15340 VGND.n5460 VGND.n5457 0.0773229
R15341 VGND.n4418 VGND.n4417 0.0753538
R15342 VGND.n3156 VGND.n3155 0.0753538
R15343 VGND.n1128 VGND.n1127 0.0753538
R15344 VGND.n2865 VGND.n2864 0.0753538
R15345 VGND.n2557 VGND.n2555 0.0685851
R15346 VGND.n3675 VGND.n3674 0.0618937
R15347 VGND.n3672 VGND.n3671 0.0618937
R15348 VGND.n368 VGND 0.0616979
R15349 VGND.n1376 VGND 0.0605028
R15350 VGND.n2523 VGND.n2522 0.0548437
R15351 VGND.n2520 VGND.n2519 0.0548437
R15352 VGND.n4297 VGND 0.0512812
R15353 VGND.n5263 VGND 0.0512812
R15354 VGND.n4599 VGND.n4598 0.0460729
R15355 VGND.n4714 VGND.n299 0.0460729
R15356 VGND.n4155 VGND.n4154 0.0460729
R15357 VGND.n594 VGND.n593 0.0460729
R15358 VGND.n3720 VGND.n3719 0.0460729
R15359 VGND.n637 VGND.n636 0.0460729
R15360 VGND.n3639 VGND.n3638 0.0460729
R15361 VGND.n989 VGND.n988 0.0460729
R15362 VGND.n3209 VGND.n3208 0.0460729
R15363 VGND.n1029 VGND.n1028 0.0460729
R15364 VGND.n3075 VGND.n3074 0.0460729
R15365 VGND.n1267 VGND.n1266 0.0460729
R15366 VGND.n2573 VGND.n1342 0.0460729
R15367 VGND.n2701 VGND.n1334 0.0460729
R15368 VGND.n2245 VGND.n2244 0.0460729
R15369 VGND.n2366 VGND.n1478 0.0460729
R15370 VGND.n2070 VGND.n2069 0.0460729
R15371 VGND.n1820 VGND.n1819 0.0460729
R15372 VGND.n5147 VGND.n5146 0.0460729
R15373 VGND.n124 VGND.n123 0.0460729
R15374 VGND.n4470 VGND.n4469 0.0460729
R15375 VGND.n4366 VGND.n4365 0.0460729
R15376 VGND.n5311 VGND.n5310 0.0460729
R15377 VGND.n5443 VGND.n5442 0.0460729
R15378 VGND.n4307 VGND.n4306 0.0421667
R15379 VGND.n4534 VGND 0.0395625
R15380 VGND VGND.n4164 0.0395625
R15381 VGND.n3711 VGND 0.0395625
R15382 VGND VGND.n3648 0.0395625
R15383 VGND.n3136 VGND 0.0395625
R15384 VGND VGND.n3084 0.0395625
R15385 VGND.n2564 VGND 0.0395625
R15386 VGND VGND.n2254 0.0395625
R15387 VGND VGND.n2079 0.0395625
R15388 VGND VGND.n5156 0.0395625
R15389 VGND.n4646 VGND 0.0343542
R15390 VGND.n1080 VGND 0.0343542
R15391 VGND.n3271 VGND 0.0343542
R15392 VGND VGND.n1156 0.0343542
R15393 VGND.n2849 VGND 0.0343542
R15394 VGND.n1276 VGND 0.0343542
R15395 VGND VGND.n1370 0.0343542
R15396 VGND VGND.n1407 0.0343542
R15397 VGND VGND.n2579 0.0343542
R15398 VGND.n2606 VGND 0.0343542
R15399 VGND.n2807 VGND 0.0343542
R15400 VGND.n2491 VGND 0.0343542
R15401 VGND.n2055 VGND 0.0343542
R15402 VGND.n4433 VGND 0.0343542
R15403 VGND.n4432 VGND 0.0343542
R15404 VGND.n4586 VGND 0.0330521
R15405 VGND VGND.n4660 0.0330521
R15406 VGND.n4803 VGND 0.0330521
R15407 VGND.n482 VGND 0.0330521
R15408 VGND.n4096 VGND 0.0330521
R15409 VGND VGND.n704 0.0330521
R15410 VGND VGND.n3802 0.0330521
R15411 VGND.n3934 VGND 0.0330521
R15412 VGND.n825 VGND 0.0330521
R15413 VGND VGND.n767 0.0330521
R15414 VGND.n3571 VGND 0.0330521
R15415 VGND VGND.n1092 0.0330521
R15416 VGND.n3267 VGND 0.0330521
R15417 VGND VGND.n1185 0.0330521
R15418 VGND.n3013 VGND 0.0330521
R15419 VGND.n2944 VGND 0.0330521
R15420 VGND.n1403 VGND 0.0330521
R15421 VGND VGND.n2649 0.0330521
R15422 VGND VGND.n2736 0.0330521
R15423 VGND.n2222 VGND 0.0330521
R15424 VGND VGND.n1487 0.0330521
R15425 VGND.n2468 VGND 0.0330521
R15426 VGND VGND.n1627 0.0330521
R15427 VGND.n2020 VGND 0.0330521
R15428 VGND.n210 VGND 0.0330521
R15429 VGND.n1928 VGND 0.0330521
R15430 VGND.n4252 VGND 0.0330521
R15431 VGND VGND.n4259 0.0330521
R15432 VGND VGND.n4296 0.0330521
R15433 VGND.n4412 VGND 0.0330521
R15434 VGND.n4965 VGND 0.0330521
R15435 VGND.n5574 VGND 0.0330521
R15436 VGND VGND.n5262 0.0330521
R15437 VGND VGND.n5367 0.0330521
R15438 VGND VGND.n5507 0.0330521
R15439 VGND.n326 VGND 0.03175
R15440 VGND.n4574 VGND 0.03175
R15441 VGND.n4661 VGND 0.03175
R15442 VGND.n429 VGND 0.03175
R15443 VGND.n465 VGND 0.03175
R15444 VGND.n4098 VGND 0.03175
R15445 VGND VGND.n547 0.03175
R15446 VGND VGND.n4026 0.03175
R15447 VGND.n4034 VGND 0.03175
R15448 VGND VGND.n678 0.03175
R15449 VGND VGND.n718 0.03175
R15450 VGND.n3742 VGND 0.03175
R15451 VGND.n3936 VGND 0.03175
R15452 VGND.n3900 VGND 0.03175
R15453 VGND.n824 VGND 0.03175
R15454 VGND.n812 VGND 0.03175
R15455 VGND.n806 VGND 0.03175
R15456 VGND.n3597 VGND 0.03175
R15457 VGND.n3581 VGND 0.03175
R15458 VGND VGND.n3507 0.03175
R15459 VGND VGND.n1059 0.03175
R15460 VGND.n3186 VGND 0.03175
R15461 VGND.n3171 VGND 0.03175
R15462 VGND VGND.n3240 0.03175
R15463 VGND.n1153 VGND 0.03175
R15464 VGND.n1229 VGND 0.03175
R15465 VGND.n2911 VGND 0.03175
R15466 VGND VGND.n1378 0.03175
R15467 VGND.n2806 VGND 0.03175
R15468 VGND VGND.n2137 0.03175
R15469 VGND VGND.n2151 0.03175
R15470 VGND.n2153 VGND 0.03175
R15471 VGND.n2333 VGND 0.03175
R15472 VGND.n2494 VGND 0.03175
R15473 VGND.n2453 VGND 0.03175
R15474 VGND VGND.n1615 0.03175
R15475 VGND VGND.n1628 0.03175
R15476 VGND.n2045 VGND 0.03175
R15477 VGND.n1722 VGND 0.03175
R15478 VGND.n1703 VGND 0.03175
R15479 VGND.n209 VGND 0.03175
R15480 VGND.n5116 VGND 0.03175
R15481 VGND.n1941 VGND 0.03175
R15482 VGND.n1905 VGND 0.03175
R15483 VGND.n4411 VGND 0.03175
R15484 VGND.n4900 VGND 0.03175
R15485 VGND VGND.n5369 0.03175
R15486 VGND.n262 VGND.n261 0.0304479
R15487 VGND.n4487 VGND.n4486 0.0304479
R15488 VGND.n4484 VGND.n4206 0.0304479
R15489 VGND.n4540 VGND.n4539 0.0304479
R15490 VGND.n4537 VGND.n4532 0.0304479
R15491 VGND.n283 VGND.n282 0.0304479
R15492 VGND.n4536 VGND.n4535 0.0304479
R15493 VGND.n4742 VGND.n4741 0.0304479
R15494 VGND.n4740 VGND.n4739 0.0304479
R15495 VGND.n385 VGND.n384 0.0304479
R15496 VGND.n4162 VGND.n4161 0.0304479
R15497 VGND.n508 VGND.n507 0.0304479
R15498 VGND.n4163 VGND.n381 0.0304479
R15499 VGND.n578 VGND.n577 0.0304479
R15500 VGND.n576 VGND.n575 0.0304479
R15501 VGND.n3700 VGND.n3699 0.0304479
R15502 VGND.n3715 VGND.n3714 0.0304479
R15503 VGND.n620 VGND.n619 0.0304479
R15504 VGND.n3713 VGND.n3712 0.0304479
R15505 VGND.n3880 VGND.n3879 0.0304479
R15506 VGND.n3878 VGND.n3877 0.0304479
R15507 VGND.n755 VGND.n754 0.0304479
R15508 VGND.n3646 VGND.n3645 0.0304479
R15509 VGND.n892 VGND.n891 0.0304479
R15510 VGND.n3647 VGND.n751 0.0304479
R15511 VGND.n973 VGND.n972 0.0304479
R15512 VGND.n971 VGND.n970 0.0304479
R15513 VGND.n3146 VGND.n3145 0.0304479
R15514 VGND.n3143 VGND.n3131 0.0304479
R15515 VGND.n1014 VGND.n1013 0.0304479
R15516 VGND.n3142 VGND.n3141 0.0304479
R15517 VGND.n3343 VGND.n3342 0.0304479
R15518 VGND.n3341 VGND.n3340 0.0304479
R15519 VGND.n1123 VGND.n1122 0.0304479
R15520 VGND.n3082 VGND.n3081 0.0304479
R15521 VGND.n1287 VGND.n1278 0.0304479
R15522 VGND.n3083 VGND.n1119 0.0304479
R15523 VGND.n1286 VGND.n1280 0.0304479
R15524 VGND.n1285 VGND.n1284 0.0304479
R15525 VGND.n2548 VGND.n2547 0.0304479
R15526 VGND.n2568 VGND.n2567 0.0304479
R15527 VGND.n1313 VGND.n1312 0.0304479
R15528 VGND.n2566 VGND.n2565 0.0304479
R15529 VGND.n2729 VGND.n2728 0.0304479
R15530 VGND.n2727 VGND.n2726 0.0304479
R15531 VGND.n2119 VGND.n2118 0.0304479
R15532 VGND.n2252 VGND.n2251 0.0304479
R15533 VGND.n2400 VGND.n2394 0.0304479
R15534 VGND.n2253 VGND.n2115 0.0304479
R15535 VGND.n2402 VGND.n2401 0.0304479
R15536 VGND.n2393 VGND.n2392 0.0304479
R15537 VGND.n1743 VGND.n1742 0.0304479
R15538 VGND.n2078 VGND.n1513 0.0304479
R15539 VGND.n2012 VGND.n2011 0.0304479
R15540 VGND.n2010 VGND.n2009 0.0304479
R15541 VGND.n1517 VGND.n1516 0.0304479
R15542 VGND.n2077 VGND.n2076 0.0304479
R15543 VGND.n1845 VGND.n1844 0.0304479
R15544 VGND.n5155 VGND.n91 0.0304479
R15545 VGND.n1854 VGND.n1853 0.0304479
R15546 VGND.n1857 VGND.n1855 0.0304479
R15547 VGND.n95 VGND.n94 0.0304479
R15548 VGND.n5154 VGND.n5153 0.0304479
R15549 VGND.n5278 VGND.n5277 0.0304479
R15550 VGND.n5296 VGND.n5295 0.0304479
R15551 VGND.n4483 VGND.n4482 0.0304479
R15552 VGND.n4355 VGND.n4354 0.0304479
R15553 VGND.n4353 VGND.n4352 0.0304479
R15554 VGND VGND.n78 0.0304479
R15555 VGND.n5298 VGND.n5297 0.0304479
R15556 VGND.n5432 VGND.n5431 0.0304479
R15557 VGND.n5430 VGND.n5429 0.0304479
R15558 VGND.n36 VGND.n35 0.0304479
R15559 VGND.n4199 VGND.n4198 0.0265417
R15560 VGND.n4603 VGND.n4602 0.0265417
R15561 VGND.n4143 VGND.n4142 0.0265417
R15562 VGND.n3789 VGND.n3788 0.0265417
R15563 VGND.n3627 VGND.n3626 0.0265417
R15564 VGND.n3213 VGND.n3212 0.0265417
R15565 VGND.n3064 VGND.n3063 0.0265417
R15566 VGND.n2636 VGND.n2635 0.0265417
R15567 VGND.n2233 VGND.n2232 0.0265417
R15568 VGND.n2058 VGND.n2057 0.0265417
R15569 VGND.n5135 VGND.n5134 0.0265417
R15570 VGND.n5288 VGND.n5287 0.0265417
R15571 VGND.n4870 VGND.n4869 0.0259094
R15572 VGND.n4871 VGND.n4870 0.0259094
R15573 VGND.n4190 VGND.n4189 0.0259094
R15574 VGND.n4189 VGND.n4188 0.0259094
R15575 VGND.n277 VGND.n276 0.0259094
R15576 VGND.n374 VGND.n373 0.0259094
R15577 VGND.n373 VGND.n372 0.0259094
R15578 VGND.n3996 VGND.n3995 0.0259094
R15579 VGND.n3681 VGND.n3680 0.0259094
R15580 VGND.n3680 VGND.n3679 0.0259094
R15581 VGND.n614 VGND.n613 0.0259094
R15582 VGND.n744 VGND.n743 0.0259094
R15583 VGND.n743 VGND.n742 0.0259094
R15584 VGND.n3463 VGND.n3462 0.0259094
R15585 VGND.n3110 VGND.n3109 0.0259094
R15586 VGND.n3109 VGND.n3108 0.0259094
R15587 VGND.n1008 VGND.n1007 0.0259094
R15588 VGND.n1112 VGND.n1111 0.0259094
R15589 VGND.n1111 VGND.n1110 0.0259094
R15590 VGND.n2840 VGND.n2839 0.0259094
R15591 VGND.n2529 VGND.n2528 0.0259094
R15592 VGND.n2528 VGND.n2527 0.0259094
R15593 VGND.n1307 VGND.n1306 0.0259094
R15594 VGND.n2108 VGND.n2107 0.0259094
R15595 VGND.n2107 VGND.n2106 0.0259094
R15596 VGND.n2513 VGND.n2512 0.0259094
R15597 VGND.n1830 VGND.n1829 0.0259094
R15598 VGND.n1506 VGND.n1505 0.0259094
R15599 VGND.n1505 VGND.n1504 0.0259094
R15600 VGND.n1983 VGND.n1982 0.0259094
R15601 VGND.n5175 VGND.n5174 0.0259094
R15602 VGND.n5174 VGND.n5173 0.0259094
R15603 VGND.n5192 VGND.n5191 0.0259094
R15604 VGND.n5191 VGND.n5190 0.0259094
R15605 VGND.n4508 VGND.n4507 0.0259094
R15606 VGND.n4507 VGND.n4506 0.0259094
R15607 VGND.n46 VGND.n45 0.0259094
R15608 VGND.n1593 VGND 0.0252396
R15609 VGND.n4457 VGND 0.0252396
R15610 VGND.n4342 VGND.n4341 0.0239375
R15611 VGND.n265 VGND.n264 0.0239375
R15612 VGND.n267 VGND.n266 0.0239375
R15613 VGND.n4488 VGND.n4487 0.0239375
R15614 VGND.n4541 VGND.n4540 0.0239375
R15615 VGND.n4722 VGND.n4721 0.0239375
R15616 VGND.n286 VGND.n285 0.0239375
R15617 VGND.n288 VGND.n287 0.0239375
R15618 VGND VGND.n356 0.0239375
R15619 VGND.n4794 VGND 0.0239375
R15620 VGND.n384 VGND.n383 0.0239375
R15621 VGND.n585 VGND.n584 0.0239375
R15622 VGND.n511 VGND.n510 0.0239375
R15623 VGND.n513 VGND.n512 0.0239375
R15624 VGND.n419 VGND 0.0239375
R15625 VGND.n463 VGND 0.0239375
R15626 VGND.n3701 VGND.n3700 0.0239375
R15627 VGND.n3860 VGND.n3859 0.0239375
R15628 VGND.n623 VGND.n622 0.0239375
R15629 VGND.n625 VGND.n624 0.0239375
R15630 VGND.n754 VGND.n753 0.0239375
R15631 VGND.n980 VGND.n979 0.0239375
R15632 VGND.n895 VGND.n894 0.0239375
R15633 VGND.n897 VGND.n896 0.0239375
R15634 VGND VGND.n921 0.0239375
R15635 VGND.n3533 VGND 0.0239375
R15636 VGND.n3147 VGND.n3146 0.0239375
R15637 VGND.n3323 VGND.n3322 0.0239375
R15638 VGND.n1017 VGND.n1016 0.0239375
R15639 VGND.n1019 VGND.n1018 0.0239375
R15640 VGND VGND.n1104 0.0239375
R15641 VGND.n3287 VGND 0.0239375
R15642 VGND.n3312 VGND 0.0239375
R15643 VGND.n3435 VGND 0.0239375
R15644 VGND.n3392 VGND 0.0239375
R15645 VGND.n1122 VGND.n1121 0.0239375
R15646 VGND.n2957 VGND.n2956 0.0239375
R15647 VGND.n1290 VGND.n1289 0.0239375
R15648 VGND.n1292 VGND.n1291 0.0239375
R15649 VGND VGND.n1188 0.0239375
R15650 VGND.n2928 VGND 0.0239375
R15651 VGND.n2549 VGND.n2548 0.0239375
R15652 VGND.n2709 VGND.n2708 0.0239375
R15653 VGND.n1316 VGND.n1315 0.0239375
R15654 VGND.n1318 VGND.n1317 0.0239375
R15655 VGND.n2608 VGND 0.0239375
R15656 VGND.n2821 VGND 0.0239375
R15657 VGND.n2818 VGND 0.0239375
R15658 VGND.n2118 VGND.n2117 0.0239375
R15659 VGND.n2374 VGND.n2373 0.0239375
R15660 VGND.n2398 VGND.n2397 0.0239375
R15661 VGND.n2396 VGND.n2395 0.0239375
R15662 VGND.n2216 VGND 0.0239375
R15663 VGND.n2441 VGND 0.0239375
R15664 VGND.n2430 VGND 0.0239375
R15665 VGND.n1811 VGND.n1810 0.0239375
R15666 VGND.n1746 VGND.n1745 0.0239375
R15667 VGND.n1748 VGND.n1747 0.0239375
R15668 VGND.n1697 VGND 0.0239375
R15669 VGND.n1516 VGND.n1515 0.0239375
R15670 VGND.n5030 VGND.n5029 0.0239375
R15671 VGND.n1848 VGND.n1847 0.0239375
R15672 VGND.n1850 VGND.n1849 0.0239375
R15673 VGND.n188 VGND 0.0239375
R15674 VGND.n94 VGND.n93 0.0239375
R15675 VGND.n5277 VGND.n5276 0.0239375
R15676 VGND.n4963 VGND 0.0239375
R15677 VGND.n60 VGND.n59 0.0239375
R15678 VGND.n39 VGND.n38 0.0239375
R15679 VGND.n41 VGND.n40 0.0239375
R15680 VGND.n4341 VGND.n4340 0.0226354
R15681 VGND.n4723 VGND.n4722 0.0226354
R15682 VGND VGND.n325 0.0226354
R15683 VGND.n336 VGND 0.0226354
R15684 VGND VGND.n353 0.0226354
R15685 VGND.n4581 VGND 0.0226354
R15686 VGND.n4570 VGND 0.0226354
R15687 VGND VGND.n359 0.0226354
R15688 VGND.n4557 VGND 0.0226354
R15689 VGND.n4552 VGND 0.0226354
R15690 VGND.n4550 VGND 0.0226354
R15691 VGND.n4616 VGND 0.0226354
R15692 VGND VGND.n4658 0.0226354
R15693 VGND VGND.n4666 0.0226354
R15694 VGND VGND.n4670 0.0226354
R15695 VGND VGND.n4672 0.0226354
R15696 VGND.n4702 VGND 0.0226354
R15697 VGND.n4851 VGND 0.0226354
R15698 VGND.n4845 VGND 0.0226354
R15699 VGND.n4837 VGND 0.0226354
R15700 VGND.n4827 VGND 0.0226354
R15701 VGND.n4822 VGND 0.0226354
R15702 VGND.n4806 VGND 0.0226354
R15703 VGND.n4797 VGND 0.0226354
R15704 VGND.n4784 VGND 0.0226354
R15705 VGND.n4781 VGND 0.0226354
R15706 VGND.n4777 VGND 0.0226354
R15707 VGND.n4775 VGND 0.0226354
R15708 VGND.n4766 VGND 0.0226354
R15709 VGND.n4765 VGND 0.0226354
R15710 VGND VGND.n4758 0.0226354
R15711 VGND.n586 VGND.n585 0.0226354
R15712 VGND VGND.n417 0.0226354
R15713 VGND VGND.n436 0.0226354
R15714 VGND.n477 VGND 0.0226354
R15715 VGND.n474 VGND 0.0226354
R15716 VGND.n468 VGND 0.0226354
R15717 VGND.n458 VGND 0.0226354
R15718 VGND.n4136 VGND 0.0226354
R15719 VGND.n4133 VGND 0.0226354
R15720 VGND.n4109 VGND 0.0226354
R15721 VGND.n4101 VGND 0.0226354
R15722 VGND.n526 VGND 0.0226354
R15723 VGND VGND.n537 0.0226354
R15724 VGND VGND.n549 0.0226354
R15725 VGND.n562 VGND 0.0226354
R15726 VGND VGND.n4016 0.0226354
R15727 VGND.n4018 VGND 0.0226354
R15728 VGND VGND.n4022 0.0226354
R15729 VGND VGND.n4031 0.0226354
R15730 VGND VGND.n4037 0.0226354
R15731 VGND.n4089 VGND 0.0226354
R15732 VGND.n4082 VGND 0.0226354
R15733 VGND.n4081 VGND 0.0226354
R15734 VGND VGND.n4043 0.0226354
R15735 VGND VGND.n4046 0.0226354
R15736 VGND.n4057 VGND 0.0226354
R15737 VGND.n3861 VGND.n3860 0.0226354
R15738 VGND.n680 VGND 0.0226354
R15739 VGND.n670 VGND 0.0226354
R15740 VGND VGND.n711 0.0226354
R15741 VGND VGND.n712 0.0226354
R15742 VGND.n658 VGND 0.0226354
R15743 VGND VGND.n720 0.0226354
R15744 VGND VGND.n727 0.0226354
R15745 VGND.n3775 VGND 0.0226354
R15746 VGND.n3751 VGND 0.0226354
R15747 VGND.n3745 VGND 0.0226354
R15748 VGND.n3728 VGND 0.0226354
R15749 VGND VGND.n3818 0.0226354
R15750 VGND.n3819 VGND 0.0226354
R15751 VGND.n3839 VGND 0.0226354
R15752 VGND.n3949 VGND 0.0226354
R15753 VGND.n3937 VGND 0.0226354
R15754 VGND.n3930 VGND 0.0226354
R15755 VGND VGND.n3894 0.0226354
R15756 VGND.n3903 VGND 0.0226354
R15757 VGND.n981 VGND.n980 0.0226354
R15758 VGND.n854 VGND 0.0226354
R15759 VGND.n861 VGND 0.0226354
R15760 VGND.n867 VGND 0.0226354
R15761 VGND.n874 VGND 0.0226354
R15762 VGND.n818 VGND 0.0226354
R15763 VGND.n813 VGND 0.0226354
R15764 VGND.n3620 VGND 0.0226354
R15765 VGND VGND.n762 0.0226354
R15766 VGND.n3596 VGND 0.0226354
R15767 VGND.n3593 VGND 0.0226354
R15768 VGND.n3591 VGND 0.0226354
R15769 VGND.n3590 VGND 0.0226354
R15770 VGND.n3578 VGND 0.0226354
R15771 VGND.n912 VGND 0.0226354
R15772 VGND.n924 VGND 0.0226354
R15773 VGND.n937 VGND 0.0226354
R15774 VGND.n944 VGND 0.0226354
R15775 VGND.n954 VGND 0.0226354
R15776 VGND.n3493 VGND 0.0226354
R15777 VGND.n3500 VGND 0.0226354
R15778 VGND.n3508 VGND 0.0226354
R15779 VGND.n3570 VGND 0.0226354
R15780 VGND.n3565 VGND 0.0226354
R15781 VGND.n3551 VGND 0.0226354
R15782 VGND.n3536 VGND 0.0226354
R15783 VGND.n3530 VGND 0.0226354
R15784 VGND.n3526 VGND 0.0226354
R15785 VGND.n3324 VGND.n3323 0.0226354
R15786 VGND VGND.n1064 0.0226354
R15787 VGND.n1074 VGND 0.0226354
R15788 VGND.n1053 VGND 0.0226354
R15789 VGND VGND.n1090 0.0226354
R15790 VGND.n3192 VGND 0.0226354
R15791 VGND VGND.n1095 0.0226354
R15792 VGND VGND.n1096 0.0226354
R15793 VGND VGND.n1101 0.0226354
R15794 VGND.n3176 VGND 0.0226354
R15795 VGND VGND.n3266 0.0226354
R15796 VGND VGND.n3286 0.0226354
R15797 VGND.n3295 VGND 0.0226354
R15798 VGND.n3304 VGND 0.0226354
R15799 VGND VGND.n3309 0.0226354
R15800 VGND VGND.n3311 0.0226354
R15801 VGND.n3443 VGND 0.0226354
R15802 VGND.n3427 VGND 0.0226354
R15803 VGND.n3416 VGND 0.0226354
R15804 VGND VGND.n1027 0.0226354
R15805 VGND.n3404 VGND 0.0226354
R15806 VGND.n3398 VGND 0.0226354
R15807 VGND.n3384 VGND 0.0226354
R15808 VGND.n3381 VGND 0.0226354
R15809 VGND.n3370 VGND 0.0226354
R15810 VGND.n3362 VGND 0.0226354
R15811 VGND.n2956 VGND.n2955 0.0226354
R15812 VGND.n1161 VGND 0.0226354
R15813 VGND.n1166 VGND 0.0226354
R15814 VGND VGND.n1177 0.0226354
R15815 VGND VGND.n1184 0.0226354
R15816 VGND VGND.n1187 0.0226354
R15817 VGND VGND.n1189 0.0226354
R15818 VGND.n1220 VGND 0.0226354
R15819 VGND.n3057 VGND 0.0226354
R15820 VGND.n3041 VGND 0.0226354
R15821 VGND.n3024 VGND 0.0226354
R15822 VGND.n3016 VGND 0.0226354
R15823 VGND.n3007 VGND 0.0226354
R15824 VGND.n3004 VGND 0.0226354
R15825 VGND.n2998 VGND 0.0226354
R15826 VGND.n2993 VGND 0.0226354
R15827 VGND.n2979 VGND 0.0226354
R15828 VGND.n2974 VGND 0.0226354
R15829 VGND VGND.n2868 0.0226354
R15830 VGND.n2869 VGND 0.0226354
R15831 VGND VGND.n2883 0.0226354
R15832 VGND.n2884 VGND 0.0226354
R15833 VGND VGND.n2893 0.0226354
R15834 VGND.n2942 VGND 0.0226354
R15835 VGND.n2939 VGND 0.0226354
R15836 VGND.n2937 VGND 0.0226354
R15837 VGND.n2931 VGND 0.0226354
R15838 VGND.n2915 VGND 0.0226354
R15839 VGND.n2710 VGND.n2709 0.0226354
R15840 VGND.n1379 VGND 0.0226354
R15841 VGND.n1384 VGND 0.0226354
R15842 VGND VGND.n1395 0.0226354
R15843 VGND VGND.n1402 0.0226354
R15844 VGND VGND.n1414 0.0226354
R15845 VGND.n1416 VGND 0.0226354
R15846 VGND VGND.n1435 0.0226354
R15847 VGND.n1436 VGND 0.0226354
R15848 VGND.n2627 VGND 0.0226354
R15849 VGND.n2612 VGND 0.0226354
R15850 VGND.n2609 VGND 0.0226354
R15851 VGND.n2604 VGND 0.0226354
R15852 VGND.n2599 VGND 0.0226354
R15853 VGND.n2596 VGND 0.0226354
R15854 VGND.n2651 VGND 0.0226354
R15855 VGND.n2657 VGND 0.0226354
R15856 VGND VGND.n2664 0.0226354
R15857 VGND.n2665 VGND 0.0226354
R15858 VGND.n2819 VGND 0.0226354
R15859 VGND VGND.n1333 0.0226354
R15860 VGND.n2795 VGND 0.0226354
R15861 VGND.n2783 VGND 0.0226354
R15862 VGND.n2775 VGND 0.0226354
R15863 VGND.n2755 VGND 0.0226354
R15864 VGND.n2375 VGND.n2374 0.0226354
R15865 VGND VGND.n2143 0.0226354
R15866 VGND.n2127 VGND 0.0226354
R15867 VGND.n2126 VGND 0.0226354
R15868 VGND VGND.n2152 0.0226354
R15869 VGND VGND.n2168 0.0226354
R15870 VGND.n2221 VGND 0.0226354
R15871 VGND.n2214 VGND 0.0226354
R15872 VGND.n2209 VGND 0.0226354
R15873 VGND.n2205 VGND 0.0226354
R15874 VGND.n2199 VGND 0.0226354
R15875 VGND.n2195 VGND 0.0226354
R15876 VGND.n2190 VGND 0.0226354
R15877 VGND.n2186 VGND 0.0226354
R15878 VGND.n2185 VGND 0.0226354
R15879 VGND.n2280 VGND 0.0226354
R15880 VGND VGND.n2287 0.0226354
R15881 VGND.n2288 VGND 0.0226354
R15882 VGND.n2297 VGND 0.0226354
R15883 VGND VGND.n2306 0.0226354
R15884 VGND.n2316 VGND 0.0226354
R15885 VGND VGND.n2326 0.0226354
R15886 VGND VGND.n2349 0.0226354
R15887 VGND.n2350 VGND 0.0226354
R15888 VGND.n2485 VGND 0.0226354
R15889 VGND.n2479 VGND 0.0226354
R15890 VGND.n2471 VGND 0.0226354
R15891 VGND.n2462 VGND 0.0226354
R15892 VGND.n2446 VGND 0.0226354
R15893 VGND.n2442 VGND 0.0226354
R15894 VGND VGND.n2417 0.0226354
R15895 VGND.n2433 VGND 0.0226354
R15896 VGND.n2427 VGND 0.0226354
R15897 VGND.n1812 VGND.n1811 0.0226354
R15898 VGND.n1610 VGND 0.0226354
R15899 VGND VGND.n1626 0.0226354
R15900 VGND.n1587 VGND 0.0226354
R15901 VGND.n1580 VGND 0.0226354
R15902 VGND.n1579 VGND 0.0226354
R15903 VGND.n1565 VGND 0.0226354
R15904 VGND.n2044 VGND 0.0226354
R15905 VGND.n2039 VGND 0.0226354
R15906 VGND.n2022 VGND 0.0226354
R15907 VGND.n1762 VGND 0.0226354
R15908 VGND VGND.n1782 0.0226354
R15909 VGND VGND.n1784 0.0226354
R15910 VGND.n1785 VGND 0.0226354
R15911 VGND.n1736 VGND 0.0226354
R15912 VGND.n1729 VGND 0.0226354
R15913 VGND.n1720 VGND 0.0226354
R15914 VGND.n1713 VGND 0.0226354
R15915 VGND.n1712 VGND 0.0226354
R15916 VGND.n1707 VGND 0.0226354
R15917 VGND.n1673 VGND 0.0226354
R15918 VGND.n1670 VGND 0.0226354
R15919 VGND.n5029 VGND.n5028 0.0226354
R15920 VGND VGND.n144 0.0226354
R15921 VGND.n145 VGND 0.0226354
R15922 VGND VGND.n158 0.0226354
R15923 VGND.n160 VGND 0.0226354
R15924 VGND.n191 VGND 0.0226354
R15925 VGND.n189 VGND 0.0226354
R15926 VGND.n5128 VGND 0.0226354
R15927 VGND.n5108 VGND 0.0226354
R15928 VGND.n5093 VGND 0.0226354
R15929 VGND.n5088 VGND 0.0226354
R15930 VGND.n5077 VGND 0.0226354
R15931 VGND.n5071 VGND 0.0226354
R15932 VGND.n5068 VGND 0.0226354
R15933 VGND.n5059 VGND 0.0226354
R15934 VGND.n1972 VGND 0.0226354
R15935 VGND.n1964 VGND 0.0226354
R15936 VGND.n1961 VGND 0.0226354
R15937 VGND.n1951 VGND 0.0226354
R15938 VGND.n1945 VGND 0.0226354
R15939 VGND.n1930 VGND 0.0226354
R15940 VGND.n1920 VGND 0.0226354
R15941 VGND.n1908 VGND 0.0226354
R15942 VGND.n1894 VGND 0.0226354
R15943 VGND.n1890 VGND 0.0226354
R15944 VGND.n4221 VGND 0.0226354
R15945 VGND VGND.n4241 0.0226354
R15946 VGND.n4253 VGND 0.0226354
R15947 VGND VGND.n4258 0.0226354
R15948 VGND VGND.n4286 0.0226354
R15949 VGND.n4289 VGND 0.0226354
R15950 VGND.n4461 VGND 0.0226354
R15951 VGND.n4448 VGND 0.0226354
R15952 VGND.n4445 VGND 0.0226354
R15953 VGND.n4436 VGND 0.0226354
R15954 VGND.n4421 VGND 0.0226354
R15955 VGND.n4413 VGND 0.0226354
R15956 VGND VGND 0.0226354
R15957 VGND.n4404 VGND 0.0226354
R15958 VGND.n4400 VGND 0.0226354
R15959 VGND.n4397 VGND 0.0226354
R15960 VGND.n4389 VGND 0.0226354
R15961 VGND.n4386 VGND 0.0226354
R15962 VGND.n4373 VGND 0.0226354
R15963 VGND VGND.n4899 0.0226354
R15964 VGND VGND.n4915 0.0226354
R15965 VGND.n4941 VGND 0.0226354
R15966 VGND.n4936 VGND 0.0226354
R15967 VGND.n4933 VGND 0.0226354
R15968 VGND.n12 VGND 0.0226354
R15969 VGND.n5588 VGND 0.0226354
R15970 VGND.n5207 VGND 0.0226354
R15971 VGND VGND.n5245 0.0226354
R15972 VGND VGND.n5261 0.0226354
R15973 VGND VGND.n5333 0.0226354
R15974 VGND.n5348 VGND 0.0226354
R15975 VGND.n5358 VGND 0.0226354
R15976 VGND VGND.n5383 0.0226354
R15977 VGND.n5404 VGND 0.0226354
R15978 VGND.n5410 VGND 0.0226354
R15979 VGND VGND.n5420 0.0226354
R15980 VGND.n5461 VGND 0.0226354
R15981 VGND VGND.n5476 0.0226354
R15982 VGND VGND.n5491 0.0226354
R15983 VGND VGND.n5506 0.0226354
R15984 VGND.n5548 VGND 0.0226354
R15985 VGND.n5534 VGND 0.0226354
R15986 VGND.n5518 VGND 0.0226354
R15987 VGND.n59 VGND.n58 0.0226354
R15988 VGND.n346 VGND 0.0213333
R15989 VGND VGND.n362 0.0213333
R15990 VGND.n4832 VGND 0.0213333
R15991 VGND.n449 VGND 0.0213333
R15992 VGND.n4117 VGND 0.0213333
R15993 VGND VGND.n693 0.0213333
R15994 VGND VGND.n725 0.0213333
R15995 VGND.n733 VGND 0.0213333
R15996 VGND.n3759 VGND 0.0213333
R15997 VGND.n3734 VGND 0.0213333
R15998 VGND VGND.n3838 0.0213333
R15999 VGND.n3977 VGND 0.0213333
R16000 VGND.n3957 VGND 0.0213333
R16001 VGND.n3940 VGND 0.0213333
R16002 VGND.n3914 VGND 0.0213333
R16003 VGND.n837 VGND 0.0213333
R16004 VGND.n791 VGND 0.0213333
R16005 VGND.n3602 VGND 0.0213333
R16006 VGND.n3485 VGND 0.0213333
R16007 VGND VGND.n3492 0.0213333
R16008 VGND.n1065 VGND 0.0213333
R16009 VGND.n3237 VGND 0.0213333
R16010 VGND.n3247 VGND 0.0213333
R16011 VGND.n3256 VGND 0.0213333
R16012 VGND.n3410 VGND 0.0213333
R16013 VGND.n1208 VGND 0.0213333
R16014 VGND.n3049 VGND 0.0213333
R16015 VGND.n2598 VGND 0.0213333
R16016 VGND.n2789 VGND 0.0213333
R16017 VGND.n2204 VGND 0.0213333
R16018 VGND VGND.n2279 0.0213333
R16019 VGND.n2307 VGND 0.0213333
R16020 VGND VGND.n2312 0.0213333
R16021 VGND VGND.n2332 0.0213333
R16022 VGND.n2342 VGND 0.0213333
R16023 VGND.n2354 VGND 0.0213333
R16024 VGND.n2495 VGND 0.0213333
R16025 VGND.n2030 VGND 0.0213333
R16026 VGND.n1778 VGND 0.0213333
R16027 VGND.n5094 VGND 0.0213333
R16028 VGND.n1959 VGND 0.0213333
R16029 VGND.n1942 VGND 0.0213333
R16030 VGND.n4332 VGND.n4331 0.0202124
R16031 VGND.n4518 VGND.n4517 0.0202124
R16032 VGND.n4177 VGND.n4176 0.0202124
R16033 VGND.n3688 VGND.n3687 0.0202124
R16034 VGND.n3664 VGND.n3663 0.0202124
R16035 VGND.n3117 VGND.n3116 0.0202124
R16036 VGND.n3097 VGND.n3096 0.0202124
R16037 VGND.n2536 VGND.n2535 0.0202124
R16038 VGND.n1498 VGND.n1497 0.0202124
R16039 VGND.n2095 VGND.n2094 0.0202124
R16040 VGND.n81 VGND.n80 0.0202124
R16041 VGND.n5196 VGND.n5195 0.0202124
R16042 VGND.n5187 VGND.n5186 0.0202124
R16043 VGND.n4495 VGND.n4494 0.0202124
R16044 VGND.n4499 VGND.n4498 0.0202124
R16045 VGND.n4343 VGND.n4342 0.0200312
R16046 VGND.n268 VGND.n267 0.0200312
R16047 VGND.n4205 VGND.n4204 0.0200312
R16048 VGND.n4203 VGND.n4202 0.0200312
R16049 VGND.n4198 VGND.n4197 0.0200312
R16050 VGND.n4196 VGND.n4195 0.0200312
R16051 VGND.n4531 VGND.n4530 0.0200312
R16052 VGND.n4529 VGND.n305 0.0200312
R16053 VGND.n4604 VGND.n4603 0.0200312
R16054 VGND.n4606 VGND.n4605 0.0200312
R16055 VGND.n4721 VGND.n4720 0.0200312
R16056 VGND.n289 VGND.n288 0.0200312
R16057 VGND.n4595 VGND.n4594 0.0200312
R16058 VGND.n4597 VGND.n4596 0.0200312
R16059 VGND.n4733 VGND.n290 0.0200312
R16060 VGND.n4160 VGND.n4159 0.0200312
R16061 VGND.n4158 VGND.n4157 0.0200312
R16062 VGND.n4144 VGND.n4143 0.0200312
R16063 VGND.n4146 VGND.n4145 0.0200312
R16064 VGND.n584 VGND.n517 0.0200312
R16065 VGND.n514 VGND.n513 0.0200312
R16066 VGND.n491 VGND.n388 0.0200312
R16067 VGND.n4153 VGND.n4152 0.0200312
R16068 VGND.n569 VGND.n506 0.0200312
R16069 VGND.n4023 VGND 0.0200312
R16070 VGND.n4067 VGND 0.0200312
R16071 VGND.n3717 VGND.n3716 0.0200312
R16072 VGND.n3792 VGND.n3718 0.0200312
R16073 VGND.n3788 VGND.n3787 0.0200312
R16074 VGND.n3786 VGND.n3785 0.0200312
R16075 VGND.n3859 VGND.n3858 0.0200312
R16076 VGND.n626 VGND.n625 0.0200312
R16077 VGND VGND.n732 0.0200312
R16078 VGND.n3722 VGND.n3721 0.0200312
R16079 VGND.n3871 VGND.n627 0.0200312
R16080 VGND.n3644 VGND.n3643 0.0200312
R16081 VGND.n3642 VGND.n3641 0.0200312
R16082 VGND.n3628 VGND.n3627 0.0200312
R16083 VGND.n3630 VGND.n3629 0.0200312
R16084 VGND.n979 VGND.n901 0.0200312
R16085 VGND.n898 VGND.n897 0.0200312
R16086 VGND.n879 VGND.n758 0.0200312
R16087 VGND.n3637 VGND.n3636 0.0200312
R16088 VGND.n966 VGND.n890 0.0200312
R16089 VGND.n3130 VGND.n3129 0.0200312
R16090 VGND.n3128 VGND.n1048 0.0200312
R16091 VGND.n3214 VGND.n3213 0.0200312
R16092 VGND.n3216 VGND.n3215 0.0200312
R16093 VGND.n3322 VGND.n3321 0.0200312
R16094 VGND.n1020 VGND.n1019 0.0200312
R16095 VGND.n3205 VGND.n3204 0.0200312
R16096 VGND.n3207 VGND.n3206 0.0200312
R16097 VGND.n3334 VGND.n1021 0.0200312
R16098 VGND.n3080 VGND.n3079 0.0200312
R16099 VGND.n3078 VGND.n3077 0.0200312
R16100 VGND.n3065 VGND.n3064 0.0200312
R16101 VGND.n3067 VGND.n3066 0.0200312
R16102 VGND.n2958 VGND.n2957 0.0200312
R16103 VGND.n1293 VGND.n1292 0.0200312
R16104 VGND.n1243 VGND.n1126 0.0200312
R16105 VGND.n3073 VGND.n3072 0.0200312
R16106 VGND VGND.n2876 0.0200312
R16107 VGND VGND.n2888 0.0200312
R16108 VGND.n2570 VGND.n2569 0.0200312
R16109 VGND.n2572 VGND.n2571 0.0200312
R16110 VGND.n2635 VGND.n2634 0.0200312
R16111 VGND.n2633 VGND.n2632 0.0200312
R16112 VGND.n2708 VGND.n2707 0.0200312
R16113 VGND.n1319 VGND.n1318 0.0200312
R16114 VGND.n2640 VGND.n2639 0.0200312
R16115 VGND.n2575 VGND.n2574 0.0200312
R16116 VGND.n2720 VGND.n1320 0.0200312
R16117 VGND.n2250 VGND.n2249 0.0200312
R16118 VGND.n2248 VGND.n2247 0.0200312
R16119 VGND.n2234 VGND.n2233 0.0200312
R16120 VGND.n2236 VGND.n2235 0.0200312
R16121 VGND.n2373 VGND.n2372 0.0200312
R16122 VGND.n2395 VGND.n1461 0.0200312
R16123 VGND.n2231 VGND.n2230 0.0200312
R16124 VGND.n2243 VGND.n2242 0.0200312
R16125 VGND.n2386 VGND.n2384 0.0200312
R16126 VGND.n1810 VGND.n1752 0.0200312
R16127 VGND.n1749 VGND.n1748 0.0200312
R16128 VGND.n1636 VGND.n1520 0.0200312
R16129 VGND.n2068 VGND.n2067 0.0200312
R16130 VGND.n2003 VGND.n2001 0.0200312
R16131 VGND.n1723 VGND 0.0200312
R16132 VGND.n2075 VGND.n2074 0.0200312
R16133 VGND.n2073 VGND.n2072 0.0200312
R16134 VGND.n2059 VGND.n2058 0.0200312
R16135 VGND.n2061 VGND.n2060 0.0200312
R16136 VGND.n5031 VGND.n5030 0.0200312
R16137 VGND.n1851 VGND.n1850 0.0200312
R16138 VGND.n218 VGND.n98 0.0200312
R16139 VGND.n5145 VGND.n5144 0.0200312
R16140 VGND.n1864 VGND.n1863 0.0200312
R16141 VGND.n5152 VGND.n5151 0.0200312
R16142 VGND.n5150 VGND.n5149 0.0200312
R16143 VGND.n5136 VGND.n5135 0.0200312
R16144 VGND.n5138 VGND.n5137 0.0200312
R16145 VGND.n5294 VGND.n5293 0.0200312
R16146 VGND.n5292 VGND.n5291 0.0200312
R16147 VGND.n5287 VGND.n5286 0.0200312
R16148 VGND.n5285 VGND.n5284 0.0200312
R16149 VGND.n4231 VGND 0.0200312
R16150 VGND.n4474 VGND.n4472 0.0200312
R16151 VGND.n4468 VGND.n4467 0.0200312
R16152 VGND.n4346 VGND.n260 0.0200312
R16153 VGND.n5308 VGND.n5307 0.0200312
R16154 VGND.n5313 VGND.n5312 0.0200312
R16155 VGND.n5423 VGND.n34 0.0200312
R16156 VGND.n61 VGND.n60 0.0200312
R16157 VGND.n42 VGND.n41 0.0200312
R16158 VGND.n4533 VGND.n367 0.0187292
R16159 VGND.n4610 VGND.n4609 0.0187292
R16160 VGND.n4713 VGND.n4712 0.0187292
R16161 VGND.n4166 VGND.n4165 0.0187292
R16162 VGND.n4149 VGND.n4141 0.0187292
R16163 VGND.n567 VGND.n566 0.0187292
R16164 VGND.n3710 VGND.n3709 0.0187292
R16165 VGND.n3782 VGND.n3781 0.0187292
R16166 VGND.n3651 VGND.n3650 0.0187292
R16167 VGND.n3633 VGND.n3625 0.0187292
R16168 VGND.n965 VGND.n964 0.0187292
R16169 VGND.n3135 VGND.n3134 0.0187292
R16170 VGND.n3220 VGND.n3219 0.0187292
R16171 VGND.n3086 VGND.n3085 0.0187292
R16172 VGND.n3070 VGND.n3062 0.0187292
R16173 VGND.n2965 VGND.n2963 0.0187292
R16174 VGND.n2563 VGND.n2560 0.0187292
R16175 VGND.n2629 VGND.n2628 0.0187292
R16176 VGND.n2700 VGND.n2699 0.0187292
R16177 VGND.n2256 VGND.n2255 0.0187292
R16178 VGND.n2365 VGND.n2364 0.0187292
R16179 VGND.n2082 VGND.n2081 0.0187292
R16180 VGND.n2064 VGND.n2056 0.0187292
R16181 VGND.n1808 VGND.n1807 0.0187292
R16182 VGND.n5159 VGND.n5158 0.0187292
R16183 VGND.n5141 VGND.n5133 0.0187292
R16184 VGND.n5035 VGND.n5034 0.0187292
R16185 VGND.n4306 VGND.n4304 0.0187292
R16186 VGND.n4463 VGND.n4462 0.0187292
R16187 VGND.n4370 VGND.n4369 0.0187292
R16188 VGND.n5265 VGND.n5264 0.0187292
R16189 VGND.n5317 VGND.n5316 0.0187292
R16190 VGND.n5282 VGND.n5281 0.0174271
R16191 VGND.n969 VGND.n966 0.0173894
R16192 VGND.n1283 VGND.n1281 0.0172616
R16193 VGND.n4874 VGND.n4873 0.0168788
R16194 VGND.n4191 VGND.n4186 0.0168788
R16195 VGND.n278 VGND.n275 0.0168788
R16196 VGND.n4864 VGND.n4863 0.0168788
R16197 VGND.n375 VGND.n370 0.0168788
R16198 VGND.n3997 VGND.n3994 0.0168788
R16199 VGND.n606 VGND.n605 0.0168788
R16200 VGND.n3682 VGND.n3677 0.0168788
R16201 VGND.n615 VGND.n612 0.0168788
R16202 VGND.n3989 VGND.n3988 0.0168788
R16203 VGND.n745 VGND.n740 0.0168788
R16204 VGND.n3464 VGND.n3461 0.0168788
R16205 VGND.n1000 VGND.n999 0.0168788
R16206 VGND.n3111 VGND.n3106 0.0168788
R16207 VGND.n1009 VGND.n1006 0.0168788
R16208 VGND.n3456 VGND.n3455 0.0168788
R16209 VGND.n1113 VGND.n1108 0.0168788
R16210 VGND.n2841 VGND.n2838 0.0168788
R16211 VGND.n1299 VGND.n1298 0.0168788
R16212 VGND.n2530 VGND.n2525 0.0168788
R16213 VGND.n1308 VGND.n1305 0.0168788
R16214 VGND.n2833 VGND.n2832 0.0168788
R16215 VGND.n2109 VGND.n2104 0.0168788
R16216 VGND.n1457 VGND.n1455 0.0168788
R16217 VGND.n2516 VGND.n2515 0.0168788
R16218 VGND.n1993 VGND.n1991 0.0168788
R16219 VGND.n1833 VGND.n1832 0.0168788
R16220 VGND.n1507 VGND.n1502 0.0168788
R16221 VGND.n1840 VGND.n1838 0.0168788
R16222 VGND.n1986 VGND.n1985 0.0168788
R16223 VGND.n5176 VGND.n5171 0.0168788
R16224 VGND.n5194 VGND.n5193 0.0168788
R16225 VGND.n5189 VGND.n5188 0.0168788
R16226 VGND.n4509 VGND.n4504 0.0168788
R16227 VGND.n5452 VGND.n5450 0.0168788
R16228 VGND.n49 VGND.n48 0.0168788
R16229 VGND.n4592 VGND.n4591 0.0166873
R16230 VGND.n3797 VGND.n3796 0.0166873
R16231 VGND.n882 VGND.n881 0.0166873
R16232 VGND.n1246 VGND.n1245 0.0166873
R16233 VGND.n2643 VGND.n2642 0.0166873
R16234 VGND.n2228 VGND.n2227 0.0166873
R16235 VGND.n1639 VGND.n1638 0.0166873
R16236 VGND.n1284 VGND.n1283 0.0166226
R16237 VGND.n970 VGND.n969 0.0164946
R16238 VGND.n4337 VGND.n4336 0.016125
R16239 VGND.n4490 VGND.n4489 0.016125
R16240 VGND.n4543 VGND.n4542 0.016125
R16241 VGND.n4727 VGND.n4726 0.016125
R16242 VGND.n4547 VGND.n4546 0.016125
R16243 VGND VGND.n4714 0.016125
R16244 VGND.n4731 VGND.n4730 0.016125
R16245 VGND.n382 VGND.n379 0.016125
R16246 VGND.n590 VGND.n589 0.016125
R16247 VGND.n4169 VGND.n4168 0.016125
R16248 VGND VGND.n594 0.016125
R16249 VGND.n583 VGND.n582 0.016125
R16250 VGND.n3703 VGND.n3702 0.016125
R16251 VGND.n3865 VGND.n3864 0.016125
R16252 VGND.n3707 VGND.n3706 0.016125
R16253 VGND VGND.n637 0.016125
R16254 VGND.n3869 VGND.n3868 0.016125
R16255 VGND.n752 VGND.n749 0.016125
R16256 VGND.n985 VGND.n984 0.016125
R16257 VGND.n3656 VGND.n3655 0.016125
R16258 VGND VGND.n989 0.016125
R16259 VGND.n978 VGND.n977 0.016125
R16260 VGND.n3149 VGND.n3148 0.016125
R16261 VGND.n3328 VGND.n3327 0.016125
R16262 VGND.n3132 VGND.n1106 0.016125
R16263 VGND VGND.n1029 0.016125
R16264 VGND.n3332 VGND.n3331 0.016125
R16265 VGND.n1120 VGND.n1117 0.016125
R16266 VGND.n1265 VGND.n1264 0.016125
R16267 VGND.n3089 VGND.n3088 0.016125
R16268 VGND.n1266 VGND 0.016125
R16269 VGND.n2951 VGND.n2950 0.016125
R16270 VGND.n2551 VGND.n2550 0.016125
R16271 VGND.n2714 VGND.n2713 0.016125
R16272 VGND.n2558 VGND.n2554 0.016125
R16273 VGND VGND.n2701 0.016125
R16274 VGND.n2718 VGND.n2717 0.016125
R16275 VGND.n2116 VGND.n2113 0.016125
R16276 VGND.n2379 VGND.n2378 0.016125
R16277 VGND.n2262 VGND.n2261 0.016125
R16278 VGND.n2239 VGND 0.016125
R16279 VGND VGND.n2366 0.016125
R16280 VGND.n2383 VGND.n2382 0.016125
R16281 VGND.n1816 VGND.n1815 0.016125
R16282 VGND.n2087 VGND.n2086 0.016125
R16283 VGND VGND.n1820 0.016125
R16284 VGND.n1809 VGND.n1642 0.016125
R16285 VGND.n1514 VGND.n1511 0.016125
R16286 VGND.n122 VGND.n121 0.016125
R16287 VGND.n5164 VGND.n5163 0.016125
R16288 VGND.n123 VGND 0.016125
R16289 VGND.n5024 VGND.n5023 0.016125
R16290 VGND.n92 VGND.n89 0.016125
R16291 VGND.n5275 VGND.n5274 0.016125
R16292 VGND.n4302 VGND.n4299 0.016125
R16293 VGND.n4363 VGND.n4362 0.016125
R16294 VGND.n4357 VGND.n4355 0.016125
R16295 VGND.n5271 VGND.n5270 0.016125
R16296 VGND.n5440 VGND.n5439 0.016125
R16297 VGND.n5434 VGND.n5432 0.016125
R16298 VGND.n55 VGND.n54 0.016125
R16299 VGND.n4344 VGND.n4343 0.0148229
R16300 VGND.n4336 VGND.n4335 0.0148229
R16301 VGND.n4880 VGND.n268 0.0148229
R16302 VGND.n4491 VGND.n4490 0.0148229
R16303 VGND.n4544 VGND.n4543 0.0148229
R16304 VGND.n4720 VGND.n4719 0.0148229
R16305 VGND.n4726 VGND.n4725 0.0148229
R16306 VGND.n4858 VGND.n289 0.0148229
R16307 VGND.n4546 VGND.n4545 0.0148229
R16308 VGND.n4718 VGND.n4715 0.0148229
R16309 VGND.n4729 VGND.n299 0.0148229
R16310 VGND.n4857 VGND.n290 0.0148229
R16311 VGND.n4171 VGND.n379 0.0148229
R16312 VGND.n599 VGND.n517 0.0148229
R16313 VGND.n589 VGND.n588 0.0148229
R16314 VGND.n4003 VGND.n514 0.0148229
R16315 VGND.n4170 VGND.n4169 0.0148229
R16316 VGND.n598 VGND.n595 0.0148229
R16317 VGND.n593 VGND.n592 0.0148229
R16318 VGND.n4004 VGND.n506 0.0148229
R16319 VGND.n3704 VGND.n3703 0.0148229
R16320 VGND.n3858 VGND.n3857 0.0148229
R16321 VGND.n3864 VGND.n3863 0.0148229
R16322 VGND.n3983 VGND.n626 0.0148229
R16323 VGND.n3706 VGND.n3705 0.0148229
R16324 VGND.n3856 VGND.n638 0.0148229
R16325 VGND.n3867 VGND.n636 0.0148229
R16326 VGND.n3982 VGND.n627 0.0148229
R16327 VGND.n3658 VGND.n749 0.0148229
R16328 VGND.n994 VGND.n901 0.0148229
R16329 VGND.n984 VGND.n983 0.0148229
R16330 VGND.n3470 VGND.n898 0.0148229
R16331 VGND.n3657 VGND.n3656 0.0148229
R16332 VGND.n993 VGND.n990 0.0148229
R16333 VGND.n988 VGND.n987 0.0148229
R16334 VGND.n3471 VGND.n890 0.0148229
R16335 VGND.n3150 VGND.n3149 0.0148229
R16336 VGND.n3321 VGND.n3320 0.0148229
R16337 VGND.n3327 VGND.n3326 0.0148229
R16338 VGND.n3450 VGND.n1020 0.0148229
R16339 VGND.n3151 VGND.n1106 0.0148229
R16340 VGND.n3319 VGND.n1030 0.0148229
R16341 VGND.n3330 VGND.n1028 0.0148229
R16342 VGND.n3449 VGND.n1021 0.0148229
R16343 VGND.n3091 VGND.n1117 0.0148229
R16344 VGND.n2959 VGND.n2958 0.0148229
R16345 VGND.n1264 VGND.n1263 0.0148229
R16346 VGND.n2847 VGND.n1293 0.0148229
R16347 VGND.n3090 VGND.n3089 0.0148229
R16348 VGND.n2962 VGND.n1259 0.0148229
R16349 VGND.n2952 VGND.n1267 0.0148229
R16350 VGND.n2848 VGND.n1277 0.0148229
R16351 VGND.n2552 VGND.n2551 0.0148229
R16352 VGND.n2707 VGND.n2706 0.0148229
R16353 VGND.n2713 VGND.n2712 0.0148229
R16354 VGND.n2827 VGND.n1319 0.0148229
R16355 VGND.n2554 VGND.n2553 0.0148229
R16356 VGND.n2705 VGND.n2702 0.0148229
R16357 VGND.n2716 VGND.n1334 0.0148229
R16358 VGND.n2826 VGND.n1320 0.0148229
R16359 VGND.n2264 VGND.n2113 0.0148229
R16360 VGND.n2372 VGND.n2371 0.0148229
R16361 VGND.n2378 VGND.n2377 0.0148229
R16362 VGND.n2509 VGND.n1461 0.0148229
R16363 VGND.n2263 VGND.n2262 0.0148229
R16364 VGND.n2370 VGND.n2367 0.0148229
R16365 VGND.n2381 VGND.n1478 0.0148229
R16366 VGND.n1825 VGND.n1752 0.0148229
R16367 VGND.n1815 VGND.n1814 0.0148229
R16368 VGND.n1999 VGND.n1749 0.0148229
R16369 VGND.n2088 VGND.n2087 0.0148229
R16370 VGND.n1824 VGND.n1821 0.0148229
R16371 VGND.n1819 VGND.n1818 0.0148229
R16372 VGND.n2001 VGND.n2000 0.0148229
R16373 VGND.n2089 VGND.n1511 0.0148229
R16374 VGND.n5032 VGND.n5031 0.0148229
R16375 VGND.n121 VGND.n120 0.0148229
R16376 VGND.n1979 VGND.n1851 0.0148229
R16377 VGND.n5165 VGND.n5164 0.0148229
R16378 VGND.n5033 VGND.n116 0.0148229
R16379 VGND.n5025 VGND.n124 0.0148229
R16380 VGND.n1978 VGND.n1864 0.0148229
R16381 VGND.n5166 VGND.n89 0.0148229
R16382 VGND.n5274 VGND.n5273 0.0148229
R16383 VGND.n4299 VGND.n4298 0.0148229
R16384 VGND.n4368 VGND.n4367 0.0148229
R16385 VGND.n4367 VGND 0.0148229
R16386 VGND.n4365 VGND.n4364 0.0148229
R16387 VGND.n4881 VGND.n260 0.0148229
R16388 VGND.n5272 VGND.n5271 0.0148229
R16389 VGND.n5445 VGND.n5444 0.0148229
R16390 VGND.n5444 VGND 0.0148229
R16391 VGND.n5442 VGND.n5441 0.0148229
R16392 VGND.n5457 VGND.n34 0.0148229
R16393 VGND.n5446 VGND.n61 0.0148229
R16394 VGND.n54 VGND.n53 0.0148229
R16395 VGND.n5456 VGND.n42 0.0148229
R16396 VGND.n4745 VGND.n4744 0.014042
R16397 VGND.n581 VGND.n580 0.014042
R16398 VGND.n3883 VGND.n3882 0.014042
R16399 VGND.n976 VGND.n975 0.014042
R16400 VGND.n3346 VGND.n3345 0.014042
R16401 VGND.n2949 VGND.n1268 0.014042
R16402 VGND.n2732 VGND.n2731 0.014042
R16403 VGND.n2405 VGND.n2404 0.014042
R16404 VGND.n2015 VGND.n2014 0.014042
R16405 VGND.n5022 VGND.n125 0.014042
R16406 VGND.n4743 VGND 0.0135208
R16407 VGND.n4737 VGND.n4735 0.0135208
R16408 VGND.n579 VGND 0.0135208
R16409 VGND.n573 VGND.n571 0.0135208
R16410 VGND.n3794 VGND 0.0135208
R16411 VGND.n3881 VGND 0.0135208
R16412 VGND.n3875 VGND.n3873 0.0135208
R16413 VGND.n974 VGND 0.0135208
R16414 VGND.n3344 VGND 0.0135208
R16415 VGND.n3338 VGND.n3336 0.0135208
R16416 VGND VGND.n1279 0.0135208
R16417 VGND.n2730 VGND 0.0135208
R16418 VGND.n2724 VGND.n2722 0.0135208
R16419 VGND.n2403 VGND 0.0135208
R16420 VGND.n2390 VGND.n2388 0.0135208
R16421 VGND.n2013 VGND 0.0135208
R16422 VGND.n2007 VGND.n2005 0.0135208
R16423 VGND VGND.n1852 0.0135208
R16424 VGND.n1861 VGND.n1859 0.0135208
R16425 VGND VGND 0.0135208
R16426 VGND.n4350 VGND.n4348 0.0135208
R16427 VGND.n5427 VGND.n5425 0.0135208
R16428 VGND.n4331 VGND.n4330 0.0130912
R16429 VGND.n4873 VGND.n4872 0.0130912
R16430 VGND.n4186 VGND.n4185 0.0130912
R16431 VGND.n4517 VGND.n4516 0.0130912
R16432 VGND.n275 VGND.n274 0.0130912
R16433 VGND.n4863 VGND.n4862 0.0130912
R16434 VGND.n370 VGND.n369 0.0130912
R16435 VGND.n4176 VGND.n4175 0.0130912
R16436 VGND.n3994 VGND.n3993 0.0130912
R16437 VGND.n605 VGND.n604 0.0130912
R16438 VGND.n3677 VGND.n3676 0.0130912
R16439 VGND.n3687 VGND.n3686 0.0130912
R16440 VGND.n612 VGND.n611 0.0130912
R16441 VGND.n3988 VGND.n3987 0.0130912
R16442 VGND.n740 VGND.n739 0.0130912
R16443 VGND.n3663 VGND.n3662 0.0130912
R16444 VGND.n3461 VGND.n3460 0.0130912
R16445 VGND.n999 VGND.n998 0.0130912
R16446 VGND.n3106 VGND.n3105 0.0130912
R16447 VGND.n3116 VGND.n3115 0.0130912
R16448 VGND.n1006 VGND.n1005 0.0130912
R16449 VGND.n3455 VGND.n3454 0.0130912
R16450 VGND.n1108 VGND.n1107 0.0130912
R16451 VGND.n3096 VGND.n3095 0.0130912
R16452 VGND.n2838 VGND.n2837 0.0130912
R16453 VGND.n1298 VGND.n1297 0.0130912
R16454 VGND.n2525 VGND.n2524 0.0130912
R16455 VGND.n2535 VGND.n2534 0.0130912
R16456 VGND.n1305 VGND.n1304 0.0130912
R16457 VGND.n2832 VGND.n2831 0.0130912
R16458 VGND.n2104 VGND.n2103 0.0130912
R16459 VGND.n1497 VGND.n1496 0.0130912
R16460 VGND.n1455 VGND.n1454 0.0130912
R16461 VGND.n2515 VGND.n2514 0.0130912
R16462 VGND.n1991 VGND.n1990 0.0130912
R16463 VGND.n1832 VGND.n1831 0.0130912
R16464 VGND.n1502 VGND.n1501 0.0130912
R16465 VGND.n2094 VGND.n2093 0.0130912
R16466 VGND.n1838 VGND.n1837 0.0130912
R16467 VGND.n1985 VGND.n1984 0.0130912
R16468 VGND.n5171 VGND.n5170 0.0130912
R16469 VGND.n80 VGND.n79 0.0130912
R16470 VGND.n5195 VGND.n5194 0.0130912
R16471 VGND.n5188 VGND.n5187 0.0130912
R16472 VGND.n4498 VGND.n4497 0.0130912
R16473 VGND.n5450 VGND.n5449 0.0130912
R16474 VGND.n48 VGND.n47 0.0130912
R16475 VGND.n489 VGND.n488 0.0122188
R16476 VGND VGND 0.0122188
R16477 VGND VGND 0.0122188
R16478 VGND.n3138 VGND.n1049 0.0122188
R16479 VGND.n1281 VGND 0.0122188
R16480 VGND.n2508 VGND 0.0122188
R16481 VGND.n216 VGND.n215 0.0122188
R16482 VGND VGND 0.0122188
R16483 VGND VGND 0.0122188
R16484 VGND.n4479 VGND.n4477 0.0122188
R16485 VGND.n4359 VGND.n4358 0.0122188
R16486 VGND.n5264 VGND 0.0122188
R16487 VGND.n5303 VGND.n5302 0.0122188
R16488 VGND.n5436 VGND.n5435 0.0122188
R16489 VGND.n4522 VGND.n4519 0.0111818
R16490 VGND.n4181 VGND.n4178 0.0111818
R16491 VGND.n3692 VGND.n3689 0.0111818
R16492 VGND.n3668 VGND.n3665 0.0111818
R16493 VGND.n3121 VGND.n3118 0.0111818
R16494 VGND.n3101 VGND.n3098 0.0111818
R16495 VGND.n2540 VGND.n2537 0.0111818
R16496 VGND.n2270 VGND.n2269 0.0111818
R16497 VGND.n2099 VGND.n2096 0.0111818
R16498 VGND.n85 VGND.n82 0.0111818
R16499 VGND.n5185 VGND.n5184 0.0111818
R16500 VGND.n4204 VGND.n4203 0.0109167
R16501 VGND.n4530 VGND.n4529 0.0109167
R16502 VGND VGND.n4599 0.0109167
R16503 VGND.n4159 VGND.n4158 0.0109167
R16504 VGND VGND.n4155 0.0109167
R16505 VGND VGND 0.0109167
R16506 VGND.n3718 VGND.n3717 0.0109167
R16507 VGND.n3719 VGND 0.0109167
R16508 VGND.n3643 VGND.n3642 0.0109167
R16509 VGND VGND 0.0109167
R16510 VGND VGND.n3639 0.0109167
R16511 VGND.n3129 VGND.n3128 0.0109167
R16512 VGND VGND.n3209 0.0109167
R16513 VGND VGND 0.0109167
R16514 VGND.n3079 VGND.n3078 0.0109167
R16515 VGND VGND.n3075 0.0109167
R16516 VGND.n2571 VGND.n2570 0.0109167
R16517 VGND VGND.n1342 0.0109167
R16518 VGND.n2249 VGND.n2248 0.0109167
R16519 VGND VGND.n2245 0.0109167
R16520 VGND VGND.n2070 0.0109167
R16521 VGND VGND 0.0109167
R16522 VGND.n2074 VGND.n2073 0.0109167
R16523 VGND VGND.n5147 0.0109167
R16524 VGND VGND 0.0109167
R16525 VGND.n5151 VGND.n5150 0.0109167
R16526 VGND.n5293 VGND.n5292 0.0109167
R16527 VGND.n4471 VGND.n4470 0.0109167
R16528 VGND VGND 0.0109167
R16529 VGND.n5310 VGND.n5309 0.0109167
R16530 VGND.n5445 VGND.n5421 0.00990278
R16531 VGND.n4333 VGND.n4332 0.00975758
R16532 VGND.n4878 VGND.n4877 0.00975758
R16533 VGND.n4526 VGND.n4525 0.00975758
R16534 VGND.n4522 VGND.n4518 0.00975758
R16535 VGND.n272 VGND.n271 0.00975758
R16536 VGND.n281 VGND.n280 0.00975758
R16537 VGND.n378 VGND.n377 0.00975758
R16538 VGND.n4181 VGND.n4177 0.00975758
R16539 VGND.n516 VGND.n515 0.00975758
R16540 VGND.n4001 VGND.n4000 0.00975758
R16541 VGND.n3696 VGND.n3695 0.00975758
R16542 VGND.n3692 VGND.n3688 0.00975758
R16543 VGND.n609 VGND.n608 0.00975758
R16544 VGND.n618 VGND.n617 0.00975758
R16545 VGND.n748 VGND.n747 0.00975758
R16546 VGND.n3668 VGND.n3664 0.00975758
R16547 VGND.n900 VGND.n899 0.00975758
R16548 VGND.n3468 VGND.n3467 0.00975758
R16549 VGND.n3125 VGND.n3124 0.00975758
R16550 VGND.n3121 VGND.n3117 0.00975758
R16551 VGND.n1003 VGND.n1002 0.00975758
R16552 VGND.n1012 VGND.n1011 0.00975758
R16553 VGND.n1116 VGND.n1115 0.00975758
R16554 VGND.n3101 VGND.n3097 0.00975758
R16555 VGND.n1261 VGND.n1260 0.00975758
R16556 VGND.n2845 VGND.n2844 0.00975758
R16557 VGND.n2544 VGND.n2543 0.00975758
R16558 VGND.n2540 VGND.n2536 0.00975758
R16559 VGND.n1302 VGND.n1301 0.00975758
R16560 VGND.n1311 VGND.n1310 0.00975758
R16561 VGND.n2112 VGND.n2111 0.00975758
R16562 VGND.n2270 VGND.n1498 0.00975758
R16563 VGND.n1452 VGND.n1451 0.00975758
R16564 VGND.n1460 VGND.n1459 0.00975758
R16565 VGND.n1751 VGND.n1750 0.00975758
R16566 VGND.n1997 VGND.n1996 0.00975758
R16567 VGND.n1510 VGND.n1509 0.00975758
R16568 VGND.n2099 VGND.n2095 0.00975758
R16569 VGND.n118 VGND.n117 0.00975758
R16570 VGND.n1843 VGND.n1842 0.00975758
R16571 VGND.n88 VGND.n87 0.00975758
R16572 VGND.n85 VGND.n81 0.00975758
R16573 VGND.n5197 VGND.n5196 0.00975758
R16574 VGND.n5186 VGND.n5185 0.00975758
R16575 VGND.n4496 VGND.n4495 0.00975758
R16576 VGND.n4502 VGND.n4499 0.00975758
R16577 VGND.n52 VGND.n51 0.00975758
R16578 VGND.n44 VGND.n43 0.00975758
R16579 VGND.n4735 VGND.n4733 0.00961458
R16580 VGND.n492 VGND.n491 0.00961458
R16581 VGND.n571 VGND.n569 0.00961458
R16582 VGND VGND 0.00961458
R16583 VGND VGND 0.00961458
R16584 VGND VGND 0.00961458
R16585 VGND.n3873 VGND.n3871 0.00961458
R16586 VGND.n3204 VGND.n3202 0.00961458
R16587 VGND.n3336 VGND.n3334 0.00961458
R16588 VGND VGND 0.00961458
R16589 VGND VGND 0.00961458
R16590 VGND.n2722 VGND.n2720 0.00961458
R16591 VGND VGND 0.00961458
R16592 VGND VGND 0.00961458
R16593 VGND.n2388 VGND.n2386 0.00961458
R16594 VGND VGND 0.00961458
R16595 VGND VGND 0.00961458
R16596 VGND.n2005 VGND.n2003 0.00961458
R16597 VGND.n219 VGND.n218 0.00961458
R16598 VGND.n1863 VGND.n1861 0.00961458
R16599 VGND.n4476 VGND.n4474 0.00961458
R16600 VGND.n4348 VGND.n4346 0.00961458
R16601 VGND.n5307 VGND.n5305 0.00961458
R16602 VGND.n5425 VGND.n5423 0.00961458
R16603 VGND.n4340 VGND.n4339 0.0083125
R16604 VGND.n4195 VGND.n4194 0.0083125
R16605 VGND.n4607 VGND.n4606 0.0083125
R16606 VGND.n4724 VGND.n4723 0.0083125
R16607 VGND.n4596 VGND.n304 0.0083125
R16608 VGND.n4744 VGND.n4743 0.0083125
R16609 VGND.n4739 VGND.n4737 0.0083125
R16610 VGND.n4147 VGND.n4146 0.0083125
R16611 VGND.n587 VGND.n586 0.0083125
R16612 VGND.n488 VGND.n486 0.0083125
R16613 VGND.n4152 VGND.n4151 0.0083125
R16614 VGND.n580 VGND.n579 0.0083125
R16615 VGND.n575 VGND.n573 0.0083125
R16616 VGND.n3785 VGND.n3784 0.0083125
R16617 VGND.n3862 VGND.n3861 0.0083125
R16618 VGND.n3723 VGND.n3722 0.0083125
R16619 VGND.n3882 VGND.n3881 0.0083125
R16620 VGND.n3877 VGND.n3875 0.0083125
R16621 VGND.n3631 VGND.n3630 0.0083125
R16622 VGND.n982 VGND.n981 0.0083125
R16623 VGND.n3636 VGND.n3635 0.0083125
R16624 VGND.n975 VGND.n974 0.0083125
R16625 VGND.n3217 VGND.n3216 0.0083125
R16626 VGND.n3325 VGND.n3324 0.0083125
R16627 VGND.n3140 VGND.n3138 0.0083125
R16628 VGND.n3206 VGND.n1047 0.0083125
R16629 VGND.n3345 VGND.n3344 0.0083125
R16630 VGND.n3340 VGND.n3338 0.0083125
R16631 VGND.n3068 VGND.n3067 0.0083125
R16632 VGND.n2955 VGND.n2954 0.0083125
R16633 VGND.n3072 VGND.n3071 0.0083125
R16634 VGND.n1279 VGND.n1268 0.0083125
R16635 VGND VGND.n1277 0.0083125
R16636 VGND.n2632 VGND.n2631 0.0083125
R16637 VGND.n2711 VGND.n2710 0.0083125
R16638 VGND.n2577 VGND.n2575 0.0083125
R16639 VGND.n2731 VGND.n2730 0.0083125
R16640 VGND.n2726 VGND.n2724 0.0083125
R16641 VGND.n2237 VGND.n2236 0.0083125
R16642 VGND.n2376 VGND.n2375 0.0083125
R16643 VGND.n2242 VGND.n2241 0.0083125
R16644 VGND.n2404 VGND.n2403 0.0083125
R16645 VGND.n2392 VGND.n2390 0.0083125
R16646 VGND.n1813 VGND.n1812 0.0083125
R16647 VGND.n2067 VGND.n2066 0.0083125
R16648 VGND.n2014 VGND.n2013 0.0083125
R16649 VGND.n2009 VGND.n2007 0.0083125
R16650 VGND.n2062 VGND.n2061 0.0083125
R16651 VGND.n5028 VGND.n5027 0.0083125
R16652 VGND.n215 VGND.n213 0.0083125
R16653 VGND.n5144 VGND.n5143 0.0083125
R16654 VGND.n1852 VGND.n125 0.0083125
R16655 VGND.n1859 VGND.n1857 0.0083125
R16656 VGND.n5139 VGND.n5138 0.0083125
R16657 VGND.n5284 VGND.n5283 0.0083125
R16658 VGND.n4481 VGND.n4479 0.0083125
R16659 VGND.n4467 VGND.n4466 0.0083125
R16660 VGND.n4358 VGND.n4357 0.0083125
R16661 VGND.n4352 VGND.n4350 0.0083125
R16662 VGND.n5302 VGND.n5300 0.0083125
R16663 VGND.n5315 VGND.n5313 0.0083125
R16664 VGND.n5435 VGND.n5434 0.0083125
R16665 VGND.n5429 VGND.n5427 0.0083125
R16666 VGND.n58 VGND.n57 0.0083125
R16667 VGND.n4339 VGND.n4338 0.00701042
R16668 VGND.n264 VGND.n263 0.00701042
R16669 VGND.n266 VGND.n265 0.00701042
R16670 VGND.n4486 VGND.n4485 0.00701042
R16671 VGND.n4201 VGND.n4200 0.00701042
R16672 VGND.n4194 VGND.n4193 0.00701042
R16673 VGND.n4539 VGND.n4538 0.00701042
R16674 VGND.n4601 VGND.n4600 0.00701042
R16675 VGND.n4608 VGND.n4607 0.00701042
R16676 VGND.n4728 VGND.n4724 0.00701042
R16677 VGND.n285 VGND.n284 0.00701042
R16678 VGND.n287 VGND.n286 0.00701042
R16679 VGND.n4609 VGND.n304 0.00701042
R16680 VGND.n386 VGND.n385 0.00701042
R16681 VGND.n4156 VGND.n387 0.00701042
R16682 VGND.n4148 VGND.n4147 0.00701042
R16683 VGND.n591 VGND.n587 0.00701042
R16684 VGND.n510 VGND.n509 0.00701042
R16685 VGND.n512 VGND.n511 0.00701042
R16686 VGND.n4151 VGND.n4149 0.00701042
R16687 VGND.n3699 VGND.n647 0.00701042
R16688 VGND.n3791 VGND.n3790 0.00701042
R16689 VGND.n3784 VGND.n3783 0.00701042
R16690 VGND.n3866 VGND.n3862 0.00701042
R16691 VGND.n622 VGND.n621 0.00701042
R16692 VGND.n624 VGND.n623 0.00701042
R16693 VGND VGND.n3793 0.00701042
R16694 VGND.n3782 VGND.n3723 0.00701042
R16695 VGND.n3781 VGND 0.00701042
R16696 VGND.n756 VGND.n755 0.00701042
R16697 VGND.n3640 VGND.n757 0.00701042
R16698 VGND.n3632 VGND.n3631 0.00701042
R16699 VGND.n986 VGND.n982 0.00701042
R16700 VGND.n894 VGND.n893 0.00701042
R16701 VGND.n896 VGND.n895 0.00701042
R16702 VGND.n3635 VGND.n3633 0.00701042
R16703 VGND.n3145 VGND.n3144 0.00701042
R16704 VGND.n3211 VGND.n3210 0.00701042
R16705 VGND.n3218 VGND.n3217 0.00701042
R16706 VGND.n3329 VGND.n3325 0.00701042
R16707 VGND.n1016 VGND.n1015 0.00701042
R16708 VGND.n1018 VGND.n1017 0.00701042
R16709 VGND.n3219 VGND.n1047 0.00701042
R16710 VGND.n1124 VGND.n1123 0.00701042
R16711 VGND.n3076 VGND.n1125 0.00701042
R16712 VGND.n3069 VGND.n3068 0.00701042
R16713 VGND.n2954 VGND.n2953 0.00701042
R16714 VGND.n1289 VGND.n1288 0.00701042
R16715 VGND.n1291 VGND.n1290 0.00701042
R16716 VGND.n3071 VGND.n3070 0.00701042
R16717 VGND.n2547 VGND.n1343 0.00701042
R16718 VGND.n2638 VGND.n2637 0.00701042
R16719 VGND.n2631 VGND.n2630 0.00701042
R16720 VGND.n2715 VGND.n2711 0.00701042
R16721 VGND.n1315 VGND.n1314 0.00701042
R16722 VGND.n1317 VGND.n1316 0.00701042
R16723 VGND.n2629 VGND.n2577 0.00701042
R16724 VGND.n2120 VGND.n2119 0.00701042
R16725 VGND.n2246 VGND.n2121 0.00701042
R16726 VGND.n2238 VGND.n2237 0.00701042
R16727 VGND.n2380 VGND.n2376 0.00701042
R16728 VGND.n2399 VGND.n2398 0.00701042
R16729 VGND.n2397 VGND.n2396 0.00701042
R16730 VGND.n2241 VGND.n2239 0.00701042
R16731 VGND.n1817 VGND.n1813 0.00701042
R16732 VGND.n1745 VGND.n1744 0.00701042
R16733 VGND.n1747 VGND.n1746 0.00701042
R16734 VGND.n2066 VGND.n2064 0.00701042
R16735 VGND.n1518 VGND.n1517 0.00701042
R16736 VGND.n2071 VGND.n1519 0.00701042
R16737 VGND.n2063 VGND.n2062 0.00701042
R16738 VGND.n5027 VGND.n5026 0.00701042
R16739 VGND.n1847 VGND.n1846 0.00701042
R16740 VGND.n1849 VGND.n1848 0.00701042
R16741 VGND.n5143 VGND.n5141 0.00701042
R16742 VGND.n96 VGND.n95 0.00701042
R16743 VGND.n5148 VGND.n97 0.00701042
R16744 VGND.n5140 VGND.n5139 0.00701042
R16745 VGND.n5279 VGND.n5278 0.00701042
R16746 VGND.n5290 VGND.n5289 0.00701042
R16747 VGND.n5283 VGND.n5282 0.00701042
R16748 VGND.n4466 VGND.n4463 0.00701042
R16749 VGND.n5316 VGND.n5315 0.00701042
R16750 VGND.n57 VGND.n56 0.00701042
R16751 VGND.n38 VGND.n37 0.00701042
R16752 VGND.n40 VGND.n39 0.00701042
R16753 VGND.n1245 VGND.n1244 0.00693178
R16754 VGND.n2229 VGND.n2228 0.00693178
R16755 VGND.n1638 VGND.n1637 0.00693178
R16756 VGND.n4593 VGND.n4592 0.00693178
R16757 VGND.n3796 VGND.n3795 0.00693178
R16758 VGND.n881 VGND.n880 0.00693178
R16759 VGND.n2642 VGND.n2641 0.00693178
R16760 VGND VGND.n4366 0.00570833
R16761 VGND VGND.n5443 0.00570833
R16762 VGND.n4594 VGND.n4593 0.00548035
R16763 VGND.n3795 VGND.n3794 0.00548035
R16764 VGND.n880 VGND.n879 0.00548035
R16765 VGND.n1244 VGND.n1243 0.00548035
R16766 VGND.n2641 VGND.n2640 0.00548035
R16767 VGND.n2230 VGND.n2229 0.00548035
R16768 VGND.n1637 VGND.n1636 0.00548035
R16769 VGND.n4591 VGND.n306 0.00484057
R16770 VGND.n3797 VGND.n646 0.00484057
R16771 VGND.n882 VGND.n878 0.00484057
R16772 VGND.n1246 VGND.n1242 0.00484057
R16773 VGND.n2643 VGND.n1341 0.00484057
R16774 VGND.n2227 VGND.n2122 0.00484057
R16775 VGND.n1639 VGND.n1635 0.00484057
R16776 VGND.n5182 VGND.n5181 0.00460158
R16777 VGND.n5178 VGND.n5177 0.00460158
R16778 VGND.n1508 VGND.n1500 0.00460158
R16779 VGND.n2110 VGND.n2102 0.00460158
R16780 VGND.n2531 VGND.n2523 0.00460158
R16781 VGND.n2532 VGND.n1114 0.00460158
R16782 VGND.n3112 VGND.n3104 0.00460158
R16783 VGND.n3113 VGND.n746 0.00460158
R16784 VGND.n3683 VGND.n3675 0.00460158
R16785 VGND.n3684 VGND.n376 0.00460158
R16786 VGND.n4192 VGND.n4184 0.00460158
R16787 VGND.n1841 VGND.n1836 0.00460158
R16788 VGND.n1994 VGND.n1989 0.00460158
R16789 VGND.n1827 VGND.n1458 0.00460158
R16790 VGND.n2519 VGND.n1309 0.00460158
R16791 VGND.n2842 VGND.n2836 0.00460158
R16792 VGND.n1294 VGND.n1010 0.00460158
R16793 VGND.n3465 VGND.n3459 0.00460158
R16794 VGND.n3671 VGND.n616 0.00460158
R16795 VGND.n3998 VGND.n3992 0.00460158
R16796 VGND.n601 VGND.n279 0.00460158
R16797 VGND.n4875 VGND.n4867 0.00460158
R16798 VGND.n5453 VGND.n5448 0.00460158
R16799 VGND.n4503 VGND.n4502 0.0045458
R16800 VGND.n4338 VGND.n4337 0.00440625
R16801 VGND.n263 VGND.n262 0.00440625
R16802 VGND.n4492 VGND.n4491 0.00440625
R16803 VGND.n4489 VGND.n4488 0.00440625
R16804 VGND.n4485 VGND.n4484 0.00440625
R16805 VGND.n4206 VGND.n4205 0.00440625
R16806 VGND.n4202 VGND.n4201 0.00440625
R16807 VGND.n4200 VGND.n4199 0.00440625
R16808 VGND.n4197 VGND.n4196 0.00440625
R16809 VGND.n4544 VGND.n4528 0.00440625
R16810 VGND.n4542 VGND.n4541 0.00440625
R16811 VGND.n4538 VGND.n4537 0.00440625
R16812 VGND.n4532 VGND.n4531 0.00440625
R16813 VGND.n4600 VGND.n305 0.00440625
R16814 VGND.n4602 VGND.n4601 0.00440625
R16815 VGND.n4605 VGND.n4604 0.00440625
R16816 VGND.n4728 VGND.n4727 0.00440625
R16817 VGND.n284 VGND.n283 0.00440625
R16818 VGND.n4545 VGND.n368 0.00440625
R16819 VGND.n4536 VGND.n4534 0.00440625
R16820 VGND.n4535 VGND.n306 0.00440625
R16821 VGND VGND.n4595 0.00440625
R16822 VGND.n4598 VGND.n4597 0.00440625
R16823 VGND.n4718 VGND.n4713 0.00440625
R16824 VGND.n4715 VGND 0.00440625
R16825 VGND.n4730 VGND.n4729 0.00440625
R16826 VGND.n4741 VGND.n4740 0.00440625
R16827 VGND.n4172 VGND.n4171 0.00440625
R16828 VGND.n383 VGND.n382 0.00440625
R16829 VGND.n4162 VGND.n386 0.00440625
R16830 VGND.n4161 VGND.n4160 0.00440625
R16831 VGND.n4157 VGND.n4156 0.00440625
R16832 VGND.n4142 VGND.n387 0.00440625
R16833 VGND.n4145 VGND.n4144 0.00440625
R16834 VGND.n591 VGND.n590 0.00440625
R16835 VGND.n509 VGND.n508 0.00440625
R16836 VGND.n4170 VGND.n380 0.00440625
R16837 VGND.n4164 VGND.n4163 0.00440625
R16838 VGND.n486 VGND.n381 0.00440625
R16839 VGND VGND.n388 0.00440625
R16840 VGND.n4154 VGND.n4153 0.00440625
R16841 VGND.n598 VGND.n567 0.00440625
R16842 VGND.n595 VGND 0.00440625
R16843 VGND.n592 VGND.n583 0.00440625
R16844 VGND.n577 VGND.n576 0.00440625
R16845 VGND.n3704 VGND.n3698 0.00440625
R16846 VGND.n3702 VGND.n3701 0.00440625
R16847 VGND.n3714 VGND.n647 0.00440625
R16848 VGND.n3716 VGND.n3715 0.00440625
R16849 VGND.n3792 VGND.n3791 0.00440625
R16850 VGND.n3790 VGND.n3789 0.00440625
R16851 VGND.n3787 VGND.n3786 0.00440625
R16852 VGND.n3866 VGND.n3865 0.00440625
R16853 VGND.n621 VGND.n620 0.00440625
R16854 VGND.n3705 VGND.n738 0.00440625
R16855 VGND.n3713 VGND.n3711 0.00440625
R16856 VGND.n3712 VGND.n646 0.00440625
R16857 VGND.n3793 VGND 0.00440625
R16858 VGND.n3721 VGND.n3720 0.00440625
R16859 VGND.n638 VGND 0.00440625
R16860 VGND.n3868 VGND.n3867 0.00440625
R16861 VGND.n3879 VGND.n3878 0.00440625
R16862 VGND.n3659 VGND.n3658 0.00440625
R16863 VGND.n753 VGND.n752 0.00440625
R16864 VGND.n3646 VGND.n756 0.00440625
R16865 VGND.n3645 VGND.n3644 0.00440625
R16866 VGND.n3641 VGND.n3640 0.00440625
R16867 VGND.n3626 VGND.n757 0.00440625
R16868 VGND.n3629 VGND.n3628 0.00440625
R16869 VGND.n986 VGND.n985 0.00440625
R16870 VGND.n893 VGND.n892 0.00440625
R16871 VGND.n3657 VGND.n750 0.00440625
R16872 VGND.n3648 VGND.n3647 0.00440625
R16873 VGND.n878 VGND.n751 0.00440625
R16874 VGND VGND.n758 0.00440625
R16875 VGND.n3638 VGND.n3637 0.00440625
R16876 VGND.n993 VGND.n965 0.00440625
R16877 VGND.n987 VGND.n978 0.00440625
R16878 VGND.n972 VGND.n971 0.00440625
R16879 VGND.n3150 VGND.n3127 0.00440625
R16880 VGND.n3148 VGND.n3147 0.00440625
R16881 VGND.n3144 VGND.n3143 0.00440625
R16882 VGND.n3131 VGND.n3130 0.00440625
R16883 VGND.n3210 VGND.n1048 0.00440625
R16884 VGND.n3212 VGND.n3211 0.00440625
R16885 VGND.n3215 VGND.n3214 0.00440625
R16886 VGND.n3329 VGND.n3328 0.00440625
R16887 VGND.n1015 VGND.n1014 0.00440625
R16888 VGND.n3152 VGND.n3151 0.00440625
R16889 VGND.n3142 VGND.n3136 0.00440625
R16890 VGND.n3141 VGND.n3140 0.00440625
R16891 VGND VGND.n3205 0.00440625
R16892 VGND.n3208 VGND.n3207 0.00440625
R16893 VGND.n1030 VGND 0.00440625
R16894 VGND.n3331 VGND.n3330 0.00440625
R16895 VGND.n3342 VGND.n3341 0.00440625
R16896 VGND.n3092 VGND.n3091 0.00440625
R16897 VGND.n1121 VGND.n1120 0.00440625
R16898 VGND.n3082 VGND.n1124 0.00440625
R16899 VGND.n3081 VGND.n3080 0.00440625
R16900 VGND.n3077 VGND.n3076 0.00440625
R16901 VGND.n3063 VGND.n1125 0.00440625
R16902 VGND.n3066 VGND.n3065 0.00440625
R16903 VGND.n2953 VGND.n1265 0.00440625
R16904 VGND.n1288 VGND.n1287 0.00440625
R16905 VGND.n3090 VGND.n1118 0.00440625
R16906 VGND.n3084 VGND.n3083 0.00440625
R16907 VGND.n1242 VGND.n1119 0.00440625
R16908 VGND VGND.n1126 0.00440625
R16909 VGND.n3074 VGND.n3073 0.00440625
R16910 VGND.n2963 VGND.n2962 0.00440625
R16911 VGND VGND.n1259 0.00440625
R16912 VGND.n2952 VGND.n2951 0.00440625
R16913 VGND.n1286 VGND.n1285 0.00440625
R16914 VGND.n2552 VGND.n2546 0.00440625
R16915 VGND.n2550 VGND.n2549 0.00440625
R16916 VGND.n2567 VGND.n1343 0.00440625
R16917 VGND.n2569 VGND.n2568 0.00440625
R16918 VGND.n2638 VGND.n2572 0.00440625
R16919 VGND.n2637 VGND.n2636 0.00440625
R16920 VGND.n2634 VGND.n2633 0.00440625
R16921 VGND.n2715 VGND.n2714 0.00440625
R16922 VGND.n1314 VGND.n1313 0.00440625
R16923 VGND.n2553 VGND.n1449 0.00440625
R16924 VGND.n2566 VGND.n2564 0.00440625
R16925 VGND.n2565 VGND.n1341 0.00440625
R16926 VGND.n2639 VGND 0.00440625
R16927 VGND.n2574 VGND.n2573 0.00440625
R16928 VGND.n2705 VGND.n2700 0.00440625
R16929 VGND.n2702 VGND 0.00440625
R16930 VGND.n2717 VGND.n2716 0.00440625
R16931 VGND.n2728 VGND.n2727 0.00440625
R16932 VGND.n2265 VGND.n2264 0.00440625
R16933 VGND.n2117 VGND.n2116 0.00440625
R16934 VGND.n2252 VGND.n2120 0.00440625
R16935 VGND.n2251 VGND.n2250 0.00440625
R16936 VGND.n2247 VGND.n2246 0.00440625
R16937 VGND.n2232 VGND.n2121 0.00440625
R16938 VGND.n2235 VGND.n2234 0.00440625
R16939 VGND.n2380 VGND.n2379 0.00440625
R16940 VGND.n2400 VGND.n2399 0.00440625
R16941 VGND.n2263 VGND.n2114 0.00440625
R16942 VGND.n2254 VGND.n2253 0.00440625
R16943 VGND.n2122 VGND.n2115 0.00440625
R16944 VGND VGND.n2231 0.00440625
R16945 VGND.n2244 VGND.n2243 0.00440625
R16946 VGND.n2370 VGND.n2365 0.00440625
R16947 VGND.n2367 VGND 0.00440625
R16948 VGND.n2382 VGND.n2381 0.00440625
R16949 VGND.n2401 VGND.n2393 0.00440625
R16950 VGND.n1817 VGND.n1816 0.00440625
R16951 VGND.n1744 VGND.n1743 0.00440625
R16952 VGND.n2088 VGND.n1512 0.00440625
R16953 VGND.n2079 VGND.n2078 0.00440625
R16954 VGND.n1635 VGND.n1513 0.00440625
R16955 VGND VGND.n1520 0.00440625
R16956 VGND.n2069 VGND.n2068 0.00440625
R16957 VGND.n1824 VGND.n1808 0.00440625
R16958 VGND.n1821 VGND 0.00440625
R16959 VGND.n1818 VGND.n1809 0.00440625
R16960 VGND.n2011 VGND.n2010 0.00440625
R16961 VGND.n2090 VGND.n2089 0.00440625
R16962 VGND.n1515 VGND.n1514 0.00440625
R16963 VGND.n2077 VGND.n1518 0.00440625
R16964 VGND.n2076 VGND.n2075 0.00440625
R16965 VGND.n2072 VGND.n2071 0.00440625
R16966 VGND.n2057 VGND.n1519 0.00440625
R16967 VGND.n2060 VGND.n2059 0.00440625
R16968 VGND.n5026 VGND.n122 0.00440625
R16969 VGND.n1846 VGND.n1845 0.00440625
R16970 VGND.n5165 VGND.n90 0.00440625
R16971 VGND.n5156 VGND.n5155 0.00440625
R16972 VGND.n213 VGND.n91 0.00440625
R16973 VGND VGND.n98 0.00440625
R16974 VGND.n5146 VGND.n5145 0.00440625
R16975 VGND.n5034 VGND.n5033 0.00440625
R16976 VGND VGND.n116 0.00440625
R16977 VGND.n5025 VGND.n5024 0.00440625
R16978 VGND.n1855 VGND.n1854 0.00440625
R16979 VGND.n5167 VGND.n5166 0.00440625
R16980 VGND.n93 VGND.n92 0.00440625
R16981 VGND.n5154 VGND.n96 0.00440625
R16982 VGND.n5153 VGND.n5152 0.00440625
R16983 VGND.n5149 VGND.n5148 0.00440625
R16984 VGND.n5134 VGND.n97 0.00440625
R16985 VGND.n5137 VGND.n5136 0.00440625
R16986 VGND.n5273 VGND.n5199 0.00440625
R16987 VGND.n5276 VGND.n5275 0.00440625
R16988 VGND.n5296 VGND.n5279 0.00440625
R16989 VGND.n5295 VGND.n5294 0.00440625
R16990 VGND.n5291 VGND.n5290 0.00440625
R16991 VGND.n5289 VGND.n5288 0.00440625
R16992 VGND.n5286 VGND.n5285 0.00440625
R16993 VGND.n4298 VGND.n4297 0.00440625
R16994 VGND.n4483 VGND.n4307 0.00440625
R16995 VGND.n4482 VGND.n4481 0.00440625
R16996 VGND.n4472 VGND.n4471 0.00440625
R16997 VGND.n4469 VGND.n4468 0.00440625
R16998 VGND.n4369 VGND.n4368 0.00440625
R16999 VGND.n4364 VGND.n4363 0.00440625
R17000 VGND.n4354 VGND.n4353 0.00440625
R17001 VGND.n5272 VGND.n5263 0.00440625
R17002 VGND.n5297 VGND.n78 0.00440625
R17003 VGND.n5300 VGND.n5298 0.00440625
R17004 VGND.n5309 VGND.n5308 0.00440625
R17005 VGND.n5312 VGND.n5311 0.00440625
R17006 VGND.n5441 VGND.n5440 0.00440625
R17007 VGND.n5431 VGND.n5430 0.00440625
R17008 VGND.n56 VGND.n55 0.00440625
R17009 VGND.n37 VGND.n36 0.00440625
R17010 VGND.n4869 VGND.n4868 0.00406061
R17011 VGND.n4874 VGND.n4871 0.00406061
R17012 VGND.n4191 VGND.n4190 0.00406061
R17013 VGND.n4188 VGND.n4187 0.00406061
R17014 VGND.n278 VGND.n277 0.00406061
R17015 VGND.n4864 VGND.n4861 0.00406061
R17016 VGND.n375 VGND.n374 0.00406061
R17017 VGND.n372 VGND.n371 0.00406061
R17018 VGND.n3997 VGND.n3996 0.00406061
R17019 VGND.n606 VGND.n603 0.00406061
R17020 VGND.n3682 VGND.n3681 0.00406061
R17021 VGND.n3679 VGND.n3678 0.00406061
R17022 VGND.n615 VGND.n614 0.00406061
R17023 VGND.n3989 VGND.n3986 0.00406061
R17024 VGND.n745 VGND.n744 0.00406061
R17025 VGND.n742 VGND.n741 0.00406061
R17026 VGND.n3464 VGND.n3463 0.00406061
R17027 VGND.n1000 VGND.n997 0.00406061
R17028 VGND.n3111 VGND.n3110 0.00406061
R17029 VGND.n3108 VGND.n3107 0.00406061
R17030 VGND.n1009 VGND.n1008 0.00406061
R17031 VGND.n3456 VGND.n3453 0.00406061
R17032 VGND.n1113 VGND.n1112 0.00406061
R17033 VGND.n1110 VGND.n1109 0.00406061
R17034 VGND.n2841 VGND.n2840 0.00406061
R17035 VGND.n1299 VGND.n1296 0.00406061
R17036 VGND.n2530 VGND.n2529 0.00406061
R17037 VGND.n2527 VGND.n2526 0.00406061
R17038 VGND.n1308 VGND.n1307 0.00406061
R17039 VGND.n2833 VGND.n2830 0.00406061
R17040 VGND.n2109 VGND.n2108 0.00406061
R17041 VGND.n2106 VGND.n2105 0.00406061
R17042 VGND.n1457 VGND.n1456 0.00406061
R17043 VGND.n2516 VGND.n2513 0.00406061
R17044 VGND.n1993 VGND.n1992 0.00406061
R17045 VGND.n1833 VGND.n1830 0.00406061
R17046 VGND.n1507 VGND.n1506 0.00406061
R17047 VGND.n1504 VGND.n1503 0.00406061
R17048 VGND.n1840 VGND.n1839 0.00406061
R17049 VGND.n1986 VGND.n1983 0.00406061
R17050 VGND.n5176 VGND.n5175 0.00406061
R17051 VGND.n5173 VGND.n5172 0.00406061
R17052 VGND.n5193 VGND.n5192 0.00406061
R17053 VGND.n5190 VGND.n5189 0.00406061
R17054 VGND.n4509 VGND.n4508 0.00406061
R17055 VGND.n4506 VGND.n4505 0.00406061
R17056 VGND.n5452 VGND.n5451 0.00406061
R17057 VGND.n49 VGND.n46 0.00406061
R17058 VGND.n1499 VGND.n86 0.00393497
R17059 VGND.n2101 VGND.n2100 0.00393497
R17060 VGND.n2268 VGND.n1450 0.00393497
R17061 VGND.n2541 VGND.n2533 0.00393497
R17062 VGND.n3103 VGND.n3102 0.00393497
R17063 VGND.n3122 VGND.n3114 0.00393497
R17064 VGND.n3670 VGND.n3669 0.00393497
R17065 VGND.n3693 VGND.n3685 0.00393497
R17066 VGND.n4183 VGND.n4182 0.00393497
R17067 VGND.n4523 VGND.n4515 0.00393497
R17068 VGND.n4511 VGND.n4510 0.00393497
R17069 VGND.n5180 VGND.n5179 0.00393497
R17070 VGND.n4514 VGND.n4513 0.00393497
R17071 VGND.n1835 VGND.n50 0.00393497
R17072 VGND.n270 VGND.n269 0.00393497
R17073 VGND.n4866 VGND.n4865 0.00393497
R17074 VGND.n607 VGND.n602 0.00393497
R17075 VGND.n3991 VGND.n3990 0.00393497
R17076 VGND.n1001 VGND.n996 0.00393497
R17077 VGND.n3458 VGND.n3457 0.00393497
R17078 VGND.n1300 VGND.n1295 0.00393497
R17079 VGND.n2835 VGND.n2834 0.00393497
R17080 VGND.n2518 VGND.n2517 0.00393497
R17081 VGND.n1834 VGND.n1828 0.00393497
R17082 VGND.n1988 VGND.n1987 0.00393497
R17083 VGND.n4496 VGND.n4493 0.00365283
R17084 VGND.n4334 VGND.n4333 0.00365283
R17085 VGND.n4167 VGND.n4166 0.00362532
R17086 VGND.n4548 VGND.n367 0.00362532
R17087 VGND.n3709 VGND.n3708 0.00362532
R17088 VGND.n2260 VGND.n2256 0.00362532
R17089 VGND VGND.n4533 0.00310417
R17090 VGND VGND.n4742 0.00310417
R17091 VGND.n4165 VGND 0.00310417
R17092 VGND VGND.n578 0.00310417
R17093 VGND VGND.n3710 0.00310417
R17094 VGND VGND.n3880 0.00310417
R17095 VGND.n3655 VGND.n3652 0.00310417
R17096 VGND.n3650 VGND 0.00310417
R17097 VGND.n990 VGND 0.00310417
R17098 VGND VGND.n973 0.00310417
R17099 VGND.n3133 VGND.n3132 0.00310417
R17100 VGND VGND.n3135 0.00310417
R17101 VGND VGND.n3343 0.00310417
R17102 VGND.n3088 VGND.n3087 0.00310417
R17103 VGND.n3085 VGND 0.00310417
R17104 VGND.n1280 VGND 0.00310417
R17105 VGND.n2559 VGND.n2558 0.00310417
R17106 VGND VGND.n2563 0.00310417
R17107 VGND VGND.n2729 0.00310417
R17108 VGND.n2255 VGND 0.00310417
R17109 VGND.n2273 VGND 0.00310417
R17110 VGND VGND.n2402 0.00310417
R17111 VGND.n2384 VGND 0.00310417
R17112 VGND.n2086 VGND.n2083 0.00310417
R17113 VGND.n2081 VGND 0.00310417
R17114 VGND VGND.n2012 0.00310417
R17115 VGND VGND 0.00310417
R17116 VGND.n5163 VGND.n5160 0.00310417
R17117 VGND.n5158 VGND 0.00310417
R17118 VGND.n1853 VGND 0.00310417
R17119 VGND.n4303 VGND.n4302 0.00310417
R17120 VGND.n4362 VGND.n4359 0.00310417
R17121 VGND.n5270 VGND.n5266 0.00310417
R17122 VGND.n5439 VGND.n5436 0.00310417
R17123 VGND.n5177 VGND.n5169 0.0028004
R17124 VGND.n2092 VGND.n1508 0.0028004
R17125 VGND.n2267 VGND.n2110 0.0028004
R17126 VGND.n2542 VGND.n2531 0.0028004
R17127 VGND.n3094 VGND.n1114 0.0028004
R17128 VGND.n3123 VGND.n3112 0.0028004
R17129 VGND.n3661 VGND.n746 0.0028004
R17130 VGND.n3694 VGND.n3683 0.0028004
R17131 VGND.n4174 VGND.n376 0.0028004
R17132 VGND.n4524 VGND.n4192 0.0028004
R17133 VGND.n5183 VGND.n5182 0.0028004
R17134 VGND.n4860 VGND.n279 0.0028004
R17135 VGND.n3999 VGND.n3998 0.0028004
R17136 VGND.n3985 VGND.n616 0.0028004
R17137 VGND.n3466 VGND.n3465 0.0028004
R17138 VGND.n3452 VGND.n1010 0.0028004
R17139 VGND.n2843 VGND.n2842 0.0028004
R17140 VGND.n2829 VGND.n1309 0.0028004
R17141 VGND.n2511 VGND.n1458 0.0028004
R17142 VGND.n1995 VGND.n1994 0.0028004
R17143 VGND.n1981 VGND.n1841 0.0028004
R17144 VGND.n4876 VGND.n4875 0.0028004
R17145 VGND.n5454 VGND.n5453 0.0028004
R17146 VGND.n5455 VGND.n44 0.00271013
R17147 VGND.n5183 VGND.n5180 0.00246749
R17148 VGND.n4513 VGND.n4512 0.00246749
R17149 VGND.n5169 VGND.n86 0.00246749
R17150 VGND.n2100 VGND.n2092 0.00246749
R17151 VGND.n2268 VGND.n2267 0.00246749
R17152 VGND.n2542 VGND.n2541 0.00246749
R17153 VGND.n3102 VGND.n3094 0.00246749
R17154 VGND.n3123 VGND.n3122 0.00246749
R17155 VGND.n3669 VGND.n3661 0.00246749
R17156 VGND.n3694 VGND.n3693 0.00246749
R17157 VGND.n4182 VGND.n4174 0.00246749
R17158 VGND.n4524 VGND.n4523 0.00246749
R17159 VGND.n4512 VGND.n4511 0.00246749
R17160 VGND.n5454 VGND.n50 0.00246749
R17161 VGND.n1987 VGND.n1981 0.00246749
R17162 VGND.n1995 VGND.n1834 0.00246749
R17163 VGND.n2517 VGND.n2511 0.00246749
R17164 VGND.n2834 VGND.n2829 0.00246749
R17165 VGND.n2843 VGND.n1300 0.00246749
R17166 VGND.n3457 VGND.n3452 0.00246749
R17167 VGND.n3466 VGND.n1001 0.00246749
R17168 VGND.n3990 VGND.n3985 0.00246749
R17169 VGND.n3999 VGND.n607 0.00246749
R17170 VGND.n4865 VGND.n4860 0.00246749
R17171 VGND.n4876 VGND.n270 0.00246749
R17172 VGND.n4859 VGND.n281 0.00237907
R17173 VGND.n4002 VGND.n4001 0.00237907
R17174 VGND.n3984 VGND.n618 0.00237907
R17175 VGND.n3469 VGND.n3468 0.00237907
R17176 VGND.n3451 VGND.n1012 0.00237907
R17177 VGND.n2846 VGND.n2845 0.00237907
R17178 VGND.n2828 VGND.n1311 0.00237907
R17179 VGND.n2510 VGND.n1460 0.00237907
R17180 VGND.n1998 VGND.n1997 0.00237907
R17181 VGND.n1980 VGND.n1843 0.00237907
R17182 VGND.n4879 VGND.n4878 0.00237907
R17183 VGND.n4527 VGND.n4526 0.00233584
R17184 VGND.n273 VGND.n272 0.00233584
R17185 VGND.n4173 VGND.n378 0.00233584
R17186 VGND.n600 VGND.n516 0.00233584
R17187 VGND.n3697 VGND.n3696 0.00233584
R17188 VGND.n610 VGND.n609 0.00233584
R17189 VGND.n3660 VGND.n748 0.00233584
R17190 VGND.n995 VGND.n900 0.00233584
R17191 VGND.n3126 VGND.n3125 0.00233584
R17192 VGND.n1004 VGND.n1003 0.00233584
R17193 VGND.n3093 VGND.n1116 0.00233584
R17194 VGND.n1262 VGND.n1261 0.00233584
R17195 VGND.n2545 VGND.n2544 0.00233584
R17196 VGND.n1303 VGND.n1302 0.00233584
R17197 VGND.n2266 VGND.n2112 0.00233584
R17198 VGND.n1453 VGND.n1452 0.00233584
R17199 VGND.n1826 VGND.n1751 0.00233584
R17200 VGND.n2091 VGND.n1510 0.00233584
R17201 VGND.n119 VGND.n118 0.00233584
R17202 VGND.n5168 VGND.n88 0.00233584
R17203 VGND.n5198 VGND.n5197 0.00233584
R17204 VGND.n5447 VGND.n52 0.00233584
R17205 VGND.n4745 VGND.n4731 0.00228056
R17206 VGND.n582 VGND.n581 0.00228056
R17207 VGND.n4168 VGND.n4167 0.00228056
R17208 VGND.n3883 VGND.n3869 0.00228056
R17209 VGND.n977 VGND.n976 0.00228056
R17210 VGND.n3346 VGND.n3332 0.00228056
R17211 VGND.n2950 VGND.n2949 0.00228056
R17212 VGND.n2732 VGND.n2718 0.00228056
R17213 VGND.n2405 VGND.n2383 0.00228056
R17214 VGND.n2015 VGND.n1642 0.00228056
R17215 VGND.n5023 VGND.n5022 0.00228056
R17216 VGND.n4548 VGND.n4547 0.00228056
R17217 VGND.n3708 VGND.n3707 0.00228056
R17218 VGND.n2261 VGND.n2260 0.00228056
R17219 VGND.n4501 VGND.n4500 0.00180208
R17220 VGND.n4521 VGND.n4520 0.00180208
R17221 VGND.n4180 VGND.n4179 0.00180208
R17222 VGND VGND 0.00180208
R17223 VGND.n492 VGND.n489 0.00180208
R17224 VGND.n3691 VGND.n3690 0.00180208
R17225 VGND VGND 0.00180208
R17226 VGND VGND 0.00180208
R17227 VGND.n3667 VGND.n3666 0.00180208
R17228 VGND VGND 0.00180208
R17229 VGND.n3652 VGND.n3651 0.00180208
R17230 VGND VGND 0.00180208
R17231 VGND.n3120 VGND.n3119 0.00180208
R17232 VGND.n3134 VGND.n3133 0.00180208
R17233 VGND.n3202 VGND.n1049 0.00180208
R17234 VGND VGND 0.00180208
R17235 VGND.n3100 VGND.n3099 0.00180208
R17236 VGND.n3087 VGND.n3086 0.00180208
R17237 VGND VGND 0.00180208
R17238 VGND.n2539 VGND.n2538 0.00180208
R17239 VGND.n2560 VGND.n2559 0.00180208
R17240 VGND VGND 0.00180208
R17241 VGND.n2272 VGND.n2271 0.00180208
R17242 VGND VGND 0.00180208
R17243 VGND.n2083 VGND.n2082 0.00180208
R17244 VGND.n2098 VGND.n2097 0.00180208
R17245 VGND.n5160 VGND.n5159 0.00180208
R17246 VGND.n219 VGND.n216 0.00180208
R17247 VGND.n84 VGND.n83 0.00180208
R17248 VGND.n5281 VGND.n5280 0.00180208
R17249 VGND.n4304 VGND.n4303 0.00180208
R17250 VGND.n4477 VGND.n4476 0.00180208
R17251 VGND.n5266 VGND.n5265 0.00180208
R17252 VGND.n5305 VGND.n5303 0.00180208
R17253 ctlp[6] ctlp[6] 13.2956
R17254 ctln[1].n0 ctln[1] 15.6555
R17255 ctln[1].n0 ctln[1] 9.6005
R17256 ctln[1] ctln[1].n0 3.2005
R17257 trim[0].n0 trim[0] 9.6005
R17258 trim[0].n0 trim[0] 6.81829
R17259 trim[0] trim[0].n0 3.2005
R17260 ctlp[7] ctlp[7].n6 30.8636
R17261 ctlp[7].n6 ctlp[7].n5 4.02551
R17262 ctlp[7].n6 ctlp[7].n0 3.89156
R17263 ctlp[7].n1 ctlp[7] 3.67837
R17264 ctlp[7].n3 ctlp[7].n2 2.25741
R17265 ctlp[7].n2 ctlp[7].n1 0.0509808
R17266 ctlp[7].n5 ctlp[7].n4 0.0389615
R17267 ctlp[7].n5 ctlp[7].n3 0.00159947
R17268 ctln[2].n0 ctln[2] 36.1406
R17269 ctln[2].n0 ctln[2] 12.424
R17270 ctln[2] ctln[2].n0 0.376971
R17271 ctln[4].n0 ctln[4] 13.3519
R17272 ctln[4].n0 ctln[4] 9.6005
R17273 ctln[4] ctln[4].n0 3.2005
R17274 trim[1].n0 trim[1] 9.6005
R17275 trim[1].n0 trim[1] 9.02802
R17276 trim[1] trim[1].n0 3.2005
R17277 result[0].n0 result[0] 9.6005
R17278 result[0].n0 result[0] 9.29247
R17279 result[0] result[0].n0 3.2005
R17280 trim[2].n0 trim[2] 9.6005
R17281 trim[2].n0 trim[2] 8.59446
R17282 trim[2] trim[2].n0 3.2005
R17283 ctln[3].n7 ctln[3].n6 26.3717
R17284 ctln[3].n7 ctln[3] 12.424
R17285 ctln[3].n6 ctln[3].n5 3.7874
R17286 ctln[3].n6 ctln[3].n0 3.62601
R17287 ctln[3].n3 ctln[3] 2.35915
R17288 ctln[3].n5 ctln[3].n3 2.24426
R17289 ctln[3] ctln[3].n7 0.376971
R17290 ctln[3].n5 ctln[3].n4 0.0389615
R17291 ctln[3].n3 ctln[3].n2 0.0141816
R17292 ctln[3].n5 ctln[3].n1 0.00290385
R17293 ctln[5].n0 ctln[5] 17.459
R17294 ctln[5].n0 ctln[5] 9.6005
R17295 ctln[5] ctln[5].n0 3.2005
R17296 result[1].n0 result[1] 9.68341
R17297 result[1].n0 result[1] 9.6005
R17298 result[1] result[1].n0 3.2005
R17299 trim[3].n0 trim[3] 9.6005
R17300 trim[3].n0 trim[3] 9.171
R17301 trim[3] trim[3].n0 3.2005
R17302 ctln[6].n0 ctln[6] 20.2269
R17303 ctln[6].n0 ctln[6] 9.6005
R17304 ctln[6] ctln[6].n0 3.2005
R17305 result[2].n0 result[2] 10.5068
R17306 result[2].n0 result[2] 9.6005
R17307 result[2] result[2].n0 3.2005
R17308 ctln[7].n0 ctln[7] 47.6537
R17309 ctln[7].n0 ctln[7] 12.424
R17310 ctln[7] ctln[7].n0 0.376971
R17311 trim[4] trim[4].n6 24.4636
R17312 trim[4].n6 trim[4].n5 4.02551
R17313 trim[4].n6 trim[4].n0 3.89156
R17314 trim[4].n3 trim[4] 3.50155
R17315 trim[4].n5 trim[4].n3 2.24426
R17316 trim[4].n5 trim[4].n4 0.0389615
R17317 trim[4].n3 trim[4].n2 0.0141816
R17318 trim[4].n5 trim[4].n1 0.00290385
R17319 ctlp[0] ctlp[0] 13.2956
R17320 trimb[0].n0 trimb[0] 9.6005
R17321 trimb[0].n0 trimb[0] 6.81829
R17322 trimb[0] trimb[0].n0 3.2005
R17323 result[3].n0 result[3] 9.6005
R17324 result[3].n0 result[3] 6.90994
R17325 result[3] result[3].n0 3.2005
R17326 ctlp[1] ctlp[1] 17.9087
R17327 result[4].n0 result[4] 11.1139
R17328 result[4].n0 result[4] 9.6005
R17329 result[4] result[4].n0 3.2005
R17330 trimb[1].n0 trimb[1] 9.6005
R17331 trimb[1].n0 trimb[1] 8.59446
R17332 trimb[1] trimb[1].n0 3.2005
R17333 ctlp[2] ctlp[2] 42.1314
R17334 trimb[2].n0 trimb[2] 9.6005
R17335 trimb[2].n0 trimb[2] 6.81829
R17336 trimb[2] trimb[2].n0 3.2005
R17337 result[5].n0 result[5] 9.6005
R17338 result[5].n0 result[5] 9.29247
R17339 result[5] result[5].n0 3.2005
R17340 clk.n0 clk.t6 184.768
R17341 clk.n1 clk.t3 184.768
R17342 clk.n2 clk.t0 184.768
R17343 clk.n3 clk.t1 184.768
R17344 clk.n0 clk.t2 146.208
R17345 clk.n1 clk.t7 146.208
R17346 clk.n2 clk.t4 146.208
R17347 clk.n3 clk.t5 146.208
R17348 clk.n5 clk 51.8509
R17349 clk.n1 clk.n0 40.6397
R17350 clk.n2 clk.n1 40.6397
R17351 clk.n3 clk.n2 40.6397
R17352 clk.n4 clk.n3 27.4116
R17353 clk.n4 clk 9.45048
R17354 clk clk.n5 2.55394
R17355 clk.n5 clk.n4 1.04526
R17356 trimb[3] trimb[3] 14.1928
R17357 ctlp[3] ctlp[3].n6 30.8636
R17358 ctlp[3].n6 ctlp[3].n5 4.02551
R17359 ctlp[3].n6 ctlp[3].n0 3.89156
R17360 ctlp[3].n1 ctlp[3] 3.67837
R17361 ctlp[3].n3 ctlp[3].n2 2.25741
R17362 ctlp[3].n2 ctlp[3].n1 0.0509808
R17363 ctlp[3].n5 ctlp[3].n4 0.0389615
R17364 ctlp[3].n5 ctlp[3].n3 0.00159947
R17365 result[6].n7 result[6].n6 26.3717
R17366 result[6].n7 result[6] 12.424
R17367 result[6].n6 result[6].n5 3.7874
R17368 result[6].n3 result[6] 3.70594
R17369 result[6].n6 result[6].n0 3.62601
R17370 result[6].n5 result[6].n3 2.24426
R17371 result[6] result[6].n7 0.376971
R17372 result[6].n5 result[6].n1 0.0389615
R17373 result[6].n3 result[6].n2 0.0141816
R17374 result[6].n5 result[6].n4 0.00290385
R17375 ctlp[4] ctlp[4] 17.9087
R17376 result[7] result[7] 16.2295
R17377 ctlp[5] ctlp[5] 19.0759
R17378 cal.n0 cal.t1 259.022
R17379 cal.n0 cal.t0 175.798
R17380 cal.n1 cal 73.8015
R17381 cal.n1 cal.n0 8.09539
R17382 cal cal.n1 2.45269
R17383 comp.n0 comp.t0 259.022
R17384 comp.n0 comp.t1 175.798
R17385 comp.n1 comp 23.7663
R17386 comp.n1 comp.n0 8.07392
R17387 comp comp.n1 2.39318
R17388 en.n0 en.t0 224.984
R17389 en.n0 en.t1 187.714
R17390 en en.n0 77.9561
R17391 en.n1 en 9.06717
R17392 en.n1 en 6.98112
R17393 en en.n1 3.02272
R17394 rstn.n0 rstn.t0 259.022
R17395 rstn.n0 rstn.t1 175.798
R17396 rstn.n1 rstn 38.3679
R17397 rstn.n1 rstn.n0 8.07414
R17398 rstn rstn.n1 2.39396
R17399 trimb[4].n0 trimb[4] 9.6005
R17400 trimb[4].n0 trimb[4] 8.59446
R17401 trimb[4] trimb[4].n0 3.2005
R17402 clkc.n0 clkc 80.1792
R17403 clkc.n0 clkc 31.412
R17404 clkc clkc.n0 2.78389
R17405 ctln[0].n0 ctln[0] 9.6005
R17406 ctln[0].n0 ctln[0] 8.73842
R17407 ctln[0] ctln[0].n0 3.2005
R17408 valid valid.n6 32.5529
R17409 valid.n1 valid 5.37628
R17410 valid.n6 valid.n5 3.7874
R17411 valid.n6 valid.n0 3.62601
R17412 valid.n3 valid.n2 2.24841
R17413 valid.n2 valid.n1 0.0509808
R17414 valid.n5 valid.n3 0.0105915
R17415 valid.n5 valid.n4 0.00290385
R17416 sample sample 14.3143
C0 _338_/D _337_/a_761_249# 1.64e-20
C1 _346_/SET_B _337_/a_193_7# 0.00628f
C2 _275_/A _319_/a_27_7# 1.18e-20
C3 _248_/A _222_/a_250_257# 0.076f
C4 _224_/a_250_257# VPWR 0.0131f
C5 _306_/S _254_/B 0.42f
C6 _216_/X _331_/a_761_249# 4.96e-20
C7 _324_/a_193_7# _217_/A 2.31e-19
C8 _324_/a_761_249# _304_/X 1.64e-20
C9 repeater43/X _316_/a_805_7# -7.61e-19
C10 _300_/a_301_257# _300_/Y 1.69e-19
C11 _147_/A _347_/a_1217_7# 9.36e-20
C12 _311_/a_27_7# _310_/D 1.36e-20
C13 _314_/a_761_249# _297_/B 8.22e-19
C14 _314_/a_193_7# _314_/D 0.00541f
C15 _311_/D _310_/a_27_7# 0.00108f
C16 _170_/a_76_159# VPWR 0.00844f
C17 _341_/a_1283_n19# _145_/A 0.0447f
C18 _322_/a_543_7# _269_/A 0.0124f
C19 _279_/Y _217_/X 3.84e-20
C20 _325_/a_543_7# _325_/D 0.0336f
C21 _319_/Q _233_/a_113_257# 0.0511f
C22 _339_/a_27_7# _340_/CLK 0.0805f
C23 _346_/Q _147_/Y 0.128f
C24 _340_/a_27_7# _337_/Q 1.71e-19
C25 _327_/a_1108_7# _217_/X 0.00851f
C26 _327_/a_651_373# _327_/Q 8.32e-19
C27 _215_/A _300_/Y 2.67e-20
C28 clkbuf_2_1_0_clk/A VPWR 4.38f
C29 _326_/a_639_7# repeater43/X 0.00458f
C30 _273_/A _222_/a_250_257# 0.0487f
C31 _326_/a_543_7# _331_/a_193_7# 1.02e-19
C32 _326_/a_27_7# _331_/a_1283_n19# 8.55e-20
C33 _206_/A _332_/Q 0.71f
C34 _326_/a_448_7# _212_/X 1.22e-19
C35 _326_/a_1108_7# _217_/X 0.0371f
C36 _310_/Q VPWR 0.206f
C37 repeater43/X _332_/D 1.28e-19
C38 _346_/a_27_7# _254_/A 1.83e-19
C39 _181_/X _146_/C 2.82e-20
C40 _308_/X _283_/A 0.00693f
C41 _345_/a_193_7# _345_/a_1032_373# -9.67e-21
C42 _222_/a_93_n19# _222_/a_250_257# -6.97e-22
C43 ctlp[6] clkbuf_2_1_0_clk/A 0.0314f
C44 _334_/D _332_/Q 0.0018f
C45 _343_/CLK _333_/Q 0.134f
C46 _300_/a_735_7# VPWR 0.00197f
C47 _300_/a_301_257# VGND 0.00648f
C48 ctln[6] _333_/a_193_7# 7.24e-20
C49 _328_/a_1108_7# _212_/X 3.26e-19
C50 _302_/a_227_7# _347_/a_1108_7# 1.65e-20
C51 _157_/A _181_/X 0.224f
C52 _344_/a_193_7# _301_/a_240_7# 1.25e-20
C53 _284_/a_121_257# VGND -4.1e-19
C54 _211_/a_373_7# _283_/A 0.00196f
C55 _294_/A _254_/B 6.71e-19
C56 _346_/a_1224_7# _346_/SET_B 6.18e-19
C57 output8/a_27_7# _273_/Y 0.0128f
C58 _342_/Q _179_/a_27_7# 1.26e-19
C59 _325_/a_1217_7# _181_/X 8.36e-20
C60 _161_/Y _297_/Y 0.00781f
C61 _173_/a_76_159# _345_/Q 0.037f
C62 _322_/a_27_7# _321_/a_27_7# 2.85e-19
C63 _339_/a_761_249# _338_/D 4.81e-19
C64 _339_/a_193_7# _346_/SET_B 0.0145f
C65 _290_/A _312_/a_1283_n19# 0.0445f
C66 repeater43/X _334_/a_1270_373# -1.54e-19
C67 _309_/a_1283_n19# _310_/D 0.00924f
C68 _309_/a_27_7# _310_/Q 5.93e-20
C69 _337_/a_1217_7# _340_/CLK 8.47e-19
C70 _326_/a_1283_n19# _217_/a_27_7# 7.51e-19
C71 _272_/a_39_257# _304_/X 4.6e-19
C72 _246_/B _224_/a_584_7# 4.55e-19
C73 _316_/Q _315_/a_448_7# 2.63e-19
C74 _297_/A _228_/A 6.18e-19
C75 result[1] _315_/a_1283_n19# 0.00389f
C76 _235_/a_199_7# _330_/Q 2.69e-19
C77 _324_/Q _304_/a_257_159# 0.0149f
C78 _215_/A VGND 1.69f
C79 _200_/a_250_257# _337_/Q 0.0634f
C80 _160_/X _346_/D 0.00221f
C81 _172_/A _301_/a_240_7# 2.02e-20
C82 _164_/Y _344_/Q 0.00603f
C83 _255_/X _305_/a_535_334# 1.66e-21
C84 _325_/a_1108_7# _216_/X 3.36e-20
C85 ctln[4] VPWR 0.415f
C86 _277_/Y VGND 1.14f
C87 _325_/Q _188_/S 6.95e-20
C88 _334_/Q _332_/D 2.66e-20
C89 _279_/Y clkbuf_0_clk/a_110_7# 0.0184f
C90 clkbuf_2_3_0_clk/A _346_/SET_B 0.011f
C91 _324_/Q _177_/A 2.49e-19
C92 _309_/a_1217_7# _265_/B 1.48e-19
C93 _345_/a_1182_221# _160_/X 1.16e-19
C94 _271_/A _227_/A 0.0413f
C95 _271_/Y en 0.00514f
C96 _337_/a_193_7# _337_/a_448_7# -0.00482f
C97 _344_/a_956_373# _297_/Y 0.00251f
C98 _235_/a_113_257# VPWR 0.0777f
C99 _299_/a_215_7# _286_/Y 0.0536f
C100 _188_/S _298_/a_27_7# 2.4e-19
C101 _227_/A _335_/a_27_7# 3.88e-20
C102 _340_/a_27_7# _339_/Q 1.1e-20
C103 _334_/a_805_7# _207_/C 0.00207f
C104 output36/a_27_7# _285_/Y 0.0113f
C105 _313_/D _257_/a_448_7# 1.5e-19
C106 _315_/a_1462_7# VGND 1.17e-19
C107 _346_/SET_B _327_/Q 0.048f
C108 _325_/Q _212_/a_27_7# 4.38e-19
C109 _331_/D _327_/D 2e-20
C110 _324_/a_1283_n19# VPWR 0.0227f
C111 _324_/a_761_249# VGND 0.011f
C112 _339_/a_448_7# _332_/Q 6.45e-21
C113 _342_/a_1108_7# _342_/Q 0.00158f
C114 _329_/a_448_7# _330_/a_27_7# 6.17e-19
C115 _329_/a_27_7# _330_/a_448_7# 6.17e-19
C116 _306_/a_76_159# clkbuf_2_1_0_clk/A 0.00629f
C117 _346_/SET_B _172_/Y 0.00464f
C118 _262_/a_199_7# VGND -3.73e-19
C119 output20/a_27_7# _330_/Q 5.71e-19
C120 _326_/a_543_7# _325_/a_1283_n19# 1.42e-20
C121 _318_/a_1283_n19# _318_/D 1.02e-20
C122 _283_/A _254_/B 0.00706f
C123 _329_/a_448_7# _318_/Q 1.98e-19
C124 _194_/X _263_/a_109_257# 1.41e-19
C125 _248_/A _331_/a_27_7# 6.96e-21
C126 _314_/a_639_7# VGND -0.00152f
C127 _314_/a_1217_7# VPWR 1.91e-19
C128 _297_/A _216_/A 1.05e-20
C129 _343_/a_543_7# VPWR 0.00708f
C130 _343_/a_193_7# VGND 0.0243f
C131 _324_/a_448_7# _297_/B 2.63e-20
C132 _346_/SET_B _313_/a_1270_373# -2.06e-19
C133 _340_/a_193_7# input1/X 4.85e-22
C134 _340_/a_761_249# cal 2.84e-21
C135 _338_/a_639_7# _337_/Q 4.16e-20
C136 _346_/SET_B _337_/a_1462_7# -8.35e-19
C137 _304_/X VGND 1.98f
C138 _157_/A _347_/a_1108_7# 0.00509f
C139 _154_/a_27_7# _204_/Y 8.71e-19
C140 _196_/A _344_/Q 8.08e-19
C141 _344_/a_27_7# _265_/B 2.04e-20
C142 _324_/Q _325_/D 4.32e-20
C143 _331_/CLK _331_/a_27_7# 0.0349f
C144 ctln[7] _204_/Y 1.25e-19
C145 repeater42/a_27_7# _324_/a_543_7# 4.55e-21
C146 _216_/A _223_/a_256_7# 1.84e-19
C147 _216_/A _164_/A 8.73e-21
C148 _236_/B _212_/X 2.82e-20
C149 _316_/D _217_/X 6.97e-20
C150 _314_/D _324_/D 3.16e-19
C151 _345_/a_1032_373# VPWR 0.00441f
C152 _278_/a_68_257# VPWR 0.0248f
C153 _318_/a_1108_7# _304_/X 2.33e-19
C154 _345_/a_476_7# VGND 0.0226f
C155 _258_/S _261_/a_109_257# 4.46e-19
C156 _322_/a_1108_7# _242_/A 8.5e-21
C157 _254_/A _338_/Q 1.64e-20
C158 _160_/A _174_/a_27_257# 1.1e-20
C159 _331_/D _283_/A 3.74e-21
C160 _200_/a_250_257# _339_/Q 1.43e-19
C161 _273_/A _331_/a_27_7# 4.43e-21
C162 _275_/A _254_/A 1.33e-19
C163 _330_/Q _279_/A 0.00125f
C164 _267_/A _312_/Q 0.00343f
C165 _283_/A _330_/a_193_7# 0.00138f
C166 repeater42/a_27_7# _217_/A 0.0115f
C167 _345_/a_381_7# _297_/B 9.95e-19
C168 clk _334_/a_27_7# 0.00946f
C169 input4/X repeater43/X 0.117f
C170 _248_/B _317_/D 7.46e-19
C171 _258_/a_76_159# _336_/Q 6.14e-22
C172 _339_/a_543_7# _337_/a_1283_n19# 8.4e-19
C173 _339_/a_761_249# _337_/a_1108_7# 3.06e-20
C174 _339_/a_1283_n19# _337_/a_543_7# 8.4e-19
C175 _339_/a_1108_7# _337_/a_761_249# 3.06e-20
C176 _217_/a_27_7# _248_/A 0.00666f
C177 _304_/a_257_159# _228_/A 5.18e-20
C178 _330_/Q _218_/a_250_257# 0.00535f
C179 _326_/D _212_/X 0.0468f
C180 _341_/a_1283_n19# _324_/Q 1.31e-21
C181 _256_/a_209_257# _228_/A 4.91e-20
C182 _145_/A _248_/A 2.37e-21
C183 _317_/Q _318_/Q 0.0128f
C184 _277_/A _320_/a_1270_373# 2.51e-20
C185 _331_/a_27_7# _222_/a_93_n19# 4.28e-21
C186 _177_/A _228_/A 0.015f
C187 _339_/a_761_249# _343_/CLK 1.97e-22
C188 _217_/a_27_7# _331_/CLK 1.49e-20
C189 _323_/a_27_7# _227_/A 4.42e-19
C190 _222_/a_256_7# _212_/X 0.0031f
C191 _222_/a_346_7# _327_/Q 0.00505f
C192 _222_/a_250_257# _217_/X 3.61e-19
C193 _218_/a_93_n19# VPWR 0.0275f
C194 _200_/a_346_7# cal 8.76e-19
C195 _272_/a_39_257# VGND 0.0223f
C196 _145_/A _331_/CLK 8.94e-22
C197 _341_/D _149_/a_27_7# 4.77e-20
C198 _254_/Y _254_/B 0.017f
C199 repeater43/X _207_/C 0.99f
C200 _300_/Y VGND 0.0208f
C201 _342_/a_761_249# _175_/Y 3.78e-19
C202 _288_/Y _345_/Q 1.87e-19
C203 output28/a_27_7# _331_/CLK 8.19e-20
C204 _303_/A _347_/a_651_373# 1.63e-19
C205 _329_/a_543_7# _331_/Q 3.19e-20
C206 _322_/a_1108_7# _322_/D 4.94e-20
C207 _338_/Q _309_/D 0.0506f
C208 valid sample 0.076f
C209 _319_/a_448_7# _217_/X 3.4e-21
C210 _255_/B _231_/a_512_7# 2.02e-19
C211 _339_/a_1462_7# _346_/SET_B -7.68e-19
C212 _226_/a_79_n19# _225_/X 0.00476f
C213 _220_/a_256_7# VPWR -2.53e-19
C214 _220_/a_93_n19# VGND 0.00324f
C215 _251_/a_79_n19# _181_/X 0.0523f
C216 _329_/Q _219_/a_250_257# 1.2e-19
C217 _320_/Q _219_/a_256_7# 3.11e-20
C218 _311_/a_27_7# VPWR 0.0762f
C219 input4/X _334_/Q 4.34e-20
C220 _188_/a_439_7# _307_/X 5.37e-22
C221 _164_/Y _306_/S 1.37e-21
C222 _325_/a_543_7# _248_/A 1.12e-19
C223 _316_/Q _315_/D 9.43e-20
C224 _313_/D _336_/a_193_7# 7.55e-20
C225 _271_/A _321_/Q 0.0339f
C226 ctln[4] ctln[3] 6.38e-20
C227 _346_/a_27_7# clkbuf_0_clk/X 6.62e-21
C228 output23/a_27_7# VPWR 0.102f
C229 _304_/a_257_159# _216_/A 0.0335f
C230 _342_/D _185_/A 3.09e-20
C231 output25/a_27_7# _322_/D 1.07e-21
C232 _325_/a_543_7# _331_/CLK 0.00105f
C233 _337_/a_193_7# _337_/D 0.0835f
C234 trimb[1] VGND 0.244f
C235 _212_/a_27_7# _326_/Q 1.3e-21
C236 _323_/a_1283_n19# _154_/A 8.46e-20
C237 _200_/a_93_n19# _267_/A 0.00831f
C238 _165_/X _299_/a_78_159# 0.044f
C239 _167_/X _299_/a_292_257# 0.00248f
C240 _227_/A _335_/a_1217_7# 3.74e-20
C241 _197_/X _336_/a_193_7# 0.00121f
C242 comp output40/a_27_7# 7.19e-19
C243 clk _207_/X 0.0328f
C244 _334_/Q _207_/C 0.0533f
C245 output22/a_27_7# _286_/Y 1.48e-19
C246 _332_/a_543_7# _207_/a_27_7# 1.25e-19
C247 input4/X _191_/B 0.00106f
C248 _255_/B _333_/a_1283_n19# 2.09e-20
C249 ctln[1] _206_/A 1.61e-20
C250 _327_/a_805_7# clkbuf_0_clk/X 4.25e-19
C251 _271_/A _318_/a_193_7# 4.38e-19
C252 _273_/A _325_/a_543_7# 1.06e-19
C253 _344_/a_27_7# clkbuf_2_1_0_clk/A 3.89e-21
C254 _328_/a_193_7# _219_/a_250_257# 2.18e-19
C255 _302_/a_227_7# _346_/SET_B 0.00532f
C256 clkbuf_2_3_0_clk/A _147_/A 0.0114f
C257 _225_/a_145_35# _254_/B 0.00175f
C258 _326_/a_1283_n19# _324_/Q 1.33e-21
C259 _254_/A _313_/a_1108_7# 0.00649f
C260 _340_/a_27_7# _336_/D 3.71e-21
C261 _313_/a_543_7# _157_/a_27_7# 0.0012f
C262 _339_/D _332_/Q 6.34e-20
C263 _281_/Y _194_/A 0.0014f
C264 repeater43/X _150_/C 0.00189f
C265 _326_/D _325_/a_193_7# 6.28e-19
C266 cal _229_/a_556_7# 9.87e-20
C267 input1/X _229_/a_226_257# 2.23e-19
C268 _344_/a_1182_221# _310_/D 9.26e-21
C269 ctln[1] _334_/D 1.08e-19
C270 _179_/a_27_7# _225_/B 1.66e-19
C271 _318_/a_1108_7# VGND -0.00548f
C272 _318_/a_651_373# VPWR -0.00799f
C273 output7/a_27_7# ctln[1] 0.00366f
C274 _191_/B _207_/C 0.00806f
C275 _343_/a_1462_7# VGND 1.97e-19
C276 _192_/B _206_/A 0.0305f
C277 _341_/a_1283_n19# _228_/A 1.05e-19
C278 _286_/B _193_/Y 0.0309f
C279 _196_/A _306_/S 1.2f
C280 _325_/a_543_7# _222_/a_93_n19# 0.0063f
C281 _325_/a_761_249# _222_/a_250_257# 2.68e-19
C282 _294_/Y _164_/A 6.07e-21
C283 _147_/A _172_/Y 9.79e-21
C284 _345_/a_381_7# _275_/Y 0.00275f
C285 _346_/a_652_n19# _301_/X 3.25e-19
C286 _294_/A _164_/Y 0.01f
C287 _307_/a_505_n19# _145_/A 0.0075f
C288 output10/a_27_7# _283_/Y 2.88e-20
C289 _321_/D result[7] 3.46e-19
C290 _211_/a_109_257# _153_/A 1.48e-20
C291 _216_/A _325_/D 0.0287f
C292 _309_/a_1283_n19# VPWR 0.0324f
C293 _309_/a_761_249# VGND -2.99e-19
C294 _188_/S _154_/A 6.47e-22
C295 repeater43/X _317_/a_193_7# 0.0333f
C296 _145_/A _145_/a_113_7# 1.68e-19
C297 _334_/D _192_/B 4.32e-20
C298 clkbuf_0_clk/X _319_/a_27_7# 1.32e-19
C299 _322_/Q _232_/A 2.25e-20
C300 _345_/a_1224_7# VGND 4.35e-20
C301 _305_/a_218_7# _225_/B 0.00133f
C302 _315_/a_27_7# _317_/D 0.0166f
C303 _145_/A _178_/a_27_7# 6.54e-20
C304 _336_/a_1108_7# _254_/B 3.6e-21
C305 _283_/Y _227_/A 1.18e-20
C306 output11/a_27_7# _281_/Y 7.5e-21
C307 _283_/A _330_/a_1462_7# 3.18e-19
C308 _197_/X _199_/a_256_7# 0.00213f
C309 clk _334_/a_1217_7# 7.13e-20
C310 _308_/X _298_/B 0.0061f
C311 _339_/D _337_/a_193_7# 3.45e-20
C312 _321_/a_27_7# _322_/Q 0.00294f
C313 _326_/D _331_/a_639_7# 7.55e-20
C314 repeater43/X _331_/a_1283_n19# 0.00209f
C315 _281_/Y _320_/Q 0.0397f
C316 _191_/a_109_257# _192_/B 8.6e-19
C317 output27/a_27_7# VGND 0.0983f
C318 _149_/a_27_7# _343_/CLK 2.71e-19
C319 _229_/a_226_7# sample 1e-19
C320 _327_/a_193_7# _281_/Y 0.00784f
C321 _309_/a_193_7# _309_/a_543_7# -0.0102f
C322 _309_/a_27_7# _309_/a_1283_n19# -7.73e-20
C323 _319_/Q _216_/X 0.00746f
C324 _295_/a_79_n19# _286_/Y 1.15e-21
C325 _331_/a_27_7# _217_/X 5.57e-20
C326 _331_/a_193_7# _212_/X 3.52e-19
C327 _263_/B _297_/Y 0.0153f
C328 _346_/a_27_7# _286_/Y 5.36e-20
C329 _157_/A _346_/SET_B 0.0127f
C330 output21/a_27_7# _283_/A 0.0386f
C331 _333_/a_543_7# _335_/Q 4.73e-21
C332 _254_/A _309_/D 1.78e-19
C333 _294_/A _196_/A 2.32e-20
C334 clkbuf_2_3_0_clk/A _337_/D 8.74e-22
C335 _192_/B _147_/A 2.66e-19
C336 _191_/B _150_/C 3.99e-20
C337 _188_/a_76_159# _146_/C 0.0161f
C338 _275_/A clkbuf_0_clk/X 0.0716f
C339 _319_/Q _329_/Q 0.0264f
C340 _276_/a_68_257# _319_/a_1283_n19# 0.00469f
C341 _306_/S _332_/a_543_7# 1.35e-21
C342 _275_/Y _311_/a_761_249# 1.68e-19
C343 _327_/a_761_249# _319_/Q 8.26e-21
C344 _330_/D _297_/B 2.65e-21
C345 _149_/A _192_/B 8.1e-20
C346 _306_/a_218_7# VPWR -4.58e-19
C347 _306_/a_218_334# VGND -6.3e-19
C348 output33/a_27_7# trim[3] 0.00247f
C349 _200_/a_93_n19# _194_/X 0.0732f
C350 _324_/Q _248_/A 0.012f
C351 _328_/D VPWR 0.123f
C352 _269_/A _268_/a_39_257# 0.00579f
C353 _251_/X _181_/X 1.01e-19
C354 _311_/a_1217_7# VPWR 2.14e-19
C355 _320_/Q _329_/D 8.81e-20
C356 _311_/a_639_7# VGND 8.73e-20
C357 _263_/B _310_/a_193_7# 3.34e-19
C358 cal _334_/a_805_7# 9.32e-20
C359 _313_/Q _336_/a_639_7# 4.3e-21
C360 _214_/a_27_257# _304_/X 1.24e-20
C361 _327_/a_193_7# _329_/D 5.42e-21
C362 _181_/X _296_/a_213_83# 0.0162f
C363 _271_/Y _335_/a_193_7# 8.72e-20
C364 _262_/a_113_257# _311_/Q 1.09e-19
C365 _290_/A _162_/A 6.51e-20
C366 _216_/X _250_/X 9.6e-21
C367 output26/a_27_7# _331_/CLK 0.00448f
C368 _346_/SET_B _202_/a_584_7# 4.91e-19
C369 _325_/Q _223_/a_93_n19# 0.0636f
C370 _324_/Q _331_/CLK 1e-19
C371 _335_/a_193_7# _335_/a_761_249# -0.0157f
C372 _335_/a_27_7# _335_/a_543_7# -0.00713f
C373 _217_/a_27_7# _217_/X 0.0103f
C374 _340_/CLK _267_/A 0.01f
C375 _337_/Q _313_/a_1283_n19# 4.17e-21
C376 _324_/Q _190_/A 8.76e-20
C377 _146_/C _143_/a_109_7# 0.00144f
C378 _337_/a_1270_373# _337_/Q 5.8e-19
C379 _345_/a_27_7# _344_/a_1032_373# 1.59e-21
C380 _345_/a_1032_373# _344_/a_27_7# 7.45e-21
C381 _255_/a_30_13# _298_/C 0.0119f
C382 _328_/a_193_7# _319_/Q 0.61f
C383 _288_/A _310_/a_1283_n19# 7.06e-19
C384 _180_/a_29_13# _286_/Y 0.0588f
C385 _265_/B _147_/Y 6.2e-21
C386 _335_/a_651_373# VGND 5.6e-19
C387 _335_/a_639_7# VPWR 6.53e-19
C388 _184_/a_439_7# VPWR -2.7e-19
C389 _184_/a_535_334# VGND -1.74e-19
C390 _309_/a_193_7# _306_/a_535_334# 6.61e-21
C391 input1/X _338_/Q 0.372f
C392 _273_/A _324_/Q 1.8e-20
C393 _343_/a_27_7# _342_/a_27_7# 2.13e-21
C394 _298_/B _254_/B 0.0146f
C395 _339_/a_193_7# _339_/D 0.0167f
C396 _287_/a_39_257# _310_/a_1283_n19# 0.0119f
C397 _292_/A _290_/Y 0.0982f
C398 _328_/a_27_7# _329_/D 0.0139f
C399 _320_/a_761_249# _279_/A 5.88e-20
C400 _346_/SET_B _260_/A 0.00782f
C401 _329_/a_27_7# _327_/a_27_7# 3.71e-19
C402 _194_/a_27_7# _254_/B 0.0222f
C403 _326_/a_1283_n19# _216_/A 0.00144f
C404 _196_/A _283_/A 0.16f
C405 _338_/a_448_7# _306_/S 1.16e-19
C406 _333_/a_1108_7# _153_/a_215_257# 2.47e-19
C407 _338_/a_1270_373# _194_/X 9.62e-20
C408 _182_/a_79_n19# _175_/Y 0.0364f
C409 _232_/X _217_/A 0.0719f
C410 _325_/a_651_373# repeater43/X 0.00128f
C411 _209_/X _333_/a_1108_7# 1.01e-19
C412 _344_/a_1296_7# _310_/D 2.62e-20
C413 _215_/A _203_/a_209_257# 2.36e-19
C414 _306_/X clkbuf_2_1_0_clk/A 5.27e-20
C415 _324_/Q _222_/a_93_n19# 2.94e-20
C416 _302_/a_227_7# _147_/A 0.00168f
C417 _277_/A ctlp[4] 0.00927f
C418 _325_/a_543_7# _217_/X 4.16e-19
C419 _275_/Y _309_/a_448_7# 0.00486f
C420 input4/X _339_/Q 5.16e-19
C421 _344_/a_476_7# _160_/X 3.69e-20
C422 _344_/a_381_7# _299_/X 1e-20
C423 output38/a_27_7# trimb[2] 0.00904f
C424 _296_/Y _145_/A 0.283f
C425 _281_/A _248_/A 2.07e-20
C426 _346_/SET_B _261_/A 1.76e-19
C427 _308_/a_505_n19# _308_/S 0.0331f
C428 _293_/a_39_257# VPWR 0.0339f
C429 _320_/a_1108_7# _220_/a_93_n19# 7.84e-20
C430 repeater43/X _317_/a_1462_7# 5.72e-19
C431 _269_/A _316_/a_27_7# 0.00611f
C432 _340_/a_639_7# _340_/Q 9.62e-19
C433 _340_/a_1108_7# _340_/D 7.76e-20
C434 _340_/a_651_373# _193_/Y 0.00352f
C435 _317_/D _242_/B 8.46e-20
C436 _313_/D _299_/X 5.15e-19
C437 ctln[5] _340_/Q 3.08e-19
C438 _279_/Y _193_/Y 0.00262f
C439 _331_/CLK _281_/A 0.484f
C440 _145_/A _146_/a_29_271# 3.37e-19
C441 _248_/A _228_/A 0.0231f
C442 _342_/Q _305_/X 4.66e-20
C443 _322_/a_761_249# _321_/Q 0.00519f
C444 _341_/a_27_7# _342_/Q 7.1e-21
C445 output13/a_27_7# VGND 0.0671f
C446 _333_/a_1108_7# _209_/a_109_257# 3.21e-19
C447 _257_/a_222_53# _194_/A 4.03e-21
C448 repeater43/X cal 0.0569f
C449 _271_/Y _323_/a_193_7# 2.04e-20
C450 _321_/a_1217_7# _322_/Q 1.36e-19
C451 _346_/a_1182_221# _346_/Q 0.00964f
C452 _307_/a_505_n19# _324_/Q 1.08e-19
C453 _311_/a_193_7# _311_/D 0.0126f
C454 _157_/A _156_/a_39_257# 0.056f
C455 _331_/CLK _228_/A 5.86e-22
C456 _145_/A clkbuf_0_clk/a_110_7# 5.05e-19
C457 _346_/a_476_7# _319_/Q 6.47e-20
C458 _322_/a_27_7# VPWR 0.0473f
C459 _330_/Q _214_/a_373_7# 3.45e-19
C460 _304_/a_591_329# _248_/B 5.18e-19
C461 _228_/A _190_/A 1.3e-20
C462 _258_/S _257_/a_222_53# 9.24e-20
C463 _170_/a_76_159# _147_/Y 0.0469f
C464 input4/a_27_7# _338_/a_27_7# 0.0116f
C465 _254_/Y _196_/A 0.0147f
C466 _320_/a_1108_7# VGND 0.0103f
C467 _320_/a_651_373# VPWR 2.32e-19
C468 _258_/S _297_/Y 0.00853f
C469 _323_/a_651_373# VGND 8.21e-19
C470 _323_/a_639_7# VPWR 8.32e-19
C471 _283_/A _332_/a_543_7# 1.1e-20
C472 _181_/a_27_7# _314_/D 2.6e-19
C473 _324_/Q _178_/a_27_7# 0.00389f
C474 output22/a_27_7# _269_/A 0.0206f
C475 _146_/C _147_/A 0.0823f
C476 _322_/a_27_7# _318_/a_543_7# 9.28e-22
C477 _322_/a_543_7# _318_/a_27_7# 2.44e-21
C478 clk _323_/Q 0.00197f
C479 _305_/a_76_159# VPWR 0.0347f
C480 _214_/a_27_257# VGND 0.00223f
C481 _214_/a_109_7# VPWR -7.96e-19
C482 _344_/a_652_n19# VGND 0.00882f
C483 _273_/A _228_/A 0.00266f
C484 _344_/a_1182_221# VPWR -0.00155f
C485 _232_/X _220_/a_250_257# 3.03e-20
C486 _294_/A trim[3] 5.68e-20
C487 _294_/Y _292_/A 0.00253f
C488 _194_/A _310_/a_193_7# 0.00126f
C489 _320_/a_639_7# _297_/B 3.98e-19
C490 _346_/SET_B _221_/a_250_257# 1.86e-19
C491 cal _337_/a_805_7# 8.74e-20
C492 _194_/X _340_/CLK 0.0165f
C493 _330_/Q _246_/a_109_257# 2.52e-19
C494 _255_/B _216_/X 5.23e-20
C495 _343_/a_761_249# _323_/D 0.00181f
C496 _157_/A _147_/A 0.133f
C497 _146_/C _149_/A 0.0952f
C498 _326_/Q _223_/a_93_n19# 0.0565f
C499 clkbuf_2_1_0_clk/A _147_/Y 0.0993f
C500 _344_/a_1602_7# _297_/B 1.38e-21
C501 _260_/A _313_/a_761_249# 1.57e-20
C502 _216_/A _248_/A 0.0903f
C503 _294_/Y _160_/A 0.0165f
C504 _227_/A _333_/a_27_7# 0.00115f
C505 _258_/a_218_7# VGND 4.03e-19
C506 cal _334_/Q 6.06e-19
C507 _325_/a_27_7# _325_/a_1108_7# -2.98e-20
C508 _258_/S _310_/a_193_7# 0.0203f
C509 ctlp[5] _220_/a_93_n19# 6.62e-23
C510 _216_/A _331_/CLK 0.00276f
C511 _342_/a_193_7# VPWR 0.0354f
C512 _290_/A _163_/a_78_159# 0.0106f
C513 _254_/A input1/X 0.344f
C514 _312_/Q _310_/a_1108_7# 6.64e-19
C515 _318_/Q _304_/X 0.139f
C516 _346_/Q _173_/a_226_257# 1.16e-20
C517 _315_/Q _247_/a_113_257# 1.09e-19
C518 _172_/A _314_/Q 1.18e-20
C519 _211_/a_109_7# VGND -0.00159f
C520 _216_/A _190_/A 0.0806f
C521 _198_/a_584_7# VPWR -8.47e-19
C522 _198_/a_256_7# VGND -1.81e-19
C523 _182_/a_79_n19# _341_/Q 0.00514f
C524 _293_/a_39_257# _306_/a_76_159# 0.00114f
C525 _260_/A _156_/a_39_257# 0.00128f
C526 _219_/a_93_n19# _212_/X 0.00605f
C527 cal _191_/B 0.151f
C528 _273_/A _216_/A 0.258f
C529 ctlp[1] _321_/a_27_7# 1.39e-19
C530 _319_/Q _319_/a_543_7# 0.00114f
C531 _240_/B _319_/a_27_7# 1.91e-21
C532 output33/a_27_7# _273_/Y 1.37e-19
C533 _232_/X _314_/Q 2.73e-19
C534 _329_/a_1283_n19# _327_/a_651_373# 5.24e-22
C535 _185_/A _334_/a_27_7# 5.31e-19
C536 _210_/a_307_257# _298_/C 3.18e-20
C537 _327_/a_448_7# _327_/D 0.0023f
C538 _309_/a_543_7# _172_/A 2.49e-20
C539 _338_/D _306_/S 0.00663f
C540 _333_/a_1283_n19# _154_/A 0.0144f
C541 _346_/SET_B _340_/Q 1.13f
C542 input1/X _226_/X 0.292f
C543 _182_/X _175_/Y 0.175f
C544 _307_/a_505_n19# _228_/A 1.1e-20
C545 _323_/a_27_7# _323_/a_543_7# -0.00353f
C546 ctlp[5] VGND 0.563f
C547 _216_/A _222_/a_93_n19# 0.0434f
C548 rstn _332_/a_1283_n19# 8.85e-20
C549 _145_/a_113_7# _228_/A 5.15e-19
C550 _332_/a_193_7# _153_/a_109_53# 0.00209f
C551 _332_/a_27_7# _153_/a_215_257# 0.00623f
C552 _260_/A _147_/A 0.432f
C553 _343_/CLK _207_/a_27_7# 1.47e-19
C554 input1/X _309_/D 4.77e-19
C555 _241_/a_199_7# _304_/X 1.85e-22
C556 _254_/A _286_/Y 0.03f
C557 _178_/a_27_7# _228_/A 1.67e-20
C558 _272_/a_39_257# _318_/Q 3.82e-21
C559 _254_/A _297_/a_27_257# 5.99e-20
C560 _269_/A _316_/a_1217_7# 1.61e-19
C561 _290_/Y _273_/A 0.105f
C562 _286_/B _298_/A 0.00445f
C563 _283_/Y _335_/a_543_7# 2.17e-19
C564 ctln[7] _335_/a_193_7# 0.545f
C565 _283_/A _204_/a_27_257# 6.61e-19
C566 _182_/a_297_257# _227_/A 6.82e-19
C567 _275_/A _240_/B 0.235f
C568 repeater43/X _284_/A 3.29e-20
C569 result[2] _316_/a_1283_n19# 0.017f
C570 _203_/a_209_257# VGND 0.00251f
C571 _203_/a_303_7# VPWR -8.22e-19
C572 _286_/B _336_/a_448_7# 0.00774f
C573 _250_/X _216_/a_27_7# 1.28e-20
C574 _339_/a_543_7# _195_/a_27_257# 3.31e-20
C575 _319_/a_27_7# _328_/Q 5.03e-19
C576 _165_/X _346_/SET_B 0.741f
C577 _175_/Y valid 0.00206f
C578 _271_/A _322_/a_1108_7# 3.46e-19
C579 _320_/Q _242_/A 1.4e-19
C580 _346_/a_1296_7# _346_/Q 5.61e-19
C581 _296_/Y _324_/Q 0.132f
C582 _327_/a_193_7# _242_/A 1.01e-19
C583 _231_/a_306_7# _315_/D 0.00256f
C584 _307_/a_505_n19# _216_/A 3.18e-19
C585 _340_/a_193_7# _336_/a_193_7# 2.08e-22
C586 _340_/a_27_7# _336_/a_761_249# 2.39e-21
C587 _162_/X _227_/A 0.147f
C588 _226_/X _286_/Y 0.0026f
C589 _322_/a_1217_7# VPWR 1.73e-19
C590 _332_/a_193_7# _209_/a_27_257# 4.2e-21
C591 _267_/B _267_/A 0.0142f
C592 _315_/a_761_249# _177_/A 5.02e-21
C593 _330_/Q _330_/a_543_7# 0.00226f
C594 _326_/a_193_7# _242_/A 0.599f
C595 _337_/Q _202_/a_93_n19# 0.0131f
C596 output36/a_27_7# _162_/A 6.35e-19
C597 _302_/a_539_257# _301_/X 0.00213f
C598 _302_/a_77_159# _303_/A 0.00121f
C599 _319_/Q _282_/a_39_257# 9.09e-19
C600 trimb[3] ctlp[3] 0.0172f
C601 _344_/a_1056_7# VGND 8.99e-20
C602 _344_/a_1296_7# VPWR 2.67e-19
C603 _342_/Q _295_/a_676_257# 5.4e-19
C604 _255_/B _295_/a_409_7# 9.88e-19
C605 _315_/Q result[2] 0.00212f
C606 _329_/a_1283_n19# _346_/SET_B 0.0491f
C607 _281_/A _217_/X 1.63e-20
C608 _330_/a_27_7# VGND 0.0293f
C609 _330_/a_761_249# VPWR 0.0182f
C610 _251_/X _346_/SET_B 2.4e-21
C611 cal _337_/Q 0.145f
C612 output18/a_27_7# _279_/A 3.27e-19
C613 _309_/a_448_7# _161_/Y 2.1e-19
C614 _275_/A _328_/Q 0.0417f
C615 _318_/Q VGND 0.742f
C616 _328_/a_27_7# _242_/A 1.5e-19
C617 result[3] VPWR 0.258f
C618 clkbuf_0_clk/a_110_7# _324_/Q 2.69e-19
C619 _308_/X _184_/a_218_334# 0.00121f
C620 _319_/Q clkbuf_2_3_0_clk/A 1.03e-20
C621 _346_/a_652_n19# _297_/Y 1.33e-21
C622 _325_/a_761_249# _324_/Q 5.81e-20
C623 _291_/a_121_257# _312_/Q 3.81e-19
C624 _320_/Q _322_/D 0.192f
C625 _193_/Y _313_/a_27_7# 1.58e-21
C626 _306_/S _313_/a_193_7# 1.73e-20
C627 _194_/X _313_/a_543_7# 4.64e-22
C628 _255_/B _332_/Q 1.62e-19
C629 _337_/a_1108_7# _306_/S 0.00128f
C630 _337_/a_651_373# _194_/X 0.0014f
C631 _337_/a_1283_n19# _193_/Y 0.0145f
C632 _318_/Q _318_/a_1108_7# 0.0738f
C633 ctln[5] rstn 0.139f
C634 _342_/a_805_7# VGND -6.36e-19
C635 _342_/a_1462_7# VPWR 1.67e-19
C636 _305_/X _225_/B 4.11e-19
C637 _194_/A _336_/Q 0.0142f
C638 _191_/B _284_/A 0.00699f
C639 _319_/Q _327_/Q 1.14e-19
C640 _343_/CLK _306_/S 3.24e-19
C641 _286_/B _300_/a_301_257# 1.41e-19
C642 _324_/Q _317_/a_651_373# 1.99e-20
C643 _196_/A _300_/a_27_257# 4.82e-20
C644 _329_/a_651_373# _331_/CLK 0.00107f
C645 _294_/A _273_/Y 5.89e-20
C646 _182_/X _341_/Q 4.81e-19
C647 _294_/Y _273_/A 0.777f
C648 _268_/a_39_257# _315_/a_651_373# 1.01e-19
C649 _196_/A _298_/B 3.92e-19
C650 _285_/A trim[0] 0.0773f
C651 _314_/a_27_7# _347_/a_193_7# 7.86e-20
C652 _314_/a_193_7# _347_/a_27_7# 0.0104f
C653 _338_/D _283_/A 0.00412f
C654 _258_/S _336_/Q 8.17e-20
C655 _297_/A _346_/D 2.75e-20
C656 _290_/A clkbuf_2_3_0_clk/A 1.86e-20
C657 _306_/a_505_n19# _254_/B 0.00108f
C658 _241_/a_199_7# VGND -2.52e-20
C659 _170_/a_226_7# _347_/a_27_7# 1.99e-22
C660 _170_/a_76_159# _347_/a_193_7# 4.53e-20
C661 _333_/D _153_/A 0.058f
C662 _217_/A _223_/a_256_7# 5.21e-19
C663 _304_/X _223_/a_346_7# 0.00131f
C664 _162_/X _347_/Q 0.158f
C665 _312_/a_543_7# _311_/a_761_249# 2.37e-20
C666 _312_/a_1283_n19# _311_/a_193_7# 2.59e-19
C667 _286_/B _215_/A 0.385f
C668 _296_/Y _228_/A 0.00792f
C669 _339_/Q _202_/a_93_n19# 9.19e-19
C670 _340_/a_543_7# _336_/Q 1.17e-20
C671 _330_/Q _331_/Q 0.218f
C672 _326_/D _327_/D 4.14e-21
C673 _341_/a_1108_7# _315_/a_193_7# 8.95e-21
C674 _341_/a_448_7# _315_/a_27_7# 3.28e-20
C675 _329_/a_27_7# repeater43/X 0.0023f
C676 _216_/A _217_/X 0.00429f
C677 _341_/a_1108_7# _298_/A 0.0484f
C678 _277_/Y _286_/B 0.00777f
C679 _332_/a_193_7# _153_/A 7.29e-19
C680 _318_/Q output27/a_27_7# 4.57e-20
C681 _229_/a_226_7# _175_/Y 0.0282f
C682 _240_/B _254_/A 5.23e-20
C683 _298_/B _298_/X 0.0017f
C684 _202_/a_93_n19# _202_/a_256_7# -3.48e-20
C685 _285_/A _311_/Q 2.5e-19
C686 _340_/Q _147_/A 1.8e-20
C687 cal _339_/Q 0.0224f
C688 _290_/A _172_/Y 5.11e-19
C689 _217_/X _221_/a_584_7# 1.77e-19
C690 _344_/a_193_7# _344_/a_476_7# -2.46e-20
C691 _344_/a_27_7# _344_/a_1182_221# -0.00103f
C692 _322_/Q VPWR 0.781f
C693 _236_/B _283_/A 2.4e-20
C694 _216_/X _326_/Q 0.00166f
C695 _294_/Y trim[4] 0.168f
C696 _346_/a_652_n19# _242_/A 1.73e-19
C697 _275_/Y _312_/a_27_7# 0.0209f
C698 _339_/D _260_/A 2.13e-19
C699 _289_/a_39_257# _311_/a_1283_n19# 0.00175f
C700 _340_/CLK _310_/a_1108_7# 2.94e-20
C701 _317_/Q _316_/D 0.011f
C702 _267_/B _194_/X 3.02e-21
C703 _324_/a_27_7# _181_/X 0.00268f
C704 _339_/a_761_249# _340_/D 5.66e-21
C705 _185_/A _226_/a_79_n19# 0.00109f
C706 clkbuf_0_clk/a_110_7# _228_/A 0.00192f
C707 _312_/a_639_7# VPWR 0.00114f
C708 _312_/a_651_373# VGND 0.0014f
C709 _299_/X _299_/a_215_7# 6.6e-19
C710 _196_/A _314_/a_1270_373# 1.4e-20
C711 output40/a_27_7# VGND 0.0734f
C712 output32/a_27_7# VGND 0.0519f
C713 _207_/X _335_/Q 0.218f
C714 _300_/a_27_257# _347_/a_1283_n19# 1.31e-19
C715 _326_/D _283_/A 2.29e-20
C716 _296_/Y _216_/A 1.31e-19
C717 _286_/B _304_/X 2.03e-21
C718 _165_/X _147_/A 7.87e-19
C719 _326_/a_761_249# _326_/Q 0.00182f
C720 clkbuf_0_clk/X _286_/Y 0.0144f
C721 _164_/Y _160_/X 0.0588f
C722 _232_/X _214_/a_109_257# 0.00274f
C723 _251_/X _156_/a_39_257# 5.12e-20
C724 _337_/Q _284_/A 0.281f
C725 rstn _346_/SET_B 2.96e-19
C726 _172_/A _308_/X 0.00265f
C727 ctlp[3] VPWR 0.0695f
C728 _162_/X _297_/B 0.32f
C729 _321_/a_543_7# _248_/A 4.99e-21
C730 clkbuf_2_1_0_clk/A _338_/a_543_7# 5.03e-21
C731 _342_/a_27_7# _172_/A 8.5e-21
C732 _304_/a_306_329# _304_/X 5.45e-19
C733 _330_/a_1217_7# VGND -4.91e-19
C734 _304_/S _296_/a_109_7# 0.00103f
C735 _227_/A _298_/C 0.018f
C736 _342_/D _271_/A 0.00748f
C737 _167_/a_27_257# clkbuf_2_3_0_clk/A 0.00753f
C738 _337_/a_1108_7# _283_/A 6.71e-20
C739 _343_/a_27_7# _298_/X 0.00997f
C740 _321_/a_543_7# _331_/CLK 0.0336f
C741 _143_/a_27_7# _248_/B 4.48e-22
C742 clkbuf_0_clk/a_110_7# _216_/A 0.0172f
C743 _346_/SET_B _310_/a_448_7# 0.00206f
C744 _325_/a_761_249# _216_/A 1.5e-19
C745 _333_/a_639_7# VPWR 8.82e-35
C746 _333_/a_651_373# VGND 0.00703f
C747 _242_/A _319_/a_761_249# 0.00176f
C748 _206_/A _205_/a_79_n19# 0.0487f
C749 _251_/X _147_/A 1.18e-20
C750 _315_/Q _315_/a_543_7# 8.53e-19
C751 _337_/D _340_/Q 0.0217f
C752 _299_/a_78_159# VPWR 0.0222f
C753 _283_/A _343_/CLK 0.0875f
C754 _343_/a_543_7# _176_/a_27_7# 6.88e-20
C755 _319_/Q _331_/a_1270_373# 7.19e-21
C756 _301_/X _267_/A 1.3e-20
C757 input1/X _286_/Y 1.22e-19
C758 _336_/a_543_7# _340_/CLK 4.37e-20
C759 _174_/a_109_257# _344_/Q 5.62e-20
C760 _326_/a_1283_n19# _224_/a_93_n19# 1.36e-20
C761 _297_/A _314_/Q 0.611f
C762 _153_/a_109_53# _190_/A 0.0222f
C763 _153_/a_297_257# _332_/Q 0.00534f
C764 _153_/a_215_257# _333_/Q 0.0694f
C765 _196_/A _160_/X 1.05e-19
C766 _286_/B _300_/Y 4.17e-19
C767 _223_/a_346_7# VGND -0.00161f
C768 _334_/D _205_/a_79_n19# 7.3e-19
C769 _209_/X _333_/Q 8.11e-19
C770 _324_/a_543_7# _325_/D 8.76e-19
C771 repeater43/X _342_/Q 0.0518f
C772 _293_/a_121_257# _313_/Q 2.14e-19
C773 _322_/a_193_7# _322_/a_448_7# -0.00482f
C774 _263_/B _311_/a_761_249# 2.84e-21
C775 _306_/a_218_7# _147_/Y 1.54e-19
C776 _283_/A _178_/a_193_257# 2.12e-21
C777 _344_/a_1602_7# _161_/Y 0.0118f
C778 _217_/A _325_/D 0.0226f
C779 _320_/D _320_/a_448_7# 0.00569f
C780 _343_/CLK _248_/B 1.47e-20
C781 _339_/Q _284_/A 0.0344f
C782 _341_/D _315_/a_27_7# 5.41e-19
C783 _172_/A _254_/B 1.4e-19
C784 _269_/A _226_/X 2.82e-20
C785 clkbuf_2_3_0_clk/A _310_/a_27_7# -4.86e-37
C786 _192_/a_150_257# VGND -3.32e-19
C787 _341_/Q _204_/a_277_7# 2.04e-21
C788 _342_/a_27_7# _244_/B 6.82e-20
C789 _183_/a_553_257# _306_/S 0.00929f
C790 _202_/a_93_n19# _336_/D 0.00157f
C791 _202_/a_256_7# _284_/A 1.41e-19
C792 _329_/a_1270_373# _212_/X 5.8e-20
C793 rstn _206_/A 2.1e-19
C794 _185_/A _323_/Q 0.00521f
C795 _209_/a_27_257# _190_/A 0.0267f
C796 _209_/a_109_257# _333_/Q 0.00482f
C797 _328_/a_761_249# clkbuf_2_1_0_clk/A 4.02e-21
C798 _339_/a_1108_7# _283_/A 0.0404f
C799 _346_/SET_B _336_/a_1283_n19# -0.00982f
C800 _210_/a_307_257# _207_/C 1.68e-19
C801 _318_/Q _214_/a_27_257# 0.0772f
C802 _279_/Y _215_/A 0.00935f
C803 _275_/Y _312_/a_1217_7# 2.47e-21
C804 _336_/Q _201_/a_27_7# 0.0541f
C805 _259_/a_113_257# VGND -0.00365f
C806 _181_/X VPWR 0.881f
C807 _286_/B VGND 1.62f
C808 cal _336_/D 8.1e-20
C809 _199_/a_584_7# _340_/CLK 2.5e-20
C810 _324_/a_1217_7# _181_/X 1.83e-19
C811 _197_/X _179_/a_27_7# 5.44e-20
C812 _339_/D _340_/Q 0.00677f
C813 _315_/a_761_249# _248_/A 0.00969f
C814 rstn _334_/D 2.62e-19
C815 _342_/a_27_7# _323_/D 4.32e-20
C816 _275_/Y _162_/X 0.00804f
C817 output7/a_27_7# rstn 0.00526f
C818 _189_/a_27_7# _192_/B 3.95e-19
C819 _319_/a_805_7# _319_/D 3.81e-19
C820 _160_/X _347_/a_1283_n19# 8.24e-20
C821 _337_/a_27_7# _199_/a_93_n19# 2.75e-21
C822 _316_/a_1108_7# _318_/D 2.93e-20
C823 _342_/Q _191_/B 0.248f
C824 _255_/B _192_/B 0.00828f
C825 _304_/a_306_329# VGND -7.24e-19
C826 _304_/a_288_7# VPWR -1.88e-19
C827 _316_/D _315_/a_193_7# 5.7e-21
C828 _283_/A _331_/a_193_7# 0.00196f
C829 _149_/A _232_/A 0.00256f
C830 output29/a_27_7# _283_/A 0.00228f
C831 _256_/a_209_7# VGND 6.84e-20
C832 _232_/X _331_/D 0.0181f
C833 _169_/Y _173_/a_76_159# 2.9e-20
C834 _279_/Y _324_/a_761_249# 3.41e-21
C835 _293_/a_39_257# _147_/Y 0.00566f
C836 _248_/A _224_/a_93_n19# 1.52e-19
C837 _309_/a_761_249# _286_/B 2.1e-20
C838 _237_/a_113_257# VPWR 0.0161f
C839 repeater43/X _204_/Y 0.0197f
C840 _225_/a_59_35# _206_/A 8.46e-19
C841 _279_/Y _314_/a_639_7# 0.00101f
C842 clkbuf_2_0_0_clk/a_75_172# _346_/SET_B 2.54e-19
C843 _342_/a_1217_7# _172_/A 4.49e-21
C844 _342_/D _186_/a_79_n19# 0.00141f
C845 _345_/a_1182_221# _292_/A 0.00307f
C846 _216_/X _324_/D 0.0135f
C847 _337_/a_27_7# _336_/Q 2.04e-20
C848 _271_/A output15/a_27_7# 0.0296f
C849 _342_/a_27_7# _342_/a_639_7# -0.0015f
C850 _346_/a_476_7# _170_/a_226_7# 9.85e-21
C851 _275_/A clkbuf_2_3_0_clk/a_75_172# 0.0179f
C852 _165_/a_78_159# _160_/X 0.0786f
C853 _343_/Q VPWR 1.14f
C854 _157_/A _250_/X 0.0694f
C855 repeater43/X _298_/a_181_7# 4.67e-20
C856 _325_/Q _327_/Q 2.37e-21
C857 _244_/B _317_/D 0.389f
C858 _345_/a_1182_221# _160_/A 6.16e-20
C859 _333_/a_1283_n19# _153_/B 0.0018f
C860 _346_/SET_B _310_/D 0.146f
C861 _338_/Q _199_/a_256_7# 4.87e-20
C862 _316_/Q _268_/a_39_257# 3.15e-19
C863 _324_/Q _251_/a_215_7# 0.00214f
C864 ctlp[1] VPWR 0.216f
C865 _251_/a_79_n19# _250_/a_78_159# 3.88e-20
C866 _341_/D _298_/B 1.04e-20
C867 _216_/a_27_7# _326_/Q 0.00114f
C868 result[0] _315_/a_1462_7# 1.93e-19
C869 _329_/a_193_7# clkbuf_0_clk/X 0.00115f
C870 clkbuf_0_clk/X _328_/Q 0.255f
C871 _346_/a_1182_221# clkbuf_2_1_0_clk/A 0.00441f
C872 _332_/a_761_249# VGND 0.00192f
C873 _332_/a_1283_n19# VPWR 0.0279f
C874 _315_/D _347_/a_639_7# 4.33e-19
C875 _329_/Q _278_/a_150_257# 6.21e-19
C876 _344_/Q _344_/D 0.203f
C877 _347_/a_1108_7# VPWR 0.00367f
C878 _347_/a_543_7# VGND 8.16e-19
C879 _326_/a_1108_7# _304_/X 0.00211f
C880 _326_/a_1283_n19# _217_/A 0.00484f
C881 _154_/A _332_/Q 0.114f
C882 _153_/A _190_/A 0.00934f
C883 ctlp[7] VGND 0.194f
C884 _167_/X _301_/X 2.54e-19
C885 _323_/D _317_/D 1.18e-20
C886 _334_/Q _204_/Y 0.0785f
C887 _338_/D _194_/a_27_7# 2.7e-22
C888 repeater43/X _321_/a_651_373# 0.00509f
C889 _308_/a_218_7# _181_/X 1.52e-19
C890 _216_/X _279_/A 2.1e-19
C891 _255_/a_30_13# cal 1.13e-19
C892 _336_/a_1283_n19# _313_/a_761_249# 6.87e-21
C893 _314_/Q _347_/a_761_249# 0.00798f
C894 _297_/B _347_/a_651_373# 0.0267f
C895 _314_/D _347_/a_448_7# 2.06e-20
C896 _267_/B _310_/a_1108_7# 0.0106f
C897 _306_/a_218_334# _286_/B 8.9e-20
C898 _263_/a_109_257# _311_/D 9.31e-19
C899 _188_/a_505_n19# _341_/Q 1.01e-19
C900 _258_/S _311_/a_761_249# 8.19e-21
C901 _216_/X _218_/a_250_257# 0.0518f
C902 _346_/a_27_7# _299_/X 0.0147f
C903 _343_/CLK _315_/a_27_7# 0.0685f
C904 _329_/Q _279_/A 0.446f
C905 repeater43/X _153_/a_487_257# 1.09e-20
C906 _165_/a_292_257# VPWR 1.88e-19
C907 _316_/a_27_7# _246_/B 0.00105f
C908 _312_/Q _311_/a_448_7# 1.16e-19
C909 _183_/a_553_257# _283_/A 0.0028f
C910 _279_/Y _300_/Y 0.004f
C911 _191_/B _204_/Y 0.0183f
C912 ctln[7] _333_/a_193_7# 1.97e-20
C913 _239_/a_113_257# _319_/Q 0.00105f
C914 _168_/a_109_7# _346_/Q 1.75e-19
C915 _250_/X _260_/A 1.65e-19
C916 _175_/Y _225_/X 0.134f
C917 _254_/A _336_/a_193_7# 6.33e-20
C918 _341_/a_1108_7# VGND -0.00465f
C919 _341_/a_651_373# VPWR 0.00172f
C920 _216_/X _220_/a_346_7# 1.48e-19
C921 _327_/a_761_249# _218_/a_250_257# 1.06e-19
C922 _284_/A _336_/D 4.06e-20
C923 _338_/a_1108_7# VGND 0.0162f
C924 _338_/a_651_373# VPWR -0.00882f
C925 _184_/a_76_159# _182_/X 0.0141f
C926 _324_/a_27_7# _346_/SET_B 2.47e-21
C927 _178_/a_109_257# _298_/A 0.00127f
C928 _346_/a_1602_7# _277_/Y 0.0035f
C929 _316_/Q _316_/a_27_7# 0.365f
C930 output23/a_27_7# _316_/a_1283_n19# 2.8e-19
C931 _329_/Q _220_/a_346_7# 9.81e-19
C932 _341_/Q _143_/a_181_7# 1.55e-19
C933 _326_/a_1108_7# _272_/a_39_257# 0.00525f
C934 clkbuf_2_1_0_clk/A _319_/a_1283_n19# 0.002f
C935 _318_/Q _330_/a_27_7# 4.53e-21
C936 _325_/a_27_7# _325_/Q 5.26e-21
C937 _331_/Q _212_/a_27_7# 1.77e-20
C938 _328_/a_193_7# _279_/A 0.00935f
C939 _281_/Y _221_/a_93_n19# 0.00856f
C940 _169_/B clkbuf_2_3_0_clk/A 0.103f
C941 _248_/A _318_/D 1.3e-19
C942 _271_/A _316_/a_761_249# 2.27e-21
C943 _285_/A _164_/Y 1.79e-19
C944 _229_/a_76_159# VPWR 0.0296f
C945 _336_/a_1283_n19# _147_/A 1.07e-20
C946 _317_/Q _317_/a_1270_373# 8.41e-20
C947 _290_/A _261_/A 0.0023f
C948 _242_/A _317_/a_1283_n19# 8.29e-20
C949 _251_/a_215_7# _228_/A 0.045f
C950 _271_/A _320_/Q 0.0134f
C951 _337_/Q _310_/a_761_249# 3.71e-19
C952 _340_/a_639_7# VPWR 8.13e-19
C953 _340_/a_651_373# VGND 6.14e-19
C954 _236_/B _242_/B 0.945f
C955 _331_/CLK _318_/D 0.0171f
C956 _255_/B _146_/C 0.259f
C957 ctln[5] VPWR 0.99f
C958 _279_/Y VGND 0.831f
C959 _283_/A _331_/a_1462_7# 4.85e-19
C960 _316_/a_448_7# VGND -2.01e-19
C961 _316_/a_1270_373# VPWR 6.65e-20
C962 input1/X _269_/A 3.28e-20
C963 _345_/a_193_7# _346_/SET_B 0.0178f
C964 _343_/a_761_249# _248_/A 1.47e-19
C965 _324_/a_543_7# _331_/CLK 1.4e-19
C966 _344_/a_193_7# _164_/Y 8.08e-20
C967 _344_/a_476_7# _164_/A 0.00297f
C968 _162_/X _171_/a_292_257# 0.00449f
C969 _258_/S _309_/a_448_7# 2.13e-19
C970 output10/a_27_7# input4/X 1.13e-19
C971 _204_/a_27_7# VPWR -0.0011f
C972 _248_/A _217_/A 0.364f
C973 _328_/Q _286_/Y 0.0694f
C974 _337_/Q _264_/a_113_257# 0.0113f
C975 _255_/B _157_/A 0.00931f
C976 _208_/a_215_7# VPWR -0.00194f
C977 _208_/a_292_257# VGND -0.00119f
C978 _326_/a_1270_373# _330_/Q 7.63e-22
C979 _326_/Q _327_/Q 0.0128f
C980 _315_/Q output23/a_27_7# 0.032f
C981 output22/a_27_7# _316_/Q 5.41e-22
C982 _255_/X clkbuf_0_clk/X 1.68e-19
C983 _313_/a_448_7# _225_/B 1.54e-20
C984 _327_/a_1108_7# VGND 0.00527f
C985 _327_/a_651_373# VPWR -0.00787f
C986 _345_/a_1296_7# _292_/A 0.00106f
C987 _342_/a_543_7# _342_/D 0.036f
C988 _346_/a_1032_373# _346_/D 1.18e-19
C989 _273_/A _324_/a_543_7# 6.88e-19
C990 _144_/A _298_/A 4.08e-19
C991 _331_/CLK _217_/A 0.0801f
C992 _316_/D _304_/X 0.0122f
C993 repeater43/X _315_/a_448_7# 1.66e-19
C994 _172_/A _164_/Y 2.97e-20
C995 _195_/a_109_257# _306_/S 0.0119f
C996 _195_/a_27_257# _193_/Y 0.0112f
C997 _195_/a_109_7# _340_/Q 8.73e-19
C998 _326_/a_651_373# VPWR -0.00938f
C999 _326_/a_1108_7# VGND -0.00412f
C1000 _215_/A _313_/a_27_7# 0.0336f
C1001 repeater43/X en 4.11e-20
C1002 input4/X _227_/A 4.31e-20
C1003 _318_/Q _241_/a_199_7# 8.72e-20
C1004 _274_/a_39_257# _279_/A 0.00422f
C1005 _306_/S _344_/D 8.37e-20
C1006 _251_/a_215_7# _216_/A 3.02e-19
C1007 _251_/a_79_n19# _250_/X 0.00415f
C1008 _341_/Q _304_/S 0.187f
C1009 _329_/a_1462_7# clkbuf_0_clk/X 5.26e-19
C1010 _273_/A _217_/A 0.0118f
C1011 _288_/A _161_/Y 5.19e-19
C1012 _346_/a_1296_7# clkbuf_2_1_0_clk/A 6.52e-19
C1013 _301_/X _301_/a_51_257# 0.00412f
C1014 result[0] VGND 0.183f
C1015 _327_/a_448_7# repeater42/a_27_7# 0.00124f
C1016 rstn _339_/D 2.04e-20
C1017 _273_/A _346_/D 1.4e-19
C1018 _328_/a_448_7# VPWR -0.00322f
C1019 _328_/a_1283_n19# VGND 4.51e-19
C1020 _275_/A _299_/X 4.32e-20
C1021 _147_/A _310_/D 3.19e-20
C1022 _346_/Q _306_/S 5.16e-19
C1023 _162_/X _161_/Y 0.107f
C1024 _227_/A _207_/C 0.00124f
C1025 _269_/A _286_/Y 0.701f
C1026 _271_/A _334_/a_27_7# 0.0559f
C1027 _191_/B _225_/B 0.00889f
C1028 _322_/D result[7] 9.33e-20
C1029 _255_/X input1/X 0.0082f
C1030 _321_/a_448_7# result[7] 2.15e-19
C1031 _217_/A _222_/a_93_n19# 0.0026f
C1032 _314_/D _347_/D 1.27e-20
C1033 _337_/Q _336_/a_27_7# 1.95e-19
C1034 _339_/Q _310_/a_761_249# 7.28e-22
C1035 _341_/Q _225_/X 0.0061f
C1036 _307_/X _341_/Q 0.322f
C1037 _334_/a_448_7# VPWR -0.00183f
C1038 _334_/a_1283_n19# VGND 0.00599f
C1039 _257_/a_79_159# _260_/A 0.011f
C1040 _172_/Y _170_/a_226_7# 7.78e-20
C1041 _272_/a_39_257# _316_/D 5.27e-19
C1042 _312_/Q _311_/D 0.00571f
C1043 _172_/A _196_/A 0.179f
C1044 cal _210_/a_307_257# 2.27e-19
C1045 _145_/A _298_/A 1.36f
C1046 _320_/Q _330_/D 0.0491f
C1047 _167_/X _166_/Y 0.0341f
C1048 _325_/Q _146_/C 2.87e-20
C1049 _317_/Q _324_/Q 5.62e-19
C1050 _216_/a_27_7# _324_/D 2.27e-20
C1051 _343_/a_27_7# _343_/CLK 0.017f
C1052 clkbuf_2_1_0_clk/A _212_/X 2.52e-19
C1053 _319_/Q _165_/X 1.03e-20
C1054 _325_/a_27_7# _326_/Q 0.00724f
C1055 _216_/A _193_/Y 1.86e-22
C1056 _273_/A _272_/a_121_257# 3.49e-19
C1057 _294_/A _344_/D 2.04e-20
C1058 _323_/a_1108_7# _343_/Q 2.42e-19
C1059 _188_/S _182_/X 0.00212f
C1060 _346_/SET_B VPWR 3.09f
C1061 _254_/A _314_/a_1283_n19# 4.69e-21
C1062 en _191_/B 1.61e-19
C1063 _316_/Q _316_/a_1217_7# 9.26e-19
C1064 _329_/a_448_7# _281_/A 0.0249f
C1065 _267_/A _297_/Y 0.00654f
C1066 input1/X _264_/a_199_7# 7.18e-21
C1067 _329_/a_543_7# _281_/Y 0.00234f
C1068 _172_/A _298_/X 6.76e-22
C1069 _342_/a_27_7# _177_/A 4.9e-20
C1070 output18/a_27_7# ctlp[4] 0.00402f
C1071 _317_/a_1108_7# _326_/Q 2.84e-19
C1072 _227_/A _150_/C 3.94e-19
C1073 _188_/a_76_159# VPWR 0.0079f
C1074 _346_/a_1602_7# VGND 0.00805f
C1075 _333_/a_193_7# _333_/a_761_249# -0.0133f
C1076 _333_/a_27_7# _333_/a_543_7# -0.00959f
C1077 _337_/Q _199_/a_250_257# 2.47e-19
C1078 _233_/a_113_257# _331_/Q 0.00382f
C1079 _309_/a_27_7# _346_/SET_B 0.0132f
C1080 _335_/a_27_7# _207_/X 6.75e-19
C1081 _335_/a_1108_7# _208_/a_215_7# 1.89e-19
C1082 _329_/a_1283_n19# _319_/Q 0.0321f
C1083 _163_/a_215_7# VGND 0.0421f
C1084 _290_/A _165_/X 0.00942f
C1085 _248_/A _314_/Q 1.98e-19
C1086 _343_/a_1108_7# _226_/a_79_n19# 9.3e-20
C1087 _192_/a_68_257# _254_/B 6.85e-20
C1088 _240_/B _328_/Q 0.0116f
C1089 _316_/D VGND 0.553f
C1090 _318_/a_448_7# _248_/A 4.04e-19
C1091 _345_/a_796_7# _346_/SET_B 5.27e-19
C1092 _300_/Y _313_/a_27_7# 2e-19
C1093 _267_/A _310_/a_193_7# 1.29e-19
C1094 _261_/A _310_/a_27_7# 1.31e-19
C1095 _339_/Q _336_/a_27_7# 6.58e-20
C1096 _283_/Y _194_/A 1.26e-21
C1097 _340_/CLK _311_/a_448_7# 2.59e-19
C1098 _328_/a_761_249# _328_/D 2.33e-20
C1099 _192_/B _154_/A 0.0061f
C1100 _331_/CLK _314_/Q 1.07e-20
C1101 _323_/a_27_7# _334_/a_27_7# 1.22e-20
C1102 _200_/a_93_n19# _311_/D 7.32e-20
C1103 _329_/a_543_7# _329_/D 0.0336f
C1104 _283_/Y _338_/a_193_7# 7.75e-19
C1105 _321_/D _318_/a_761_249# 2.02e-19
C1106 _318_/a_448_7# _331_/CLK 6.51e-21
C1107 _286_/B _203_/a_209_257# 3.79e-19
C1108 _196_/A _203_/a_80_n19# 2.24e-20
C1109 output38/a_27_7# trimb[3] 0.00292f
C1110 _337_/Q _225_/B 2.09e-21
C1111 _336_/a_761_249# _202_/a_93_n19# 0.00291f
C1112 _336_/a_193_7# _202_/a_250_257# 1.11e-19
C1113 _255_/B _251_/a_79_n19# 5.73e-20
C1114 output37/a_27_7# _288_/Y 0.0105f
C1115 _143_/a_109_7# VPWR -2.8e-19
C1116 _219_/a_346_7# _319_/D 3.03e-20
C1117 repeater43/X _315_/D 0.00526f
C1118 _306_/S _340_/D 0.166f
C1119 repeater43/a_27_7# VGND 0.0266f
C1120 output14/a_27_7# _322_/a_448_7# 8.29e-19
C1121 ctlp[0] _322_/a_27_7# 7.87e-20
C1122 _254_/A _299_/X 0.327f
C1123 _273_/A _314_/Q 1.05e-19
C1124 repeater43/X _324_/a_651_373# -5.55e-35
C1125 _305_/a_218_334# _194_/A 0.00206f
C1126 cal _336_/a_761_249# 3.59e-21
C1127 input1/X _336_/a_193_7# 0.607f
C1128 _251_/X _250_/X 3.1e-20
C1129 _222_/a_346_7# VPWR -9.97e-19
C1130 _222_/a_250_257# VGND -0.00285f
C1131 _332_/a_805_7# _153_/B 5.18e-19
C1132 trim[0] _292_/A 6.68e-20
C1133 _324_/a_1283_n19# _212_/X 0.00108f
C1134 _324_/a_1108_7# _327_/Q 1.31e-21
C1135 _144_/A _304_/X 3.27e-20
C1136 _250_/X _296_/a_213_83# 1.36e-20
C1137 _343_/a_448_7# repeater43/X 3.15e-19
C1138 _329_/a_27_7# _329_/a_761_249# -0.0166f
C1139 output11/a_27_7# _283_/Y 2.3e-19
C1140 _177_/A _317_/D 0.0037f
C1141 _206_/A VPWR 1.26f
C1142 _145_/A _215_/A 0.037f
C1143 _271_/A _334_/a_1217_7# 1.01e-19
C1144 _331_/a_27_7# _304_/X 2.89e-21
C1145 _326_/D repeater42/a_27_7# 6.51e-20
C1146 _319_/a_448_7# VGND 0.00411f
C1147 _319_/a_1270_373# VPWR 1.16e-19
C1148 _313_/a_761_249# VPWR 0.0018f
C1149 _313_/a_27_7# VGND -0.0805f
C1150 _346_/SET_B _311_/a_651_373# 0.00252f
C1151 _338_/Q _311_/a_1283_n19# 5.76e-19
C1152 _337_/a_448_7# VPWR -8.01e-19
C1153 _337_/a_1283_n19# VGND -0.0172f
C1154 _217_/A _217_/X 0.0715f
C1155 _297_/B _345_/Q 0.00628f
C1156 _324_/D _327_/Q 1.04e-19
C1157 _342_/a_761_249# _341_/a_761_249# 1.8e-21
C1158 _342_/a_193_7# _341_/a_543_7# 9.01e-19
C1159 _342_/a_543_7# _341_/a_193_7# 1.7e-20
C1160 _339_/Q _199_/a_250_257# 0.111f
C1161 _344_/a_1032_373# _162_/A 7.9e-19
C1162 _197_/X _305_/X 3.09e-20
C1163 _343_/CLK ctln[0] 5.52e-19
C1164 _334_/D VPWR 0.395f
C1165 _320_/Q _322_/a_761_249# 0.0187f
C1166 _166_/Y _301_/a_51_257# 2.66e-19
C1167 _333_/D _254_/B 0.0152f
C1168 _292_/A _311_/Q 0.154f
C1169 _212_/X _278_/a_68_257# 0.00114f
C1170 output7/a_27_7# VPWR 0.0978f
C1171 _190_/a_27_7# _153_/B 1.39e-20
C1172 _310_/a_1283_n19# _284_/A 1.57e-20
C1173 _197_/X _338_/a_27_7# 1.93e-21
C1174 _307_/a_218_7# VPWR -4.66e-19
C1175 _307_/a_218_334# VGND -4.17e-19
C1176 _323_/D _298_/X 0.00955f
C1177 _254_/a_109_257# VGND -7.75e-19
C1178 _345_/a_1140_373# _345_/Q 7.87e-19
C1179 _156_/a_39_257# VPWR 0.0574f
C1180 _165_/X _167_/a_27_257# 0.00683f
C1181 _317_/Q _216_/A 3.98e-19
C1182 _167_/X _167_/a_109_257# 0.00256f
C1183 rstn _195_/a_109_7# 0.00301f
C1184 _324_/a_805_7# _304_/S 0.0021f
C1185 _325_/a_1217_7# _326_/Q 7.95e-20
C1186 _309_/a_543_7# trim[4] 3.28e-20
C1187 input1/X _199_/a_256_7# 7.58e-19
C1188 _271_/A _226_/a_79_n19# 0.0159f
C1189 _217_/a_27_7# _304_/X 0.0239f
C1190 _191_/a_109_257# VPWR 7.37e-19
C1191 _319_/Q _234_/a_109_257# 0.0013f
C1192 _178_/a_109_257# VGND -5.25e-19
C1193 _327_/Q _279_/A 0.0331f
C1194 _304_/S _314_/D 4.88e-20
C1195 _319_/Q _321_/a_27_7# 1.44e-19
C1196 _324_/Q _315_/a_193_7# 7.58e-20
C1197 _340_/a_761_249# _197_/X 0.00567f
C1198 _324_/Q _298_/A 0.0565f
C1199 _194_/X _310_/a_193_7# 2.68e-20
C1200 _183_/a_471_7# _227_/A 6.92e-21
C1201 _218_/a_93_n19# _212_/X 0.00148f
C1202 _147_/A VPWR 0.599f
C1203 _343_/a_1108_7# _323_/Q 0.00233f
C1204 clkbuf_2_3_0_clk/A _311_/a_193_7# 2.89e-20
C1205 _328_/a_1283_n19# _320_/a_1108_7# 0.00177f
C1206 _328_/a_1108_7# _320_/a_1283_n19# 0.00177f
C1207 _302_/a_77_159# _347_/Q 4.83e-20
C1208 _325_/a_193_7# _324_/a_1283_n19# 0.0157f
C1209 _325_/a_27_7# _324_/a_1108_7# 0.00111f
C1210 _167_/X _297_/Y 0.00599f
C1211 _283_/Y _334_/a_27_7# 2.12e-19
C1212 _157_/A _314_/a_193_7# 0.00209f
C1213 _255_/a_30_13# _342_/Q 0.0336f
C1214 _255_/a_184_257# _255_/B 7.15e-19
C1215 _320_/a_27_7# _319_/a_27_7# 1.62e-20
C1216 _165_/a_215_7# _161_/Y 0.0651f
C1217 _149_/A VPWR 0.743f
C1218 _169_/B _260_/A 0.0886f
C1219 _309_/a_1217_7# _346_/SET_B -3.08e-19
C1220 _335_/a_1217_7# _207_/X 5.2e-19
C1221 _343_/a_651_373# _226_/X 5.87e-20
C1222 _212_/X _220_/a_256_7# 9.4e-19
C1223 _341_/a_1283_n19# _317_/D 9.29e-20
C1224 _339_/a_448_7# VPWR 0.0028f
C1225 _339_/a_1283_n19# VGND -0.00193f
C1226 _327_/a_448_7# _232_/X 0.00278f
C1227 _339_/Q _336_/a_1217_7# 3.38e-20
C1228 _308_/a_218_7# _206_/A 3.65e-21
C1229 _265_/B _344_/Q 0.0867f
C1230 _153_/B _332_/Q 0.446f
C1231 _199_/a_93_n19# _267_/A 4.84e-20
C1232 _258_/a_505_n19# _340_/CLK 1.56e-20
C1233 _340_/CLK _311_/D 0.346f
C1234 _325_/a_543_7# _304_/X 0.0357f
C1235 _325_/a_761_249# _217_/A 7.46e-19
C1236 _325_/a_27_7# _324_/D 1.66e-19
C1237 _277_/Y input1/a_75_172# 1.84e-19
C1238 _294_/Y output5/a_27_7# 2.86e-19
C1239 _283_/Y _338_/a_1462_7# 2.3e-19
C1240 _283_/A _340_/D 0.00734f
C1241 _326_/a_448_7# _232_/X 0.0014f
C1242 output38/a_27_7# VPWR 0.161f
C1243 _309_/a_27_7# _147_/A 1.63e-20
C1244 input4/X _335_/a_543_7# 3.73e-19
C1245 repeater43/X _335_/a_193_7# -0.00481f
C1246 _336_/a_27_7# _336_/D 0.0449f
C1247 _336_/a_761_249# _284_/A 0.00275f
C1248 _330_/Q _331_/a_543_7# 0.0107f
C1249 _255_/B _251_/X 1.99e-20
C1250 _258_/S _312_/a_27_7# 1.44e-20
C1251 _288_/A _263_/B 0.00101f
C1252 _144_/A VGND 0.167f
C1253 _318_/a_193_7# _317_/a_193_7# 1.36e-19
C1254 _318_/a_761_249# _317_/a_27_7# 6.27e-20
C1255 _255_/B _296_/a_213_83# 9.62e-19
C1256 _312_/a_1283_n19# _312_/Q 0.0624f
C1257 _267_/A _336_/Q 2.94e-20
C1258 _260_/a_27_257# _284_/A 2.13e-19
C1259 cal _227_/A 0.0118f
C1260 _331_/a_27_7# VGND -0.0312f
C1261 _331_/a_761_249# VPWR 0.00532f
C1262 _287_/a_39_257# _263_/B 3.23e-20
C1263 _200_/a_346_7# _197_/X 6.48e-19
C1264 _320_/a_543_7# _346_/SET_B 0.0239f
C1265 _275_/Y _345_/Q 0.00877f
C1266 _343_/D _269_/A 0.615f
C1267 _275_/A _320_/a_27_7# 7e-21
C1268 _335_/a_1108_7# _206_/A 0.00255f
C1269 _335_/a_543_7# _207_/C 1.27e-20
C1270 _164_/A _164_/Y 0.0255f
C1271 _294_/Y comp 1.23e-19
C1272 repeater43/X _318_/a_805_7# 0.00115f
C1273 _344_/a_27_7# _346_/SET_B 0.0114f
C1274 _316_/a_651_373# _244_/B 1.23e-20
C1275 _302_/a_77_159# _297_/B 0.0256f
C1276 _260_/A _314_/a_193_7# 3.19e-20
C1277 _181_/X _330_/a_639_7# 4.29e-20
C1278 _313_/a_1217_7# VGND -3.65e-19
C1279 _341_/D _172_/A 4.25e-20
C1280 _258_/a_218_334# _346_/SET_B 5.45e-19
C1281 _328_/a_1283_n19# ctlp[5] 5.86e-20
C1282 _344_/a_1224_7# _292_/A 3.77e-19
C1283 _283_/Y _207_/X 6e-20
C1284 _335_/a_448_7# _343_/CLK 8.08e-19
C1285 _335_/D _334_/a_1108_7# 3.56e-36
C1286 _335_/a_193_7# _334_/Q 0.00157f
C1287 _337_/D VPWR 0.307f
C1288 clkbuf_0_clk/X _299_/X 2.11e-20
C1289 _315_/a_193_7# _228_/A 3.73e-19
C1290 _228_/A _298_/A 0.0133f
C1291 _217_/a_27_7# VGND 0.0595f
C1292 _297_/A _196_/A 3.87e-20
C1293 _344_/a_1032_373# _163_/a_78_159# 2.86e-19
C1294 output13/a_27_7# repeater43/a_27_7# 0.00137f
C1295 _214_/a_109_257# _331_/CLK 7.48e-19
C1296 trim[0] _273_/A 9.23e-19
C1297 _247_/a_199_7# _232_/A 1.58e-19
C1298 _247_/a_113_257# _248_/B 0.0671f
C1299 _271_/A _323_/Q 0.0253f
C1300 _145_/A VGND 0.147f
C1301 _324_/Q _215_/A 0.00446f
C1302 _346_/SET_B _198_/a_93_n19# 0.0117f
C1303 _186_/a_79_n19# _226_/a_79_n19# 8.51e-20
C1304 output28/a_27_7# VGND 0.103f
C1305 _147_/Y _347_/a_1108_7# 5.47e-19
C1306 _308_/X _248_/A 4.28e-21
C1307 result[3] _316_/a_1283_n19# 9.05e-19
C1308 _320_/Q _330_/a_1283_n19# 0.0376f
C1309 _342_/a_27_7# _248_/A 0.0229f
C1310 _209_/X _306_/S 0.224f
C1311 _326_/Q _221_/a_250_257# 7.23e-21
C1312 _146_/a_112_13# VGND 5.6e-20
C1313 _343_/a_27_7# output30/a_27_7# 5.52e-19
C1314 repeater43/a_27_7# _323_/a_651_373# 4.93e-22
C1315 repeater43/X _323_/a_193_7# 0.0173f
C1316 _346_/SET_B _171_/a_215_7# 4.42e-21
C1317 _255_/B _232_/A 0.00932f
C1318 _225_/B _336_/D 4.18e-20
C1319 _184_/a_76_159# _225_/X 0.00123f
C1320 _184_/a_505_n19# _147_/A 0.00222f
C1321 _188_/a_505_n19# _188_/S 0.0344f
C1322 _307_/X _184_/a_76_159# 4.33e-20
C1323 _301_/a_51_257# _297_/Y 0.113f
C1324 _331_/a_1108_7# _246_/B 3.56e-36
C1325 _316_/Q _317_/a_761_249# 1.02e-20
C1326 _216_/A _298_/A 2.67e-19
C1327 _183_/a_1241_257# VPWR 0.00692f
C1328 _273_/A _311_/Q 0.00404f
C1329 _199_/a_93_n19# _194_/X 0.0325f
C1330 _324_/a_761_249# _324_/Q 7.77e-19
C1331 clk _269_/Y 0.0176f
C1332 _328_/a_1108_7# _320_/D 4.41e-20
C1333 _325_/a_543_7# VGND 0.00187f
C1334 _325_/a_1108_7# VPWR 0.0101f
C1335 _236_/B _232_/X 0.55f
C1336 _172_/A _143_/a_27_7# 5.47e-21
C1337 _271_/A _317_/a_1283_n19# 0.00759f
C1338 _286_/B _192_/a_150_257# 9.54e-19
C1339 _323_/a_1108_7# _206_/A 6.76e-20
C1340 _207_/a_109_7# _153_/A 1.09e-19
C1341 _339_/a_193_7# _153_/B 2.72e-20
C1342 _290_/A trimb[0] 9.63e-19
C1343 _212_/X _328_/D 0.108f
C1344 _341_/D _244_/B 0.0063f
C1345 _339_/D VPWR 0.198f
C1346 _324_/Q _304_/X 0.199f
C1347 _168_/a_109_7# clkbuf_2_1_0_clk/A 0.00204f
C1348 _194_/X _336_/Q 0.139f
C1349 _333_/a_1283_n19# _332_/a_1108_7# 9.4e-21
C1350 _313_/Q _340_/CLK 2.06e-19
C1351 _317_/a_805_7# VPWR 2.99e-19
C1352 _323_/a_1108_7# _334_/D 8.01e-21
C1353 _323_/a_448_7# _343_/CLK 0.0158f
C1354 _326_/D _232_/X 0.00416f
C1355 _227_/A _284_/A 3.96e-19
C1356 _271_/A result[7] 0.00468f
C1357 _297_/A _347_/a_1283_n19# 0.00304f
C1358 repeater43/X _335_/a_1462_7# -9.14e-19
C1359 _258_/a_505_n19# _313_/a_543_7# 0.00214f
C1360 _337_/Q _311_/a_543_7# 4.53e-20
C1361 _216_/X _331_/Q 0.108f
C1362 _258_/S _288_/A 0.0121f
C1363 _292_/A _312_/a_1270_373# 9.87e-20
C1364 _172_/A _313_/a_193_7# 4.6e-20
C1365 input1/a_75_172# VGND 0.0591f
C1366 _276_/a_150_257# VPWR -4.41e-19
C1367 _299_/X _286_/Y 0.0294f
C1368 _248_/A _317_/D 0.285f
C1369 _330_/Q _280_/a_68_257# 0.0239f
C1370 _331_/a_1217_7# VGND 7.96e-19
C1371 _304_/a_306_329# _286_/B 9.46e-20
C1372 _258_/S _162_/X 1.49e-19
C1373 _325_/Q _230_/a_27_7# 8.11e-21
C1374 _303_/A _315_/D 0.00651f
C1375 _258_/S _287_/a_39_257# 1.28e-20
C1376 _185_/A _175_/Y 0.0137f
C1377 _215_/A _228_/A 0.2f
C1378 _169_/B _165_/X 0.0269f
C1379 _211_/a_27_257# _206_/A 0.0248f
C1380 _323_/a_27_7# _323_/Q 0.00592f
C1381 _256_/a_80_n19# _181_/X 2.25e-19
C1382 _256_/a_209_257# _196_/A 0.047f
C1383 clkbuf_2_3_0_clk/a_75_172# _328_/Q 5.05e-20
C1384 _344_/a_586_7# _346_/SET_B 4.73e-19
C1385 _236_/B _244_/B 2.67e-20
C1386 _343_/a_1270_373# cal 8.78e-20
C1387 _331_/CLK _317_/D 0.0116f
C1388 _189_/a_27_7# _225_/a_59_35# 0.00543f
C1389 _290_/A _310_/D 0.498f
C1390 _190_/A _203_/a_209_7# 0.00116f
C1391 _308_/S _191_/B 0.0456f
C1392 _283_/Y _339_/a_27_7# 2.43e-20
C1393 _336_/a_639_7# _340_/Q 1.09e-20
C1394 _336_/a_651_373# _193_/Y 4.66e-20
C1395 _254_/B _190_/A 0.00992f
C1396 _172_/A _307_/a_535_334# 1.44e-19
C1397 _242_/A clkbuf_1_1_0_clk/a_75_172# 8.35e-19
C1398 _294_/A _265_/B 0.00838f
C1399 _323_/a_761_249# _226_/X 2.32e-21
C1400 _272_/a_39_257# _324_/Q 2.76e-20
C1401 _174_/a_109_7# VPWR -6.75e-19
C1402 _174_/a_27_257# VGND -0.00227f
C1403 _150_/a_27_7# VPWR 0.0764f
C1404 _306_/X _346_/SET_B 0.0123f
C1405 _335_/D _343_/CLK 0.00287f
C1406 _306_/S _314_/a_27_7# 9.14e-21
C1407 _325_/a_1270_373# _246_/B 1.04e-20
C1408 _331_/D _248_/A 2.32e-21
C1409 _325_/Q _232_/A 0.119f
C1410 _310_/a_27_7# _310_/a_448_7# -0.00297f
C1411 _323_/a_1108_7# _149_/A 4.88e-19
C1412 _248_/A _330_/a_193_7# 4.02e-20
C1413 _324_/a_761_249# _228_/A 9.27e-19
C1414 _196_/A _333_/D 3e-21
C1415 _281_/A _304_/X 0.00394f
C1416 _247_/a_113_257# _315_/a_27_7# 1.06e-19
C1417 _308_/X _178_/a_27_7# 5.17e-20
C1418 _219_/a_256_7# _330_/Q 0.00208f
C1419 _344_/a_1602_7# _158_/Y 5.14e-20
C1420 _258_/a_218_334# _147_/A 2.15e-19
C1421 _331_/D _331_/CLK 0.00469f
C1422 _188_/S _304_/S 0.0209f
C1423 _283_/A _153_/a_215_257# 2.31e-19
C1424 _316_/D _330_/a_27_7# 5.22e-21
C1425 _331_/CLK _330_/a_193_7# 0.108f
C1426 _209_/X _283_/A 6.64e-20
C1427 output41/a_27_7# valid 0.0129f
C1428 _216_/A _215_/A 2.34f
C1429 _228_/A _304_/X 0.00407f
C1430 _324_/a_1270_373# _286_/Y 1.39e-19
C1431 _318_/Q _316_/D 0.00791f
C1432 _340_/CLK _312_/a_1283_n19# 1.24e-20
C1433 _219_/a_250_257# VPWR 0.026f
C1434 _309_/a_761_249# _174_/a_27_257# 1.74e-19
C1435 _309_/a_193_7# _174_/a_109_257# 4.33e-21
C1436 _277_/Y _216_/A 0.0063f
C1437 repeater43/X _322_/a_543_7# 9.49e-20
C1438 _267_/B _311_/D 0.00656f
C1439 _342_/a_1217_7# _248_/A 1.15e-19
C1440 _347_/Q _284_/A 0.00544f
C1441 _192_/B _153_/B 1.61e-20
C1442 _339_/Q _311_/a_543_7# 3.73e-20
C1443 clkbuf_2_1_0_clk/A _306_/S 0.0118f
C1444 _161_/Y _345_/Q 0.0221f
C1445 _292_/A _164_/Y 0.335f
C1446 _255_/X _336_/a_193_7# 1.23e-21
C1447 result[6] _318_/a_805_7# 2.48e-20
C1448 clk _335_/a_1283_n19# 4.38e-20
C1449 _337_/a_543_7# _254_/B 1.11e-21
C1450 _188_/S _225_/X 2.85e-20
C1451 _345_/a_27_7# _166_/Y 5.64e-19
C1452 _307_/X _188_/S 0.0178f
C1453 _330_/D _331_/a_651_373# 1.4e-19
C1454 output26/a_27_7# VGND 0.106f
C1455 _176_/a_27_7# _343_/Q 0.0445f
C1456 _308_/a_505_n19# input1/X 0.0297f
C1457 _214_/a_27_257# _331_/a_27_7# 7.63e-19
C1458 _164_/Y _160_/A 0.0973f
C1459 _324_/Q VGND 1.36f
C1460 _167_/X _170_/a_489_373# 0.00277f
C1461 _250_/a_78_159# VPWR 0.035f
C1462 _324_/a_761_249# _216_/A 0.00106f
C1463 _321_/a_193_7# _234_/B 9.62e-20
C1464 _331_/D _222_/a_93_n19# 6.9e-20
C1465 _214_/a_109_7# _212_/X 5.98e-19
C1466 _343_/CLK _244_/B 0.0157f
C1467 _268_/a_39_257# _316_/a_193_7# 0.00269f
C1468 _160_/X _344_/D 5.23e-20
C1469 _216_/A _304_/X 0.238f
C1470 _251_/X _314_/a_193_7# 0.00107f
C1471 _342_/a_1283_n19# repeater43/X 0.012f
C1472 _236_/B _241_/a_113_257# 0.00766f
C1473 _346_/SET_B _147_/Y 0.426f
C1474 _346_/SET_B _312_/a_1108_7# 0.0208f
C1475 _340_/a_27_7# _194_/A 2.39e-20
C1476 _300_/Y _228_/A 0.00142f
C1477 _323_/D _343_/CLK 0.0317f
C1478 _346_/Q _160_/X 0.204f
C1479 _332_/a_27_7# _332_/a_1283_n19# -1.19e-19
C1480 _283_/Y _323_/Q 3.68e-20
C1481 _332_/a_193_7# _332_/a_543_7# -8.58e-19
C1482 _279_/Y _192_/a_150_257# 1.32e-19
C1483 _313_/Q _313_/a_543_7# 4.26e-19
C1484 _313_/D _313_/a_448_7# 0.00436f
C1485 _275_/Y cal 7.95e-21
C1486 _345_/a_193_7# _290_/A 0.0051f
C1487 _340_/a_193_7# _338_/a_27_7# 1.88e-21
C1488 _175_/Y _335_/Q 8.86e-22
C1489 _232_/X _331_/a_193_7# 9.2e-19
C1490 _217_/a_27_7# _214_/a_27_257# 2.95e-20
C1491 ctln[4] _306_/S 1.59e-20
C1492 _347_/a_27_7# _347_/a_448_7# -0.00346f
C1493 _347_/a_193_7# _347_/a_1108_7# -0.00656f
C1494 _294_/A clkbuf_2_1_0_clk/A 0.116f
C1495 _297_/B _284_/A 1.82e-19
C1496 _325_/Q _243_/a_199_7# 0.00183f
C1497 _340_/a_448_7# _196_/A 0.0245f
C1498 _261_/A _311_/a_193_7# 0.0158f
C1499 _267_/A _311_/a_761_249# 0.00456f
C1500 _269_/A _315_/a_651_373# 7.9e-19
C1501 _279_/Y _286_/B 0.00919f
C1502 _289_/a_121_257# _338_/Q 8.47e-19
C1503 _281_/Y _330_/Q 0.0304f
C1504 _323_/a_1217_7# _323_/Q 2.56e-19
C1505 _260_/B _181_/X 4.92e-20
C1506 _294_/A _310_/Q 0.00335f
C1507 output26/a_27_7# output27/a_27_7# 0.0246f
C1508 _277_/A _242_/A 0.586f
C1509 _305_/a_505_n19# _192_/B 4.03e-22
C1510 _232_/A _326_/Q 0.192f
C1511 _195_/a_27_257# VGND -0.00162f
C1512 _195_/a_109_7# VPWR -6.55e-19
C1513 _281_/A VGND 1.82f
C1514 _254_/Y _265_/B 1.13e-19
C1515 _324_/a_1283_n19# _306_/S 9.73e-21
C1516 _346_/a_652_n19# _162_/X 1.24e-19
C1517 clkbuf_0_clk/X _320_/a_27_7# 2.87e-22
C1518 _345_/D _172_/B 0.00121f
C1519 _323_/a_1283_n19# clk 5.43e-19
C1520 _281_/Y _324_/a_805_7# 2.96e-19
C1521 _272_/a_39_257# _216_/A 0.00496f
C1522 _294_/Y _284_/a_121_257# 1.05e-19
C1523 _216_/A _300_/Y 2.04e-20
C1524 output22/a_27_7# _341_/a_27_7# 0.00852f
C1525 _325_/a_543_7# _214_/a_27_257# 1.09e-21
C1526 _316_/a_27_7# _316_/a_193_7# -0.0576f
C1527 _279_/Y _256_/a_209_7# 2.79e-19
C1528 _326_/a_543_7# _181_/X 6.82e-19
C1529 _310_/a_27_7# _310_/D 0.485f
C1530 _228_/A VGND 2.58f
C1531 _281_/Y _314_/D 0.0104f
C1532 _308_/X _146_/a_29_271# 7.76e-20
C1533 _299_/X _328_/Q 1.01e-24
C1534 _229_/a_76_159# _176_/a_27_7# 4.69e-21
C1535 _329_/D _330_/Q 0.0299f
C1536 _336_/a_27_7# _336_/a_761_249# -0.0166f
C1537 _319_/Q VPWR 4.68f
C1538 _306_/X _147_/A 1.95e-19
C1539 _162_/a_27_7# _171_/a_78_159# 5.29e-20
C1540 _237_/a_199_7# _329_/Q 0.00161f
C1541 _197_/X _191_/B 2.28e-20
C1542 _168_/a_397_257# VGND -0.00343f
C1543 _207_/a_181_7# VGND 3.39e-19
C1544 clkbuf_2_1_0_clk/A _283_/A 7e-19
C1545 _248_/B _314_/a_27_7# 9.72e-20
C1546 output10/a_27_7# input4/a_27_7# 2.45e-20
C1547 _342_/a_1108_7# _226_/X 4.01e-19
C1548 _319_/Q _318_/a_543_7# 6.46e-22
C1549 _309_/a_1283_n19# _344_/Q 1e-19
C1550 _309_/a_193_7# _344_/D 6.54e-20
C1551 _154_/A _205_/a_79_n19# 4.15e-19
C1552 _346_/a_193_7# _299_/a_215_7# 1.84e-20
C1553 _346_/a_1182_221# _299_/a_78_159# 0.0013f
C1554 _206_/A _147_/Y 3.55e-19
C1555 _313_/a_761_249# _147_/Y 9.74e-20
C1556 output36/a_27_7# trimb[0] 0.00903f
C1557 output25/a_27_7# _317_/a_193_7# 2.37e-19
C1558 _342_/Q _227_/A 0.00882f
C1559 _333_/a_1270_373# _190_/A 1.44e-19
C1560 _323_/a_543_7# cal 0.00579f
C1561 _254_/Y _336_/a_1270_373# 5.43e-19
C1562 output21/a_27_7# _331_/CLK 1.33e-20
C1563 _144_/a_27_7# _227_/A 2.97e-20
C1564 _345_/a_586_7# _166_/Y 6.07e-20
C1565 _329_/a_27_7# _321_/Q 9.05e-23
C1566 _162_/X _173_/a_226_7# 1.3e-19
C1567 _258_/a_76_159# _202_/a_93_n19# 5.89e-19
C1568 _345_/a_193_7# _167_/a_27_257# 6.97e-20
C1569 _345_/a_27_7# _167_/a_109_257# 9.55e-20
C1570 _277_/Y _240_/a_109_257# 1.66e-19
C1571 repeater43/X _330_/a_1108_7# 0.0186f
C1572 _279_/Y _347_/a_543_7# 7.71e-19
C1573 _216_/A VGND 1.5f
C1574 _250_/X VPWR 0.526f
C1575 _294_/Y _262_/a_199_7# 1.43e-19
C1576 _331_/a_27_7# _330_/a_27_7# 9.42e-21
C1577 _332_/a_27_7# _208_/a_215_7# 7e-21
C1578 _332_/a_193_7# _208_/a_493_257# 1.16e-21
C1579 _331_/D _217_/X 1.16e-19
C1580 _290_/A VPWR 1.1f
C1581 _164_/Y _163_/a_493_257# 4.23e-19
C1582 _211_/a_27_257# _339_/D 4.1e-20
C1583 _197_/X _339_/a_805_7# 8.8e-20
C1584 output37/a_27_7# input2/a_27_7# 0.0109f
C1585 _292_/A _165_/a_78_159# 0.00737f
C1586 _345_/a_381_7# _167_/X 1.64e-21
C1587 _339_/D _198_/a_93_n19# 0.00235f
C1588 _318_/Q _331_/a_27_7# 8.22e-20
C1589 _251_/a_510_7# VGND -0.00222f
C1590 repeater43/X _333_/a_193_7# -0.00136f
C1591 _221_/a_584_7# VGND -7.84e-19
C1592 _341_/Q _335_/Q 1.07e-20
C1593 _329_/a_27_7# _297_/B 4.19e-21
C1594 _273_/A _164_/Y 0.101f
C1595 _275_/Y _284_/A 0.0097f
C1596 _338_/D _312_/D 0.0017f
C1597 _251_/X _324_/D 3.63e-19
C1598 ctln[4] _283_/A 2.3e-20
C1599 _322_/a_543_7# result[6] 0.00868f
C1600 _333_/a_1108_7# _206_/A 0.0581f
C1601 _333_/a_543_7# _207_/C 0.00202f
C1602 _290_/A _309_/a_27_7# 0.00507f
C1603 _254_/Y clkbuf_2_1_0_clk/A 0.00785f
C1604 _231_/a_512_7# _304_/S 0.00431f
C1605 output16/a_27_7# output38/a_27_7# 0.0246f
C1606 _232_/X _331_/a_1462_7# 3.67e-19
C1607 _290_/Y VGND 0.448f
C1608 rstn _154_/A 1.8e-20
C1609 _292_/A trim[3] 0.00641f
C1610 _147_/A _147_/Y 0.187f
C1611 _347_/a_27_7# _347_/D 0.0523f
C1612 _341_/D _177_/A 0.0056f
C1613 _181_/X _295_/a_512_7# 0.00807f
C1614 _172_/A _174_/a_109_257# 0.0262f
C1615 _336_/a_543_7# _336_/Q 3.15e-21
C1616 _318_/Q _217_/a_27_7# 0.0398f
C1617 _254_/Y _310_/Q 4.51e-20
C1618 _322_/Q _282_/a_121_257# 3.91e-19
C1619 _331_/Q _282_/a_39_257# 0.0101f
C1620 _343_/CLK _333_/a_448_7# 2.63e-20
C1621 _334_/Q _333_/a_193_7# 2.7e-19
C1622 _317_/Q _318_/D 1.44e-20
C1623 _157_/A _181_/a_27_7# 4.88e-20
C1624 _267_/B _312_/a_1283_n19# 5.37e-20
C1625 _197_/X _337_/Q 1.21f
C1626 _231_/a_409_7# _150_/C 0.00272f
C1627 _181_/X _333_/Q 2.44e-19
C1628 trim[4] _164_/Y 1.43e-19
C1629 _196_/A _190_/A 0.0735f
C1630 _227_/A _204_/Y 0.0482f
C1631 _288_/A _158_/Y 0.00113f
C1632 _269_/A _318_/a_27_7# 0.0178f
C1633 clkbuf_2_3_0_clk/A _263_/a_109_257# 0.0013f
C1634 _317_/a_651_373# _317_/D 0.00178f
C1635 _248_/A _298_/X 2.04e-20
C1636 _158_/Y _162_/X 0.0897f
C1637 _315_/a_193_7# _315_/a_761_249# -0.00517f
C1638 _315_/Q _341_/a_651_373# 2.2e-21
C1639 result[0] _341_/a_1108_7# 3.59e-19
C1640 _333_/a_193_7# _191_/B 0.486f
C1641 _329_/a_1283_n19# _218_/a_250_257# 4.95e-19
C1642 _218_/a_93_n19# _327_/D 0.00101f
C1643 _317_/Q _217_/A 0.0123f
C1644 _331_/Q _327_/Q 0.00403f
C1645 _294_/A _311_/a_27_7# 8.43e-22
C1646 _338_/a_761_249# _340_/CLK 0.0194f
C1647 _256_/a_303_7# _190_/A 0.00345f
C1648 _167_/a_27_257# VPWR 0.0981f
C1649 _325_/a_543_7# _318_/Q 4.7e-22
C1650 _247_/a_199_7# VPWR -1.13e-19
C1651 _169_/a_109_257# clkbuf_2_1_0_clk/A 0.00183f
C1652 _298_/C _295_/a_306_7# 9.39e-20
C1653 _346_/SET_B _347_/a_193_7# -0.00122f
C1654 _219_/a_93_n19# _232_/X 0.00684f
C1655 _324_/a_1283_n19# _248_/B 4.35e-20
C1656 _333_/a_1283_n19# _225_/X 4.89e-21
C1657 _162_/a_27_7# _172_/B 1.21e-20
C1658 _208_/a_78_159# _204_/a_27_257# 1.68e-19
C1659 _343_/a_639_7# _185_/A 0.00129f
C1660 _234_/B _242_/B 3.63e-20
C1661 _167_/a_109_7# _297_/B 0.00166f
C1662 _224_/a_93_n19# _298_/A 4.42e-20
C1663 _189_/a_27_7# VPWR 0.0951f
C1664 _342_/D _150_/C 1.47e-20
C1665 _321_/a_1283_n19# _242_/B 5.21e-20
C1666 _143_/a_27_7# _177_/A 5.73e-19
C1667 _286_/B _313_/a_27_7# 0.00413f
C1668 _343_/Q _333_/Q 9.41e-20
C1669 _258_/S output35/a_27_7# 3.43e-21
C1670 _255_/B VPWR 1.47f
C1671 result[3] _317_/a_448_7# 8.66e-20
C1672 _284_/a_39_257# _265_/B 9.07e-20
C1673 _340_/a_1283_n19# _340_/CLK 6.07e-20
C1674 _257_/a_79_159# VPWR 0.00835f
C1675 _341_/a_1283_n19# _341_/D 0.057f
C1676 _216_/X _347_/D 1.02e-20
C1677 _294_/Y VGND 0.254f
C1678 _329_/a_805_7# _330_/Q 1.8e-19
C1679 _153_/A _298_/A 5.06e-20
C1680 _258_/a_76_159# _284_/A 0.00147f
C1681 _331_/D _331_/a_805_7# 5.87e-19
C1682 _269_/A _246_/B 2.82e-20
C1683 _332_/a_1108_7# _332_/Q 0.00346f
C1684 _332_/a_1283_n19# _333_/Q 0.00367f
C1685 _332_/a_543_7# _190_/A 6.37e-21
C1686 _197_/X _339_/Q 0.143f
C1687 _162_/X _313_/a_651_373# 4.62e-20
C1688 _305_/a_505_n19# _260_/A 0.00172f
C1689 _328_/a_651_373# _329_/Q 0.00272f
C1690 _328_/a_1108_7# _238_/B 0.00251f
C1691 _317_/Q _272_/a_121_257# 1.81e-21
C1692 _307_/a_505_n19# _196_/A 2.9e-20
C1693 repeater43/X _333_/a_1462_7# -9.14e-19
C1694 _329_/a_651_373# VGND 4.27e-19
C1695 _329_/a_639_7# VPWR 5.2e-19
C1696 _338_/a_543_7# _346_/SET_B 0.0269f
C1697 _338_/a_1283_n19# _338_/D 0.0497f
C1698 _338_/a_27_7# _338_/Q 2.3e-20
C1699 _180_/a_183_257# _298_/C 5.51e-19
C1700 _244_/B output30/a_27_7# 0.00141f
C1701 _244_/a_109_257# _286_/Y 0.00122f
C1702 _197_/X _202_/a_256_7# 5.4e-19
C1703 _310_/a_27_7# VPWR 0.117f
C1704 _240_/a_109_257# VGND -2.85e-19
C1705 _325_/Q _245_/a_113_257# 2.22e-19
C1706 _289_/a_39_257# _337_/Q 1.62e-20
C1707 _306_/a_218_7# _306_/S 4.94e-20
C1708 _344_/a_1182_221# _344_/Q 0.0276f
C1709 _344_/a_193_7# _344_/D 0.0498f
C1710 _341_/a_448_7# _248_/A 0.00239f
C1711 _342_/a_448_7# cal 1.34e-19
C1712 _342_/a_1108_7# input1/X 0.0017f
C1713 _182_/a_79_n19# _192_/B 0.02f
C1714 _196_/A _178_/a_27_7# 0.00193f
C1715 _316_/Q _269_/A 0.063f
C1716 _294_/A _309_/a_1283_n19# 0.057f
C1717 _343_/CLK _177_/A 0.0025f
C1718 _326_/D _325_/D 5.23e-20
C1719 _290_/A _309_/a_1217_7# 1.61e-19
C1720 repeater43/X _268_/a_39_257# 0.0113f
C1721 _271_/Y _269_/A 0.101f
C1722 _340_/a_1108_7# _346_/SET_B -0.00722f
C1723 _323_/D output30/a_27_7# 0.00245f
C1724 _273_/A _165_/a_78_159# 8.94e-19
C1725 _227_/A _225_/B 2.33e-20
C1726 _332_/a_27_7# _206_/A 8.51e-19
C1727 _172_/A _344_/D 0.00604f
C1728 _260_/B _346_/SET_B 2.09e-19
C1729 _330_/Q _242_/A 5.89e-19
C1730 _309_/a_27_7# _310_/a_27_7# 5.85e-19
C1731 _343_/CLK _333_/D 9.83e-19
C1732 _172_/A _346_/Q 1.3e-19
C1733 _271_/A _270_/a_121_257# 4.47e-19
C1734 _327_/a_543_7# _346_/SET_B 0.0289f
C1735 _324_/a_27_7# _326_/Q 9.43e-19
C1736 output23/a_27_7# _248_/B 7.66e-20
C1737 _308_/S _255_/a_30_13# 8.82e-19
C1738 _346_/a_27_7# _346_/a_193_7# -0.0853f
C1739 _288_/A _160_/a_27_7# 2.88e-20
C1740 _343_/CLK _332_/a_193_7# 4.37e-20
C1741 _339_/Q _312_/a_193_7# 0.00107f
C1742 _271_/Y _343_/D 7.27e-20
C1743 _316_/a_651_373# _248_/A 9.07e-20
C1744 _251_/a_79_n19# _181_/a_27_7# 0.0115f
C1745 _340_/CLK _190_/a_27_7# 0.00114f
C1746 _343_/a_1108_7# _175_/Y 0.0654f
C1747 _185_/A _184_/a_76_159# 0.00224f
C1748 _162_/X _160_/a_27_7# 6.28e-19
C1749 input4/X _338_/a_193_7# 9.6e-19
C1750 _340_/a_27_7# _339_/a_27_7# 5.3e-19
C1751 _325_/Q VPWR 0.278f
C1752 _216_/A _214_/a_27_257# 1.19e-20
C1753 _286_/B _144_/A 1.59e-20
C1754 _342_/a_543_7# sample 0.00102f
C1755 _342_/a_1108_7# _286_/Y 4.62e-21
C1756 trim[3] _273_/A 0.00465f
C1757 _292_/A _273_/Y 0.0262f
C1758 _242_/A _318_/a_761_249# 0.012f
C1759 _320_/a_27_7# _328_/Q 3.61e-19
C1760 _316_/a_448_7# _316_/D 0.00196f
C1761 _344_/a_27_7# _290_/A 0.00317f
C1762 _294_/A _306_/a_218_7# 0.00191f
C1763 _318_/Q output26/a_27_7# 5.55e-20
C1764 _161_/Y _284_/A 2.68e-20
C1765 _298_/a_27_7# VPWR 0.0366f
C1766 _329_/a_543_7# _330_/D 0.00995f
C1767 clkbuf_2_3_0_clk/A _312_/Q 3.53e-21
C1768 en _227_/A 0.00643f
C1769 _298_/C _226_/a_79_n19# 1.87e-19
C1770 output39/a_27_7# trimb[3] 0.00995f
C1771 ctln[5] _333_/Q 3.38e-20
C1772 _301_/a_240_7# VGND -0.00443f
C1773 _328_/a_761_249# _346_/SET_B -0.00735f
C1774 _346_/SET_B _347_/a_1462_7# 8.79e-19
C1775 _289_/a_39_257# _339_/Q 3.99e-19
C1776 _326_/a_448_7# _248_/A 5.98e-21
C1777 _334_/a_193_7# _334_/a_651_373# -0.00701f
C1778 input1/X _312_/a_761_249# 3.54e-20
C1779 clkbuf_2_1_0_clk/A _194_/a_27_7# 0.00219f
C1780 _181_/X _212_/X 0.531f
C1781 _293_/a_39_257# _306_/S 0.00541f
C1782 _200_/a_346_7# _338_/Q 0.00232f
C1783 _204_/a_27_257# _190_/A 1.37e-20
C1784 clk _333_/a_1283_n19# 0.0136f
C1785 _327_/a_448_7# _331_/CLK 0.0165f
C1786 _274_/a_39_257# _347_/D 1.25e-19
C1787 _208_/a_215_7# _333_/Q 2.12e-19
C1788 output36/a_27_7# VPWR 0.136f
C1789 _343_/a_761_249# _298_/A 6.19e-20
C1790 _329_/a_1108_7# _328_/D 7.62e-19
C1791 _255_/B _184_/a_505_n19# 7.75e-21
C1792 _217_/A _298_/A 7.68e-19
C1793 _326_/a_448_7# _331_/CLK 4.31e-19
C1794 _326_/a_1108_7# _316_/D 1.08e-19
C1795 _326_/a_1283_n19# _236_/B 2.16e-19
C1796 _172_/B _286_/Y 1.34e-19
C1797 repeater43/X _316_/a_27_7# 0.0115f
C1798 _341_/a_1283_n19# _343_/CLK 1.24e-19
C1799 _258_/S _313_/a_1283_n19# 1.76e-20
C1800 output11/a_27_7# input4/X 4.04e-19
C1801 _147_/A _347_/a_193_7# 0.00125f
C1802 _286_/B _313_/a_1217_7# 1.07e-19
C1803 _321_/a_1108_7# VPWR 0.0306f
C1804 _321_/a_543_7# VGND 6.8e-20
C1805 _283_/Y _194_/X 0.0327f
C1806 _338_/a_1283_n19# _343_/CLK 5.12e-19
C1807 result[5] _269_/A 8.18e-19
C1808 _169_/Y _347_/Q 0.0111f
C1809 _325_/a_1108_7# _223_/a_250_257# 8.7e-20
C1810 _234_/B _318_/a_1283_n19# 8.53e-20
C1811 _313_/D _336_/D 2.46e-19
C1812 clkbuf_2_1_0_clk/a_75_172# _242_/A 3.56e-19
C1813 _153_/a_297_257# VPWR -0.0029f
C1814 _153_/a_109_53# VGND -0.00326f
C1815 _224_/a_93_n19# _304_/X 0.0669f
C1816 _340_/CLK _332_/Q 0.00548f
C1817 _340_/a_651_373# _337_/a_1283_n19# 8.38e-19
C1818 _340_/a_1283_n19# _337_/a_651_373# 8.38e-19
C1819 _267_/A _312_/a_27_7# 0.00271f
C1820 _326_/a_1283_n19# _326_/D 9.29e-21
C1821 _296_/Y _196_/A 8.44e-20
C1822 _145_/A _286_/B 0.00891f
C1823 _275_/Y _310_/a_761_249# 0.00136f
C1824 _290_/A _171_/a_215_7# 1.26e-19
C1825 _287_/a_121_257# _337_/Q 4.96e-19
C1826 _305_/a_76_159# _306_/S 1.22e-20
C1827 _274_/a_121_257# _346_/SET_B 2.06e-19
C1828 _238_/B _319_/a_651_373# 0.00145f
C1829 _281_/A _330_/a_27_7# 0.00628f
C1830 _197_/X _336_/D 0.00403f
C1831 _310_/a_1217_7# VPWR 1.7e-19
C1832 output22/a_27_7# repeater43/X 0.00527f
C1833 _318_/Q _281_/A 1.44e-20
C1834 _165_/a_215_7# _158_/Y 0.0118f
C1835 _341_/D _248_/A 0.0103f
C1836 _342_/D cal 3.95e-19
C1837 _182_/X _192_/B 0.00211f
C1838 _275_/Y _264_/a_113_257# 0.00712f
C1839 _294_/A _293_/a_39_257# 0.00495f
C1840 _296_/Y _304_/a_591_329# 1.27e-19
C1841 _343_/CLK _208_/a_78_159# 0.00115f
C1842 _216_/X _304_/S 0.0984f
C1843 _346_/a_1182_221# _346_/SET_B 0.0632f
C1844 _216_/A _203_/a_209_257# 5.07e-20
C1845 _271_/A _175_/Y 0.0112f
C1846 _346_/a_193_7# _275_/A 2.46e-21
C1847 _271_/A _243_/a_113_257# 0.0063f
C1848 clkbuf_0_clk/a_110_7# _196_/A 0.00195f
C1849 _325_/a_193_7# _181_/X 0.016f
C1850 _169_/B VPWR 0.0182f
C1851 _209_/a_109_7# VPWR -5.45e-19
C1852 _209_/a_27_257# VGND -0.00707f
C1853 _347_/Q _314_/a_543_7# 2.97e-20
C1854 _339_/a_543_7# _338_/a_448_7# 2.45e-19
C1855 input4/X _334_/a_27_7# 0.0116f
C1856 trim[0] output5/a_27_7# 7.65e-22
C1857 _337_/a_193_7# _340_/CLK 0.0273f
C1858 _272_/a_39_257# _224_/a_93_n19# 4.23e-20
C1859 _335_/a_1283_n19# _335_/Q 0.0415f
C1860 _335_/a_543_7# _204_/Y 1.49e-19
C1861 _169_/Y _297_/B 6.5e-20
C1862 _297_/B _225_/B 1.67e-19
C1863 _326_/Q VPWR 0.553f
C1864 _160_/X _170_/a_76_159# 0.0456f
C1865 _324_/a_543_7# _215_/A 1.73e-19
C1866 _319_/a_27_7# _319_/a_193_7# -9.38e-20
C1867 _324_/a_1217_7# _326_/Q 6.2e-20
C1868 _325_/a_1108_7# _304_/a_79_n19# 2.87e-19
C1869 _309_/Q _310_/D 3.75e-20
C1870 _346_/a_193_7# _346_/a_586_7# -7.91e-19
C1871 repeater43/X _341_/a_805_7# -0.00125f
C1872 _266_/a_199_7# _310_/Q 3.06e-20
C1873 _236_/B _248_/A 0.262f
C1874 _309_/a_193_7# _265_/B 0.0113f
C1875 _260_/B _147_/A 0.049f
C1876 _298_/C _323_/Q 0.00835f
C1877 _185_/A _188_/S 8.11e-19
C1878 _334_/a_761_249# _206_/A 3.77e-21
C1879 _334_/a_27_7# _207_/C 0.223f
C1880 _181_/a_27_7# _296_/a_213_83# 1.99e-19
C1881 cal _263_/B 0.00317f
C1882 _236_/a_109_257# _321_/D 7e-20
C1883 _236_/B _331_/CLK 4.64e-19
C1884 _315_/a_761_249# VGND 0.00247f
C1885 _315_/a_1283_n19# VPWR 0.024f
C1886 clkbuf_2_1_0_clk/A _160_/X 0.0128f
C1887 _227_/A _315_/D 0.0113f
C1888 input3/a_27_7# VGND 0.0712f
C1889 output39/a_27_7# VPWR 0.131f
C1890 _318_/Q _216_/A 6.04e-21
C1891 _336_/a_639_7# VPWR 2.35e-19
C1892 _324_/a_651_373# _227_/A 0.00687f
C1893 _336_/a_651_373# VGND 0.0032f
C1894 _317_/a_761_249# _316_/a_193_7# 1.6e-19
C1895 _324_/a_193_7# _324_/a_1283_n19# -7.59e-20
C1896 _277_/Y _346_/D 3.28e-21
C1897 _326_/D _248_/A 0.0187f
C1898 _334_/a_543_7# _343_/CLK 1.58e-20
C1899 _334_/a_761_249# _334_/D 0.043f
C1900 repeater43/X _229_/a_226_257# 2.74e-19
C1901 _315_/D _314_/a_1108_7# 0.00873f
C1902 _314_/a_193_7# VPWR 0.0571f
C1903 _346_/SET_B _319_/a_1283_n19# -0.00597f
C1904 _338_/D _337_/a_543_7# 4.55e-20
C1905 _346_/SET_B _337_/a_761_249# -7.09e-19
C1906 _275_/A _319_/a_193_7# 2.12e-20
C1907 _326_/D _331_/CLK 0.00276f
C1908 _224_/a_93_n19# VGND 0.0351f
C1909 _224_/a_256_7# VPWR -7.75e-19
C1910 _193_/Y _254_/B 0.174f
C1911 _216_/X _331_/a_543_7# 4.87e-20
C1912 repeater43/X _316_/a_1217_7# -3.08e-19
C1913 _300_/a_735_7# _160_/X 1.12e-19
C1914 _324_/a_27_7# _324_/D 0.477f
C1915 _324_/a_543_7# _304_/X 2.81e-19
C1916 _314_/a_543_7# _297_/B 0.00835f
C1917 _314_/a_761_249# _314_/D 2.33e-20
C1918 _311_/D _310_/a_193_7# 5.37e-19
C1919 _311_/a_193_7# _310_/D 1.58e-21
C1920 _286_/B _174_/a_27_257# 0.00198f
C1921 _170_/a_226_7# VPWR -0.00385f
C1922 _273_/A _273_/Y 0.0899f
C1923 _322_/a_1283_n19# _269_/A 6.19e-20
C1924 _341_/a_1108_7# _145_/A 0.00368f
C1925 input4/X _207_/X 9.16e-20
C1926 _325_/a_1283_n19# _325_/D 0.058f
C1927 _339_/a_27_7# _332_/D 1.69e-20
C1928 _339_/a_193_7# _340_/CLK 0.0249f
C1929 _326_/D _273_/A 0.0264f
C1930 rstn _153_/B 0.0814f
C1931 _323_/a_27_7# _175_/Y 7.14e-19
C1932 _154_/A VPWR 1.24f
C1933 _153_/A VGND 0.745f
C1934 _304_/X _217_/A 0.568f
C1935 _340_/a_193_7# _337_/Q 0.0118f
C1936 _340_/a_1108_7# _337_/D 3.99e-20
C1937 _327_/a_1270_373# _327_/Q 5.8e-20
C1938 _327_/a_651_373# _212_/X 0.00387f
C1939 _326_/a_805_7# repeater43/X 0.00128f
C1940 _247_/a_113_257# _244_/B 0.00778f
C1941 _343_/CLK _248_/A 0.0248f
C1942 _288_/A _267_/A 0.00655f
C1943 _326_/a_27_7# _331_/a_1108_7# 3.29e-21
C1944 _326_/a_193_7# _331_/a_1283_n19# 8.23e-20
C1945 _206_/A _333_/Q 0.254f
C1946 clkbuf_2_3_0_clk/A _340_/CLK 0.0518f
C1947 _207_/X _207_/C 0.472f
C1948 _326_/a_448_7# _217_/X 0.0162f
C1949 _326_/D _222_/a_93_n19# 0.00312f
C1950 _293_/a_39_257# _254_/Y 0.0255f
C1951 _271_/A _341_/Q 0.618f
C1952 _162_/X _267_/A 1.07e-19
C1953 _343_/CLK _331_/CLK 3.06e-21
C1954 _182_/X _146_/C 7.36e-19
C1955 _346_/a_193_7# _254_/A 7.31e-20
C1956 _345_/a_193_7# _345_/a_1602_7# -4.7e-21
C1957 _345_/a_27_7# _345_/a_381_7# -0.00438f
C1958 _347_/Q _315_/D 4.77e-20
C1959 _222_/a_93_n19# _222_/a_256_7# -3.48e-20
C1960 _334_/D _333_/Q 1.45e-19
C1961 _343_/CLK _190_/A 0.0174f
C1962 _275_/Y _169_/Y 1.01e-20
C1963 _300_/a_383_7# VGND 0.00129f
C1964 _281_/Y _333_/a_1283_n19# 1.01e-19
C1965 _328_/a_448_7# _212_/X 0.0228f
C1966 _308_/a_76_159# _227_/A 0.0522f
C1967 _327_/Q _347_/D -1.01e-24
C1968 _301_/X _347_/a_27_7# 2.46e-20
C1969 _324_/Q _286_/B 0.0451f
C1970 _191_/B _295_/a_79_n19# 8.18e-20
C1971 _346_/a_1296_7# _346_/SET_B 6.78e-19
C1972 _309_/a_193_7# clkbuf_2_1_0_clk/A 2.12e-21
C1973 _177_/a_27_7# _286_/Y 8.85e-20
C1974 _290_/A _147_/Y 1.97e-20
C1975 _322_/a_193_7# _321_/a_27_7# 9.14e-20
C1976 _173_/a_76_159# _345_/D 0.00316f
C1977 _173_/a_226_7# _345_/Q 0.0266f
C1978 _266_/a_113_257# _309_/Q 8.06e-19
C1979 _339_/a_543_7# _338_/D 0.00877f
C1980 _339_/a_761_249# _346_/SET_B -0.00113f
C1981 _290_/A _312_/a_1108_7# 0.00312f
C1982 repeater43/X _334_/a_639_7# -1.78e-19
C1983 _194_/A _202_/a_93_n19# 0.0559f
C1984 _326_/a_1108_7# _217_/a_27_7# 0.00173f
C1985 result[1] _315_/a_1108_7# 5.16e-19
C1986 _309_/a_1108_7# _310_/D 0.00622f
C1987 _309_/a_193_7# _310_/Q 7.61e-20
C1988 _337_/a_1462_7# _340_/CLK 0.00188f
C1989 _258_/a_76_159# _336_/a_27_7# 3.28e-20
C1990 _272_/a_39_257# _217_/A 0.00578f
C1991 _324_/Q _304_/a_306_329# 2.59e-19
C1992 _300_/Y _346_/D 1.18e-20
C1993 clk _216_/X 1.18e-21
C1994 _164_/A _344_/D 1.27e-19
C1995 _263_/B _284_/A 2.67e-20
C1996 _254_/Y _305_/a_76_159# 4.41e-19
C1997 cal _194_/A 0.0101f
C1998 _258_/S _202_/a_93_n19# 2.94e-20
C1999 _345_/a_1032_373# _160_/X 0.012f
C2000 _337_/a_193_7# _337_/a_651_373# -0.00504f
C2001 _344_/a_1140_373# _297_/Y 0.00155f
C2002 _215_/A _314_/Q 4.53e-21
C2003 _235_/a_199_7# VPWR -2.56e-19
C2004 _225_/X _332_/Q 1e-19
C2005 result[0] _145_/A 2.18e-20
C2006 _227_/A _335_/a_193_7# 6.84e-20
C2007 _242_/A _212_/a_27_7# 1.57e-19
C2008 _334_/a_1217_7# _207_/C 8.12e-19
C2009 _197_/a_27_7# _194_/A 3.06e-19
C2010 _327_/a_27_7# clkbuf_0_clk/X 0.178f
C2011 _318_/D VGND 0.0197f
C2012 _149_/A _333_/Q 1.38e-21
C2013 _258_/S cal 1.75e-20
C2014 _346_/SET_B _212_/X 0.717f
C2015 output6/a_27_7# _269_/Y 0.0188f
C2016 _324_/a_1108_7# VPWR 0.00338f
C2017 _324_/a_543_7# VGND 0.00217f
C2018 _180_/a_29_13# _191_/B 8.46e-19
C2019 _342_/a_448_7# _342_/Q 7.3e-22
C2020 _340_/CLK _192_/B 1.14e-20
C2021 _306_/a_505_n19# clkbuf_2_1_0_clk/A 6.71e-19
C2022 _315_/D _297_/B 0.0621f
C2023 _318_/a_651_373# _242_/B 2.1e-20
C2024 _318_/a_1108_7# _318_/D 8.95e-20
C2025 _285_/A _265_/B 0.00856f
C2026 _234_/B _232_/X 0.00168f
C2027 _314_/a_805_7# VGND -7.01e-19
C2028 _314_/a_1462_7# VPWR 3.65e-19
C2029 _321_/a_1283_n19# _232_/X 0.0115f
C2030 _248_/A _331_/a_193_7# 2.67e-20
C2031 _346_/SET_B _313_/a_639_7# 0.00102f
C2032 _344_/a_1224_7# comp 4.04e-22
C2033 _343_/a_1283_n19# VPWR 0.0402f
C2034 _343_/a_761_249# VGND 0.0061f
C2035 _216_/a_27_7# _304_/S 0.00105f
C2036 _144_/A _316_/D 2.3e-19
C2037 _340_/a_543_7# cal 1.09e-20
C2038 _338_/a_805_7# _337_/Q 6.56e-21
C2039 _172_/A _209_/X 1.89e-21
C2040 _272_/a_39_257# _272_/a_121_257# 8.88e-34
C2041 _217_/A VGND 0.341f
C2042 _324_/D VPWR 0.412f
C2043 _317_/Q _317_/D 0.0216f
C2044 result[2] _244_/B 1.31e-19
C2045 output20/a_27_7# VPWR 0.0854f
C2046 input4/X _339_/a_27_7# 1.63e-20
C2047 _254_/B _205_/a_297_7# 1.94e-19
C2048 _344_/a_193_7# _265_/B 1.61e-20
C2049 _331_/CLK _331_/a_193_7# 0.0054f
C2050 _346_/D VGND 0.172f
C2051 _216_/A _223_/a_346_7# 1.05e-19
C2052 _236_/B _217_/X 1.28e-20
C2053 _293_/a_39_257# _336_/a_1108_7# 7.75e-20
C2054 _276_/a_68_257# _238_/B 7.41e-20
C2055 _341_/a_27_7# _286_/Y 0.502f
C2056 _286_/B _228_/A 0.00813f
C2057 _278_/a_150_257# VPWR -4.42e-19
C2058 _345_/a_1602_7# VPWR 0.0047f
C2059 _345_/a_1182_221# VGND 0.00166f
C2060 _158_/Y _345_/Q 0.0154f
C2061 _323_/a_1217_7# _175_/Y 6.96e-20
C2062 _273_/A _331_/a_193_7# 4.53e-22
C2063 _167_/a_27_257# _147_/Y 2.91e-19
C2064 _309_/Q VPWR 0.429f
C2065 output20/a_27_7# ctlp[6] 0.00862f
C2066 _340_/a_1462_7# _337_/Q 1.92e-19
C2067 _283_/A _330_/a_761_249# 0.00109f
C2068 _261_/A _312_/Q 0.0059f
C2069 _172_/A _265_/B 0.00392f
C2070 clk _334_/a_193_7# 0.00887f
C2071 _186_/a_79_n19# _341_/Q 3.39e-19
C2072 _220_/a_93_n19# _220_/a_250_257# -6.97e-22
C2073 _168_/a_397_257# _286_/B 3.77e-20
C2074 _339_/a_543_7# _337_/a_1108_7# 0.00203f
C2075 _339_/a_1108_7# _337_/a_543_7# 0.00203f
C2076 _330_/Q _218_/a_256_7# 5.44e-19
C2077 _307_/a_76_159# _147_/A 0.0403f
C2078 _326_/D _217_/X 0.0208f
C2079 _279_/A VPWR 0.497f
C2080 _277_/A _238_/a_109_257# 3.99e-19
C2081 _339_/a_543_7# _343_/CLK 1.66e-21
C2082 _323_/a_193_7# _227_/A 3.71e-20
C2083 _257_/a_79_159# _147_/Y 5.03e-21
C2084 _222_/a_346_7# _212_/X 0.00311f
C2085 _222_/a_584_7# _327_/Q 0.00295f
C2086 _218_/a_250_257# VPWR 0.0468f
C2087 _167_/X _162_/X 0.0409f
C2088 _272_/a_121_257# VGND 4.94e-20
C2089 _145_/A _316_/D 4.74e-21
C2090 _309_/a_27_7# _309_/Q -1.85e-21
C2091 _308_/S _227_/A 0.161f
C2092 _312_/a_1283_n19# _297_/Y 0.00125f
C2093 _286_/B _216_/A 0.372f
C2094 _260_/A _347_/a_448_7# 1.44e-20
C2095 _322_/a_448_7# _322_/D 0.00243f
C2096 _319_/a_651_373# _217_/X 8.15e-22
C2097 _300_/Y _314_/Q 7.68e-19
C2098 _294_/Y output40/a_27_7# 0.012f
C2099 _294_/Y output32/a_27_7# 0.00762f
C2100 _226_/a_382_257# _225_/X 0.00167f
C2101 _226_/a_297_7# _147_/A 0.00905f
C2102 _226_/a_79_n19# _150_/C 8.33e-19
C2103 _220_/a_346_7# VPWR -4.56e-19
C2104 _320_/Q _219_/a_346_7# 2.71e-21
C2105 _220_/a_250_257# VGND -0.00482f
C2106 _251_/a_297_257# _181_/X 2.33e-20
C2107 _311_/a_193_7# VPWR 0.0745f
C2108 _327_/a_27_7# _286_/Y 1.81e-20
C2109 _194_/A _284_/A 0.0574f
C2110 cal _334_/a_27_7# 0.00153f
C2111 _271_/A _330_/Q 1.03e-19
C2112 _325_/a_1283_n19# _248_/A 2.07e-19
C2113 _313_/D _336_/a_761_249# 5.37e-19
C2114 clk _295_/a_409_7# 1.53e-19
C2115 _327_/a_1283_n19# _219_/a_93_n19# 0.00457f
C2116 _308_/X _298_/A 0.00482f
C2117 repeater42/a_27_7# _218_/a_93_n19# 0.00123f
C2118 _346_/a_193_7# clkbuf_0_clk/X 1.95e-19
C2119 _342_/a_27_7# _298_/A 6.44e-20
C2120 _279_/Y _324_/Q 1.43e-20
C2121 _292_/Y output17/a_27_7# 8.5e-19
C2122 _325_/a_1283_n19# _331_/CLK 3.58e-21
C2123 _271_/A _269_/Y 5.23e-20
C2124 _318_/Q _321_/a_543_7# 1.63e-19
C2125 _146_/a_29_271# _143_/a_27_7# 1.84e-20
C2126 _258_/S _284_/A 1.19f
C2127 _337_/a_761_249# _337_/D 5.97e-19
C2128 _200_/a_250_257# _267_/A 1.44e-19
C2129 _323_/a_1108_7# _154_/A 8.81e-22
C2130 _165_/X _299_/a_292_257# 4.86e-19
C2131 clk _332_/Q 0.159f
C2132 _197_/X _336_/a_761_249# 9.14e-19
C2133 _320_/a_1283_n19# clkbuf_2_1_0_clk/A 3.58e-20
C2134 output9/a_27_7# VPWR 0.157f
C2135 _293_/a_39_257# _194_/a_27_7# 0.00969f
C2136 input4/X _323_/Q 3e-19
C2137 _317_/a_639_7# _248_/A 1.69e-19
C2138 _304_/S _327_/Q 2.14e-19
C2139 _332_/a_1283_n19# _207_/a_27_7# 0.00319f
C2140 _255_/B _333_/a_1108_7# 1.91e-20
C2141 _285_/A _310_/Q 3.08e-20
C2142 _327_/a_1217_7# clkbuf_0_clk/X 1.32e-19
C2143 _322_/Q _283_/A 0.0322f
C2144 _271_/A _318_/a_761_249# 2.37e-19
C2145 _344_/a_193_7# clkbuf_2_1_0_clk/A 4.28e-21
C2146 _328_/a_761_249# _219_/a_250_257# 0.00122f
C2147 _273_/A _325_/a_1283_n19# 1.54e-19
C2148 _340_/a_193_7# _336_/D 3e-21
C2149 _342_/D _342_/Q 0.252f
C2150 _289_/a_39_257# _310_/a_1283_n19# 0.00114f
C2151 repeater43/X _226_/X 0.0106f
C2152 _169_/Y _161_/Y 3.88e-20
C2153 _344_/a_1032_373# _310_/D 4.41e-20
C2154 _314_/Q VGND 0.361f
C2155 clkbuf_2_3_0_clk/A _267_/B 0.00343f
C2156 _318_/a_1270_373# VPWR -1.47e-19
C2157 _318_/a_448_7# VGND 6.39e-19
C2158 _341_/a_1108_7# _228_/A 4.15e-20
C2159 _196_/A _193_/Y 1.61e-19
C2160 _323_/Q _207_/C 3.93e-19
C2161 _157_/A _340_/CLK 7.58e-20
C2162 _181_/X _306_/S 0.0414f
C2163 _325_/a_543_7# _222_/a_250_257# 1.91e-20
C2164 _338_/Q _337_/Q 0.0434f
C2165 _157_/A _347_/D 5.93e-19
C2166 _172_/A clkbuf_2_1_0_clk/A 0.121f
C2167 _276_/a_68_257# _331_/CLK 0.0135f
C2168 _346_/a_476_7# _301_/X 1.43e-19
C2169 _211_/a_27_257# _154_/A 1.22e-19
C2170 _292_/A _344_/D 3.46e-20
C2171 _321_/a_1283_n19# _241_/a_113_257# 7.41e-21
C2172 _309_/a_1108_7# VPWR 0.0136f
C2173 _309_/a_543_7# VGND 0.0135f
C2174 _313_/a_639_7# _147_/A 0.005f
C2175 _331_/Q _232_/A 1.68e-21
C2176 repeater43/X _317_/a_761_249# 0.02f
C2177 _306_/a_218_7# _160_/X 2.07e-20
C2178 _340_/a_27_7# _194_/X 2.17e-19
C2179 clkbuf_0_clk/X _319_/a_193_7# 1.09e-19
C2180 _345_/a_1296_7# VGND 1.31e-19
C2181 _160_/a_27_7# _345_/Q 3.29e-20
C2182 _269_/A _177_/a_27_7# 0.00388f
C2183 cal _201_/a_27_7# 0.0208f
C2184 _279_/Y _195_/a_27_257# 1.66e-19
C2185 _254_/B _298_/A 0.0882f
C2186 _315_/a_193_7# _317_/D 0.0121f
C2187 _160_/A _344_/D 0.0021f
C2188 _317_/D _298_/A 0.152f
C2189 _281_/Y _216_/X 1.42f
C2190 _316_/Q _246_/B 0.0124f
C2191 _197_/X _199_/a_346_7# 6.45e-19
C2192 _322_/D _233_/a_113_257# 1.09e-20
C2193 clk _334_/a_1462_7# 1.31e-19
C2194 _313_/Q _336_/Q 0.0146f
C2195 _164_/Y comp 2.82e-20
C2196 _321_/a_193_7# _322_/Q 0.00527f
C2197 _321_/a_27_7# _331_/Q 2.9e-21
C2198 _326_/D _331_/a_805_7# 1.19e-20
C2199 repeater43/X _331_/a_1108_7# -8.77e-19
C2200 _281_/Y _329_/Q 6.21e-20
C2201 _330_/Q _330_/D 0.0132f
C2202 _283_/A _333_/a_639_7# 0.00447f
C2203 _279_/Y _228_/A 0.0103f
C2204 _324_/a_27_7# _181_/a_27_7# 3.29e-21
C2205 _229_/a_489_373# sample 5.6e-20
C2206 _248_/A output30/a_27_7# 0.00141f
C2207 _301_/a_51_257# _162_/X 0.0295f
C2208 _331_/a_193_7# _217_/X 3.48e-19
C2209 _331_/a_761_249# _212_/X 6.57e-20
C2210 _219_/a_93_n19# _248_/A 6.81e-20
C2211 _325_/a_27_7# _304_/S 3.66e-19
C2212 _346_/a_193_7# _286_/Y 4.52e-21
C2213 _183_/a_553_257# _178_/a_27_7# 9.5e-21
C2214 _333_/a_1283_n19# _335_/Q 5.81e-19
C2215 _192_/B _225_/X 0.00713f
C2216 _188_/a_505_n19# _146_/C 5.01e-19
C2217 _307_/X _192_/B 1.56e-20
C2218 _260_/A _340_/CLK 0.2f
C2219 _329_/D _216_/X 0.223f
C2220 _276_/a_68_257# _319_/a_1108_7# 9.99e-20
C2221 _275_/Y _311_/a_543_7# 5.9e-19
C2222 _219_/a_93_n19# _331_/CLK 1.61e-20
C2223 _340_/D _332_/a_193_7# 6.28e-21
C2224 cal _337_/a_27_7# 9.25e-19
C2225 _343_/a_1283_n19# _323_/a_1108_7# 5.48e-20
C2226 _343_/a_1108_7# _323_/a_1283_n19# 1.78e-21
C2227 _343_/a_651_373# _323_/a_761_249# 1.61e-20
C2228 _255_/B _304_/a_79_n19# 1.35e-19
C2229 _306_/a_439_7# VPWR -3.62e-19
C2230 trim[1] clkc 0.00909f
C2231 _306_/a_535_334# VGND -2.3e-19
C2232 _200_/a_250_257# _194_/X 0.00701f
C2233 _339_/Q _338_/Q 0.145f
C2234 _200_/a_93_n19# _340_/Q 0.0138f
C2235 _329_/Q _329_/D 0.0215f
C2236 _269_/A _268_/a_121_257# 3.75e-19
C2237 _181_/X _327_/D 7.39e-20
C2238 _311_/a_1462_7# VPWR 4.21e-19
C2239 _256_/a_80_n19# _255_/B 2.15e-19
C2240 _263_/B _310_/a_761_249# 1.24e-20
C2241 _242_/A _223_/a_93_n19# 2.22e-20
C2242 _145_/A _144_/A 3.63e-20
C2243 cal _334_/a_1217_7# 2.97e-20
C2244 _313_/Q _336_/a_805_7# 2.46e-21
C2245 _327_/a_761_249# _329_/D 5.76e-21
C2246 _214_/a_27_257# _217_/A 0.0311f
C2247 _262_/a_199_7# _311_/Q 1.47e-19
C2248 _271_/A _184_/a_76_159# 0.00486f
C2249 result[0] _228_/A 0.00209f
C2250 _235_/a_113_257# _232_/X 5.55e-19
C2251 _149_/a_27_7# _147_/A 1.12e-19
C2252 _324_/a_1283_n19# _172_/A 2.12e-21
C2253 _324_/Q _316_/D 0.477f
C2254 _325_/Q _223_/a_250_257# 4.21e-20
C2255 _279_/Y _216_/A 0.00856f
C2256 _335_/a_193_7# _335_/a_543_7# -0.0231f
C2257 _340_/CLK _261_/A 0.0666f
C2258 output9/a_27_7# ctln[3] 0.0156f
C2259 _345_/a_476_7# _344_/a_476_7# 1.67e-19
C2260 _345_/a_1032_373# _344_/a_193_7# 1.95e-20
C2261 _146_/C _143_/a_181_7# 0.00167f
C2262 _255_/a_112_257# _298_/C 2.77e-19
C2263 _288_/A _310_/a_1108_7# 6.14e-19
C2264 _328_/a_761_249# _319_/Q 0.0436f
C2265 _149_/a_27_7# _149_/A 0.0316f
C2266 _335_/a_1270_373# VGND 5.26e-20
C2267 _335_/a_805_7# VPWR 3.06e-19
C2268 _341_/a_27_7# _269_/A 0.0164f
C2269 _180_/a_111_257# _286_/Y 6.08e-19
C2270 _184_/a_218_7# VGND 6.69e-20
C2271 _320_/D clkbuf_2_1_0_clk/A 1.22e-19
C2272 _291_/a_39_257# _289_/a_39_257# 5.11e-19
C2273 _302_/a_227_7# _304_/S 1.36e-19
C2274 _343_/a_193_7# _342_/a_27_7# 5.12e-20
C2275 _343_/a_27_7# _342_/a_193_7# 2.61e-20
C2276 output35/a_27_7# _267_/A 0.0738f
C2277 _281_/Y _190_/a_27_7# 0.0058f
C2278 _329_/a_27_7# _320_/Q 1.26e-20
C2279 _169_/B _147_/Y 1.64e-19
C2280 _287_/a_39_257# _310_/a_1108_7# 6.87e-19
C2281 _339_/a_761_249# _339_/D 6.85e-20
C2282 _153_/B VPWR 0.644f
C2283 _328_/a_193_7# _329_/D 2.45e-19
C2284 _320_/a_543_7# _279_/A 1.3e-20
C2285 _329_/a_27_7# _327_/a_193_7# 7.57e-22
C2286 _329_/a_193_7# _327_/a_27_7# 2.93e-19
C2287 _327_/a_27_7# _328_/Q 1.03e-19
C2288 _326_/a_1108_7# _216_/A 5.72e-19
C2289 _181_/X _283_/A 0.0236f
C2290 _338_/a_448_7# _193_/Y 1.37e-19
C2291 _338_/a_639_7# _194_/X 0.00129f
C2292 _254_/A _337_/Q 1.4e-19
C2293 output16/a_27_7# output39/a_27_7# 3.1e-20
C2294 repeater43/X clkbuf_0_clk/X 0.00214f
C2295 cal _226_/a_79_n19# 0.00539f
C2296 _325_/a_1270_373# repeater43/X -6.51e-20
C2297 _182_/a_297_257# _175_/Y 0.00203f
C2298 _341_/Q _231_/a_79_n19# 0.00121f
C2299 _324_/Q _222_/a_250_257# 2.15e-20
C2300 _215_/A _254_/B 0.00807f
C2301 _346_/SET_B _344_/Q 0.0259f
C2302 _325_/a_1283_n19# _217_/X 3.67e-21
C2303 _277_/Y _254_/B 1.29e-19
C2304 _275_/Y _309_/a_651_373# 0.00178f
C2305 _341_/a_1283_n19# _247_/a_113_257# 1.39e-21
C2306 _284_/A _201_/a_27_7# 0.037f
C2307 _285_/A _311_/a_27_7# 5.47e-21
C2308 _344_/a_381_7# _347_/Q 1.35e-21
C2309 _304_/a_288_7# _283_/A 1.38e-19
C2310 cal _339_/a_27_7# 1.31e-21
C2311 output19/a_27_7# _297_/B 0.00224f
C2312 _293_/a_121_257# VPWR -5.37e-19
C2313 _157_/A _313_/a_543_7# 5.57e-19
C2314 _320_/a_1108_7# _220_/a_250_257# 9.62e-20
C2315 _329_/a_27_7# _328_/a_27_7# 1.35e-19
C2316 _269_/A _316_/a_193_7# 0.00798f
C2317 _340_/a_805_7# _340_/Q 6.94e-19
C2318 _340_/a_448_7# _340_/D 0.00445f
C2319 _340_/a_639_7# _306_/S 0.00173f
C2320 ctln[5] _306_/S 5e-19
C2321 _316_/D _281_/A 5.51e-21
C2322 _336_/a_639_7# _147_/Y 0.00441f
C2323 _181_/X _248_/B 0.0098f
C2324 _322_/a_543_7# _321_/Q 0.00318f
C2325 _342_/Q _194_/A 3.12e-20
C2326 _255_/X _305_/X 0.00627f
C2327 _283_/Y _269_/Y 8.33e-19
C2328 _146_/C _304_/S 0.043f
C2329 _270_/a_39_257# _316_/a_27_7# 3.62e-21
C2330 _337_/Q _309_/D 0.00999f
C2331 repeater43/X input1/X 0.00414f
C2332 clkbuf_2_3_0_clk/A _301_/X 3.95e-20
C2333 ctln[1] clk 0.0376f
C2334 _271_/A _323_/a_1283_n19# 0.00114f
C2335 _321_/a_1462_7# _322_/Q 4.42e-19
C2336 _346_/a_1032_373# _346_/Q 0.00992f
C2337 _346_/a_476_7# _166_/Y 1.76e-19
C2338 _281_/Y _332_/Q 0.00772f
C2339 _339_/Q _337_/a_639_7# 8.3e-19
C2340 _322_/a_639_7# _318_/D 3.69e-20
C2341 _311_/a_761_249# _311_/D 4.6e-21
C2342 _157_/A _156_/a_121_257# 5.51e-19
C2343 _181_/a_27_7# VPWR 0.138f
C2344 _343_/a_193_7# _317_/D 5.41e-22
C2345 _218_/a_93_n19# _232_/X 0.0036f
C2346 trim[0] VGND 0.137f
C2347 _322_/a_193_7# VPWR -0.237f
C2348 _157_/A _304_/S 0.00209f
C2349 _188_/a_218_7# _286_/Y 0.00134f
C2350 _164_/A _265_/B 0.136f
C2351 _258_/S _257_/a_544_257# 3.52e-20
C2352 _170_/a_226_7# _147_/Y 0.043f
C2353 _273_/A _344_/D 2.02e-21
C2354 _337_/a_27_7# _284_/A 2.84e-20
C2355 _320_/a_448_7# VGND 0.00402f
C2356 _320_/a_1270_373# VPWR 4.09e-20
C2357 input4/a_27_7# _338_/a_193_7# 7.99e-20
C2358 _323_/a_805_7# VPWR 4.63e-19
C2359 _283_/A _332_/a_1283_n19# 1.91e-20
C2360 output33/a_27_7# _346_/SET_B 2.37e-19
C2361 clk _192_/B 0.0085f
C2362 clkbuf_0_clk/X _191_/B 7.14e-21
C2363 _322_/a_1283_n19# _318_/a_27_7# 3.34e-22
C2364 _214_/a_109_257# VGND -7.53e-19
C2365 _214_/a_373_7# VPWR -5.47e-19
C2366 _307_/X _146_/C 0.114f
C2367 trim[3] output5/a_27_7# 0.00358f
C2368 _305_/a_505_n19# VPWR 0.0626f
C2369 _344_/a_476_7# VGND 0.0196f
C2370 _344_/a_1032_373# VPWR -0.00368f
C2371 _232_/X _220_/a_256_7# 1.96e-19
C2372 _301_/X _172_/Y 2.09e-21
C2373 _318_/Q _318_/D 0.0394f
C2374 _273_/A _346_/Q 7.51e-20
C2375 result[3] _242_/B 0.00264f
C2376 _320_/a_805_7# _297_/B 2.33e-19
C2377 _346_/SET_B _221_/a_256_7# 1.56e-19
C2378 _340_/Q _340_/CLK 0.0106f
C2379 _343_/a_543_7# _323_/D 0.00689f
C2380 _326_/Q _223_/a_250_257# 0.0286f
C2381 _186_/a_79_n19# _184_/a_76_159# 7.15e-19
C2382 _344_/a_381_7# _297_/B 5.05e-19
C2383 _162_/A _297_/Y 0.00802f
C2384 _227_/A _333_/a_193_7# 7.72e-20
C2385 _260_/B _255_/B 4.74e-20
C2386 _258_/a_439_7# VGND 1.18e-19
C2387 _311_/Q VGND 0.347f
C2388 _285_/A _309_/a_1283_n19# 2.08e-19
C2389 _250_/X _295_/a_512_7# 5.78e-19
C2390 _257_/a_79_159# _260_/B 0.0751f
C2391 _325_/a_27_7# _325_/a_448_7# -0.00642f
C2392 _258_/S _310_/a_761_249# 3.71e-21
C2393 _331_/D _304_/X 2.13e-20
C2394 _246_/a_109_257# VPWR -0.00147f
C2395 _337_/a_1283_n19# _195_/a_27_257# 2.97e-21
C2396 _308_/X VGND 0.0965f
C2397 _271_/A _188_/S 0.00789f
C2398 ctlp[5] _220_/a_250_257# 1.12e-20
C2399 _342_/a_27_7# VGND -0.0655f
C2400 _342_/a_761_249# VPWR 0.00332f
C2401 repeater43/X _286_/Y 0.165f
C2402 _216_/A _316_/D 0.00602f
C2403 _318_/Q _217_/A 0.721f
C2404 _315_/Q _247_/a_199_7# 1.17e-19
C2405 _297_/A _314_/a_27_7# 0.00135f
C2406 _281_/Y _216_/a_27_7# 1.92e-21
C2407 _258_/S _264_/a_113_257# 0.013f
C2408 _211_/a_373_7# VGND -0.00132f
C2409 _254_/A _303_/A 1.28e-19
C2410 _198_/a_346_7# VGND -7.51e-19
C2411 _182_/a_297_257# _341_/Q 2.88e-19
C2412 _260_/A _156_/a_121_257# 1.03e-19
C2413 _267_/A _313_/a_1283_n19# 1.37e-19
C2414 input1/X _191_/B 0.00975f
C2415 cal _323_/Q 0.0498f
C2416 _219_/a_93_n19# _217_/X 0.0315f
C2417 _219_/a_250_257# _212_/X 0.00431f
C2418 _339_/Q _309_/D 2.09e-19
C2419 _240_/B _319_/a_193_7# 3.64e-22
C2420 _319_/Q _319_/a_1283_n19# 0.0708f
C2421 ctlp[1] _321_/a_193_7# 6.45e-20
C2422 _324_/Q _144_/A 0.00463f
C2423 _297_/A _170_/a_76_159# 1.8e-20
C2424 _207_/a_27_7# _206_/A 1.26e-21
C2425 _338_/D _193_/Y 0.0584f
C2426 _346_/SET_B _306_/S 0.0541f
C2427 _333_/a_1108_7# _154_/A 1.9e-19
C2428 _341_/Q _162_/X 1.18e-19
C2429 _209_/X _333_/D 0.0147f
C2430 _323_/a_193_7# _323_/a_543_7# -0.00424f
C2431 _332_/a_193_7# _153_/a_215_257# 8.01e-19
C2432 _336_/a_27_7# _194_/A 4.04e-20
C2433 _322_/Q _242_/B 0.00212f
C2434 ctln[7] _271_/Y 3.23e-20
C2435 _320_/a_1283_n19# _328_/D 1.31e-19
C2436 _304_/a_79_n19# _326_/Q 4.55e-19
C2437 _216_/A _313_/a_27_7# 0.609f
C2438 _329_/a_1108_7# _328_/a_448_7# 5.75e-21
C2439 _269_/A _316_/a_1462_7# 2.57e-19
C2440 _251_/X _347_/D 8.46e-21
C2441 _344_/Q _147_/A 0.0196f
C2442 _196_/A _298_/A 0.0157f
C2443 _216_/X _242_/A 0.00457f
C2444 _283_/Y _335_/a_1283_n19# 2.64e-19
C2445 ctln[7] _335_/a_761_249# 0.0186f
C2446 _182_/a_215_7# _227_/A 0.00635f
C2447 _258_/S _336_/a_27_7# 6.11e-19
C2448 result[2] _316_/a_1108_7# 0.00343f
C2449 _309_/a_1108_7# _171_/a_215_7# 7.88e-21
C2450 _283_/A _208_/a_215_7# 2.28e-20
C2451 _203_/a_209_7# VGND 6.94e-19
C2452 _286_/B _336_/a_651_373# 0.00167f
C2453 _345_/a_956_373# _172_/B 0.0013f
C2454 _339_/a_543_7# _195_/a_109_257# 7.6e-21
C2455 _339_/a_1283_n19# _195_/a_27_257# 6.31e-20
C2456 _319_/a_193_7# _328_/Q 2.95e-19
C2457 _254_/B VGND 4.3f
C2458 _191_/B _286_/Y 4.32e-20
C2459 _317_/D VGND 0.161f
C2460 _340_/D _190_/A 0.00183f
C2461 _329_/Q _242_/A 1.45e-19
C2462 _164_/A _310_/Q 2.02e-20
C2463 _346_/a_1224_7# _166_/Y 7.52e-20
C2464 _327_/a_761_249# _242_/A 7.09e-20
C2465 _145_/A _324_/Q 0.00177f
C2466 _311_/a_639_7# _311_/Q 1.55e-19
C2467 _298_/C _175_/Y 0.147f
C2468 _231_/a_409_7# _315_/D 0.00151f
C2469 _307_/a_76_159# _250_/X 8.93e-19
C2470 _307_/a_218_334# _216_/A 2.28e-20
C2471 _340_/a_27_7# _336_/a_543_7# 2.63e-21
C2472 _340_/a_543_7# _336_/a_27_7# 5.1e-22
C2473 _340_/a_761_249# _336_/a_193_7# 5.7e-21
C2474 _346_/a_1182_221# _167_/a_27_257# 1.68e-20
C2475 _332_/a_193_7# _209_/a_109_257# 5.83e-21
C2476 _322_/a_1462_7# VPWR 3.96e-19
C2477 _267_/B _261_/A 0.156f
C2478 _315_/a_543_7# _177_/A 1.45e-20
C2479 _313_/a_651_373# _284_/A 0.00177f
C2480 _315_/a_651_373# _177_/a_27_7# 7.93e-21
C2481 _330_/Q _330_/a_1283_n19# 0.00477f
C2482 _294_/A _346_/SET_B 0.412f
C2483 _326_/a_761_249# _242_/A 0.0437f
C2484 _344_/a_381_7# _275_/Y 0.00301f
C2485 _337_/Q _202_/a_250_257# 0.00774f
C2486 _346_/a_1140_373# _167_/X 9.57e-19
C2487 input4/X _194_/X 0.00269f
C2488 _298_/A _298_/X 3.82e-19
C2489 _183_/a_27_7# _146_/C 1.07e-20
C2490 _302_/a_227_7# _301_/X 0.0145f
C2491 _319_/Q _282_/a_121_257# 1.39e-19
C2492 _250_/a_215_7# _191_/B 0.00251f
C2493 _281_/A _331_/a_27_7# 4.37e-20
C2494 ctln[6] repeater43/X 0.00292f
C2495 _331_/D VGND 0.292f
C2496 _344_/a_1224_7# VGND 8.23e-20
C2497 _232_/X _328_/D 0.00232f
C2498 _255_/B _295_/a_512_7# 7.93e-19
C2499 _342_/Q _295_/a_306_7# 6.35e-19
C2500 _330_/a_193_7# VGND 0.0293f
C2501 _330_/a_543_7# VPWR 0.0143f
C2502 _144_/A _228_/A 0.023f
C2503 _286_/B _153_/A 4.19e-19
C2504 _346_/SET_B _327_/D 0.0104f
C2505 _329_/a_1108_7# _346_/SET_B -0.0051f
C2506 input1/X _337_/Q 0.0252f
C2507 clkbuf_2_3_0_clk/A _166_/Y 0.422f
C2508 _183_/a_27_7# _157_/A 0.00992f
C2509 _328_/a_193_7# _242_/A 2.53e-20
C2510 _281_/Y _327_/Q 0.0248f
C2511 _345_/a_27_7# _288_/A 1.84e-20
C2512 _164_/Y _215_/A 0.00167f
C2513 clk _157_/A 2.86e-19
C2514 _189_/a_27_7# _333_/Q 1.11e-19
C2515 _308_/X _184_/a_535_334# 0.00117f
C2516 _186_/a_79_n19# _188_/S 4.74e-19
C2517 _325_/a_543_7# _324_/Q 6.07e-19
C2518 _157_/a_27_7# _284_/A 0.0318f
C2519 _315_/Q _325_/Q 6.34e-21
C2520 _306_/S _206_/A 0.00876f
C2521 clkbuf_2_1_0_clk/A _312_/D 2.46e-20
C2522 _163_/a_78_159# _297_/Y 5.73e-20
C2523 _345_/a_27_7# _162_/X 9.68e-21
C2524 _306_/S _313_/a_761_249# 7.1e-20
C2525 _194_/X _313_/a_1283_n19# 3.49e-21
C2526 _255_/B _333_/Q 2.11e-21
C2527 _337_/a_1108_7# _193_/Y 0.00568f
C2528 _318_/Q _318_/a_448_7# 0.0164f
C2529 _342_/a_1217_7# VGND -4.44e-19
C2530 _194_/A _225_/B 0.00534f
C2531 _335_/a_639_7# _335_/D 0.00132f
C2532 _319_/Q _212_/X 0.514f
C2533 _166_/Y _172_/Y 1.62e-19
C2534 _312_/Q _310_/D 0.00187f
C2535 _252_/a_109_257# _297_/B 5.21e-19
C2536 _211_/a_27_257# _153_/B 0.0395f
C2537 _343_/CLK _193_/Y 3.08e-19
C2538 _286_/B _300_/a_383_7# 4.74e-19
C2539 _196_/A _300_/a_301_257# 3.89e-21
C2540 _273_/Y output5/a_27_7# 0.0126f
C2541 _334_/a_27_7# _204_/Y 2.48e-21
C2542 _217_/a_27_7# _281_/A 1.47e-19
C2543 _181_/X _298_/B 0.00826f
C2544 ctln[6] _334_/Q 3.64e-36
C2545 _292_/A _265_/B 0.0111f
C2546 _314_/a_193_7# _347_/a_193_7# 5.49e-19
C2547 _314_/a_761_249# _347_/a_27_7# 2.73e-19
C2548 _329_/D _327_/Q 2.67e-20
C2549 _258_/S _169_/Y 1.18e-20
C2550 _258_/S _225_/B 2.54e-20
C2551 _346_/SET_B _283_/A 0.419f
C2552 _216_/A _144_/A 2.43e-19
C2553 _265_/B _160_/A 0.0442f
C2554 _217_/A _223_/a_346_7# 9.29e-19
C2555 _304_/X _223_/a_584_7# 4.76e-19
C2556 _312_/a_543_7# _311_/a_543_7# 1.87e-20
C2557 _312_/a_27_7# _311_/a_448_7# 3.09e-20
C2558 _216_/A _331_/a_27_7# 1.33e-20
C2559 _339_/Q _202_/a_250_257# 4.87e-19
C2560 _274_/a_39_257# _242_/A 0.0589f
C2561 _271_/A _233_/a_113_257# 0.0072f
C2562 _196_/A _215_/A 0.00957f
C2563 _145_/A _228_/A 0.0711f
C2564 _157_/A _301_/X 0.0275f
C2565 _340_/a_1283_n19# _336_/Q 2.49e-20
C2566 _341_/a_448_7# _315_/a_193_7# 2.69e-20
C2567 repeater43/X _328_/Q 1.47e-21
C2568 ctln[6] _191_/B 2.85e-20
C2569 _281_/Y _192_/B 0.153f
C2570 _329_/a_193_7# repeater43/X 7.66e-19
C2571 _341_/a_448_7# _298_/A 3.56e-19
C2572 rstn _340_/CLK 4.6e-19
C2573 _277_/Y _196_/A 0.00974f
C2574 clkbuf_0_clk/X _303_/A 1.73e-20
C2575 _332_/a_761_249# _153_/A 5.17e-19
C2576 _332_/a_27_7# _154_/A 3.4e-19
C2577 clk _260_/A 1.47e-20
C2578 _229_/a_489_373# _175_/Y 0.00836f
C2579 ctlp[4] VPWR 0.121f
C2580 _345_/a_1032_373# _164_/A 4.61e-19
C2581 _202_/a_93_n19# _202_/a_346_7# -5.12e-20
C2582 result[2] _248_/A 1.65e-19
C2583 _306_/S _147_/A 0.296f
C2584 input1/X _339_/Q 0.0253f
C2585 _344_/a_27_7# _344_/a_1032_373# -0.00889f
C2586 _344_/a_193_7# _344_/a_1182_221# -2.22e-21
C2587 _331_/Q VPWR 0.769f
C2588 _200_/a_93_n19# clkbuf_2_0_0_clk/a_75_172# 3.06e-21
C2589 _263_/a_109_257# VPWR 8.28e-19
C2590 _346_/a_476_7# _242_/A 5.68e-20
C2591 _346_/SET_B _248_/B 1.26e-19
C2592 _281_/Y _325_/a_27_7# 0.00163f
C2593 _298_/B _343_/Q 1.1e-19
C2594 _275_/Y _312_/a_193_7# 0.02f
C2595 _341_/Q _298_/C 0.101f
C2596 _289_/a_39_257# _311_/a_1108_7# 0.00525f
C2597 _149_/A _306_/S 6.58e-22
C2598 _340_/CLK _310_/a_448_7# 1.08e-19
C2599 _182_/a_79_n19# VPWR 0.0606f
C2600 _317_/Q _236_/B 1.91e-19
C2601 _267_/B _340_/Q 3.98e-21
C2602 result[2] _331_/CLK 3.79e-19
C2603 _324_/a_193_7# _181_/X 0.00278f
C2604 _339_/a_543_7# _340_/D 0.00293f
C2605 _339_/a_1108_7# _193_/Y 9.86e-21
C2606 _339_/a_651_373# _340_/Q 9.07e-20
C2607 _339_/a_448_7# _306_/S 0.00257f
C2608 _339_/a_1270_373# _194_/X 1.29e-19
C2609 _312_/a_805_7# VPWR 0.00221f
C2610 _160_/X _299_/a_78_159# 0.00414f
C2611 _319_/a_27_7# _319_/D 0.0548f
C2612 _217_/a_27_7# _216_/A 1.63e-19
C2613 _335_/Q _332_/Q 0.23f
C2614 _207_/X _204_/Y 0.00421f
C2615 _300_/a_301_257# _347_/a_1283_n19# 3.93e-20
C2616 _300_/a_27_257# _347_/a_1108_7# 2.85e-20
C2617 _258_/a_76_159# _313_/D 0.00561f
C2618 _145_/A _216_/A 1.8e-19
C2619 _316_/a_193_7# _315_/a_651_373# 3.54e-21
C2620 _316_/a_1283_n19# _315_/a_1283_n19# 1.76e-21
C2621 _316_/a_651_373# _315_/a_193_7# 1.39e-20
C2622 _316_/a_1108_7# _315_/a_543_7# 2.33e-20
C2623 _324_/a_1283_n19# _304_/a_257_159# 8.83e-19
C2624 _254_/Y _346_/SET_B 0.0164f
C2625 repeater43/X _269_/A 0.0712f
C2626 _326_/a_543_7# _326_/Q 0.00139f
C2627 _232_/X _214_/a_109_7# 3.4e-19
C2628 _325_/a_639_7# _286_/Y 1.35e-19
C2629 _326_/D _317_/Q 2.08e-20
C2630 _234_/B _248_/A 2.67e-20
C2631 _251_/X _304_/S 1.34e-19
C2632 _301_/X _260_/A 1.44e-20
C2633 _342_/Q _226_/a_79_n19# 1.39e-20
C2634 _321_/a_1283_n19# _248_/A 3.29e-22
C2635 _162_/X _314_/D 2.98e-19
C2636 clkbuf_2_1_0_clk/A _338_/a_1283_n19# 3.56e-19
C2637 _342_/a_1108_7# _186_/a_297_7# 2.3e-20
C2638 _342_/a_193_7# _172_/A 6e-21
C2639 _258_/a_76_159# _197_/X 2.24e-19
C2640 _304_/a_591_329# _304_/X 1.71e-19
C2641 _304_/a_79_n19# _324_/D 1.81e-19
C2642 _330_/a_1462_7# VGND 0.00184f
C2643 _283_/A _206_/A 0.0347f
C2644 _321_/D _234_/a_109_257# 4.76e-19
C2645 _234_/B _331_/CLK 6.82e-20
C2646 _344_/a_1032_373# _171_/a_215_7# 9.59e-20
C2647 _294_/A _147_/A 4.19e-19
C2648 _343_/a_193_7# _298_/X 1.05e-19
C2649 _167_/a_109_257# clkbuf_2_3_0_clk/A 0.0051f
C2650 _321_/D _321_/a_27_7# 0.148f
C2651 _321_/a_1283_n19# _331_/CLK 0.0589f
C2652 repeater43/X _343_/D 4.51e-19
C2653 _346_/SET_B _310_/a_651_373# 0.00383f
C2654 _338_/Q _310_/a_1283_n19# 3.36e-19
C2655 _325_/a_543_7# _216_/A 0.00178f
C2656 _333_/a_805_7# VPWR 5.98e-20
C2657 _333_/a_1270_373# VGND 5.97e-20
C2658 cal _267_/A 7.36e-19
C2659 _275_/A _319_/D 0.103f
C2660 _242_/A _319_/a_543_7# 4.22e-19
C2661 _206_/A _205_/a_382_257# 5.26e-19
C2662 _299_/a_292_257# VPWR -8e-19
C2663 _315_/Q _315_/a_1283_n19# 0.0251f
C2664 clk _251_/a_79_n19# 0.00976f
C2665 _337_/D _306_/S 7.01e-21
C2666 _343_/a_27_7# _343_/Q 1.6e-19
C2667 _166_/Y _302_/a_227_7# 1.11e-19
C2668 output21/a_27_7# VGND 0.0819f
C2669 _292_/A _310_/Q 0.152f
C2670 output31/a_27_7# _338_/Q 2.98e-19
C2671 _153_/a_297_257# _333_/Q 0.00203f
C2672 _153_/a_215_257# _190_/A 0.00204f
C2673 _153_/a_403_257# _332_/Q 0.00224f
C2674 _196_/A _300_/Y 2.95e-19
C2675 _343_/CLK _205_/a_297_7# 1.33e-19
C2676 _223_/a_584_7# VGND -0.00126f
C2677 _303_/A _286_/Y 5.23e-20
C2678 _164_/Y VGND 0.102f
C2679 _209_/X _190_/A 0.00477f
C2680 clkbuf_2_3_0_clk/A _297_/Y 0.00933f
C2681 _238_/B clkbuf_2_1_0_clk/A 1.01e-19
C2682 _322_/a_193_7# _322_/a_651_373# -0.00701f
C2683 _306_/a_439_7# _147_/Y 1.01e-19
C2684 _269_/A _191_/B 2.42e-20
C2685 _261_/a_109_257# _261_/A 0.00129f
C2686 _312_/a_27_7# _311_/D 5.41e-19
C2687 _312_/D _311_/a_27_7# 4.17e-20
C2688 _346_/a_652_n19# _169_/Y 7.09e-22
C2689 _283_/A _147_/A 0.00738f
C2690 _323_/a_639_7# _323_/D 8.62e-19
C2691 _171_/a_78_159# _172_/B 0.00828f
C2692 _172_/Y _297_/Y 7.69e-20
C2693 _341_/D _315_/a_193_7# 8.41e-19
C2694 clkbuf_2_3_0_clk/A _310_/a_193_7# 2.28e-20
C2695 _233_/a_113_257# _232_/a_27_7# 4.99e-21
C2696 _341_/D _298_/A 0.0188f
C2697 _309_/a_1283_n19# _164_/A 0.014f
C2698 _342_/a_193_7# _244_/B 1.18e-19
C2699 _248_/B _156_/a_39_257# 7.62e-20
C2700 _183_/a_1241_257# _306_/S 2.66e-20
C2701 _202_/a_346_7# _284_/A 4.08e-19
C2702 _214_/a_27_257# _331_/D 0.0196f
C2703 clkbuf_2_0_0_clk/a_75_172# _340_/CLK 0.032f
C2704 _329_/a_1270_373# _217_/X 3.11e-20
C2705 _304_/S _232_/A 9.74e-20
C2706 _149_/A _283_/A 1.84e-21
C2707 _281_/Y _157_/A 0.00886f
C2708 _273_/A _265_/B 0.00752f
C2709 _185_/A _192_/B 1.12e-19
C2710 _343_/D _191_/B 3.19e-19
C2711 _209_/a_109_7# _333_/Q 8.44e-19
C2712 _209_/a_109_257# _190_/A 0.0471f
C2713 _209_/a_373_7# _332_/Q 1.72e-19
C2714 output14/a_27_7# VPWR 0.103f
C2715 _339_/a_448_7# _283_/A 0.0218f
C2716 _346_/SET_B _336_/a_1108_7# -0.0185f
C2717 _318_/Q _214_/a_109_257# 0.00201f
C2718 _210_/a_27_7# _207_/C 1.93e-19
C2719 _259_/a_199_7# VGND -3.88e-19
C2720 _340_/CLK _310_/D 0.00818f
C2721 _182_/X VPWR 0.132f
C2722 _196_/A VGND 3.63f
C2723 input1/X _336_/D 0.0294f
C2724 _324_/Q _228_/A 0.0313f
C2725 _279_/A _347_/a_193_7# 9.79e-21
C2726 _324_/a_1462_7# _181_/X 2.71e-19
C2727 _345_/a_27_7# _165_/a_215_7# 7.36e-20
C2728 _226_/a_297_7# _298_/a_27_7# 1.2e-20
C2729 _339_/D _306_/S 0.604f
C2730 _315_/a_543_7# _248_/A 0.00586f
C2731 _312_/Q VPWR 0.462f
C2732 _342_/a_193_7# _323_/D 6.44e-20
C2733 _248_/B _147_/A 1.08e-20
C2734 ctln[2] _297_/Y 1.44e-19
C2735 _230_/a_27_7# _317_/a_27_7# 3.69e-19
C2736 _227_/A _295_/a_79_n19# 0.00323f
C2737 _160_/X _347_/a_1108_7# 8.6e-20
C2738 _300_/Y _347_/a_1283_n19# 3.7e-19
C2739 _337_/a_193_7# _199_/a_93_n19# 9.26e-20
C2740 _194_/X _202_/a_93_n19# 0.00654f
C2741 _304_/a_591_329# VGND -2.58e-19
C2742 _304_/a_578_7# VPWR -3.07e-19
C2743 _255_/X _191_/B 0.0274f
C2744 _331_/CLK _315_/a_543_7# 5.47e-20
C2745 _324_/a_448_7# _216_/X 2.82e-20
C2746 _248_/A _314_/a_27_7# 2.76e-21
C2747 clkbuf_2_3_0_clk/A _242_/A 0.00154f
C2748 _283_/A _331_/a_761_249# 0.00175f
C2749 _343_/a_27_7# _229_/a_76_159# 1.02e-19
C2750 _256_/a_303_7# VGND -9.17e-20
C2751 repeater42/a_27_7# _181_/X 0.00214f
C2752 _169_/Y _173_/a_226_7# 7.78e-20
C2753 _279_/Y _324_/a_543_7# 2.22e-21
C2754 _248_/A _224_/a_250_257# 3.74e-20
C2755 _293_/a_121_257# _147_/Y 2.16e-19
C2756 trim[4] _265_/B 1.59e-19
C2757 _309_/a_543_7# _286_/B 5.95e-20
C2758 cal _194_/X 0.03f
C2759 _237_/a_199_7# VPWR -3.24e-19
C2760 VPWR valid 0.292f
C2761 VGND _298_/X 1.39f
C2762 _291_/a_39_257# _338_/Q 0.001f
C2763 _279_/Y _314_/a_805_7# 4.56e-19
C2764 _342_/a_1462_7# _172_/A 5.16e-21
C2765 clkbuf_0_clk/X clkbuf_1_0_0_clk/a_75_172# 0.0439f
C2766 _260_/B _314_/a_1462_7# 4.83e-20
C2767 _345_/a_1032_373# _292_/A 0.00823f
C2768 _317_/a_27_7# _232_/A 0.00954f
C2769 _254_/Y _147_/A 4.14e-19
C2770 _337_/a_193_7# _336_/Q 2.67e-20
C2771 _203_/a_80_n19# _203_/a_303_7# 8.88e-34
C2772 _242_/A _327_/Q 0.0849f
C2773 _267_/A _284_/A 0.0757f
C2774 _143_/a_27_7# _298_/A 4.58e-20
C2775 _165_/a_292_257# _160_/X 0.00307f
C2776 _279_/Y _217_/A 6.2e-21
C2777 _316_/D _224_/a_93_n19# 3.33e-19
C2778 _324_/Q _216_/A 0.0437f
C2779 _175_/Y _207_/C 4.53e-21
C2780 _337_/D _283_/A 5.08e-19
C2781 _281_/Y _260_/A 0.0118f
C2782 _345_/a_1032_373# _160_/A 0.0104f
C2783 _325_/Q _212_/X 2.22e-22
C2784 _333_/a_1108_7# _153_/B 5.27e-19
C2785 _320_/a_543_7# ctlp[4] 5.5e-19
C2786 _338_/Q _199_/a_346_7# 6.02e-19
C2787 _324_/Q _251_/a_510_7# 4.88e-19
C2788 _327_/a_448_7# _304_/X 0.00882f
C2789 _327_/a_1108_7# _217_/A 1.1e-20
C2790 _332_/a_543_7# VGND 0.00589f
C2791 _332_/a_1108_7# VPWR -0.00466f
C2792 _346_/a_1032_373# clkbuf_2_1_0_clk/A 0.0125f
C2793 _300_/a_27_257# _346_/SET_B 0.00413f
C2794 _315_/D _347_/a_805_7# 1.82e-19
C2795 _347_/a_1283_n19# VGND 0.0292f
C2796 _347_/a_448_7# VPWR -0.00229f
C2797 _346_/SET_B _284_/a_39_257# 8.03e-22
C2798 _200_/a_93_n19# VPWR 0.0197f
C2799 _326_/a_448_7# _304_/X 1.13e-20
C2800 _326_/a_1108_7# _217_/A 3.69e-19
C2801 trim[0] output32/a_27_7# 4.26e-20
C2802 clkbuf_2_1_0_clk/A _331_/CLK 0.0829f
C2803 _154_/A _333_/Q 0.221f
C2804 _165_/X _301_/X 2.53e-20
C2805 _305_/a_505_n19# _147_/Y 1.99e-19
C2806 repeater43/X _321_/a_1270_373# -1.24e-19
C2807 result[6] _269_/A 0.0664f
C2808 _308_/a_439_7# _181_/X 3.24e-19
C2809 _316_/Q _341_/a_27_7# 7.61e-22
C2810 _314_/Q _347_/a_543_7# 0.00935f
C2811 _297_/B _347_/a_1270_373# 5.54e-19
C2812 _336_/a_1108_7# _313_/a_761_249# 6.78e-22
C2813 _336_/a_1283_n19# _313_/a_543_7# 4.01e-20
C2814 _306_/a_535_334# _286_/B 1.39e-19
C2815 _188_/a_76_159# _298_/B 4.18e-20
C2816 _273_/A clkbuf_2_1_0_clk/A 0.00637f
C2817 _346_/a_193_7# _299_/X 0.0107f
C2818 _346_/a_27_7# _347_/Q 0.00689f
C2819 _343_/CLK _315_/a_193_7# 0.559f
C2820 _318_/Q _317_/D 2.21e-19
C2821 _343_/CLK _298_/A 1.02e-19
C2822 _225_/X _225_/a_59_35# 2.2e-19
C2823 _277_/Y _338_/D 3.39e-20
C2824 _292_/A _311_/a_27_7# 1.94e-20
C2825 _165_/a_78_159# VGND 0.0125f
C2826 _165_/a_493_257# VPWR 3.39e-20
C2827 _316_/a_193_7# _246_/B 2.27e-20
C2828 _183_/a_1241_257# _283_/A 0.00536f
C2829 _192_/B _335_/Q 0.00248f
C2830 _273_/A _310_/Q 0.023f
C2831 _323_/a_27_7# output41/a_27_7# 9.3e-19
C2832 _328_/a_543_7# _278_/a_68_257# 8.57e-20
C2833 _168_/a_109_257# _346_/Q 2.9e-19
C2834 _322_/Q _232_/X 0.0153f
C2835 _325_/a_1108_7# _283_/A 3.56e-36
C2836 _254_/A _336_/a_761_249# 4.1e-20
C2837 clkbuf_2_3_0_clk/A _199_/a_93_n19# 0.00106f
C2838 _175_/Y _150_/C 0.266f
C2839 _341_/a_1270_373# VPWR -1.59e-19
C2840 _341_/a_448_7# VGND -0.00361f
C2841 _342_/a_1462_7# _244_/B 1.03e-19
C2842 _339_/a_27_7# _225_/B 2.02e-20
C2843 _258_/a_505_n19# _162_/X 1.16e-20
C2844 _303_/A _328_/Q 2.67e-20
C2845 _338_/a_448_7# VGND 7.92e-19
C2846 _338_/a_1270_373# VPWR -2.18e-19
C2847 _184_/a_505_n19# _182_/X 0.00123f
C2848 _331_/D _330_/a_27_7# 2.38e-20
C2849 _325_/a_27_7# _242_/A 1.6e-20
C2850 _337_/Q clkc -1.05e-36
C2851 _178_/a_193_257# _298_/A 5.76e-19
C2852 _339_/D _283_/A 0.189f
C2853 _324_/a_193_7# _346_/SET_B 2.97e-21
C2854 _330_/a_27_7# _330_/a_193_7# -0.0552f
C2855 _329_/Q _220_/a_584_7# 0.00183f
C2856 _318_/Q _331_/D 0.0156f
C2857 _288_/A _285_/Y 8.75e-20
C2858 _316_/Q _316_/a_193_7# 0.0429f
C2859 _326_/a_27_7# _246_/B 1.73e-20
C2860 _290_/A _344_/Q 0.376f
C2861 clkbuf_2_1_0_clk/A _319_/a_1108_7# 9.85e-22
C2862 _318_/Q _330_/a_193_7# 1.04e-19
C2863 _325_/a_193_7# _325_/Q 3.46e-20
C2864 _328_/a_761_249# _279_/A 0.00687f
C2865 _216_/A _228_/A 0.0401f
C2866 clkbuf_2_3_0_clk/A _336_/Q 8.36e-21
C2867 trim[3] VGND 0.154f
C2868 _271_/A _316_/a_543_7# 1.68e-21
C2869 _229_/a_226_7# VPWR 0.00547f
C2870 _188_/S _162_/X 0.0514f
C2871 _251_/a_510_7# _228_/A 0.00423f
C2872 _325_/a_1108_7# _248_/B 2.46e-21
C2873 _149_/A _315_/a_27_7# 1.62e-19
C2874 _340_/a_805_7# VPWR 4.29e-19
C2875 _340_/a_1270_373# VGND 3.55e-20
C2876 _337_/Q _310_/a_543_7# 7.08e-19
C2877 _194_/X _284_/A 0.141f
C2878 _327_/a_639_7# _330_/Q 5.45e-19
C2879 _345_/a_652_n19# _346_/SET_B 0.0116f
C2880 _316_/a_639_7# VPWR 4.15e-19
C2881 _316_/a_651_373# VGND 0.00193f
C2882 _343_/a_543_7# _248_/A 0.00111f
C2883 _344_/a_1182_221# _164_/A 1.19e-19
C2884 _300_/a_27_257# _313_/a_761_249# 2.34e-20
C2885 _298_/B _206_/A 8.43e-20
C2886 _341_/Q _207_/C 4.58e-20
C2887 _346_/a_27_7# _297_/B 0.0109f
C2888 _162_/X _171_/a_493_257# 8.12e-19
C2889 _258_/S _309_/a_651_373# 2.26e-19
C2890 _204_/a_27_257# VGND -0.00748f
C2891 _204_/a_277_7# VPWR 0.00141f
C2892 _337_/Q _264_/a_199_7# 0.00111f
C2893 _208_/a_493_257# VGND -2.49e-19
C2894 _326_/Q _212_/X 0.0566f
C2895 _184_/a_76_159# _298_/C 2.84e-20
C2896 _309_/a_1283_n19# _292_/A 0.0116f
C2897 _279_/Y _314_/Q 0.0379f
C2898 _313_/a_651_373# _225_/B 2.27e-20
C2899 _296_/a_493_257# _286_/Y 3.67e-20
C2900 _327_/a_1270_373# VPWR 1.9e-19
C2901 _327_/a_448_7# VGND 4.68e-19
C2902 _157_/A _297_/Y 9.78e-20
C2903 _342_/a_1283_n19# _342_/D 0.0831f
C2904 _346_/a_1602_7# _346_/D 2.24e-20
C2905 _316_/D _217_/A 0.91f
C2906 _236_/B _304_/X 2.02e-20
C2907 _283_/A _150_/a_27_7# 0.00362f
C2908 repeater43/X _315_/a_651_373# 0.00351f
C2909 clk rstn 0.292f
C2910 _195_/a_109_257# _193_/Y 0.00201f
C2911 _195_/a_373_7# _340_/Q 2.21e-19
C2912 _326_/a_448_7# VGND -0.00248f
C2913 _326_/a_1270_373# VPWR -2.28e-19
C2914 _215_/A _313_/a_193_7# 0.548f
C2915 _167_/X _284_/A 2.26e-21
C2916 _274_/a_121_257# _279_/A 2.04e-19
C2917 output33/a_27_7# _290_/A 0.0319f
C2918 _339_/Q clkc 1.09e-20
C2919 _169_/Y _157_/a_27_7# 3.4e-20
C2920 _332_/a_27_7# _153_/B 0.0187f
C2921 _160_/X _346_/SET_B 0.652f
C2922 _340_/CLK VPWR 4.42f
C2923 _275_/A _347_/Q 8.1e-20
C2924 _328_/a_651_373# VPWR 0.00216f
C2925 _328_/a_1108_7# VGND -0.00286f
C2926 _347_/D VPWR 0.101f
C2927 clkbuf_0_clk/X _319_/D 0.00817f
C2928 _326_/D _304_/X 6.77e-20
C2929 clkbuf_2_3_0_clk/A _170_/a_489_373# 2.58e-19
C2930 _277_/Y _343_/CLK 0.0221f
C2931 _345_/a_1032_373# _273_/A 0.00197f
C2932 _271_/A _334_/a_193_7# 0.554f
C2933 _192_/B _336_/Q 0.159f
C2934 _217_/A _222_/a_250_257# 0.00497f
C2935 _300_/a_27_257# _147_/A 0.00678f
C2936 _267_/B _310_/D 0.0142f
C2937 _337_/Q _336_/a_193_7# 0.0113f
C2938 _341_/Q _150_/C 0.306f
C2939 _298_/B _147_/A 0.00759f
C2940 _319_/a_27_7# _297_/B 0.0217f
C2941 _346_/a_796_7# _299_/X 3.31e-19
C2942 _346_/a_586_7# _347_/Q 1.98e-20
C2943 _258_/a_439_7# _286_/B 1.8e-19
C2944 _216_/X _330_/D 0.014f
C2945 _334_/a_651_373# VPWR -0.0064f
C2946 _334_/a_1108_7# VGND -0.00764f
C2947 _257_/a_222_53# _260_/A 0.0049f
C2948 _218_/a_93_n19# _331_/CLK 0.00514f
C2949 _309_/a_27_7# _340_/CLK 0.0086f
C2950 _298_/B _149_/A 6.31e-20
C2951 _296_/a_109_7# _284_/A 1.6e-20
C2952 _308_/X _286_/B 0.0038f
C2953 _172_/A _181_/X 0.164f
C2954 cal _210_/a_27_7# 1.49e-19
C2955 result[4] _269_/A 0.0821f
C2956 _345_/a_27_7# _345_/Q 0.0031f
C2957 _165_/X _166_/Y 0.0787f
C2958 _341_/D VGND 1.47f
C2959 clkbuf_2_1_0_clk/A _217_/X 3.79e-20
C2960 _343_/a_193_7# _343_/CLK 0.00117f
C2961 _325_/a_193_7# _326_/Q 0.0171f
C2962 _250_/X _306_/S 1.8e-21
C2963 _273_/A _218_/a_93_n19# 1.96e-21
C2964 _324_/a_27_7# _304_/S 0.0652f
C2965 _181_/X _232_/X 0.0815f
C2966 _313_/Q _162_/X 1.91e-20
C2967 _338_/D VGND 0.323f
C2968 en _323_/Q 1.66e-19
C2969 _316_/Q _316_/a_1462_7# 0.00204f
C2970 output23/a_27_7# _331_/CLK 1.92e-20
C2971 _322_/Q _241_/a_113_257# 8.25e-19
C2972 _326_/D _272_/a_39_257# 9.7e-20
C2973 _329_/a_1283_n19# _281_/Y 0.00395f
C2974 _281_/Y _251_/X 0.196f
C2975 _183_/a_553_257# _298_/A 0.00608f
C2976 _273_/A _311_/a_27_7# 2.01e-21
C2977 _346_/a_27_7# _275_/Y 8.09e-21
C2978 _342_/Q sample 7.32e-20
C2979 _275_/A _297_/B 0.202f
C2980 _342_/a_193_7# _177_/A 1.57e-19
C2981 _227_/A _226_/X 1.04e-20
C2982 _188_/a_505_n19# VPWR 0.0743f
C2983 _271_/A _332_/Q 8.91e-20
C2984 _346_/a_381_7# VGND 0.00913f
C2985 repeater42/a_27_7# _346_/SET_B 0.00525f
C2986 _233_/a_199_7# _331_/Q 0.00133f
C2987 _172_/B trimb[4] 2.29e-20
C2988 _333_/a_193_7# _333_/a_543_7# -0.0233f
C2989 _335_/a_27_7# _332_/Q 2.88e-19
C2990 _237_/a_113_257# _232_/X 0.0128f
C2991 clkbuf_0_clk/a_110_7# _314_/a_27_7# 3.02e-19
C2992 _309_/a_193_7# _346_/SET_B 0.00767f
C2993 _335_/a_193_7# _207_/X 9.02e-19
C2994 _343_/a_27_7# _147_/A 1.73e-19
C2995 _321_/D VPWR 0.347f
C2996 _236_/B VGND 0.362f
C2997 _329_/a_1108_7# _319_/Q 0.0642f
C2998 _319_/Q _327_/D 3.06e-20
C2999 cal _175_/Y 0.0172f
C3000 _347_/Q _313_/a_1108_7# 4.69e-21
C3001 _299_/X _313_/a_448_7# 7.66e-20
C3002 _300_/Y _313_/a_193_7# 1.45e-19
C3003 _261_/A _310_/a_193_7# 2.14e-20
C3004 _339_/Q _336_/a_193_7# 1.02e-19
C3005 _328_/a_543_7# _328_/D 2.39e-19
C3006 _343_/a_27_7# _149_/A 1.88e-21
C3007 _200_/a_250_257# _311_/D 5.46e-20
C3008 _329_/a_1283_n19# _329_/D 0.0448f
C3009 _188_/S _298_/C 0.0116f
C3010 _283_/Y _338_/a_761_249# 7.03e-19
C3011 _323_/a_27_7# _334_/a_193_7# 1.21e-21
C3012 _321_/D _318_/a_543_7# 0.00267f
C3013 _236_/B _318_/a_1108_7# 1.78e-36
C3014 _318_/a_651_373# _331_/CLK 2.55e-20
C3015 _319_/D _286_/Y 6.44e-20
C3016 _273_/Y VGND 0.531f
C3017 _336_/a_543_7# _202_/a_93_n19# 6.11e-19
C3018 _172_/A _347_/a_1108_7# 2.63e-20
C3019 _286_/B _254_/B 0.428f
C3020 _143_/a_27_7# VGND 0.0265f
C3021 _143_/a_181_7# VPWR -1.55e-19
C3022 _219_/a_584_7# _319_/D 4.84e-20
C3023 _320_/Q output19/a_27_7# 8.2e-19
C3024 _294_/A _290_/A 0.00856f
C3025 _193_/Y _340_/D 0.00443f
C3026 _326_/D VGND 0.212f
C3027 input4/X _269_/Y 1.21e-20
C3028 ctlp[0] _322_/a_193_7# 2.48e-19
C3029 _254_/A _347_/Q 0.742f
C3030 repeater43/X _324_/a_1270_373# -2.06e-19
C3031 cal _336_/a_543_7# 9.44e-21
C3032 input1/X _336_/a_761_249# 0.0432f
C3033 _305_/a_535_334# _194_/A 0.00105f
C3034 _305_/a_218_7# _305_/X 6.02e-19
C3035 _222_/a_584_7# VPWR -6.78e-19
C3036 _222_/a_256_7# VGND 3.87e-19
C3037 _324_/a_1108_7# _212_/X 2.85e-19
C3038 _324_/a_1283_n19# _217_/X 5.16e-21
C3039 _319_/Q _283_/A 0.00808f
C3040 _289_/a_39_257# _263_/B 0.023f
C3041 repeater43/X _318_/a_27_7# 0.116f
C3042 _267_/B _266_/a_113_257# 0.00663f
C3043 _343_/a_651_373# repeater43/X 0.00109f
C3044 _329_/a_27_7# _329_/a_543_7# -0.00936f
C3045 _329_/a_193_7# _329_/a_761_249# -0.0157f
C3046 _313_/D _194_/A 3e-21
C3047 _309_/a_1283_n19# _273_/A 0.0037f
C3048 _167_/a_27_257# _306_/S 8.48e-19
C3049 _207_/C _269_/Y 0.00131f
C3050 _239_/a_113_257# _242_/A 0.0368f
C3051 _271_/A _334_/a_1462_7# 2.44e-19
C3052 _319_/a_639_7# VPWR 8.82e-35
C3053 _319_/a_651_373# VGND 0.0125f
C3054 _331_/a_27_7# _217_/A 0.0107f
C3055 _313_/a_543_7# VPWR -0.00664f
C3056 _313_/a_193_7# VGND 0.0217f
C3057 _344_/a_1182_221# _292_/A 0.00374f
C3058 _337_/a_1108_7# VGND -0.00735f
C3059 _337_/a_651_373# VPWR -0.00518f
C3060 _346_/SET_B _311_/a_1270_373# 1.37e-19
C3061 _297_/B _345_/D 0.0172f
C3062 _231_/a_512_7# _162_/X 1.44e-19
C3063 _183_/a_1241_257# _298_/B 1.63e-19
C3064 _183_/a_471_7# _341_/Q 1.5e-19
C3065 _160_/X _147_/A 2.6e-20
C3066 _324_/D _212_/X 8.38e-20
C3067 _342_/a_761_249# _341_/a_543_7# 1.35e-19
C3068 _342_/a_543_7# _341_/a_761_249# 1.53e-20
C3069 _258_/S _313_/D 0.0341f
C3070 _189_/a_27_7# _306_/S 0.0433f
C3071 _308_/S _295_/a_306_7# 8.73e-19
C3072 _344_/a_1602_7# _162_/A 2.91e-20
C3073 _197_/X _194_/A 0.0456f
C3074 _320_/Q _322_/a_543_7# 0.0316f
C3075 _343_/CLK VGND 1.43f
C3076 _346_/Q _301_/a_149_7# 4.31e-19
C3077 _212_/X _278_/a_150_257# 4.27e-20
C3078 _217_/X _278_/a_68_257# 0.00276f
C3079 _255_/B _306_/S 0.459f
C3080 _250_/X _283_/A 8.12e-22
C3081 _257_/a_79_159# _306_/S 0.00329f
C3082 _197_/X _338_/a_193_7# 1.39e-21
C3083 _260_/B _305_/a_505_n19# 1.86e-20
C3084 _307_/a_439_7# VPWR -3.8e-19
C3085 _307_/a_535_334# VGND -9.35e-20
C3086 _324_/a_1283_n19# _296_/Y 9.74e-21
C3087 _156_/a_121_257# VPWR -2.59e-19
C3088 _275_/Y _338_/Q 0.00742f
C3089 _317_/a_27_7# _245_/a_113_257# 3.55e-19
C3090 _165_/X _167_/a_109_257# 0.00357f
C3091 _304_/S VPWR 2.38f
C3092 rstn _195_/a_373_7# 0.00236f
C3093 input4/a_27_7# _194_/X 0.00252f
C3094 _258_/S _197_/X 4.75e-19
C3095 _275_/Y _275_/A 0.0939f
C3096 _325_/a_1462_7# _326_/Q 1.31e-19
C3097 _324_/a_1217_7# _304_/S 8.73e-19
C3098 _331_/CLK _328_/D 3.16e-20
C3099 _309_/a_1283_n19# trim[4] 6.45e-19
C3100 input1/X _199_/a_346_7# 0.00185f
C3101 _323_/D _343_/Q 0.00353f
C3102 _254_/A _297_/B 0.159f
C3103 _281_/Y rstn 1.44e-20
C3104 _271_/A _226_/a_382_257# 5.56e-19
C3105 _217_/a_27_7# _217_/A 0.0365f
C3106 _212_/X _279_/A 0.0136f
C3107 _178_/a_193_257# VGND -1.57e-19
C3108 _319_/Q _321_/a_193_7# 9.36e-20
C3109 repeater43/X _246_/B 0.00734f
C3110 _188_/S _229_/a_489_373# 1.4e-20
C3111 _164_/Y output40/a_27_7# 1.36e-19
C3112 _324_/Q _315_/a_761_249# 5.86e-19
C3113 _340_/a_543_7# _197_/X 0.00184f
C3114 _341_/Q cal 0.0668f
C3115 _340_/Q _310_/a_193_7# 6.28e-21
C3116 _218_/a_93_n19# _217_/X 0.0144f
C3117 _218_/a_250_257# _212_/X 0.00709f
C3118 _225_/X VPWR 2.56f
C3119 clkbuf_0_clk/X _227_/A 0.0122f
C3120 _162_/X _223_/a_93_n19# 3.11e-21
C3121 _307_/X VPWR 1.39f
C3122 _328_/a_193_7# _238_/a_109_257# 3.12e-20
C3123 _250_/X _248_/B 7.61e-21
C3124 _271_/A _282_/a_39_257# 0.00109f
C3125 _165_/X _297_/Y 0.00841f
C3126 _325_/a_448_7# _324_/a_27_7# 6.33e-19
C3127 _325_/a_193_7# _324_/a_1108_7# 5.86e-21
C3128 _325_/a_761_249# _324_/a_1283_n19# 0.00131f
C3129 _283_/Y _334_/a_193_7# 1.15e-19
C3130 _157_/A _314_/a_761_249# 7.58e-19
C3131 _320_/a_193_7# _319_/a_27_7# 1.52e-21
C3132 _255_/a_30_13# _255_/X 0.00604f
C3133 _335_/D _204_/a_27_7# 0.00116f
C3134 _316_/Q repeater43/X 0.426f
C3135 _267_/B VPWR 0.944f
C3136 _309_/a_1462_7# _346_/SET_B -9.14e-19
C3137 _335_/D _208_/a_215_7# 5.15e-19
C3138 _335_/a_1462_7# _207_/X 0.00211f
C3139 _260_/A _336_/Q 0.0869f
C3140 _339_/a_1108_7# VGND -0.00561f
C3141 _339_/a_651_373# VPWR 0.00166f
C3142 _212_/X _220_/a_346_7# 0.00223f
C3143 _217_/X _220_/a_256_7# 5.36e-19
C3144 _341_/a_1108_7# _317_/D 0.00725f
C3145 _324_/Q _224_/a_93_n19# 0.0526f
C3146 _308_/a_439_7# _206_/A 4.63e-20
C3147 _327_/a_651_373# _232_/X 0.00178f
C3148 _199_/a_93_n19# _261_/A 3.15e-21
C3149 _153_/B _333_/Q 0.0781f
C3150 _199_/a_250_257# _267_/A 3.67e-20
C3151 _341_/Q _150_/a_193_257# 1.72e-21
C3152 _258_/a_218_334# _340_/CLK 2.25e-19
C3153 _298_/B _150_/a_27_7# 0.0167f
C3154 _325_/a_1283_n19# _304_/X 0.0868f
C3155 _325_/a_193_7# _324_/D 2.55e-20
C3156 _325_/a_543_7# _217_/A 0.0109f
C3157 _240_/B _319_/D 0.00384f
C3158 _276_/a_68_257# _277_/Y 5.28e-21
C3159 _317_/a_27_7# VPWR 0.112f
C3160 repeater43/X _271_/Y 0.886f
C3161 _281_/Y _225_/a_59_35# 0.00225f
C3162 _343_/a_1283_n19# _149_/a_27_7# 1.91e-19
C3163 _343_/a_1217_7# _149_/A 2.71e-20
C3164 _169_/B _344_/Q 5.12e-20
C3165 _326_/a_651_373# _232_/X 0.00154f
C3166 output24/a_27_7# _269_/A 0.0131f
C3167 input4/X _335_/a_1283_n19# 4.56e-19
C3168 repeater43/X _335_/a_761_249# 7.91e-22
C3169 _309_/a_193_7# _147_/A 9.67e-21
C3170 _336_/a_193_7# _336_/D -0.0108f
C3171 _336_/a_543_7# _284_/A 9.44e-19
C3172 _330_/Q _331_/a_1283_n19# 0.018f
C3173 _321_/Q _331_/a_1108_7# 9.24e-21
C3174 _258_/S _312_/a_193_7# 9.79e-21
C3175 _271_/A _327_/Q 0.0128f
C3176 _318_/a_543_7# _317_/a_27_7# 0.00102f
C3177 _318_/a_27_7# _317_/a_543_7# 4.77e-21
C3178 _285_/A _346_/SET_B 0.00231f
C3179 _169_/Y _267_/A 0.0222f
C3180 _211_/a_27_257# _340_/CLK 0.0122f
C3181 _267_/A _225_/B 3.67e-20
C3182 _312_/a_1108_7# _312_/Q 0.0353f
C3183 _198_/a_93_n19# _340_/CLK 1.29e-21
C3184 input1/X _227_/A 0.265f
C3185 _309_/a_27_7# _267_/B 7.82e-19
C3186 _328_/a_448_7# _232_/X 7e-19
C3187 _331_/a_193_7# VGND 0.0372f
C3188 _331_/a_543_7# VPWR 0.0271f
C3189 output29/a_27_7# VGND 0.13f
C3190 _200_/a_584_7# _197_/X 3.45e-19
C3191 _320_/a_1283_n19# _346_/SET_B 1.71e-19
C3192 _325_/Q _306_/S 1.07e-20
C3193 _275_/Y _345_/D 0.185f
C3194 _275_/A _320_/a_193_7# 6.28e-21
C3195 _169_/B _168_/a_109_7# 0.00137f
C3196 _294_/A _310_/a_27_7# 3.05e-21
C3197 _335_/a_1283_n19# _207_/C 0.0022f
C3198 repeater43/X _318_/a_1217_7# 7.48e-19
C3199 _279_/Y _254_/B 0.0586f
C3200 _344_/a_193_7# _346_/SET_B 0.0173f
C3201 _316_/a_448_7# _317_/D 0.002f
C3202 _258_/S _289_/a_39_257# 0.0226f
C3203 _336_/a_27_7# _194_/X 1.55e-19
C3204 _302_/a_227_257# _297_/B 2.26e-20
C3205 _303_/A _314_/a_1283_n19# 7.98e-21
C3206 _260_/A _314_/a_761_249# 1.47e-19
C3207 _331_/a_1462_7# _304_/X 2.29e-19
C3208 _271_/Y _334_/Q 4.55e-19
C3209 _313_/a_1462_7# VGND -2.42e-20
C3210 _283_/Y _332_/Q 6.43e-19
C3211 _323_/D _229_/a_76_159# 9.84e-19
C3212 _319_/D _328_/Q 0.0102f
C3213 _181_/X _330_/a_805_7# 6.77e-21
C3214 ctln[1] _271_/A 0.0015f
C3215 _344_/a_1296_7# _292_/A 0.00106f
C3216 _258_/a_535_334# _346_/SET_B 3.83e-19
C3217 _335_/a_651_373# _343_/CLK 0.00123f
C3218 _335_/a_761_249# _334_/Q 2.36e-19
C3219 _322_/a_27_7# _331_/CLK 0.0329f
C3220 ctln[1] _335_/a_27_7# 0.00541f
C3221 _255_/B _283_/A 0.0084f
C3222 _172_/A _346_/SET_B 0.025f
C3223 _275_/Y _254_/A 2.62e-20
C3224 _214_/a_109_7# _331_/CLK 2.02e-19
C3225 _247_/a_199_7# _248_/B 6.43e-20
C3226 _315_/a_1270_373# _286_/Y 9.97e-21
C3227 _271_/Y _191_/B 1.37e-21
C3228 _271_/A _192_/B 0.0119f
C3229 _346_/SET_B _198_/a_250_257# 0.00649f
C3230 _232_/X _346_/SET_B 0.104f
C3231 _227_/A _286_/Y 0.398f
C3232 _188_/a_76_159# _172_/A 4.3e-21
C3233 result[0] _317_/D 0.00158f
C3234 _320_/Q _330_/a_1108_7# 0.0537f
C3235 _342_/a_193_7# _248_/A 0.0173f
C3236 _286_/B _164_/Y 1.56e-21
C3237 _146_/a_184_13# VGND -4.28e-19
C3238 result[6] _318_/a_27_7# 9.07e-20
C3239 repeater43/X _323_/a_761_249# 0.0105f
C3240 _314_/a_1108_7# _297_/a_27_257# 1.55e-19
C3241 _329_/a_1283_n19# _242_/A 5.34e-21
C3242 _184_/a_218_334# _147_/A 0.00122f
C3243 _184_/a_76_159# _150_/C 0.00305f
C3244 result[4] _242_/a_109_257# 3.41e-19
C3245 _255_/B _248_/B 0.0655f
C3246 _326_/D _214_/a_27_257# 6.26e-20
C3247 _307_/X _184_/a_505_n19# 2.8e-20
C3248 _301_/a_245_257# _297_/Y 0.00262f
C3249 _237_/a_113_257# _297_/A 3.34e-20
C3250 _183_/a_27_7# VPWR 0.00331f
C3251 _183_/a_553_257# VGND 0.0101f
C3252 _199_/a_250_257# _194_/X 0.0125f
C3253 _330_/D _327_/Q 6.44e-20
C3254 _324_/a_543_7# _324_/Q 5.26e-19
C3255 clk VPWR 2.94f
C3256 _333_/a_1283_n19# _298_/C 2.65e-19
C3257 _325_/a_1283_n19# VGND 0.0381f
C3258 _325_/a_448_7# VPWR -0.00504f
C3259 _275_/Y _309_/D 0.0342f
C3260 output13/a_27_7# _343_/CLK 0.0685f
C3261 _271_/A _317_/a_1108_7# 0.00177f
C3262 _181_/X _192_/a_68_257# 7.06e-22
C3263 _323_/a_1283_n19# _207_/C 1.12e-20
C3264 clkbuf_0_clk/X _297_/B 0.459f
C3265 _197_/X _201_/a_27_7# 6.92e-19
C3266 _217_/X _328_/D 0.0013f
C3267 _324_/Q _217_/A 0.058f
C3268 _257_/a_79_159# _254_/Y 0.00902f
C3269 _216_/A _224_/a_93_n19# 0.0187f
C3270 _169_/B _306_/S 3.67e-19
C3271 _306_/S _209_/a_109_7# 0.00388f
C3272 _194_/X _225_/B 7.01e-21
C3273 _340_/Q _336_/Q 0.0548f
C3274 _333_/a_1108_7# _332_/a_1108_7# 3.63e-20
C3275 _306_/X _340_/CLK 1.71e-19
C3276 _317_/a_1217_7# VPWR 8.58e-19
C3277 _317_/a_639_7# VGND -0.00139f
C3278 _323_/a_651_373# _343_/CLK 0.00344f
C3279 _286_/B _196_/A 0.11f
C3280 _297_/A _347_/a_1108_7# 0.00751f
C3281 output22/a_27_7# _342_/D 3.88e-19
C3282 _317_/Q result[2] 0.0043f
C3283 _337_/Q _311_/a_1283_n19# 1.01e-20
C3284 _325_/Q _283_/A 0.00621f
C3285 output21/a_27_7# ctlp[7] 0.0104f
C3286 _230_/a_27_7# _242_/A 0.0349f
C3287 _341_/a_27_7# _177_/a_27_7# 6.68e-20
C3288 _232_/a_27_7# _327_/Q 9.56e-20
C3289 _172_/A _313_/a_761_249# 0.00111f
C3290 _314_/a_448_7# _284_/A 4.62e-21
C3291 _347_/Q _286_/Y 0.0662f
C3292 _205_/a_79_n19# _335_/Q 0.0254f
C3293 _276_/a_68_257# VGND 0.0085f
C3294 _330_/Q _280_/a_150_257# 6.02e-19
C3295 _331_/a_1462_7# VGND 2.52e-19
C3296 _347_/Q _297_/a_27_257# 0.0103f
C3297 _304_/a_257_159# _181_/X 0.00102f
C3298 _277_/Y _344_/D 5.07e-20
C3299 _320_/D _346_/SET_B 0.0684f
C3300 _211_/a_109_257# _206_/A 7.24e-19
C3301 _323_/a_193_7# _323_/Q 0.00987f
C3302 _301_/X VPWR 0.406f
C3303 _169_/Y _167_/X 0.0183f
C3304 _335_/D _206_/A 0.0244f
C3305 _344_/a_796_7# _346_/SET_B 4.72e-19
C3306 _327_/a_543_7# _331_/Q 1.24e-19
C3307 _288_/A _162_/A 0.00625f
C3308 _197_/X _337_/a_27_7# 0.00783f
C3309 _316_/D _317_/D 7.88e-19
C3310 _343_/a_639_7# cal 5.58e-19
C3311 _190_/A _203_/a_303_7# 0.00203f
C3312 _277_/Y _346_/Q 0.0153f
C3313 _280_/a_68_257# VPWR 0.0311f
C3314 _283_/Y _339_/a_193_7# 3.51e-20
C3315 _219_/a_93_n19# _220_/a_93_n19# 0.00117f
C3316 _242_/A _232_/A 0.00228f
C3317 _162_/X _162_/A 0.00278f
C3318 _172_/A _307_/a_218_7# 9.5e-19
C3319 output31/a_27_7# clkc 0.00171f
C3320 _323_/a_543_7# _226_/X 3.73e-21
C3321 _281_/Y _324_/a_27_7# 0.0102f
C3322 _172_/A _156_/a_39_257# 3.39e-20
C3323 _150_/a_109_257# VPWR -5.31e-20
C3324 _174_/a_373_7# VPWR -7.11e-20
C3325 _216_/X _162_/X 2.59e-19
C3326 _174_/a_109_257# VGND -0.00171f
C3327 _335_/D _334_/D 0.153f
C3328 _321_/a_1108_7# _283_/A 7.82e-21
C3329 _294_/A _169_/B 2.67e-20
C3330 _322_/a_651_373# _321_/D 1.2e-19
C3331 _325_/Q _248_/B 6.84e-20
C3332 output7/a_27_7# _335_/D 0.00273f
C3333 _310_/a_193_7# _310_/a_448_7# -0.00297f
C3334 _323_/a_448_7# _149_/A 4.42e-20
C3335 _248_/A _330_/a_761_249# 1.2e-21
C3336 _324_/a_543_7# _228_/A 0.011f
C3337 _342_/Q _175_/Y 1.61e-20
C3338 _281_/A _217_/A 6.01e-19
C3339 _319_/Q _242_/B 3.09e-20
C3340 _181_/X _333_/D 2.42e-20
C3341 _283_/Y clkbuf_2_3_0_clk/A 1.56e-19
C3342 _261_/a_109_257# VPWR 0.00177f
C3343 result[3] _248_/A 1.65e-19
C3344 _321_/a_27_7# _242_/A 0.00561f
C3345 _219_/a_346_7# _330_/Q 6.49e-19
C3346 ctln[7] repeater43/X 0.00476f
C3347 _271_/A _146_/C 0.183f
C3348 _316_/D _330_/a_193_7# 3.59e-20
C3349 _331_/CLK _330_/a_761_249# 0.00196f
C3350 VGND output30/a_27_7# 0.11f
C3351 _340_/CLK _147_/Y 0.0843f
C3352 repeater43/X _179_/a_27_7# 7.07e-19
C3353 _324_/a_639_7# _286_/Y 5.72e-19
C3354 _172_/A _147_/A 0.273f
C3355 _318_/Q _236_/B 0.00602f
C3356 result[3] _331_/CLK 0.111f
C3357 _228_/A _217_/A 6.76e-22
C3358 _340_/CLK _312_/a_1108_7# 8.02e-20
C3359 _219_/a_256_7# VPWR -3.43e-19
C3360 _219_/a_93_n19# VGND -0.00267f
C3361 _309_/a_543_7# _174_/a_27_257# 5.8e-20
C3362 _306_/S _154_/A 0.00521f
C3363 repeater43/X _322_/a_1283_n19# 0.0567f
C3364 rstn _335_/Q 0.247f
C3365 _181_/X _325_/D 0.00946f
C3366 _255_/B _315_/a_27_7# 4.16e-21
C3367 _206_/A _203_/a_80_n19# 0.00974f
C3368 _339_/Q _311_/a_1283_n19# 2.79e-19
C3369 _176_/a_27_7# valid 2.25e-19
C3370 _298_/C output41/a_27_7# 2.3e-19
C3371 clkbuf_2_1_0_clk/A _193_/Y 0.106f
C3372 _297_/B _286_/Y 0.0148f
C3373 _326_/Q _327_/D 2.47e-19
C3374 _172_/A _149_/A 6.19e-19
C3375 _161_/Y _345_/D 0.00185f
C3376 _313_/a_27_7# _254_/B 1.97e-22
C3377 _297_/B _297_/a_27_257# 0.0124f
C3378 _219_/a_584_7# _297_/B 0.00183f
C3379 clk _335_/a_1108_7# 9.68e-21
C3380 _333_/a_27_7# _332_/Q 6.09e-19
C3381 _188_/S _150_/C 0.29f
C3382 _333_/a_193_7# _207_/X 1.11e-20
C3383 _345_/a_193_7# _166_/Y 0.00272f
C3384 _275_/Y clkbuf_0_clk/X 1.8e-21
C3385 _308_/a_218_334# input1/X 0.00203f
C3386 _214_/a_27_257# _331_/a_193_7# 0.00753f
C3387 _214_/a_109_257# _331_/a_27_7# 5.4e-20
C3388 _250_/a_292_257# VPWR -9.07e-19
C3389 _326_/D _318_/Q 6.44e-20
C3390 _234_/a_109_257# _322_/D 0.00391f
C3391 _324_/a_543_7# _216_/A 7.73e-19
C3392 _324_/a_193_7# _250_/X 1.41e-19
C3393 _334_/Q _154_/a_27_7# 4.71e-19
C3394 _214_/a_373_7# _212_/X 0.00157f
C3395 _197_/X _339_/a_27_7# 0.00313f
C3396 _321_/a_27_7# _322_/D 5e-20
C3397 _315_/D _221_/a_93_n19# 2.93e-19
C3398 _339_/a_651_373# _198_/a_93_n19# 1.84e-21
C3399 _321_/a_27_7# _321_/a_448_7# -0.00642f
C3400 ctln[7] _334_/Q 7.34e-20
C3401 _290_/A _262_/a_113_257# 2.49e-19
C3402 _268_/a_39_257# _316_/a_761_249# 0.00101f
C3403 _227_/A _328_/Q 3.63e-20
C3404 cal _311_/a_448_7# 3.63e-20
C3405 result[4] _318_/a_27_7# 0.00769f
C3406 ctln[1] _283_/Y 0.0257f
C3407 _323_/D _206_/A 0.0044f
C3408 output14/a_27_7# ctlp[0] 0.00541f
C3409 _216_/A _217_/A 0.0181f
C3410 _342_/a_1108_7# repeater43/X -8.76e-20
C3411 _236_/B _241_/a_199_7# 1.41e-19
C3412 _239_/a_199_7# _279_/A 1.82e-19
C3413 _283_/A _326_/Q 0.0345f
C3414 _346_/SET_B _312_/a_448_7# 2.49e-19
C3415 _338_/Q _312_/a_543_7# 3.21e-21
C3416 _191_/B _154_/a_27_7# 1.89e-20
C3417 _340_/a_193_7# _194_/A 5.52e-21
C3418 _322_/Q _248_/A 3.01e-19
C3419 _346_/Q _300_/Y 5.09e-20
C3420 ctln[7] _191_/B 3.39e-21
C3421 result[5] result[6] 0.0569f
C3422 _332_/a_193_7# _332_/a_1283_n19# -7.11e-33
C3423 _184_/a_76_159# cal 0.00267f
C3424 _313_/Q _313_/a_1283_n19# 0.00605f
C3425 _306_/X _313_/a_543_7# 4.51e-19
C3426 _275_/Y input1/X 1.39e-20
C3427 _340_/a_761_249# _338_/a_27_7# 3.37e-21
C3428 _232_/X _331_/a_761_249# 8.29e-19
C3429 _345_/a_652_n19# _290_/A 1.05e-19
C3430 _240_/B _347_/Q 1.05e-19
C3431 _179_/a_27_7# _191_/B 0.0324f
C3432 _341_/a_651_373# _177_/A 8.54e-19
C3433 ctln[4] _193_/Y 2.91e-20
C3434 _347_/a_193_7# _347_/a_448_7# -0.00482f
C3435 _169_/Y _301_/a_51_257# 0.00502f
C3436 _314_/D _284_/A 6.42e-20
C3437 _322_/Q _331_/CLK 0.00958f
C3438 _267_/A _311_/a_543_7# 0.0142f
C3439 _269_/A _315_/a_1270_373# 1.39e-19
C3440 _310_/D _297_/Y 0.00464f
C3441 _227_/A _269_/A 0.0224f
C3442 _323_/a_1462_7# _323_/Q 5.11e-19
C3443 _304_/S _227_/a_113_7# 7.41e-19
C3444 _279_/Y _196_/A 0.0188f
C3445 _149_/A _244_/B 0.0328f
C3446 _275_/A output17/a_27_7# 0.0249f
C3447 _197_/X _337_/a_1217_7# 4.35e-20
C3448 _195_/a_109_257# VGND -0.00267f
C3449 _195_/a_373_7# VPWR -5.39e-19
C3450 _182_/a_79_n19# _333_/Q 2.46e-19
C3451 _248_/B _326_/Q 0.00115f
C3452 _342_/Q _341_/Q 0.0323f
C3453 _255_/B _298_/B 3.52e-19
C3454 _161_/Y _309_/D 6.55e-20
C3455 _308_/X _145_/A 4.51e-21
C3456 _281_/Y VPWR 0.69f
C3457 _346_/a_476_7# _162_/X 2.98e-19
C3458 _325_/Q _315_/a_27_7# 1.25e-21
C3459 _341_/Q _144_/a_27_7# 7.46e-21
C3460 _254_/Y _169_/B 9.79e-21
C3461 _323_/a_1108_7# clk 9.08e-19
C3462 _344_/D VGND 0.347f
C3463 _163_/a_78_159# _162_/X 0.0288f
C3464 output22/a_27_7# _341_/a_193_7# 8.64e-19
C3465 _290_/A _160_/X 0.0155f
C3466 _310_/a_193_7# _310_/D 0.52f
C3467 _279_/Y _256_/a_303_7# 1.97e-20
C3468 _326_/a_1283_n19# _181_/X 6.12e-20
C3469 _297_/A _346_/SET_B 0.404f
C3470 _317_/Q _224_/a_250_257# 1.53e-20
C3471 _343_/D _227_/A 0.0311f
C3472 clkbuf_2_3_0_clk/A _312_/a_27_7# 4.86e-22
C3473 _323_/D _149_/A 2.12e-21
C3474 _306_/S _324_/D 2.04e-20
C3475 _209_/a_27_257# _153_/a_109_53# 9.12e-22
C3476 _346_/Q VGND 0.49f
C3477 _166_/Y VPWR 0.0706f
C3478 _186_/a_79_n19# _146_/C 1.22e-19
C3479 _275_/Y _286_/Y 1.1e-19
C3480 _342_/a_1283_n19# _323_/Q 7.18e-20
C3481 _210_/a_27_7# _225_/B 9.14e-21
C3482 _336_/a_193_7# _336_/a_761_249# -0.0157f
C3483 _336_/a_27_7# _336_/a_543_7# -0.00951f
C3484 _314_/Q _228_/A 1.06e-20
C3485 _283_/A _154_/A 0.0189f
C3486 _237_/a_113_257# _238_/B 0.00669f
C3487 _164_/A _346_/SET_B 0.0903f
C3488 _168_/a_481_7# VGND -8.12e-19
C3489 _248_/B _314_/a_193_7# 4.32e-20
C3490 _240_/B _297_/B 0.0157f
C3491 _329_/D VPWR 0.494f
C3492 _309_/a_1108_7# _344_/Q 3.78e-20
C3493 _309_/a_761_249# _344_/D 2.02e-19
C3494 _319_/Q _318_/a_1283_n19# 3.77e-20
C3495 _194_/a_27_7# _310_/a_27_7# 8.3e-22
C3496 _322_/a_543_7# result[7] 1.66e-21
C3497 _313_/a_543_7# _147_/Y 4.25e-21
C3498 _188_/S _183_/a_471_7# 0.00897f
C3499 _323_/a_1283_n19# cal 0.00893f
C3500 _333_/a_1217_7# _332_/Q 6.43e-20
C3501 repeater42/a_27_7# _319_/Q 6.5e-21
C3502 _345_/a_796_7# _166_/Y 3.32e-20
C3503 _200_/a_93_n19# _340_/a_1108_7# 2.9e-20
C3504 _256_/a_80_n19# _340_/CLK 2.83e-20
C3505 _329_/a_27_7# _330_/Q 0.00944f
C3506 _345_/a_193_7# _167_/a_109_257# 8.98e-20
C3507 _162_/X _173_/a_489_373# 4.66e-19
C3508 repeater43/X _330_/a_448_7# 4.17e-19
C3509 _331_/D _331_/a_27_7# 0.179f
C3510 _225_/a_59_35# _336_/Q 0.0041f
C3511 _331_/a_193_7# _330_/a_27_7# 5.06e-21
C3512 _164_/Y _163_/a_215_7# 0.00414f
C3513 _211_/a_109_257# _339_/D 6.75e-20
C3514 _197_/X _339_/a_1217_7# 3.56e-20
C3515 _292_/A _165_/a_292_257# 0.00251f
C3516 _316_/D _223_/a_584_7# 0.00169f
C3517 _344_/a_27_7# _301_/X 2.8e-20
C3518 _273_/A _299_/a_78_159# 0.0629f
C3519 _318_/Q _331_/a_193_7# 8.03e-20
C3520 _330_/a_543_7# _212_/X 1.99e-19
C3521 clkbuf_2_1_0_clk/A _301_/a_149_7# 0.0033f
C3522 repeater43/X _333_/a_761_249# -0.00336f
C3523 cal _311_/D 5.36e-20
C3524 _258_/a_76_159# input1/X 9.33e-20
C3525 _162_/a_27_7# _161_/Y 0.00141f
C3526 _315_/D _296_/a_109_7# 0.0282f
C3527 _145_/A _317_/D 9.8e-21
C3528 _338_/Q _263_/B 0.209f
C3529 _341_/Q _204_/Y 3.58e-19
C3530 _340_/a_27_7# _190_/a_27_7# 3.17e-20
C3531 _344_/a_476_7# _174_/a_27_257# 1.26e-20
C3532 _329_/a_193_7# _297_/B 5.38e-20
C3533 _297_/B _328_/Q 0.24f
C3534 _346_/SET_B _312_/D 0.00468f
C3535 _298_/B _298_/a_27_7# 0.00873f
C3536 _322_/a_1283_n19# result[6] 5.49e-19
C3537 _290_/A _309_/a_193_7# 0.00597f
C3538 _333_/a_448_7# _206_/A 0.0142f
C3539 _332_/a_27_7# _340_/CLK 0.0301f
C3540 _188_/S cal 0.0026f
C3541 _167_/a_27_257# _160_/X 0.00851f
C3542 _345_/a_1056_7# _290_/A 6.66e-19
C3543 _217_/a_27_7# _331_/D 3.97e-20
C3544 _294_/A _309_/Q 0.00499f
C3545 _321_/Q _269_/A 0.0545f
C3546 _172_/a_109_257# _172_/B 3.91e-19
C3547 _181_/X _248_/A 0.00845f
C3548 _153_/a_109_53# _153_/A 0.00207f
C3549 _347_/a_193_7# _347_/D 0.0577f
C3550 _334_/a_193_7# _298_/C 3.75e-21
C3551 _172_/A _150_/a_27_7# 0.0594f
C3552 _172_/A _174_/a_109_7# 0.00236f
C3553 _336_/a_1283_n19# _336_/Q 0.00858f
C3554 _331_/Q _282_/a_121_257# 6.94e-20
C3555 _324_/a_1108_7# _283_/A 1.17e-20
C3556 _181_/X _331_/CLK 0.0565f
C3557 result[2] _315_/a_1462_7# 2.2e-19
C3558 result[4] result[5] 0.0797f
C3559 _231_/a_512_7# _150_/C 0.0059f
C3560 _181_/X _190_/A 0.129f
C3561 _340_/D VGND 0.441f
C3562 _324_/a_27_7# _242_/A 1.37e-21
C3563 _325_/Q _242_/B 2.42e-20
C3564 clkbuf_2_0_0_clk/a_75_172# _199_/a_93_n19# 5.17e-19
C3565 _269_/A _318_/a_193_7# 0.0131f
C3566 _297_/A _156_/a_39_257# 1.94e-21
C3567 _317_/a_1270_373# _317_/D 3.74e-20
C3568 _188_/a_76_159# _177_/A 0.0035f
C3569 _273_/A _181_/X 0.00842f
C3570 _283_/A _324_/D 0.00936f
C3571 output24/a_27_7# _318_/a_27_7# 7.71e-21
C3572 _315_/a_193_7# _315_/a_543_7# -0.0129f
C3573 result[0] _341_/a_448_7# 5.06e-19
C3574 _333_/a_761_249# _191_/B 0.0143f
C3575 _333_/a_27_7# _192_/B 0.0124f
C3576 _310_/a_1462_7# _310_/D 8.56e-19
C3577 _185_/A VPWR 0.337f
C3578 _218_/a_250_257# _327_/D 1.29e-19
C3579 _331_/Q _212_/X 0.067f
C3580 _209_/a_27_257# _153_/A 0.0476f
C3581 _338_/a_543_7# _340_/CLK 0.0303f
C3582 _294_/A _311_/a_193_7# 7.75e-21
C3583 _248_/A _343_/Q 7.7e-21
C3584 _237_/a_113_257# _331_/CLK 0.0638f
C3585 _167_/a_109_257# VPWR 0.00183f
C3586 _247_/a_113_257# VGND -0.00229f
C3587 _327_/a_639_7# _216_/X 4.87e-19
C3588 _346_/SET_B _347_/a_761_249# -0.00726f
C3589 _219_/a_250_257# _232_/X 0.00215f
C3590 _181_/X _222_/a_93_n19# 0.00857f
C3591 _207_/a_27_7# _153_/B 5.09e-19
C3592 _343_/a_805_7# _185_/A 6.71e-19
C3593 clkbuf_2_3_0_clk/A _162_/X 0.303f
C3594 _297_/A _147_/A 0.0113f
C3595 _172_/A _250_/a_78_159# 2.39e-20
C3596 _224_/a_250_257# _298_/A 2.69e-20
C3597 _321_/a_1108_7# _242_/B 4.01e-20
C3598 _298_/C _332_/Q 4.1e-19
C3599 _286_/B _313_/a_193_7# 0.00527f
C3600 _196_/A _313_/a_27_7# 1.39e-20
C3601 _314_/a_1283_n19# _260_/a_27_257# 8.51e-20
C3602 _248_/B _324_/D 1.12e-19
C3603 repeater43/X _177_/a_27_7# 0.00514f
C3604 ctlp[1] _331_/CLK 1.48e-20
C3605 _340_/a_1108_7# _340_/CLK 1.1e-20
C3606 _324_/a_1462_7# _255_/B 1.79e-20
C3607 _164_/A _147_/A 9.05e-20
C3608 _257_/a_222_53# VPWR 0.00378f
C3609 _297_/Y VPWR 2.78f
C3610 _341_/a_1108_7# _341_/D 0.0393f
C3611 _329_/a_1217_7# _330_/Q 1.09e-19
C3612 _260_/B _340_/CLK 0.142f
C3613 _311_/D _284_/A 1.8e-20
C3614 _162_/X _172_/Y 1e-19
C3615 _313_/Q _202_/a_93_n19# 7.52e-21
C3616 _258_/a_505_n19# _284_/A 0.0263f
C3617 rstn output6/a_27_7# 0.0121f
C3618 _332_/a_448_7# _332_/Q 7.66e-19
C3619 _332_/a_1283_n19# _190_/A 3.37e-19
C3620 _332_/a_1108_7# _333_/Q 0.00998f
C3621 _340_/a_27_7# _337_/a_193_7# 0.00102f
C3622 _340_/a_193_7# _337_/a_27_7# 0.00102f
C3623 _338_/Q _194_/A 8.19e-19
C3624 output35/a_27_7# _162_/A 6.35e-19
C3625 _254_/A _263_/B 5.52e-21
C3626 _215_/A _265_/B 1.11e-19
C3627 output24/a_27_7# _246_/B 1.72e-19
C3628 _307_/a_505_n19# _181_/X 0.00228f
C3629 _329_/a_805_7# VPWR 2.99e-19
C3630 _338_/a_1283_n19# _346_/SET_B -0.00169f
C3631 _338_/a_193_7# _338_/Q -1.36e-19
C3632 _338_/a_1108_7# _338_/D 0.0492f
C3633 _313_/Q cal 9.33e-20
C3634 _277_/Y _265_/B 3.77e-20
C3635 _320_/Q _319_/a_27_7# 1.09e-19
C3636 _197_/X _202_/a_346_7# -6.1e-21
C3637 _310_/a_193_7# VPWR 0.0612f
C3638 _258_/S _338_/Q 0.327f
C3639 _325_/Q _245_/a_199_7# 0.00142f
C3640 _270_/a_39_257# _246_/B 3.39e-20
C3641 _306_/a_439_7# _306_/S 2.32e-19
C3642 _344_/a_1032_373# _344_/Q 0.0352f
C3643 _344_/a_652_n19# _344_/D 0.0018f
C3644 _341_/a_651_373# _248_/A 0.00539f
C3645 _342_/a_651_373# cal 4.56e-19
C3646 _248_/B _279_/A 2.35e-19
C3647 _292_/A _346_/SET_B 0.0302f
C3648 _181_/X _178_/a_27_7# 0.00126f
C3649 _294_/A _309_/a_1108_7# 0.0397f
C3650 _316_/Q output24/a_27_7# 4.07e-19
C3651 _304_/a_79_n19# _304_/S 0.0542f
C3652 _333_/D _206_/A 0.0612f
C3653 _290_/A _309_/a_1462_7# 1.83e-19
C3654 repeater43/X _268_/a_121_257# 8.92e-19
C3655 _346_/SET_B _160_/A 3.1e-19
C3656 _340_/a_448_7# _346_/SET_B -1.22e-19
C3657 ctlp[2] trimb[2] 0.00294f
C3658 _182_/X _226_/a_297_7# 0.0175f
C3659 _324_/Q _317_/D 0.00977f
C3660 _328_/a_27_7# _328_/a_639_7# -0.0015f
C3661 _316_/Q _270_/a_39_257# 0.0036f
C3662 _332_/a_193_7# _206_/A 0.001f
C3663 _271_/A _230_/a_27_7# 3.29e-19
C3664 _146_/C _231_/a_79_n19# 0.0429f
C3665 _309_/D _263_/B 0.242f
C3666 _271_/A _205_/a_79_n19# 0.00254f
C3667 _229_/a_76_159# _248_/A 0.0414f
C3668 _313_/D _267_/A 6.54e-20
C3669 _326_/Q _242_/B 7.7e-21
C3670 _238_/B _346_/SET_B 0.473f
C3671 _281_/Y _211_/a_27_257# 0.00115f
C3672 _275_/A _320_/Q 1.89e-19
C3673 _327_/a_1283_n19# _346_/SET_B 0.0814f
C3674 _324_/a_193_7# _326_/Q 0.00117f
C3675 _306_/S _153_/B 0.17f
C3676 result[2] VGND 0.208f
C3677 _285_/A _290_/A 0.00111f
C3678 _318_/Q _219_/a_93_n19# 3.65e-19
C3679 _346_/a_27_7# _346_/a_652_n19# -0.00237f
C3680 _242_/A VPWR 3.23f
C3681 repeater43/X _341_/a_27_7# 0.00392f
C3682 _316_/a_1270_373# _248_/A 1.25e-19
C3683 _335_/Q VPWR 1.29f
C3684 _177_/A _147_/A 0.00117f
C3685 _215_/A _314_/a_27_7# 4.11e-20
C3686 input4/X _338_/a_761_249# 1.36e-19
C3687 _343_/a_448_7# _175_/Y 3.78e-20
C3688 _197_/X _267_/A 2.94e-19
C3689 _271_/A _232_/A 0.604f
C3690 _340_/a_193_7# _339_/a_27_7# 0.00145f
C3691 _340_/a_27_7# _339_/a_193_7# 0.00138f
C3692 _342_/a_1283_n19# sample 3.96e-19
C3693 _216_/A _214_/a_109_257# 5.37e-21
C3694 _342_/a_448_7# _286_/Y 0.00846f
C3695 result[0] _341_/D 0.00252f
C3696 _298_/B _154_/A 8.05e-20
C3697 _320_/a_193_7# _328_/Q 3.85e-20
C3698 _242_/A _318_/a_543_7# 0.0172f
C3699 _319_/Q _232_/X 0.00672f
C3700 _344_/a_193_7# _290_/A 0.00325f
C3701 _294_/A _306_/a_439_7# 0.0021f
C3702 _298_/a_109_7# VPWR -6.73e-20
C3703 clkbuf_0_clk/X _330_/a_651_373# 2.43e-19
C3704 _149_/A _177_/A 1.15f
C3705 _328_/a_543_7# _346_/SET_B -9.86e-19
C3706 input1/X _312_/a_543_7# 1.12e-19
C3707 _334_/a_27_7# _334_/a_639_7# -0.0015f
C3708 _271_/A _321_/a_27_7# 1.1e-20
C3709 _181_/X _217_/X 0.0284f
C3710 _293_/a_39_257# _193_/Y 8.31e-19
C3711 clk _333_/a_1108_7# 4.61e-20
C3712 _327_/a_651_373# _331_/CLK 0.0268f
C3713 _204_/a_277_7# _333_/Q 0.00194f
C3714 _301_/X _147_/Y 0.171f
C3715 _208_/a_215_7# _190_/A 5.98e-20
C3716 _172_/A _250_/X 0.117f
C3717 _342_/Q _184_/a_76_159# 3.46e-20
C3718 _290_/A _172_/A 3.18e-19
C3719 _338_/a_448_7# _337_/a_1283_n19# 2.65e-21
C3720 _338_/a_651_373# _337_/a_543_7# 1.15e-20
C3721 _338_/a_543_7# _337_/a_651_373# 6.56e-21
C3722 _326_/a_1108_7# _236_/B 5.05e-20
C3723 clkbuf_2_1_0_clk/A _215_/A 0.0077f
C3724 _322_/D VPWR 1.08f
C3725 _234_/B VGND 0.403f
C3726 _326_/a_651_373# _331_/CLK 1.93e-20
C3727 repeater43/X _316_/a_193_7# 0.00661f
C3728 _305_/a_218_7# _336_/D 1.68e-19
C3729 _311_/a_1283_n19# _310_/a_1283_n19# 2.44e-19
C3730 _321_/a_448_7# VPWR 0.00332f
C3731 _321_/a_1283_n19# VGND 0.00602f
C3732 _314_/a_1283_n19# _314_/a_1108_7# 5.68e-32
C3733 _314_/a_27_7# _314_/a_639_7# -0.0015f
C3734 _283_/Y _340_/Q 3.31e-19
C3735 _277_/Y clkbuf_2_1_0_clk/A 0.00938f
C3736 rstn _335_/a_27_7# 0.513f
C3737 _338_/a_1108_7# _343_/CLK 3.33e-19
C3738 _254_/A _194_/A 6.03e-20
C3739 _169_/B _160_/X 3.94e-20
C3740 _162_/A _345_/Q 6.03e-20
C3741 _234_/B _318_/a_1108_7# 3.09e-19
C3742 _322_/D _318_/a_543_7# 4.55e-19
C3743 _181_/a_27_7# _306_/S 7.1e-20
C3744 _313_/Q _284_/A 0.268f
C3745 _224_/a_93_n19# _217_/A 0.00889f
C3746 _224_/a_250_257# _304_/X 0.00104f
C3747 _228_/A _317_/D 0.00958f
C3748 _153_/a_403_257# VPWR -0.00123f
C3749 _153_/a_215_257# VGND 0.00985f
C3750 _332_/D _332_/Q 0.154f
C3751 _340_/a_651_373# _337_/a_1108_7# 5.28e-20
C3752 _340_/a_1108_7# _337_/a_651_373# 5.28e-20
C3753 _267_/A _312_/a_193_7# 0.00108f
C3754 _261_/A _312_/a_27_7# 5.44e-20
C3755 _209_/X VGND 0.176f
C3756 _326_/a_1108_7# _326_/D 3.83e-21
C3757 _326_/a_27_7# repeater43/X 0.218f
C3758 _258_/S _254_/A 0.0139f
C3759 _279_/Y _313_/a_193_7# 2.49e-21
C3760 _296_/Y _181_/X 0.0106f
C3761 _260_/B _313_/a_543_7# 1.34e-19
C3762 _145_/A _196_/A 3.61e-20
C3763 _275_/Y _310_/a_543_7# 0.00547f
C3764 _305_/a_505_n19# _306_/S 0.0274f
C3765 _331_/D _281_/A 6.03e-20
C3766 _281_/A _330_/a_193_7# 0.00147f
C3767 _310_/a_1462_7# VPWR 2.28e-19
C3768 clkbuf_2_3_0_clk/a_75_172# _297_/B 0.00975f
C3769 _199_/a_93_n19# VPWR 0.0183f
C3770 repeater43/X _332_/a_1270_373# 7.85e-20
C3771 _279_/Y _343_/CLK 2.68e-19
C3772 _342_/D input1/X 5.21e-21
C3773 _343_/D _323_/a_543_7# 0.00212f
C3774 _187_/a_27_7# _341_/Q 0.0126f
C3775 _346_/SET_B _248_/A 4.45e-20
C3776 _341_/Q _315_/D 0.00976f
C3777 _341_/a_1283_n19# _149_/A 0.00267f
C3778 _334_/D _208_/a_78_159# 0.00277f
C3779 _343_/CLK _208_/a_292_257# 1.36e-20
C3780 _265_/B VGND 0.172f
C3781 _309_/D _194_/A 1.94e-19
C3782 ctlp[7] output29/a_27_7# 6.08e-19
C3783 _302_/a_77_159# _347_/a_27_7# 5.64e-19
C3784 _183_/a_553_257# _286_/B 0.00529f
C3785 _346_/a_1032_373# _346_/SET_B 0.099f
C3786 _255_/a_30_13# _179_/a_27_7# 5.22e-19
C3787 _271_/A _243_/a_199_7# 4.97e-19
C3788 _277_/Y ctln[4] 0.00457f
C3789 _209_/a_373_7# VPWR -6.14e-19
C3790 _209_/a_109_257# VGND -0.00329f
C3791 _325_/a_761_249# _181_/X 0.00596f
C3792 _216_/A _254_/B 0.0644f
C3793 _336_/Q VPWR 0.645f
C3794 _346_/SET_B _331_/CLK 0.0473f
C3795 _347_/Q _314_/a_1283_n19# 9.02e-20
C3796 _146_/C _162_/X 2.37e-19
C3797 input4/X _334_/a_193_7# 0.00729f
C3798 _283_/A _153_/B 0.204f
C3799 _197_/X _194_/X 0.252f
C3800 _337_/a_761_249# _340_/CLK 0.022f
C3801 _232_/a_27_7# _230_/a_27_7# 8.38e-21
C3802 _272_/a_39_257# _224_/a_250_257# 1.26e-20
C3803 _258_/S _309_/D 0.38f
C3804 _346_/SET_B _190_/A 1.21e-19
C3805 _294_/Y trim[0] 0.00272f
C3806 _335_/a_1283_n19# _204_/Y 8.36e-19
C3807 _335_/a_1108_7# _335_/Q 0.0279f
C3808 _157_/A _162_/X 0.709f
C3809 _160_/X _170_/a_226_7# 0.0307f
C3810 _338_/Q _201_/a_27_7# 1.75e-19
C3811 _319_/a_27_7# _319_/a_761_249# -6.54e-19
C3812 _324_/a_1462_7# _326_/Q 1.06e-19
C3813 _273_/A _346_/SET_B 0.0127f
C3814 result[0] _343_/CLK 0.187f
C3815 repeater43/X _341_/a_1217_7# -1.47e-19
C3816 _309_/a_761_249# _265_/B 0.00898f
C3817 _344_/a_27_7# _297_/Y 0.551f
C3818 _298_/C _192_/B 0.0847f
C3819 _334_/a_543_7# _206_/A 1.7e-20
C3820 _334_/a_193_7# _207_/C 0.0251f
C3821 _216_/A _331_/D 5.08e-21
C3822 _342_/D _286_/Y 0.0259f
C3823 _285_/A _310_/a_27_7# 6.57e-22
C3824 _232_/a_27_7# _232_/A 0.0141f
C3825 _315_/Q _304_/S 1.34e-19
C3826 input1/X _263_/B 1.36e-19
C3827 _236_/B _316_/D 0.0128f
C3828 ctln[5] _339_/a_543_7# 1.71e-19
C3829 _315_/a_543_7# VGND 0.0194f
C3830 _315_/a_1108_7# VPWR -0.0014f
C3831 _284_/a_39_257# _309_/Q 0.0115f
C3832 en _269_/Y 6.11e-19
C3833 repeater42/a_27_7# _326_/Q 0.00401f
C3834 _255_/B _172_/A 0.0395f
C3835 _294_/Y _311_/Q 3.21e-20
C3836 _336_/a_805_7# VPWR 1.03e-19
C3837 _336_/a_1270_373# VGND 1.8e-19
C3838 _324_/a_27_7# _324_/a_448_7# -0.00972f
C3839 _324_/a_193_7# _324_/a_1108_7# 1.42e-32
C3840 _334_/a_1283_n19# _343_/CLK 4.77e-19
C3841 _334_/a_543_7# _334_/D 0.0336f
C3842 repeater43/X _229_/a_556_7# 2.95e-19
C3843 _315_/D _314_/a_448_7# 0.0249f
C3844 _291_/a_39_257# _311_/a_1283_n19# 0.0013f
C3845 _314_/a_27_7# VGND -0.0714f
C3846 _314_/a_761_249# VPWR 0.017f
C3847 _344_/a_1182_221# comp 9.73e-20
C3848 _346_/SET_B _319_/a_1108_7# -0.00977f
C3849 _342_/Q _188_/S 0.269f
C3850 _338_/D _337_/a_1283_n19# 1.76e-21
C3851 _338_/Q _337_/a_27_7# 2.25e-21
C3852 _338_/a_27_7# _337_/Q 2.26e-20
C3853 _346_/SET_B _337_/a_543_7# 0.00688f
C3854 trim[4] _346_/SET_B 4.72e-19
C3855 _224_/a_250_257# VGND 0.00426f
C3856 _224_/a_346_7# VPWR -8.77e-19
C3857 clk _332_/a_27_7# 0.00328f
C3858 _326_/D _316_/D 7.04e-21
C3859 _299_/X _347_/Q 0.0663f
C3860 repeater43/X _316_/a_1462_7# -9.14e-19
C3861 _324_/a_193_7# _324_/D 0.513f
C3862 _324_/a_543_7# _217_/A 3.95e-20
C3863 _324_/a_1283_n19# _304_/X 8.43e-19
C3864 _311_/D _310_/a_761_249# 1.09e-19
C3865 _311_/a_761_249# _310_/D 2.5e-21
C3866 _281_/Y _147_/Y 0.00717f
C3867 _314_/a_1283_n19# _297_/B 2.02e-20
C3868 _314_/a_543_7# _314_/D 0.00149f
C3869 _286_/B _174_/a_109_257# 3.47e-19
C3870 _170_/a_76_159# VGND 0.00734f
C3871 _170_/a_489_373# VPWR 0.0286f
C3872 input4/X _332_/Q 0.00121f
C3873 _341_/a_448_7# _145_/A 3.71e-21
C3874 _322_/a_1108_7# _269_/A 0.00166f
C3875 _162_/X _260_/A 2.22e-19
C3876 cal output41/a_27_7# 0.0119f
C3877 _325_/a_1108_7# _325_/D 0.0576f
C3878 _320_/Q _331_/a_1108_7# 2.83e-21
C3879 _339_/a_761_249# _340_/CLK 7.35e-19
C3880 _163_/a_78_159# _345_/Q 0.0517f
C3881 _166_/Y _147_/Y 9.65e-20
C3882 _323_/a_193_7# _175_/Y 4.9e-19
C3883 _169_/B _306_/a_505_n19# 1.09e-19
C3884 _340_/a_761_249# _337_/Q 1.43e-19
C3885 clkbuf_2_1_0_clk/A VGND 1.58f
C3886 _326_/a_1217_7# repeater43/X 7.16e-19
C3887 _247_/a_199_7# _244_/B 4.28e-19
C3888 _309_/Q _262_/a_113_257# 5.3e-19
C3889 _326_/a_193_7# _331_/a_1108_7# 2.17e-19
C3890 _207_/C _332_/Q 0.123f
C3891 _206_/A _190_/A 0.391f
C3892 output25/a_27_7# _269_/A 0.0109f
C3893 _326_/a_651_373# _217_/X 0.0266f
C3894 _310_/Q VGND 1.01f
C3895 _293_/a_121_257# _254_/Y 0.00129f
C3896 _281_/Y _330_/a_639_7# 1.19e-19
C3897 _283_/A _246_/a_109_257# 0.00204f
C3898 _346_/a_652_n19# _254_/A 1.84e-21
C3899 _343_/CLK _316_/D 7.54e-21
C3900 _345_/a_193_7# _345_/a_381_7# -0.00202f
C3901 _277_/Y _311_/a_27_7# 5.7e-19
C3902 _334_/D _190_/A 1.12e-20
C3903 _342_/a_448_7# _269_/A 0.00617f
C3904 _300_/a_735_7# VGND 0.00543f
C3905 _281_/Y _333_/a_1108_7# 2.39e-20
C3906 _328_/a_651_373# _212_/X 0.00179f
C3907 _328_/a_448_7# _217_/X 2.57e-19
C3908 _301_/X _347_/a_193_7# 0.00932f
C3909 _308_/a_505_n19# _227_/A 0.0621f
C3910 _324_/Q _196_/A 4.1e-19
C3911 _191_/B _295_/a_676_257# 1.57e-19
C3912 output21/a_27_7# _281_/A 2.26e-20
C3913 _173_/a_226_7# _345_/D 2.25e-19
C3914 _173_/a_489_373# _345_/Q 0.00122f
C3915 _299_/X _297_/B 0.0109f
C3916 _283_/Y rstn 0.0695f
C3917 _339_/Q _338_/a_27_7# 0.00126f
C3918 _339_/a_1283_n19# _338_/D 3.17e-19
C3919 _339_/a_543_7# _346_/SET_B 0.00367f
C3920 trim[2] _312_/a_1283_n19# 2.82e-19
C3921 _248_/A _147_/A 7.98e-21
C3922 repeater43/X _334_/a_805_7# -1e-18
C3923 repeater43/a_27_7# _343_/CLK 0.0266f
C3924 _218_/a_93_n19# _304_/X 0.0112f
C3925 _309_/a_761_249# _310_/Q 5.74e-20
C3926 _194_/A _202_/a_250_257# 0.0679f
C3927 _258_/a_76_159# _336_/a_193_7# 1.06e-19
C3928 _258_/a_505_n19# _336_/a_27_7# 0.00142f
C3929 _272_/a_121_257# _217_/A 2.75e-20
C3930 result[1] _315_/a_448_7# 6.14e-20
C3931 _324_/Q _304_/a_591_329# 1.38e-19
C3932 _313_/a_27_7# _313_/a_193_7# -0.33f
C3933 _149_/A _248_/A 2.49e-19
C3934 ctln[4] VGND 0.116f
C3935 _254_/Y _305_/a_505_n19# 6.52e-20
C3936 input1/X _194_/A 2.03e-19
C3937 _271_/Y _227_/A 1.05e-19
C3938 _337_/a_27_7# _337_/a_639_7# -0.0015f
C3939 _309_/a_1108_7# _284_/a_39_257# 7.75e-20
C3940 _235_/a_113_257# VGND 5.21e-19
C3941 _251_/a_79_n19# _162_/X 0.081f
C3942 _146_/C _298_/C 3.14e-20
C3943 _225_/X _333_/Q 3.09e-20
C3944 _147_/A _190_/A 0.0427f
C3945 _320_/Q clkbuf_0_clk/X 0.114f
C3946 _340_/a_448_7# _339_/D 0.00344f
C3947 _334_/a_1462_7# _207_/C 0.00183f
C3948 _273_/A _147_/A 2.32e-20
C3949 _327_/a_193_7# clkbuf_0_clk/X 0.204f
C3950 _258_/S input1/X 0.00338f
C3951 _220_/a_93_n19# _278_/a_68_257# 4.42e-19
C3952 _346_/SET_B _217_/X 0.438f
C3953 output6/a_27_7# VPWR 0.126f
C3954 _340_/a_1283_n19# _202_/a_93_n19# 2.17e-20
C3955 _324_/a_448_7# VPWR -0.00313f
C3956 _324_/a_1283_n19# VGND -0.00818f
C3957 _306_/a_218_334# clkbuf_2_1_0_clk/A 1.06e-19
C3958 _309_/D _201_/a_27_7# 7.33e-20
C3959 _318_/a_1270_373# _242_/B 1.58e-20
C3960 _318_/a_448_7# _318_/D 0.0023f
C3961 _315_/D _314_/D 0.0732f
C3962 _277_/A output19/a_27_7# 2.19e-19
C3963 ctln[1] _334_/a_1270_373# 3.8e-20
C3964 _314_/a_1217_7# VGND 5.56e-20
C3965 _344_/a_1296_7# comp 3.86e-20
C3966 _343_/a_543_7# VGND 0.0217f
C3967 _346_/SET_B _313_/a_805_7# -8.08e-19
C3968 _343_/a_1108_7# VPWR 0.028f
C3969 _340_/a_1283_n19# cal 3.77e-21
C3970 input4/X _339_/a_193_7# 1.72e-20
C3971 _328_/a_27_7# clkbuf_0_clk/X 1.3e-21
C3972 _147_/A _173_/a_556_7# 8.57e-20
C3973 _286_/B _344_/D 1.13e-19
C3974 _344_/a_652_n19# _265_/B 1.64e-19
C3975 _316_/D _331_/a_193_7# 1.21e-20
C3976 _331_/CLK _331_/a_761_249# 2.82e-19
C3977 _273_/A output38/a_27_7# 0.02f
C3978 _236_/B _331_/a_27_7# 3.32e-21
C3979 _340_/a_27_7# _260_/A 2.56e-19
C3980 output29/a_27_7# _316_/D 1.31e-19
C3981 _318_/a_27_7# _318_/a_193_7# -0.0355f
C3982 _216_/A _164_/Y 8.59e-21
C3983 _308_/S _341_/Q 4.2e-20
C3984 _341_/D _145_/A 0.0264f
C3985 _276_/a_150_257# _238_/B 3.57e-20
C3986 _325_/Q _244_/B 0.0419f
C3987 _290_/A _164_/A 0.873f
C3988 _341_/a_193_7# _286_/Y 0.541f
C3989 _345_/a_381_7# VPWR 0.00703f
C3990 _278_/a_68_257# VGND 0.0138f
C3991 _345_/a_1032_373# VGND 0.00904f
C3992 _196_/A _228_/A 1.64e-19
C3993 clkbuf_2_2_0_clk/a_75_172# clkbuf_2_3_0_clk/A 0.0135f
C3994 _143_/a_27_7# _144_/A 8.42e-19
C3995 _346_/Q _286_/B 3.05e-19
C3996 _158_/Y _345_/D 5.62e-20
C3997 _314_/Q _346_/D 5.17e-20
C3998 repeater42/a_27_7# _324_/D 4.82e-19
C3999 _283_/A _330_/a_543_7# 8.19e-19
C4000 _281_/Y _256_/a_80_n19# 0.0086f
C4001 clk _334_/a_761_249# 0.00158f
C4002 _168_/a_481_7# _286_/B 7.22e-20
C4003 _220_/a_93_n19# _220_/a_256_7# -3.48e-20
C4004 _339_/a_1283_n19# _337_/a_1108_7# 7.33e-19
C4005 _339_/a_1108_7# _337_/a_1283_n19# 7.33e-19
C4006 _326_/D _331_/a_27_7# 1.8e-20
C4007 _284_/A _347_/a_27_7# 2.91e-22
C4008 _172_/A _169_/B 0.0181f
C4009 _330_/Q _218_/a_346_7# 5.77e-19
C4010 _307_/a_505_n19# _147_/A 0.0183f
C4011 _321_/Q _246_/B 0.00973f
C4012 _307_/X _307_/a_76_159# 0.00227f
C4013 _275_/Y _299_/X 1.97e-20
C4014 _231_/a_79_n19# _232_/A 0.00251f
C4015 _339_/a_1283_n19# _343_/CLK 9.79e-21
C4016 _323_/a_761_249# _227_/A 6.67e-21
C4017 _257_/a_222_53# _147_/Y 7.54e-20
C4018 _222_/a_346_7# _217_/X 4.26e-19
C4019 _218_/a_256_7# VPWR -3.99e-19
C4020 _218_/a_93_n19# VGND -0.00312f
C4021 _200_/a_584_7# input1/X 7.67e-19
C4022 _333_/a_27_7# _205_/a_79_n19# 4.2e-21
C4023 _198_/a_93_n19# _336_/Q 0.0626f
C4024 _342_/D _269_/A 0.00896f
C4025 _165_/X _162_/X 0.333f
C4026 _147_/Y _297_/Y 0.00762f
C4027 _178_/a_27_7# _147_/A 0.0818f
C4028 _188_/a_76_159# _146_/a_29_271# 6.63e-19
C4029 _342_/a_1283_n19# _175_/Y 0.00135f
C4030 _309_/a_193_7# _309_/Q 1.66e-19
C4031 _329_/a_1108_7# _331_/Q 4.75e-19
C4032 _196_/A _216_/A 0.00965f
C4033 _331_/Q _327_/D 1.86e-19
C4034 _320_/Q _286_/Y 2.32e-20
C4035 _345_/Q _172_/Y 0.0677f
C4036 _281_/Y _332_/a_27_7# 4.32e-19
C4037 _232_/X _326_/Q 0.101f
C4038 _318_/a_193_7# _246_/B 1.81e-21
C4039 _226_/a_297_7# _225_/X 1.57e-19
C4040 _226_/a_382_257# _150_/C -6.49e-21
C4041 _226_/a_79_n19# _226_/X 0.0029f
C4042 _220_/a_256_7# VGND -2.02e-19
C4043 _220_/a_584_7# VPWR -2.88e-19
C4044 _251_/a_215_7# _181_/X 2.61e-20
C4045 _290_/A _312_/D 1.18e-20
C4046 output33/a_27_7# _312_/Q 1.85e-19
C4047 _311_/a_761_249# VPWR 0.0352f
C4048 _327_/a_193_7# _286_/Y 1.06e-20
C4049 _311_/a_27_7# VGND -0.0525f
C4050 repeater43/X _334_/Q 0.138f
C4051 _305_/X _336_/D 0.00259f
C4052 cal _334_/a_193_7# 6.13e-19
C4053 _313_/Q _336_/a_27_7# 7.7e-20
C4054 _325_/a_1108_7# _248_/A 3.4e-20
C4055 _231_/a_512_7# _144_/a_27_7# 4.09e-19
C4056 result[1] _315_/D 1.72e-19
C4057 _313_/D _336_/a_543_7# 5.47e-19
C4058 _145_/A _143_/a_27_7# 1.41e-20
C4059 clk _295_/a_512_7# 0.00603f
C4060 ctln[1] input4/X 0.0702f
C4061 _283_/Y clkbuf_2_0_0_clk/a_75_172# 0.00297f
C4062 repeater42/a_27_7# _218_/a_250_257# 8.13e-21
C4063 output23/a_27_7# VGND 0.102f
C4064 _342_/a_193_7# _298_/A 2.48e-19
C4065 _342_/D _343_/D 1.44e-20
C4066 _318_/Q _234_/B 7.93e-20
C4067 _325_/a_1108_7# _331_/CLK 2.79e-21
C4068 _271_/A VPWR 2.43f
C4069 _337_/a_543_7# _337_/D 3.95e-19
C4070 _318_/Q _321_/a_1283_n19# 3.91e-20
C4071 _200_/a_256_7# _267_/A 4.56e-19
C4072 _167_/X _299_/a_215_7# 5.35e-19
C4073 _165_/X _299_/a_493_257# 2.42e-19
C4074 _316_/Q _318_/a_193_7# 1.77e-21
C4075 _251_/X _162_/X 0.308f
C4076 clk _333_/Q 0.38f
C4077 _335_/a_27_7# VPWR 0.052f
C4078 _197_/X _336_/a_543_7# 0.00871f
C4079 _320_/a_1108_7# clkbuf_2_1_0_clk/A 2.13e-20
C4080 input4/X _192_/B 1.49e-19
C4081 _332_/a_1108_7# _207_/a_27_7# 2.1e-20
C4082 repeater43/X _191_/B 0.0145f
C4083 _304_/S _212_/X 0.0032f
C4084 _342_/Q _333_/a_1283_n19# 6.47e-20
C4085 ctln[1] _207_/C 3.63e-20
C4086 _331_/Q _283_/A 0.0315f
C4087 _327_/a_1462_7# clkbuf_0_clk/X 1.07e-19
C4088 _339_/a_27_7# _339_/a_639_7# -0.0015f
C4089 _271_/A _318_/a_543_7# 1.46e-19
C4090 _273_/A _325_/a_1108_7# 2.13e-20
C4091 _172_/A _170_/a_226_7# 9.73e-19
C4092 _162_/A _284_/A 2.04e-20
C4093 _340_/a_1283_n19# _284_/A 8.15e-20
C4094 _339_/D _190_/A 3.7e-21
C4095 _317_/Q _322_/Q 0.00187f
C4096 _182_/a_79_n19# _283_/A 5.87e-20
C4097 _289_/a_39_257# _310_/a_1108_7# 4.2e-19
C4098 _216_/X _284_/A 1.01e-19
C4099 _318_/a_651_373# VGND 0.00316f
C4100 _318_/a_639_7# VPWR 8.76e-19
C4101 _192_/B _207_/C 5e-19
C4102 _286_/B _340_/D 1.07e-19
C4103 _244_/B _326_/Q 0.00426f
C4104 _145_/A _343_/CLK 4.9e-21
C4105 _144_/a_27_7# _223_/a_93_n19# 8.18e-21
C4106 _276_/a_150_257# _331_/CLK 8.78e-19
C4107 _294_/Y _164_/Y 0.00341f
C4108 _346_/a_193_7# _303_/A 9.16e-21
C4109 _307_/a_535_334# _145_/A 3.88e-19
C4110 cal _332_/Q 1.18e-19
C4111 repeater43/X _317_/a_543_7# 0.0395f
C4112 _309_/a_448_7# VPWR 0.00387f
C4113 _309_/a_1283_n19# VGND -4.05e-19
C4114 _334_/Q _191_/B 5.67e-20
C4115 _340_/a_27_7# _340_/Q 0.0112f
C4116 _340_/a_193_7# _194_/X 0.00111f
C4117 _313_/a_805_7# _147_/A 0.00237f
C4118 clkbuf_0_clk/X _319_/a_761_249# 1.01e-20
C4119 input1/X _201_/a_27_7# 2.16e-20
C4120 _315_/a_761_249# _317_/D 8e-20
C4121 _258_/a_76_159# _299_/X 1.42e-20
C4122 _227_/A _154_/a_27_7# 0.00529f
C4123 _255_/B _192_/a_68_257# 1.99e-20
C4124 result[5] _321_/Q 6.24e-20
C4125 output11/a_27_7# ctln[6] 0.00515f
C4126 ctln[7] _227_/A 4.53e-21
C4127 _281_/Y _260_/B 0.00224f
C4128 _164_/A _310_/a_27_7# 3.23e-20
C4129 _306_/X _336_/Q 3.09e-20
C4130 _220_/a_93_n19# _328_/D 0.0327f
C4131 _342_/a_1283_n19# _341_/Q 5.56e-20
C4132 _321_/a_761_249# _322_/Q 0.00282f
C4133 _321_/a_193_7# _331_/Q 2.67e-20
C4134 _307_/a_76_159# _183_/a_27_7# 1.38e-21
C4135 repeater43/X _331_/a_448_7# 9.11e-19
C4136 _327_/a_448_7# _281_/A 4.63e-22
C4137 _296_/Y _147_/A 0.0163f
C4138 _316_/a_651_373# _228_/A 2.72e-21
C4139 _341_/D _324_/Q 6.28e-21
C4140 _283_/A _333_/a_805_7# 0.00216f
C4141 _331_/a_27_7# _331_/a_193_7# -0.301f
C4142 _324_/a_193_7# _181_/a_27_7# 1.2e-20
C4143 ctlp[5] clkbuf_2_1_0_clk/A 0.0546f
C4144 _229_/a_226_257# sample 3.59e-20
C4145 _327_/a_543_7# _281_/Y 0.00174f
C4146 _309_/a_27_7# _309_/a_448_7# -0.00642f
C4147 _331_/a_1283_n19# _327_/Q 6.46e-21
C4148 _331_/a_543_7# _212_/X 5.63e-20
C4149 _162_/X _232_/A 1.37e-19
C4150 _263_/B clkc 9.59e-20
C4151 _325_/a_193_7# _304_/S 5.28e-19
C4152 _323_/a_27_7# VPWR 0.0802f
C4153 _330_/D VPWR 0.262f
C4154 _183_/a_1241_257# _178_/a_27_7# 1.77e-21
C4155 _333_/a_1108_7# _335_/Q 3.5e-19
C4156 _323_/Q _226_/X 2.61e-20
C4157 _192_/B _150_/C 1.14e-19
C4158 _146_/a_29_271# _147_/A 0.0349f
C4159 _188_/a_218_334# _146_/C 6.25e-19
C4160 _319_/Q _238_/B 0.104f
C4161 _149_/a_27_7# _304_/S 7.41e-19
C4162 _320_/a_27_7# _297_/B 0.619f
C4163 input1/X _337_/a_27_7# 2.54e-21
C4164 cal _337_/a_193_7# 4.14e-19
C4165 _294_/A _312_/Q 1.11e-19
C4166 _185_/A _176_/a_27_7# 0.00998f
C4167 _254_/B _153_/A 0.0369f
C4168 _146_/a_29_271# _149_/A 4.86e-19
C4169 _306_/a_218_7# VGND -7.49e-19
C4170 _290_/A _292_/A 1.12f
C4171 _328_/D VGND 0.224f
C4172 _256_/a_209_257# _255_/B 2.31e-19
C4173 clkbuf_0_clk/a_110_7# _147_/A 1.23e-19
C4174 output37/a_27_7# _285_/Y 0.0302f
C4175 _311_/a_1217_7# VGND 5.4e-20
C4176 cal _334_/a_1462_7# 5.68e-20
C4177 _313_/Q _336_/a_1217_7# 4.61e-21
C4178 ctlp[6] _330_/D 0.0041f
C4179 _326_/a_1283_n19# _319_/Q 8.76e-22
C4180 _214_/a_109_257# _217_/A 0.0459f
C4181 _255_/B _177_/A 3.05e-19
C4182 _290_/A _160_/A 2.06e-19
C4183 _186_/a_79_n19# VPWR 0.03f
C4184 _235_/a_199_7# _232_/X 0.00146f
C4185 _325_/Q _223_/a_256_7# 0.00317f
C4186 _324_/a_1108_7# _172_/A 3.03e-21
C4187 _335_/a_193_7# _335_/a_1283_n19# -6.53e-19
C4188 repeater43/X result[6] 0.00659f
C4189 _285_/A _309_/Q 0.0251f
C4190 clkbuf_1_1_0_clk/a_75_172# _299_/a_215_7# 4.39e-19
C4191 _326_/Q _241_/a_113_257# 1.32e-21
C4192 _329_/a_27_7# _216_/X 2.69e-19
C4193 _188_/S _315_/D 8.1e-20
C4194 trim[1] _310_/a_1283_n19# 2.52e-19
C4195 _250_/a_78_159# _190_/A 0.00874f
C4196 _328_/a_543_7# _319_/Q 0.0338f
C4197 _232_/a_27_7# VPWR 0.148f
C4198 _180_/a_183_257# _286_/Y 4.04e-19
C4199 _335_/a_639_7# VGND 3.11e-19
C4200 _335_/a_1217_7# VPWR 9.35e-20
C4201 _184_/a_439_7# VGND 3.17e-19
C4202 _341_/a_193_7# _269_/A 0.0134f
C4203 _343_/a_193_7# _342_/a_193_7# 4.66e-20
C4204 _343_/a_761_249# _342_/a_27_7# 5.16e-21
C4205 _329_/a_193_7# _320_/Q 3.82e-20
C4206 _329_/a_27_7# _329_/Q 5.03e-20
C4207 _324_/Q _143_/a_27_7# 5.96e-19
C4208 _183_/a_553_257# _144_/A 3.18e-19
C4209 _320_/Q _328_/Q 0.782f
C4210 _339_/a_543_7# _339_/D 0.00639f
C4211 _336_/Q _147_/Y 0.196f
C4212 _328_/a_761_249# _329_/D 2.41e-20
C4213 clkbuf_2_1_0_clk/A _330_/a_27_7# 9.24e-20
C4214 _320_/a_1283_n19# _279_/A 3.96e-19
C4215 _326_/D _324_/Q 1.3e-20
C4216 output31/a_27_7# trim[1] 5.93e-20
C4217 _329_/a_761_249# _327_/a_27_7# 0.00111f
C4218 _329_/a_193_7# _327_/a_193_7# 8.38e-19
C4219 _327_/a_193_7# _328_/Q 1.22e-19
C4220 _338_/a_639_7# _340_/Q 0.00108f
C4221 _338_/D _195_/a_27_257# 8.44e-19
C4222 _338_/a_805_7# _194_/X 6.71e-19
C4223 cal _226_/a_382_257# 3.97e-19
C4224 input1/X _226_/a_79_n19# 4.93e-20
C4225 _182_/a_215_7# _175_/Y 0.0135f
C4226 _325_/a_639_7# repeater43/X -5.17e-19
C4227 _341_/Q _231_/a_676_257# 3.48e-20
C4228 _209_/X _333_/a_651_373# 5.97e-20
C4229 _317_/a_27_7# _317_/a_448_7# -0.00346f
C4230 _341_/a_543_7# _185_/A 1.51e-20
C4231 _341_/D _228_/A 1.45e-19
C4232 _325_/a_651_373# _327_/Q 9.03e-20
C4233 _178_/a_27_7# _150_/a_27_7# 0.00699f
C4234 _285_/A _311_/a_193_7# 2.64e-20
C4235 _344_/a_1032_373# _160_/X 5.54e-20
C4236 _338_/Q _267_/A 0.2f
C4237 _293_/a_39_257# VGND 0.0247f
C4238 _329_/a_27_7# _328_/a_193_7# 2.35e-21
C4239 _329_/a_193_7# _328_/a_27_7# 1.88e-21
C4240 _328_/a_27_7# _328_/Q 0.00924f
C4241 _269_/A _316_/a_761_249# 0.00181f
C4242 _340_/a_1217_7# _340_/Q 0.00103f
C4243 _340_/a_805_7# _306_/S 6.43e-19
C4244 _340_/a_639_7# _193_/Y 8.12e-19
C4245 _340_/a_1462_7# _194_/X 4.65e-19
C4246 ctln[5] _193_/Y 8.74e-19
C4247 _279_/Y _340_/D 0.123f
C4248 _320_/Q _269_/A 0.17f
C4249 _336_/a_805_7# _147_/Y 0.00215f
C4250 _294_/Y _165_/a_78_159# 4.28e-20
C4251 clkbuf_2_3_0_clk/A cal 0.014f
C4252 _255_/X _194_/A 0.0104f
C4253 _322_/a_1283_n19# _321_/Q 0.016f
C4254 _324_/Q _343_/CLK 0.0124f
C4255 _341_/a_1283_n19# _255_/B 1.49e-20
C4256 _283_/Y VPWR 0.355f
C4257 _232_/X _279_/A 0.214f
C4258 ctlp[5] _278_/a_68_257# 0.0169f
C4259 _164_/A _310_/a_1217_7# 3.14e-20
C4260 _270_/a_39_257# _316_/a_193_7# 1.65e-19
C4261 _271_/A _323_/a_1108_7# 6.26e-19
C4262 _339_/Q _337_/a_805_7# 4.44e-19
C4263 _319_/Q _248_/A 0.00773f
C4264 _346_/a_1602_7# _346_/Q 0.0244f
C4265 _346_/a_1182_221# _166_/Y 0.00401f
C4266 _281_/Y _333_/Q 5.82e-20
C4267 _311_/a_543_7# _311_/D 2.07e-19
C4268 _325_/Q _177_/A 1.09e-19
C4269 ctln[6] _207_/X 4.49e-19
C4270 _322_/a_27_7# VGND 0.0073f
C4271 _322_/a_761_249# VPWR 0.0184f
C4272 _325_/a_1108_7# _296_/Y 3.28e-20
C4273 _188_/a_439_7# _286_/Y 1.61e-19
C4274 _258_/S _255_/X 1.45e-21
C4275 _258_/S _257_/a_448_7# 2.99e-20
C4276 _346_/a_27_7# _167_/X 0.00339f
C4277 _170_/a_489_373# _147_/Y 3.2e-19
C4278 _337_/a_193_7# _284_/A 3.87e-20
C4279 _308_/a_76_159# _188_/S 1.91e-19
C4280 _319_/Q _331_/CLK 0.778f
C4281 _320_/a_639_7# VPWR 1.48e-19
C4282 _320_/a_651_373# VGND 0.0112f
C4283 _323_/a_1217_7# VPWR 2.06e-19
C4284 _323_/a_639_7# VGND 2.63e-19
C4285 _238_/a_109_257# VPWR 3.11e-19
C4286 _258_/S clkc 0.00118f
C4287 _283_/A _332_/a_1108_7# 9.57e-21
C4288 _322_/a_1283_n19# _318_/a_193_7# 5.9e-22
C4289 _146_/C _150_/C 0.0942f
C4290 _305_/a_218_334# VPWR 6.55e-20
C4291 _305_/a_76_159# VGND 0.0184f
C4292 _214_/a_109_7# VGND 3.84e-19
C4293 _344_/a_1182_221# VGND -0.00158f
C4294 _344_/a_1602_7# VPWR 0.00546f
C4295 _200_/a_93_n19# _283_/A 4.06e-20
C4296 _232_/X _220_/a_346_7# 1.88e-19
C4297 _294_/Y trim[3] 2.99e-20
C4298 _280_/a_68_257# _212_/X 3.67e-21
C4299 _143_/a_27_7# _228_/A 0.0796f
C4300 _346_/SET_B _221_/a_346_7# 5.82e-21
C4301 _320_/a_1217_7# _297_/B 1.88e-19
C4302 _306_/S _340_/CLK 0.0865f
C4303 _273_/A _319_/Q 1.13e-19
C4304 _332_/a_27_7# _335_/Q 0.0103f
C4305 _286_/B _209_/X 0.0207f
C4306 _157_/A _150_/C 0.00833f
C4307 _326_/Q _223_/a_256_7# 4.63e-19
C4308 _260_/A _313_/a_1283_n19# 2.05e-20
C4309 _285_/A _309_/a_1108_7# 6.87e-20
C4310 _227_/A _333_/a_761_249# 6.43e-21
C4311 _216_/X _144_/a_27_7# 2.85e-20
C4312 _257_/a_222_53# _260_/B 0.0399f
C4313 _325_/a_193_7# _325_/a_448_7# -0.00831f
C4314 _277_/A _299_/a_215_7# 1.6e-19
C4315 _331_/D _217_/A 0.0151f
C4316 _252_/a_27_7# _227_/A 5.12e-20
C4317 _337_/a_1108_7# _195_/a_27_257# 1.1e-21
C4318 output25/a_27_7# _318_/a_27_7# 2.21e-20
C4319 output12/a_27_7# _206_/A 0.00854f
C4320 _325_/Q _325_/D 0.0472f
C4321 _292_/A _310_/a_27_7# 1.1e-20
C4322 _342_/a_193_7# VGND 0.00381f
C4323 _342_/a_543_7# VPWR 0.0121f
C4324 _329_/a_1217_7# _216_/X 9.91e-20
C4325 _297_/A _314_/a_193_7# 3.35e-19
C4326 _343_/CLK _195_/a_27_257# 1.74e-19
C4327 _258_/S _264_/a_199_7# 0.00172f
C4328 _250_/X _190_/A 2.18e-19
C4329 _288_/A _310_/D 0.00506f
C4330 output32/a_27_7# _310_/Q 4.03e-19
C4331 _286_/B _265_/B 1.42e-20
C4332 _182_/a_79_n19# _298_/B 0.00374f
C4333 _198_/a_584_7# VGND 1.39e-19
C4334 _182_/a_215_7# _341_/Q 0.00535f
C4335 _267_/A _313_/a_1108_7# 2.1e-21
C4336 _219_/a_250_257# _217_/X 0.0456f
C4337 input1/X _323_/Q 1.81e-20
C4338 cal _192_/B 0.0108f
C4339 _162_/X _310_/D 1.68e-20
C4340 _322_/a_27_7# output27/a_27_7# 0.00187f
C4341 ctlp[1] _321_/a_761_249# 7.58e-20
C4342 _319_/Q _319_/a_1108_7# 0.0538f
C4343 _329_/a_1217_7# _329_/Q 1.05e-19
C4344 _290_/A _273_/A 0.0251f
C4345 _287_/a_39_257# _310_/D 0.00939f
C4346 repeater43/X result[4] 3.3e-19
C4347 _343_/CLK _228_/A 7.15e-20
C4348 _326_/D _216_/A 0.111f
C4349 ctlp[2] trimb[3] 0.0941f
C4350 _338_/Q _194_/X 0.358f
C4351 _346_/SET_B _193_/Y 0.506f
C4352 _320_/a_27_7# _320_/a_193_7# -0.328f
C4353 _323_/a_193_7# _323_/a_1283_n19# -7.11e-33
C4354 _157_/A _302_/a_77_159# 0.017f
C4355 _294_/A _340_/CLK 0.00229f
C4356 _216_/A _222_/a_256_7# 6.48e-19
C4357 _254_/A _267_/A 0.0251f
C4358 _332_/a_761_249# _153_/a_215_257# 0.00322f
C4359 _297_/B _172_/B 2.51e-20
C4360 _336_/a_193_7# _194_/A 5.97e-20
C4361 _256_/a_80_n19# _336_/Q 2.97e-19
C4362 clkbuf_2_3_0_clk/A _284_/A 0.00807f
C4363 _320_/a_1108_7# _328_/D 8.5e-20
C4364 _304_/a_257_159# _326_/Q 7.48e-19
C4365 _216_/A _313_/a_193_7# 0.587f
C4366 _328_/a_1217_7# _328_/Q 0.00103f
C4367 _157_/a_27_7# _297_/a_27_257# 1.81e-20
C4368 _181_/X _298_/A 0.1f
C4369 ctln[7] _335_/a_543_7# 0.0297f
C4370 _283_/Y _335_/a_1108_7# 1.21e-19
C4371 _182_/a_510_7# _227_/A 0.00123f
C4372 _258_/S _336_/a_193_7# 4.42e-19
C4373 result[2] _316_/a_448_7# 3.09e-20
C4374 _290_/A trim[4] 4.75e-20
C4375 _203_/a_303_7# VGND 4e-19
C4376 _286_/B _336_/a_1270_373# 8.78e-20
C4377 _242_/A _316_/a_1283_n19# 1.06e-20
C4378 _319_/a_761_249# _328_/Q 1.16e-19
C4379 _312_/a_27_7# VPWR 0.103f
C4380 _275_/A _167_/X 4.77e-21
C4381 _267_/B _344_/Q 9.06e-21
C4382 ctlp[0] _322_/D 0.00119f
C4383 _346_/a_1296_7# _166_/Y 6.42e-19
C4384 _339_/Q _337_/Q 0.0328f
C4385 _311_/a_805_7# _311_/Q 9.65e-20
C4386 _292_/A output36/a_27_7# 2.83e-19
C4387 _326_/a_1270_373# _283_/A 1.06e-19
C4388 _231_/a_512_7# _315_/D 0.0429f
C4389 _307_/a_505_n19# _250_/X 0.00216f
C4390 _307_/a_535_334# _216_/A 2.63e-20
C4391 _340_/a_193_7# _336_/a_543_7# 4.64e-22
C4392 _340_/a_543_7# _336_/a_193_7# 3.67e-19
C4393 _340_/a_1283_n19# _336_/a_27_7# 1.56e-21
C4394 _346_/a_1032_373# _167_/a_27_257# 0.00142f
C4395 _172_/A _306_/a_439_7# 2.41e-22
C4396 _231_/a_79_n19# VPWR 0.0224f
C4397 _226_/X sample 5.54e-20
C4398 _332_/a_543_7# _209_/a_27_257# 4.68e-21
C4399 _309_/D _267_/A 0.00574f
C4400 _313_/a_1270_373# _284_/A 1.12e-19
C4401 _330_/Q _330_/a_1108_7# 0.00121f
C4402 _225_/B _347_/a_27_7# 1.64e-19
C4403 _326_/a_543_7# _242_/A 0.0337f
C4404 _316_/D _247_/a_113_257# 1.39e-19
C4405 input4/X _340_/Q 7.67e-19
C4406 _337_/Q _202_/a_256_7# 7.67e-19
C4407 _308_/S _188_/S 0.00339f
C4408 _283_/A _340_/CLK 0.0468f
C4409 _183_/a_471_7# _146_/C 6.89e-20
C4410 input3/a_27_7# _298_/X 4.24e-21
C4411 en output41/a_27_7# 0.00129f
C4412 _250_/a_493_257# _192_/B 6.84e-20
C4413 _281_/A _331_/a_193_7# 1.72e-20
C4414 _250_/X _178_/a_27_7# 7.05e-21
C4415 _344_/a_1296_7# VGND 7.71e-20
C4416 _326_/a_1283_n19# _325_/Q 4.06e-21
C4417 result[0] result[2] 0.002f
C4418 _196_/A _153_/A 9.79e-21
C4419 _330_/a_761_249# VGND 0.0057f
C4420 _330_/a_1283_n19# VPWR 0.0431f
C4421 _343_/Q _298_/A 2.09e-21
C4422 _183_/a_553_257# _324_/Q 0.0112f
C4423 _183_/a_471_7# _157_/A 3.63e-19
C4424 _281_/Y _212_/X 0.0492f
C4425 result[3] VGND 0.144f
C4426 _345_/a_193_7# _288_/A 2.17e-20
C4427 _286_/B clkbuf_2_1_0_clk/A 0.0513f
C4428 _326_/Q _325_/D 0.0231f
C4429 _186_/a_382_257# _188_/S 1.93e-19
C4430 clkbuf_0_clk/a_110_7# _250_/a_78_159# 5.01e-19
C4431 _189_/a_27_7# _190_/A 0.074f
C4432 _333_/a_27_7# VPWR 0.0567f
C4433 comp _346_/SET_B 7.13e-21
C4434 _345_/a_193_7# _162_/X 1.39e-20
C4435 _306_/S _313_/a_543_7# 1.84e-19
C4436 _288_/A _266_/a_113_257# 0.00236f
C4437 _255_/B _190_/A 0.0279f
C4438 _337_/a_1283_n19# _340_/D 8.28e-21
C4439 _337_/a_448_7# _193_/Y 2.56e-21
C4440 _318_/Q _318_/a_651_373# 0.0266f
C4441 _257_/a_79_159# _190_/A 8.27e-19
C4442 _335_/a_805_7# _335_/D 5.87e-19
C4443 _342_/a_1462_7# VGND -8.49e-19
C4444 _192_/B _284_/A 2.78e-20
C4445 _319_/Q _217_/X 0.0063f
C4446 _211_/a_109_257# _153_/B 0.00129f
C4447 _252_/a_27_7# _297_/B 0.00359f
C4448 _248_/B _347_/D 8.54e-19
C4449 _286_/B _300_/a_735_7# 3.92e-19
C4450 _196_/A _300_/a_383_7# 2.38e-21
C4451 _294_/Y _273_/Y 0.00183f
C4452 _182_/X _298_/B 0.00951f
C4453 _329_/a_639_7# _331_/CLK 6.21e-19
C4454 repeater43/X clkbuf_1_0_0_clk/a_75_172# 0.00134f
C4455 _329_/D _212_/X 0.00574f
C4456 _314_/a_543_7# _347_/a_27_7# 0.00197f
C4457 _254_/A _194_/X 1.49e-20
C4458 _165_/X _345_/Q 0.00127f
C4459 _167_/X _345_/D 1.85e-21
C4460 _325_/a_27_7# _284_/A 8.06e-21
C4461 _275_/Y _172_/B 0.0334f
C4462 _304_/S _306_/S 4.71e-19
C4463 ctlp[2] VPWR 0.0612f
C4464 _333_/D _154_/A 0.0136f
C4465 _254_/Y _340_/CLK 0.00848f
C4466 _162_/a_27_7# _267_/A 4.48e-19
C4467 _274_/a_121_257# _242_/A 9.54e-19
C4468 _216_/A _331_/a_193_7# 4.67e-21
C4469 _181_/X _215_/A 0.00986f
C4470 _271_/A _233_/a_199_7# 2.24e-19
C4471 _171_/a_78_159# _171_/a_292_257# -1.09e-21
C4472 _273_/A _310_/a_27_7# 2.33e-21
C4473 _340_/a_1108_7# _336_/Q 4.43e-20
C4474 _341_/a_651_373# _298_/A 0.00722f
C4475 rstn _332_/D 2.12e-19
C4476 _332_/a_543_7# _153_/A 0.00278f
C4477 _332_/a_193_7# _154_/A 7.37e-20
C4478 _229_/a_226_257# _175_/Y 8.21e-19
C4479 _345_/a_1182_221# _164_/Y 0.0132f
C4480 trim[0] _311_/Q 4.37e-19
C4481 _306_/S _225_/X 0.0442f
C4482 _193_/Y _147_/A 0.00185f
C4483 _329_/a_27_7# _327_/Q 2.6e-20
C4484 _344_/a_193_7# _344_/a_1032_373# -9.67e-21
C4485 _344_/a_27_7# _344_/a_1602_7# -2.39e-19
C4486 _307_/X _306_/S 0.0127f
C4487 _322_/Q VGND 0.97f
C4488 _254_/A _167_/X 0.0147f
C4489 _200_/a_250_257# clkbuf_2_0_0_clk/a_75_172# 1.13e-20
C4490 _301_/a_149_7# _346_/SET_B 1.41e-20
C4491 ctlp[7] clkbuf_2_1_0_clk/A 2.07e-19
C4492 _281_/Y _325_/a_193_7# 4.85e-19
C4493 ctln[3] _312_/a_27_7# 4.14e-20
C4494 _275_/Y _312_/a_761_249# 0.00503f
C4495 input2/a_27_7# _288_/Y 1.34e-21
C4496 _153_/B _203_/a_80_n19# 3.15e-20
C4497 _325_/Q _248_/A 1.91e-19
C4498 _182_/a_297_257# VPWR -0.00288f
C4499 _275_/A clkbuf_1_1_0_clk/a_75_172# 0.0366f
C4500 result[2] _316_/D 2.98e-19
C4501 _309_/D _194_/X 2.09e-20
C4502 output8/a_27_7# _297_/Y 0.00995f
C4503 _339_/a_651_373# _306_/S 0.00437f
C4504 _255_/B _307_/a_505_n19# 0.0142f
C4505 _312_/a_1217_7# VPWR 2.06e-20
C4506 _229_/a_76_159# _298_/A 1.67e-19
C4507 _160_/X _299_/a_292_257# 7.89e-19
C4508 clkbuf_0_clk/X _267_/A 2e-19
C4509 _319_/a_193_7# _319_/D 0.00551f
C4510 _346_/a_27_7# _277_/A 2.67e-20
C4511 _288_/A VPWR 0.849f
C4512 _325_/Q _331_/CLK 0.0158f
C4513 _204_/Y _332_/Q 0.142f
C4514 _335_/Q _333_/Q 0.233f
C4515 repeater42/a_27_7# _331_/Q 4.09e-20
C4516 _300_/a_301_257# _347_/a_1108_7# 1.78e-20
C4517 _258_/a_505_n19# _313_/D 2.11e-20
C4518 result[4] result[6] 6.22e-19
C4519 _161_/Y _171_/a_78_159# 0.0343f
C4520 _296_/Y _250_/X 1.36e-19
C4521 _255_/a_30_13# _191_/B 1.66e-19
C4522 _181_/X _304_/X 0.01f
C4523 _316_/a_1283_n19# _315_/a_1108_7# 4.22e-19
C4524 _162_/X VPWR 6.11f
C4525 ctln[2] trim[2] 0.00175f
C4526 _326_/a_1283_n19# _326_/Q 0.027f
C4527 clk _207_/a_27_7# 6.14e-21
C4528 _287_/a_39_257# VPWR 0.0341f
C4529 _232_/X _214_/a_373_7# 3.78e-19
C4530 cal _260_/A 0.00839f
C4531 output24/a_27_7# repeater43/X 0.00108f
C4532 _298_/A _204_/a_27_7# 2.55e-20
C4533 _337_/Q _336_/D 1.17e-19
C4534 _273_/A _325_/Q 3.96e-20
C4535 _200_/a_93_n19# _194_/a_27_7# 2.92e-21
C4536 ctlp[3] VGND 0.182f
C4537 _197_/a_27_7# _260_/A 0.0201f
C4538 _321_/a_1108_7# _248_/A 1.8e-20
C4539 _279_/Y _314_/a_27_7# 0.0145f
C4540 clkbuf_2_1_0_clk/A _338_/a_1108_7# 6.06e-20
C4541 _197_/X _311_/D 0.00244f
C4542 _304_/a_257_159# _324_/D 3.75e-21
C4543 _335_/a_1108_7# _333_/a_27_7# 1.3e-20
C4544 _234_/B _316_/D 5.09e-21
C4545 _343_/a_1283_n19# _177_/A 2.89e-21
C4546 _321_/D _321_/a_193_7# 0.0044f
C4547 _232_/X _246_/a_109_257# 1.77e-19
C4548 _343_/a_761_249# _298_/X 2.27e-20
C4549 _343_/a_27_7# valid 0.02f
C4550 _321_/a_1108_7# _331_/CLK 0.0574f
C4551 _346_/SET_B _310_/a_1270_373# -2.06e-19
C4552 _338_/Q _310_/a_1108_7# 0.00143f
C4553 _325_/a_1283_n19# _216_/A 4.98e-19
C4554 _333_/a_1217_7# VPWR 2.92e-20
C4555 _333_/a_639_7# VGND 0.00128f
C4556 _273_/A output36/a_27_7# 0.018f
C4557 cal _261_/A 1.04e-20
C4558 input1/X _267_/A 0.632f
C4559 _242_/A _319_/a_1283_n19# 0.0097f
C4560 _206_/A _205_/a_297_7# 4.92e-19
C4561 _294_/A _267_/B 3.23e-19
C4562 _251_/X _150_/C 3.58e-21
C4563 _337_/D _193_/Y 0.00461f
C4564 _299_/a_78_159# VGND 6.28e-19
C4565 _299_/a_493_257# VPWR -3.53e-19
C4566 _315_/Q _315_/a_1108_7# 0.00728f
C4567 _343_/a_193_7# _343_/Q 1.87e-19
C4568 clkbuf_0_clk/X _221_/a_93_n19# 0.00625f
C4569 _315_/D _347_/a_27_7# 0.019f
C4570 _174_/a_27_257# _344_/D 0.05f
C4571 _174_/a_373_7# _344_/Q 0.00157f
C4572 input1/X sample 0.00181f
C4573 _336_/a_1108_7# _340_/CLK 1.05e-20
C4574 _258_/S _299_/X 2.12e-21
C4575 _153_/a_403_257# _333_/Q 6.99e-19
C4576 _153_/a_487_257# _332_/Q 0.00145f
C4577 _277_/A _319_/a_27_7# 0.00252f
C4578 _304_/S _283_/A 0.071f
C4579 _324_/a_1108_7# _325_/D 8.31e-19
C4580 _157_/A _284_/A 0.203f
C4581 _263_/B _311_/a_1283_n19# 1.07e-19
C4582 _269_/A _323_/Q 1.28e-20
C4583 input4/X rstn 0.13f
C4584 _346_/D _347_/a_1283_n19# 6.31e-21
C4585 _324_/D _325_/D 2.08e-21
C4586 _312_/D _311_/a_193_7# 8.44e-21
C4587 _346_/a_476_7# _169_/Y 5.6e-19
C4588 _283_/A _225_/X 0.00526f
C4589 _341_/D _315_/a_761_249# 1.52e-20
C4590 _307_/X _283_/A 0.00789f
C4591 _318_/Q _322_/a_27_7# 3.8e-22
C4592 _254_/A _301_/a_51_257# 0.0118f
C4593 _309_/a_1108_7# _164_/A 0.00157f
C4594 _145_/A _247_/a_113_257# 2.31e-19
C4595 _342_/a_761_249# _244_/B 5.12e-20
C4596 _254_/Y _313_/a_543_7# 8.85e-21
C4597 _342_/a_27_7# _317_/D 1.6e-19
C4598 _248_/A _326_/Q 0.341f
C4599 _183_/a_27_7# _306_/S 0.00609f
C4600 _202_/a_584_7# _284_/A 5.98e-19
C4601 _214_/a_109_257# _331_/D 4.71e-20
C4602 clk _306_/S 0.0387f
C4603 _304_/S _248_/B 0.674f
C4604 _150_/C _205_/a_79_n19# 1.53e-20
C4605 rstn _207_/C 0.102f
C4606 _343_/D _323_/Q 1.75e-19
C4607 _328_/a_1283_n19# clkbuf_2_1_0_clk/A 1.07e-20
C4608 _277_/A _275_/A 0.0773f
C4609 _286_/Y sample 0.178f
C4610 _346_/SET_B _336_/a_448_7# 0.00126f
C4611 output18/a_27_7# output19/a_27_7# 3.81e-21
C4612 _331_/CLK _326_/Q 0.0313f
C4613 output37/a_27_7# _162_/A 0.0117f
C4614 _181_/X VGND 0.943f
C4615 _339_/D _193_/Y 0.0191f
C4616 _345_/a_1182_221# _165_/a_78_159# 1.58e-19
C4617 _255_/B _296_/Y 0.234f
C4618 _315_/a_1283_n19# _248_/A 2.86e-21
C4619 _188_/a_76_159# _298_/A 0.0292f
C4620 _196_/A _314_/Q 2.04e-20
C4621 _230_/a_27_7# _317_/a_193_7# 9.72e-19
C4622 _260_/A _284_/A 0.692f
C4623 _232_/A _150_/C 0.00609f
C4624 _273_/A _326_/Q 0.205f
C4625 _216_/X _315_/D 2.83e-19
C4626 output35/a_27_7# _310_/D 2.56e-19
C4627 _340_/a_27_7# VPWR 0.0575f
C4628 _300_/Y _347_/a_1108_7# 0.00948f
C4629 _337_/a_193_7# _199_/a_250_257# 1.02e-19
C4630 _340_/Q _202_/a_93_n19# 1.41e-19
C4631 _194_/X _202_/a_250_257# 0.0017f
C4632 _185_/A _149_/a_27_7# 8.11e-21
C4633 _313_/D _313_/Q 5.73e-19
C4634 _304_/a_288_7# VGND 2.65e-19
C4635 _161_/Y _172_/B 0.103f
C4636 _255_/B _146_/a_29_271# 1.6e-19
C4637 _342_/Q _192_/B 0.0891f
C4638 _248_/A _314_/a_193_7# 5.42e-21
C4639 _167_/X clkbuf_0_clk/X 0.0168f
C4640 _283_/A _331_/a_543_7# 6.41e-19
C4641 _343_/a_193_7# _229_/a_76_159# 4.03e-19
C4642 _343_/a_27_7# _229_/a_226_7# 5.24e-20
C4643 _340_/CLK _194_/a_27_7# 3.75e-19
C4644 result[7] _269_/A 0.0035f
C4645 _271_/A _176_/a_27_7# 1.96e-21
C4646 cal _340_/Q 0.0326f
C4647 _237_/a_113_257# VGND 5.12e-19
C4648 _221_/a_93_n19# _286_/Y 0.0817f
C4649 input1/X _194_/X 0.254f
C4650 _326_/Q _222_/a_93_n19# 0.0159f
C4651 _309_/a_193_7# _312_/Q 2.88e-20
C4652 _342_/D _186_/a_297_7# 2.03e-19
C4653 _325_/a_27_7# _342_/Q 3.94e-22
C4654 _317_/a_193_7# _232_/A 1.13e-19
C4655 _325_/a_761_249# _255_/B 2.39e-20
C4656 _313_/Q _197_/X 0.00194f
C4657 _242_/A _212_/X 0.0193f
C4658 _301_/X _306_/S 1.49e-20
C4659 _273_/A output39/a_27_7# 0.00274f
C4660 _197_/a_27_7# _340_/Q 5.61e-20
C4661 _346_/a_1182_221# _170_/a_489_373# 2.15e-21
C4662 _165_/a_493_257# _160_/X 7.76e-19
C4663 _344_/a_956_373# _172_/B 9.04e-19
C4664 _316_/D _224_/a_250_257# 1.32e-19
C4665 _343_/Q VGND 0.298f
C4666 _320_/Q _318_/a_27_7# 2.77e-19
C4667 _298_/C VPWR 1.74f
C4668 _292_/A _309_/Q 0.00538f
C4669 _345_/a_1602_7# _160_/A 3.53e-19
C4670 _338_/Q _199_/a_584_7# 0.00213f
C4671 result[1] _268_/a_39_257# 1.14e-19
C4672 _254_/a_109_257# _265_/B 8.8e-20
C4673 ctlp[1] VGND 0.32f
C4674 _309_/Q _160_/A 1.61e-20
C4675 _327_/a_448_7# _217_/A 2.87e-20
C4676 _327_/a_651_373# _304_/X 5.14e-21
C4677 _329_/a_543_7# clkbuf_0_clk/X 9.68e-22
C4678 _332_/a_1283_n19# VGND 0.0485f
C4679 _332_/a_448_7# VPWR 0.0014f
C4680 _300_/a_301_257# _346_/SET_B 0.00723f
C4681 _347_/a_1108_7# VGND 0.00409f
C4682 _347_/a_651_373# VPWR -0.0085f
C4683 _326_/a_651_373# _304_/X 0.00245f
C4684 _200_/a_250_257# VPWR 0.0346f
C4685 _292_/Y trimb[2] 5.96e-20
C4686 _206_/A _298_/A 2.75e-20
C4687 _154_/A _190_/A 0.418f
C4688 _277_/A _319_/a_1217_7# 1.27e-19
C4689 repeater43/X _321_/a_639_7# 3.01e-19
C4690 ctln[1] _204_/Y 3.74e-20
C4691 _336_/a_193_7# _313_/a_651_373# 9.52e-22
C4692 _336_/a_1108_7# _313_/a_543_7# 1.87e-20
C4693 _306_/a_218_7# _286_/B 1.25e-19
C4694 _188_/a_505_n19# _298_/B 0.0089f
C4695 _258_/S _311_/a_1283_n19# 3.53e-19
C4696 _215_/A _346_/SET_B 0.0126f
C4697 _216_/X _218_/a_346_7# 7.79e-20
C4698 _346_/a_193_7# _347_/Q 0.00306f
C4699 _346_/a_652_n19# _299_/X 0.00669f
C4700 _251_/a_79_n19# _284_/A 0.00501f
C4701 _343_/CLK _315_/a_761_249# 0.0191f
C4702 _334_/D _298_/A 9.79e-21
C4703 _238_/B _279_/A 1.65e-19
C4704 input3/a_27_7# _343_/CLK 0.0135f
C4705 _292_/A _311_/a_193_7# 6.48e-20
C4706 _277_/Y _346_/SET_B 0.0163f
C4707 _165_/a_215_7# VPWR -0.00196f
C4708 _165_/a_292_257# VGND -9.02e-19
C4709 _312_/Q _311_/a_1270_373# 1.91e-19
C4710 _327_/a_1283_n19# _279_/A 0.00151f
C4711 _344_/a_27_7# _162_/X 3.06e-19
C4712 _183_/a_27_7# _283_/A 0.00179f
C4713 _192_/B _204_/Y 0.0148f
C4714 clk _283_/A 0.00704f
C4715 _331_/Q _232_/X 0.568f
C4716 _168_/a_397_257# _346_/Q 4.01e-20
C4717 _304_/S _315_/a_27_7# 0.00161f
C4718 _320_/Q _246_/B 0.0255f
C4719 clkbuf_2_3_0_clk/A _199_/a_250_257# 0.00402f
C4720 _341_/a_651_373# VGND 7.52e-19
C4721 _175_/Y _226_/X 0.245f
C4722 _254_/A _336_/a_543_7# 1.33e-20
C4723 _336_/a_193_7# _157_/a_27_7# 1.52e-19
C4724 _341_/a_639_7# VPWR 4.88e-19
C4725 _342_/a_1217_7# _317_/D 7.57e-20
C4726 _338_/a_639_7# VPWR 4.72e-19
C4727 _338_/a_651_373# VGND 8.72e-19
C4728 _323_/a_27_7# _176_/a_27_7# 4.08e-20
C4729 _325_/a_193_7# _242_/A 2.28e-21
C4730 _331_/D _330_/a_193_7# 6.02e-19
C4731 _274_/a_39_257# _315_/D 8.8e-19
C4732 _168_/a_397_257# _168_/a_481_7# -1.71e-20
C4733 _167_/X _286_/Y 0.0611f
C4734 output9/a_27_7# _292_/A 6.73e-19
C4735 _316_/Q _316_/a_761_249# 0.0225f
C4736 _325_/a_761_249# _325_/Q 3.55e-20
C4737 clkbuf_2_1_0_clk/A _313_/a_27_7# 1.31e-21
C4738 _328_/a_543_7# _279_/A 0.00845f
C4739 _346_/SET_B _314_/a_639_7# -7.75e-19
C4740 _169_/Y clkbuf_2_3_0_clk/A 7.37e-19
C4741 _345_/Q _310_/D 3.57e-22
C4742 _318_/Q result[3] 0.00954f
C4743 _147_/A _298_/A 0.0389f
C4744 _343_/CLK _153_/A 5.93e-19
C4745 _235_/a_113_257# _316_/D 0.00656f
C4746 _324_/Q _247_/a_113_257# 0.0125f
C4747 _229_/a_76_159# VGND 0.00444f
C4748 _229_/a_489_373# VPWR 0.0386f
C4749 _346_/SET_B _304_/X 0.008f
C4750 _242_/A _317_/a_448_7# 0.00126f
C4751 _324_/a_1108_7# _248_/A 1.28e-21
C4752 clk _248_/B 2.95e-22
C4753 clkbuf_0_clk/X clkbuf_1_1_0_clk/a_75_172# 0.0106f
C4754 _337_/Q _310_/a_1283_n19# 0.00107f
C4755 _340_/a_1217_7# VPWR 1.38e-20
C4756 _340_/a_639_7# VGND 5.12e-19
C4757 _149_/A _298_/A 0.00729f
C4758 _340_/Q _284_/A 0.00784f
C4759 _236_/B _318_/D 0.00539f
C4760 _321_/D _242_/B 0.0641f
C4761 _342_/Q _146_/C 0.0172f
C4762 _316_/a_805_7# VPWR 2.26e-19
C4763 _316_/a_1270_373# VGND 4.72e-20
C4764 ctln[5] VGND 0.0805f
C4765 _327_/a_805_7# _330_/Q 3.13e-19
C4766 _345_/a_476_7# _346_/SET_B 0.0141f
C4767 _344_/a_1032_373# _164_/A 0.00446f
C4768 _169_/Y _172_/Y 0.00201f
C4769 _300_/a_301_257# _313_/a_761_249# 1.01e-20
C4770 _293_/a_39_257# _286_/B 0.00429f
C4771 _346_/a_193_7# _297_/B 0.0012f
C4772 _162_/X _171_/a_215_7# 0.00136f
C4773 _258_/S _309_/a_1270_373# 8.96e-21
C4774 _204_/a_27_7# VGND 0.00233f
C4775 _248_/A _324_/D 2.79e-20
C4776 _342_/Q _157_/A 0.00712f
C4777 _208_/a_215_7# VGND 0.0469f
C4778 cal _205_/a_79_n19# 0.00272f
C4779 _326_/Q _217_/X 0.161f
C4780 result[0] output23/a_27_7# 0.00264f
C4781 _309_/a_1108_7# _292_/A 0.00168f
C4782 _327_/a_651_373# VGND 0.00191f
C4783 _283_/A _280_/a_68_257# 0.00734f
C4784 _327_/a_639_7# VPWR 6.48e-19
C4785 _317_/a_1462_7# _232_/A 1.01e-19
C4786 _342_/a_1108_7# _342_/D 0.0406f
C4787 _346_/a_381_7# _346_/D 0.00318f
C4788 _273_/A _324_/a_1108_7# 1.11e-21
C4789 _236_/B _217_/A 2.54e-20
C4790 _331_/CLK _324_/D 3.1e-20
C4791 repeater43/X _315_/a_1270_373# -3.58e-20
C4792 _195_/a_373_7# _306_/S 1.83e-19
C4793 _195_/a_27_257# _340_/D 0.00316f
C4794 _326_/a_651_373# VGND 0.00703f
C4795 _215_/A _313_/a_761_249# 0.0184f
C4796 repeater43/X _227_/A 0.0332f
C4797 _312_/a_193_7# _312_/a_1283_n19# -6.53e-19
C4798 _320_/D ctlp[4] 4.32e-20
C4799 _281_/Y _306_/S 0.0347f
C4800 _345_/a_1032_373# _163_/a_215_7# 9.59e-20
C4801 _298_/B _304_/S 0.00428f
C4802 _273_/A _324_/D 0.00134f
C4803 _332_/a_193_7# _153_/B 0.0167f
C4804 _330_/Q _319_/a_27_7# 7.05e-20
C4805 _161_/Y trimb[4] 7.68e-19
C4806 _300_/Y _346_/SET_B 0.0173f
C4807 _324_/a_1108_7# _222_/a_93_n19# 2.81e-21
C4808 _332_/D VPWR 0.374f
C4809 _301_/X _248_/B 2.72e-21
C4810 _285_/A _312_/Q 4.06e-22
C4811 _328_/a_1270_373# VPWR 8.21e-20
C4812 _328_/a_448_7# VGND -0.00614f
C4813 _221_/a_93_n19# _328_/Q 0.033f
C4814 _326_/D _217_/A 1.22e-19
C4815 _166_/Y _306_/S 0.00552f
C4816 _248_/A _279_/A 0.0142f
C4817 _181_/X _214_/a_27_257# 0.0106f
C4818 _305_/a_76_159# _286_/B 0.0329f
C4819 _318_/Q _322_/Q 2.68e-19
C4820 _345_/a_1602_7# _273_/A 0.00971f
C4821 _271_/A _334_/a_761_249# 0.0203f
C4822 _271_/Y _334_/a_27_7# 1.78e-19
C4823 _269_/A sample 0.00292f
C4824 _192_/B _225_/B 0.00719f
C4825 _346_/SET_B _220_/a_93_n19# 0.00198f
C4826 _297_/B _173_/a_76_159# 0.0285f
C4827 output35/a_27_7# VPWR 0.0642f
C4828 _300_/a_301_257# _147_/A 0.00223f
C4829 _331_/CLK _279_/A 0.00943f
C4830 _337_/Q _336_/a_761_249# 0.00115f
C4831 _273_/A _309_/Q 0.0573f
C4832 _341_/Q _226_/X 0.0016f
C4833 _298_/B _225_/X 0.00986f
C4834 _307_/X _298_/B 0.0121f
C4835 _319_/a_193_7# _297_/B 0.00308f
C4836 _346_/a_1056_7# _299_/X 7.56e-19
C4837 _251_/X _284_/A 2.9e-19
C4838 _320_/Q result[5] 0.00783f
C4839 _334_/a_448_7# VGND -0.00614f
C4840 _334_/a_1270_373# VPWR -1.44e-19
C4841 _227_/A _334_/Q 5.32e-19
C4842 _292_/A _311_/a_1462_7# 4.85e-19
C4843 _321_/a_193_7# _280_/a_68_257# 8.83e-21
C4844 _218_/a_250_257# _331_/CLK 3.52e-19
C4845 _309_/a_193_7# _340_/CLK 0.00284f
C4846 _296_/a_213_83# _284_/A 0.00503f
C4847 _172_/A _182_/X 5.64e-20
C4848 _308_/X _196_/A 0.00703f
C4849 _320_/Q _320_/a_27_7# 2.67e-19
C4850 output16/a_27_7# ctlp[2] 0.0205f
C4851 _273_/A _279_/A 0.04f
C4852 _345_/a_27_7# _345_/D 0.139f
C4853 _345_/a_193_7# _345_/Q 6.38e-19
C4854 _215_/A _147_/A 0.0281f
C4855 _343_/a_761_249# _343_/CLK 4.24e-19
C4856 _324_/a_193_7# _304_/S 0.018f
C4857 _325_/a_761_249# _326_/Q 0.00471f
C4858 clkbuf_1_1_0_clk/a_75_172# _286_/Y 2.45e-20
C4859 _283_/Y _332_/a_27_7# 1.16e-20
C4860 _344_/Q _297_/Y 0.241f
C4861 _277_/Y _147_/A 0.289f
C4862 _346_/SET_B VGND 2.21f
C4863 en _192_/B 2.51e-20
C4864 _227_/A _191_/B 0.022f
C4865 _331_/Q _241_/a_113_257# 1.08e-20
C4866 trim[4] _309_/Q 0.00286f
C4867 _267_/A clkc 0.259f
C4868 _281_/Y _327_/D 0.00559f
C4869 _329_/a_1108_7# _281_/Y 0.0123f
C4870 _183_/a_1241_257# _298_/A 8.92e-19
C4871 _340_/a_27_7# _198_/a_93_n19# 6.21e-19
C4872 _273_/A _311_/a_193_7# 1.03e-20
C4873 _277_/A clkbuf_0_clk/X 0.0429f
C4874 _342_/a_761_249# _177_/A 4.32e-19
C4875 _342_/a_27_7# _298_/X 7.38e-22
C4876 _188_/a_76_159# VGND -0.00217f
C4877 _188_/a_218_334# VPWR -0.00162f
C4878 cal _225_/a_59_35# 0.0385f
C4879 _168_/a_109_7# _297_/Y 1.12e-19
C4880 _271_/A _333_/Q 5.62e-20
C4881 _346_/a_1140_373# VPWR 4.97e-20
C4882 _346_/a_562_373# VGND 8.84e-19
C4883 _271_/Y _207_/X 4.91e-20
C4884 _335_/a_193_7# _332_/Q 3.28e-19
C4885 _237_/a_199_7# _232_/X 3.34e-20
C4886 clkbuf_0_clk/a_110_7# _314_/a_193_7# 0.00166f
C4887 _309_/a_761_249# _346_/SET_B 0.00277f
C4888 _335_/a_761_249# _207_/X 0.00157f
C4889 _197_/a_27_7# _225_/a_59_35# 1.85e-20
C4890 _342_/a_543_7# _176_/a_27_7# 2.59e-20
C4891 _329_/a_448_7# _319_/Q 0.0162f
C4892 _343_/a_193_7# _147_/A 2.46e-20
C4893 _343_/a_1108_7# _226_/a_297_7# 3.09e-20
C4894 _306_/a_505_n19# _340_/CLK 5.65e-20
C4895 input1/X _175_/Y 0.0344f
C4896 _300_/Y _313_/a_761_249# 2.22e-20
C4897 _317_/a_27_7# _242_/B 1.17e-19
C4898 _265_/B _174_/a_27_257# 6.44e-19
C4899 _339_/Q _336_/a_761_249# 7.46e-20
C4900 _267_/B _262_/a_113_257# 1.04e-19
C4901 _346_/a_381_7# _314_/Q 1.97e-20
C4902 _328_/a_1283_n19# _328_/D 9.79e-21
C4903 _343_/a_193_7# _149_/A 9.34e-20
C4904 _329_/D _327_/D 2.04e-20
C4905 _323_/a_761_249# _334_/a_27_7# 1.68e-21
C4906 _200_/a_256_7# _311_/D 6.44e-21
C4907 _329_/a_1108_7# _329_/D 0.0482f
C4908 repeater43/X _321_/Q 0.459f
C4909 _283_/Y _338_/a_543_7# 3.55e-19
C4910 _236_/B _318_/a_448_7# 6.05e-20
C4911 _336_/a_543_7# _202_/a_250_257# 5.26e-20
C4912 _342_/Q _251_/a_79_n19# 0.00413f
C4913 _196_/A _254_/B 0.177f
C4914 _281_/Y _283_/A 0.123f
C4915 clkbuf_2_2_0_clk/a_75_172# VPWR 0.0882f
C4916 output33/a_27_7# _297_/Y 0.0114f
C4917 _290_/A output5/a_27_7# 7.41e-20
C4918 _143_/a_109_7# VGND 2.36e-19
C4919 _329_/Q output19/a_27_7# 6.23e-19
C4920 input4/X VPWR 4.35f
C4921 _299_/X _157_/a_27_7# 9.76e-19
C4922 _300_/Y _156_/a_39_257# 2.24e-19
C4923 repeater43/X _324_/a_639_7# -7.75e-19
C4924 _305_/a_439_7# _305_/X 2.68e-19
C4925 cal _336_/a_1283_n19# 2.69e-21
C4926 input1/X _336_/a_543_7# 0.0338f
C4927 _275_/A clkbuf_2_1_0_clk/a_75_172# 6.32e-19
C4928 _315_/D _327_/Q 0.0244f
C4929 _275_/Y _173_/a_76_159# 0.00351f
C4930 _222_/a_346_7# VGND -0.00177f
C4931 _162_/X _147_/Y 0.0202f
C4932 _324_/a_651_373# _327_/Q 1.47e-19
C4933 repeater43/X _297_/B -9.05e-20
C4934 _324_/a_1108_7# _217_/X 3.57e-21
C4935 _289_/a_121_257# _263_/B 8.96e-19
C4936 repeater43/X _318_/a_193_7# 0.0314f
C4937 _343_/a_1270_373# repeater43/X -7.59e-20
C4938 _336_/a_27_7# _260_/A 9.95e-20
C4939 _345_/Q VPWR 0.906f
C4940 _329_/a_193_7# _329_/a_543_7# -0.0231f
C4941 _291_/a_39_257# _339_/Q 0.0548f
C4942 _290_/A comp 9.17e-21
C4943 _254_/B _298_/X 0.00243f
C4944 _207_/C VPWR 0.366f
C4945 _206_/A VGND 1.06f
C4946 _239_/a_199_7# _242_/A 5.43e-19
C4947 _298_/A _150_/a_27_7# 0.0197f
C4948 _331_/a_193_7# _217_/A 5.87e-20
C4949 _244_/B valid 9.13e-19
C4950 _175_/Y _286_/Y 8.67e-19
C4951 _319_/a_1270_373# VGND 6.33e-20
C4952 _181_/X _330_/a_27_7# 9.79e-21
C4953 _313_/a_1283_n19# VPWR 0.0254f
C4954 _313_/a_761_249# VGND 0.00208f
C4955 _281_/Y _248_/B 0.00512f
C4956 _338_/Q _311_/a_448_7# 9.11e-22
C4957 _346_/SET_B _311_/a_639_7# 0.00103f
C4958 _328_/a_193_7# output19/a_27_7# 9.27e-20
C4959 _344_/a_1032_373# _292_/A 0.011f
C4960 _337_/a_1270_373# VPWR -1.13e-19
C4961 _337_/a_448_7# VGND -0.00223f
C4962 _300_/Y _147_/A 0.625f
C4963 _324_/D _217_/X 3.42e-21
C4964 _342_/a_543_7# _341_/a_543_7# 6.3e-19
C4965 _318_/Q _181_/X 0.0706f
C4966 _207_/a_27_7# _335_/Q 1.83e-19
C4967 _339_/Q _199_/a_346_7# 0.00244f
C4968 _169_/Y _157_/A 4.72e-21
C4969 _308_/S _295_/a_409_7# 1.57e-19
C4970 _314_/Q _313_/a_193_7# 2.47e-20
C4971 _157_/A _225_/B 0.0821f
C4972 _344_/a_1032_373# _160_/A 0.0144f
C4973 _340_/a_448_7# _305_/a_505_n19# 2.6e-20
C4974 _320_/Q _322_/a_1283_n19# 0.0351f
C4975 _334_/D VGND 0.0784f
C4976 _336_/a_193_7# _267_/A 6.42e-22
C4977 output7/a_27_7# VGND 0.091f
C4978 _279_/Y _305_/a_76_159# 0.00674f
C4979 clkbuf_2_0_0_clk/a_75_172# cal 2.04e-19
C4980 _257_/a_222_53# _306_/S 0.00168f
C4981 _277_/A _286_/Y 1.58e-19
C4982 _307_/a_218_7# VGND -5.84e-19
C4983 _323_/D valid 0.00228f
C4984 _306_/S _297_/Y 0.0102f
C4985 _156_/a_39_257# VGND 0.0172f
C4986 _317_/a_193_7# _245_/a_113_257# 7.71e-19
C4987 _254_/Y _281_/Y 1.28e-20
C4988 _165_/X _167_/a_109_7# 7.38e-20
C4989 _308_/S _332_/Q 0.0016f
C4990 input4/a_27_7# _340_/Q 4.84e-21
C4991 _324_/a_1462_7# _304_/S 0.00201f
C4992 _309_/a_1108_7# trim[4] 1.58e-19
C4993 _329_/D _248_/B 1.35e-19
C4994 _271_/A _226_/a_297_7# 3.07e-19
C4995 _191_/a_109_257# VGND -0.00128f
C4996 _217_/X _279_/A 0.295f
C4997 _319_/Q _321_/a_761_249# 2.15e-19
C4998 _296_/Y _324_/D 1.61e-20
C4999 _324_/Q _315_/a_543_7# 1.13e-19
C5000 _218_/a_93_n19# _331_/a_27_7# 2.75e-21
C5001 _340_/a_1283_n19# _197_/X 0.0279f
C5002 _188_/S _295_/a_79_n19# 6.6e-20
C5003 _341_/Q input1/X 0.00454f
C5004 _342_/D _177_/a_27_7# 1.04e-19
C5005 _218_/a_250_257# _217_/X 0.0215f
C5006 _325_/a_27_7# _315_/D 6.53e-21
C5007 _147_/A VGND 5.24f
C5008 _150_/C VPWR 1.08f
C5009 repeater42/a_27_7# _304_/S 8.43e-21
C5010 _325_/a_543_7# _324_/a_1283_n19# 0.0102f
C5011 _325_/a_27_7# _324_/a_651_373# 1.17e-19
C5012 _325_/a_761_249# _324_/a_1108_7# 0.00823f
C5013 _325_/a_448_7# _324_/a_193_7# 5.24e-21
C5014 _174_/a_27_257# _310_/Q 8.01e-21
C5015 ctln[7] _334_/a_27_7# 7.49e-21
C5016 _157_/A _314_/a_543_7# 3.09e-19
C5017 _255_/a_112_257# _255_/X 7.08e-20
C5018 _340_/Q _264_/a_113_257# 1.99e-20
C5019 _320_/a_193_7# _319_/a_193_7# 3.89e-21
C5020 _320_/a_761_249# _319_/a_27_7# 1.02e-21
C5021 _320_/a_27_7# _319_/a_761_249# 1.1e-21
C5022 _149_/A VGND 0.681f
C5023 _169_/Y _260_/A 0.0269f
C5024 clkbuf_0_clk/X _314_/a_448_7# 0.00261f
C5025 _260_/A _225_/B 0.565f
C5026 _217_/X _220_/a_346_7# 6.02e-19
C5027 _339_/a_1270_373# VPWR 7.38e-20
C5028 _339_/a_448_7# VGND -0.00607f
C5029 _324_/Q _224_/a_250_257# 0.0726f
C5030 _327_/a_1270_373# _232_/X 1.04e-19
C5031 _153_/B _190_/A 0.154f
C5032 _298_/B _150_/a_109_257# 9.65e-19
C5033 _258_/a_535_334# _340_/CLK 3.81e-21
C5034 _325_/a_1108_7# _304_/X 0.0421f
C5035 _325_/a_1283_n19# _217_/A 1.04e-19
C5036 _325_/a_761_249# _324_/D 1.29e-20
C5037 _317_/a_193_7# VPWR 0.06f
C5038 _294_/A _297_/Y 0.00699f
C5039 _281_/Y _225_/a_145_35# 6.26e-19
C5040 _343_/a_1108_7# _149_/a_27_7# 4.79e-21
C5041 _343_/a_1462_7# _149_/A 2.3e-19
C5042 _326_/a_1270_373# _232_/X 6.38e-20
C5043 _172_/A _340_/CLK 3.6e-19
C5044 output38/a_27_7# VGND 0.0661f
C5045 input4/X _335_/a_1108_7# 2.15e-19
C5046 repeater43/X _335_/a_543_7# 2.08e-19
C5047 _336_/a_761_249# _336_/D 1.25e-20
C5048 _336_/a_1283_n19# _284_/A 0.00794f
C5049 _330_/Q _331_/a_1108_7# 0.0121f
C5050 _342_/Q _251_/X 1.18e-19
C5051 _271_/A _212_/X 2.23e-20
C5052 _318_/a_543_7# _317_/a_193_7# 2.21e-21
C5053 _318_/a_193_7# _317_/a_543_7# 1.26e-19
C5054 _211_/a_27_257# _332_/D 0.00193f
C5055 _211_/a_109_257# _340_/CLK 0.00175f
C5056 _342_/Q _296_/a_213_83# 0.00547f
C5057 _306_/S _335_/Q 5.92e-21
C5058 _312_/a_448_7# _312_/Q 6.16e-21
C5059 _188_/S _180_/a_29_13# 0.00938f
C5060 _309_/a_193_7# _267_/B 4.69e-19
C5061 _331_/a_1283_n19# VPWR 0.0444f
C5062 _331_/a_761_249# VGND 0.0314f
C5063 _340_/a_27_7# _147_/Y 3.72e-21
C5064 _328_/a_651_373# _232_/X 0.00109f
C5065 _232_/X _347_/D 1.02e-19
C5066 _320_/a_1108_7# _346_/SET_B -0.00685f
C5067 _341_/Q _286_/Y 0.307f
C5068 _294_/A _310_/a_193_7# 7.75e-21
C5069 _302_/a_77_159# VPWR 0.0136f
C5070 _335_/a_1108_7# _207_/C 9.43e-19
C5071 _214_/a_27_257# _346_/SET_B 1.39e-19
C5072 repeater43/X _318_/a_1462_7# 0.0014f
C5073 _344_/a_652_n19# _346_/SET_B 0.0107f
C5074 _316_/a_651_373# _317_/D 0.00435f
C5075 _290_/A _310_/a_1270_373# 1.79e-19
C5076 _308_/a_76_159# _192_/B 0.0427f
C5077 _336_/a_193_7# _194_/X 0.00112f
C5078 _336_/a_27_7# _340_/Q 7.47e-21
C5079 _254_/B _204_/a_27_257# 1.37e-19
C5080 _302_/a_323_257# _297_/B 1.56e-19
C5081 _260_/A _314_/a_543_7# 1.96e-19
C5082 _304_/a_79_n19# _162_/X 6.06e-19
C5083 _283_/Y _333_/Q 1.76e-19
C5084 _323_/D _229_/a_226_7# 3.19e-20
C5085 _338_/Q _311_/D 0.00682f
C5086 _258_/a_218_7# _346_/SET_B 7.09e-19
C5087 _335_/a_651_373# _334_/D 1.02e-19
C5088 ctln[7] _207_/X 4.5e-19
C5089 _335_/a_1270_373# _343_/CLK 1.39e-19
C5090 _335_/a_543_7# _334_/Q 0.00156f
C5091 _337_/D VGND 0.143f
C5092 _315_/a_543_7# _228_/A 0.0013f
C5093 _342_/D _341_/a_27_7# 2.29e-20
C5094 _197_/X _190_/a_27_7# 0.0144f
C5095 _322_/a_193_7# _331_/CLK 0.00344f
C5096 ctln[1] _335_/a_193_7# 0.00123f
C5097 _298_/C _147_/Y 3.61e-21
C5098 _181_/a_27_7# _190_/A 8.85e-22
C5099 _321_/Q result[6] 0.117f
C5100 _277_/A _240_/B 1.57e-19
C5101 _344_/a_1182_221# _163_/a_215_7# 2.94e-19
C5102 _314_/a_27_7# _228_/A 1.85e-20
C5103 _310_/D _284_/A 0.00878f
C5104 ctlp[7] _322_/Q 2.39e-19
C5105 _251_/a_79_n19# _225_/B 4.21e-21
C5106 _271_/Y _323_/Q 1.61e-20
C5107 _275_/A _285_/Y 6.87e-20
C5108 _340_/CLK _203_/a_80_n19# 3.64e-21
C5109 _346_/SET_B _198_/a_256_7# 0.00221f
C5110 _250_/a_78_159# _215_/A 0.0222f
C5111 _317_/a_1283_n19# _246_/B 2.15e-19
C5112 _187_/a_27_7# _146_/C 0.00121f
C5113 _320_/Q _330_/a_448_7# 0.0161f
C5114 _342_/a_761_249# _248_/A 0.0103f
C5115 _327_/a_448_7# _331_/D 7.67e-20
C5116 _146_/C _315_/D 0.238f
C5117 _344_/a_1032_373# _273_/A 7.5e-20
C5118 _252_/a_109_257# _216_/X 4.19e-19
C5119 output12/a_27_7# _154_/A 9.24e-21
C5120 clkbuf_2_1_0_clk/A _281_/A 0.0147f
C5121 result[6] _318_/a_193_7# 3.82e-20
C5122 input4/X _323_/a_1108_7# 3.51e-20
C5123 repeater43/X _323_/a_543_7# 0.00516f
C5124 clkbuf_0_clk/X _330_/Q 0.0593f
C5125 _242_/A _327_/D 0.00461f
C5126 _342_/Q _232_/A 0.00387f
C5127 _184_/a_505_n19# _150_/C 0.0592f
C5128 _184_/a_76_159# _226_/X 0.00258f
C5129 _184_/a_535_334# _147_/A 7.89e-20
C5130 _157_/A _315_/D 1.06e-19
C5131 _301_/a_512_257# _297_/Y 0.00217f
C5132 _271_/A _149_/a_27_7# 8.86e-21
C5133 _183_/a_471_7# VPWR -0.00198f
C5134 _183_/a_1241_257# VGND -1.84e-20
C5135 _144_/a_27_7# _232_/A 1.1e-19
C5136 _250_/X _298_/A 1.05e-19
C5137 _316_/Q _317_/a_1283_n19# 1.85e-20
C5138 _330_/D _212_/X 5.15e-20
C5139 _324_/a_1283_n19# _324_/Q 0.0155f
C5140 clk ctln[0] 0.00419f
C5141 _303_/A _347_/Q 2.54e-20
C5142 _325_/a_651_373# VPWR 2.05e-19
C5143 _301_/X _160_/X 0.232f
C5144 _325_/a_1108_7# VGND 0.0165f
C5145 _333_/a_1108_7# _298_/C 2.43e-20
C5146 _277_/A _328_/Q 0.21f
C5147 output13/a_27_7# _334_/D 9.34e-20
C5148 _308_/X _143_/a_27_7# 1.1e-21
C5149 _271_/A _317_/a_448_7# 6.75e-20
C5150 _197_/X _332_/Q 0.0111f
C5151 _344_/a_27_7# _345_/Q 7.63e-19
C5152 clkbuf_0_clk/X _314_/D 0.155f
C5153 _341_/D _317_/D 0.00783f
C5154 _257_/a_222_53# _254_/Y 0.00404f
C5155 _339_/D VGND 0.337f
C5156 _168_/a_397_257# clkbuf_2_1_0_clk/A 0.00281f
C5157 _216_/A _224_/a_250_257# 0.00795f
C5158 _306_/S _209_/a_373_7# 0.002f
C5159 _306_/S _336_/Q 0.228f
C5160 _333_/a_651_373# _332_/a_1283_n19# 2e-20
C5161 _333_/a_1283_n19# _332_/a_651_373# 2.06e-20
C5162 _275_/Y _172_/a_109_257# 7.92e-19
C5163 _269_/A _175_/Y 7.15e-20
C5164 _317_/a_1462_7# VPWR 3.75e-19
C5165 _317_/a_805_7# VGND -6.39e-19
C5166 _242_/A _283_/A 0.00818f
C5167 _286_/B _181_/X 0.137f
C5168 _202_/a_93_n19# VPWR 0.0163f
C5169 _297_/A _347_/a_448_7# 0.025f
C5170 _283_/A _335_/Q 5.16e-19
C5171 _299_/X _267_/A 5.38e-20
C5172 output36/a_27_7# comp 0.0114f
C5173 input4/a_27_7# rstn 0.0524f
C5174 ctln[4] _195_/a_27_257# 1.14e-19
C5175 _341_/a_193_7# _177_/a_27_7# 1.21e-19
C5176 _258_/S trim[1] 0.0138f
C5177 _232_/X _222_/a_584_7# 2.11e-19
C5178 _314_/a_651_373# _284_/A 4.88e-21
C5179 _312_/D _312_/Q 8.91e-20
C5180 cal VPWR 5.29f
C5181 _276_/a_150_257# VGND -2.14e-19
C5182 _216_/A clkbuf_2_1_0_clk/A 0.00766f
C5183 _205_/a_79_n19# _204_/Y 0.00322f
C5184 _238_/B ctlp[4] 1.21e-19
C5185 _317_/Q _325_/Q 0.668f
C5186 _304_/a_288_7# _286_/B 2.41e-19
C5187 _260_/A _315_/D 0.00202f
C5188 _343_/D _175_/Y 0.00245f
C5189 _169_/Y _165_/X 9.39e-19
C5190 _323_/a_761_249# _323_/Q 0.00262f
C5191 _197_/a_27_7# VPWR 0.093f
C5192 _256_/a_209_7# _181_/X 1.17e-19
C5193 _197_/X _337_/a_193_7# 0.00445f
C5194 _236_/B _317_/D 1.07e-19
C5195 _343_/a_805_7# cal 2.74e-19
C5196 _258_/a_505_n19# _254_/A 1.5e-19
C5197 _254_/A _311_/D 7.15e-19
C5198 _280_/a_150_257# VPWR -5.5e-19
C5199 _308_/S _192_/B 0.00346f
C5200 clkbuf_0_clk/X clkbuf_2_1_0_clk/a_75_172# 1.36e-21
C5201 _342_/a_27_7# _343_/CLK 0.0239f
C5202 _275_/Y _337_/Q 0.0277f
C5203 _283_/Y _339_/a_761_249# 8.47e-21
C5204 _242_/A _248_/B 1.98e-19
C5205 _318_/Q _346_/SET_B 0.185f
C5206 _303_/A _297_/B 2.37e-19
C5207 _172_/A _307_/a_439_7# 9.5e-20
C5208 _277_/Y _319_/Q 0.00188f
C5209 _326_/a_1283_n19# _331_/Q 1.12e-19
C5210 _294_/Y _265_/B 0.0107f
C5211 _150_/a_193_257# VPWR -1.54e-19
C5212 _281_/Y _324_/a_193_7# 0.00945f
C5213 _174_/a_109_7# VGND 1.65e-19
C5214 _150_/a_27_7# VGND 0.0919f
C5215 _285_/A _267_/B 4.96e-20
C5216 _172_/A _304_/S 6.94e-20
C5217 _266_/a_113_257# _284_/A 0.0196f
C5218 _286_/B _343_/Q 3.13e-21
C5219 _165_/a_78_159# _164_/Y 0.0159f
C5220 _260_/B _162_/X 6.44e-20
C5221 _248_/A _330_/a_543_7# 1e-20
C5222 _330_/Q _286_/Y 6.4e-21
C5223 _324_/a_1283_n19# _228_/A 7.74e-20
C5224 _219_/a_584_7# _330_/Q 3.49e-19
C5225 _321_/a_193_7# _242_/A 9.19e-19
C5226 _258_/a_218_7# _147_/A 5.34e-19
C5227 output23/a_27_7# _324_/Q 1.29e-19
C5228 _251_/X _225_/B 1.95e-20
C5229 _331_/CLK _330_/a_543_7# 0.00432f
C5230 _250_/X _215_/A 0.00589f
C5231 _172_/A _225_/X 1.27e-20
C5232 _196_/A _347_/a_1283_n19# 2.86e-21
C5233 _324_/a_805_7# _286_/Y 3.41e-19
C5234 _290_/A _215_/A 2.62e-20
C5235 _307_/X _172_/A 4.39e-19
C5236 _340_/CLK _312_/a_448_7# 0.00193f
C5237 _219_/a_346_7# VPWR -2.03e-19
C5238 _219_/a_250_257# VGND -0.00542f
C5239 repeater43/X _322_/a_1108_7# 0.00433f
C5240 rstn _204_/Y 9.06e-20
C5241 _309_/D _311_/D 0.00628f
C5242 _255_/B _298_/A 0.376f
C5243 _339_/Q _311_/a_1108_7# 4.13e-19
C5244 _314_/D _286_/Y 1.2e-21
C5245 _319_/Q _304_/X 2.04e-19
C5246 _346_/Q _346_/D 0.00673f
C5247 _313_/a_193_7# _254_/B 2.15e-20
C5248 _335_/D _225_/X 4.53e-21
C5249 _333_/a_193_7# _332_/Q 0.00197f
C5250 _333_/a_27_7# _333_/Q 0.0159f
C5251 _188_/S _226_/X 9.24e-19
C5252 _345_/a_652_n19# _166_/Y 2.97e-20
C5253 _341_/a_27_7# _341_/a_193_7# -0.292f
C5254 _305_/X _194_/A 0.0731f
C5255 _176_/a_27_7# _298_/C 0.00208f
C5256 _167_/X _170_/a_556_7# 4.45e-19
C5257 _308_/a_535_334# input1/X 0.00104f
C5258 _250_/a_493_257# VPWR -2.68e-20
C5259 _250_/a_78_159# VGND -0.00729f
C5260 _324_/a_1283_n19# _216_/A 2.43e-20
C5261 repeater43/X output25/a_27_7# 6.86e-19
C5262 _343_/CLK _254_/B 2.57e-20
C5263 _197_/X _339_/a_193_7# 7.06e-20
C5264 _321_/a_543_7# _234_/B 2.61e-19
C5265 _321_/a_193_7# _322_/D 1.27e-20
C5266 _306_/a_76_159# cal 5.67e-20
C5267 _251_/a_79_n19# _315_/D 5.03e-21
C5268 _343_/CLK _317_/D 0.0127f
C5269 _315_/D _221_/a_250_257# 7.71e-19
C5270 _321_/a_193_7# _321_/a_448_7# -0.00297f
C5271 _275_/Y _339_/Q 0.00742f
C5272 _218_/a_93_n19# _281_/A 1.57e-19
C5273 _338_/a_27_7# _338_/a_193_7# -0.298f
C5274 _275_/A output18/a_27_7# 1.51e-19
C5275 result[4] _318_/a_193_7# 0.00134f
C5276 _268_/a_39_257# _316_/a_543_7# 3.28e-19
C5277 _283_/A _336_/Q 2.74e-20
C5278 _304_/S _244_/B 0.00807f
C5279 _342_/a_448_7# repeater43/X 1.84e-21
C5280 _158_/Y _172_/B 9.72e-20
C5281 clkbuf_2_3_0_clk/A _197_/X 5.15e-20
C5282 _323_/Q _154_/a_27_7# 4.78e-20
C5283 _338_/Q _312_/a_1283_n19# 4.29e-20
C5284 _296_/Y _181_/a_27_7# 3.33e-20
C5285 _331_/Q _248_/A 0.0124f
C5286 _166_/Y _160_/X 0.0225f
C5287 _284_/A VPWR 1.59f
C5288 _322_/a_27_7# output28/a_27_7# 0.00236f
C5289 _297_/A _347_/D 0.0231f
C5290 ctln[7] _323_/Q 1.18e-19
C5291 _332_/a_193_7# _332_/a_1108_7# -0.00656f
C5292 output32/a_27_7# _346_/SET_B 1.79e-19
C5293 _317_/Q _326_/Q 0.0332f
C5294 _313_/Q _313_/a_1108_7# 1.35e-19
C5295 _306_/X _313_/a_1283_n19# 6.09e-20
C5296 _184_/a_505_n19# cal 0.00141f
C5297 _184_/a_76_159# input1/X 0.0505f
C5298 ctlp[7] ctlp[1] 2.69e-20
C5299 _345_/a_476_7# _290_/A 6.29e-19
C5300 _340_/a_543_7# _338_/a_27_7# 3.06e-21
C5301 _232_/X _331_/a_543_7# 0.00221f
C5302 _319_/Q _300_/Y 7.96e-22
C5303 _258_/a_76_159# _337_/Q 1.89e-19
C5304 _347_/a_193_7# _347_/a_651_373# -0.00701f
C5305 _292_/A _312_/Q 0.0505f
C5306 _169_/B _301_/a_149_7# 2.75e-21
C5307 _322_/Q _316_/D 0.0011f
C5308 _331_/Q _331_/CLK 0.324f
C5309 _167_/X _299_/X 1.13f
C5310 _267_/A _311_/a_1283_n19# 1.63e-19
C5311 _319_/Q _220_/a_93_n19# 3.54e-20
C5312 _294_/Y _310_/Q 7.25e-20
C5313 clkbuf_0_clk/a_110_7# _181_/a_27_7# 2.65e-19
C5314 _273_/A _331_/Q 7.26e-22
C5315 _313_/Q _254_/A 0.436f
C5316 _195_/a_109_7# VGND 6.85e-20
C5317 _309_/a_27_7# _284_/A 0.623f
C5318 _340_/a_193_7# _340_/a_1283_n19# -6.53e-19
C5319 _291_/a_39_257# _310_/a_1283_n19# 2.31e-20
C5320 _277_/Y _167_/a_27_257# 0.00488f
C5321 _346_/a_1182_221# _162_/X 1.82e-19
C5322 _325_/Q _298_/A 3.08e-20
C5323 _177_/A _229_/a_226_7# 4.1e-21
C5324 _317_/a_27_7# _244_/B 2.73e-19
C5325 _323_/a_448_7# clk 3.36e-19
C5326 _163_/a_292_257# _162_/X 4.11e-19
C5327 _254_/Y _336_/Q 0.0193f
C5328 _308_/S _157_/A 3.28e-20
C5329 _298_/a_27_7# _298_/A 0.00896f
C5330 _316_/a_27_7# _316_/a_543_7# -0.00505f
C5331 _310_/a_761_249# _310_/D 0.0432f
C5332 _326_/a_1108_7# _181_/X 2.04e-19
C5333 clkbuf_2_3_0_clk/A _312_/a_193_7# 3.78e-20
C5334 _331_/Q _222_/a_93_n19# 3.8e-20
C5335 _209_/a_109_257# _153_/a_109_53# 1.37e-21
C5336 _308_/X _146_/a_184_13# 9.35e-20
C5337 _255_/B _215_/A 0.00868f
C5338 _232_/A _315_/a_448_7# 7.67e-20
C5339 _186_/a_382_257# _146_/C 2.59e-20
C5340 _209_/X _209_/a_27_257# 0.00134f
C5341 _336_/a_193_7# _336_/a_543_7# -0.0231f
C5342 _336_/a_27_7# _336_/a_1283_n19# -9.15e-20
C5343 _319_/Q VGND 1.25f
C5344 _281_/Y repeater42/a_27_7# 0.0043f
C5345 _172_/A _183_/a_27_7# 0.00604f
C5346 _343_/a_27_7# _185_/A 0.0121f
C5347 _282_/a_39_257# _330_/a_1108_7# 6.24e-21
C5348 _345_/Q _147_/Y 0.202f
C5349 _248_/B _314_/a_761_249# 1.24e-19
C5350 _172_/A clk 0.0867f
C5351 _327_/a_1108_7# _237_/a_113_257# 1.36e-19
C5352 _327_/a_27_7# _320_/Q 3.52e-21
C5353 _340_/CLK _312_/D 0.09f
C5354 _194_/a_27_7# _310_/a_193_7# 1.99e-20
C5355 _313_/Q _309_/D 1.18e-20
C5356 _154_/A _205_/a_297_7# 4.41e-20
C5357 _327_/a_27_7# _327_/a_193_7# -0.138f
C5358 _322_/a_1283_n19# result[7] 0.00279f
C5359 _313_/a_1283_n19# _147_/Y 0.00181f
C5360 _290_/A trimb[1] 3e-20
C5361 _301_/a_149_7# _170_/a_226_7# 4.38e-19
C5362 _333_/a_1462_7# _332_/Q 1.83e-19
C5363 _323_/a_1108_7# cal 0.00654f
C5364 _306_/a_76_159# _284_/A 0.045f
C5365 clk _335_/D 0.00972f
C5366 _215_/A _310_/a_27_7# 3.59e-21
C5367 _200_/a_250_257# _340_/a_1108_7# 3.1e-20
C5368 _292_/Y trimb[3] 0.0115f
C5369 _256_/a_209_257# _340_/CLK 7.23e-20
C5370 _330_/Q _328_/Q 0.00253f
C5371 _329_/a_193_7# _330_/Q 0.00872f
C5372 _345_/a_193_7# _167_/a_109_7# 9.7e-20
C5373 _331_/D _331_/a_193_7# 0.00428f
C5374 _262_/a_113_257# _297_/Y 0.0037f
C5375 _250_/X VGND 0.0823f
C5376 _331_/a_193_7# _330_/a_193_7# 1.5e-20
C5377 _225_/a_59_35# _225_/B 0.0283f
C5378 trim[2] VPWR 0.263f
C5379 _290_/A VGND 1.02f
C5380 _332_/a_1108_7# _208_/a_78_159# 8.41e-20
C5381 _211_/a_109_7# _339_/D 5.75e-20
C5382 _277_/A clkbuf_2_3_0_clk/a_75_172# 8.92e-20
C5383 repeater42/a_27_7# _329_/D 1.09e-21
C5384 _326_/a_27_7# _326_/a_193_7# -0.327f
C5385 _251_/X _315_/D 0.0088f
C5386 _273_/A _299_/a_292_257# 0.00376f
C5387 _255_/B _304_/X 3.95e-20
C5388 _339_/D _198_/a_256_7# 5.39e-19
C5389 clkbuf_2_1_0_clk/A _301_/a_240_7# 0.00171f
C5390 _308_/S _260_/A 2.31e-21
C5391 repeater43/X _333_/a_543_7# 3.32e-19
C5392 _329_/a_27_7# VPWR 0.0411f
C5393 input1/X _311_/D 2.45e-19
C5394 _258_/a_505_n19# input1/X 1.07e-20
C5395 _315_/D _296_/a_213_83# 0.0676f
C5396 _198_/a_93_n19# _202_/a_93_n19# 1.68e-19
C5397 _340_/a_193_7# _190_/a_27_7# 1.42e-19
C5398 _286_/B _346_/SET_B 0.154f
C5399 _329_/a_761_249# _297_/B 3.58e-20
C5400 _342_/D repeater43/X 0.414f
C5401 _319_/Q output27/a_27_7# 5.45e-20
C5402 _182_/a_79_n19# _178_/a_27_7# 1.11e-20
C5403 _281_/A _328_/D 3.4e-20
C5404 _172_/A _301_/X 2.16e-20
C5405 _193_/Y _311_/a_193_7# 6.47e-21
C5406 _322_/a_1108_7# result[6] 0.0055f
C5407 _333_/a_651_373# _206_/A 8.49e-19
C5408 _332_/a_193_7# _340_/CLK 2.92e-19
C5409 _332_/a_27_7# _332_/D 0.0552f
C5410 cal _198_/a_93_n19# 0.0101f
C5411 _301_/a_51_257# _299_/X 0.0423f
C5412 _290_/A _309_/a_761_249# 0.00181f
C5413 _188_/S input1/X 0.365f
C5414 _167_/a_109_257# _160_/X 5.32e-19
C5415 _345_/a_1224_7# _290_/A 3.74e-20
C5416 _182_/X _248_/A 2.34e-20
C5417 _153_/a_215_257# _153_/A 0.0148f
C5418 clk _203_/a_80_n19# 0.00122f
C5419 _347_/a_761_249# _347_/D 0.00117f
C5420 _334_/a_1283_n19# _343_/Q 1.42e-19
C5421 _209_/X _153_/A 0.261f
C5422 _336_/a_1108_7# _336_/Q 7.63e-20
C5423 output14/a_27_7# _331_/CLK 2.03e-21
C5424 _269_/A _269_/Y 0.0862f
C5425 _326_/Q _298_/A 4.92e-21
C5426 output26/a_27_7# _322_/a_27_7# 1.99e-19
C5427 _242_/A _242_/B 0.373f
C5428 _158_/Y trimb[4] 2.84e-19
C5429 _160_/X _297_/Y 0.00998f
C5430 output12/a_27_7# _153_/B 2.42e-19
C5431 _346_/a_1296_7# _162_/X 1.92e-19
C5432 _323_/D clk 6.86e-19
C5433 clkbuf_2_1_0_clk/a_75_172# _328_/Q 1.85e-19
C5434 _297_/A _304_/S 4.81e-20
C5435 _342_/a_27_7# output30/a_27_7# 1.86e-19
C5436 _248_/A valid 2.19e-19
C5437 _333_/a_193_7# _192_/B 5.71e-19
C5438 _333_/a_543_7# _191_/B 0.0308f
C5439 _233_/a_113_257# _331_/a_1108_7# 5.81e-20
C5440 _273_/A _312_/Q 3.06e-20
C5441 _279_/Y ctln[5] 0.257f
C5442 _187_/a_27_7# _232_/A 0.00139f
C5443 _310_/a_639_7# _310_/Q 1.76e-19
C5444 _329_/a_651_373# _218_/a_93_n19# 2.1e-19
C5445 _343_/D _269_/Y 0.00183f
C5446 _331_/Q _217_/X 0.0213f
C5447 _209_/a_109_257# _153_/A 0.0037f
C5448 _294_/Y _311_/a_27_7# 3.45e-21
C5449 _232_/A _315_/D 0.281f
C5450 _338_/a_1283_n19# _340_/CLK 0.0375f
C5451 _167_/a_109_7# VPWR -8.08e-19
C5452 _167_/a_27_257# VGND -0.00535f
C5453 _188_/S _286_/Y 0.0819f
C5454 _342_/a_1283_n19# _146_/C 1.63e-20
C5455 _247_/a_199_7# VGND -3.13e-19
C5456 _313_/D _157_/A 8.5e-19
C5457 _346_/SET_B _347_/a_543_7# -9.49e-19
C5458 _219_/a_256_7# _232_/X 5.29e-19
C5459 _181_/X _222_/a_250_257# 0.00777f
C5460 _309_/a_448_7# _306_/S 2.93e-20
C5461 _347_/Q _319_/D 0.00388f
C5462 _325_/Q _304_/X 0.61f
C5463 _207_/a_109_7# _153_/B 1.41e-19
C5464 _322_/D _242_/B 1.61e-20
C5465 _292_/A _340_/CLK 1.31e-20
C5466 _338_/a_27_7# _337_/a_27_7# 8.92e-20
C5467 _189_/a_27_7# VGND 0.121f
C5468 _286_/B _206_/A 0.00769f
C5469 _286_/B _313_/a_761_249# 0.00312f
C5470 _196_/A _313_/a_193_7# 5.13e-20
C5471 _298_/C _333_/Q 2.49e-19
C5472 _255_/B VGND 0.567f
C5473 _342_/Q VPWR 2.2f
C5474 _340_/a_448_7# _340_/CLK 0.0115f
C5475 _257_/a_544_257# VPWR -7.83e-19
C5476 _257_/a_79_159# VGND 0.0165f
C5477 _292_/Y VPWR 0.252f
C5478 _144_/a_27_7# VPWR 0.0765f
C5479 _341_/a_448_7# _341_/D 0.0275f
C5480 _329_/a_1462_7# _330_/Q 3.27e-19
C5481 _154_/A _298_/A 2.44e-19
C5482 _258_/a_76_159# _336_/D 1.45e-20
C5483 _313_/Q _202_/a_250_257# 7.39e-21
C5484 _306_/X _202_/a_93_n19# 1.11e-20
C5485 input4/a_27_7# VPWR 0.0865f
C5486 _224_/a_93_n19# _224_/a_250_257# -6.97e-22
C5487 _332_/a_1108_7# _190_/A 2.15e-19
C5488 _340_/a_193_7# _337_/a_193_7# 0.0045f
C5489 _194_/a_27_7# _336_/Q 4.05e-19
C5490 _164_/A _267_/B 3.26e-20
C5491 _305_/a_535_334# _260_/A 3.1e-19
C5492 _328_/a_639_7# _329_/Q 0.00466f
C5493 _329_/a_639_7# VGND -0.00152f
C5494 _329_/a_1217_7# VPWR 2.02e-19
C5495 clkbuf_2_3_0_clk/A _299_/a_215_7# 0.00329f
C5496 _338_/a_1108_7# _346_/SET_B -0.00919f
C5497 _338_/a_448_7# _338_/D 0.0145f
C5498 _338_/a_761_249# _338_/Q 4.87e-20
C5499 _306_/X cal 1.43e-22
C5500 _313_/Q input1/X 0.0865f
C5501 _169_/B _215_/A 1.4e-19
C5502 _329_/Q _319_/a_27_7# 0.00378f
C5503 _320_/Q _319_/a_193_7# 5.13e-20
C5504 _244_/a_109_257# sample 0.00156f
C5505 _310_/a_27_7# VGND 0.0361f
C5506 _310_/a_761_249# VPWR 0.025f
C5507 _198_/a_93_n19# _284_/A 8.06e-19
C5508 _272_/a_39_257# _325_/Q 3.3e-19
C5509 _277_/Y _169_/B 9.29e-20
C5510 input4/X _332_/a_27_7# 1.52e-20
C5511 _283_/Y _207_/a_27_7# 1.1e-19
C5512 _188_/a_76_159# _341_/a_1108_7# 3.31e-20
C5513 _344_/a_1602_7# _344_/Q 0.0271f
C5514 _344_/a_476_7# _344_/D 0.00312f
C5515 _313_/D _260_/A 1e-19
C5516 _342_/a_1270_373# cal 2.6e-20
C5517 _182_/a_215_7# _192_/B 4.55e-19
C5518 _309_/a_193_7# _297_/Y 2.12e-20
C5519 result[1] _269_/A 0.00627f
C5520 _294_/A _309_/a_448_7# 0.0248f
C5521 _277_/A _299_/X 0.00183f
C5522 _334_/a_1108_7# _204_/a_27_257# 1.61e-19
C5523 _343_/CLK _298_/X 0.0162f
C5524 _297_/B _319_/D 0.00303f
C5525 _304_/a_257_159# _304_/S 0.04f
C5526 _264_/a_113_257# VPWR 0.0395f
C5527 _340_/a_651_373# _346_/SET_B 0.00164f
C5528 _286_/B _147_/A 0.041f
C5529 _273_/A _165_/a_493_257# 2.5e-19
C5530 _281_/Y _172_/A 0.0108f
C5531 _197_/X _260_/A 0.088f
C5532 _304_/S _177_/A 0.0107f
C5533 _275_/A _216_/X 7.98e-21
C5534 _279_/Y _346_/SET_B 0.0124f
C5535 _332_/a_761_249# _206_/A 4.16e-21
C5536 _332_/a_27_7# _207_/C 5.4e-19
C5537 _339_/a_27_7# _338_/a_27_7# 3.23e-19
C5538 _271_/A _205_/a_382_257# 1.81e-19
C5539 _309_/a_761_249# _310_/a_27_7# 4.89e-21
C5540 _229_/a_226_7# _248_/A 0.034f
C5541 _307_/a_76_159# _298_/C 2.26e-19
C5542 _281_/Y _211_/a_109_257# 6.56e-20
C5543 _172_/A _166_/Y 1.16e-19
C5544 _281_/Y _232_/X 0.029f
C5545 _275_/A _329_/Q 2.45e-19
C5546 _304_/a_79_n19# _150_/C 0.00251f
C5547 _327_/a_1108_7# _346_/SET_B 0.0183f
C5548 _324_/a_761_249# _326_/Q 0.00115f
C5549 _346_/a_193_7# _346_/a_652_n19# -0.00373f
C5550 _346_/a_27_7# _346_/a_476_7# -0.00544f
C5551 repeater43/X _341_/a_193_7# 0.00118f
C5552 _343_/CLK _332_/a_543_7# 1.9e-20
C5553 _339_/Q _312_/a_543_7# 5.39e-20
C5554 _309_/a_27_7# _264_/a_113_257# 2.65e-19
C5555 _204_/Y VPWR 0.0967f
C5556 _215_/A _314_/a_193_7# 1.16e-19
C5557 _307_/X _177_/A 4.48e-20
C5558 _197_/X _261_/A 5.25e-21
C5559 _147_/Y _202_/a_93_n19# 1.72e-19
C5560 _271_/A _248_/B 0.00876f
C5561 _340_/a_761_249# _339_/a_27_7# 1.73e-21
C5562 _340_/a_193_7# _339_/a_193_7# 3.19e-19
C5563 _343_/a_651_373# _175_/Y 3.06e-20
C5564 _325_/Q VGND 2.79f
C5565 _342_/a_1108_7# sample 4.84e-19
C5566 _181_/X _144_/A 8.16e-19
C5567 trim[3] _273_/Y 0.013f
C5568 _242_/A _318_/a_1283_n19# 0.00527f
C5569 _254_/A _347_/a_27_7# 1.12e-21
C5570 _320_/a_761_249# _328_/Q 3.19e-21
C5571 _326_/Q _304_/X 0.156f
C5572 _344_/a_652_n19# _290_/A 1.05e-19
C5573 output36/a_27_7# trimb[1] 4.29e-20
C5574 trimb[0] output37/a_27_7# 2.76e-20
C5575 _298_/a_181_7# VPWR -6.03e-20
C5576 _298_/a_27_7# VGND 0.0495f
C5577 _308_/a_505_n19# _210_/a_27_7# 8.53e-21
C5578 cal _147_/Y 4.32e-20
C5579 _298_/C _226_/a_297_7# 1.34e-20
C5580 _181_/X _331_/a_27_7# 0.00729f
C5581 _336_/a_27_7# VPWR 0.0258f
C5582 _328_/a_1283_n19# _346_/SET_B 0.0429f
C5583 repeater42/a_27_7# _242_/A 0.0596f
C5584 _304_/S _325_/D 2.46e-19
C5585 _329_/D _232_/X 0.00438f
C5586 _267_/A _172_/B 2.04e-20
C5587 _333_/D _225_/X 0.00469f
C5588 _271_/A _321_/a_193_7# 9.64e-20
C5589 _327_/a_1270_373# _331_/CLK 6.4e-19
C5590 _321_/a_639_7# _321_/Q 0.0047f
C5591 _197_/a_27_7# _147_/Y 2.87e-21
C5592 output36/a_27_7# VGND 0.0997f
C5593 _319_/Q ctlp[5] 4.7e-19
C5594 _258_/S _313_/a_448_7# 1.28e-20
C5595 repeater43/X _316_/a_761_249# 0.00515f
C5596 _337_/Q _263_/B 0.0613f
C5597 _281_/Y _203_/a_80_n19# 0.00283f
C5598 _305_/a_439_7# _336_/D 3.18e-19
C5599 _311_/a_651_373# _310_/a_761_249# 4.5e-21
C5600 _311_/a_1108_7# _310_/a_1283_n19# 9.8e-21
C5601 _311_/a_761_249# _310_/a_651_373# 6.62e-21
C5602 _311_/a_1283_n19# _310_/a_1108_7# 2.04e-19
C5603 _321_/a_651_373# VPWR 0.00771f
C5604 _321_/a_1108_7# VGND -0.00653f
C5605 _248_/A _347_/D 0.0333f
C5606 _283_/Y _306_/S 2.44e-19
C5607 rstn _335_/a_193_7# 0.55f
C5608 repeater43/X _320_/Q 0.141f
C5609 _341_/a_1283_n19# _304_/S 0.00132f
C5610 _331_/CLK _347_/D 4.53e-21
C5611 _330_/D _283_/A 1.67e-19
C5612 _306_/X _284_/A 0.0348f
C5613 _153_/a_297_257# VGND -0.00156f
C5614 _153_/a_487_257# VPWR -0.00117f
C5615 _224_/a_250_257# _217_/A 0.00246f
C5616 output31/a_27_7# _311_/a_1108_7# 7.66e-20
C5617 _332_/D _333_/Q 3.41e-20
C5618 _340_/CLK _190_/A 0.00332f
C5619 _246_/B _243_/a_113_257# 0.0425f
C5620 _279_/Y _206_/A 5.6e-20
C5621 _326_/a_448_7# _326_/D 0.00458f
C5622 _272_/a_39_257# _326_/Q 0.0246f
C5623 _326_/a_193_7# repeater43/X 0.0377f
C5624 _145_/A _181_/X 0.00681f
C5625 _170_/a_76_159# _346_/D 0.00255f
C5626 cal _333_/a_1108_7# 2.26e-21
C5627 _305_/a_505_n19# _193_/Y 2.48e-19
C5628 _273_/A _347_/D 6.44e-20
C5629 _281_/A _330_/a_761_249# 2.59e-19
C5630 _274_/a_39_257# _275_/A 0.00354f
C5631 _310_/a_1217_7# VGND 9.41e-20
C5632 _199_/a_250_257# VPWR 0.0256f
C5633 _307_/X _341_/a_1283_n19# 2.58e-19
C5634 _182_/X _146_/a_29_271# 4.48e-20
C5635 _185_/A _323_/a_448_7# 0.00195f
C5636 _297_/A _301_/X 8.7e-19
C5637 _296_/Y _304_/a_578_7# 1.65e-19
C5638 _343_/CLK _204_/a_27_257# 0.00384f
C5639 _341_/a_1108_7# _149_/A 6.7e-19
C5640 clkbuf_2_1_0_clk/A _346_/D 1.31e-20
C5641 _343_/CLK _208_/a_493_257# 1.74e-19
C5642 _279_/Y _156_/a_39_257# 0.00441f
C5643 _302_/a_77_159# _347_/a_193_7# 6.82e-19
C5644 _346_/a_1602_7# _346_/SET_B 0.065f
C5645 _325_/a_543_7# _181_/X 0.0138f
C5646 _169_/B VGND 0.166f
C5647 _169_/Y VPWR 0.123f
C5648 _325_/a_1108_7# _286_/B 7.61e-21
C5649 _209_/a_109_7# VGND -0.0011f
C5650 _163_/a_215_7# _346_/SET_B 3.34e-19
C5651 _347_/Q _314_/a_1108_7# 1.29e-19
C5652 _225_/B VPWR 0.907f
C5653 _300_/Y _314_/a_193_7# 1.73e-20
C5654 _339_/a_1283_n19# _338_/a_651_373# 1.05e-19
C5655 output33/a_27_7# _312_/a_27_7# 9.67e-21
C5656 _197_/X _340_/Q 0.4f
C5657 _319_/Q _318_/Q 5.23e-19
C5658 repeater43/X _334_/a_27_7# 0.0204f
C5659 _339_/Q _263_/B 0.00197f
C5660 _285_/A _297_/Y 8.61e-19
C5661 _337_/a_543_7# _340_/CLK 0.0358f
C5662 _335_/a_448_7# _335_/Q 1.26e-19
C5663 _335_/a_1108_7# _204_/Y 8.41e-19
C5664 _172_/A _185_/A 9.57e-19
C5665 _292_/A _267_/B 0.00816f
C5666 _326_/Q VGND 0.851f
C5667 _160_/X _170_/a_489_373# 0.0241f
C5668 _279_/Y _147_/A 0.00933f
C5669 _271_/A _315_/a_27_7# 1.76e-19
C5670 repeater43/X _341_/a_1462_7# -9.14e-19
C5671 _321_/D _248_/A 0.00248f
C5672 _309_/a_543_7# _265_/B 0.00281f
C5673 _344_/a_193_7# _297_/Y 0.0196f
C5674 output15/a_27_7# result[6] 4.11e-20
C5675 ctlp[1] output28/a_27_7# 6.2e-19
C5676 _147_/Y _284_/A 0.111f
C5677 _334_/a_761_249# _207_/C 0.0219f
C5678 _215_/A _324_/D 2.32e-20
C5679 _285_/A _310_/a_193_7# 6.04e-21
C5680 _321_/D _331_/CLK 0.327f
C5681 _315_/a_1283_n19# VGND 0.0197f
C5682 _344_/a_1056_7# _290_/A 4.13e-19
C5683 _315_/a_448_7# VPWR -6.06e-19
C5684 _284_/a_121_257# _309_/Q 3.27e-20
C5685 en VPWR 0.239f
C5686 output39/a_27_7# VGND 0.0983f
C5687 _320_/a_193_7# _319_/D 1.94e-19
C5688 _336_/a_1217_7# VPWR 7.39e-21
C5689 _336_/a_639_7# VGND -0.00112f
C5690 _324_/a_639_7# _227_/A 8.48e-19
C5691 _324_/a_193_7# _324_/a_448_7# -0.00831f
C5692 _235_/a_113_257# _217_/A 7.29e-19
C5693 _346_/a_27_7# clkbuf_2_3_0_clk/A 7.4e-20
C5694 _172_/A _297_/Y 0.00903f
C5695 _334_/a_1108_7# _343_/CLK 1.38e-20
C5696 _334_/a_1283_n19# _334_/D 0.0534f
C5697 _334_/a_27_7# _334_/Q 2.17e-20
C5698 clk _333_/D 1.61e-20
C5699 _291_/a_39_257# _311_/a_1108_7# 6.55e-19
C5700 _337_/Q _194_/A 0.0901f
C5701 output7/a_27_7# _334_/a_1283_n19# 0.0111f
C5702 _314_/a_193_7# VGND -0.00277f
C5703 _227_/A _297_/B 0.0435f
C5704 _314_/a_543_7# VPWR 0.0239f
C5705 _346_/SET_B _319_/a_448_7# 0.00235f
C5706 _344_/a_1032_373# comp 2.75e-19
C5707 _346_/SET_B _313_/a_27_7# 0.0126f
C5708 _283_/Y _283_/A 0.0186f
C5709 _338_/a_193_7# _337_/Q 1.89e-20
C5710 _338_/a_1108_7# _337_/D 4.71e-20
C5711 _338_/D _337_/a_1108_7# 8.27e-20
C5712 _346_/SET_B _337_/a_1283_n19# 0.00277f
C5713 clk _332_/a_193_7# 0.215f
C5714 _224_/a_256_7# VGND 4.17e-19
C5715 _224_/a_584_7# VPWR -5.99e-19
C5716 _340_/D _254_/B 2.43e-21
C5717 _341_/D _343_/CLK 0.00454f
C5718 _324_/a_761_249# _324_/D 0.043f
C5719 _324_/a_1108_7# _304_/X 1.31e-19
C5720 _341_/Q _246_/B 1.44e-20
C5721 _314_/a_27_7# _314_/Q 7.86e-20
C5722 _314_/a_1283_n19# _314_/D 1.29e-20
C5723 _314_/a_1108_7# _297_/B 3.88e-21
C5724 _311_/D _310_/a_543_7# 2.16e-19
C5725 _170_/a_226_7# VGND 0.014f
C5726 _170_/a_226_257# VPWR -7.89e-19
C5727 _258_/S _337_/Q 0.306f
C5728 input4/X _333_/Q 2.96e-19
C5729 _338_/D _343_/CLK 0.05f
C5730 _322_/a_448_7# _269_/A 0.00399f
C5731 _341_/a_651_373# _145_/A 1.5e-20
C5732 repeater43/X _207_/X 0.296f
C5733 _346_/a_27_7# _172_/Y 1.27e-20
C5734 _334_/a_27_7# _191_/B 7.41e-20
C5735 _325_/a_448_7# _325_/D 0.0145f
C5736 _339_/a_543_7# _340_/CLK 0.00171f
C5737 _288_/A _344_/Q 0.00254f
C5738 _163_/a_292_257# _345_/Q 4.2e-19
C5739 _163_/a_78_159# _345_/D 1.69e-19
C5740 _185_/A _244_/B 1.61e-20
C5741 _323_/a_761_249# _175_/Y 1.82e-19
C5742 _154_/A VGND 0.292f
C5743 _304_/X _324_/D 0.144f
C5744 _169_/Y _306_/a_76_159# 1.33e-19
C5745 cal _176_/a_27_7# 0.00918f
C5746 _340_/a_543_7# _337_/Q 1.02e-19
C5747 _327_/a_639_7# _212_/X 0.00103f
C5748 _326_/a_1462_7# repeater43/X 0.00116f
C5749 _162_/X _344_/Q 0.473f
C5750 _326_/a_761_249# _331_/a_1108_7# 5.73e-21
C5751 _326_/a_651_373# _331_/a_27_7# 5.74e-20
C5752 _207_/C _333_/Q 0.211f
C5753 _162_/a_27_7# _162_/A 0.0366f
C5754 _326_/a_1270_373# _217_/X 5.91e-19
C5755 _326_/D _222_/a_256_7# 6.2e-19
C5756 _149_/A _334_/a_1283_n19# 1.14e-19
C5757 output24/a_27_7# output25/a_27_7# 0.0246f
C5758 _271_/A _298_/B 0.0211f
C5759 _277_/A _320_/a_27_7# 0.0197f
C5760 _281_/Y _330_/a_805_7# 5.18e-20
C5761 _346_/a_476_7# _254_/A 2.18e-19
C5762 _304_/S _248_/A 4.04e-19
C5763 _185_/A _323_/D 0.159f
C5764 _277_/Y _311_/a_193_7# 7.32e-20
C5765 _168_/a_109_7# _162_/X 0.0312f
C5766 _342_/a_651_373# _269_/A 0.00187f
C5767 repeater43/a_27_7# _206_/A 3.48e-21
C5768 _334_/Q _207_/X 0.0465f
C5769 ctln[6] _333_/a_1283_n19# 6.27e-21
C5770 _328_/a_1270_373# _212_/X 2.78e-20
C5771 _328_/a_651_373# _217_/X 0.00178f
C5772 _308_/a_218_334# _227_/A 7.68e-20
C5773 _324_/Q _181_/X 0.411f
C5774 _339_/Q _194_/A 2.83e-19
C5775 _304_/S _331_/CLK 7.6e-19
C5776 _281_/Y _297_/A 1.88e-20
C5777 _320_/Q result[6] 0.045f
C5778 _173_/a_489_373# _345_/D 4.64e-19
C5779 _173_/a_226_257# _345_/Q 0.00118f
C5780 output41/a_27_7# _286_/Y 7.12e-20
C5781 _347_/Q _297_/B 0.0741f
C5782 _339_/Q _338_/a_193_7# 3.12e-19
C5783 _339_/a_1283_n19# _346_/SET_B -6.5e-19
C5784 _339_/a_1108_7# _338_/D 5.07e-20
C5785 trim[2] _312_/a_1108_7# 4.32e-19
C5786 repeater43/a_27_7# _334_/D 0.0059f
C5787 repeater43/X _334_/a_1217_7# -2.64e-19
C5788 _194_/A _202_/a_256_7# 5.76e-19
C5789 _218_/a_250_257# _304_/X 8.76e-19
C5790 _232_/X _242_/A 0.265f
C5791 _258_/a_76_159# _336_/a_761_249# 7.92e-19
C5792 _258_/a_505_n19# _336_/a_193_7# 0.00442f
C5793 output7/a_27_7# repeater43/a_27_7# 2.93e-20
C5794 _277_/Y output9/a_27_7# 0.00104f
C5795 output10/a_27_7# _275_/Y 5.03e-21
C5796 _335_/D _335_/Q 0.0116f
C5797 _258_/S _339_/Q 0.0609f
C5798 _273_/A _304_/S 0.00306f
C5799 _324_/Q _304_/a_288_7# 1.44e-19
C5800 _200_/a_584_7# _337_/Q 8.95e-19
C5801 _210_/a_27_7# _179_/a_27_7# 7.78e-20
C5802 clkbuf_0_clk/X _216_/X 0.222f
C5803 _313_/a_27_7# _313_/a_761_249# -0.0166f
C5804 _164_/Y _344_/D 2.26e-20
C5805 _271_/A _242_/B 0.102f
C5806 clkbuf_1_0_0_clk/a_75_172# _330_/a_651_373# 8.6e-19
C5807 clkbuf_2_3_0_clk/A _338_/Q 0.659f
C5808 output37/a_27_7# VPWR 0.149f
C5809 _251_/a_297_257# _162_/X 0.00567f
C5810 _275_/A clkbuf_2_3_0_clk/A 0.0901f
C5811 _235_/a_199_7# VGND 2.85e-20
C5812 _225_/X _190_/A 0.0123f
C5813 _340_/a_651_373# _339_/D 1.44e-20
C5814 _329_/Q clkbuf_0_clk/X 0.0456f
C5815 clk _208_/a_78_159# 0.0698f
C5816 _317_/a_27_7# _248_/A 0.00127f
C5817 _304_/S _222_/a_93_n19# 7.74e-20
C5818 _187_/a_27_7# VPWR 0.0767f
C5819 _327_/a_761_249# clkbuf_0_clk/X 0.0373f
C5820 _315_/D VPWR 0.61f
C5821 _279_/Y _339_/D 3.17e-19
C5822 _220_/a_250_257# _278_/a_68_257# 4.46e-19
C5823 output6/a_27_7# ctln[0] 0.00443f
C5824 _343_/a_27_7# _271_/A 3.94e-21
C5825 _321_/Q _318_/a_193_7# 2.81e-21
C5826 _340_/a_1283_n19# _202_/a_250_257# 5.35e-20
C5827 _340_/a_1108_7# _202_/a_93_n19# 4.98e-20
C5828 _275_/A _327_/Q 0.0059f
C5829 _324_/a_1108_7# VGND 0.00957f
C5830 _324_/a_651_373# VPWR 0.00166f
C5831 _281_/Y _192_/a_68_257# 6.91e-19
C5832 _317_/a_27_7# _331_/CLK 0.0267f
C5833 repeater43/X _226_/a_79_n19# 3.24e-19
C5834 _306_/a_535_334# clkbuf_2_1_0_clk/A 2.21e-19
C5835 _322_/D _232_/X 3.76e-21
C5836 _273_/A _267_/B 0.0609f
C5837 _275_/A _172_/Y 4.32e-20
C5838 _283_/A _312_/a_27_7# 1.02e-19
C5839 _314_/a_1462_7# VGND 2.24e-19
C5840 _346_/SET_B _313_/a_1217_7# -3.08e-19
C5841 _343_/a_448_7# VPWR 0.00285f
C5842 _343_/a_1283_n19# VGND 0.034f
C5843 _181_/X _281_/A 1.72e-20
C5844 _340_/a_1283_n19# input1/X 1.29e-21
C5845 _340_/a_1108_7# cal 3.96e-20
C5846 result[2] _317_/D 6.6e-20
C5847 _324_/D VGND 0.264f
C5848 _242_/A _244_/B 1.8e-20
C5849 _220_/a_93_n19# _279_/A 0.00254f
C5850 output20/a_27_7# VGND 0.125f
C5851 _252_/a_109_257# _251_/X 3.86e-19
C5852 input4/X _339_/a_761_249# 2.19e-22
C5853 _328_/a_193_7# clkbuf_0_clk/X 4.46e-21
C5854 _314_/a_1217_7# _314_/Q 1.43e-19
C5855 _344_/a_476_7# _265_/B 2.46e-19
C5856 rstn _197_/X 2.32e-20
C5857 _236_/B _331_/a_193_7# 0.00158f
C5858 _196_/A _344_/D 1.22e-19
C5859 _340_/a_193_7# _260_/A 3.55e-19
C5860 _331_/CLK _331_/a_543_7# 0.00123f
C5861 _231_/a_79_n19# _283_/A 4.9e-19
C5862 _158_/Y _288_/Y 2.9e-19
C5863 _313_/a_27_7# _147_/A 0.226f
C5864 _341_/a_761_249# _286_/Y 0.0431f
C5865 _341_/a_27_7# sample 0.00267f
C5866 _344_/a_27_7# _169_/Y 1.37e-21
C5867 _278_/a_150_257# VGND -3.64e-19
C5868 _345_/a_1602_7# VGND 0.0241f
C5869 _345_/a_562_373# VPWR 0.00236f
C5870 _181_/X _228_/A 0.17f
C5871 _260_/B _197_/a_27_7# 1.07e-21
C5872 _346_/Q _196_/A 9.79e-21
C5873 _162_/X _306_/S 0.0182f
C5874 _292_/Y output16/a_27_7# 2.67e-19
C5875 _160_/A _174_/a_373_7# 2.63e-21
C5876 _309_/Q VGND 0.183f
C5877 _292_/A _261_/a_109_257# 5.6e-20
C5878 _283_/A _330_/a_1283_n19# 0.0087f
C5879 _320_/D _242_/A 0.0795f
C5880 _281_/Y _256_/a_209_257# 0.00429f
C5881 _214_/a_27_257# _326_/Q 0.00103f
C5882 clk _334_/a_543_7# 0.00335f
C5883 _186_/a_297_7# _341_/Q 1.85e-19
C5884 _220_/a_93_n19# _220_/a_346_7# -3.48e-20
C5885 _326_/D _331_/a_193_7# 1.44e-20
C5886 _330_/Q _218_/a_584_7# 5.4e-19
C5887 _307_/a_76_159# _150_/C 9.02e-22
C5888 _283_/A _333_/a_27_7# 0.0865f
C5889 _172_/A _336_/Q 1.45e-20
C5890 _330_/Q _246_/B 0.0356f
C5891 _341_/a_651_373# _324_/Q 2.69e-21
C5892 _307_/X _307_/a_505_n19# 2.23e-19
C5893 _188_/a_76_159# _145_/A 0.0409f
C5894 clkbuf_2_3_0_clk/A _345_/D 2e-20
C5895 _279_/A VGND 0.488f
C5896 _275_/Y _347_/Q 7.98e-21
C5897 _231_/a_79_n19# _248_/B 4.84e-20
C5898 _326_/a_1283_n19# _280_/a_68_257# 2.41e-21
C5899 _337_/Q _201_/a_27_7# 1.84e-19
C5900 _222_/a_584_7# _217_/X 0.00168f
C5901 _197_/X _225_/a_59_35# 2.42e-19
C5902 _218_/a_346_7# VPWR -4.95e-19
C5903 _218_/a_250_257# VGND -0.00585f
C5904 _216_/X _286_/Y 0.0814f
C5905 _333_/a_193_7# _205_/a_79_n19# 2.96e-20
C5906 _318_/Q _325_/Q 1.97e-21
C5907 _198_/a_93_n19# _225_/B 9.5e-20
C5908 _198_/a_250_257# _336_/Q 0.00359f
C5909 _342_/a_1108_7# _175_/Y 0.0014f
C5910 _178_/a_27_7# _225_/X 2.7e-21
C5911 _309_/a_761_249# _309_/Q 6.18e-20
C5912 _307_/X _178_/a_27_7# 0.0828f
C5913 _308_/a_76_159# VPWR 0.0183f
C5914 _286_/B _250_/X 2.68e-20
C5915 _181_/X _216_/A 0.0378f
C5916 _259_/a_113_257# _290_/A 1.04e-20
C5917 _329_/Q _286_/Y 1.8e-20
C5918 _343_/a_27_7# _323_/a_27_7# 6.95e-19
C5919 _345_/D _172_/Y 2.83e-19
C5920 _209_/X _254_/B 0.00879f
C5921 _294_/A _288_/A 0.00736f
C5922 _226_/a_297_7# _150_/C 0.00141f
C5923 _220_/a_346_7# VGND 1.39e-20
C5924 _311_/a_543_7# VPWR 0.033f
C5925 _157_/A _295_/a_79_n19# 9.2e-20
C5926 _311_/a_193_7# VGND 0.00857f
C5927 _194_/A _336_/D 0.0298f
C5928 cal _334_/a_761_249# 2.63e-19
C5929 _306_/X _336_/a_27_7# 0.00496f
C5930 _313_/Q _336_/a_193_7# 9e-19
C5931 _325_/a_448_7# _248_/A 4.06e-20
C5932 _254_/A clkbuf_2_3_0_clk/A 0.0153f
C5933 _294_/A _162_/X 2.26e-21
C5934 _281_/Y _325_/D 4.97e-19
C5935 _304_/a_288_7# _216_/A 8.42e-19
C5936 _294_/A _287_/a_39_257# 4.05e-19
C5937 _342_/a_761_249# _298_/A 6.96e-19
C5938 _346_/Q _347_/a_1283_n19# 1.76e-20
C5939 _232_/a_27_7# _242_/B 0.00772f
C5940 _325_/a_448_7# _331_/CLK 2.63e-20
C5941 _325_/a_1108_7# _316_/D 5.84e-21
C5942 _258_/S _336_/D 8.1e-20
C5943 _271_/A ctln[0] 1.8e-20
C5944 _271_/Y _269_/Y 0.0306f
C5945 _318_/Q _321_/a_1108_7# 1.44e-20
C5946 _337_/a_27_7# _337_/Q 0.00356f
C5947 _337_/a_1283_n19# _337_/D 3.61e-20
C5948 _200_/a_346_7# _267_/A 9.56e-19
C5949 _242_/A _241_/a_113_257# 1.88e-19
C5950 _316_/Q _318_/a_761_249# 6.34e-21
C5951 output32/a_27_7# _310_/a_27_7# 1.28e-20
C5952 _165_/X _299_/a_215_7# 1.86e-19
C5953 _335_/a_193_7# VPWR -0.307f
C5954 clk _190_/A 0.0276f
C5955 output9/a_27_7# VGND 0.0684f
C5956 repeater43/X _323_/Q 0.263f
C5957 _304_/S _217_/X 2.35e-20
C5958 _342_/Q _333_/a_1108_7# 4.15e-21
C5959 _265_/B _254_/B 3.99e-20
C5960 _341_/Q _154_/a_27_7# 0.0109f
C5961 _271_/A _318_/a_1283_n19# 0.00202f
C5962 _336_/Q _203_/a_80_n19# 0.0433f
C5963 _144_/A _147_/A 1.18e-20
C5964 _340_/a_1108_7# _284_/A 3.49e-19
C5965 _340_/a_543_7# _336_/D 1.28e-19
C5966 _327_/a_27_7# _221_/a_93_n19# 3.21e-20
C5967 _275_/Y _297_/B 1.08f
C5968 _254_/A _313_/a_1270_373# 9.87e-20
C5969 _317_/Q _331_/Q 1.09e-20
C5970 _297_/A _297_/Y 0.00112f
C5971 _338_/a_27_7# _194_/X 0.0114f
C5972 _346_/Q _165_/a_78_159# 1.9e-20
C5973 _158_/Y _172_/a_109_257# 8.43e-21
C5974 _339_/Q _201_/a_27_7# 0.00101f
C5975 _260_/B _284_/A 0.096f
C5976 _144_/A _149_/A 0.00169f
C5977 _318_/a_805_7# VPWR 3.1e-19
C5978 _318_/a_1270_373# VGND 3.66e-20
C5979 clkbuf_2_3_0_clk/A _309_/D 0.0102f
C5980 _341_/a_651_373# _228_/A 9.64e-20
C5981 _196_/A _340_/D 0.0109f
C5982 _346_/SET_B _174_/a_27_257# 0.00612f
C5983 _144_/a_27_7# _223_/a_250_257# 1.21e-21
C5984 _164_/A _297_/Y 0.00553f
C5985 _307_/a_439_7# _296_/Y 5.37e-22
C5986 _311_/Q _310_/Q 0.00335f
C5987 _280_/a_68_257# _248_/A 0.00516f
C5988 _162_/X _283_/A 0.0101f
C5989 _181_/a_27_7# _215_/A 0.0292f
C5990 _309_/a_651_373# VPWR 0.0113f
C5991 _309_/a_1108_7# VGND -0.00196f
C5992 cal _333_/Q 6.44e-20
C5993 _313_/a_1217_7# _147_/A 9.92e-19
C5994 repeater43/X _317_/a_1283_n19# 0.00303f
C5995 _296_/Y _304_/S 0.00107f
C5996 clkbuf_2_0_0_clk/a_75_172# _197_/X 9.64e-21
C5997 _340_/a_193_7# _340_/Q 0.0168f
C5998 _340_/a_27_7# _306_/S 0.00956f
C5999 _340_/a_761_249# _194_/X 5.58e-19
C6000 _258_/a_505_n19# _299_/X 1.68e-22
C6001 _315_/a_543_7# _317_/D 0.00542f
C6002 ctln[5] _195_/a_27_257# 0.0021f
C6003 _331_/CLK _280_/a_68_257# 0.0577f
C6004 _167_/a_27_257# _286_/B 7.88e-20
C6005 _269_/A output41/a_27_7# 0.0186f
C6006 _336_/a_27_7# _147_/Y 0.223f
C6007 _273_/A _301_/X 2.32e-20
C6008 _305_/a_505_n19# _215_/A 4.06e-22
C6009 _220_/a_250_257# _328_/D 2.93e-19
C6010 _321_/a_543_7# _322_/Q 0.00155f
C6011 _339_/D _337_/a_1283_n19# 1.92e-19
C6012 _339_/Q _337_/a_27_7# 0.042f
C6013 _322_/a_27_7# _318_/D 4.53e-21
C6014 _307_/a_76_159# _183_/a_471_7# 9.38e-22
C6015 repeater43/X _331_/a_651_373# 0.00359f
C6016 repeater43/X result[7] 0.00209f
C6017 _191_/B _323_/Q 0.0398f
C6018 _318_/Q _326_/Q 0.00282f
C6019 _145_/A _147_/A 0.013f
C6020 _283_/A _333_/a_1217_7# 8.61e-19
C6021 _331_/a_27_7# _331_/a_761_249# -0.0166f
C6022 _307_/X _296_/Y 6.95e-19
C6023 _306_/S _298_/C 0.539f
C6024 _309_/a_193_7# _309_/a_448_7# -0.00297f
C6025 _331_/a_543_7# _217_/X 3.33e-22
C6026 _331_/a_1108_7# _327_/Q 1.3e-20
C6027 _331_/a_1283_n19# _212_/X 2.75e-20
C6028 _162_/X _248_/B 6.56e-20
C6029 _185_/A _177_/A 3.61e-20
C6030 _255_/B _286_/B 0.642f
C6031 _325_/a_761_249# _304_/S 0.00136f
C6032 _257_/a_79_159# _286_/B 0.00147f
C6033 _346_/a_476_7# _286_/Y 1.93e-20
C6034 _316_/Q result[1] 0.0104f
C6035 _343_/D output41/a_27_7# 0.00209f
C6036 _323_/a_193_7# VPWR 0.0441f
C6037 _145_/A _149_/A 0.00711f
C6038 _183_/a_27_7# _178_/a_27_7# 1.51e-20
C6039 _333_/a_448_7# _335_/Q 1.9e-20
C6040 _146_/a_112_13# _147_/A 3.87e-19
C6041 _297_/A _242_/A 1.44e-20
C6042 _307_/X _146_/a_29_271# 0.0109f
C6043 _308_/S VPWR 0.316f
C6044 _320_/a_193_7# _297_/B 0.589f
C6045 cal _337_/a_761_249# 6.9e-20
C6046 _306_/a_439_7# VGND -3.8e-19
C6047 _328_/a_448_7# _281_/A 3.79e-21
C6048 output12/a_27_7# _340_/CLK 7.22e-19
C6049 _200_/a_346_7# _194_/X 8.79e-19
C6050 _200_/a_256_7# _340_/Q 7.43e-19
C6051 _200_/a_93_n19# _193_/Y 0.0229f
C6052 clkbuf_2_1_0_clk/A _254_/B 0.00698f
C6053 _256_/a_80_n19# _342_/Q 1.98e-19
C6054 _254_/Y _162_/X 1.92e-21
C6055 _304_/a_79_n19# _144_/a_27_7# 5.09e-21
C6056 _311_/a_1462_7# VGND 1.14e-19
C6057 _263_/B _310_/a_1283_n19# 3.18e-19
C6058 _313_/Q _336_/a_1462_7# 3.43e-21
C6059 _259_/a_113_257# _310_/a_27_7# 2.65e-19
C6060 _327_/a_1283_n19# _329_/D 7.11e-19
C6061 _186_/a_382_257# VPWR 7.53e-21
C6062 repeater42/a_27_7# _330_/D 8.24e-20
C6063 _320_/Q clkbuf_1_0_0_clk/a_75_172# 2.46e-20
C6064 _149_/a_27_7# _150_/C 0.00619f
C6065 _325_/Q _223_/a_346_7# 0.00422f
C6066 _335_/a_27_7# _335_/a_448_7# -0.00972f
C6067 _335_/a_193_7# _335_/a_1108_7# -0.0069f
C6068 _329_/a_193_7# _216_/X 0.0011f
C6069 _216_/X _328_/Q 0.0486f
C6070 _345_/a_1032_373# _344_/a_476_7# 2.35e-20
C6071 trim[1] _310_/a_1108_7# 2.62e-19
C6072 _250_/a_292_257# _190_/A 2.31e-20
C6073 _328_/a_1283_n19# _319_/Q 0.00429f
C6074 _254_/A _302_/a_227_7# 0.00588f
C6075 _335_/a_805_7# VGND 1.67e-19
C6076 _335_/a_1462_7# VPWR 5.65e-20
C6077 _341_/a_761_249# _269_/A 1.62e-19
C6078 _343_/a_193_7# _342_/a_761_249# 1.17e-20
C6079 _343_/a_761_249# _342_/a_193_7# 9.63e-20
C6080 _343_/a_543_7# _342_/a_27_7# 3.98e-21
C6081 _343_/a_27_7# _342_/a_543_7# 3.58e-21
C6082 _329_/a_193_7# _329_/Q -8.97e-20
C6083 _329_/Q _328_/Q 0.236f
C6084 _169_/Y _147_/Y 0.167f
C6085 _183_/a_1241_257# _144_/A 0.0045f
C6086 _339_/a_27_7# _339_/Q 1.9e-19
C6087 _153_/B VGND 0.483f
C6088 clkbuf_2_1_0_clk/A _331_/D 5.41e-20
C6089 _268_/a_39_257# _232_/A 8.68e-21
C6090 _225_/B _147_/Y 0.688f
C6091 _328_/a_543_7# _329_/D 9.92e-20
C6092 clkbuf_2_1_0_clk/A _330_/a_193_7# 1.08e-21
C6093 _320_/a_1108_7# _279_/A 1.65e-19
C6094 clkbuf_0_clk/X clkbuf_2_3_0_clk/A 0.00819f
C6095 _329_/a_543_7# _327_/a_27_7# 1.53e-20
C6096 _329_/a_27_7# _327_/a_543_7# 8.4e-21
C6097 _327_/a_761_249# _328_/Q 1.33e-19
C6098 _338_/D _195_/a_109_257# 6.84e-20
C6099 _338_/a_805_7# _340_/Q 4.47e-19
C6100 _338_/a_1217_7# _194_/X 1.84e-19
C6101 _346_/SET_B _195_/a_27_257# 0.00123f
C6102 _289_/a_39_257# _310_/D 3.72e-19
C6103 _346_/SET_B _281_/A 0.185f
C6104 _345_/a_381_7# _172_/A 6.7e-20
C6105 cal _226_/a_297_7# 0.00114f
C6106 _325_/a_805_7# repeater43/X -0.00104f
C6107 output19/a_27_7# VPWR 0.0927f
C6108 _216_/a_27_7# _286_/Y 0.0122f
C6109 clkbuf_0_clk/X _327_/Q 0.108f
C6110 _325_/a_651_373# _212_/X 0.00151f
C6111 _343_/CLK output30/a_27_7# 0.0156f
C6112 _275_/Y _309_/a_639_7# 5.97e-19
C6113 _340_/a_27_7# _283_/A 2.04e-20
C6114 trim[0] _311_/a_27_7# 2.42e-20
C6115 _293_/a_121_257# VGND -1.87e-19
C6116 _338_/Q _261_/A 0.0329f
C6117 _281_/Y _248_/A 0.00541f
C6118 _328_/a_193_7# _328_/Q 0.00857f
C6119 _269_/A _316_/a_543_7# 4.01e-19
C6120 _340_/a_805_7# _193_/Y 6.41e-19
C6121 _340_/a_1462_7# _340_/Q 0.00218f
C6122 _174_/a_27_257# _147_/A 4.88e-19
C6123 _182_/a_79_n19# _298_/A 0.00441f
C6124 _274_/a_39_257# _240_/B 1.59e-19
C6125 _275_/A _239_/a_113_257# 0.0629f
C6126 _313_/Q _299_/X 1.8e-20
C6127 _230_/a_27_7# _316_/a_27_7# 5.58e-21
C6128 _345_/a_27_7# _172_/B 0.0129f
C6129 _336_/a_1217_7# _147_/Y 9.39e-19
C6130 _188_/a_76_159# _228_/A 1.23e-21
C6131 clkbuf_2_3_0_clk/A input1/X 0.176f
C6132 _322_/a_1108_7# _321_/Q 0.0166f
C6133 _341_/a_1108_7# _255_/B 4.22e-22
C6134 _281_/Y _331_/CLK 0.0157f
C6135 _283_/Y ctln[0] 0.0198f
C6136 ctln[7] _269_/Y 9.86e-20
C6137 _270_/a_121_257# _316_/a_193_7# 8.88e-20
C6138 _283_/A _298_/C 1.16f
C6139 _346_/a_1032_373# _166_/Y 0.011f
C6140 ctln[6] _332_/Q 0.0393f
C6141 _296_/Y _183_/a_27_7# 0.0039f
C6142 _281_/Y _190_/A 0.164f
C6143 _311_/a_27_7# _311_/Q 7.06e-20
C6144 _254_/A _157_/A 3.51e-19
C6145 _181_/a_27_7# VGND 0.0892f
C6146 _296_/Y clk 4.83e-21
C6147 _218_/a_256_7# _232_/X 4.9e-19
C6148 _343_/a_543_7# _317_/D 1.39e-20
C6149 _322_/a_193_7# VGND 0.00695f
C6150 _322_/a_543_7# VPWR 0.0225f
C6151 _166_/Y _331_/CLK 3.09e-20
C6152 _281_/Y _273_/A 0.0256f
C6153 _161_/Y _297_/B 0.0027f
C6154 _164_/Y _265_/B 0.00911f
C6155 _170_/a_226_257# _147_/Y 6.85e-19
C6156 _337_/a_761_249# _284_/A 4.17e-21
C6157 _308_/S _184_/a_505_n19# 2.92e-20
C6158 _308_/a_505_n19# _188_/S 1.33e-20
C6159 _320_/a_1270_373# VGND 6.61e-20
C6160 _346_/a_193_7# _167_/X 0.00258f
C6161 _346_/a_27_7# _165_/X 0.00144f
C6162 _329_/D _248_/A 1.05e-20
C6163 _316_/a_27_7# _232_/A 0.0106f
C6164 _319_/Q _316_/D 0.00761f
C6165 _323_/a_1462_7# VPWR 4.51e-19
C6166 _323_/a_805_7# VGND 1.41e-19
C6167 _216_/A _346_/SET_B 0.118f
C6168 ctlp[5] _279_/A 0.244f
C6169 _333_/D _335_/Q 0.00502f
C6170 clkbuf_0_clk/X _192_/B 3.43e-19
C6171 _322_/a_1283_n19# _318_/a_761_249# 5.61e-22
C6172 _214_/a_373_7# VGND -2.54e-19
C6173 _322_/a_448_7# _318_/a_27_7# 3.29e-21
C6174 _305_/a_535_334# VPWR 7.41e-20
C6175 _344_/a_1032_373# VGND 0.00403f
C6176 _344_/a_381_7# VPWR 0.00488f
C6177 _305_/a_505_n19# VGND 0.0659f
C6178 _291_/a_39_257# _263_/B 3.28e-21
C6179 _232_/X _220_/a_584_7# 2.12e-19
C6180 _292_/A _297_/Y 0.257f
C6181 _280_/a_68_257# _217_/X 2e-20
C6182 _273_/A _166_/Y 0.00867f
C6183 result[3] _318_/D 0.0021f
C6184 _143_/a_109_7# _228_/A 7.8e-21
C6185 _320_/a_1462_7# _297_/B 5.26e-19
C6186 _329_/D _331_/CLK 0.0436f
C6187 _306_/S _332_/D 1.44e-20
C6188 _193_/Y _340_/CLK 0.0201f
C6189 _172_/A _271_/A 0.0155f
C6190 _196_/A _209_/X 1.35e-20
C6191 _212_/a_27_7# _246_/B 2.01e-21
C6192 _332_/a_27_7# _204_/Y 4.99e-21
C6193 _332_/a_193_7# _335_/Q 4.09e-19
C6194 _274_/a_39_257# _328_/Q 0.0256f
C6195 _324_/Q _147_/A 6.65e-19
C6196 _254_/Y _340_/a_27_7# 1.08e-21
C6197 _326_/Q _223_/a_346_7# 2.62e-20
C6198 _248_/B _298_/C 4.53e-21
C6199 _186_/a_297_7# _184_/a_76_159# 1.3e-20
C6200 _160_/A _297_/Y 0.00757f
C6201 _162_/A clkc 0.0135f
C6202 _260_/A _313_/a_1108_7# 6.55e-20
C6203 _227_/A _333_/a_543_7# 4.16e-21
C6204 _313_/D VPWR 0.119f
C6205 clkbuf_0_clk/a_110_7# clk 0.00989f
C6206 _279_/Y _257_/a_79_159# 8.08e-20
C6207 _257_/a_544_257# _260_/B 0.0016f
C6208 _344_/Q _345_/Q 0.00421f
C6209 clkbuf_2_3_0_clk/A _286_/Y 0.0098f
C6210 _258_/S _310_/a_1283_n19# 8.98e-20
C6211 _271_/A _232_/X 0.00642f
C6212 _246_/a_109_257# VGND -9.02e-19
C6213 _324_/Q _149_/A 8.41e-20
C6214 _271_/A _335_/D 0.03f
C6215 _292_/A _310_/a_193_7# 9.64e-20
C6216 _342_/a_761_249# VGND 0.0106f
C6217 _342_/a_1283_n19# VPWR 0.056f
C6218 _335_/a_27_7# _335_/D 0.183f
C6219 repeater43/X sample 1.77e-19
C6220 input4/X _207_/a_27_7# 1.94e-19
C6221 _290_/A _163_/a_215_7# 0.00171f
C6222 _199_/a_93_n19# _312_/D 2.94e-19
C6223 result[6] result[7] 0.143f
C6224 _297_/A _314_/a_761_249# 1.1e-19
C6225 _197_/X VPWR 1.54f
C6226 _327_/Q _286_/Y 0.398f
C6227 _254_/A _260_/A 0.00916f
C6228 output31/a_27_7# _258_/S 4.05e-19
C6229 input1/X _192_/B 0.0169f
C6230 _219_/a_346_7# _212_/X 0.00182f
C6231 _319_/Q _319_/a_448_7# 2.83e-19
C6232 _322_/a_193_7# output27/a_27_7# 1.29e-20
C6233 _172_/Y _286_/Y 0.00207f
C6234 _169_/B _286_/B 0.00203f
C6235 _286_/B _209_/a_109_7# 5.66e-19
C6236 _309_/a_1283_n19# _311_/Q 7.28e-21
C6237 _329_/a_1462_7# _329_/Q 4.9e-19
C6238 _248_/a_109_257# _315_/D 5.84e-19
C6239 _287_/a_121_257# _310_/D 4.73e-19
C6240 _207_/a_27_7# _207_/C 0.0163f
C6241 _288_/A _284_/a_39_257# 1.38e-19
C6242 _320_/Q _319_/D 4.48e-20
C6243 _338_/Q _340_/Q 6.42e-19
C6244 _320_/a_27_7# _320_/a_761_249# -0.0166f
C6245 _162_/X _300_/a_27_257# 0.0984f
C6246 _323_/a_27_7# _323_/a_448_7# -0.00297f
C6247 _323_/a_193_7# _323_/a_1108_7# 1.42e-32
C6248 _157_/A _302_/a_227_257# 0.00316f
C6249 _228_/A _156_/a_39_257# 7.01e-20
C6250 _332_/a_543_7# _153_/a_215_257# 0.00145f
C6251 _332_/a_1283_n19# _153_/a_109_53# 0.00321f
C6252 _318_/Q _279_/A 0.00102f
C6253 _218_/a_93_n19# _331_/D 7.37e-21
C6254 _336_/a_761_249# _194_/A 3.18e-21
C6255 _256_/a_209_257# _336_/Q 5.97e-19
C6256 output21/a_27_7# clkbuf_2_1_0_clk/A 7.78e-20
C6257 _271_/A _244_/B 0.0104f
C6258 _294_/A output35/a_27_7# 0.0423f
C6259 _304_/a_306_329# _326_/Q 2.04e-19
C6260 _216_/A _313_/a_761_249# 0.0428f
C6261 _236_/a_109_257# _269_/A 6.1e-19
C6262 _328_/a_1462_7# _328_/Q 0.00226f
C6263 _182_/X _298_/A 8.04e-19
C6264 _283_/Y _335_/a_448_7# 1.6e-21
C6265 ctln[7] _335_/a_1283_n19# 0.022f
C6266 _258_/S _336_/a_761_249# 1.58e-19
C6267 _286_/B _336_/a_639_7# 6.89e-19
C6268 _275_/Y _161_/Y 0.161f
C6269 _228_/A _147_/A 4.13e-20
C6270 _312_/a_193_7# VPWR 0.0461f
C6271 _185_/A _248_/A 0.222f
C6272 _275_/A _165_/X 1.37e-19
C6273 _331_/Q _304_/X 0.0864f
C6274 _164_/Y _310_/Q 2.03e-21
C6275 _238_/B _242_/A 0.129f
C6276 _196_/A _314_/a_27_7# 7.22e-19
C6277 output8/a_27_7# trim[2] 3.73e-20
C6278 _325_/Q _316_/a_448_7# 4.89e-19
C6279 _208_/a_78_159# _335_/Q 0.0151f
C6280 _327_/a_1283_n19# _242_/A 1.04e-19
C6281 _149_/A _228_/A 0.284f
C6282 _311_/a_1217_7# _311_/Q 1.27e-19
C6283 _307_/a_218_334# _250_/X 1.94e-19
C6284 _145_/A _250_/a_78_159# 1.66e-19
C6285 _288_/A _262_/a_113_257# 5.07e-19
C6286 _340_/a_1283_n19# _336_/a_193_7# 2.88e-21
C6287 _340_/a_1108_7# _336_/a_27_7# 2.29e-19
C6288 _346_/a_1602_7# _167_/a_27_257# 9.48e-20
C6289 _346_/a_1032_373# _167_/a_109_257# 1.46e-19
C6290 _318_/a_651_373# _317_/D 7.21e-20
C6291 _216_/A _156_/a_39_257# 2.2e-21
C6292 _330_/D _232_/X 0.00147f
C6293 _346_/a_193_7# clkbuf_1_1_0_clk/a_75_172# 2.04e-21
C6294 _231_/a_676_257# VPWR -3.37e-19
C6295 _332_/a_543_7# _209_/a_109_257# 7.64e-21
C6296 _309_/D _261_/A 0.0136f
C6297 _325_/a_27_7# _286_/Y 0.0166f
C6298 _313_/a_639_7# _284_/A 1.32e-19
C6299 _330_/Q _330_/a_448_7# 9.9e-19
C6300 _294_/Y _346_/SET_B 8.57e-20
C6301 _260_/B _336_/a_27_7# 5.48e-19
C6302 _326_/a_1283_n19# _242_/A 0.0413f
C6303 _337_/Q _202_/a_346_7# 0.00122f
C6304 input4/X _306_/S 6.58e-19
C6305 _283_/A _332_/D 0.00586f
C6306 _289_/a_39_257# VPWR 0.0368f
C6307 _186_/a_79_n19# _172_/A 0.0522f
C6308 _250_/a_215_7# _192_/B 4e-19
C6309 _342_/Q _295_/a_512_7# 0.00439f
C6310 _330_/a_543_7# VGND 0.0185f
C6311 _330_/a_1108_7# VPWR -0.00625f
C6312 _181_/X _153_/A 5.69e-20
C6313 _258_/S _291_/a_39_257# 8.48e-21
C6314 _183_/a_1241_257# _324_/Q 0.0089f
C6315 _196_/A clkbuf_2_1_0_clk/A 0.0108f
C6316 _281_/Y _217_/X 0.0232f
C6317 _306_/S _345_/Q 0.00854f
C6318 _216_/A _147_/A 0.92f
C6319 clkbuf_0_clk/X _157_/A 0.0116f
C6320 _255_/B _316_/D 5.23e-20
C6321 _346_/SET_B _240_/a_109_257# 6.78e-19
C6322 _240_/B clkbuf_2_3_0_clk/A 4.52e-21
C6323 _325_/a_1108_7# _324_/Q 1.3e-20
C6324 _186_/a_297_7# _188_/S 0.0252f
C6325 _333_/a_193_7# VPWR -0.255f
C6326 _306_/S _207_/C 0.0165f
C6327 _306_/S _313_/a_1283_n19# 1.13e-19
C6328 _341_/a_27_7# _341_/Q -6.5e-21
C6329 _288_/A _266_/a_199_7# 5.65e-20
C6330 output32/a_27_7# _309_/Q 2.8e-19
C6331 _252_/a_109_257# VPWR 1.92e-20
C6332 _337_/a_1108_7# _340_/D 3.56e-36
C6333 _318_/Q _318_/a_1270_373# 5.47e-19
C6334 _257_/a_222_53# _190_/A 0.00108f
C6335 _319_/Q _331_/a_27_7# 1.5e-19
C6336 _232_/a_27_7# _232_/X 0.0137f
C6337 _335_/a_1217_7# _335_/D 1.14e-19
C6338 _240_/B _327_/Q 7.8e-20
C6339 _252_/a_27_7# _314_/D 0.0459f
C6340 _343_/CLK _340_/D 6.44e-20
C6341 _211_/a_109_7# _153_/B 6.1e-19
C6342 _196_/A _300_/a_735_7# 3.6e-22
C6343 _273_/A _297_/Y 1.88f
C6344 _271_/A _241_/a_113_257# 0.00891f
C6345 _314_/a_1283_n19# _347_/a_27_7# 5.44e-19
C6346 _329_/D _217_/X 0.172f
C6347 _146_/C input1/X 1.68e-20
C6348 _165_/X _345_/D 2.87e-19
C6349 _254_/A _340_/Q 0.00503f
C6350 _337_/Q _267_/A 0.257f
C6351 _325_/a_193_7# _284_/A 2.08e-21
C6352 _288_/A _160_/X 0.0075f
C6353 _343_/Q _153_/A 3.18e-20
C6354 clkbuf_2_3_0_clk/A _328_/Q 3.35e-20
C6355 _162_/X _160_/X 0.722f
C6356 _312_/a_1283_n19# _311_/a_1283_n19# 1.6e-19
C6357 _343_/CLK _247_/a_113_257# 1.1e-19
C6358 _323_/a_27_7# _323_/D 0.046f
C6359 _273_/A _310_/a_193_7# 1.21e-20
C6360 _319_/Q _217_/a_27_7# 3.41e-21
C6361 _341_/a_651_373# _315_/a_761_249# 1.59e-21
C6362 _341_/a_761_249# _315_/a_651_373# 2.64e-21
C6363 _341_/a_1270_373# _298_/A 4.54e-19
C6364 _332_/a_1283_n19# _153_/A 3.49e-21
C6365 _332_/a_761_249# _154_/A 1.31e-19
C6366 clkbuf_0_clk/X _260_/A 0.00605f
C6367 _229_/a_556_7# _175_/Y 0.0011f
C6368 ctlp[4] VGND 0.35f
C6369 _345_/a_1032_373# _164_/Y 0.00606f
C6370 repeater43/X _296_/a_109_7# 3.3e-22
C6371 _260_/B _225_/B 0.00656f
C6372 _277_/Y _312_/Q 8.5e-21
C6373 _329_/a_193_7# _327_/Q 3.09e-20
C6374 _329_/a_27_7# _212_/X 2.37e-19
C6375 _306_/S _150_/C 0.0175f
C6376 _327_/Q _328_/Q 0.316f
C6377 _344_/a_193_7# _344_/a_1602_7# -4.7e-21
C6378 _344_/a_27_7# _344_/a_381_7# -0.00844f
C6379 trim[4] _297_/Y 3.32e-19
C6380 _242_/A _248_/A 1.33f
C6381 _331_/Q VGND 0.971f
C6382 _254_/A _165_/X 0.00297f
C6383 _301_/a_240_7# _346_/SET_B 1.38e-20
C6384 _324_/Q _150_/a_27_7# 3.57e-19
C6385 output12/a_27_7# clk 2e-21
C6386 _290_/Y output38/a_27_7# 0.0306f
C6387 _281_/Y clkbuf_0_clk/a_110_7# 0.0332f
C6388 _263_/a_109_257# VGND -5.38e-19
C6389 ctln[3] _312_/a_193_7# 2.13e-19
C6390 _275_/Y _312_/a_543_7# 0.0104f
C6391 _298_/B _298_/C 0.195f
C6392 _283_/Y _335_/D 3.18e-19
C6393 _153_/B _203_/a_209_257# 1.52e-21
C6394 _182_/a_215_7# VPWR 0.00354f
C6395 _182_/a_79_n19# VGND 0.0373f
C6396 _267_/B _193_/Y 3.1e-20
C6397 _309_/D _340_/Q 4.17e-20
C6398 _183_/a_1241_257# _228_/A 3.15e-19
C6399 _324_/a_543_7# _181_/X 8.53e-21
C6400 _242_/A _331_/CLK 0.559f
C6401 _339_/a_651_373# _193_/Y 0.00357f
C6402 _312_/a_1462_7# VPWR 4.29e-19
C6403 _146_/C _286_/Y 0.0118f
C6404 _160_/X _299_/a_493_257# 6.54e-19
C6405 _335_/Q _190_/A 0.00604f
C6406 _204_/Y _333_/Q 0.295f
C6407 _319_/a_761_249# _319_/D 6.23e-19
C6408 _325_/Q _316_/D 0.371f
C6409 _304_/a_79_n19# _315_/D 3.17e-19
C6410 _300_/a_383_7# _347_/a_1108_7# 9.61e-21
C6411 _157_/A _286_/Y 0.00597f
C6412 _145_/A _250_/X 6.25e-19
C6413 _273_/A _242_/A 5.93e-19
C6414 input4/X _283_/A 1.63e-20
C6415 _181_/X _217_/A 0.296f
C6416 _286_/B _324_/D 2.71e-20
C6417 _246_/B _223_/a_93_n19# 0.0128f
C6418 _157_/A _297_/a_27_257# 5.14e-20
C6419 _326_/a_1108_7# _326_/Q 0.00439f
C6420 _287_/a_121_257# VPWR -5.08e-19
C6421 input1/X _260_/A 0.00648f
C6422 _339_/Q _267_/A 0.106f
C6423 _298_/A _204_/a_277_7# 5.95e-20
C6424 _322_/D _248_/A 1.18e-20
C6425 _293_/a_39_257# _254_/B 3.88e-19
C6426 _321_/a_448_7# _248_/A 7.62e-20
C6427 _279_/Y _314_/a_193_7# 0.0174f
C6428 _258_/a_218_334# _197_/X 6.44e-20
C6429 _342_/a_27_7# _342_/a_193_7# -4.92e-19
C6430 _283_/A _207_/C 0.314f
C6431 output15/a_27_7# _321_/Q 7.04e-19
C6432 _288_/A _309_/a_193_7# 1.73e-20
C6433 _322_/D _331_/CLK 0.108f
C6434 _236_/B _234_/B 0.0132f
C6435 _183_/a_1241_257# _216_/A 2.21e-19
C6436 _324_/Q _250_/a_78_159# 3.08e-21
C6437 _343_/a_193_7# valid 0.00235f
C6438 _167_/a_373_7# clkbuf_2_3_0_clk/A 4.21e-19
C6439 _321_/D _321_/a_761_249# 3.32e-20
C6440 _321_/a_448_7# _331_/CLK 0.0138f
C6441 _236_/B _321_/a_1283_n19# 4.43e-19
C6442 _320_/a_27_7# output18/a_27_7# 0.0105f
C6443 _346_/SET_B _310_/a_639_7# 0.00117f
C6444 _325_/a_1108_7# _216_/A 7.43e-20
C6445 _333_/a_1462_7# VPWR 7.25e-20
C6446 _333_/a_805_7# VGND 8.59e-20
C6447 input1/X _261_/A 1.96e-21
C6448 _342_/a_1108_7# _188_/S 1.83e-20
C6449 _242_/A _319_/a_1108_7# 0.0181f
C6450 _211_/a_27_257# _197_/X 0.0106f
C6451 _299_/a_215_7# VPWR -0.00103f
C6452 _299_/a_292_257# VGND -0.00102f
C6453 clk _251_/a_215_7# 0.00155f
C6454 result[0] _315_/a_1283_n19# 0.00389f
C6455 _343_/a_761_249# _343_/Q 2.72e-19
C6456 _337_/Q _194_/X 1.82f
C6457 clkbuf_0_clk/X _221_/a_250_257# 0.00818f
C6458 _197_/X _198_/a_93_n19# 0.0523f
C6459 _315_/D _347_/a_193_7# 0.00661f
C6460 _174_/a_109_257# _344_/D 4.53e-19
C6461 _336_/a_448_7# _340_/CLK 7.73e-19
C6462 result[2] _343_/CLK 3.45e-19
C6463 _255_/B _144_/A 0.0577f
C6464 _153_/a_487_257# _333_/Q 0.00114f
C6465 _277_/A _319_/a_193_7# 0.00154f
C6466 _308_/S _147_/Y 7.48e-21
C6467 _305_/a_76_159# _254_/B 0.0241f
C6468 _268_/a_39_257# VPWR 0.0531f
C6469 _232_/a_27_7# _241_/a_113_257# 8.91e-19
C6470 _317_/Q _304_/S 2.1e-20
C6471 _227_/A _334_/a_27_7# 2e-19
C6472 _346_/D _347_/a_1108_7# 4.47e-20
C6473 _316_/a_27_7# _245_/a_113_257# 1.54e-19
C6474 _283_/A _150_/C 0.0122f
C6475 _250_/a_215_7# _260_/A 0.00447f
C6476 _318_/Q _322_/a_193_7# 2.97e-21
C6477 _254_/Y _313_/a_1283_n19# 9.33e-21
C6478 _309_/a_1283_n19# _164_/Y 8.99e-19
C6479 _183_/a_471_7# _306_/S 0.00542f
C6480 _342_/a_193_7# _317_/D 3.04e-19
C6481 _275_/Y _263_/B 0.00707f
C6482 _214_/a_109_7# _331_/D 4.9e-19
C6483 _302_/a_227_7# _328_/Q 3.8e-20
C6484 _328_/a_1108_7# clkbuf_2_1_0_clk/A 4.92e-21
C6485 _343_/D _192_/B 0.00281f
C6486 output14/a_27_7# VGND 0.103f
C6487 _336_/Q _190_/A 0.133f
C6488 _206_/A _153_/a_109_53# 3.54e-19
C6489 _346_/SET_B _336_/a_651_373# 0.00399f
C6490 _316_/D _326_/Q 0.0121f
C6491 _182_/X VGND 0.521f
C6492 _279_/A _347_/a_543_7# 4.08e-20
C6493 _345_/a_1032_373# _165_/a_78_159# 2.86e-19
C6494 _255_/B _145_/A 0.11f
C6495 _339_/Q _194_/X 0.867f
C6496 _315_/a_1108_7# _248_/A 5.14e-19
C6497 _188_/a_505_n19# _298_/A 0.0214f
C6498 _312_/Q VGND 0.426f
C6499 _342_/a_543_7# _323_/D 0.00125f
C6500 _343_/CLK _153_/a_215_257# 2.56e-21
C6501 _319_/Q output26/a_27_7# 0.0416f
C6502 _317_/Q _317_/a_27_7# 0.00103f
C6503 _230_/a_27_7# _317_/a_761_249# 0.00388f
C6504 _248_/B _150_/C 1.21e-19
C6505 _271_/A _177_/A 0.215f
C6506 _340_/a_193_7# VPWR 0.0361f
C6507 _340_/Q _202_/a_250_257# 0.00113f
C6508 _306_/S _202_/a_93_n19# 8.39e-19
C6509 _320_/Q _321_/Q 0.0105f
C6510 _313_/D _306_/X 0.0046f
C6511 _304_/a_578_7# VGND -2.04e-19
C6512 _255_/X _192_/B 0.0324f
C6513 _165_/X clkbuf_0_clk/X 1.54e-19
C6514 _270_/a_39_257# _317_/a_1283_n19# 8.1e-19
C6515 repeater43/X _175_/Y 0.553f
C6516 _327_/a_27_7# _330_/Q 0.00282f
C6517 _283_/A _331_/a_1283_n19# 0.0172f
C6518 _316_/a_27_7# VPWR 0.0896f
C6519 _343_/a_27_7# _229_/a_489_373# 4.1e-20
C6520 _343_/a_193_7# _229_/a_226_7# 0.0105f
C6521 _343_/a_761_249# _229_/a_76_159# 5.81e-19
C6522 _344_/Q _284_/A 1.86e-20
C6523 _251_/a_79_n19# _286_/Y 0.0102f
C6524 _221_/a_250_257# _286_/Y 0.00299f
C6525 _248_/A _224_/a_346_7# 1.97e-19
C6526 cal _306_/S 0.618f
C6527 _237_/a_199_7# VGND -4.25e-19
C6528 input1/X _340_/Q 0.0964f
C6529 VGND valid 0.215f
C6530 _325_/Q _144_/A 0.00151f
C6531 output35/a_27_7# _284_/a_39_257# 0.0234f
C6532 _209_/a_27_257# _206_/A 2.29e-20
C6533 _326_/a_27_7# _330_/Q 7.22e-21
C6534 _326_/Q _222_/a_250_257# 0.00594f
C6535 _279_/Y _314_/a_1462_7# 9.2e-20
C6536 clkbuf_2_1_0_clk/A _338_/D 0.226f
C6537 clkbuf_2_0_0_clk/a_75_172# _338_/Q 0.0142f
C6538 _215_/A _340_/CLK 0.0177f
C6539 _317_/a_761_249# _232_/A 6.16e-20
C6540 _306_/X _197_/X 4.92e-22
C6541 _242_/A _217_/X 0.826f
C6542 _337_/a_543_7# _336_/Q 1.58e-21
C6543 _335_/D _333_/a_27_7# 3.77e-21
C6544 _197_/a_27_7# _306_/S 0.0405f
C6545 _165_/a_215_7# _160_/X 3.83e-19
C6546 _277_/Y _340_/CLK 0.43f
C6547 _320_/Q _297_/B 0.0206f
C6548 _237_/a_113_257# _314_/Q 6.93e-20
C6549 _279_/Y _324_/D 2.09e-20
C6550 _324_/Q _250_/X 0.00832f
C6551 _250_/a_78_159# _216_/A 0.0537f
C6552 _342_/Q _149_/a_27_7# 0.00707f
C6553 _338_/Q _310_/D 4.74e-19
C6554 output14/a_27_7# output27/a_27_7# 1.26e-20
C6555 _283_/Y _312_/a_448_7# 9.57e-21
C6556 _157_/A _328_/Q 0.00183f
C6557 _327_/a_651_373# _217_/A 3.65e-20
C6558 clkbuf_0_clk/X _251_/X 0.0673f
C6559 _315_/Q _315_/D 6.54e-20
C6560 output12/a_27_7# _281_/Y 0.0486f
C6561 _329_/a_1283_n19# clkbuf_0_clk/X 0.0176f
C6562 _300_/a_383_7# _346_/SET_B 0.00548f
C6563 output22/a_27_7# VPWR 0.114f
C6564 _332_/a_1108_7# VGND 0.00504f
C6565 _332_/a_651_373# VPWR -0.00288f
C6566 _331_/Q _214_/a_27_257# 0.0112f
C6567 _347_/a_448_7# VGND -0.00288f
C6568 _347_/a_1270_373# VPWR -2.05e-19
C6569 _200_/a_256_7# VPWR -6.86e-19
C6570 _285_/A _288_/A 1.74f
C6571 _200_/a_93_n19# VGND 0.00237f
C6572 _277_/A _319_/a_1462_7# 2.64e-19
C6573 input3/a_27_7# _206_/A 0.00116f
C6574 repeater43/X _321_/a_805_7# -7.69e-19
C6575 _319_/Q _281_/A 0.0367f
C6576 _328_/a_27_7# _297_/B 0.00677f
C6577 _314_/Q _347_/a_1108_7# 9.86e-21
C6578 _314_/D _347_/a_639_7# 1.49e-20
C6579 _285_/A _162_/X 0.0203f
C6580 _267_/B _310_/a_1270_373# 1.37e-19
C6581 _279_/Y _279_/A 0.0136f
C6582 _306_/a_439_7# _286_/B 2.74e-19
C6583 _258_/S _311_/a_1108_7# 5.11e-20
C6584 _288_/A _344_/a_193_7# 2.17e-20
C6585 _346_/a_476_7# _299_/X 0.00794f
C6586 _346_/a_652_n19# _347_/Q 7.8e-21
C6587 _304_/X _347_/D 0.00131f
C6588 _251_/a_297_257# _284_/A 2.88e-19
C6589 _343_/CLK _315_/a_543_7# 0.0301f
C6590 _294_/A cal 4.98e-19
C6591 _175_/Y _191_/B 1.18e-21
C6592 _216_/X _218_/a_584_7# 7.13e-19
C6593 result[3] _317_/D 0.00271f
C6594 clkbuf_2_3_0_clk/a_75_172# clkbuf_2_3_0_clk/A 0.0159f
C6595 _313_/D _147_/Y 3.21e-20
C6596 ctln[4] _338_/D 5.35e-20
C6597 _165_/a_493_257# VGND -7.55e-20
C6598 _327_/a_1108_7# _279_/A 2.19e-19
C6599 _344_/a_193_7# _162_/X 1.81e-19
C6600 _183_/a_471_7# _283_/A 0.00648f
C6601 _239_/a_113_257# _240_/B 0.0102f
C6602 _345_/a_27_7# _173_/a_76_159# 1.37e-19
C6603 _304_/S _298_/A 0.00247f
C6604 _254_/A _336_/a_1283_n19# 8.61e-19
C6605 _341_/a_1270_373# VGND 3.71e-20
C6606 _336_/a_761_249# _157_/a_27_7# 9.26e-21
C6607 _341_/a_805_7# VPWR 2.79e-19
C6608 _188_/a_505_n19# _215_/A 6.01e-20
C6609 _179_/a_27_7# _333_/a_1283_n19# 5.13e-20
C6610 _197_/X _147_/Y 8.41e-19
C6611 _258_/S _275_/Y 0.506f
C6612 _338_/a_805_7# VPWR 1.55e-19
C6613 _338_/a_1270_373# VGND 6.82e-20
C6614 _323_/a_193_7# _176_/a_27_7# 8.17e-19
C6615 _331_/D _330_/a_761_249# 4.39e-20
C6616 _274_/a_121_257# _315_/D 1.71e-19
C6617 _206_/A _153_/A 0.0127f
C6618 _165_/X _286_/Y 0.162f
C6619 clkbuf_2_3_0_clk/a_75_172# _172_/Y 3.7e-19
C6620 _330_/a_193_7# _330_/a_761_249# -0.00517f
C6621 _275_/A trimb[3] 4.22e-20
C6622 _316_/Q _316_/a_543_7# 0.0416f
C6623 _172_/A _162_/X 0.0325f
C6624 _286_/B _153_/B 5.25e-20
C6625 ctlp[4] ctlp[5] 0.00198f
C6626 clkbuf_2_1_0_clk/A _313_/a_193_7# 1.21e-20
C6627 _325_/a_543_7# _325_/Q 3.39e-20
C6628 _328_/a_1283_n19# _279_/A 2.81e-20
C6629 _346_/SET_B _314_/a_805_7# -0.00125f
C6630 _186_/a_79_n19# _177_/A 2.94e-19
C6631 repeater43/X _341_/Q -0.0014f
C6632 _250_/X _228_/A 0.0065f
C6633 _225_/X _298_/A 0.00583f
C6634 _307_/X _298_/A 0.0517f
C6635 _236_/B _235_/a_113_257# 0.00667f
C6636 _235_/a_199_7# _316_/D 5.98e-19
C6637 _324_/Q _247_/a_199_7# 0.00201f
C6638 _229_/a_226_7# VGND -0.0119f
C6639 _229_/a_226_257# VPWR -1.28e-19
C6640 _346_/SET_B _217_/A 8.35e-19
C6641 _336_/a_651_373# _147_/A 3.65e-19
C6642 _295_/a_79_n19# VPWR -0.00267f
C6643 clkbuf_2_1_0_clk/A _343_/CLK 0.00262f
C6644 _346_/a_27_7# VPWR 0.0645f
C6645 _337_/Q _310_/a_1108_7# 0.0043f
C6646 _300_/Y _347_/D 4.71e-20
C6647 _340_/a_1462_7# VPWR 7.03e-20
C6648 _194_/X _336_/D 2.33e-19
C6649 _340_/a_805_7# VGND 2.92e-19
C6650 _346_/SET_B _346_/D 0.0972f
C6651 _306_/S _284_/A 0.663f
C6652 _144_/A _326_/Q 1.88e-20
C6653 cal _283_/A 0.0509f
C6654 _335_/a_27_7# _208_/a_78_159# 0.00133f
C6655 _239_/a_113_257# _328_/Q 0.011f
C6656 _345_/a_1182_221# _346_/SET_B -1.39e-21
C6657 _316_/a_639_7# VGND -0.00141f
C6658 _316_/a_1217_7# VPWR 6.88e-20
C6659 _343_/a_1108_7# _248_/A 4.11e-19
C6660 _344_/a_1182_221# _164_/Y 0.0122f
C6661 _300_/a_383_7# _313_/a_761_249# 3.48e-20
C6662 _346_/a_652_n19# _297_/B 3.53e-20
C6663 _293_/a_121_257# _286_/B 1.2e-19
C6664 _331_/a_27_7# _326_/Q 1.15e-20
C6665 _251_/X _286_/Y 6.51e-20
C6666 _255_/X _157_/A 9.79e-21
C6667 _204_/a_277_7# VGND -0.00392f
C6668 _255_/B _324_/Q 0.15f
C6669 _338_/Q _266_/a_113_257# 7.1e-21
C6670 _296_/a_213_83# _286_/Y 0.00103f
C6671 _327_/a_805_7# VPWR 3.7e-19
C6672 _342_/a_448_7# _342_/D 0.0275f
C6673 _273_/A _324_/a_448_7# 5.57e-19
C6674 _341_/Q _334_/Q 2.15e-19
C6675 repeater43/X _315_/a_639_7# 0.00195f
C6676 _216_/A _250_/X 0.00257f
C6677 _195_/a_373_7# _193_/Y 8.02e-19
C6678 _326_/a_1270_373# VGND 7.49e-20
C6679 _215_/A _313_/a_543_7# 0.0296f
C6680 _312_/a_193_7# _312_/a_1108_7# -3.36e-19
C6681 output33/a_27_7# trim[2] 0.00874f
C6682 _283_/Y _312_/D 7.92e-20
C6683 _251_/a_510_7# _250_/X 8.53e-19
C6684 _149_/A _153_/A 1.96e-20
C6685 _180_/a_29_13# VPWR 0.0306f
C6686 _332_/a_761_249# _153_/B 0.00426f
C6687 _330_/Q _319_/a_193_7# 1.65e-20
C6688 _324_/a_1108_7# _222_/a_250_257# 1.99e-21
C6689 _301_/X _301_/a_149_7# 0.00115f
C6690 _340_/CLK VGND 2.88f
C6691 _328_/a_639_7# VPWR 5.25e-19
C6692 _328_/a_651_373# VGND 0.00139f
C6693 _347_/D VGND 0.19f
C6694 _254_/Y _202_/a_93_n19# 1.26e-20
C6695 _221_/a_250_257# _328_/Q 0.0581f
C6696 _331_/Q _330_/a_27_7# 2.29e-19
C6697 _217_/a_27_7# _326_/Q 0.00157f
C6698 _341_/Q _191_/B 0.00131f
C6699 _258_/a_76_159# _194_/A 5.17e-21
C6700 ctln[4] _343_/CLK 0.0323f
C6701 _318_/Q _331_/Q 0.0668f
C6702 _181_/X _214_/a_109_257# 0.00936f
C6703 _305_/a_505_n19# _286_/B 0.0415f
C6704 _294_/A _284_/A 0.119f
C6705 _271_/Y _334_/a_193_7# 1.72e-20
C6706 _271_/A _334_/a_543_7# 0.0311f
C6707 _319_/a_27_7# VPWR 0.0627f
C6708 _328_/a_1217_7# _297_/B 1.58e-20
C6709 _297_/B _173_/a_226_7# 3.93e-19
C6710 _321_/a_639_7# result[7] 1.47e-19
C6711 _215_/A _304_/S 1.68e-20
C6712 _300_/a_383_7# _147_/A 4.43e-19
C6713 _254_/Y cal 2.32e-20
C6714 _309_/D _310_/D 7.16e-19
C6715 _337_/Q _336_/a_543_7# 0.00129f
C6716 _298_/B _150_/C 0.584f
C6717 _258_/S _258_/a_76_159# 0.0396f
C6718 _319_/a_761_249# _297_/B 2.87e-19
C6719 _255_/X _260_/A 8.38e-20
C6720 _290_/A _290_/Y 0.0122f
C6721 _334_/a_639_7# VPWR 7.25e-19
C6722 _334_/a_651_373# VGND 0.0014f
C6723 _254_/Y _197_/a_27_7# 1.87e-21
C6724 _257_/a_448_7# _260_/A 0.00363f
C6725 clkbuf_0_clk/a_110_7# _336_/Q 6.22e-20
C6726 _218_/a_256_7# _331_/CLK 5.59e-19
C6727 _309_/a_761_249# _340_/CLK 3.33e-20
C6728 _329_/Q _320_/a_27_7# 1.14e-20
C6729 _320_/Q _320_/a_193_7# 7.57e-19
C6730 _345_/a_193_7# _345_/D 0.0868f
C6731 _345_/a_652_n19# _345_/Q 7e-19
C6732 _343_/a_543_7# _343_/CLK 2.91e-20
C6733 _325_/a_543_7# _326_/Q 0.00584f
C6734 _232_/A _286_/Y 1.97e-22
C6735 _324_/a_761_249# _304_/S 0.022f
C6736 _283_/Y _332_/a_193_7# 3.61e-20
C6737 _273_/A _218_/a_256_7# 3.48e-21
C6738 _255_/B _228_/A 0.021f
C6739 _338_/Q VPWR 1.18f
C6740 _227_/A _323_/Q 0.00298f
C6741 clkbuf_2_3_0_clk/A _299_/X 0.00509f
C6742 _275_/A VPWR 2.59f
C6743 _271_/A _248_/A 0.0143f
C6744 _325_/Q _324_/Q 0.0652f
C6745 _329_/a_639_7# _281_/A 0.00462f
C6746 _277_/Y _267_/B 0.00883f
C6747 _183_/a_27_7# _298_/A 0.00384f
C6748 _346_/SET_B _314_/Q 0.124f
C6749 _304_/S _304_/X 0.274f
C6750 _340_/a_193_7# _198_/a_93_n19# 6.25e-19
C6751 _340_/a_27_7# _198_/a_250_257# 4.93e-20
C6752 _283_/A _284_/A 1.86e-20
C6753 _342_/a_651_373# _177_/a_27_7# 8.8e-20
C6754 _342_/a_543_7# _177_/A 1.16e-19
C6755 _271_/A _331_/CLK 0.00942f
C6756 _188_/a_505_n19# VGND 0.0682f
C6757 _188_/a_535_334# VPWR -7.21e-19
C6758 _342_/a_193_7# _298_/X 2.51e-21
C6759 _346_/a_956_373# VGND 8.77e-19
C6760 _299_/X _172_/Y 1.48e-20
C6761 _160_/X _345_/Q 0.891f
C6762 _333_/a_27_7# _333_/a_448_7# -0.00972f
C6763 _172_/A _298_/C 0.0066f
C6764 _335_/a_761_249# _332_/Q 3.56e-21
C6765 _279_/Y _153_/B 2.82e-19
C6766 _309_/a_543_7# _346_/SET_B 0.0073f
C6767 _335_/a_543_7# _207_/X 8.34e-19
C6768 _343_/a_193_7# _225_/X 3.77e-20
C6769 _343_/a_761_249# _147_/A 7e-22
C6770 _342_/a_27_7# _343_/Q 1.31e-21
C6771 _321_/D VGND 0.337f
C6772 _329_/a_651_373# _319_/Q 0.0266f
C6773 _273_/A _271_/A 9.17e-21
C6774 _347_/Q _313_/a_651_373# 7.17e-21
C6775 _339_/Q _336_/a_543_7# 5.16e-19
C6776 _317_/a_193_7# _242_/B 1.55e-20
C6777 _162_/a_27_7# _310_/D 3.27e-20
C6778 _265_/B _174_/a_109_257# 8.14e-19
C6779 _319_/Q _240_/a_109_257# 4.52e-19
C6780 _328_/a_1108_7# _328_/D 5.47e-21
C6781 _147_/A _346_/D 2.4e-21
C6782 _158_/Y _297_/B 7.51e-21
C6783 _255_/B _216_/A 3.38e-19
C6784 _335_/D _298_/C 1.44e-20
C6785 _200_/a_346_7# _311_/D 6.57e-20
C6786 _329_/a_448_7# _329_/D 0.0145f
C6787 repeater43/X _330_/Q 0.0814f
C6788 _283_/Y _338_/a_1283_n19# 0.00529f
C6789 _321_/D _318_/a_1108_7# 6.03e-20
C6790 _326_/a_1283_n19# _232_/a_27_7# 1.49e-20
C6791 _263_/B _312_/a_543_7# 1.89e-21
C6792 _336_/a_1283_n19# _202_/a_250_257# 6.76e-20
C6793 _235_/a_113_257# _331_/a_193_7# 1.7e-19
C6794 _248_/B _284_/A 5.13e-20
C6795 _342_/Q _251_/a_297_257# 0.00262f
C6796 _143_/a_181_7# VGND 1.6e-19
C6797 _294_/A trim[2] 0.00223f
C6798 _294_/Y _290_/A 4.01e-19
C6799 input4/X ctln[0] 1.81e-20
C6800 repeater43/X _269_/Y 3.9e-19
C6801 _312_/a_27_7# _312_/D 0.0548f
C6802 _347_/Q _157_/a_27_7# 0.0115f
C6803 _300_/Y _156_/a_121_257# 1.74e-21
C6804 repeater43/X _324_/a_805_7# -0.00125f
C6805 input1/X _336_/a_1283_n19# 0.0602f
C6806 _315_/D _212_/X 0.004f
C6807 _300_/Y _304_/S 5.84e-20
C6808 _275_/Y _173_/a_226_7# 2.39e-20
C6809 _222_/a_584_7# VGND -8.39e-19
C6810 output23/a_27_7# _343_/CLK 1.36e-19
C6811 _336_/a_193_7# _260_/A 2.24e-20
C6812 repeater43/X _318_/a_761_249# 0.0191f
C6813 _343_/a_639_7# repeater43/X 7.5e-19
C6814 _345_/D VPWR 0.271f
C6815 _329_/a_193_7# _329_/a_1283_n19# -5.93e-19
C6816 _251_/X _328_/Q 7.18e-20
C6817 _254_/Y _284_/A 0.0106f
C6818 _329_/a_27_7# _327_/D 1.8e-20
C6819 _291_/a_121_257# _339_/Q 0.001f
C6820 _306_/a_76_159# _338_/Q 3.62e-20
C6821 _181_/X _331_/D 0.00458f
C6822 _318_/a_27_7# _327_/Q 3.12e-21
C6823 _319_/a_1217_7# VPWR 6.22e-20
C6824 _319_/a_639_7# VGND 0.00458f
C6825 _313_/a_1108_7# VPWR -0.00143f
C6826 _313_/a_543_7# VGND 0.0169f
C6827 _323_/a_27_7# _248_/A 1.47e-19
C6828 _283_/Y _208_/a_78_159# 2.95e-21
C6829 _337_/a_639_7# VPWR 3.31e-19
C6830 _337_/a_651_373# VGND 0.00108f
C6831 _346_/SET_B _311_/a_805_7# 5.85e-19
C6832 _183_/a_471_7# _298_/B 8.45e-19
C6833 _321_/D output27/a_27_7# 5.94e-19
C6834 _342_/a_651_373# _341_/a_27_7# 2.28e-20
C6835 _298_/C _203_/a_80_n19# 0.0266f
C6836 _343_/Q _254_/B 9.52e-20
C6837 _297_/B _313_/a_651_373# 4.76e-20
C6838 _231_/a_79_n19# _177_/A 3.64e-19
C6839 output21/a_27_7# _322_/Q 7.76e-19
C6840 _344_/a_1602_7# _160_/A 0.0116f
C6841 _320_/Q _322_/a_1108_7# 0.0532f
C6842 _321_/a_1108_7# _281_/A 7.21e-21
C6843 _330_/D _331_/CLK 0.179f
C6844 _342_/Q _306_/S 0.0199f
C6845 _197_/X _338_/a_543_7# 4.98e-21
C6846 _276_/a_68_257# clkbuf_2_1_0_clk/A 5.28e-19
C6847 _282_/a_39_257# _246_/B 9.15e-19
C6848 _238_/a_109_257# _238_/B 0.00285f
C6849 _307_/a_439_7# VGND -3.52e-19
C6850 _254_/A VPWR 0.858f
C6851 _324_/Q _326_/Q 0.00205f
C6852 _156_/a_121_257# VGND -4.61e-19
C6853 _267_/A _260_/a_27_257# 0.0171f
C6854 clk _215_/A 0.0521f
C6855 _308_/X _229_/a_76_159# 2.74e-21
C6856 _304_/S VGND 1.71f
C6857 input4/a_27_7# _306_/S 2.41e-19
C6858 _342_/a_27_7# _229_/a_76_159# 8.42e-19
C6859 _323_/D _298_/C 6.91e-19
C6860 ctln[6] rstn 0.0115f
C6861 _297_/B _157_/a_27_7# 1.75e-19
C6862 _313_/D _260_/B 0.00231f
C6863 _297_/A _162_/X 1.05e-19
C6864 _319_/Q _321_/a_543_7# 3.1e-19
C6865 _325_/Q _216_/A 0.182f
C6866 _232_/a_27_7# _248_/A 0.0598f
C6867 _288_/A _164_/A 1.22e-20
C6868 _218_/a_93_n19# _331_/a_193_7# 9.26e-20
C6869 _340_/a_1108_7# _197_/X 0.0352f
C6870 _298_/B cal 0.162f
C6871 _218_/a_256_7# _217_/X 3.61e-20
C6872 _325_/a_193_7# _315_/D 1.82e-21
C6873 _225_/X VGND 0.0553f
C6874 _246_/B _327_/Q 0.00641f
C6875 _226_/X VPWR 0.276f
C6876 _164_/A _162_/X 0.203f
C6877 _307_/X VGND 0.0954f
C6878 _275_/Y _158_/Y 1.2e-21
C6879 _232_/a_27_7# _331_/CLK 7.28e-23
C6880 _324_/a_27_7# clkbuf_0_clk/X 0.00542f
C6881 cal _194_/a_27_7# 1.38e-20
C6882 _325_/a_543_7# _324_/a_1108_7# 5.1e-20
C6883 _285_/A output35/a_27_7# 0.00829f
C6884 ctln[7] _334_/a_193_7# 6.27e-21
C6885 _283_/Y _334_/a_543_7# 3.56e-22
C6886 _157_/A _314_/a_1283_n19# 0.00339f
C6887 _320_/a_193_7# _319_/a_761_249# 8.57e-22
C6888 _320_/a_761_249# _319_/a_193_7# 1.3e-21
C6889 _333_/a_27_7# _333_/D 0.191f
C6890 _255_/a_184_257# _255_/X 7.52e-20
C6891 _314_/Q _147_/A 3.65e-19
C6892 clkbuf_0_clk/X _314_/a_651_373# 8.59e-19
C6893 result[1] repeater43/X 0.00472f
C6894 _267_/B VGND 0.231f
C6895 _309_/D VPWR 0.339f
C6896 _339_/a_639_7# VPWR 5.14e-19
C6897 _339_/a_651_373# VGND 5.86e-19
C6898 _217_/X _220_/a_584_7# 0.00138f
C6899 _341_/a_651_373# _317_/D 5.47e-19
C6900 _183_/a_1241_257# _217_/A 1.96e-19
C6901 _327_/a_639_7# _232_/X 5.86e-19
C6902 _163_/a_78_159# _171_/a_78_159# 5.04e-19
C6903 _265_/B _344_/D 8.85e-19
C6904 _199_/a_346_7# _267_/A 6.34e-20
C6905 _298_/B _150_/a_193_257# 4.47e-19
C6906 _325_/a_448_7# _304_/X 0.025f
C6907 _325_/a_1108_7# _217_/A 3.5e-19
C6908 _325_/a_543_7# _324_/D 6.44e-21
C6909 output5/a_27_7# _297_/Y 0.0185f
C6910 _317_/a_27_7# VGND -0.0716f
C6911 _317_/a_761_249# VPWR 0.0185f
C6912 _301_/X _215_/A 4.53e-21
C6913 _182_/a_79_n19# _286_/B 0.0676f
C6914 _326_/a_639_7# _232_/X 3.56e-19
C6915 repeater43/X _335_/a_1283_n19# 0.0328f
C6916 _252_/a_27_7# _347_/a_27_7# 9.11e-21
C6917 _277_/Y _301_/X 2.09e-20
C6918 _336_/a_543_7# _336_/D 2.27e-19
C6919 _336_/a_1108_7# _284_/A 0.0119f
C6920 _330_/Q _331_/a_448_7# 0.00449f
C6921 _258_/S _312_/a_543_7# 6.05e-21
C6922 _321_/Q result[7] 0.00806f
C6923 _271_/A _217_/X 1.12e-20
C6924 _292_/A _312_/a_27_7# 3e-19
C6925 trim[0] _346_/SET_B 1.33e-19
C6926 _211_/a_109_257# _332_/D 0.00255f
C6927 _312_/a_651_373# _312_/Q 1.47e-19
C6928 _188_/S _180_/a_111_257# 4.18e-19
C6929 _308_/S _307_/a_76_159# 0.00118f
C6930 _229_/a_76_159# _317_/D 5.76e-20
C6931 _229_/a_489_373# _244_/B 7.31e-20
C6932 _309_/a_27_7# _309_/D 0.147f
C6933 _309_/a_761_249# _267_/B 5.82e-19
C6934 _340_/a_193_7# _147_/Y 6.57e-22
C6935 _331_/a_1108_7# VPWR 0.0147f
C6936 _331_/a_543_7# VGND 0.0174f
C6937 _320_/a_448_7# _346_/SET_B 0.00329f
C6938 _290_/Y output36/a_27_7# 4.44e-19
C6939 _302_/a_227_257# VPWR 4.35e-19
C6940 _169_/B _168_/a_397_257# 2.33e-19
C6941 _294_/Y _310_/a_27_7# 3.94e-21
C6942 _254_/A _306_/a_76_159# 1.07e-20
C6943 _269_/A _232_/A 2.92e-21
C6944 _344_/a_476_7# _346_/SET_B 0.013f
C6945 _343_/a_27_7# cal 0.00961f
C6946 _308_/a_505_n19# _192_/B 7.38e-19
C6947 _336_/a_761_249# _194_/X 7.24e-20
C6948 _336_/a_27_7# _306_/S 0.0126f
C6949 _336_/a_193_7# _340_/Q 1.1e-20
C6950 _254_/B _204_/a_27_7# 1.42e-19
C6951 _302_/a_539_257# _297_/B 0.00404f
C6952 _260_/A _314_/a_1283_n19# 3.16e-19
C6953 _294_/A _264_/a_113_257# 6.31e-20
C6954 _157_/A _299_/X 0.0553f
C6955 _304_/a_257_159# _162_/X 7.4e-20
C6956 ctln[1] _271_/Y 0.223f
C6957 ctln[7] _332_/Q 0.00865f
C6958 _283_/Y _190_/A 1.12e-20
C6959 _346_/SET_B _311_/Q 2.51e-19
C6960 _258_/a_439_7# _346_/SET_B 8.96e-19
C6961 _335_/a_1283_n19# _334_/Q 0.0099f
C6962 _322_/a_761_249# _331_/CLK 9.01e-21
C6963 _325_/a_27_7# _246_/B 2.22e-20
C6964 _342_/D _341_/a_193_7# 5.98e-21
C6965 _342_/Q _283_/A 0.00818f
C6966 ctln[1] _335_/a_761_249# 6.55e-20
C6967 _321_/a_27_7# _269_/A 4.64e-19
C6968 _162_/X _177_/A 0.00173f
C6969 _169_/B _216_/A 8.1e-20
C6970 _162_/a_27_7# VPWR 0.117f
C6971 _144_/a_27_7# _283_/A 2.45e-19
C6972 _344_/a_1032_373# _163_/a_215_7# 8.34e-19
C6973 _314_/a_193_7# _228_/A 5.13e-20
C6974 rstn _269_/A 0.00239f
C6975 _271_/A _146_/a_29_271# 0.00629f
C6976 _346_/SET_B _198_/a_346_7# 0.00109f
C6977 _216_/A _326_/Q 0.167f
C6978 _250_/a_292_257# _215_/A 5.15e-20
C6979 _317_/a_1108_7# _246_/B 1.07e-20
C6980 _306_/a_76_159# _309_/D 4.58e-20
C6981 _188_/a_76_159# _308_/X 1.99e-21
C6982 _324_/a_27_7# _286_/Y 0.0114f
C6983 _320_/Q _330_/a_651_373# 0.0262f
C6984 _342_/a_543_7# _248_/A 0.0107f
C6985 _252_/a_27_7# _216_/X 0.0112f
C6986 _344_/a_1602_7# _273_/A 0.00398f
C6987 _284_/a_39_257# _284_/A 0.0257f
C6988 _346_/Q _170_/a_76_159# 0.0127f
C6989 result[6] _318_/a_761_249# 3.41e-20
C6990 repeater43/X _323_/a_1283_n19# -4.49e-19
C6991 _342_/Q _248_/B 5.23e-20
C6992 _184_/a_218_7# _147_/A 0.0013f
C6993 _184_/a_218_334# _150_/C 2.58e-20
C6994 _184_/a_505_n19# _226_/X 2.53e-20
C6995 _194_/a_27_7# _284_/A 1.15e-20
C6996 clkbuf_2_1_0_clk/A _344_/D 1.3e-20
C6997 _285_/A _345_/Q 0.00101f
C6998 _144_/a_27_7# _248_/B 0.0403f
C6999 _294_/A _336_/a_27_7# 2e-21
C7000 _183_/a_27_7# VGND 0.0394f
C7001 _199_/a_93_n19# _193_/Y 0.0353f
C7002 _330_/D _217_/X 0.00326f
C7003 _324_/a_1108_7# _324_/Q 0.00346f
C7004 clkbuf_0_clk/X VPWR 2.08f
C7005 _301_/X _300_/Y 0.0282f
C7006 clk VGND 0.494f
C7007 _325_/a_448_7# VGND -0.00395f
C7008 _346_/Q clkbuf_2_1_0_clk/A 0.0105f
C7009 _299_/X _260_/A 7.1e-20
C7010 _263_/B _194_/A 1.4e-19
C7011 _219_/a_93_n19# _278_/a_68_257# 1.51e-20
C7012 _344_/a_27_7# _345_/D 0.00105f
C7013 _344_/a_193_7# _345_/Q 5.83e-20
C7014 _216_/A _314_/a_193_7# 2.28e-20
C7015 _257_/a_544_257# _254_/Y 0.00114f
C7016 _324_/Q _324_/D 0.598f
C7017 _168_/a_481_7# clkbuf_2_1_0_clk/A 9.45e-19
C7018 _216_/A _224_/a_256_7# 0.00266f
C7019 _169_/Y _306_/S 9.2e-20
C7020 _163_/a_78_159# _172_/B 0.00257f
C7021 _193_/Y _336_/Q 0.68f
C7022 _258_/S _263_/B 0.0387f
C7023 _306_/S _225_/B 0.334f
C7024 _346_/SET_B _254_/B 0.0196f
C7025 clkbuf_1_1_0_clk/a_75_172# _319_/D 6.23e-20
C7026 ctlp[6] clkbuf_0_clk/X 0.07f
C7027 _323_/a_639_7# _343_/CLK 4.14e-19
C7028 _286_/B _182_/X 6.23e-19
C7029 _196_/A _181_/X 0.043f
C7030 _202_/a_250_257# VPWR 0.0394f
C7031 input4/X _335_/D 4.89e-19
C7032 _283_/A _204_/Y 0.00121f
C7033 _297_/A _347_/a_651_373# 9.07e-20
C7034 _172_/A _345_/Q 0.00444f
C7035 _288_/Y _285_/Y 0.0338f
C7036 _347_/Q _267_/A 8.06e-21
C7037 _324_/a_193_7# _284_/A 2.45e-21
C7038 _337_/Q _311_/a_448_7# 2.09e-20
C7039 _290_/Y output39/a_27_7# 6.45e-19
C7040 _317_/Q _242_/A 7.36e-20
C7041 _341_/a_761_249# _177_/a_27_7# 4.33e-19
C7042 _281_/Y _215_/A 0.144f
C7043 output10/a_27_7# _194_/X 3.63e-21
C7044 ctln[4] _195_/a_109_257# 2.14e-19
C7045 _232_/a_27_7# _217_/X 2.04e-20
C7046 _172_/A _313_/a_1283_n19# 3.27e-20
C7047 _344_/a_27_7# _254_/A 5.65e-21
C7048 _205_/a_382_257# _204_/Y 3.25e-19
C7049 _205_/a_297_7# _335_/Q 0.0334f
C7050 input1/X VPWR 3.15f
C7051 _288_/A _292_/A 0.0203f
C7052 _323_/a_543_7# _323_/Q 9.4e-19
C7053 _323_/a_1283_n19# _191_/B 0.0011f
C7054 repeater43/X _212_/a_27_7# 9.04e-20
C7055 _301_/X VGND 0.316f
C7056 _256_/a_303_7# _181_/X 1.43e-19
C7057 _292_/A _162_/X 0.382f
C7058 _331_/D _346_/SET_B 0.00148f
C7059 _335_/D _207_/C 0.0106f
C7060 _162_/A trimb[4] 0.0931f
C7061 _288_/A _160_/A 0.00775f
C7062 _292_/A _287_/a_39_257# 0.00748f
C7063 _197_/X _337_/a_761_249# 9e-19
C7064 _343_/a_1217_7# cal 5.25e-20
C7065 _189_/a_27_7# _209_/a_27_257# 4.12e-20
C7066 _258_/a_76_159# _157_/a_27_7# 3.62e-21
C7067 _342_/a_193_7# _343_/CLK 0.00334f
C7068 _254_/Y _264_/a_113_257# 3.16e-19
C7069 _277_/Y _166_/Y 0.00563f
C7070 _280_/a_68_257# VGND 0.0151f
C7071 _158_/Y _161_/Y 0.0465f
C7072 _283_/Y _339_/a_543_7# 6.04e-22
C7073 _162_/X _160_/A 0.0103f
C7074 _255_/B _209_/a_27_257# 2.05e-19
C7075 _281_/Y _324_/a_761_249# 0.00121f
C7076 _150_/a_109_257# VGND -2.69e-19
C7077 _174_/a_373_7# VGND -0.00129f
C7078 _266_/a_199_7# _284_/A 0.00114f
C7079 _196_/A _343_/Q 3.25e-21
C7080 _322_/a_639_7# _321_/D 2.61e-19
C7081 _294_/A _169_/Y 5.06e-20
C7082 _185_/A _298_/A 4.53e-21
C7083 _273_/A _312_/a_27_7# 1.75e-21
C7084 _248_/A _330_/a_1283_n19# 5.88e-19
C7085 _324_/a_1108_7# _228_/A 3.26e-19
C7086 _319_/Q _318_/D 6.44e-20
C7087 _261_/a_109_257# VGND -0.00128f
C7088 output20/a_27_7# _281_/A 0.0284f
C7089 _281_/Y _304_/X 0.924f
C7090 _331_/CLK _330_/a_1283_n19# 7.89e-19
C7091 VPWR _286_/Y 0.884f
C7092 _297_/B _267_/A 1.61e-20
C7093 _308_/X _147_/A 0.174f
C7094 _172_/A _150_/C 0.0144f
C7095 _318_/Q _321_/D 0.00598f
C7096 _324_/a_1217_7# _286_/Y 1.59e-19
C7097 _297_/a_27_257# VPWR 0.127f
C7098 _228_/A _324_/D 0.0269f
C7099 _188_/S _191_/B 0.00425f
C7100 _219_/a_256_7# VGND -4.66e-19
C7101 _219_/a_584_7# VPWR -2.31e-19
C7102 repeater43/X _322_/a_448_7# 7.3e-22
C7103 _342_/Q _315_/a_27_7# 0.00869f
C7104 _206_/A _203_/a_209_7# 0.00182f
C7105 _343_/Q _298_/X 0.436f
C7106 _308_/X _149_/A 1.18e-19
C7107 _254_/B _206_/A 0.0104f
C7108 _319_/Q _217_/A 9.64e-20
C7109 _319_/Q _346_/D 4.53e-21
C7110 _333_/a_761_249# _332_/Q 8e-20
C7111 _333_/a_27_7# _190_/A 0.0218f
C7112 _333_/a_193_7# _333_/Q 9.11e-19
C7113 _254_/Y _336_/a_27_7# 0.0265f
C7114 _345_/a_476_7# _166_/Y 1.42e-19
C7115 _341_/a_27_7# _341_/a_761_249# -0.0166f
C7116 _320_/Q output15/a_27_7# 1.33e-19
C7117 _329_/D _304_/X 1.33e-19
C7118 _214_/a_27_257# _331_/a_543_7# 5.74e-19
C7119 _250_/a_215_7# VPWR 0.00105f
C7120 _250_/a_292_257# VGND -0.00119f
C7121 _324_/a_1108_7# _216_/A 6.83e-19
C7122 _334_/D _254_/B 4.3e-20
C7123 _333_/D _298_/C 0.0329f
C7124 _197_/X _339_/a_761_249# 4.4e-19
C7125 _258_/S _194_/A 2.68e-20
C7126 _218_/a_250_257# _281_/A 3.39e-19
C7127 _283_/A _225_/B 6.63e-21
C7128 _338_/a_27_7# _338_/a_761_249# -0.0166f
C7129 result[4] _318_/a_761_249# 2.84e-19
C7130 ctln[1] ctln[7] 0.0103f
C7131 _324_/a_27_7# _328_/Q 2.75e-19
C7132 _277_/A _319_/D 2e-19
C7133 _227_/A _296_/a_109_7# 0.00103f
C7134 _189_/a_27_7# _153_/A 1.18e-19
C7135 _216_/A _324_/D 6.56e-19
C7136 _342_/a_651_373# repeater43/X 5.73e-19
C7137 _297_/B _221_/a_93_n19# 9.48e-21
C7138 _255_/B _153_/A 0.00313f
C7139 _192_/B _154_/a_27_7# 2.15e-20
C7140 _340_/a_543_7# _194_/A 1.45e-20
C7141 _281_/Y _220_/a_93_n19# 3.6e-21
C7142 _166_/Y _300_/Y 5.37e-20
C7143 _322_/a_193_7# output28/a_27_7# 0.00473f
C7144 _184_/a_218_334# cal 8.28e-20
C7145 _184_/a_505_n19# input1/X 0.0275f
C7146 _313_/Q _313_/a_448_7# 8.92e-21
C7147 _306_/X _313_/a_1108_7# 5.5e-36
C7148 _232_/X _331_/a_1283_n19# 0.00555f
C7149 _345_/a_1182_221# _290_/A 0.00161f
C7150 _273_/A ctlp[2] 0.0317f
C7151 _337_/Q _311_/D 0.0553f
C7152 _179_/a_27_7# _192_/B 1.49e-20
C7153 _347_/a_27_7# _347_/a_639_7# -0.0015f
C7154 _169_/Y _301_/a_512_257# 0.00115f
C7155 _169_/B _301_/a_240_7# 4.79e-21
C7156 _147_/A _254_/B 0.0449f
C7157 _236_/B _322_/Q 0.00109f
C7158 _331_/Q _316_/D 0.0322f
C7159 _165_/X _299_/X 0.00888f
C7160 _167_/X _347_/Q 0.00109f
C7161 _244_/B _150_/C 0.00501f
C7162 _340_/a_639_7# _196_/A 0.00142f
C7163 _248_/B _225_/B 0.00206f
C7164 output13/a_27_7# clk 0.00599f
C7165 _315_/Q _268_/a_39_257# 0.0383f
C7166 _267_/A _311_/a_1108_7# 3.81e-19
C7167 _252_/a_27_7# _216_/a_27_7# 9.16e-20
C7168 _310_/D clkc 5.2e-19
C7169 _149_/A _254_/B 0.00232f
C7170 _149_/A _317_/D 3.34e-19
C7171 _306_/S _315_/D 0.257f
C7172 _305_/a_218_7# _192_/B 2.62e-21
C7173 _306_/X _254_/A 0.00749f
C7174 _195_/a_373_7# VGND -4.52e-19
C7175 _335_/Q _298_/A 2.21e-20
C7176 _342_/Q _298_/B 0.13f
C7177 _309_/a_193_7# _284_/A 0.607f
C7178 _291_/a_39_257# _310_/a_1108_7# 3.04e-19
C7179 _340_/a_193_7# _340_/a_1108_7# -3.36e-19
C7180 _340_/a_27_7# _340_/a_448_7# -0.00733f
C7181 _219_/a_93_n19# _328_/D 4.72e-19
C7182 _277_/Y _167_/a_109_257# 0.00481f
C7183 ctln[6] VPWR 0.252f
C7184 _281_/Y VGND 0.527f
C7185 _172_/Y _172_/B 0.0108f
C7186 _346_/a_1032_373# _162_/X 0.0109f
C7187 _317_/a_193_7# _244_/B 0.00127f
C7188 _323_/a_651_373# clk 4.61e-19
C7189 _229_/a_76_159# _298_/X 1.69e-21
C7190 _254_/Y _225_/B 0.214f
C7191 _275_/Y _267_/A 0.361f
C7192 _310_/a_543_7# _310_/D 0.0337f
C7193 _326_/a_448_7# _181_/X 2.34e-19
C7194 _166_/Y VGND 0.714f
C7195 _288_/A _273_/A 0.656f
C7196 _186_/a_297_7# _146_/C 0.00203f
C7197 _257_/a_222_53# _215_/A 7.21e-22
C7198 _336_/a_27_7# _336_/a_1108_7# -2.98e-20
C7199 _336_/a_193_7# _336_/a_1283_n19# -4.76e-19
C7200 _327_/a_27_7# _216_/X 0.0107f
C7201 _240_/B VPWR 0.223f
C7202 _215_/A _297_/Y 2.05e-21
C7203 _273_/A _162_/X 0.00744f
C7204 _259_/a_113_257# _340_/CLK 9.94e-19
C7205 _325_/Q _224_/a_93_n19# 0.0274f
C7206 _162_/a_27_7# _171_/a_215_7# 1.35e-19
C7207 _273_/A _287_/a_39_257# 0.00415f
C7208 _286_/B _340_/CLK 0.113f
C7209 _277_/Y _297_/Y 0.00842f
C7210 _330_/Q clkbuf_1_0_0_clk/a_75_172# 5.15e-19
C7211 _164_/Y _346_/SET_B 0.0101f
C7212 _165_/a_78_159# _165_/a_292_257# -1.09e-21
C7213 _172_/A _183_/a_471_7# 1.28e-19
C7214 _343_/a_193_7# _185_/A 0.0156f
C7215 _248_/B _314_/a_543_7# 3.74e-19
C7216 _327_/a_193_7# _320_/Q 3.88e-21
C7217 _327_/a_27_7# _329_/Q 2.31e-20
C7218 _345_/D _147_/Y 0.00264f
C7219 _329_/D VGND 0.0891f
C7220 _306_/X _309_/D 8.22e-21
C7221 _346_/a_1182_221# _299_/a_215_7# 9.92e-20
C7222 _327_/a_27_7# _327_/a_761_249# -0.00751f
C7223 _258_/a_505_n19# _339_/Q 2.33e-20
C7224 _339_/Q _311_/D 0.00567f
C7225 _322_/a_1108_7# result[7] 0.00144f
C7226 _167_/X _297_/B 0.166f
C7227 _313_/a_1108_7# _147_/Y 1.93e-19
C7228 _318_/Q _317_/a_27_7# 4.06e-19
C7229 _301_/a_240_7# _170_/a_226_7# 4.01e-19
C7230 _324_/a_193_7# _342_/Q 3.17e-21
C7231 _323_/a_448_7# cal 0.00285f
C7232 _342_/a_1283_n19# _149_/a_27_7# 0.00789f
C7233 _333_/a_1217_7# _190_/A 3.47e-19
C7234 _306_/a_505_n19# _284_/A 0.0275f
C7235 _315_/Q _316_/a_27_7# 3.64e-20
C7236 output22/a_27_7# _316_/a_1283_n19# 1.11e-21
C7237 _329_/a_761_249# _330_/Q 0.00238f
C7238 _277_/Y _310_/a_193_7# 5.13e-20
C7239 repeater43/X _330_/a_1270_373# -3.58e-20
C7240 _262_/a_199_7# _297_/Y 1.72e-19
C7241 _331_/D _331_/a_761_249# 6.11e-19
C7242 _288_/A trim[4] 5.16e-19
C7243 _227_/A _210_/a_27_7# 1.42e-20
C7244 _326_/a_27_7# _326_/a_761_249# -0.0166f
C7245 _211_/a_373_7# _339_/D 8.91e-22
C7246 _328_/a_27_7# _320_/Q 0.00935f
C7247 _292_/A _165_/a_215_7# 0.00233f
C7248 _273_/A _299_/a_493_257# 3.37e-19
C7249 _315_/D _327_/D 9.3e-21
C7250 _255_/B _217_/A 4.17e-20
C7251 _339_/D _198_/a_346_7# 2.5e-19
C7252 repeater43/X _333_/a_1283_n19# -0.0114f
C7253 _329_/a_193_7# VPWR -0.31f
C7254 _328_/Q VPWR 0.519f
C7255 _254_/A _147_/Y 0.56f
C7256 _308_/a_76_159# _306_/S 0.0127f
C7257 _296_/a_295_257# VPWR -4.51e-19
C7258 _298_/B _204_/Y 0.00217f
C7259 _198_/a_250_257# _202_/a_93_n19# 0.00113f
C7260 _172_/A cal 2.23e-19
C7261 _196_/A _346_/SET_B 0.0116f
C7262 _329_/a_543_7# _297_/B 1.15e-20
C7263 _252_/a_109_257# _212_/X 4.8e-20
C7264 _307_/a_505_n19# _162_/X 6.89e-21
C7265 repeater43/X _223_/a_93_n19# 5.02e-19
C7266 _322_/a_448_7# result[6] 0.00323f
C7267 output22/a_27_7# _315_/Q 0.0383f
C7268 _290_/A _309_/a_543_7# 3.35e-19
C7269 _333_/a_448_7# _207_/C 0.007f
C7270 _333_/a_1270_373# _206_/A 3.05e-19
C7271 _332_/a_193_7# _332_/D 0.058f
C7272 cal _335_/D 0.00131f
C7273 cal _198_/a_250_257# 0.0757f
C7274 _301_/a_245_257# _299_/X 5.17e-19
C7275 _301_/a_51_257# _347_/Q 0.039f
C7276 _167_/a_109_7# _160_/X 7.84e-19
C7277 _266_/a_113_257# clkc 1.42e-20
C7278 _294_/Y _309_/Q 0.0019f
C7279 _313_/Q _337_/Q 9.78e-19
C7280 _277_/Y _242_/A 0.0368f
C7281 _153_/a_109_53# _154_/A 2.4e-19
C7282 _153_/a_297_257# _153_/A 5.77e-19
C7283 _347_/a_543_7# _347_/D 0.00208f
C7284 _334_/a_1108_7# _343_/Q 2.27e-19
C7285 _308_/X _150_/a_27_7# 4.94e-19
C7286 _283_/A _315_/D 0.0116f
C7287 _194_/A _201_/a_27_7# 7.76e-19
C7288 _164_/A _345_/Q 0.0595f
C7289 _275_/Y _194_/X 4.35e-21
C7290 _309_/D _147_/Y 2.09e-21
C7291 _269_/A VPWR 1.15f
C7292 _227_/A _175_/Y 4.11e-19
C7293 _258_/S _201_/a_27_7# 6.57e-21
C7294 _300_/Y _297_/Y 1.42e-19
C7295 _342_/a_193_7# output30/a_27_7# 0.00128f
C7296 _315_/a_193_7# _315_/a_1108_7# -0.00656f
C7297 _333_/a_761_249# _192_/B 2.23e-20
C7298 _333_/a_1283_n19# _191_/B 7.12e-19
C7299 _331_/Q _331_/a_27_7# 0.632f
C7300 _230_/a_27_7# _318_/a_27_7# 0.00104f
C7301 output29/a_27_7# _322_/Q 0.0404f
C7302 _326_/Q _224_/a_93_n19# 0.00444f
C7303 _340_/a_27_7# _190_/A 3.05e-19
C7304 _310_/a_805_7# _310_/Q 1.11e-19
C7305 clkbuf_2_1_0_clk/A _265_/B 9.17e-21
C7306 _326_/D _181_/X 0.00166f
C7307 _187_/a_27_7# _248_/B 0.0385f
C7308 _343_/D VPWR 0.546f
C7309 clkbuf_0_clk/X _227_/a_113_7# 9.73e-20
C7310 _185_/A VGND 1.33f
C7311 _242_/A _304_/X 0.0129f
C7312 _209_/a_27_257# _154_/A 0.0575f
C7313 _209_/a_109_7# _153_/A 4.6e-19
C7314 _248_/B _315_/D 0.742f
C7315 _338_/a_1108_7# _340_/CLK 0.0659f
C7316 _294_/Y _311_/a_193_7# 8.89e-21
C7317 _167_/a_373_7# VPWR -6.09e-19
C7318 _167_/a_109_257# VGND 4.2e-19
C7319 _275_/Y _167_/X 2.02e-20
C7320 _342_/D _323_/Q 8.11e-22
C7321 _346_/SET_B _347_/a_1283_n19# 0.0391f
C7322 _235_/a_113_257# _234_/B 4.01e-20
C7323 _285_/A _284_/A 0.155f
C7324 _219_/a_346_7# _232_/X 8.06e-19
C7325 _181_/X _222_/a_256_7# 6.21e-19
C7326 _337_/a_27_7# _194_/A 5.07e-21
C7327 _325_/Q _217_/A 0.215f
C7328 _265_/B _310_/Q 0.00245f
C7329 _309_/a_651_373# _306_/S 2.16e-21
C7330 _207_/a_181_7# _153_/B 1.13e-19
C7331 _301_/a_51_257# _297_/B 1.12e-19
C7332 _338_/a_193_7# _337_/a_27_7# 3.6e-22
C7333 _338_/a_27_7# _337_/a_193_7# 5.26e-19
C7334 _196_/A _206_/A 1.49e-20
C7335 _298_/C _190_/A 0.00574f
C7336 _286_/B _313_/a_543_7# 0.00325f
C7337 _196_/A _313_/a_761_249# 9.96e-21
C7338 _255_/X VPWR 0.723f
C7339 _340_/a_651_373# _340_/CLK 2.63e-21
C7340 _164_/Y _147_/A 1.21e-21
C7341 _257_/a_448_7# VPWR 0.00321f
C7342 _257_/a_222_53# VGND 0.00135f
C7343 _323_/D cal 0.0414f
C7344 _217_/a_27_7# _331_/Q 8.56e-20
C7345 _165_/a_78_159# _346_/SET_B 0.00106f
C7346 _297_/Y VGND 0.678f
C7347 clkc VPWR 0.658f
C7348 _279_/Y _340_/CLK 0.821f
C7349 _306_/X _202_/a_250_257# 1.17e-20
C7350 _258_/a_535_334# _284_/A 1.21e-19
C7351 _279_/Y _347_/D 0.101f
C7352 _224_/a_93_n19# _224_/a_256_7# -6.6e-20
C7353 _332_/a_651_373# _333_/Q 0.00164f
C7354 _332_/a_1270_373# _332_/Q 3.11e-20
C7355 clkbuf_0_clk/X _248_/a_109_257# 3.29e-19
C7356 _210_/a_109_257# VPWR 2.59e-20
C7357 _308_/a_76_159# _283_/A 1.61e-19
C7358 _330_/Q _319_/D 0.00151f
C7359 _172_/A _284_/A 0.302f
C7360 _305_/a_218_7# _260_/A 1.66e-19
C7361 _328_/a_1217_7# _320_/Q 6.31e-21
C7362 _328_/a_805_7# _329_/Q 0.00261f
C7363 _230_/a_27_7# _246_/B 1.75e-20
C7364 _196_/A _156_/a_39_257# 0.00909f
C7365 _161_/Y _267_/A 6.64e-20
C7366 _329_/a_1462_7# VPWR 4.44e-19
C7367 _329_/a_805_7# VGND -7.11e-19
C7368 _272_/a_39_257# _242_/A 1.88e-20
C7369 _300_/Y _242_/A 3.48e-21
C7370 _338_/a_651_373# _338_/D 8.49e-19
C7371 _338_/a_543_7# _338_/Q 2.68e-20
C7372 _338_/a_448_7# _346_/SET_B 0.00349f
C7373 _306_/X input1/X 1.04e-20
C7374 _181_/a_27_7# _228_/A 0.00778f
C7375 _206_/A _298_/X 1.58e-21
C7376 _286_/B _304_/S 0.011f
C7377 _308_/S _306_/S 0.00928f
C7378 _329_/Q _319_/a_193_7# 1.02e-19
C7379 _215_/A _336_/Q 2.26e-19
C7380 _310_/a_193_7# VGND 0.0209f
C7381 _310_/a_543_7# VPWR 0.0424f
C7382 _198_/a_250_257# _284_/A 0.00138f
C7383 input4/X _332_/a_193_7# 4.94e-20
C7384 _344_/a_381_7# _344_/Q 3.32e-20
C7385 _344_/a_1182_221# _344_/D 6.28e-20
C7386 _341_/a_639_7# _248_/A 0.00114f
C7387 _182_/a_510_7# _192_/B 2.73e-19
C7388 _297_/A _302_/a_77_159# 0.00732f
C7389 _294_/Y _309_/a_1108_7# 1.48e-20
C7390 _258_/a_76_159# _194_/X 3.29e-20
C7391 _296_/Y _162_/X 0.0222f
C7392 _334_/a_1108_7# _204_/a_27_7# 8.13e-20
C7393 _319_/Q _320_/a_448_7# 1.83e-19
C7394 output23/a_27_7# result[2] 0.0111f
C7395 clkbuf_2_1_0_clk/A _170_/a_76_159# 4.57e-19
C7396 _304_/a_306_329# _304_/S 0.00563f
C7397 _264_/a_199_7# VPWR -3.16e-19
C7398 _316_/Q _230_/a_27_7# 6.17e-21
C7399 _341_/Q _227_/A 0.00109f
C7400 _333_/D _207_/C 0.425f
C7401 _232_/A _246_/B 0.144f
C7402 _340_/a_1270_373# _346_/SET_B 7.91e-20
C7403 _340_/a_1108_7# _338_/Q 5.27e-21
C7404 _286_/B _225_/X 0.485f
C7405 _196_/A _147_/A 0.0348f
C7406 _307_/X _286_/B 0.00974f
C7407 _273_/A _165_/a_215_7# 9.72e-19
C7408 _153_/A _154_/A 0.277f
C7409 _317_/Q _271_/A 0.289f
C7410 _332_/a_193_7# _207_/C 0.00173f
C7411 _332_/a_543_7# _206_/A 8.85e-19
C7412 _339_/a_27_7# _338_/a_193_7# 0.00934f
C7413 _339_/a_193_7# _338_/a_27_7# 0.00524f
C7414 _343_/CLK _343_/Q 1.6e-19
C7415 _271_/A _205_/a_297_7# 1.15e-19
C7416 _309_/a_193_7# _310_/a_761_249# 5.17e-21
C7417 _196_/A _149_/A 7.4e-21
C7418 _259_/a_113_257# _267_/B 0.0347f
C7419 _229_/a_489_373# _248_/A 1.97e-19
C7420 _307_/a_505_n19# _298_/C 1.24e-19
C7421 ctln[6] _211_/a_27_257# 0.00465f
C7422 _196_/A _339_/a_448_7# 1.46e-19
C7423 _321_/a_27_7# _246_/B 3.05e-21
C7424 _342_/a_761_249# _228_/A 1.08e-20
C7425 _181_/a_27_7# _216_/A 0.0126f
C7426 _327_/a_448_7# _346_/SET_B 0.0019f
C7427 _324_/a_543_7# _326_/Q 4.91e-19
C7428 _316_/Q _232_/A 0.00717f
C7429 _285_/A trim[2] 2.74e-20
C7430 trim[0] _290_/A 4.08e-20
C7431 _346_/a_193_7# _346_/a_476_7# -0.0132f
C7432 clkbuf_0_clk/a_110_7# _162_/X 3.5e-19
C7433 _343_/CLK _332_/a_1283_n19# 7.6e-20
C7434 _339_/Q _312_/a_1283_n19# 9.72e-19
C7435 _242_/A VGND 1.95f
C7436 repeater43/X _341_/a_761_249# -0.00437f
C7437 _335_/Q VGND 0.261f
C7438 _177_/A _150_/C 0.154f
C7439 _203_/a_80_n19# _284_/A 4.84e-20
C7440 _178_/a_27_7# _298_/C 0.0914f
C7441 _343_/a_1270_373# _175_/Y 3.27e-19
C7442 _340_/a_193_7# _339_/a_761_249# 5.17e-21
C7443 _340_/a_761_249# _339_/a_193_7# 7.54e-21
C7444 _340_/a_543_7# _339_/a_27_7# 3.45e-20
C7445 _147_/A _298_/X 5.35e-19
C7446 _340_/a_27_7# _339_/a_543_7# 2.16e-20
C7447 _342_/a_448_7# sample 4.88e-19
C7448 _305_/a_505_n19# _216_/A 5.34e-21
C7449 _315_/a_27_7# _315_/D 0.154f
C7450 _320_/a_543_7# _328_/Q 1.88e-20
C7451 _242_/A _318_/a_1108_7# 0.0065f
C7452 _254_/A _347_/a_193_7# 1.03e-20
C7453 _326_/Q _217_/A 0.193f
C7454 _298_/a_109_7# VGND 0.00107f
C7455 _275_/Y clkbuf_1_1_0_clk/a_75_172# 1.12e-20
C7456 _329_/a_448_7# _330_/D 0.00274f
C7457 _149_/A _298_/X 0.0106f
C7458 input1/X _147_/Y 0.13f
C7459 _336_/a_193_7# VPWR -0.319f
C7460 _181_/X _331_/a_193_7# 2.94e-19
C7461 _328_/a_1108_7# _346_/SET_B -0.00474f
C7462 cal _312_/a_448_7# 1.41e-21
C7463 _290_/A _311_/Q 0.00244f
C7464 _277_/A _297_/B 0.0216f
C7465 _321_/a_805_7# _321_/Q 0.00216f
C7466 _343_/a_27_7# en 1.01e-20
C7467 repeater43/X _216_/X 1.01e-19
C7468 _322_/D VGND 0.0815f
C7469 _292_/A _345_/Q 0.74f
C7470 _258_/S _313_/a_651_373# 8.9e-21
C7471 repeater43/X _316_/a_543_7# 0.0052f
C7472 _271_/Y rstn 0.0104f
C7473 _288_/Y _162_/A 0.146f
C7474 _147_/A _347_/a_1283_n19# 0.011f
C7475 _324_/a_1108_7# _224_/a_93_n19# 2.26e-20
C7476 _321_/a_448_7# VGND -0.00451f
C7477 _321_/a_1270_373# VPWR 1.24e-19
C7478 _283_/Y _193_/Y 1.93e-19
C7479 rstn _335_/a_761_249# 0.0441f
C7480 input4/X _208_/a_78_159# 3.91e-21
C7481 _160_/A _345_/Q 0.00515f
C7482 _169_/Y _160_/X 0.487f
C7483 _341_/a_1108_7# _304_/S 0.00303f
C7484 _329_/a_27_7# _232_/X 2.15e-20
C7485 _321_/a_651_373# _318_/a_1283_n19# 6.19e-20
C7486 _224_/a_346_7# _304_/X -8.88e-34
C7487 _224_/a_93_n19# _324_/D 0.00254f
C7488 _153_/a_403_257# VGND -0.00106f
C7489 _332_/D _190_/A 1.61e-20
C7490 output14/a_27_7# output28/a_27_7# 3.1e-20
C7491 input2/a_27_7# _285_/Y 0.00908f
C7492 _272_/a_121_257# _326_/Q 1.94e-19
C7493 _308_/S _283_/A 2.01e-19
C7494 _267_/A _312_/a_543_7# 8.61e-19
C7495 _305_/X _192_/B 0.0278f
C7496 _327_/a_27_7# _327_/Q 0.143f
C7497 _326_/a_761_249# repeater43/X 0.0181f
C7498 clkbuf_2_3_0_clk/a_75_172# VPWR 0.0948f
C7499 _258_/S _157_/a_27_7# 7.49e-21
C7500 _343_/CLK _229_/a_76_159# 1.46e-20
C7501 _338_/D _346_/SET_B 0.119f
C7502 _147_/Y _286_/Y 3.15e-21
C7503 _170_/a_226_7# _346_/D 3.35e-22
C7504 _206_/A _204_/a_27_257# 3.1e-19
C7505 ctln[2] output34/a_27_7# 3.34e-19
C7506 _326_/a_27_7# _327_/Q 1.34e-19
C7507 _281_/A _330_/a_543_7# 3.64e-19
C7508 output15/a_27_7# result[7] 0.00816f
C7509 _341_/a_1283_n19# _150_/C 6.36e-19
C7510 _310_/a_1462_7# VGND 1.37e-19
C7511 _199_/a_93_n19# VGND 0.00294f
C7512 _199_/a_256_7# VPWR -5.91e-19
C7513 _307_/a_76_159# _295_/a_79_n19# 2.3e-20
C7514 _281_/Y _330_/a_27_7# 4.01e-19
C7515 _167_/X _161_/Y 2.09e-19
C7516 _188_/a_76_159# _341_/D 0.00264f
C7517 _307_/X _341_/a_1108_7# 4.69e-22
C7518 ctln[5] _343_/CLK 0.011f
C7519 _337_/a_27_7# _201_/a_27_7# 8.21e-21
C7520 _185_/A _323_/a_651_373# 0.00556f
C7521 _273_/A output35/a_27_7# 4.6e-20
C7522 _281_/Y _318_/Q 0.00441f
C7523 _313_/D _306_/S 0.0733f
C7524 _334_/D _204_/a_27_257# 0.00366f
C7525 _343_/CLK _208_/a_215_7# 0.00521f
C7526 _279_/Y _156_/a_121_257# 1.86e-19
C7527 output12/a_27_7# _333_/a_27_7# 2.01e-21
C7528 _302_/a_77_159# _347_/a_761_249# 1.63e-19
C7529 _183_/a_27_7# _286_/B 0.00621f
C7530 _183_/a_553_257# _181_/X 0.0327f
C7531 _346_/a_381_7# _346_/SET_B 0.0269f
C7532 _279_/Y _304_/S 0.0233f
C7533 clk _286_/B 0.156f
C7534 _250_/a_215_7# _147_/Y 6.53e-21
C7535 result[5] _234_/a_109_257# 8.2e-20
C7536 output27/a_27_7# _322_/D 0.0183f
C7537 _319_/Q _331_/D 1.81e-19
C7538 clkbuf_2_1_0_clk/A _278_/a_68_257# 0.0435f
C7539 _346_/a_1182_221# _275_/A 2.76e-21
C7540 _325_/a_1283_n19# _181_/X 4.42e-19
C7541 _209_/a_373_7# VGND -0.00112f
C7542 _336_/Q VGND 0.781f
C7543 result[5] _321_/a_27_7# 1.32e-19
C7544 _319_/Q _330_/a_193_7# 2.7e-20
C7545 _339_/a_1108_7# _338_/a_651_373# 2.91e-19
C7546 _340_/CLK _313_/a_27_7# 0.0273f
C7547 _317_/Q _232_/a_27_7# 0.00157f
C7548 input4/X _334_/a_543_7# 0.00217f
C7549 repeater43/X _334_/a_193_7# 0.0119f
C7550 _197_/X _306_/S 0.262f
C7551 _337_/a_1283_n19# _340_/CLK 0.068f
C7552 _296_/Y _298_/C 0.0026f
C7553 _335_/a_651_373# _335_/Q 1.48e-19
C7554 _196_/A _339_/D 0.115f
C7555 _329_/D _330_/a_27_7# 5.85e-19
C7556 _160_/X _170_/a_226_257# 0.00153f
C7557 _318_/Q _329_/D 1.57e-19
C7558 _279_/Y _225_/X 1.37e-21
C7559 _271_/A _315_/a_193_7# 1.53e-20
C7560 _333_/a_193_7# _207_/a_27_7# 5.69e-20
C7561 _271_/A _298_/A 0.0103f
C7562 _309_/a_1283_n19# _265_/B 1.22e-19
C7563 _344_/a_652_n19# _297_/Y 0.0338f
C7564 output35/a_27_7# trim[4] 0.0119f
C7565 _326_/D _346_/SET_B 2.42e-20
C7566 _334_/a_543_7# _207_/C 0.0356f
C7567 _342_/D sample 0.0141f
C7568 result[0] _304_/S 5.06e-20
C7569 _242_/a_109_257# VPWR 2.82e-19
C7570 _344_/a_1224_7# _290_/A 3.76e-19
C7571 _315_/a_1108_7# VGND 0.00207f
C7572 _315_/a_651_373# VPWR -0.00819f
C7573 _324_/a_193_7# _315_/D 2.36e-20
C7574 en ctln[0] 4.36e-22
C7575 _255_/B _308_/X 4.53e-21
C7576 _227_/A _269_/Y 2.04e-20
C7577 _342_/Q _172_/A 0.388f
C7578 _188_/a_76_159# _143_/a_27_7# 0.00233f
C7579 _324_/a_805_7# _227_/A 4.3e-19
C7580 _336_/a_1462_7# VPWR 1.82e-20
C7581 _336_/a_805_7# VGND -4.94e-19
C7582 _317_/a_27_7# _316_/a_448_7# 1.68e-20
C7583 _317_/a_448_7# _316_/a_27_7# 3.72e-20
C7584 cal _312_/D 8.38e-20
C7585 _331_/Q _281_/A 2.36e-19
C7586 _346_/a_193_7# clkbuf_2_3_0_clk/A 3.21e-22
C7587 _326_/a_27_7# _325_/a_27_7# 1.84e-20
C7588 _286_/B _301_/X 1.28e-20
C7589 _334_/a_448_7# _343_/CLK 2.63e-20
C7590 _334_/a_1108_7# _334_/D 0.0517f
C7591 _334_/a_193_7# _334_/Q 0.00355f
C7592 clkbuf_2_1_0_clk/A _311_/a_27_7# 2.25e-21
C7593 _314_/a_1283_n19# VPWR 0.0202f
C7594 _314_/a_761_249# VGND 0.00641f
C7595 _227_/A _314_/D 0.00482f
C7596 _344_/a_1602_7# comp 2.22e-19
C7597 _346_/SET_B _319_/a_651_373# 0.00363f
C7598 _346_/SET_B _313_/a_193_7# 0.00466f
C7599 _338_/a_761_249# _337_/Q 2.43e-19
C7600 _338_/D _337_/a_448_7# 3.05e-20
C7601 _346_/SET_B _337_/a_1108_7# 5.84e-19
C7602 _275_/A _319_/a_1283_n19# 8.6e-21
C7603 _165_/X _172_/B 0.0154f
C7604 clk _332_/a_761_249# 0.0184f
C7605 _224_/a_346_7# VGND 4.63e-19
C7606 _294_/A _197_/X 3.99e-20
C7607 _216_/X _331_/a_448_7# 2.32e-20
C7608 repeater43/X _236_/a_109_257# 5.18e-19
C7609 _324_/a_448_7# _304_/X 2.97e-19
C7610 _324_/a_543_7# _324_/D 0.0335f
C7611 _324_/a_1108_7# _217_/A 3.95e-19
C7612 _311_/a_1283_n19# _310_/D 5.79e-19
C7613 _196_/A _150_/a_27_7# 0.0108f
C7614 _314_/a_193_7# _314_/Q 1.22e-19
C7615 _314_/a_448_7# _297_/B 2.63e-20
C7616 _314_/a_1108_7# _314_/D 5.47e-21
C7617 _196_/A _174_/a_109_7# 6.56e-20
C7618 _170_/a_489_373# VGND -8.03e-20
C7619 _170_/a_556_7# VPWR -4.88e-19
C7620 input4/X _190_/A 2.21e-20
C7621 repeater43/X _332_/Q 0.239f
C7622 _346_/SET_B _343_/CLK 2.14e-19
C7623 _322_/a_651_373# _269_/A 0.00247f
C7624 _334_/a_193_7# _191_/B 0.00584f
C7625 _334_/a_27_7# _323_/Q 0.0058f
C7626 _263_/B _267_/A 0.0194f
C7627 _325_/a_651_373# _325_/D 8.49e-19
C7628 _320_/Q result[7] 0.00245f
C7629 _339_/a_1283_n19# _340_/CLK 6e-19
C7630 _163_/a_292_257# _345_/D 8.16e-20
C7631 _153_/a_109_53# _153_/B 1.66e-20
C7632 _323_/a_543_7# _175_/Y 6.18e-22
C7633 _217_/A _324_/D 6.65e-20
C7634 _340_/a_1283_n19# _337_/Q 0.0377f
C7635 _345_/a_27_7# _297_/B 0.0479f
C7636 _327_/a_639_7# _217_/X 1.17e-19
C7637 _327_/a_805_7# _212_/X 4.67e-19
C7638 _172_/A _264_/a_113_257# 8.8e-20
C7639 _326_/a_1283_n19# _331_/a_1283_n19# 6.99e-20
C7640 _326_/a_543_7# _331_/a_1108_7# 5.46e-20
C7641 _248_/a_109_257# _328_/Q 1.86e-19
C7642 _339_/a_27_7# _337_/a_27_7# 3.77e-20
C7643 cal _333_/D 0.213f
C7644 _214_/a_27_257# _242_/A 1.77e-20
C7645 _207_/C _190_/A 0.0168f
C7646 _273_/A _345_/Q 0.0837f
C7647 _326_/D _222_/a_346_7# 1.03e-19
C7648 _149_/A _334_/a_1108_7# 1.44e-19
C7649 _189_/a_27_7# _254_/B 1.59e-19
C7650 _164_/A _284_/A 1.33e-19
C7651 _277_/A _320_/a_193_7# 0.00775f
C7652 output14/a_27_7# output26/a_27_7# 4.94e-21
C7653 _255_/B _254_/B 1.3e-19
C7654 _216_/A _331_/Q 1.19e-21
C7655 _306_/S _333_/a_193_7# 7.39e-20
C7656 _286_/a_113_7# _286_/Y 2.88e-19
C7657 _342_/Q _244_/B 0.111f
C7658 _334_/Q _332_/Q 0.902f
C7659 _168_/a_109_257# _162_/X 0.00423f
C7660 _257_/a_79_159# _254_/B 0.00689f
C7661 _299_/X VPWR 0.523f
C7662 _341_/D _149_/A 0.00705f
C7663 ctln[6] _333_/a_1108_7# 8.13e-20
C7664 _303_/A _347_/a_27_7# 4.32e-20
C7665 _308_/a_535_334# _227_/A 8.82e-20
C7666 input4/X _337_/a_543_7# 2.12e-20
C7667 _197_/X _283_/A 0.0842f
C7668 _304_/S _316_/D 0.00774f
C7669 _209_/a_27_257# _153_/B 0.00581f
C7670 _322_/a_1283_n19# _321_/a_27_7# 0.0112f
C7671 _173_/a_76_159# _172_/Y 0.00539f
C7672 ctln[7] rstn 0.0778f
C7673 _339_/Q _338_/a_761_249# 1.3e-19
C7674 _339_/a_1108_7# _346_/SET_B 0.0133f
C7675 _248_/A _150_/C 0.00232f
C7676 repeater43/X _334_/a_1462_7# -8.62e-19
C7677 _218_/a_256_7# _304_/X 0.00107f
C7678 _309_/a_1283_n19# _310_/Q 6.49e-19
C7679 _258_/a_76_159# _336_/a_543_7# 5.06e-19
C7680 _308_/X _298_/a_27_7# 1.15e-19
C7681 _335_/D _204_/Y 0.0438f
C7682 _191_/B _332_/Q 0.0355f
C7683 _321_/Q _330_/Q 0.0794f
C7684 _324_/Q _304_/a_578_7# 4.88e-19
C7685 _313_/a_27_7# _313_/a_543_7# -0.00941f
C7686 _313_/a_193_7# _313_/a_761_249# -0.0157f
C7687 _310_/a_27_7# _254_/B 2.84e-20
C7688 _293_/a_39_257# _265_/B 1.61e-20
C7689 output21/a_27_7# _319_/Q 1.02e-20
C7690 _294_/A _289_/a_39_257# 2.03e-21
C7691 _260_/B clkbuf_0_clk/X 3.72e-20
C7692 clk _208_/a_292_257# 0.00419f
C7693 _340_/a_1283_n19# _339_/Q 0.0166f
C7694 _184_/a_76_159# _227_/A 1.29e-19
C7695 _343_/CLK _206_/A 0.151f
C7696 _260_/A _305_/X 1.13e-19
C7697 _198_/a_93_n19# _336_/a_193_7# 3.72e-20
C7698 _198_/a_250_257# _336_/a_27_7# 9.53e-21
C7699 _317_/a_193_7# _248_/A 0.00511f
C7700 _255_/a_30_13# _333_/a_1283_n19# 1.78e-20
C7701 _327_/a_543_7# clkbuf_0_clk/X 0.0115f
C7702 _313_/D _254_/Y 1.43e-19
C7703 _330_/Q _297_/B 0.0308f
C7704 _343_/a_193_7# _271_/A 1.03e-20
C7705 output6/a_27_7# VGND 0.101f
C7706 _188_/a_505_n19# _144_/A 6.34e-19
C7707 _340_/a_1108_7# _202_/a_250_257# 7.19e-20
C7708 _275_/A _212_/X 4.64e-19
C7709 _324_/a_448_7# VGND -0.00539f
C7710 _324_/a_1270_373# VPWR 6.69e-20
C7711 _271_/A _304_/X 3.49e-20
C7712 _317_/a_193_7# _331_/CLK 4.14e-19
C7713 _317_/a_27_7# _316_/D 6.96e-19
C7714 _304_/a_257_159# _284_/A 6.19e-19
C7715 _306_/a_218_7# clkbuf_2_1_0_clk/A 1.42e-19
C7716 _326_/a_651_373# _325_/a_1283_n19# 7.83e-21
C7717 _343_/CLK _334_/D 0.00982f
C7718 output7/a_27_7# _343_/CLK 0.0114f
C7719 _194_/X _263_/B 6.62e-20
C7720 clkbuf_2_1_0_clk/A _328_/D 7.83e-20
C7721 _143_/a_27_7# _149_/A 0.0485f
C7722 _283_/A _312_/a_193_7# 6.33e-20
C7723 _248_/A _331_/a_1283_n19# 6.01e-19
C7724 _318_/a_27_7# VPWR 0.0718f
C7725 _343_/a_651_373# VPWR 0.00167f
C7726 _343_/a_1108_7# VGND 6.21e-19
C7727 _346_/SET_B _313_/a_1462_7# -9.14e-19
C7728 _254_/Y _197_/X 3.9e-19
C7729 _338_/D _337_/D 0.00182f
C7730 _245_/a_113_257# _246_/B 0.0489f
C7731 _267_/A _194_/A 0.00916f
C7732 _252_/a_27_7# _251_/X 0.00721f
C7733 _281_/Y _286_/B 0.00578f
C7734 _220_/a_250_257# _279_/A 0.00593f
C7735 input4/X _339_/a_543_7# 1.81e-21
C7736 _345_/a_27_7# _275_/Y 0.0195f
C7737 _328_/a_761_249# clkbuf_0_clk/X 1.47e-21
C7738 _314_/a_1462_7# _314_/Q 6.13e-19
C7739 _297_/B _314_/D 0.0107f
C7740 _260_/B input1/X 8.1e-20
C7741 repeater43/X _282_/a_39_257# 1.53e-20
C7742 _331_/CLK _331_/a_1283_n19# 2.28e-20
C7743 _318_/a_193_7# _318_/a_761_249# -0.00517f
C7744 _318_/a_27_7# _318_/a_543_7# -0.00714f
C7745 _231_/a_676_257# _283_/A 1.84e-19
C7746 _308_/S _298_/B 5.82e-23
C7747 _325_/Q _317_/D 0.00106f
C7748 _279_/Y _301_/X 1.45e-20
C7749 _290_/A _164_/Y 0.0154f
C7750 _313_/a_193_7# _147_/A 0.0442f
C7751 _341_/a_543_7# _286_/Y 0.0338f
C7752 _345_/a_381_7# VGND 0.00395f
C7753 _345_/a_956_373# VPWR 2.49e-19
C7754 _166_/Y _286_/B 2.42e-19
C7755 _258_/S _267_/A 0.00759f
C7756 _254_/B _298_/a_27_7# 8.19e-19
C7757 _153_/A _153_/B 0.0535f
C7758 _283_/A _330_/a_1108_7# 0.0036f
C7759 _281_/Y _256_/a_209_7# 0.00101f
C7760 clk _334_/a_1283_n19# 0.00512f
C7761 _339_/a_651_373# _337_/a_1283_n19# 1.27e-19
C7762 _339_/a_1283_n19# _337_/a_651_373# 1.27e-19
C7763 _326_/D _331_/a_761_249# 3e-19
C7764 _172_/A _169_/Y 0.027f
C7765 _172_/A _225_/B 0.00748f
C7766 _283_/A _333_/a_193_7# 0.0299f
C7767 repeater43/X _327_/Q 0.0216f
C7768 _307_/X _307_/a_218_334# 8.5e-19
C7769 _188_/a_505_n19# _145_/A 0.0298f
C7770 _149_/A _343_/CLK 2.05e-21
C7771 result[2] result[3] 0.0637f
C7772 _325_/D _284_/A 3e-21
C7773 _318_/Q _242_/A 1.01f
C7774 _165_/X trimb[4] 1.12e-19
C7775 _231_/a_306_7# _232_/A 3.58e-19
C7776 input1/a_75_172# _340_/CLK 6.03e-19
C7777 _255_/X _147_/Y 0.00876f
C7778 _310_/D _171_/a_78_159# 9.68e-20
C7779 _197_/X _225_/a_145_35# 2.27e-19
C7780 _218_/a_256_7# VGND -4.18e-19
C7781 _218_/a_584_7# VPWR -3.47e-19
C7782 _333_/a_27_7# _205_/a_297_7# 9.73e-21
C7783 _333_/a_193_7# _205_/a_382_257# 1.17e-20
C7784 _198_/a_250_257# _225_/B 9.8e-21
C7785 _246_/B VPWR 1.97f
C7786 clkbuf_2_1_0_clk/a_75_172# _297_/B 4.41e-19
C7787 _178_/a_193_257# _147_/A 2.55e-20
C7788 _178_/a_27_7# _150_/C 3.47e-19
C7789 _309_/a_543_7# _309_/Q 2.1e-20
C7790 _308_/a_505_n19# VPWR 0.0562f
C7791 _293_/a_39_257# clkbuf_2_1_0_clk/A 0.00364f
C7792 _307_/X _178_/a_109_257# 0.00244f
C7793 _343_/a_193_7# _323_/a_27_7# 3.82e-19
C7794 output32/a_27_7# _297_/Y 0.00104f
C7795 _318_/a_543_7# _246_/B 2.34e-21
C7796 ctln[6] _332_/a_27_7# 0.0128f
C7797 _220_/a_584_7# VGND 5.26e-19
C7798 _226_/a_297_7# _226_/X 9.09e-19
C7799 _327_/a_543_7# _286_/Y 9.19e-22
C7800 _311_/a_1283_n19# VPWR 0.0305f
C7801 _311_/a_761_249# VGND 0.00352f
C7802 _330_/D _304_/X 0.0026f
C7803 cal _334_/a_543_7# 4.88e-19
C7804 _306_/X _336_/a_193_7# 7.79e-19
C7805 _313_/Q _336_/a_761_249# 4.25e-19
C7806 _325_/a_651_373# _248_/A 1.93e-20
C7807 ctln[1] repeater43/X 0.226f
C7808 _316_/Q VPWR 0.484f
C7809 _304_/a_578_7# _216_/A 7.11e-20
C7810 _304_/S _144_/A 0.672f
C7811 _342_/a_543_7# _298_/A 0.00132f
C7812 _252_/a_109_257# _248_/B 0.0012f
C7813 _318_/Q _322_/D 3.09e-20
C7814 _271_/Y VPWR 0.622f
C7815 _337_/a_193_7# _337_/Q 0.124f
C7816 _337_/a_1108_7# _337_/D 1.13e-19
C7817 _271_/A VGND 0.879f
C7818 _200_/a_584_7# _267_/A 0.00288f
C7819 output32/a_27_7# _310_/a_193_7# 8.24e-20
C7820 _316_/Q _318_/a_543_7# 2.51e-19
C7821 _242_/A _241_/a_199_7# 4.21e-21
C7822 _158_/Y _160_/a_27_7# 4.12e-19
C7823 _288_/A comp 8.01e-20
C7824 _335_/a_27_7# VGND -0.0287f
C7825 _335_/a_761_249# VPWR 0.00895f
C7826 _276_/a_68_257# _346_/SET_B 1.3e-19
C7827 _188_/S _227_/A 0.0482f
C7828 _315_/Q _286_/Y 5.47e-19
C7829 _292_/A _284_/A 0.014f
C7830 repeater43/X _192_/B 0.00261f
C7831 _162_/X comp 4.29e-20
C7832 _194_/X _194_/A 0.854f
C7833 _271_/A _318_/a_1108_7# 7.55e-19
C7834 _336_/Q _203_/a_209_257# 6.7e-20
C7835 _225_/B _203_/a_80_n19# 0.0184f
C7836 _160_/A _284_/A 1.8e-20
C7837 _307_/X _144_/A 8.19e-20
C7838 _327_/a_193_7# _221_/a_93_n19# 5.09e-22
C7839 _327_/a_27_7# _221_/a_250_257# 8.97e-21
C7840 _313_/a_651_373# _157_/a_27_7# 8.81e-19
C7841 _338_/a_27_7# _340_/Q 0.0157f
C7842 _338_/a_193_7# _194_/X 0.0179f
C7843 repeater43/a_27_7# clk 0.035f
C7844 _326_/D _325_/a_1108_7# 5.01e-19
C7845 _325_/a_27_7# repeater43/X 0.0068f
C7846 cal _248_/A 0.00182f
C7847 _258_/S _194_/X 5.04e-20
C7848 _318_/a_1217_7# VPWR 1.3e-19
C7849 _318_/a_639_7# VGND 1.31e-19
C7850 _346_/SET_B _174_/a_109_257# 0.00268f
C7851 _345_/a_586_7# _275_/Y 2.97e-19
C7852 _344_/a_27_7# _299_/X 1.34e-19
C7853 _307_/a_439_7# _145_/A 8.05e-20
C7854 _277_/Y _283_/Y 0.00336f
C7855 _280_/a_150_257# _248_/A 3.75e-19
C7856 cal _190_/A 0.0117f
C7857 repeater43/X _317_/a_1108_7# 0.0153f
C7858 _145_/A _304_/S 0.08f
C7859 _309_/a_448_7# VGND -0.00289f
C7860 _309_/a_1270_373# VPWR 6.24e-20
C7861 _334_/Q _192_/B 4.71e-20
C7862 _313_/a_1462_7# _147_/A 0.00217f
C7863 _340_/a_761_249# _340_/Q 0.0221f
C7864 _340_/a_193_7# _306_/S 0.00999f
C7865 _340_/a_27_7# _193_/Y 0.00629f
C7866 _340_/a_543_7# _194_/X 3.74e-19
C7867 clkbuf_0_clk/X _319_/a_1283_n19# 4.02e-19
C7868 _330_/D _220_/a_93_n19# 1.41e-20
C7869 ctln[1] _191_/B 1.44e-20
C7870 _315_/a_448_7# _244_/B 0.00392f
C7871 _315_/a_1283_n19# _317_/D 1.15e-21
C7872 _258_/a_505_n19# _347_/Q 1.35e-19
C7873 ctln[5] _195_/a_109_257# 0.00299f
C7874 _197_/a_27_7# _190_/A 1.07e-21
C7875 _336_/a_193_7# _147_/Y 0.0272f
C7876 _331_/CLK _280_/a_150_257# 9.54e-19
C7877 _285_/A output37/a_27_7# 0.00558f
C7878 _342_/Q _192_/a_68_257# 7.72e-20
C7879 _219_/a_93_n19# _346_/SET_B 0.026f
C7880 _279_/Y _281_/Y 0.063f
C7881 _258_/S _167_/X 1.05e-21
C7882 _331_/D _326_/Q 5.09e-19
C7883 _234_/B _322_/Q 0.0549f
C7884 _220_/a_256_7# _328_/D 0.00134f
C7885 _290_/A _165_/a_78_159# 0.0094f
C7886 _339_/D _337_/a_1108_7# 1.88e-19
C7887 _339_/a_193_7# _337_/Q 9.64e-21
C7888 _339_/Q _337_/a_193_7# 0.389f
C7889 _321_/a_1283_n19# _322_/Q 0.011f
C7890 _322_/a_193_7# _318_/D 1.94e-21
C7891 repeater43/X _331_/a_1270_373# -9.44e-20
C7892 _172_/Y _172_/a_109_257# 0.00301f
C7893 _296_/Y _150_/C 6.29e-20
C7894 _189_/a_27_7# _196_/A 0.0233f
C7895 _231_/a_79_n19# _298_/A 0.00235f
C7896 _191_/B _192_/B 1.33f
C7897 _283_/A _333_/a_1462_7# 0.0019f
C7898 _331_/a_193_7# _331_/a_761_249# -0.0105f
C7899 _331_/a_27_7# _331_/a_543_7# -0.00728f
C7900 _307_/X _145_/A 0.0448f
C7901 result[5] VPWR 0.361f
C7902 _301_/a_149_7# _162_/X 0.00253f
C7903 _255_/B _196_/A 0.193f
C7904 _331_/a_1108_7# _212_/X 3.86e-20
C7905 _331_/a_1283_n19# _217_/X 1.91e-19
C7906 _295_/a_512_7# _286_/Y 2.04e-19
C7907 _325_/a_543_7# _304_/S 4.86e-19
C7908 _337_/a_543_7# _202_/a_93_n19# 3.8e-21
C7909 _320_/a_27_7# VPWR 0.0661f
C7910 _346_/a_1182_221# _286_/Y 1.45e-20
C7911 _257_/a_222_53# _286_/B 7.46e-19
C7912 _277_/A output17/a_27_7# 1.5e-19
C7913 _257_/a_79_159# _196_/A 0.0862f
C7914 _323_/a_761_249# VPWR 0.0154f
C7915 _323_/a_27_7# VGND 0.0236f
C7916 _330_/D VGND 0.332f
C7917 _286_/B _297_/Y 0.00961f
C7918 _197_/X _194_/a_27_7# 1.49e-21
C7919 _183_/a_471_7# _178_/a_27_7# 1.06e-19
C7920 clkbuf_2_3_0_clk/A _337_/Q 0.00985f
C7921 _146_/a_184_13# _147_/A 0.00219f
C7922 _146_/a_29_271# _150_/C 0.0763f
C7923 _188_/a_218_7# _146_/C 0.00124f
C7924 _342_/D _175_/Y 7.72e-20
C7925 _320_/a_761_249# _297_/B 0.0443f
C7926 _195_/a_27_257# _340_/CLK 1.36e-20
C7927 _275_/Y _311_/a_448_7# 0.00745f
C7928 cal _337_/a_543_7# 2.79e-19
C7929 _343_/D _176_/a_27_7# 4.32e-20
C7930 _345_/a_27_7# _161_/Y 4.95e-19
C7931 _254_/B _154_/A 0.0475f
C7932 trim[2] _292_/A 4.27e-20
C7933 _290_/A trim[3] 0.00139f
C7934 _200_/a_250_257# _193_/Y 0.0025f
C7935 _200_/a_346_7# _340_/Q 8.31e-19
C7936 _291_/a_39_257# _312_/a_1283_n19# 0.0119f
C7937 _256_/a_80_n19# _255_/X 0.00251f
C7938 _304_/a_257_159# _144_/a_27_7# 2.95e-19
C7939 _263_/B _310_/a_1108_7# 1.23e-19
C7940 _172_/A _315_/D 4.62e-21
C7941 _342_/Q _177_/A 0.0921f
C7942 _186_/a_297_7# VPWR 4.47e-20
C7943 _186_/a_79_n19# VGND 0.0135f
C7944 output26/a_27_7# _321_/D 4.83e-20
C7945 _149_/a_27_7# _226_/X 1.07e-20
C7946 _325_/Q _223_/a_584_7# 0.00419f
C7947 _228_/A _347_/D 5.04e-20
C7948 _335_/a_193_7# _335_/a_448_7# -0.00779f
C7949 _329_/a_761_249# _216_/X 1.36e-19
C7950 _232_/X _315_/D 9.08e-19
C7951 _345_/a_1032_373# _344_/a_1182_221# 3.86e-20
C7952 _345_/a_1182_221# _344_/a_1032_373# 7.25e-20
C7953 _328_/a_1108_7# _319_/Q 0.0336f
C7954 _232_/a_27_7# VGND 0.0542f
C7955 _335_/a_1217_7# VGND 9.02e-20
C7956 _341_/a_543_7# _269_/A 0.00573f
C7957 repeater43/X _146_/C 0.00682f
C7958 _343_/a_27_7# _342_/a_1283_n19# 1.17e-20
C7959 _343_/a_543_7# _342_/a_193_7# 8.25e-19
C7960 _343_/a_193_7# _342_/a_543_7# 1.83e-20
C7961 _343_/a_761_249# _342_/a_761_249# 7.88e-21
C7962 input2/a_27_7# _162_/A 0.0135f
C7963 _342_/Q _333_/D 2.47e-21
C7964 _285_/Y _297_/B 6.2e-21
C7965 _321_/Q _212_/a_27_7# 0.00174f
C7966 _329_/a_543_7# _320_/Q 3.14e-20
C7967 _339_/a_1108_7# _339_/D 6.56e-21
C7968 _339_/a_193_7# _339_/Q 7.3e-19
C7969 _268_/a_39_257# _248_/B 1.94e-19
C7970 _328_/a_1283_n19# _329_/D 3.12e-21
C7971 ctlp[0] _269_/A 0.011f
C7972 _327_/a_543_7# _328_/Q 1.35e-19
C7973 _329_/a_1283_n19# _327_/a_27_7# 1.82e-21
C7974 _329_/a_193_7# _327_/a_543_7# 1.53e-20
C7975 _338_/a_1462_7# _194_/X 2.52e-19
C7976 _346_/SET_B _195_/a_109_257# 9.06e-19
C7977 _171_/a_78_159# VPWR 0.0329f
C7978 _325_/a_1217_7# repeater43/X -1.57e-19
C7979 _309_/Q _311_/Q 3.1e-20
C7980 _346_/SET_B _344_/D 0.0967f
C7981 _341_/a_1108_7# _185_/A 9.46e-22
C7982 clkbuf_2_3_0_clk/A _339_/Q 0.00786f
C7983 _190_/A _284_/A 0.064f
C7984 clkbuf_0_clk/X _212_/X 0.366f
C7985 _216_/A _340_/CLK 0.0753f
C7986 _286_/B _335_/Q 9.44e-22
C7987 _340_/a_193_7# _283_/A 1.57e-20
C7988 cal _267_/a_109_257# 1.89e-19
C7989 _275_/Y _309_/a_805_7# 2.53e-19
C7990 _277_/Y _312_/a_27_7# 0.0058f
C7991 trim[0] _311_/a_193_7# 0.00168f
C7992 _273_/A _284_/A 0.0534f
C7993 _346_/Q _346_/SET_B 0.0535f
C7994 _157_/A _313_/a_448_7# 6.63e-20
C7995 _328_/a_761_249# _328_/Q 0.00118f
C7996 _346_/a_27_7# _306_/S 1.84e-20
C7997 _269_/A _316_/a_1283_n19# 0.0113f
C7998 _182_/a_297_257# _298_/A 0.00305f
C7999 output13/a_27_7# _335_/a_27_7# 1.1e-19
C8000 _274_/a_121_257# _240_/B 5.66e-20
C8001 _230_/a_27_7# _316_/a_193_7# 2.42e-21
C8002 _315_/D _244_/B 0.0174f
C8003 _306_/X _299_/X 2.91e-19
C8004 ctln[5] _340_/D 0.00546f
C8005 _345_/a_193_7# _172_/B 0.0101f
C8006 _154_/a_27_7# VPWR 0.0478f
C8007 _336_/a_1462_7# _147_/Y 0.00215f
C8008 _244_/a_109_257# VPWR 5.13e-19
C8009 _341_/a_1283_n19# _342_/Q 0.0139f
C8010 ctln[7] VPWR 1.82f
C8011 _283_/Y VGND 0.174f
C8012 _342_/D _341_/Q 2.08e-21
C8013 _346_/a_1602_7# _166_/Y 0.0117f
C8014 _145_/A _183_/a_27_7# 5.96e-19
C8015 _296_/Y _183_/a_471_7# 5.85e-21
C8016 ctln[6] _333_/Q 0.00559f
C8017 _194_/X _201_/a_27_7# 0.0042f
C8018 _311_/a_193_7# _311_/Q 1.36e-19
C8019 _179_/a_27_7# VPWR 0.0877f
C8020 _297_/A _225_/B 2.32e-20
C8021 _162_/X _298_/A 0.0111f
C8022 _146_/C _191_/B 0.00155f
C8023 _145_/A clk 6.39e-19
C8024 _322_/a_1283_n19# VPWR 0.00389f
C8025 _322_/a_761_249# VGND 0.00338f
C8026 _218_/a_346_7# _232_/X 5.22e-19
C8027 _324_/Q _304_/S 0.235f
C8028 _346_/a_193_7# _165_/X 0.0059f
C8029 _316_/a_193_7# _232_/A 7.07e-19
C8030 _170_/a_556_7# _147_/Y 3.04e-19
C8031 rstn _338_/a_27_7# 1.65e-19
C8032 input4/a_27_7# _338_/a_1283_n19# 5.15e-19
C8033 _337_/a_543_7# _284_/A 3.75e-19
C8034 _319_/Q _236_/B 0.134f
C8035 _320_/a_1217_7# VPWR 8.54e-20
C8036 _320_/a_639_7# VGND 0.00328f
C8037 trim[4] _284_/A 0.00589f
C8038 _298_/a_27_7# _298_/X 0.00211f
C8039 _238_/a_109_257# VGND -0.00108f
C8040 _323_/a_1217_7# VGND 5.4e-20
C8041 _157_/A _191_/B 6.75e-21
C8042 output33/a_27_7# _338_/Q 1.55e-20
C8043 _315_/Q _269_/A 0.124f
C8044 _333_/D _204_/Y 2.04e-20
C8045 _322_/a_1283_n19# _318_/a_543_7# 8.9e-21
C8046 _322_/a_27_7# _318_/a_651_373# 7.68e-22
C8047 _305_/a_218_7# VPWR -3.78e-19
C8048 _305_/a_218_334# VGND -6.08e-19
C8049 _292_/Y _292_/A 0.0573f
C8050 _344_/a_1602_7# VGND 0.0201f
C8051 _344_/a_562_373# VPWR 5.56e-19
C8052 _143_/a_181_7# _228_/A 1.6e-19
C8053 _275_/Y _311_/D 0.0118f
C8054 _332_/a_193_7# _204_/Y 7.04e-21
C8055 _181_/X _209_/X 1.09e-19
C8056 _343_/a_448_7# _323_/D 0.0101f
C8057 _326_/Q _223_/a_584_7# 9.53e-19
C8058 _307_/X _324_/Q 8.35e-19
C8059 _307_/a_505_n19# _284_/A 2.63e-19
C8060 _260_/B _255_/X 0.0149f
C8061 _326_/a_27_7# _232_/A 2.48e-21
C8062 _326_/D _319_/Q 9.79e-21
C8063 _257_/a_448_7# _260_/B 0.00533f
C8064 _325_/a_27_7# _325_/a_639_7# -0.0015f
C8065 _258_/S _310_/a_1108_7# 1.31e-20
C8066 _344_/Q _345_/D 2.28e-20
C8067 _255_/a_30_13# _332_/Q 2.76e-19
C8068 _337_/a_27_7# _194_/X 0.00941f
C8069 _275_/Y _285_/Y 4.87e-20
C8070 _324_/a_27_7# _252_/a_27_7# 2.07e-20
C8071 _342_/a_543_7# VGND -0.00116f
C8072 _342_/a_1108_7# VPWR 0.0153f
C8073 _335_/a_193_7# _335_/D 8.28e-19
C8074 _297_/A _314_/a_543_7# 2.52e-19
C8075 trim[1] _310_/D 0.00213f
C8076 _324_/Q _317_/a_27_7# 2.23e-21
C8077 _212_/X _286_/Y 0.05f
C8078 _299_/X _147_/Y 0.016f
C8079 _182_/a_215_7# _298_/B 1.65e-20
C8080 _217_/a_27_7# _280_/a_68_257# 5.64e-19
C8081 _329_/a_27_7# _331_/CLK 0.212f
C8082 _268_/a_39_257# _315_/a_27_7# 7.83e-20
C8083 ctlp[1] _234_/B 4.18e-21
C8084 _216_/X _319_/D 1.57e-21
C8085 ctlp[3] clkbuf_2_1_0_clk/A 2.05e-19
C8086 _169_/B _196_/A 0.104f
C8087 _290_/A _273_/Y 0.00145f
C8088 trim[2] _273_/A 0.037f
C8089 _286_/B _336_/Q 0.0109f
C8090 _260_/A _191_/B 1.9e-19
C8091 _329_/Q _319_/D 1.05e-19
C8092 _346_/SET_B _340_/D 2.94e-19
C8093 _338_/Q _306_/S 2.93e-20
C8094 _172_/B VPWR 0.505f
C8095 _320_/a_27_7# _320_/a_543_7# -0.0117f
C8096 _320_/a_193_7# _320_/a_761_249# -0.0105f
C8097 _162_/X _300_/a_301_257# 0.0964f
C8098 _275_/A _306_/S 1.98e-19
C8099 _323_/a_193_7# _323_/a_448_7# -0.00297f
C8100 _157_/A _302_/a_323_257# 0.00129f
C8101 _304_/S _228_/A 0.822f
C8102 _267_/A _157_/a_27_7# 0.028f
C8103 _332_/a_1283_n19# _153_/a_215_257# 0.00151f
C8104 _332_/a_1108_7# _153_/a_109_53# 0.00104f
C8105 _149_/a_27_7# input1/X 2.08e-20
C8106 clkbuf_2_1_0_clk/A _299_/a_78_159# 0.00976f
C8107 _218_/a_250_257# _331_/D 6.8e-20
C8108 _336_/a_543_7# _194_/A 2.39e-20
C8109 _209_/X _332_/a_1283_n19# 1.93e-20
C8110 _254_/A _168_/a_109_7# 3.64e-20
C8111 _304_/a_591_329# _326_/Q 1.12e-19
C8112 _216_/A _313_/a_543_7# 0.0334f
C8113 _215_/A _162_/X 0.0073f
C8114 output18/a_27_7# _297_/B 0.00879f
C8115 ctln[7] _335_/a_1108_7# 0.0424f
C8116 _309_/a_27_7# _172_/B 4.81e-20
C8117 _258_/S _336_/a_543_7# 0.00112f
C8118 _277_/Y _162_/X 0.00875f
C8119 _279_/Y _242_/A 4.32e-20
C8120 _286_/B _336_/a_805_7# 2.96e-19
C8121 _339_/a_651_373# _195_/a_27_257# 8.98e-21
C8122 _339_/a_27_7# _194_/X 1.5e-19
C8123 _319_/a_1283_n19# _328_/Q 3.52e-19
C8124 _345_/a_796_7# _172_/B 5.54e-19
C8125 _307_/X _228_/A 9.6e-20
C8126 _312_/a_761_249# VPWR 0.038f
C8127 _312_/a_27_7# VGND 0.0663f
C8128 _346_/Q _147_/A 3.64e-20
C8129 _341_/D _255_/B 0.00485f
C8130 _309_/D _344_/Q 4.73e-21
C8131 _331_/Q _217_/A 0.0544f
C8132 _196_/A _314_/a_193_7# 0.00216f
C8133 _181_/X _314_/a_27_7# 1.63e-19
C8134 _308_/S _172_/A 0.0271f
C8135 _333_/D _225_/B 1.07e-20
C8136 _208_/a_78_159# _204_/Y 0.0101f
C8137 _208_/a_292_257# _335_/Q 0.00249f
C8138 _311_/a_1462_7# _311_/Q 5.79e-19
C8139 _307_/a_535_334# _250_/X 1.73e-19
C8140 _340_/a_1283_n19# _336_/a_761_249# 2.39e-21
C8141 _340_/a_543_7# _336_/a_543_7# 5.74e-21
C8142 _340_/a_1108_7# _336_/a_193_7# 5.24e-20
C8143 _346_/a_1602_7# _167_/a_109_257# 7.76e-21
C8144 _231_/a_79_n19# VGND 0.00284f
C8145 _231_/a_306_7# VPWR -3.26e-19
C8146 _216_/A _304_/S 0.0557f
C8147 _313_/a_805_7# _284_/A 4.25e-19
C8148 _325_/a_193_7# _286_/Y 0.0147f
C8149 _330_/Q _330_/a_651_373# 4.57e-19
C8150 _196_/A _170_/a_226_7# 3.39e-21
C8151 _315_/a_448_7# _177_/A 1.18e-20
C8152 _260_/B _336_/a_193_7# 1.05e-19
C8153 _326_/a_1108_7# _242_/A 0.0574f
C8154 _346_/a_1056_7# _167_/X 2.74e-19
C8155 input4/X _193_/Y 4.66e-19
C8156 _337_/Q _202_/a_584_7# 0.00174f
C8157 _318_/Q _271_/A 0.0154f
C8158 _180_/a_29_13# _283_/A 0.0125f
C8159 _302_/a_227_7# _303_/A 0.00222f
C8160 input3/a_27_7# valid 4.57e-20
C8161 _289_/a_121_257# VPWR -4.48e-19
C8162 _186_/a_382_257# _172_/A 5.78e-20
C8163 _149_/a_27_7# _286_/Y 1.44e-19
C8164 clkbuf_2_0_0_clk/a_75_172# _338_/a_27_7# 1.04e-20
C8165 _342_/Q _248_/A 2.37e-20
C8166 _281_/Y _331_/a_27_7# 3.99e-20
C8167 _330_/a_448_7# VPWR -0.00267f
C8168 _330_/a_1283_n19# VGND 0.0427f
C8169 _162_/X _304_/X 4.53e-21
C8170 _329_/a_1270_373# _346_/SET_B -2.06e-19
C8171 _320_/a_1283_n19# output19/a_27_7# 0.00844f
C8172 _344_/a_27_7# _171_/a_78_159# 2.45e-19
C8173 _251_/a_79_n19# _191_/B 1.02e-20
C8174 _183_/a_27_7# _324_/Q 0.00555f
C8175 _298_/C _298_/A 0.324f
C8176 _328_/a_1283_n19# _242_/A 1.77e-19
C8177 _306_/S _345_/D 7.68e-20
C8178 repeater43/a_27_7# _185_/A 8.12e-19
C8179 clk _324_/Q 0.0128f
C8180 _296_/Y _284_/A 0.0464f
C8181 _342_/Q _331_/CLK 0.0024f
C8182 _307_/X _216_/A 3.64e-20
C8183 _333_/a_27_7# VGND -0.0517f
C8184 _333_/a_761_249# VPWR 0.00955f
C8185 _337_/Q _260_/A 7.62e-21
C8186 _274_/a_39_257# _319_/D 6.66e-21
C8187 _297_/A _315_/D 0.0102f
C8188 _194_/X _313_/a_651_373# 3.84e-22
C8189 output13/a_27_7# _283_/Y 0.0192f
C8190 _341_/a_193_7# _341_/Q -2e-19
C8191 _342_/Q _190_/A 0.15f
C8192 _252_/a_27_7# VPWR 0.00121f
C8193 _337_/a_1217_7# _194_/X 1.32e-19
C8194 output22/a_27_7# _315_/a_27_7# 1.72e-19
C8195 _319_/Q _331_/a_193_7# 4.7e-20
C8196 _192_/B _336_/D 1.06e-21
C8197 _211_/a_373_7# _153_/B 0.00164f
C8198 _255_/B _143_/a_27_7# 0.00487f
C8199 _292_/Y _273_/A 0.0576f
C8200 _334_/a_1283_n19# _335_/Q 3.19e-20
C8201 _329_/D _331_/a_27_7# 1.87e-19
C8202 _271_/A _241_/a_199_7# 6.99e-19
C8203 _308_/S _203_/a_80_n19# 1.85e-19
C8204 _314_/a_1108_7# _347_/a_27_7# 9.74e-20
C8205 _314_/a_1283_n19# _347_/a_193_7# 3.66e-19
C8206 _162_/a_27_7# _344_/Q 4.97e-21
C8207 _254_/A _306_/S 0.00736f
C8208 clkbuf_0_clk/a_110_7# _284_/A 0.229f
C8209 _338_/Q _283_/A 2.07e-19
C8210 _325_/a_761_249# _284_/A 4.53e-21
C8211 _337_/Q _261_/A 1.88e-20
C8212 _281_/Y _145_/A 1.17e-20
C8213 ctlp[2] VGND 0.207f
C8214 _170_/a_226_7# _347_/a_1283_n19# 1.06e-20
C8215 _170_/a_76_159# _347_/a_1108_7# 4.97e-20
C8216 _162_/X _300_/Y 0.0858f
C8217 _312_/a_1283_n19# _311_/a_1108_7# 1.85e-19
C8218 _312_/a_1108_7# _311_/a_1283_n19# 1.24e-20
C8219 _312_/a_651_373# _311_/a_761_249# 4.5e-21
C8220 _339_/Q _202_/a_584_7# 2.09e-19
C8221 _323_/a_193_7# _323_/D -0.00415f
C8222 _157_/A _303_/A 0.00157f
C8223 _332_/a_543_7# _154_/A 6.77e-19
C8224 _332_/a_1108_7# _153_/A 2.65e-19
C8225 _279_/Y _336_/Q 0.0109f
C8226 repeater43/X _296_/a_213_83# 3.16e-22
C8227 _345_/a_1602_7# _164_/Y 9.14e-20
C8228 _330_/D _330_/a_27_7# 0.149f
C8229 _329_/a_761_249# _327_/Q 4.42e-20
C8230 _329_/a_193_7# _212_/X 7.89e-20
C8231 _212_/X _328_/Q 0.398f
C8232 _344_/a_27_7# _344_/a_562_373# -0.0012f
C8233 _344_/a_193_7# _344_/a_381_7# -0.00218f
C8234 _318_/Q _330_/D 9.79e-21
C8235 _161_/Y _285_/Y 5.28e-19
C8236 _255_/B _343_/CLK 0.00148f
C8237 _275_/Y _312_/a_1283_n19# 5.22e-19
C8238 _339_/Q _260_/A 2.04e-20
C8239 _182_/a_510_7# VPWR -0.00126f
C8240 _153_/B _203_/a_209_7# 1.2e-19
C8241 _182_/a_297_257# VGND -0.00115f
C8242 _183_/a_27_7# _228_/A 0.149f
C8243 _309_/D _306_/S 0.0914f
C8244 _242_/A _316_/D 0.00803f
C8245 _254_/B _153_/B 2.64e-19
C8246 _219_/a_93_n19# _219_/a_250_257# -6.97e-22
C8247 _324_/a_1283_n19# _181_/X 0.0141f
C8248 _339_/a_1217_7# _194_/X 1.36e-19
C8249 _339_/a_639_7# _306_/S 0.00104f
C8250 _339_/a_448_7# _340_/D 0.00489f
C8251 _255_/B _307_/a_535_334# 3.37e-19
C8252 _342_/Q _307_/a_505_n19# 2.5e-20
C8253 clk _228_/A 5.23e-19
C8254 comp _345_/Q 1.36e-20
C8255 _312_/a_1217_7# VGND -5.03e-19
C8256 _160_/X _299_/a_215_7# 2.8e-20
C8257 _325_/Q _236_/B 2.87e-20
C8258 _319_/a_543_7# _319_/D 0.00226f
C8259 _346_/a_652_n19# _277_/A 1.94e-19
C8260 _288_/A VGND 0.45f
C8261 trimb[4] VPWR 0.183f
C8262 trim[1] VPWR 0.354f
C8263 _204_/Y _190_/A 0.00292f
C8264 _294_/A _254_/A 0.0358f
C8265 _347_/Q _347_/a_27_7# 1.73e-20
C8266 _299_/X _347_/a_193_7# 2.3e-19
C8267 _316_/a_27_7# _242_/B 1.46e-21
C8268 _258_/a_76_159# _313_/Q 0.00187f
C8269 _216_/X _227_/A 0.146f
C8270 _161_/Y _171_/a_493_257# 1.79e-19
C8271 _215_/A _298_/C 0.0193f
C8272 _254_/Y _338_/Q 1.44e-20
C8273 _255_/a_30_13# _192_/B 0.0572f
C8274 _162_/X VGND 0.519f
C8275 _246_/B _223_/a_250_257# 0.0675f
C8276 _342_/Q _178_/a_27_7# 3.13e-19
C8277 _326_/a_448_7# _326_/Q 0.00148f
C8278 _287_/a_39_257# VGND 0.0205f
C8279 _315_/D _177_/A 0.0235f
C8280 _313_/D _172_/A 8.69e-20
C8281 _339_/Q _261_/A 0.424f
C8282 repeater43/X _230_/a_27_7# 0.00268f
C8283 _177_/a_27_7# VPWR 0.124f
C8284 _318_/Q _232_/a_27_7# 3.6e-19
C8285 _279_/Y _314_/a_761_249# 0.0102f
C8286 _342_/a_1283_n19# _172_/A 1.11e-19
C8287 _260_/B _314_/a_1283_n19# 2.22e-19
C8288 _344_/a_27_7# _172_/B 0.0114f
C8289 _321_/D _321_/a_543_7# 7.69e-19
C8290 _343_/a_1283_n19# _298_/X 3.22e-20
C8291 _321_/a_651_373# _331_/CLK 8.49e-19
C8292 _280_/a_68_257# _281_/A 0.00142f
C8293 clk _216_/A 0.0059f
C8294 _346_/SET_B _310_/a_805_7# 6.41e-19
C8295 _320_/a_193_7# output18/a_27_7# 2.53e-20
C8296 _165_/X _172_/a_109_257# 1.07e-21
C8297 _309_/a_761_249# _162_/X 3.53e-22
C8298 _333_/a_1217_7# VGND -4.7e-19
C8299 repeater43/X _232_/A 0.147f
C8300 _294_/Y _267_/B 0.00184f
C8301 _294_/A _309_/D 0.23f
C8302 _276_/a_68_257# _319_/Q 0.0294f
C8303 _211_/a_109_257# _197_/X 4.9e-19
C8304 _337_/Q _340_/Q 0.0378f
C8305 _299_/a_493_257# VGND -1.65e-19
C8306 _315_/Q _315_/a_651_373# 1.4e-19
C8307 result[0] _315_/a_1108_7# 0.00279f
C8308 clk _251_/a_510_7# 7.21e-20
C8309 _343_/a_193_7# _298_/C 1.86e-20
C8310 _343_/a_651_373# _176_/a_27_7# 2.42e-19
C8311 _343_/a_543_7# _343_/Q 5.56e-19
C8312 _197_/X _198_/a_250_257# 0.0109f
C8313 _315_/D _347_/a_761_249# 2.36e-19
C8314 _346_/SET_B _265_/B 0.599f
C8315 _174_/a_109_7# _344_/D 8.6e-19
C8316 repeater43/X _234_/a_109_257# 5.77e-19
C8317 _334_/Q _205_/a_79_n19# 2.19e-19
C8318 repeater43/X _321_/a_27_7# 0.0158f
C8319 _305_/a_505_n19# _254_/B 0.0486f
C8320 _297_/B _347_/a_27_7# 0.111f
C8321 _268_/a_121_257# VPWR 3.16e-19
C8322 repeater43/X rstn 0.647f
C8323 _227_/A _334_/a_193_7# 1.47e-19
C8324 _312_/a_543_7# _311_/D 2.04e-21
C8325 _191_/B _205_/a_79_n19# 0.0311f
C8326 _341_/D _315_/a_1283_n19# 1.61e-19
C8327 _171_/a_215_7# _172_/B 6.58e-19
C8328 _175_/Y _226_/a_79_n19# 0.0617f
C8329 clkbuf_2_3_0_clk/A _319_/D 3.67e-20
C8330 _341_/a_27_7# VPWR 0.089f
C8331 _305_/X VPWR 0.165f
C8332 _342_/a_1283_n19# _244_/B 5.84e-19
C8333 _202_/a_584_7# _336_/D 4.76e-20
C8334 _214_/a_373_7# _331_/D 7.87e-19
C8335 _292_/A output37/a_27_7# 1.51e-19
C8336 _338_/a_27_7# VPWR 0.015f
C8337 _319_/Q _219_/a_93_n19# 4.2e-20
C8338 _281_/Y _324_/Q 2.77e-19
C8339 _206_/A _153_/a_215_257# 0.0121f
C8340 _225_/B _190_/A 0.0272f
C8341 _339_/a_639_7# _283_/A 0.00422f
C8342 _346_/SET_B _336_/a_1270_373# -9.44e-20
C8343 _209_/X _206_/A 7.21e-20
C8344 _319_/D _327_/Q 3.48e-21
C8345 _236_/B _326_/Q 2.68e-19
C8346 _346_/SET_B _314_/a_27_7# -2.33e-19
C8347 output34/a_27_7# VPWR 0.13f
C8348 _339_/D _340_/D 0.188f
C8349 _339_/Q _340_/Q 0.0406f
C8350 _294_/A _162_/a_27_7# 7.51e-19
C8351 _342_/Q _296_/Y 1.06e-19
C8352 _308_/a_76_159# _333_/D 6.33e-20
C8353 _188_/a_218_334# _298_/A 0.00243f
C8354 rstn _334_/Q 0.00116f
C8355 _254_/Y _254_/A 0.531f
C8356 _317_/Q _317_/a_193_7# 0.00171f
C8357 _260_/A _336_/D 8.04e-20
C8358 _246_/a_109_257# _330_/a_193_7# 6.05e-20
C8359 _230_/a_27_7# _317_/a_543_7# 2.4e-19
C8360 _298_/B _180_/a_29_13# 0.00453f
C8361 _340_/a_761_249# VPWR 0.0141f
C8362 _340_/a_27_7# VGND -0.0668f
C8363 _346_/SET_B _170_/a_76_159# 5.1e-20
C8364 _193_/Y _202_/a_93_n19# 0.0311f
C8365 _306_/S _202_/a_250_257# 9.52e-20
C8366 _320_/Q _330_/Q 0.0456f
C8367 _326_/D _326_/Q 0.0135f
C8368 _327_/a_193_7# _330_/Q 0.00145f
C8369 _283_/A _331_/a_1108_7# 0.00797f
C8370 _316_/a_193_7# VPWR 0.0405f
C8371 _343_/a_761_249# _229_/a_226_7# 8.29e-19
C8372 _343_/a_193_7# _229_/a_489_373# 1.66e-20
C8373 _343_/a_543_7# _229_/a_76_159# 1.76e-19
C8374 _279_/Y _324_/a_448_7# 5.5e-21
C8375 _251_/a_297_257# _286_/Y 3.02e-19
C8376 _309_/a_448_7# _286_/B 8.66e-20
C8377 _227_/A _332_/Q 2.7e-19
C8378 cal _193_/Y 1.59f
C8379 _216_/X _297_/B 0.286f
C8380 _221_/a_256_7# _286_/Y 0.00429f
C8381 input1/X _306_/S 0.017f
C8382 rstn _191_/B -1.32e-38
C8383 _242_/A _331_/a_27_7# 2.76e-20
C8384 _326_/a_193_7# _330_/Q 6.53e-21
C8385 _326_/Q _222_/a_256_7# 4.83e-19
C8386 _313_/a_27_7# _336_/Q 5.23e-20
C8387 _342_/Q clkbuf_0_clk/a_110_7# 0.0102f
C8388 _327_/a_27_7# VPWR 0.0767f
C8389 clkbuf_2_1_0_clk/A _346_/SET_B 0.044f
C8390 _317_/a_543_7# _232_/A 6.72e-19
C8391 _317_/a_761_249# _248_/B 4.95e-21
C8392 _335_/D _333_/a_193_7# 1.05e-20
C8393 _197_/a_27_7# _193_/Y 1.23e-19
C8394 _329_/Q _297_/B 0.208f
C8395 _298_/C VGND 0.766f
C8396 _250_/a_292_257# _216_/A 0.00443f
C8397 _326_/a_27_7# VPWR 0.0674f
C8398 _322_/a_27_7# _322_/Q 5.9e-19
C8399 _346_/SET_B _310_/Q 0.0176f
C8400 _254_/Y _309_/D 3.67e-20
C8401 _328_/a_27_7# _330_/Q 3.78e-20
C8402 _342_/D _188_/S 6.6e-20
C8403 _281_/Y _281_/A 0.136f
C8404 ctlp[7] _271_/A 2.67e-20
C8405 _329_/a_1108_7# clkbuf_0_clk/X 0.00607f
C8406 clkbuf_0_clk/X _327_/D 0.00393f
C8407 _332_/a_1270_373# VPWR -2.18e-19
C8408 _332_/a_448_7# VGND 0.00146f
C8409 _331_/Q _214_/a_109_257# 0.00133f
C8410 _300_/a_735_7# _346_/SET_B 0.00223f
C8411 _338_/Q _284_/a_39_257# 2.21e-22
C8412 _347_/a_651_373# VGND 0.00132f
C8413 _347_/a_639_7# VPWR 5.41e-19
C8414 _200_/a_346_7# VPWR -7.53e-19
C8415 _200_/a_250_257# VGND -0.0043f
C8416 _326_/a_639_7# _304_/X 6.64e-19
C8417 _194_/X _267_/A 0.00631f
C8418 _281_/Y _228_/A 0.706f
C8419 _207_/C _298_/A 5.84e-20
C8420 _217_/a_27_7# _242_/A 6.32e-20
C8421 _191_/B _225_/a_59_35# 0.00115f
C8422 repeater43/X _321_/a_1217_7# -2.1e-19
C8423 _328_/a_193_7# _297_/B 0.00124f
C8424 _314_/Q _347_/a_448_7# 0.0018f
C8425 _314_/D _347_/a_805_7# 1.02e-20
C8426 _306_/S _286_/Y 0.0667f
C8427 _265_/B _147_/A 8.84e-20
C8428 _263_/B _311_/D 0.0426f
C8429 _341_/Q _226_/a_79_n19# 6.41e-21
C8430 output28/a_27_7# _242_/A 1.57e-20
C8431 _216_/a_27_7# _227_/A 0.024f
C8432 _329_/D _281_/A 0.011f
C8433 _346_/a_27_7# _160_/X 7.93e-20
C8434 _346_/a_476_7# _347_/Q 3.08e-19
C8435 _217_/A _347_/D 7.77e-20
C8436 _251_/a_215_7# _284_/A 0.00368f
C8437 _343_/CLK _315_/a_1283_n19# 0.0278f
C8438 _294_/A input1/X 0.0503f
C8439 ctln[6] _207_/a_27_7# 0.00185f
C8440 _175_/Y _323_/Q 0.0233f
C8441 _165_/a_215_7# VGND 0.0284f
C8442 _344_/a_652_n19# _162_/X 9.28e-20
C8443 _239_/a_199_7# _240_/B -2.22e-34
C8444 clkbuf_0_clk/X _283_/A 0.00229f
C8445 _254_/A _336_/a_1108_7# 2.31e-19
C8446 _167_/X _267_/A 2.15e-19
C8447 _341_/a_639_7# VGND -0.00153f
C8448 _341_/a_1217_7# VPWR 1.18e-19
C8449 _179_/a_27_7# _333_/a_1108_7# 1.56e-20
C8450 _174_/a_27_257# _297_/Y 1.01e-20
C8451 _184_/a_218_7# _182_/X 8.05e-19
C8452 _325_/a_543_7# _242_/A 2.46e-21
C8453 _338_/a_639_7# VGND 4.72e-19
C8454 _338_/a_1217_7# VPWR 6.07e-20
C8455 _331_/D _330_/a_543_7# 1.89e-19
C8456 _314_/a_27_7# _156_/a_39_257# 0.00214f
C8457 _281_/Y _216_/A 0.0139f
C8458 _330_/a_193_7# _330_/a_543_7# -0.0129f
C8459 _316_/Q _316_/a_1283_n19# 0.0844f
C8460 ctln[3] output34/a_27_7# 2.08e-19
C8461 output9/a_27_7# trim[3] 2.75e-19
C8462 _338_/Q _262_/a_113_257# 0.0146f
C8463 _290_/A _344_/D 5.95e-20
C8464 _196_/A _153_/B 0.00125f
C8465 _325_/a_1283_n19# _325_/Q 0.00146f
C8466 _328_/a_1108_7# _279_/A 3.48e-21
C8467 _346_/SET_B _314_/a_1217_7# 3.36e-21
C8468 _304_/S _224_/a_93_n19# 1.77e-19
C8469 _321_/a_27_7# result[6] 0.00217f
C8470 _315_/D _248_/A 0.294f
C8471 _150_/C _298_/A 0.124f
C8472 _271_/A _316_/a_448_7# 3.94e-21
C8473 _172_/B _147_/Y 3.5e-20
C8474 _290_/A _346_/Q 5.85e-21
C8475 _343_/CLK _154_/A 1.24e-19
C8476 _229_/a_556_7# VPWR -5.97e-19
C8477 _229_/a_489_373# VGND 6.2e-19
C8478 _295_/a_676_257# VPWR -4.89e-19
C8479 clkbuf_0_clk/X _248_/B 0.0686f
C8480 _346_/a_193_7# VPWR 0.0265f
C8481 _337_/Q _310_/a_448_7# 0.00121f
C8482 _340_/a_1217_7# VGND -4.9e-19
C8483 _340_/Q _336_/D 1.84e-19
C8484 _193_/Y _284_/A 0.0607f
C8485 _321_/D _318_/D 0.218f
C8486 _331_/CLK _315_/D 4.64e-20
C8487 input1/X _283_/A 0.0105f
C8488 _335_/a_193_7# _208_/a_78_159# 0.00913f
C8489 _277_/Y clkbuf_2_2_0_clk/a_75_172# 0.00599f
C8490 _239_/a_199_7# _328_/Q 0.00126f
C8491 _316_/a_805_7# VGND -6.33e-19
C8492 _316_/a_1462_7# VPWR 9.93e-20
C8493 _273_/A output37/a_27_7# 0.015f
C8494 _346_/SET_B _278_/a_68_257# 7.07e-21
C8495 _345_/a_1032_373# _346_/SET_B -8.05e-19
C8496 _344_/a_1032_373# _164_/Y 0.0157f
C8497 _300_/a_301_257# _313_/a_1283_n19# 2.19e-20
C8498 _324_/a_651_373# _331_/CLK 4.9e-20
C8499 _346_/a_476_7# _297_/B 4.24e-20
C8500 _331_/a_193_7# _326_/Q 2.79e-21
C8501 _277_/Y input4/X 2.99e-20
C8502 _327_/D _286_/Y 0.12f
C8503 cal _205_/a_297_7# 3.62e-19
C8504 _315_/Q _316_/Q 0.0449f
C8505 _313_/a_1217_7# _336_/Q 3.05e-20
C8506 _273_/A _315_/D 0.19f
C8507 _327_/a_639_7# VGND -0.00134f
C8508 _327_/a_1217_7# VPWR 4.39e-19
C8509 repeater43/X _315_/a_805_7# 6.21e-19
C8510 _195_/a_109_7# _340_/D 3.22e-19
C8511 _277_/Y _345_/Q 0.0122f
C8512 _225_/X _153_/A 2.05e-19
C8513 _326_/a_1217_7# VPWR 1.91e-20
C8514 _326_/a_639_7# VGND 9.99e-19
C8515 _215_/A _313_/a_1283_n19# 0.0267f
C8516 clk _153_/a_109_53# 1.87e-20
C8517 _254_/A _300_/a_27_257# 3.98e-21
C8518 repeater43/X _324_/a_27_7# -0.00149f
C8519 clkbuf_2_1_0_clk/A _147_/A 0.00775f
C8520 _345_/a_27_7# _158_/Y 1.11e-19
C8521 _227_/A _327_/Q 0.00266f
C8522 _218_/a_93_n19# _346_/SET_B 0.00281f
C8523 _332_/a_543_7# _153_/B 0.0148f
C8524 _180_/a_111_257# VPWR -4.77e-19
C8525 _254_/A _194_/a_27_7# 8.71e-21
C8526 _332_/D VGND 0.0812f
C8527 _331_/Q _331_/D 0.101f
C8528 _301_/X _301_/a_240_7# 0.00298f
C8529 trim[0] _312_/Q 3.54e-20
C8530 rstn _339_/Q 2.67e-20
C8531 _331_/Q _330_/a_193_7# 3.24e-19
C8532 _328_/a_805_7# VPWR 2.79e-19
C8533 _328_/a_1270_373# VGND 4.74e-20
C8534 _173_/a_76_159# VPWR 0.00547f
C8535 _275_/A _160_/X 1.79e-20
C8536 _147_/A _310_/Q 4.96e-19
C8537 _326_/D _324_/D 1.44e-20
C8538 _283_/A _286_/Y 0.0085f
C8539 _194_/A _311_/D 1.93e-19
C8540 _305_/a_505_n19# _196_/A 0.00742f
C8541 _181_/X _214_/a_109_7# 2.97e-20
C8542 _271_/A _334_/a_1283_n19# 0.0396f
C8543 _319_/a_193_7# VPWR 0.0487f
C8544 _346_/SET_B _311_/a_27_7# 0.0211f
C8545 _328_/a_1462_7# _297_/B 4.37e-19
C8546 _321_/a_805_7# result[7] 2.89e-20
C8547 _314_/Q _347_/D 0.0321f
C8548 _217_/A _222_/a_584_7# 6.38e-19
C8549 output35/a_27_7# VGND 0.0309f
C8550 _335_/a_27_7# _334_/a_1283_n19# 1.91e-21
C8551 _300_/a_735_7# _147_/A 1.58e-20
C8552 _337_/Q _336_/a_1283_n19# 3.1e-19
C8553 _254_/Y input1/X 0.472f
C8554 _216_/X _320_/a_193_7# 1.87e-20
C8555 _258_/S _311_/D 0.00317f
C8556 _258_/S _258_/a_505_n19# 0.0422f
C8557 _319_/a_543_7# _297_/B 1.66e-19
C8558 _334_/a_805_7# VPWR 3.7e-19
C8559 clk _209_/a_27_257# 0.00596f
C8560 clkbuf_0_clk/a_110_7# _225_/B 0.00123f
C8561 _167_/a_27_257# _346_/Q 0.0383f
C8562 _301_/a_51_257# _267_/A 1.16e-20
C8563 ctln[1] _227_/A 2.32e-20
C8564 _309_/a_543_7# _340_/CLK 4.37e-20
C8565 _312_/Q _311_/Q 0.00599f
C8566 _308_/X _182_/X 0.00496f
C8567 _320_/Q _320_/a_761_249# 5.48e-19
C8568 _329_/Q _320_/a_193_7# 2.36e-20
C8569 _216_/a_27_7# _297_/B 1.46e-19
C8570 _345_/a_652_n19# _345_/D 0.00167f
C8571 _345_/a_476_7# _345_/Q 9.67e-19
C8572 _215_/A _150_/C 2.56e-19
C8573 output26/a_27_7# _242_/A 5.76e-20
C8574 _248_/B _286_/Y 0.1f
C8575 _324_/a_543_7# _304_/S 0.0356f
C8576 _325_/a_1283_n19# _326_/Q 0.00758f
C8577 _344_/Q clkc 1.11e-19
C8578 input1/a_75_172# _199_/a_93_n19# 6.84e-20
C8579 _227_/A _192_/B 0.599f
C8580 clkbuf_2_3_0_clk/A _347_/Q 7.03e-20
C8581 _197_/X _312_/D 2.62e-20
C8582 _329_/a_805_7# _281_/A 0.00259f
C8583 _329_/a_651_373# _281_/Y 0.00112f
C8584 _183_/a_471_7# _298_/A 0.0033f
C8585 clkbuf_2_0_0_clk/a_75_172# _337_/Q 1.76e-21
C8586 clkbuf_2_1_0_clk/A _337_/D 1.56e-19
C8587 _304_/S _217_/A 0.00195f
C8588 _340_/a_193_7# _198_/a_250_257# 1.17e-19
C8589 _340_/a_761_249# _198_/a_93_n19# 4.94e-20
C8590 _342_/a_1283_n19# _177_/A 8.8e-20
C8591 _271_/A _316_/D 0.136f
C8592 clk input3/a_27_7# 0.00295f
C8593 _188_/a_218_7# VPWR -3.66e-19
C8594 _188_/a_218_334# VGND -6.97e-19
C8595 _342_/a_27_7# valid 0.00356f
C8596 _325_/a_27_7# _227_/A 0.00157f
C8597 _346_/a_1140_373# VGND 3.13e-19
C8598 _337_/Q _310_/D 0.00992f
C8599 _160_/X _345_/D 0.0985f
C8600 _333_/a_193_7# _333_/a_448_7# -0.00779f
C8601 _335_/a_543_7# _332_/Q 2.63e-19
C8602 _275_/A repeater42/a_27_7# 5.02e-20
C8603 clkbuf_0_clk/a_110_7# _314_/a_543_7# 2.35e-20
C8604 _309_/a_1283_n19# _346_/SET_B -0.0131f
C8605 _335_/a_1283_n19# _207_/X 0.0658f
C8606 _342_/a_193_7# _343_/Q 6.78e-21
C8607 _343_/a_193_7# _150_/C 1.86e-20
C8608 _343_/a_543_7# _147_/A 7.33e-22
C8609 _343_/a_27_7# _226_/X 1.01e-19
C8610 _329_/a_1270_373# _319_/Q 6.24e-19
C8611 output26/a_27_7# _322_/D 0.0355f
C8612 _160_/X _313_/a_1108_7# 1.07e-20
C8613 _150_/C _304_/X 8.22e-20
C8614 _328_/a_448_7# _328_/D 0.00355f
C8615 _239_/a_113_257# _319_/D 1.03e-19
C8616 repeater43/a_27_7# _271_/A 2.5e-19
C8617 _323_/a_1283_n19# _334_/a_27_7# 1.4e-20
C8618 _200_/a_584_7# _311_/D 1.25e-19
C8619 _329_/a_651_373# _329_/D 8.49e-19
C8620 _283_/Y _338_/a_1108_7# 0.00237f
C8621 _257_/a_222_53# _216_/A 1.09e-21
C8622 _321_/D _318_/a_448_7# 0.00922f
C8623 _326_/a_1108_7# _232_/a_27_7# 4.49e-19
C8624 _342_/Q _251_/a_215_7# 0.00504f
C8625 ctln[6] _283_/A 0.277f
C8626 clkbuf_2_2_0_clk/a_75_172# VGND 0.0676f
C8627 output33/a_27_7# clkc 0.00593f
C8628 trim[2] output5/a_27_7# 1.32e-19
C8629 _321_/Q _327_/Q 7.32e-20
C8630 cal _298_/A 0.0358f
C8631 input4/X VGND 0.184f
C8632 clk _153_/A 0.0202f
C8633 repeater43/X VPWR 1.97f
C8634 _254_/A _160_/X 0.333f
C8635 _312_/a_193_7# _312_/D 0.00637f
C8636 repeater43/X _324_/a_1217_7# -3.08e-19
C8637 _317_/a_27_7# _217_/A 1.58e-21
C8638 input1/X _336_/a_1108_7# 0.0522f
C8639 clkbuf_2_3_0_clk/A _297_/B 0.0258f
C8640 _315_/D _217_/X 6.53e-19
C8641 _288_/Y VPWR 0.054f
C8642 _288_/A output40/a_27_7# 1.21e-19
C8643 output32/a_27_7# _288_/A 0.0328f
C8644 _324_/a_639_7# _327_/Q 1.67e-19
C8645 repeater43/X _318_/a_543_7# 0.0343f
C8646 _343_/a_805_7# repeater43/X 5.41e-19
C8647 _161_/Y _162_/A 0.00403f
C8648 _316_/a_27_7# _244_/B 0.019f
C8649 _345_/Q VGND 0.496f
C8650 _329_/a_27_7# _329_/a_448_7# -0.00642f
C8651 _329_/a_193_7# _329_/a_1108_7# -0.00817f
C8652 _329_/a_193_7# _327_/D 2.69e-20
C8653 _328_/Q _327_/D 0.0034f
C8654 _279_/Y _283_/Y 2.04e-19
C8655 clkbuf_2_0_0_clk/a_75_172# _339_/Q 2.5e-21
C8656 _313_/Q _194_/A 4.83e-19
C8657 _297_/B _327_/Q 1.04e-19
C8658 _207_/C VGND 2.92f
C8659 _331_/a_1283_n19# _304_/X 7.68e-19
C8660 _260_/A _260_/a_27_257# 0.044f
C8661 _317_/D valid 5.36e-19
C8662 _175_/Y sample 1.66e-19
C8663 _319_/a_1462_7# VPWR 1.04e-19
C8664 _319_/a_805_7# VGND 0.00227f
C8665 _313_/a_1283_n19# VGND 0.0363f
C8666 _313_/a_448_7# VPWR -0.00348f
C8667 _323_/a_193_7# _248_/A 2.3e-20
C8668 _346_/SET_B _328_/D 0.05f
C8669 _181_/X _330_/a_761_249# 1.13e-19
C8670 _346_/SET_B _311_/a_1217_7# 2.37e-19
C8671 _337_/a_805_7# VPWR 1.67e-19
C8672 _337_/a_1270_373# VGND 4.37e-20
C8673 _297_/B _172_/Y 0.0134f
C8674 _342_/a_1283_n19# _341_/a_1283_n19# 0.00144f
C8675 _342_/a_1108_7# _341_/a_543_7# 5.16e-21
C8676 _342_/a_651_373# _341_/a_193_7# 5.06e-22
C8677 output9/a_27_7# _343_/CLK 4.03e-19
C8678 _298_/C _203_/a_209_257# 8.23e-19
C8679 output15/a_27_7# _233_/a_113_257# 2.77e-20
C8680 _339_/Q _310_/D 2.65e-21
C8681 _189_/a_27_7# _340_/D 8e-21
C8682 _258_/S _313_/Q 0.0874f
C8683 _231_/a_676_257# _177_/A 1.8e-21
C8684 output21/a_27_7# _331_/Q 4.33e-21
C8685 _320_/Q _322_/a_448_7# 0.0289f
C8686 _334_/Q VPWR 1.03f
C8687 _255_/X _306_/S 8.48e-20
C8688 _296_/Y _315_/D 0.0249f
C8689 _257_/a_448_7# _306_/S 6.06e-19
C8690 _315_/a_27_7# _286_/Y 1.12e-20
C8691 _345_/a_1224_7# _345_/Q 8.54e-19
C8692 _272_/a_39_257# _317_/a_193_7# 1.76e-20
C8693 _167_/X _301_/a_51_257# 0.00643f
C8694 _308_/X _229_/a_226_7# 3.82e-21
C8695 output22/a_27_7# _244_/B 0.00107f
C8696 _308_/S _190_/A 0.00184f
C8697 _329_/a_193_7# _283_/A 6.28e-21
C8698 _167_/X clkbuf_1_1_0_clk/a_75_172# 9.92e-19
C8699 _216_/A _242_/A 1.94e-19
C8700 _172_/A _295_/a_79_n19# 8.12e-19
C8701 _342_/a_193_7# _229_/a_76_159# 6.07e-19
C8702 _342_/a_27_7# _229_/a_226_7# 1.33e-19
C8703 _346_/a_27_7# _172_/A 1.08e-20
C8704 _210_/a_109_257# _306_/S 8.37e-19
C8705 _319_/Q _234_/B 0.486f
C8706 _191_/B VPWR 1.65f
C8707 _304_/S _314_/Q 3.55e-20
C8708 _319_/Q _321_/a_1283_n19# 0.00132f
C8709 _184_/a_76_159# _226_/a_79_n19# 6.4e-19
C8710 _337_/Q _266_/a_113_257# 6.92e-20
C8711 _218_/a_250_257# _331_/a_193_7# 4.91e-20
C8712 _340_/a_448_7# _197_/X 1.22e-19
C8713 _298_/B input1/X 0.0057f
C8714 _157_/A _227_/A 0.00964f
C8715 clkbuf_0_clk/a_110_7# _315_/D 3.35e-20
C8716 _218_/a_584_7# _212_/X 7.26e-19
C8717 _218_/a_346_7# _217_/X 3.77e-20
C8718 _150_/C VGND 0.612f
C8719 _246_/B _212_/X 0.00626f
C8720 _342_/D output41/a_27_7# 1.1e-21
C8721 _302_/a_77_159# _300_/Y 0.0428f
C8722 _324_/a_193_7# clkbuf_0_clk/X 0.00133f
C8723 _325_/a_1217_7# _227_/A 3.05e-20
C8724 _232_/a_27_7# _316_/D 1.75e-19
C8725 input1/X _194_/a_27_7# 1.95e-20
C8726 _283_/Y _334_/a_1283_n19# 7.12e-22
C8727 _157_/A _314_/a_1108_7# 0.00222f
C8728 _333_/a_193_7# _333_/D 0.0123f
C8729 _293_/a_39_257# _346_/SET_B 5.38e-20
C8730 _320_/a_761_249# _319_/a_761_249# 4.11e-21
C8731 _320_/a_1283_n19# _319_/a_27_7# 4.58e-20
C8732 _320_/a_27_7# _319_/a_1283_n19# 5.66e-20
C8733 _344_/a_27_7# _173_/a_76_159# 1.2e-19
C8734 _248_/B _328_/Q 5.99e-19
C8735 _343_/a_1217_7# _226_/X 3.56e-20
C8736 _339_/a_805_7# VPWR 2.83e-19
C8737 _339_/a_1270_373# VGND 4.82e-20
C8738 _341_/a_1270_373# _317_/D 1.37e-19
C8739 _327_/a_805_7# _232_/X 3.28e-19
C8740 _325_/a_448_7# _217_/A 0.018f
C8741 _277_/Y cal 2.67e-19
C8742 _317_/a_543_7# VPWR 0.011f
C8743 _317_/a_193_7# VGND 0.00192f
C8744 _294_/Y _297_/Y 3.68e-19
C8745 _275_/Y clkbuf_2_3_0_clk/A 0.00289f
C8746 _294_/A clkc 1.14f
C8747 _298_/A _284_/A 6.46e-21
C8748 _182_/a_297_257# _286_/B 5.66e-20
C8749 _182_/a_79_n19# _196_/A 0.0411f
C8750 _169_/B _344_/D 3.12e-20
C8751 _326_/a_805_7# _232_/X 1.8e-19
C8752 repeater43/X _335_/a_1108_7# -0.00674f
C8753 _172_/a_109_257# VPWR -0.00157f
C8754 _330_/Q _331_/a_651_373# 0.00267f
C8755 _330_/Q result[7] 4.39e-19
C8756 _258_/S _312_/a_1283_n19# 5.3e-22
C8757 _318_/a_1108_7# _317_/a_193_7# 3.15e-21
C8758 _169_/B _346_/Q 9.77e-21
C8759 _292_/A _312_/a_193_7# 1.64e-19
C8760 _285_/A _338_/Q 1.15e-20
C8761 _188_/S _180_/a_183_257# 5.74e-19
C8762 _285_/A _275_/A 7.33e-20
C8763 _309_/a_193_7# _309_/D 0.0035f
C8764 _308_/S _307_/a_505_n19# 0.0106f
C8765 _229_/a_226_7# _317_/D 1.18e-19
C8766 _328_/a_639_7# _232_/X 2.02e-19
C8767 _331_/a_1283_n19# VGND 0.0248f
C8768 _331_/a_448_7# VPWR 0.00308f
C8769 _298_/B _286_/Y 0.229f
C8770 _275_/Y _172_/Y 0.0126f
C8771 _286_/B _162_/X 0.161f
C8772 _169_/B _168_/a_481_7# 1.48e-19
C8773 _294_/Y _310_/a_193_7# 1.03e-20
C8774 _302_/a_77_159# VGND 0.0164f
C8775 _302_/a_323_257# VPWR -0.00138f
C8776 _214_/a_109_7# _346_/SET_B 6.83e-20
C8777 _324_/a_27_7# _303_/A 3.11e-22
C8778 _344_/a_1182_221# _346_/SET_B -0.00733f
C8779 _269_/A _248_/B 0.00141f
C8780 _316_/a_639_7# _317_/D 0.00104f
C8781 _343_/a_193_7# cal 0.0082f
C8782 _163_/a_78_159# _161_/Y 7.99e-20
C8783 output24/a_27_7# _232_/A 4.46e-21
C8784 _308_/S _178_/a_27_7# 2.57e-19
C8785 _336_/a_761_249# _340_/Q 2.9e-21
C8786 _336_/a_193_7# _306_/S 0.013f
C8787 _336_/a_27_7# _193_/Y 2.02e-19
C8788 _154_/a_27_7# _333_/Q 3.7e-19
C8789 _302_/a_227_7# _297_/B 0.00896f
C8790 _292_/A _289_/a_39_257# 0.0132f
C8791 _260_/A _314_/a_1108_7# 2.38e-20
C8792 ctln[7] _333_/Q 1.41e-20
C8793 _304_/a_306_329# _162_/X 1.16e-19
C8794 _157_/A _347_/Q 9.22e-20
C8795 _335_/a_639_7# _334_/D 2.38e-19
C8796 _335_/a_1108_7# _334_/Q 0.00129f
C8797 _337_/Q VPWR 1.53f
C8798 _342_/a_761_249# _341_/D 2.8e-21
C8799 _325_/a_193_7# _246_/B 4.89e-21
C8800 _342_/D _341_/a_761_249# 1.08e-20
C8801 _290_/A _265_/B 0.153f
C8802 _322_/a_543_7# _331_/CLK 4.44e-20
C8803 _270_/a_39_257# _232_/A 0.015f
C8804 _255_/X _283_/A 8.46e-21
C8805 _145_/A _271_/A 0.00677f
C8806 ctln[1] _335_/a_543_7# 4.86e-19
C8807 ctlp[1] _322_/Q 0.00105f
C8808 _179_/a_27_7# _333_/Q 0.0127f
C8809 _321_/a_193_7# _269_/A 3.36e-20
C8810 _301_/X _346_/D 0.181f
C8811 _271_/A output28/a_27_7# 2.93e-19
C8812 _280_/a_68_257# _217_/A 3.24e-20
C8813 _343_/CLK _153_/B 6.44e-20
C8814 _216_/A _336_/Q 4.26e-20
C8815 _275_/A _172_/A 4.25e-19
C8816 _283_/Y repeater43/a_27_7# 0.00174f
C8817 output13/a_27_7# input4/X 0.0332f
C8818 _271_/A _146_/a_112_13# 2.59e-20
C8819 _250_/a_493_257# _215_/A 0.00102f
C8820 result[6] VPWR 0.435f
C8821 _324_/a_193_7# _286_/Y 0.0143f
C8822 _340_/CLK _254_/B 0.381f
C8823 _306_/a_505_n19# _309_/D 5.76e-20
C8824 _275_/A _232_/X 0.0173f
C8825 _320_/Q _330_/a_1270_373# 3.5e-19
C8826 _342_/a_1283_n19# _248_/A 0.00131f
C8827 _309_/a_27_7# _337_/Q 0.00945f
C8828 _284_/a_121_257# _284_/A 9.5e-19
C8829 _346_/Q _170_/a_226_7# 8.99e-19
C8830 _281_/Y _153_/A 3.61e-21
C8831 result[6] _318_/a_543_7# 4.92e-20
C8832 repeater43/X _323_/a_1108_7# 0.00625f
C8833 _343_/a_27_7# _286_/Y 0.0131f
C8834 _313_/D _190_/A 4.95e-20
C8835 _188_/S _226_/a_79_n19# 1.55e-19
C8836 _184_/a_535_334# _150_/C 1.68e-19
C8837 _330_/D _331_/a_27_7# 0.0017f
C8838 _301_/a_240_7# _297_/Y 2.33e-19
C8839 _320_/a_27_7# _212_/X 2.2e-21
C8840 _313_/Q _201_/a_27_7# 4.85e-21
C8841 _294_/A _336_/a_193_7# 1.85e-20
C8842 _158_/Y _285_/Y 2.78e-21
C8843 _183_/a_471_7# VGND -0.0233f
C8844 _316_/Q _317_/a_448_7# 0.00148f
C8845 _199_/a_250_257# _193_/Y 4.6e-19
C8846 _199_/a_584_7# _194_/X 0.00183f
C8847 _324_/a_448_7# _324_/Q 1.03e-20
C8848 _325_/a_651_373# VGND 0.00401f
C8849 _325_/a_639_7# VPWR 9.63e-20
C8850 _347_/Q _260_/A 9.15e-21
C8851 _215_/A _284_/A 0.155f
C8852 _251_/a_79_n19# _227_/A 5.61e-20
C8853 _157_/A _297_/B 0.0165f
C8854 _277_/Y _284_/A 0.00808f
C8855 _197_/X _190_/A 0.00854f
C8856 _319_/Q clkbuf_2_1_0_clk/A 0.0187f
C8857 _219_/a_250_257# _278_/a_68_257# 6.6e-21
C8858 _344_/a_652_n19# _345_/Q 2.43e-20
C8859 _344_/a_193_7# _345_/D 0.0012f
C8860 _320_/D _319_/a_27_7# 3.44e-19
C8861 _254_/Y _255_/X 2.46e-20
C8862 _339_/Q VPWR 2.75f
C8863 _257_/a_448_7# _254_/Y 0.00538f
C8864 _193_/Y _225_/B 4.74e-21
C8865 _189_/a_27_7# _209_/X 7.36e-21
C8866 _317_/a_1462_7# VGND 1.95e-19
C8867 _196_/A _182_/X 0.00467f
C8868 _202_/a_256_7# VPWR -6.36e-19
C8869 _202_/a_93_n19# VGND -0.00588f
C8870 _306_/a_76_159# _337_/Q 1.31e-21
C8871 trimb[0] input2/a_27_7# 0.00403f
C8872 _172_/A _345_/D 4.79e-19
C8873 _259_/a_199_7# _312_/Q 4.45e-20
C8874 _258_/a_505_n19# _313_/a_651_373# 9.43e-20
C8875 _219_/a_93_n19# _279_/A 0.00563f
C8876 _341_/a_543_7# _177_/a_27_7# 1.83e-19
C8877 _168_/a_109_7# _299_/X 0.00424f
C8878 cal VGND 0.842f
C8879 _160_/X _286_/Y 0.0157f
C8880 _205_/a_297_7# _204_/Y 0.00318f
C8881 _308_/S _296_/Y 0.0122f
C8882 result[2] _325_/Q 4.86e-20
C8883 _269_/A _315_/a_27_7# 0.0132f
C8884 _304_/X _284_/A 3.69e-21
C8885 _323_/a_1108_7# _191_/B 1.77e-19
C8886 _323_/a_1283_n19# _323_/Q 0.0676f
C8887 _303_/A VPWR 0.319f
C8888 _197_/a_27_7# VGND 0.0915f
C8889 _197_/X _337_/a_543_7# 9.33e-19
C8890 _327_/a_448_7# _331_/Q 1.32e-20
C8891 _292_/A _287_/a_121_257# 6.1e-20
C8892 _258_/a_505_n19# _157_/a_27_7# 0.00124f
C8893 _343_/a_1462_7# cal 2.24e-19
C8894 _342_/a_761_249# _343_/CLK 2.86e-19
C8895 _280_/a_150_257# VGND -3.06e-19
C8896 _290_/A _310_/Q 0.0103f
C8897 _283_/Y _339_/a_1283_n19# 1.37e-19
C8898 _301_/X _314_/Q 2.3e-20
C8899 _260_/A _297_/B 1.8e-20
C8900 _172_/A _254_/A 0.00896f
C8901 _255_/B _209_/a_109_257# 7.03e-21
C8902 _150_/a_193_257# VGND -1.48e-19
C8903 _281_/Y _324_/a_543_7# 0.00299f
C8904 _211_/a_27_257# _334_/Q 2.27e-20
C8905 _319_/Q _235_/a_113_257# 4.48e-19
C8906 _279_/Y _162_/X 0.0115f
C8907 _181_/X _343_/Q 2.83e-21
C8908 _286_/B _298_/C 0.651f
C8909 _322_/a_805_7# _321_/D 4.12e-20
C8910 _165_/a_493_257# _164_/Y 1.67e-19
C8911 _185_/A input3/a_27_7# 3.03e-19
C8912 _323_/a_639_7# _149_/A 9.53e-20
C8913 _322_/a_1108_7# _282_/a_39_257# 1.69e-20
C8914 _248_/A _330_/a_1108_7# 8.68e-20
C8915 _324_/a_448_7# _228_/A 0.0182f
C8916 clkbuf_2_3_0_clk/A _161_/Y 2.81e-20
C8917 _321_/a_543_7# _242_/A 5.46e-21
C8918 _281_/Y _217_/A 0.00472f
C8919 _265_/B _310_/a_27_7# 5.23e-20
C8920 _331_/CLK _330_/a_1108_7# 8.41e-19
C8921 _298_/X valid 0.00471f
C8922 _308_/X _225_/X 0.00106f
C8923 _196_/A _347_/a_448_7# 1.54e-19
C8924 _239_/a_113_257# _297_/B 0.00322f
C8925 _173_/a_76_159# _147_/Y 0.0276f
C8926 _307_/X _308_/X 2.14e-20
C8927 _219_/a_346_7# VGND 4.13e-20
C8928 _267_/B _311_/Q 5.75e-20
C8929 _346_/a_27_7# _297_/A 3.99e-20
C8930 _300_/Y _284_/A 1.72e-19
C8931 _153_/a_109_53# _335_/Q 0.0145f
C8932 _271_/A _324_/Q 0.322f
C8933 _342_/Q _315_/a_193_7# 4.73e-19
C8934 _342_/Q _298_/A 0.0169f
C8935 _206_/A _203_/a_303_7# 0.00123f
C8936 _166_/Y _346_/D 0.00799f
C8937 _161_/Y _172_/Y 1.32e-20
C8938 _172_/A _309_/D 2.67e-20
C8939 _333_/a_543_7# _332_/Q 9.52e-20
C8940 _333_/a_193_7# _190_/A 0.0135f
C8941 _342_/a_193_7# _149_/A 2.01e-21
C8942 _254_/Y _336_/a_193_7# 0.551f
C8943 _341_/a_27_7# _341_/a_543_7# -0.00936f
C8944 _341_/a_193_7# _341_/a_761_249# -0.0144f
C8945 _330_/Q _221_/a_93_n19# 1.93e-20
C8946 result[4] VPWR 0.278f
C8947 _255_/B _314_/a_27_7# 7.83e-20
C8948 repeater42/a_27_7# _286_/Y 8.68e-19
C8949 _319_/Q _278_/a_68_257# 9.41e-21
C8950 output32/a_27_7# output35/a_27_7# 4.25e-20
C8951 _250_/a_493_257# VGND -2.35e-19
C8952 _197_/X _339_/a_543_7# 7.82e-20
C8953 _321_/a_1108_7# _234_/B 0.00159f
C8954 _345_/a_27_7# _167_/X 3.81e-19
C8955 _273_/A _252_/a_109_257# 8.7e-20
C8956 _306_/a_505_n19# input1/X 2.15e-19
C8957 _321_/a_27_7# _321_/a_639_7# -0.0015f
C8958 _251_/X _227_/A 2.08e-19
C8959 _338_/a_27_7# _338_/a_543_7# -0.0117f
C8960 _338_/a_193_7# _338_/a_761_249# -0.0157f
C8961 result[4] _318_/a_543_7# 4.3e-19
C8962 _167_/a_27_257# clkbuf_2_1_0_clk/A 0.00364f
C8963 _268_/a_39_257# _316_/a_1108_7# 5.82e-19
C8964 _299_/X _306_/S 1.15e-19
C8965 _227_/A _296_/a_213_83# 8.91e-20
C8966 _304_/S _317_/D 2.54e-19
C8967 _285_/A _162_/a_27_7# 0.00735f
C8968 _342_/a_1270_373# repeater43/X 1.41e-19
C8969 _297_/B _221_/a_250_257# 7.5e-20
C8970 _209_/a_27_257# _335_/Q 2.02e-20
C8971 _346_/SET_B _312_/a_639_7# 8.67e-19
C8972 _340_/a_1283_n19# _194_/A 8.85e-21
C8973 _329_/a_27_7# _304_/X 7.11e-20
C8974 _284_/A VGND 1.58f
C8975 _336_/D VPWR 0.132f
C8976 _332_/a_193_7# _332_/a_651_373# -0.00334f
C8977 _319_/Q _218_/a_93_n19# 7.71e-20
C8978 _184_/a_535_334# cal 4.44e-20
C8979 _184_/a_218_334# input1/X 0.00226f
C8980 _306_/X _313_/a_448_7# 5.61e-19
C8981 _345_/a_1032_373# _290_/A 0.012f
C8982 _232_/X _331_/a_1108_7# 7.76e-19
C8983 _225_/X _254_/B 0.0378f
C8984 _236_/B _331_/Q 0.235f
C8985 _165_/X _347_/Q 0.00179f
C8986 _340_/a_805_7# _196_/A 5.2e-19
C8987 _269_/A _242_/B 0.00844f
C8988 _267_/A _311_/a_448_7# 0.0323f
C8989 _269_/A _315_/a_1217_7# 3.33e-19
C8990 result[2] _315_/a_1283_n19# 0.00329f
C8991 _182_/a_510_7# _333_/Q 4.89e-21
C8992 _305_/a_439_7# _192_/B 1.79e-21
C8993 _313_/Q _157_/a_27_7# 7.95e-21
C8994 _204_/Y _298_/A 3.78e-20
C8995 _337_/Q _198_/a_93_n19# 0.00461f
C8996 _309_/a_761_249# _284_/A 0.0431f
C8997 _271_/A _228_/A 0.0064f
C8998 _227_/A _205_/a_79_n19# 0.0571f
C8999 _219_/a_250_257# _328_/D 7.42e-19
C9000 _277_/Y _167_/a_109_7# 0.0021f
C9001 _294_/A _299_/X 1.3e-20
C9002 _284_/a_39_257# clkc 9.55e-21
C9003 _326_/D _331_/Q 1.61e-20
C9004 _343_/a_27_7# _269_/A 0.0165f
C9005 _323_/D _226_/X 3.6e-19
C9006 _317_/a_27_7# _317_/D 0.0549f
C9007 _317_/a_761_249# _244_/B 5.5e-36
C9008 _323_/a_1270_373# clk 2.18e-20
C9009 _279_/Y _340_/a_27_7# 0.0143f
C9010 _163_/a_215_7# _162_/X 0.0404f
C9011 _275_/Y _261_/A 0.234f
C9012 _315_/Q _341_/a_27_7# 3.11e-20
C9013 _310_/a_1283_n19# _310_/D 0.0211f
C9014 _310_/a_27_7# _310_/Q 2.43e-19
C9015 _326_/a_651_373# _181_/X 4.46e-19
C9016 _320_/Q _216_/X 0.108f
C9017 _346_/SET_B _299_/a_78_159# 0.00347f
C9018 _275_/A _297_/A 1.18e-20
C9019 _342_/Q _215_/A 0.0166f
C9020 _229_/a_76_159# _343_/Q 8.7e-19
C9021 _327_/a_193_7# _216_/X 0.0137f
C9022 _336_/a_27_7# _336_/a_448_7# -0.00642f
C9023 _336_/a_193_7# _336_/a_1108_7# -0.00677f
C9024 _259_/a_199_7# _340_/CLK 1.99e-20
C9025 _290_/A _311_/a_27_7# 3.34e-20
C9026 _325_/Q _224_/a_250_257# 0.00149f
C9027 _283_/Y input1/a_75_172# 2.83e-19
C9028 _320_/Q _329_/Q 1f
C9029 _196_/A _340_/CLK 1.1f
C9030 _343_/a_27_7# _343_/D 0.0519f
C9031 _343_/a_761_249# _185_/A 0.0111f
C9032 _231_/a_79_n19# _144_/A 0.00387f
C9033 _196_/A _347_/D 5.82e-20
C9034 _172_/A clkbuf_0_clk/X 0.224f
C9035 _327_/a_193_7# _329_/Q 5.36e-21
C9036 output10/a_27_7# rstn 4.16e-19
C9037 _277_/Y input4/a_27_7# 2.23e-20
C9038 _153_/A _335_/Q 0.0176f
C9039 _346_/a_1032_373# _299_/a_215_7# 3.51e-20
C9040 _327_/a_27_7# _327_/a_543_7# -0.00385f
C9041 _327_/a_193_7# _327_/a_761_249# -0.0118f
C9042 _271_/A _216_/A 1.52e-19
C9043 _165_/X _297_/B 0.0121f
C9044 _255_/a_30_13# VPWR 0.0726f
C9045 clkbuf_1_0_0_clk/a_75_172# VPWR 0.0817f
C9046 _318_/Q _317_/a_193_7# 2.17e-19
C9047 _324_/a_1283_n19# _255_/B 1.58e-19
C9048 _323_/a_651_373# cal 0.00132f
C9049 _342_/a_1108_7# _149_/a_27_7# 8.68e-19
C9050 clkbuf_0_clk/X _232_/X 0.139f
C9051 _306_/a_218_334# _284_/A 0.00111f
C9052 _328_/a_27_7# _216_/X 0.00149f
C9053 _315_/Q _316_/a_193_7# 2.75e-19
C9054 _329_/a_543_7# _330_/Q 0.00408f
C9055 _268_/a_39_257# _248_/A 0.00828f
C9056 _227_/A rstn 1.21e-19
C9057 repeater43/X _330_/a_639_7# 8.67e-19
C9058 _331_/D _331_/a_543_7# 0.0105f
C9059 _262_/a_113_257# clkc 1.13e-20
C9060 _331_/a_27_7# _330_/a_1283_n19# 2.37e-20
C9061 trim[2] VGND 0.151f
C9062 _326_/a_27_7# _326_/a_543_7# -0.00936f
C9063 _326_/a_193_7# _326_/a_761_249# -0.0157f
C9064 _162_/X _313_/a_27_7# 1.01e-20
C9065 _328_/a_193_7# _320_/Q 0.0108f
C9066 _328_/a_27_7# _329_/Q 0.197f
C9067 _339_/Q _198_/a_93_n19# 0.00261f
C9068 output37/a_27_7# comp 0.0121f
C9069 _273_/A _299_/a_215_7# 5.09e-20
C9070 _215_/A _264_/a_113_257# 1.02e-20
C9071 _341_/Q _175_/Y 0.0174f
C9072 _318_/Q _331_/a_1283_n19# 2.21e-21
C9073 _341_/Q _243_/a_113_257# 8.26e-20
C9074 _330_/D _281_/A 0.0657f
C9075 ctlp[6] clkbuf_1_0_0_clk/a_75_172# 5.77e-19
C9076 repeater43/X _333_/a_1108_7# -0.0219f
C9077 _329_/a_761_249# VPWR 0.0152f
C9078 _329_/a_27_7# VGND -0.084f
C9079 _268_/a_39_257# _331_/CLK 1.66e-19
C9080 _144_/a_27_7# _304_/X 4.31e-20
C9081 _308_/a_505_n19# _306_/S 0.00216f
C9082 _296_/a_493_257# VPWR 2.47e-20
C9083 _172_/A input1/X 9.45e-20
C9084 _181_/X _346_/SET_B 7.84e-19
C9085 input2/a_27_7# VPWR 0.0822f
C9086 _251_/X _297_/B 0.148f
C9087 _341_/a_1108_7# _229_/a_489_373# 1.24e-20
C9088 _329_/a_1283_n19# _297_/B 1.1e-19
C9089 _191_/B _147_/Y 4.87e-20
C9090 _252_/a_27_7# _212_/X 8.86e-21
C9091 _338_/Q _312_/D 1.71e-19
C9092 _322_/a_651_373# result[6] 0.00368f
C9093 _332_/a_543_7# _340_/CLK 3.33e-22
C9094 _333_/a_639_7# _206_/A 7.55e-19
C9095 _332_/a_761_249# _332_/D 7.16e-19
C9096 _301_/a_245_257# _347_/Q 2.87e-19
C9097 _290_/A _309_/a_1283_n19# 0.0051f
C9098 _329_/a_193_7# repeater42/a_27_7# 2.76e-19
C9099 _306_/X _337_/Q 7.66e-20
C9100 _328_/a_27_7# _328_/a_193_7# -0.329f
C9101 _153_/a_403_257# _153_/A 0.00196f
C9102 _153_/a_215_257# _154_/A 0.0105f
C9103 _347_/a_1283_n19# _347_/D 4.1e-20
C9104 clk _254_/B 0.00978f
C9105 _308_/X _150_/a_109_257# 4.27e-20
C9106 _209_/X _154_/A 0.0249f
C9107 _164_/A _345_/D 1.87e-19
C9108 _267_/A _311_/D 0.289f
C9109 _258_/a_505_n19# _267_/A 6.49e-21
C9110 _334_/Q _333_/a_1108_7# 2.43e-19
C9111 _319_/Q _328_/D 0.0294f
C9112 _269_/A ctln[0] 0.00182f
C9113 _242_/A _318_/D 0.0385f
C9114 output24/a_27_7# VPWR 0.0998f
C9115 _291_/a_39_257# _310_/D 1.4e-21
C9116 _316_/a_27_7# _248_/A 0.00964f
C9117 _254_/A _297_/A 1.36e-19
C9118 clkbuf_2_3_0_clk/A _263_/B 0.114f
C9119 _172_/A _286_/Y 0.101f
C9120 _270_/a_39_257# VPWR 0.0469f
C9121 _230_/a_27_7# _318_/a_193_7# 5.68e-19
C9122 _315_/a_193_7# _315_/a_448_7# -0.00482f
C9123 result[0] _341_/a_639_7# 2.99e-19
C9124 _333_/a_543_7# _192_/B 9.28e-20
C9125 _333_/a_1108_7# _191_/B 0.00484f
C9126 _331_/Q _331_/a_193_7# 0.31f
C9127 _326_/Q _224_/a_250_257# 0.00174f
C9128 _316_/a_27_7# _331_/CLK 0.0244f
C9129 _344_/Q _171_/a_78_159# 0.0355f
C9130 _340_/a_193_7# _190_/A 1.06e-19
C9131 _310_/a_1217_7# _310_/Q 1.58e-19
C9132 _242_/A _217_/A 0.0114f
C9133 _209_/a_373_7# _153_/A 0.0016f
C9134 _209_/a_109_257# _154_/A 0.047f
C9135 _232_/X _286_/Y 0.0027f
C9136 output11/a_27_7# _332_/Q 0.00213f
C9137 _338_/a_448_7# _340_/CLK 0.0165f
C9138 input1/X _203_/a_80_n19# 0.0322f
C9139 _275_/Y _165_/X 0.00797f
C9140 _167_/a_109_7# VGND 4.04e-19
C9141 _169_/B clkbuf_2_1_0_clk/A 0.145f
C9142 _242_/A _346_/D 2.67e-20
C9143 _346_/SET_B _347_/a_1108_7# 0.012f
C9144 input1/a_75_172# _312_/a_27_7# 7.27e-21
C9145 _219_/a_584_7# _232_/X 6.98e-19
C9146 _334_/a_27_7# _334_/a_193_7# -0.293f
C9147 _328_/a_27_7# _274_/a_39_257# 3.41e-21
C9148 _181_/X _222_/a_346_7# 5.01e-19
C9149 _321_/a_27_7# _321_/Q 0.141f
C9150 _162_/X _144_/A 4.32e-19
C9151 _286_/B _345_/Q 0.00531f
C9152 _322_/D _318_/D 6.36e-20
C9153 repeater43/X _304_/a_79_n19# 5.3e-19
C9154 _338_/a_761_249# _337_/a_27_7# 1e-20
C9155 _338_/a_193_7# _337_/a_193_7# 4.55e-20
C9156 _318_/a_193_7# _232_/A 2.89e-19
C9157 output22/a_27_7# _248_/A 0.00122f
C9158 _181_/X _206_/A 5.64e-20
C9159 _286_/B _207_/C 2.41e-19
C9160 _161_/Y _260_/A 1.11e-19
C9161 _314_/a_27_7# _314_/a_193_7# -0.00228f
C9162 _286_/B _313_/a_1283_n19# 0.00319f
C9163 _311_/a_27_7# _310_/a_27_7# 2.01e-21
C9164 _283_/Y _195_/a_27_257# 2.45e-19
C9165 output10/a_27_7# clkbuf_2_0_0_clk/a_75_172# 0.0127f
C9166 _306_/X _339_/Q 5.78e-22
C9167 _342_/Q VGND 0.824f
C9168 _257_/a_544_257# VGND -0.00117f
C9169 _337_/Q _147_/Y 7.02e-19
C9170 _323_/D input1/X 3.75e-19
C9171 _292_/Y VGND 0.305f
C9172 _144_/a_27_7# VGND 0.058f
C9173 _279_/Y _332_/D 2.69e-19
C9174 _321_/a_27_7# _318_/a_193_7# 3.7e-21
C9175 _321_/a_193_7# _318_/a_27_7# 2.91e-20
C9176 input4/a_27_7# VGND 0.0487f
C9177 _283_/A _246_/B 0.0721f
C9178 _277_/Y _199_/a_250_257# 9.84e-20
C9179 _224_/a_93_n19# _224_/a_346_7# -3.48e-20
C9180 _332_/a_1270_373# _333_/Q 1.27e-19
C9181 repeater43/X _176_/a_27_7# 8.22e-20
C9182 output8/a_27_7# output34/a_27_7# 3.1e-20
C9183 _340_/a_27_7# _337_/a_1283_n19# 0.00383f
C9184 _340_/a_1283_n19# _337_/a_27_7# 0.00383f
C9185 _210_/a_307_257# VPWR -2.5e-19
C9186 _314_/Q _297_/Y 4.04e-19
C9187 _305_/a_439_7# _260_/A 7.03e-19
C9188 _303_/A _227_/a_113_7# 2.88e-21
C9189 _338_/a_651_373# _346_/SET_B 0.00215f
C9190 _338_/a_1270_373# _338_/D 2.49e-19
C9191 _338_/a_1283_n19# _338_/Q 0.00128f
C9192 _169_/Y _215_/A 8.1e-20
C9193 _329_/Q _319_/a_761_249# 3.77e-21
C9194 _238_/B _319_/a_27_7# 0.0193f
C9195 _215_/A _225_/B 0.127f
C9196 _244_/B _286_/Y 0.018f
C9197 _310_/a_1283_n19# VPWR 0.0326f
C9198 _310_/a_761_249# VGND 0.00517f
C9199 _319_/D VPWR 0.297f
C9200 _277_/Y _169_/Y 6.63e-20
C9201 ctln[7] _207_/a_27_7# 2.39e-20
C9202 repeater43/X _332_/a_27_7# 0.00182f
C9203 _344_/a_1032_373# _344_/D 7.17e-20
C9204 _344_/a_562_373# _344_/Q 1.68e-20
C9205 _341_/a_805_7# _248_/A 7.43e-19
C9206 _309_/a_193_7# clkc 6.82e-21
C9207 _319_/Q _322_/a_27_7# 1.57e-20
C9208 _292_/A _338_/Q 0.0152f
C9209 _297_/A _302_/a_227_257# 0.00116f
C9210 _343_/Q _206_/A 8.1e-20
C9211 _258_/a_76_159# _340_/Q 1.28e-20
C9212 _194_/X _311_/D 0.00283f
C9213 _258_/a_505_n19# _194_/X 1.03e-21
C9214 _334_/a_27_7# _332_/Q 6.5e-21
C9215 _275_/A _292_/A 0.0211f
C9216 _145_/A _162_/X 4.79e-20
C9217 _343_/CLK valid 0.309f
C9218 _304_/a_591_329# _304_/S 0.00309f
C9219 _264_/a_113_257# VGND 0.00162f
C9220 output31/a_27_7# VPWR 0.142f
C9221 _196_/A _225_/X 0.00381f
C9222 _181_/X _147_/A 0.00608f
C9223 _286_/B _150_/C 0.0126f
C9224 _307_/X _196_/A 3.63e-20
C9225 _323_/D _286_/Y 7.33e-19
C9226 _334_/D _343_/Q 1.8e-20
C9227 _332_/a_1283_n19# _206_/A 0.0625f
C9228 _339_/a_761_249# _338_/a_27_7# 0.00344f
C9229 _339_/a_193_7# _338_/a_193_7# 7.1e-19
C9230 _256_/a_80_n19# _191_/B 0.017f
C9231 _309_/a_761_249# _310_/a_761_249# 0.00117f
C9232 _229_/a_226_257# _248_/A 2.6e-19
C9233 _313_/Q _267_/A 2.7e-19
C9234 ctln[6] _211_/a_109_257# 0.00123f
C9235 output12/a_27_7# _197_/X 0.00737f
C9236 clkbuf_2_3_0_clk/A _194_/A 6.46e-20
C9237 _321_/a_193_7# _246_/B 7.75e-21
C9238 _275_/A _238_/B 7.51e-19
C9239 _339_/Q _147_/Y 2.32e-20
C9240 _323_/Q output41/a_27_7# 5.42e-21
C9241 _324_/Q _231_/a_79_n19# 8.1e-19
C9242 _342_/a_543_7# _228_/A 1.1e-19
C9243 _327_/a_651_373# _346_/SET_B 0.00203f
C9244 _324_/a_1283_n19# _326_/Q 0.00421f
C9245 _316_/Q _248_/B 3.15e-20
C9246 _346_/a_193_7# _346_/a_1182_221# -1.52e-19
C9247 repeater43/X _341_/a_543_7# -4.24e-19
C9248 _339_/Q _312_/a_1108_7# 0.00408f
C9249 _204_/Y VGND 0.0757f
C9250 clkbuf_2_2_0_clk/a_75_172# _338_/a_1108_7# 2.39e-20
C9251 _316_/a_1217_7# _248_/A 1.48e-19
C9252 _177_/A _226_/X 4.77e-20
C9253 _158_/Y _162_/A 5.22e-20
C9254 _185_/A _184_/a_218_7# 5.9e-19
C9255 _203_/a_209_257# _284_/A 3.33e-19
C9256 _258_/S clkbuf_2_3_0_clk/A 0.00813f
C9257 input4/X _338_/a_1108_7# 4e-19
C9258 _340_/a_543_7# _339_/a_193_7# 2.3e-19
C9259 _340_/a_761_249# _339_/a_761_249# 7.15e-19
C9260 _340_/a_193_7# _339_/a_543_7# 2.44e-20
C9261 _242_/a_109_257# _242_/B 1.07e-20
C9262 _242_/A _314_/Q 1.8e-20
C9263 _190_/A _295_/a_79_n19# 0.0011f
C9264 _164_/A _162_/a_27_7# 6.65e-20
C9265 _242_/A _318_/a_448_7# 7.26e-19
C9266 _315_/a_193_7# _315_/D 0.00926f
C9267 _309_/Q _265_/B 5.51e-21
C9268 _320_/a_1283_n19# _328_/Q 0.00814f
C9269 _315_/D _298_/A 0.212f
C9270 _240_/B _232_/X 1.15e-19
C9271 _344_/a_1182_221# _290_/A 0.00223f
C9272 _344_/Q _172_/B 0.104f
C9273 _149_/a_27_7# _177_/a_27_7# 3.1e-20
C9274 _298_/a_181_7# VGND 2.71e-19
C9275 _329_/a_651_373# _330_/D 0.00405f
C9276 _343_/Q _147_/A 5.88e-19
C9277 _329_/a_27_7# _214_/a_27_257# 1.1e-20
C9278 _338_/D _340_/CLK 0.537f
C9279 _336_/a_761_249# VPWR 0.00169f
C9280 _346_/a_27_7# _273_/A 1.95e-19
C9281 _324_/a_27_7# _227_/A 0.334f
C9282 _336_/a_27_7# VGND -0.115f
C9283 _328_/a_448_7# _346_/SET_B 0.00157f
C9284 input1/X _312_/a_448_7# 1.19e-19
C9285 _320_/Q _282_/a_39_257# 0.0281f
C9286 _321_/a_1217_7# _321_/Q 8.83e-19
C9287 _207_/X _332_/Q 0.0309f
C9288 _149_/A _343_/Q 0.262f
C9289 _260_/a_27_257# VPWR 0.106f
C9290 clkbuf_0_clk/X _297_/A 0.00875f
C9291 _292_/A _345_/D 3.39e-20
C9292 _168_/a_109_7# _172_/B 2.55e-21
C9293 _279_/Y input4/X 3.55e-19
C9294 repeater43/X _316_/a_1283_n19# -0.00619f
C9295 _324_/a_1108_7# _224_/a_250_257# 1.76e-20
C9296 _300_/a_27_257# _299_/X 0.00333f
C9297 _147_/A _347_/a_1108_7# 0.0105f
C9298 _321_/a_651_373# VGND 0.00142f
C9299 _321_/a_639_7# VPWR 6.63e-19
C9300 _281_/Y _254_/B 0.01f
C9301 rstn _335_/a_543_7# 0.0343f
C9302 _160_/A _345_/D 5.82e-20
C9303 _179_/a_27_7# _306_/S 0.00335f
C9304 _300_/Y _225_/B 6.03e-21
C9305 _163_/a_78_159# _173_/a_226_7# 1.54e-20
C9306 _232_/X _328_/Q 0.19f
C9307 _320_/Q _327_/Q 9.54e-21
C9308 _329_/a_193_7# _232_/X 8.22e-21
C9309 _153_/a_487_257# VGND -8.69e-19
C9310 _224_/a_346_7# _217_/A 8.36e-19
C9311 _224_/a_250_257# _324_/D 4.28e-21
C9312 _291_/a_39_257# VPWR 0.0463f
C9313 _194_/A _192_/B 4.24e-19
C9314 _327_/a_193_7# _327_/Q 0.0229f
C9315 _327_/a_27_7# _212_/X 0.00654f
C9316 _319_/a_27_7# _331_/CLK 8.25e-20
C9317 _326_/a_543_7# repeater43/X 0.0446f
C9318 _162_/X _174_/a_27_257# 6.96e-20
C9319 _260_/B _313_/a_448_7# 6.27e-19
C9320 _275_/Y _310_/a_448_7# 0.00564f
C9321 _206_/A _204_/a_27_7# 1.39e-19
C9322 _305_/a_505_n19# _340_/D 0.00106f
C9323 _231_/a_79_n19# _228_/A 1.1e-19
C9324 _281_/A _330_/a_1283_n19# 6.09e-20
C9325 _326_/a_27_7# _212_/X 0.00624f
C9326 _326_/a_193_7# _327_/Q 1.11e-19
C9327 _277_/A clkbuf_2_1_0_clk/a_75_172# 5.66e-19
C9328 _281_/Y _331_/D 1e-20
C9329 _199_/a_250_257# VGND -0.00251f
C9330 _199_/a_346_7# VPWR -5.69e-19
C9331 _307_/a_505_n19# _295_/a_79_n19# 0.0023f
C9332 repeater43/X _332_/a_1217_7# 1.88e-19
C9333 _165_/X _161_/Y 0.0148f
C9334 _315_/Q repeater43/X 0.0215f
C9335 _281_/Y _330_/a_193_7# 2.86e-19
C9336 _343_/D _323_/a_448_7# 0.00239f
C9337 _337_/a_193_7# _201_/a_27_7# 4.5e-21
C9338 _313_/Q _194_/X 0.00503f
C9339 output20/a_27_7# clkbuf_2_1_0_clk/A 0.035f
C9340 _313_/D _193_/Y 2.53e-19
C9341 _343_/CLK _204_/a_277_7# 2.36e-20
C9342 output12/a_27_7# _333_/a_193_7# 5.29e-20
C9343 _328_/a_27_7# _327_/Q 3.88e-21
C9344 _302_/a_77_159# _347_/a_543_7# 0.00301f
C9345 _183_/a_1241_257# _181_/X 0.00335f
C9346 _183_/a_471_7# _286_/B 0.00391f
C9347 _346_/a_562_373# _346_/SET_B 6.82e-19
C9348 clk _196_/A 0.00618f
C9349 clkbuf_2_1_0_clk/A _278_/a_150_257# 0.00128f
C9350 _254_/A _238_/B 0.0029f
C9351 _169_/Y VGND 0.258f
C9352 _346_/a_1032_373# _275_/A 3.34e-21
C9353 _325_/a_1108_7# _181_/X 0.00291f
C9354 result[5] _321_/a_193_7# 0.0018f
C9355 _225_/B VGND 0.327f
C9356 _184_/a_76_159# _175_/Y 1.14e-20
C9357 _340_/CLK _313_/a_193_7# 2.89e-19
C9358 _197_/X _193_/Y 0.42f
C9359 _260_/B _191_/B 4.16e-19
C9360 _275_/A _331_/CLK 7.16e-20
C9361 repeater43/X _334_/a_761_249# -0.00425f
C9362 input4/X _334_/a_1283_n19# 8.76e-22
C9363 _316_/Q _315_/a_27_7# 1.8e-20
C9364 output23/a_27_7# _315_/a_1283_n19# 0.0131f
C9365 trim[0] _297_/Y 2.3e-19
C9366 _337_/a_1108_7# _340_/CLK 0.0402f
C9367 _285_/A clkc 0.927f
C9368 _215_/A _315_/D 0.0437f
C9369 _145_/A _298_/C 0.0863f
C9370 _308_/X _185_/A 9.08e-19
C9371 _329_/D _330_/a_193_7# 0.00143f
C9372 _324_/Q _162_/X 0.165f
C9373 _342_/a_27_7# _185_/A 4.8e-19
C9374 _324_/a_651_373# _215_/A 1.67e-19
C9375 _273_/A _338_/Q 0.0143f
C9376 output10/a_27_7# VPWR 0.0981f
C9377 _309_/Q _310_/Q 2.53e-19
C9378 _343_/CLK _340_/CLK 0.016f
C9379 _309_/a_1108_7# _265_/B 0.00603f
C9380 clkbuf_2_1_0_clk/A _279_/A 0.305f
C9381 _271_/A input3/a_27_7# 6.36e-20
C9382 _160_/a_27_7# _162_/A 0.013f
C9383 _337_/a_27_7# _337_/a_193_7# -0.0518f
C9384 _344_/a_476_7# _297_/Y 0.0338f
C9385 _297_/A _286_/Y 3.87e-20
C9386 _286_/B _202_/a_93_n19# 0.00229f
C9387 _306_/S _172_/B 1.04e-20
C9388 _147_/Y _336_/D 0.0807f
C9389 _297_/A _297_/a_27_257# 0.00984f
C9390 _334_/a_448_7# _206_/A 5.12e-21
C9391 _334_/a_1283_n19# _207_/C 0.0492f
C9392 _163_/a_78_159# _158_/Y 0.0116f
C9393 _236_/B _321_/D 0.00416f
C9394 _320_/D _328_/Q 0.00229f
C9395 _344_/a_1296_7# _290_/A 3.35e-19
C9396 _315_/a_448_7# VGND 0.00139f
C9397 _315_/a_1270_373# VPWR -1.77e-19
C9398 _311_/Q _297_/Y 0.0572f
C9399 _255_/X _172_/A 2.67e-20
C9400 en VGND 0.156f
C9401 _286_/B cal 0.209f
C9402 _227_/A VPWR 0.919f
C9403 _336_/a_1217_7# VGND -3.75e-19
C9404 _180_/a_29_13# _178_/a_27_7# 0.00714f
C9405 _339_/a_27_7# _332_/Q 5.58e-20
C9406 _317_/a_193_7# _316_/a_448_7# 2.02e-20
C9407 _271_/A _224_/a_93_n19# 7.63e-21
C9408 _329_/a_27_7# _330_/a_27_7# 0.00512f
C9409 _324_/a_27_7# _324_/a_639_7# -0.0015f
C9410 _326_/a_27_7# _325_/a_193_7# 1.96e-19
C9411 _326_/a_193_7# _325_/a_27_7# 2.98e-20
C9412 _334_/a_448_7# _334_/D 0.0145f
C9413 _334_/a_761_249# _334_/Q 3.07e-20
C9414 input1/X _312_/D 1.16e-19
C9415 _318_/a_27_7# _242_/B 1.52e-19
C9416 _315_/D _314_/a_639_7# 0.00462f
C9417 _196_/A _301_/X 1.8e-20
C9418 _286_/B _197_/a_27_7# 3.5e-19
C9419 _329_/a_27_7# _318_/Q 1.8e-20
C9420 ctln[1] _334_/a_27_7# 6.35e-21
C9421 _314_/a_543_7# VGND -0.00412f
C9422 _314_/a_1108_7# VPWR 0.0131f
C9423 clkbuf_2_1_0_clk/A _311_/a_193_7# 2.49e-21
C9424 _187_/a_27_7# _304_/X 1.15e-20
C9425 _269_/A _244_/B 0.00807f
C9426 _346_/SET_B _319_/a_1270_373# 1.39e-19
C9427 _324_/a_27_7# _297_/B 0.0229f
C9428 _346_/SET_B _313_/a_761_249# -0.00247f
C9429 ctln[7] _283_/A 0.0016f
C9430 _315_/D _304_/X 1.15e-19
C9431 _346_/SET_B _337_/a_448_7# 2.63e-21
C9432 _338_/a_543_7# _337_/Q 2.8e-20
C9433 _275_/A _319_/a_1108_7# 8.9e-37
C9434 clk _332_/a_543_7# 0.0055f
C9435 _224_/a_584_7# VGND 3.37e-19
C9436 _299_/X _160_/X 0.23f
C9437 _324_/a_1283_n19# _324_/D 0.0583f
C9438 _314_/a_761_249# _314_/Q 8.24e-21
C9439 _314_/a_448_7# _314_/D 0.00377f
C9440 _271_/A _153_/A 6.2e-21
C9441 _311_/D _310_/a_1108_7# 6.99e-20
C9442 _196_/A _150_/a_109_257# 1.27e-20
C9443 _181_/X _150_/a_27_7# 1.05e-19
C9444 _170_/a_226_257# VGND -4.16e-19
C9445 repeater43/X _333_/Q 0.122f
C9446 _322_/a_1270_373# _269_/A 4.66e-20
C9447 input1/X _177_/A 3.47e-20
C9448 clkbuf_0_clk/X _325_/D 1.25e-20
C9449 _346_/a_1602_7# _345_/Q 5.39e-21
C9450 _334_/a_193_7# _323_/Q 0.00115f
C9451 _334_/a_27_7# _192_/B 1.53e-19
C9452 _279_/Y _302_/a_77_159# 0.00125f
C9453 _325_/a_1270_373# _325_/D 3.05e-19
C9454 _263_/B _261_/A 0.144f
C9455 _319_/Q _322_/Q 0.0132f
C9456 _339_/a_1108_7# _340_/CLK 3.94e-19
C9457 _341_/D _304_/S 9.48e-20
C9458 _163_/a_215_7# _345_/Q 0.00124f
C9459 _163_/a_493_257# _345_/D 7.35e-21
C9460 _153_/a_215_257# _153_/B 0.0151f
C9461 _323_/D _269_/A 0.0962f
C9462 _343_/D _244_/B 4.53e-21
C9463 _185_/A _317_/D 2.35e-20
C9464 _323_/a_1283_n19# _175_/Y 9.12e-19
C9465 _294_/A _172_/B 1.3e-20
C9466 ctlp[0] result[6] 0.00767f
C9467 _340_/a_1108_7# _337_/Q 0.025f
C9468 _320_/a_448_7# _242_/A 1.16e-19
C9469 _345_/a_193_7# _297_/B 0.00647f
C9470 repeater43/a_27_7# input4/X 0.0176f
C9471 _275_/Y _310_/D 0.0187f
C9472 _339_/a_193_7# _337_/a_27_7# 0.00143f
C9473 _339_/a_27_7# _337_/a_193_7# 0.00143f
C9474 _326_/a_1108_7# _331_/a_1283_n19# 1e-20
C9475 input1/X _333_/D 5.35e-21
C9476 _162_/X _228_/A 0.0071f
C9477 _273_/A _345_/D 4.17e-20
C9478 _326_/D _222_/a_584_7# 5.27e-20
C9479 _254_/A _248_/A 9.06e-21
C9480 _296_/Y _295_/a_79_n19# 0.00161f
C9481 _277_/A _320_/a_761_249# 0.00108f
C9482 _307_/X _341_/D 5.25e-19
C9483 _255_/X _203_/a_80_n19# 5.6e-20
C9484 _246_/B _242_/B 4.16e-20
C9485 _343_/D _323_/D 0.431f
C9486 _184_/a_76_159# _341_/Q 2.04e-20
C9487 _323_/a_27_7# input3/a_27_7# 5.21e-19
C9488 _300_/Y _315_/D 1.85e-20
C9489 _346_/SET_B _147_/A 0.936f
C9490 _334_/Q _333_/Q 0.0211f
C9491 clkbuf_2_3_0_clk/A _337_/a_27_7# 2.43e-37
C9492 _168_/a_397_257# _162_/X 0.0451f
C9493 _257_/a_222_53# _254_/B 0.0205f
C9494 _342_/a_639_7# _269_/A 7.77e-19
C9495 _254_/A _331_/CLK 2.04e-20
C9496 repeater43/a_27_7# _207_/C 1.05e-19
C9497 _347_/Q VPWR 0.674f
C9498 _308_/S _298_/A 4.74e-20
C9499 _328_/a_639_7# _217_/X 7.76e-19
C9500 _308_/a_218_7# _227_/A 2.46e-19
C9501 _303_/A _347_/a_193_7# 6.44e-20
C9502 _301_/X _347_/a_1283_n19# 3.19e-19
C9503 ctln[1] _207_/X 7.04e-21
C9504 _209_/a_109_257# _153_/B 1.29e-20
C9505 _177_/A _286_/Y 0.00574f
C9506 _322_/a_1108_7# _321_/a_27_7# 8.52e-21
C9507 _173_/a_226_7# _172_/Y 0.0146f
C9508 output41/a_27_7# sample 8.39e-22
C9509 valid output30/a_27_7# 0.00763f
C9510 _319_/a_27_7# _217_/X 1.56e-19
C9511 _318_/a_193_7# _245_/a_113_257# 3.15e-20
C9512 _290_/Y ctlp[2] 2.81e-19
C9513 _339_/a_448_7# _346_/SET_B -2.34e-19
C9514 _339_/Q _338_/a_543_7# 5.26e-19
C9515 _188_/S _175_/Y 4.09e-21
C9516 _248_/A _226_/X 0.199f
C9517 _316_/Q _242_/B 6.5e-20
C9518 _273_/A _254_/A 0.0802f
C9519 _188_/a_76_159# _147_/A 1.17e-20
C9520 _218_/a_346_7# _304_/X 7.16e-19
C9521 _309_/a_1108_7# _310_/Q 1.45e-19
C9522 output37/a_27_7# trimb[1] 0.0085f
C9523 _279_/A _278_/a_68_257# 0.00672f
C9524 ctln[4] output9/a_27_7# 4.39e-20
C9525 output10/a_27_7# ctln[3] 1.62e-19
C9526 _191_/B _333_/Q 0.0085f
C9527 _304_/S _143_/a_27_7# 0.0373f
C9528 _172_/A _336_/a_193_7# 7.06e-22
C9529 _216_/A _162_/X 0.00915f
C9530 _313_/a_193_7# _313_/a_543_7# -0.0231f
C9531 _188_/a_76_159# _149_/A 4.25e-19
C9532 _326_/D _304_/S 4.53e-21
C9533 _316_/D _150_/C 3.33e-20
C9534 _341_/a_1283_n19# input1/X 3.78e-22
C9535 _267_/A _347_/a_27_7# 1.02e-20
C9536 output37/a_27_7# VGND 0.072f
C9537 _321_/Q VPWR 0.432f
C9538 _286_/B _284_/A 0.179f
C9539 _227_/A _335_/a_1108_7# 7.78e-20
C9540 _163_/a_78_159# _160_/a_27_7# 5.29e-20
C9541 _340_/a_639_7# _339_/D 3.06e-19
C9542 _340_/a_1108_7# _339_/Q 0.0014f
C9543 _184_/a_505_n19# _227_/A 5.22e-19
C9544 _238_/B clkbuf_0_clk/X 0.29f
C9545 clk _208_/a_493_257# 4.81e-19
C9546 _334_/D _206_/A 3.17e-19
C9547 _198_/a_93_n19# _336_/a_761_249# 2.54e-21
C9548 _198_/a_250_257# _336_/a_193_7# 3.7e-20
C9549 _260_/A _194_/A 0.00663f
C9550 _187_/a_27_7# VGND 0.074f
C9551 _255_/a_30_13# _333_/a_1108_7# 9.24e-21
C9552 _327_/a_1283_n19# clkbuf_0_clk/X 0.0448f
C9553 _315_/D VGND 3.44f
C9554 ctln[5] _339_/D 0.00202f
C9555 _339_/a_27_7# _339_/a_193_7# -0.00704f
C9556 _324_/Q _298_/C 0.0104f
C9557 _321_/Q _318_/a_543_7# 2.6e-21
C9558 _325_/D _286_/Y 0.0159f
C9559 _275_/A _217_/X 0.00183f
C9560 _324_/a_639_7# VPWR 4.63e-19
C9561 _324_/a_651_373# VGND 0.00308f
C9562 _271_/A _217_/A 8.1e-20
C9563 _236_/B _317_/a_27_7# 1.54e-19
C9564 _317_/a_193_7# _316_/D 4.77e-20
C9565 _317_/a_761_249# _331_/CLK 8.12e-19
C9566 repeater43/X _226_/a_297_7# 1.09e-19
C9567 _306_/a_439_7# clkbuf_2_1_0_clk/A 3.89e-19
C9568 _258_/S _260_/A 1.02e-19
C9569 _143_/a_109_7# _149_/A 3.29e-20
C9570 output7/a_27_7# _334_/D 2.76e-19
C9571 _297_/B VPWR 4.89f
C9572 _318_/a_193_7# VPWR -0.284f
C9573 _343_/a_1270_373# VPWR 9.95e-20
C9574 _343_/a_448_7# VGND 0.00299f
C9575 _218_/a_93_n19# _218_/a_250_257# -6.97e-22
C9576 _346_/SET_B _337_/D 2.24e-19
C9577 _242_/A _317_/D 6.8e-19
C9578 _172_/A clkbuf_2_3_0_clk/a_75_172# 2.52e-19
C9579 _297_/A _328_/Q 2.04e-20
C9580 input4/X _339_/a_1283_n19# 1.08e-20
C9581 _281_/Y _196_/A 0.0256f
C9582 _304_/S _343_/CLK 0.00842f
C9583 _279_/Y cal 0.00774f
C9584 _254_/B _335_/Q 6.31e-20
C9585 _345_/a_193_7# _275_/Y 0.00863f
C9586 _344_/a_1032_373# _265_/B 1.41e-20
C9587 _331_/CLK _331_/a_1108_7# 8.22e-20
C9588 _318_/a_193_7# _318_/a_543_7# -0.0129f
C9589 _147_/A _206_/A 4.53e-21
C9590 _313_/a_761_249# _147_/A 0.0228f
C9591 _341_/a_1283_n19# _286_/Y 0.106f
C9592 _279_/Y _197_/a_27_7# 8.09e-19
C9593 _345_/a_562_373# VGND -5.84e-35
C9594 _345_/a_1140_373# VPWR 1.85e-19
C9595 _258_/S _261_/A 0.263f
C9596 _158_/Y _172_/Y 0.00225f
C9597 _254_/B _298_/a_109_7# 1.77e-19
C9598 _149_/A _206_/A 5.23e-20
C9599 _307_/a_76_159# _191_/B 0.0533f
C9600 _319_/Q _181_/X 3.27e-20
C9601 _316_/Q _245_/a_199_7# 2.57e-19
C9602 _283_/A _330_/a_448_7# 1.82e-19
C9603 _343_/CLK _225_/X 1.05e-20
C9604 _281_/Y _256_/a_303_7# 0.00165f
C9605 clk _334_/a_1108_7# 0.00466f
C9606 _308_/S _215_/A 7.77e-20
C9607 _326_/D _331_/a_543_7# 2.7e-20
C9608 _339_/a_651_373# _337_/a_1108_7# 1.23e-20
C9609 _339_/a_1108_7# _337_/a_651_373# 1.23e-20
C9610 _331_/D _242_/A 5.4e-20
C9611 _311_/a_27_7# _311_/a_193_7# -0.00496f
C9612 _162_/A _267_/A 0.00916f
C9613 _307_/a_218_7# _147_/A 0.0018f
C9614 _283_/A _333_/a_761_249# 0.0213f
C9615 _307_/X _307_/a_535_334# 1.23e-19
C9616 _188_/a_218_334# _145_/A 0.00111f
C9617 repeater43/X _212_/X 0.258f
C9618 _149_/A _334_/D 1.44e-20
C9619 _229_/a_226_7# output30/a_27_7# 5.51e-20
C9620 _310_/D _171_/a_292_257# 9.1e-20
C9621 _188_/S _341_/Q 0.0295f
C9622 _181_/a_27_7# _314_/a_27_7# 4.09e-21
C9623 _218_/a_346_7# VGND -3.17e-19
C9624 _198_/a_346_7# _336_/Q 9.35e-19
C9625 _309_/a_1283_n19# _309_/Q 0.0078f
C9626 _239_/a_113_257# _320_/Q 0.00164f
C9627 _307_/X _178_/a_193_257# 6.93e-19
C9628 _308_/a_218_334# VPWR -2.02e-19
C9629 _308_/a_76_159# VGND 0.0216f
C9630 _293_/a_121_257# clkbuf_2_1_0_clk/A 1.35e-19
C9631 _181_/X _250_/X 0.456f
C9632 _298_/C _228_/A 1.99e-19
C9633 _238_/B _286_/Y 3.09e-20
C9634 _343_/a_761_249# _323_/a_27_7# 3.84e-21
C9635 _343_/a_27_7# _323_/a_761_249# 3.5e-21
C9636 ctln[6] _332_/a_193_7# 0.00814f
C9637 _294_/Y _288_/A 0.0254f
C9638 _294_/A trim[1] 0.0185f
C9639 _339_/D _346_/SET_B 0.0206f
C9640 _283_/Y _153_/A 9.79e-21
C9641 _311_/a_1108_7# VPWR 0.0238f
C9642 _311_/a_543_7# VGND 0.0252f
C9643 _330_/D _217_/A 1.13e-21
C9644 clkbuf_0_clk/X _248_/A 0.0123f
C9645 cal _334_/a_1283_n19# 0.00118f
C9646 _313_/Q _336_/a_543_7# 0.00678f
C9647 _306_/X _336_/a_761_249# 8.63e-20
C9648 _294_/Y _162_/X 0.00756f
C9649 _346_/a_1032_373# clkbuf_0_clk/X 4.32e-20
C9650 _342_/a_1283_n19# _298_/A 7.11e-21
C9651 _149_/A _147_/A 4.15e-19
C9652 _319_/Q ctlp[1] 9.04e-21
C9653 _252_/a_27_7# _248_/B 5.25e-19
C9654 _199_/a_93_n19# _254_/B 2.16e-21
C9655 clkbuf_0_clk/X _331_/CLK 0.975f
C9656 _271_/Y ctln[0] 2.07e-20
C9657 _216_/X _221_/a_93_n19# 0.0263f
C9658 _337_/a_448_7# _337_/D 0.00197f
C9659 _337_/a_761_249# _337_/Q 0.0199f
C9660 _172_/A _314_/a_1283_n19# 3.35e-21
C9661 _161_/Y _310_/D 1.58e-19
C9662 clkbuf_0_clk/X _190_/A 1.8e-20
C9663 _335_/a_193_7# VGND 3.25e-19
C9664 _335_/a_543_7# VPWR 2.35e-19
C9665 _197_/X _336_/a_448_7# 5.81e-19
C9666 _267_/a_109_257# _309_/D 0.00427f
C9667 _275_/Y VPWR 0.888f
C9668 _298_/B _154_/a_27_7# 5.91e-19
C9669 trim[4] _162_/a_27_7# 2e-19
C9670 _273_/A clkbuf_0_clk/X 0.048f
C9671 _306_/S _305_/X 0.00147f
C9672 _225_/B _203_/a_209_257# 0.00369f
C9673 _336_/Q _203_/a_209_7# 2.75e-19
C9674 _340_/Q _194_/A 0.247f
C9675 _216_/A _298_/C 7.07e-20
C9676 _144_/A _150_/C 0.273f
C9677 _336_/Q _254_/B 0.736f
C9678 _327_/a_193_7# _221_/a_250_257# 5.77e-22
C9679 _333_/a_27_7# _153_/a_109_53# 2.72e-19
C9680 _338_/a_27_7# _306_/S 0.0148f
C9681 _338_/a_193_7# _340_/Q 0.00795f
C9682 _338_/a_761_249# _194_/X 0.00843f
C9683 _325_/a_193_7# repeater43/X 0.00189f
C9684 _279_/Y _284_/A 0.0108f
C9685 input1/X _248_/A 0.006f
C9686 _260_/B _336_/D 0.00477f
C9687 _258_/S _340_/Q 1.27e-19
C9688 _318_/a_805_7# VGND -7.08e-19
C9689 _318_/a_1462_7# VPWR 2.28e-19
C9690 repeater43/X _149_/a_27_7# 0.00546f
C9691 _277_/A output18/a_27_7# 0.0293f
C9692 _275_/Y _309_/a_27_7# 0.017f
C9693 _164_/A clkc 2.29e-20
C9694 _328_/D _279_/A 1.05e-19
C9695 _164_/Y _297_/Y 0.00736f
C9696 _344_/a_193_7# _299_/X 0.00232f
C9697 _344_/a_27_7# _347_/Q 4.21e-20
C9698 result[7] _282_/a_39_257# 0.00259f
C9699 _309_/a_639_7# VPWR 0.00289f
C9700 _309_/a_651_373# VGND 9.33e-19
C9701 repeater43/X _317_/a_448_7# 0.0266f
C9702 input1/X _190_/A 0.00742f
C9703 _340_/a_543_7# _340_/Q 0.00495f
C9704 _340_/a_193_7# _193_/Y 0.0117f
C9705 _340_/a_761_249# _306_/S 0.00412f
C9706 _340_/a_1283_n19# _194_/X 0.0505f
C9707 _269_/A _177_/A 0.00205f
C9708 _336_/a_761_249# _147_/Y 0.0222f
C9709 _255_/X _192_/a_68_257# 0.0137f
C9710 _219_/a_250_257# _346_/SET_B 0.0805f
C9711 _172_/A _299_/X 0.00706f
C9712 _339_/D _206_/A 2.24e-21
C9713 _260_/A _201_/a_27_7# 2.72e-21
C9714 _234_/B _331_/Q 0.0064f
C9715 clk _343_/CLK 0.0618f
C9716 _333_/a_27_7# _209_/a_27_257# 0.00366f
C9717 _321_/a_1283_n19# _331_/Q 0.00348f
C9718 _321_/a_1108_7# _322_/Q 0.0156f
C9719 _220_/a_346_7# _328_/D 0.00129f
C9720 _339_/a_761_249# _337_/Q 4.55e-21
C9721 _339_/Q _337_/a_761_249# 0.00752f
C9722 repeater43/X _331_/a_639_7# 0.00117f
C9723 _231_/a_676_257# _298_/A 1.62e-19
C9724 _145_/A _150_/C 0.009f
C9725 _323_/Q _192_/B 0.0226f
C9726 _331_/a_193_7# _331_/a_543_7# -0.0102f
C9727 _327_/a_448_7# _281_/Y 0.00623f
C9728 _248_/A _286_/Y 0.162f
C9729 _301_/a_240_7# _162_/X 3.67e-19
C9730 _309_/a_27_7# _309_/a_639_7# -0.0015f
C9731 _331_/a_448_7# _212_/X 0.00168f
C9732 _331_/a_1108_7# _217_/X 7.13e-21
C9733 _313_/D _215_/A 0.0205f
C9734 _342_/Q _286_/B 0.685f
C9735 _255_/B _181_/X 0.812f
C9736 _337_/a_543_7# _202_/a_250_257# 2.71e-21
C9737 _320_/a_193_7# VPWR 0.0287f
C9738 _257_/a_544_257# _286_/B 3.82e-20
C9739 _257_/a_222_53# _196_/A 0.0117f
C9740 _346_/a_1032_373# _286_/Y 5.03e-20
C9741 _185_/A _298_/X 0.0102f
C9742 _323_/a_543_7# VPWR 0.0228f
C9743 _323_/a_193_7# VGND 0.0045f
C9744 _146_/a_112_13# _150_/C 5.79e-20
C9745 _188_/a_439_7# _146_/C 2.59e-19
C9746 _240_/B _238_/B 1.05e-19
C9747 _331_/CLK _286_/Y 0.114f
C9748 _308_/S VGND 0.41f
C9749 _320_/a_543_7# _297_/B 0.0347f
C9750 _227_/A _227_/a_113_7# 6.36e-20
C9751 _190_/A _286_/Y 2.04e-20
C9752 _345_/a_193_7# _161_/Y 5.93e-20
C9753 _200_/a_256_7# _193_/Y 7.08e-19
C9754 _344_/a_27_7# _297_/B 0.0103f
C9755 _277_/Y _197_/X 2.35e-20
C9756 _291_/a_39_257# _312_/a_1108_7# 6.87e-19
C9757 _256_/a_209_257# _255_/X 0.00653f
C9758 _258_/a_76_159# VPWR 0.00667f
C9759 _273_/A _286_/Y 0.587f
C9760 _344_/Q _173_/a_76_159# 2.84e-21
C9761 _183_/a_1241_257# _149_/A 4.76e-20
C9762 _186_/a_382_257# VGND -5.47e-19
C9763 _217_/a_27_7# _331_/a_1283_n19# 0.0117f
C9764 _335_/a_193_7# _335_/a_651_373# -0.00701f
C9765 _275_/Y ctln[3] 0.00943f
C9766 _329_/a_543_7# _216_/X 0.00254f
C9767 _345_/a_1032_373# _344_/a_1032_373# 0.00204f
C9768 _250_/a_215_7# _190_/A 0.00764f
C9769 _328_/a_448_7# _319_/Q 0.0139f
C9770 _222_/a_93_n19# _286_/Y 3.54e-20
C9771 _335_/a_1462_7# VGND -8.37e-19
C9772 _343_/a_193_7# _342_/a_1283_n19# 7.21e-21
C9773 _343_/a_761_249# _342_/a_543_7# 8.8e-19
C9774 _343_/a_27_7# _342_/a_1108_7# 2.47e-19
C9775 _338_/a_27_7# _283_/A 5.16e-20
C9776 input1/X _178_/a_27_7# 4.39e-20
C9777 _329_/a_1283_n19# _320_/Q 2.77e-20
C9778 _238_/B _328_/Q 0.0611f
C9779 _330_/Q _212_/a_27_7# 0.0151f
C9780 _183_/a_471_7# _144_/A 4.19e-19
C9781 _339_/a_448_7# _339_/D 0.0144f
C9782 _339_/a_761_249# _339_/Q 4.13e-19
C9783 _268_/a_121_257# _248_/B 2.24e-20
C9784 _328_/a_1108_7# _329_/D 1.37e-20
C9785 _320_/a_651_373# _279_/A 4.31e-20
C9786 _327_/a_1283_n19# _328_/Q 3.72e-20
C9787 _329_/a_1283_n19# _327_/a_193_7# 1.12e-20
C9788 _329_/a_1108_7# _327_/a_27_7# 2.18e-20
C9789 _327_/a_27_7# _327_/D 0.0518f
C9790 _346_/SET_B _195_/a_109_7# 7.72e-19
C9791 _171_/a_292_257# VPWR -3.26e-19
C9792 _333_/a_27_7# _153_/A 6.33e-19
C9793 _325_/a_1462_7# repeater43/X -6.42e-19
C9794 _210_/a_109_257# _333_/D 9.57e-19
C9795 output19/a_27_7# VGND 0.104f
C9796 _326_/a_27_7# _327_/D 1.8e-21
C9797 _297_/Y _347_/a_1283_n19# 1.65e-19
C9798 _317_/a_27_7# _317_/a_639_7# -0.0015f
C9799 clkbuf_0_clk/X _217_/X 0.287f
C9800 _196_/A _335_/Q 5.79e-20
C9801 _325_/a_639_7# _212_/X 4.94e-20
C9802 _340_/a_761_249# _283_/A 4.89e-21
C9803 _277_/Y _312_/a_193_7# 1.83e-19
C9804 trim[0] _311_/a_761_249# 4.89e-20
C9805 _285_/A _311_/a_1283_n19# 1.63e-19
C9806 cal _339_/a_1283_n19# 2.23e-19
C9807 _325_/Q _181_/X 2.37e-20
C9808 _307_/a_505_n19# _286_/Y 4.08e-20
C9809 _329_/a_1283_n19# _328_/a_27_7# 7.17e-21
C9810 _328_/a_543_7# _328_/Q 2.16e-19
C9811 _269_/A _316_/a_1108_7# 0.0178f
C9812 _147_/A _150_/a_27_7# 3.37e-19
C9813 _319_/Q _346_/SET_B 0.472f
C9814 _339_/a_27_7# _260_/A 7.69e-21
C9815 _182_/a_215_7# _298_/A 0.0041f
C9816 output13/a_27_7# _335_/a_193_7# 7.22e-20
C9817 _317_/Q _316_/a_27_7# 2.95e-20
C9818 output24/a_27_7# _316_/a_1283_n19# 0.00235f
C9819 _286_/B _336_/a_27_7# 0.0154f
C9820 _345_/a_652_n19# _172_/B 0.0073f
C9821 _175_/Y output41/a_27_7# 9.6e-20
C9822 _294_/Y _165_/a_215_7# 2.36e-19
C9823 _322_/a_651_373# _321_/Q 6.97e-19
C9824 _341_/a_1108_7# _342_/Q 2.94e-19
C9825 _178_/a_27_7# _286_/Y 6.05e-20
C9826 ctln[7] ctln[0] 1.39e-19
C9827 _308_/a_505_n19# _172_/A 2.03e-19
C9828 _161_/Y VPWR 0.17f
C9829 _271_/Y _323_/a_448_7# 1.96e-19
C9830 _339_/D _337_/D 6.2e-21
C9831 ctln[6] _190_/A 0.00498f
C9832 _340_/Q _201_/a_27_7# 2.68e-19
C9833 _311_/a_448_7# _311_/D 0.00197f
C9834 _311_/a_761_249# _311_/Q 2.13e-19
C9835 _326_/a_27_7# _283_/A 0.00822f
C9836 _157_/A _157_/a_27_7# 0.0172f
C9837 _318_/a_27_7# _244_/B 9.72e-20
C9838 _218_/a_584_7# _232_/X 4.95e-19
C9839 _346_/a_562_373# _319_/Q 4.51e-20
C9840 _322_/a_1108_7# VPWR -7.86e-19
C9841 _232_/X _246_/B 0.227f
C9842 _322_/a_543_7# VGND 0.00622f
C9843 _313_/a_27_7# _284_/A 0.00992f
C9844 _315_/a_27_7# _177_/a_27_7# 2.01e-21
C9845 _344_/a_27_7# _275_/Y 0.0205f
C9846 _320_/a_1462_7# VPWR 1.79e-19
C9847 _320_/a_805_7# VGND 0.00227f
C9848 input4/a_27_7# _338_/a_1108_7# 1.9e-19
C9849 input4/X _195_/a_27_257# 0.00128f
C9850 rstn _338_/a_193_7# 7.07e-19
C9851 _298_/a_109_7# _298_/X 3.66e-19
C9852 _323_/a_1462_7# VGND 1.14e-19
C9853 ctlp[4] clkbuf_2_1_0_clk/A 0.126f
C9854 output39/a_27_7# ctlp[3] 2.08e-19
C9855 trimb[3] output17/a_27_7# 1.33e-19
C9856 _290_/A _346_/SET_B 0.0989f
C9857 _331_/Q clkbuf_2_1_0_clk/A 2.78e-20
C9858 _305_/a_439_7# VPWR -1.27e-19
C9859 _305_/a_535_334# VGND -2.65e-19
C9860 _344_/a_381_7# VGND 0.00301f
C9861 _344_/a_956_373# VPWR -6.78e-19
C9862 _292_/A clkc 2.06e-19
C9863 trim[3] _297_/Y 0.00386f
C9864 _315_/Q output24/a_27_7# 9.36e-21
C9865 _343_/Q _298_/a_27_7# 0.00109f
C9866 _318_/Q _315_/D 1.36e-19
C9867 _160_/X _172_/B 0.0181f
C9868 _309_/a_27_7# _161_/Y 1.8e-20
C9869 _308_/X _271_/A 4.26e-19
C9870 _340_/D _340_/CLK 0.41f
C9871 _332_/a_761_249# _204_/Y 1.08e-20
C9872 output25/a_27_7# VPWR 0.124f
C9873 clkbuf_2_3_0_clk/A _267_/A 0.176f
C9874 _343_/a_651_373# _323_/D 0.00153f
C9875 _306_/S _173_/a_76_159# 0.00707f
C9876 _324_/Q _150_/C 0.101f
C9877 _250_/a_78_159# _147_/A 0.0232f
C9878 _160_/A clkc 2.53e-19
C9879 _313_/D VGND 0.244f
C9880 clkbuf_0_clk/a_110_7# clkbuf_0_clk/X 0.0177f
C9881 _263_/B _310_/D 2.73e-19
C9882 _320_/Q _321_/a_27_7# 3.02e-20
C9883 _258_/S _310_/a_448_7# 2.94e-20
C9884 _255_/a_30_13# _333_/Q 1.13e-20
C9885 _271_/Y _335_/D 0.0017f
C9886 _337_/a_27_7# _340_/Q 2.67e-19
C9887 _337_/a_193_7# _194_/X 0.0122f
C9888 _248_/A _328_/Q 0.00471f
C9889 output11/a_27_7# rstn 0.0382f
C9890 _342_/a_1283_n19# VGND 0.0362f
C9891 _342_/a_448_7# VPWR 0.00151f
C9892 _335_/a_761_249# _335_/D 0.00154f
C9893 _296_/Y input1/X 3.19e-20
C9894 repeater43/X _207_/a_27_7# 0.00362f
C9895 _184_/a_76_159# _188_/S 2.89e-19
C9896 _199_/a_256_7# _312_/D 5.77e-20
C9897 _297_/A _314_/a_1283_n19# 0.00403f
C9898 _324_/Q _317_/a_193_7# 4.01e-21
C9899 _197_/X VGND 1.6f
C9900 _217_/X _286_/Y 0.426f
C9901 _329_/a_193_7# _331_/CLK 0.0308f
C9902 _347_/Q _147_/Y 0.0079f
C9903 _331_/CLK _328_/Q 0.0101f
C9904 _268_/a_39_257# _315_/a_193_7# 3.26e-20
C9905 _260_/A _157_/a_27_7# 0.0399f
C9906 _246_/B _244_/B 0.646f
C9907 _265_/B _312_/Q 1.3e-20
C9908 ctlp[1] _321_/a_1108_7# 8.13e-20
C9909 _169_/Y _286_/B 0.00109f
C9910 _196_/A _336_/Q 0.00837f
C9911 _286_/B _225_/B 0.0094f
C9912 trim[1] _284_/a_39_257# 1.88e-21
C9913 _273_/A _328_/Q 0.0399f
C9914 _338_/Q _193_/Y 0.0176f
C9915 _320_/a_193_7# _320_/a_543_7# -0.0102f
C9916 _162_/X _300_/a_383_7# 1.78e-33
C9917 clkbuf_0_clk/a_110_7# input1/X 3.41e-21
C9918 _181_/X _326_/Q 0.0744f
C9919 _235_/a_113_257# _331_/Q 0.0143f
C9920 _341_/a_27_7# _315_/a_27_7# 1.62e-20
C9921 _316_/Q _244_/B 0.107f
C9922 _269_/A _248_/A 0.707f
C9923 clkbuf_2_1_0_clk/A _299_/a_292_257# 7.27e-20
C9924 _336_/a_1283_n19# _194_/A 8.77e-20
C9925 _209_/X _332_/a_1108_7# 2.87e-20
C9926 _271_/A _254_/B 0.0136f
C9927 _327_/Q _221_/a_93_n19# 0.0124f
C9928 _222_/a_93_n19# _328_/Q 5.4e-20
C9929 _271_/A _317_/D 1.94e-19
C9930 _296_/Y _286_/Y 0.0067f
C9931 _294_/Y output35/a_27_7# 0.0128f
C9932 _250_/X _206_/A 9.54e-25
C9933 _216_/A _313_/a_1283_n19# 0.0418f
C9934 _167_/a_27_257# _346_/SET_B 0.00606f
C9935 _269_/A _331_/CLK 0.194f
C9936 ctln[7] _335_/a_448_7# 0.0162f
C9937 _258_/S _336_/a_1283_n19# 0.00562f
C9938 _309_/a_193_7# _172_/B 4.27e-20
C9939 _286_/B _336_/a_1217_7# 6.79e-20
C9940 _345_/a_1056_7# _172_/B 6.53e-19
C9941 _339_/a_193_7# _194_/X 7.22e-19
C9942 _339_/a_27_7# _340_/Q 0.00898f
C9943 _319_/a_1108_7# _328_/Q 1.68e-20
C9944 _298_/C _209_/a_27_257# 2.22e-19
C9945 _228_/A _150_/C 0.631f
C9946 _312_/a_193_7# VGND 0.041f
C9947 _312_/a_543_7# VPWR 0.038f
C9948 _146_/a_29_271# _286_/Y 1.68e-20
C9949 rstn _334_/a_27_7# 1.78e-20
C9950 _297_/A _299_/X 6.82e-20
C9951 _181_/X _314_/a_193_7# 1.65e-19
C9952 _196_/A _314_/a_761_249# 7.72e-19
C9953 _335_/Q _204_/a_27_257# 0.0519f
C9954 _319_/Q _147_/A 5.27e-20
C9955 _297_/B _147_/Y 0.00404f
C9956 _271_/Y _323_/D 7.71e-20
C9957 _208_/a_493_257# _335_/Q 9.28e-20
C9958 _208_/a_292_257# _204_/Y 9.45e-19
C9959 input1/a_75_172# cal 0.0439f
C9960 _326_/a_1217_7# _283_/A 2.76e-19
C9961 _340_/a_27_7# _336_/a_651_373# 2.18e-21
C9962 _340_/a_1283_n19# _336_/a_543_7# 1.97e-19
C9963 _316_/a_193_7# _315_/a_27_7# 1.57e-20
C9964 _304_/a_79_n19# _227_/A 0.0191f
C9965 _316_/a_27_7# _315_/a_193_7# 3.18e-21
C9966 _231_/a_676_257# VGND -3.88e-19
C9967 _231_/a_409_7# VPWR -6.53e-19
C9968 clkbuf_2_3_0_clk/A _194_/X 0.012f
C9969 clkbuf_0_clk/a_110_7# _286_/Y 0.00142f
C9970 _313_/a_1217_7# _284_/A 1.32e-19
C9971 _315_/a_651_373# _177_/A 1.27e-20
C9972 _279_/Y _336_/a_27_7# 9.66e-21
C9973 _330_/Q _330_/a_1270_373# 9.01e-21
C9974 _326_/a_448_7# _242_/A 0.0137f
C9975 _344_/a_586_7# _275_/Y 2.97e-19
C9976 _346_/a_1224_7# _167_/X 3.74e-20
C9977 _180_/a_111_257# _283_/A 2.91e-19
C9978 repeater43/X _306_/S 2.32e-20
C9979 _186_/a_79_n19# _308_/X 0.00379f
C9980 _186_/a_297_7# _172_/A 0.0417f
C9981 _289_/a_39_257# VGND 0.00154f
C9982 output17/a_27_7# VPWR 0.132f
C9983 _165_/X _158_/Y 2.31e-20
C9984 clkbuf_2_0_0_clk/a_75_172# _338_/a_193_7# 1.59e-20
C9985 _188_/a_76_159# _255_/B 0.00562f
C9986 _342_/a_27_7# _186_/a_79_n19# 2.71e-21
C9987 _260_/B _260_/a_27_257# 0.0101f
C9988 _330_/a_651_373# VPWR -0.0088f
C9989 _330_/a_1108_7# VGND 0.0413f
C9990 _258_/a_76_159# _198_/a_93_n19# 2.82e-21
C9991 _329_/a_639_7# _346_/SET_B -7.75e-19
C9992 _281_/Y _331_/a_193_7# 2.97e-21
C9993 _162_/X _217_/A 3.18e-19
C9994 _251_/a_297_257# _191_/B 4.61e-20
C9995 _344_/a_193_7# _171_/a_78_159# 0.00765f
C9996 _183_/a_471_7# _324_/Q 0.00739f
C9997 _343_/a_27_7# _177_/a_27_7# 1.23e-21
C9998 _328_/a_1108_7# _242_/A 5.05e-20
C9999 _250_/X _147_/A 0.0152f
C10000 _162_/X _346_/D 0.0203f
C10001 _216_/A _150_/C 4.26e-20
C10002 _342_/Q _316_/D 2.32e-20
C10003 clkbuf_0_clk/a_110_7# _250_/a_215_7# 2.12e-19
C10004 _145_/A _284_/A 0.00268f
C10005 _346_/SET_B _310_/a_27_7# 0.015f
C10006 _333_/a_193_7# VGND 0.026f
C10007 _333_/a_543_7# VPWR 0.0184f
C10008 _345_/a_1182_221# _162_/X 7.88e-20
C10009 _167_/X clkbuf_2_3_0_clk/A 0.0171f
C10010 _341_/a_761_249# _341_/Q 3.89e-20
C10011 _252_/a_109_257# VGND -3.31e-19
C10012 _302_/a_77_159# _228_/A 4.89e-20
C10013 _144_/a_27_7# _316_/D 1.25e-19
C10014 _258_/S _310_/D 0.00419f
C10015 _255_/X _190_/A 0.0497f
C10016 output22/a_27_7# _315_/a_193_7# 0.00169f
C10017 _337_/a_1217_7# _340_/Q 4.27e-20
C10018 _218_/a_93_n19# _331_/Q 0.0485f
C10019 _257_/a_448_7# _190_/A 0.0143f
C10020 _342_/D VPWR 0.223f
C10021 _240_/B _217_/X 0.00149f
C10022 _312_/Q _310_/Q 0.00158f
C10023 rstn _207_/X 0.0212f
C10024 _334_/a_1108_7# _335_/Q 1.16e-20
C10025 _273_/A clkc 0.118f
C10026 _273_/Y _297_/Y 0.229f
C10027 _210_/a_27_7# _332_/Q 6.07e-20
C10028 _308_/S _203_/a_209_257# 7.83e-20
C10029 _314_/a_1283_n19# _347_/a_761_249# 0.00226f
C10030 _314_/a_1108_7# _347_/a_193_7# 0.0106f
C10031 _167_/X _172_/Y 2.3e-20
C10032 _254_/A _193_/Y 2.32e-20
C10033 _322_/a_27_7# _322_/a_193_7# -0.00111f
C10034 _325_/a_543_7# _284_/A 2.53e-19
C10035 _160_/X trimb[4] 2.28e-19
C10036 _344_/a_27_7# _161_/Y 9.47e-19
C10037 _343_/Q _154_/A 0.00282f
C10038 _298_/C _153_/A 3.23e-19
C10039 _185_/A _343_/CLK 0.274f
C10040 _189_/a_27_7# _206_/A 6.05e-19
C10041 _170_/a_226_7# _347_/a_1108_7# 8.54e-19
C10042 _312_/a_543_7# _311_/a_651_373# 5.67e-20
C10043 _312_/a_1108_7# _311_/a_1108_7# 5.35e-21
C10044 _320_/D _320_/a_27_7# 0.0461f
C10045 _306_/S _191_/B 0.151f
C10046 _323_/a_761_249# _323_/D 1.56e-20
C10047 repeater43/X _327_/D 5.15e-20
C10048 _255_/B _206_/A 1.93e-19
C10049 _294_/Y _345_/Q 1.48e-19
C10050 _332_/a_1283_n19# _154_/A 4.68e-21
C10051 _340_/CLK _153_/a_215_257# 4.67e-21
C10052 _329_/a_27_7# _331_/a_27_7# 0.0054f
C10053 _330_/D _331_/D 2.21e-19
C10054 _279_/Y _225_/B 1.1f
C10055 _330_/D _330_/a_193_7# 0.00253f
C10056 _304_/S _247_/a_113_257# 2.58e-21
C10057 _329_/a_193_7# _217_/X 0.00111f
C10058 _329_/a_761_249# _212_/X 2.14e-19
C10059 _217_/X _328_/Q 0.0283f
C10060 output19/a_27_7# ctlp[5] 0.0052f
C10061 _329_/a_543_7# _327_/Q 3.69e-20
C10062 _344_/a_27_7# _344_/a_956_373# -0.00135f
C10063 trim[4] clkc 0.0865f
C10064 _275_/Y _147_/Y 6.99e-19
C10065 _200_/a_93_n19# clkbuf_2_1_0_clk/A 0.00595f
C10066 _263_/B VPWR 2f
C10067 _286_/B _315_/D 0.116f
C10068 ctln[3] _312_/a_543_7# 2.21e-19
C10069 _275_/Y _312_/a_1108_7# 0.00204f
C10070 ctln[7] _335_/D 0.0208f
C10071 _182_/a_215_7# VGND 0.00259f
C10072 _309_/D _193_/Y 0.00299f
C10073 _236_/B _242_/A 0.374f
C10074 _324_/a_1108_7# _181_/X 0.0136f
C10075 _183_/a_471_7# _228_/A 0.176f
C10076 _219_/a_93_n19# _219_/a_256_7# -6.6e-20
C10077 _339_/a_651_373# _340_/D 1.08e-20
C10078 _339_/a_805_7# _306_/S 4.26e-19
C10079 _339_/a_639_7# _193_/Y 5.49e-19
C10080 _339_/a_1217_7# _340_/Q 3.05e-20
C10081 _339_/a_1462_7# _194_/X 4.04e-19
C10082 _157_/A _267_/A 0.005f
C10083 _265_/B _340_/CLK 0.00197f
C10084 _347_/Q _347_/a_193_7# 6.48e-20
C10085 _258_/a_218_7# _313_/D 8.85e-19
C10086 _258_/a_505_n19# _313_/Q 0.0481f
C10087 _258_/a_76_159# _306_/X 0.00323f
C10088 repeater43/X _283_/A 0.522f
C10089 _161_/Y _171_/a_215_7# 0.0871f
C10090 _181_/X _324_/D 0.00969f
C10091 _326_/a_651_373# _326_/Q 3.49e-19
C10092 _287_/a_121_257# VGND -3.99e-19
C10093 _174_/a_27_257# _284_/A 1.95e-20
C10094 _326_/D _242_/A 0.0279f
C10095 _286_/a_113_7# _297_/B 1.48e-19
C10096 _162_/X _314_/Q 6.44e-20
C10097 _296_/Y _296_/a_295_257# 6.95e-19
C10098 _279_/Y _314_/a_543_7# 0.0116f
C10099 _255_/B _147_/A 0.0063f
C10100 _260_/B _314_/a_1108_7# 3.9e-19
C10101 _342_/a_1108_7# _172_/A 1.65e-20
C10102 _336_/a_1283_n19# _201_/a_27_7# 6.06e-19
C10103 _258_/S _266_/a_113_257# 0.00399f
C10104 _342_/a_27_7# _342_/a_543_7# -0.00482f
C10105 _321_/D _234_/B 0.0023f
C10106 _344_/a_193_7# _172_/B 0.00717f
C10107 _183_/a_471_7# _216_/A 1.63e-20
C10108 _255_/B _149_/A 2.11e-19
C10109 clkbuf_2_3_0_clk/A _301_/a_51_257# 0.00595f
C10110 _343_/a_1108_7# _298_/X 1.6e-20
C10111 _321_/a_1270_373# _331_/CLK 3.05e-19
C10112 _345_/a_27_7# _162_/A 9.3e-21
C10113 clkbuf_2_3_0_clk/A clkbuf_1_1_0_clk/a_75_172# 0.00478f
C10114 _338_/D _199_/a_93_n19# 0.00373f
C10115 _325_/a_651_373# _216_/A 5.16e-20
C10116 _333_/a_1462_7# VGND -8.77e-19
C10117 repeater43/X _248_/B 1.43e-19
C10118 output15/a_27_7# VPWR 0.108f
C10119 _271_/A _223_/a_584_7# 9e-20
C10120 _180_/a_29_13# _298_/A 0.00648f
C10121 _211_/a_109_7# _197_/X 0.00109f
C10122 _283_/A _334_/Q 1.63e-19
C10123 _343_/a_1283_n19# _343_/Q 0.00136f
C10124 _337_/Q _306_/S 0.0187f
C10125 _299_/a_215_7# VGND 0.0488f
C10126 _346_/Q _301_/X 0.00826f
C10127 _197_/X _198_/a_256_7# 0.00283f
C10128 rstn _339_/a_27_7# 3.52e-20
C10129 _315_/D _347_/a_543_7# 0.00146f
C10130 _260_/A _267_/A 1.28f
C10131 _172_/A _172_/B 0.0145f
C10132 _174_/a_373_7# _344_/D 0.00211f
C10133 _154_/A _204_/a_27_7# 1.33e-20
C10134 clkbuf_2_3_0_clk/a_75_172# _331_/CLK 1.62e-19
C10135 _343_/CLK _335_/Q 0.205f
C10136 repeater43/X _321_/a_193_7# 0.0137f
C10137 _308_/a_76_159# _286_/B 0.00369f
C10138 _324_/Q _284_/A 0.0236f
C10139 _144_/a_27_7# _144_/A 0.0105f
C10140 _305_/a_218_334# _254_/B 3.77e-19
C10141 _336_/a_27_7# _313_/a_27_7# 7.65e-19
C10142 _268_/a_39_257# VGND 0.00577f
C10143 _297_/B _347_/a_193_7# 0.574f
C10144 _314_/a_27_7# _347_/D 0.00118f
C10145 _314_/D _347_/a_27_7# 6.2e-20
C10146 _283_/A _191_/B 0.0243f
C10147 _237_/a_113_257# _279_/A 5.15e-19
C10148 _258_/a_76_159# _147_/Y 4.41e-20
C10149 _267_/A _261_/A 0.0221f
C10150 _312_/Q _311_/a_27_7# 0.00424f
C10151 _191_/B _205_/a_382_257# 0.00113f
C10152 ctlp[0] _321_/Q 2.4e-19
C10153 _341_/D _315_/a_1108_7# 4.95e-20
C10154 _332_/D _153_/A 9.64e-20
C10155 _175_/Y _226_/a_382_257# 0.00119f
C10156 _194_/A VPWR 1.79f
C10157 _265_/a_109_257# _267_/A 0.0013f
C10158 _341_/a_193_7# VPWR -0.0776f
C10159 _271_/A _196_/A 1.78e-20
C10160 _341_/Q _332_/Q 4.54e-19
C10161 _342_/a_543_7# _317_/D 1.55e-20
C10162 _342_/a_1108_7# _244_/B 0.00108f
C10163 clkbuf_2_1_0_clk/A _340_/CLK 0.043f
C10164 _338_/a_193_7# VPWR -0.313f
C10165 _207_/C _153_/a_109_53# 1.92e-19
C10166 _294_/A _337_/Q 1.44e-19
C10167 _339_/a_805_7# _283_/A 0.00205f
C10168 _346_/SET_B _336_/a_639_7# 5.38e-19
C10169 _346_/a_27_7# _277_/Y 2.92e-20
C10170 _319_/D _212_/X 4.59e-20
C10171 _258_/S VPWR 2.57f
C10172 _340_/CLK _310_/Q 8.86e-19
C10173 _346_/SET_B _314_/a_193_7# -6.5e-19
C10174 _219_/a_93_n19# _329_/D 4.22e-19
C10175 _345_/a_1182_221# _165_/a_215_7# 2.94e-19
C10176 _342_/Q _145_/A 0.17f
C10177 _339_/Q _306_/S 2.05e-20
C10178 _147_/A _298_/a_27_7# 0.00613f
C10179 _330_/Q _216_/X 0.527f
C10180 _248_/A _242_/a_109_257# 3.7e-20
C10181 _308_/a_505_n19# _333_/D 8.78e-20
C10182 _315_/a_651_373# _248_/A 0.00516f
C10183 _188_/a_535_334# _298_/A 0.00107f
C10184 _317_/Q _317_/a_761_249# 0.0013f
C10185 _271_/A _298_/X 0.0158f
C10186 _340_/a_543_7# VPWR 0.0164f
C10187 _193_/Y _202_/a_250_257# 1.12e-19
C10188 _340_/a_193_7# VGND -0.00182f
C10189 _329_/Q _330_/Q 5.46e-19
C10190 _300_/Y _347_/a_1270_373# 1.44e-19
C10191 _331_/CLK _242_/a_109_257# 0.00287f
C10192 _279_/Y _315_/D 0.117f
C10193 _246_/B _325_/D 5.96e-19
C10194 output11/a_27_7# VPWR 0.158f
C10195 _254_/Y _191_/B 2.88e-21
C10196 _327_/a_761_249# _330_/Q 0.00126f
C10197 _316_/a_761_249# VPWR 0.025f
C10198 _316_/a_27_7# VGND -0.0745f
C10199 _343_/a_543_7# _229_/a_226_7# 0.00284f
C10200 _279_/Y _324_/a_651_373# 5.54e-21
C10201 _258_/S _309_/a_27_7# 0.00287f
C10202 _251_/a_215_7# _286_/Y 0.002f
C10203 _227_/A _333_/Q 0.16f
C10204 _216_/X _314_/D 0.118f
C10205 _221_/a_346_7# _286_/Y 0.00596f
C10206 input1/X _193_/Y 0.00114f
C10207 _320_/Q VPWR 6.34f
C10208 _228_/A _284_/A 0.00515f
C10209 _242_/A _331_/a_193_7# 7.36e-22
C10210 _326_/Q _222_/a_346_7# 3.2e-19
C10211 _180_/a_29_13# _215_/A 0.0024f
C10212 _255_/X clkbuf_0_clk/a_110_7# 4.22e-19
C10213 _313_/a_193_7# _336_/Q 9.13e-20
C10214 _313_/a_27_7# _225_/B 5.46e-20
C10215 _210_/a_27_7# _192_/B 3.17e-20
C10216 _327_/a_193_7# VPWR -0.273f
C10217 _317_/a_1283_n19# _232_/A 8.12e-19
C10218 _277_/A clkbuf_2_3_0_clk/A 1.96e-19
C10219 ctln[4] _340_/CLK 4.43e-20
C10220 _344_/a_796_7# _172_/B 5.54e-19
C10221 repeater43/X _315_/a_27_7# 0.0162f
C10222 _250_/a_493_257# _216_/A 2.83e-19
C10223 _250_/a_78_159# _250_/X 0.00183f
C10224 _337_/Q _283_/A 8.53e-20
C10225 _326_/a_193_7# VPWR -0.307f
C10226 _322_/a_193_7# _322_/Q 3.75e-19
C10227 _209_/X _225_/X 4.57e-19
C10228 _328_/a_193_7# _330_/Q 4.49e-21
C10229 ctlp[6] _320_/Q 1.06e-19
C10230 _277_/Y _319_/a_27_7# 9.47e-21
C10231 _345_/a_27_7# _163_/a_78_159# 2.45e-19
C10232 output12/a_27_7# ctln[6] 0.00328f
C10233 _294_/A _339_/Q 0.00224f
C10234 _157_/A _296_/a_109_7# 3.06e-21
C10235 output22/a_27_7# VGND 0.102f
C10236 _332_/a_651_373# VGND 7.23e-19
C10237 _332_/a_639_7# VPWR 6.43e-19
C10238 _327_/a_27_7# repeater42/a_27_7# 0.00661f
C10239 _331_/Q _214_/a_109_7# 0.00289f
C10240 _328_/a_27_7# VPWR 0.0463f
C10241 _347_/a_1270_373# VGND 9.31e-20
C10242 _221_/a_93_n19# _221_/a_250_257# -6.97e-22
C10243 _347_/a_805_7# VPWR 2.64e-19
C10244 _326_/a_805_7# _304_/X 3.87e-19
C10245 _340_/Q _267_/A 0.00531f
C10246 _194_/X _261_/A 1.71e-19
C10247 _200_/a_584_7# VPWR -7.15e-19
C10248 _285_/A trimb[4] 6.97e-19
C10249 _285_/A trim[1] 0.0356f
C10250 _200_/a_256_7# VGND -3.56e-20
C10251 repeater43/X _321_/a_1462_7# -8.37e-19
C10252 _326_/a_27_7# repeater42/a_27_7# 6.77e-21
C10253 _167_/X _260_/A 1.04e-19
C10254 _308_/S _286_/B 0.0284f
C10255 _336_/a_1283_n19# _313_/a_651_373# 1.43e-20
C10256 _328_/a_761_249# _297_/B 5.9e-20
C10257 _314_/Q _347_/a_651_373# 0.00302f
C10258 _297_/B _347_/a_1462_7# 3.77e-19
C10259 _314_/a_1217_7# _347_/D 1.56e-19
C10260 _216_/A _284_/A 0.641f
C10261 _321_/a_27_7# result[7] 5.06e-19
C10262 _258_/S _306_/a_76_159# 0.0293f
C10263 _164_/A _171_/a_78_159# 0.0556f
C10264 _322_/Q _246_/a_109_257# 3.08e-19
C10265 _343_/CLK _315_/a_1108_7# 0.0561f
C10266 _175_/Y _192_/B 1.31e-21
C10267 _346_/Q _166_/Y 0.451f
C10268 _346_/a_1032_373# _299_/X 0.00539f
C10269 _346_/a_193_7# _160_/X 3.45e-20
C10270 _169_/B _147_/A 3.1e-19
C10271 input4/X _153_/A 1.18e-20
C10272 _334_/a_27_7# VPWR 0.0782f
C10273 _277_/Y _338_/Q 0.00738f
C10274 _292_/A _311_/a_1283_n19# 0.0198f
C10275 _267_/B _265_/B 1.26e-19
C10276 _299_/X _331_/CLK 2.04e-20
C10277 _312_/Q _311_/a_1217_7# 2.56e-19
C10278 _186_/a_79_n19# _196_/A 1.59e-20
C10279 _344_/a_476_7# _162_/X 7.01e-21
C10280 _277_/Y _275_/A 0.659f
C10281 _307_/a_76_159# _227_/A 0.0105f
C10282 _323_/a_27_7# _298_/X 6.3e-19
C10283 _328_/a_651_373# _278_/a_68_257# 5.54e-22
C10284 _288_/A _311_/Q 3.39e-19
C10285 _255_/B _150_/a_27_7# 3.07e-20
C10286 _165_/X _267_/A 5.81e-20
C10287 clkbuf_2_3_0_clk/A _199_/a_584_7# 0.00103f
C10288 _341_/a_805_7# VGND -7.05e-19
C10289 _341_/a_1462_7# VPWR 2.15e-19
C10290 _254_/Y _337_/Q 6.52e-20
C10291 _273_/A _299_/X 0.153f
C10292 _338_/a_805_7# VGND 2.5e-19
C10293 _323_/a_543_7# _176_/a_27_7# 4.16e-19
C10294 _184_/a_439_7# _182_/X 0.00104f
C10295 _325_/a_1283_n19# _242_/A 4.84e-21
C10296 _287_/a_39_257# _311_/Q 0.00106f
C10297 _314_/a_193_7# _156_/a_39_257# 0.00423f
C10298 _206_/A _154_/A 0.391f
C10299 _207_/C _153_/A 0.112f
C10300 _339_/Q _283_/A 0.0785f
C10301 _325_/Q _183_/a_1241_257# 2.93e-20
C10302 _316_/Q _316_/a_1108_7# 0.0413f
C10303 _304_/S _314_/a_27_7# 8.01e-21
C10304 _329_/a_27_7# _281_/A 0.155f
C10305 _326_/a_1283_n19# _246_/B 0.00992f
C10306 _338_/Q _262_/a_199_7# 3.45e-19
C10307 _325_/a_1108_7# _325_/Q 1.17e-19
C10308 _346_/SET_B _314_/a_1462_7# 2.34e-21
C10309 _186_/a_297_7# _177_/A 1.94e-19
C10310 _226_/X _298_/A 1.07e-20
C10311 _271_/A _316_/a_651_373# 2.81e-21
C10312 _229_/a_226_257# VGND -3.01e-19
C10313 _346_/SET_B _324_/D 7.4e-21
C10314 _336_/a_639_7# _147_/A 1.24e-19
C10315 _295_/a_79_n19# VGND 0.0122f
C10316 _295_/a_306_7# VPWR -7.05e-19
C10317 _275_/A _304_/X 6.2e-21
C10318 _271_/A _204_/a_27_257# 2.71e-19
C10319 _346_/a_652_n19# VPWR 8.4e-19
C10320 _346_/a_27_7# VGND 0.0581f
C10321 _271_/Y _208_/a_78_159# 1.87e-19
C10322 _306_/S _336_/D 0.153f
C10323 _340_/a_1462_7# VGND -8.35e-19
C10324 _160_/X _173_/a_76_159# 0.0623f
C10325 _335_/a_27_7# _204_/a_27_257# 5.22e-20
C10326 _314_/a_193_7# _147_/A 1.43e-20
C10327 _316_/D _315_/D 1.88e-20
C10328 _318_/a_27_7# _248_/A 0.00333f
C10329 _345_/a_1602_7# _346_/SET_B 1.36e-20
C10330 _316_/a_1217_7# VGND -4.43e-19
C10331 _344_/a_1602_7# _164_/Y 9.14e-20
C10332 _346_/a_1182_221# _297_/B 5.3e-20
C10333 _340_/CLK _311_/a_27_7# 0.0248f
C10334 _276_/a_68_257# _242_/A 0.00916f
C10335 _342_/Q _324_/Q 0.0795f
C10336 _207_/X VPWR 0.12f
C10337 _346_/SET_B _309_/Q -7.64e-19
C10338 _318_/a_27_7# _331_/CLK 0.0278f
C10339 _201_/a_27_7# VPWR 0.135f
C10340 _327_/a_805_7# VGND -7.08e-19
C10341 _327_/a_1462_7# VPWR 1.61e-19
C10342 _324_/Q _144_/a_27_7# 9.01e-19
C10343 repeater43/X _242_/B 0.0117f
C10344 _277_/Y _345_/D 4.04e-20
C10345 _195_/a_373_7# _340_/D 4.91e-19
C10346 _346_/SET_B _279_/A 0.0541f
C10347 _326_/a_1462_7# VPWR 4.71e-20
C10348 _326_/a_805_7# VGND 5.65e-19
C10349 _194_/X _340_/Q 0.41f
C10350 _215_/A _313_/a_1108_7# 0.0476f
C10351 clk _153_/a_215_257# 0.0155f
C10352 output14/a_27_7# _322_/a_27_7# 6.26e-19
C10353 _254_/A _300_/a_301_257# 0.00322f
C10354 repeater43/X _324_/a_193_7# -0.00451f
C10355 _254_/Y _339_/Q 1.3e-20
C10356 _281_/Y _340_/D 2.46e-20
C10357 clk _209_/X 0.00549f
C10358 _345_/a_193_7# _158_/Y 1.25e-19
C10359 _277_/Y _313_/a_1108_7# 8.9e-37
C10360 _181_/X _181_/a_27_7# 0.00288f
C10361 _149_/A _154_/A 3.32e-19
C10362 _218_/a_250_257# _346_/SET_B 2.33e-19
C10363 _227_/A _212_/X 8.73e-20
C10364 _180_/a_29_13# VGND 0.0573f
C10365 _180_/a_183_257# VPWR -6.6e-19
C10366 _343_/a_27_7# repeater43/X 0.0165f
C10367 _303_/A _248_/B 3.94e-19
C10368 _328_/a_1217_7# VPWR 1.35e-20
C10369 _328_/a_639_7# VGND -0.00153f
C10370 _251_/X _221_/a_93_n19# 9.64e-21
C10371 _298_/B _191_/B 4.03e-20
C10372 clkbuf_2_1_0_clk/A _267_/B 7.98e-21
C10373 _341_/Q _192_/B 1.81e-19
C10374 _173_/a_226_7# VPWR 0.0187f
C10375 _221_/a_346_7# _328_/Q 6.65e-19
C10376 _177_/a_27_7# _244_/B 0.0418f
C10377 _181_/X _214_/a_373_7# 2.96e-19
C10378 _254_/A _215_/A 0.00914f
C10379 _294_/Y _284_/A 0.33f
C10380 _271_/A _334_/a_1108_7# 0.0534f
C10381 _319_/a_761_249# VPWR 0.0146f
C10382 _319_/a_27_7# VGND 0.0342f
C10383 _345_/a_27_7# clkbuf_2_3_0_clk/A 3.65e-21
C10384 _337_/a_27_7# VPWR 0.0689f
C10385 _346_/SET_B _311_/a_193_7# 0.024f
C10386 _335_/a_193_7# _334_/a_1283_n19# 2.34e-21
C10387 _277_/Y _254_/A 0.00487f
C10388 _321_/a_1217_7# result[7] 2.89e-20
C10389 _248_/A _246_/B 0.446f
C10390 _164_/A _172_/B 0.478f
C10391 _267_/B _310_/Q 0.031f
C10392 _258_/S _258_/a_218_334# 0.0034f
C10393 _219_/a_93_n19# _242_/A 1.53e-21
C10394 _319_/a_1283_n19# _297_/B 1.46e-20
C10395 _341_/D _271_/A 0.0106f
C10396 _313_/D _286_/B 0.0263f
C10397 _343_/CLK output6/a_27_7# 0.00269f
C10398 _334_/a_639_7# VGND -0.00169f
C10399 _334_/a_1217_7# VPWR 1.62e-19
C10400 clk _209_/a_109_257# 2.97e-19
C10401 _167_/a_109_257# _346_/Q 0.00402f
C10402 _255_/a_30_13# _306_/S 3.52e-19
C10403 _331_/CLK _246_/B 0.0885f
C10404 _323_/D _177_/a_27_7# 3.91e-20
C10405 _320_/Q _320_/a_543_7# 2.9e-19
C10406 _238_/B _320_/a_27_7# 9.27e-20
C10407 _216_/a_27_7# _314_/D 2.09e-20
C10408 _200_/a_93_n19# _293_/a_39_257# 1.5e-20
C10409 output12/a_27_7# _255_/X 1.64e-20
C10410 _345_/a_1182_221# _345_/Q 0.0368f
C10411 _345_/a_476_7# _345_/D 0.00316f
C10412 _345_/a_27_7# _172_/Y 9.95e-20
C10413 _316_/Q _248_/A 0.00649f
C10414 input4/a_27_7# _195_/a_27_257# 1.13e-19
C10415 _179_/a_27_7# _333_/D 4.45e-20
C10416 _325_/a_1108_7# _326_/Q 0.00674f
C10417 _324_/a_1283_n19# _304_/S 0.0826f
C10418 _283_/Y _332_/a_543_7# 1.64e-20
C10419 _286_/B _197_/X 0.00511f
C10420 _258_/S _198_/a_93_n19# 3.7e-21
C10421 _273_/A _246_/B 3.15e-19
C10422 _344_/D _297_/Y 0.0135f
C10423 _342_/Q _228_/A 0.0187f
C10424 input1/a_75_172# _199_/a_250_257# 2.98e-21
C10425 _258_/a_76_159# _260_/B 5.59e-19
C10426 _338_/Q VGND 0.954f
C10427 _167_/X _165_/X 0.329f
C10428 _275_/A VGND 0.784f
C10429 _316_/Q _331_/CLK 0.11f
C10430 _215_/A _309_/D 6.62e-20
C10431 _329_/a_1217_7# _281_/A 3.71e-19
C10432 _285_/Y _162_/A 0.135f
C10433 _346_/Q _297_/Y 5.23e-20
C10434 _277_/Y _309_/D 0.103f
C10435 _329_/a_1270_373# _281_/Y 1.39e-19
C10436 _340_/a_543_7# _198_/a_93_n19# 0.00302f
C10437 _342_/a_1108_7# _177_/A 1.12e-19
C10438 _271_/A _236_/B 0.535f
C10439 _226_/a_79_n19# VPWR 0.0201f
C10440 _188_/a_535_334# VGND -2.78e-19
C10441 _188_/a_439_7# VPWR -2.67e-19
C10442 _342_/a_193_7# valid 9.91e-19
C10443 _325_/a_193_7# _227_/A 1.1e-19
C10444 _292_/A _171_/a_78_159# 0.00892f
C10445 _346_/a_586_7# VGND -8.32e-19
C10446 _322_/Q _331_/Q 0.0408f
C10447 _333_/a_193_7# _333_/a_651_373# -0.00701f
C10448 _308_/X _298_/C 0.0127f
C10449 _335_/a_1283_n19# _332_/Q 7.71e-19
C10450 ctln[5] _153_/B 1.16e-19
C10451 _158_/Y VPWR 0.191f
C10452 _309_/a_1108_7# _346_/SET_B -0.0235f
C10453 _335_/a_1108_7# _207_/X 0.0195f
C10454 _342_/a_761_249# _343_/Q 4.47e-21
C10455 _342_/a_27_7# _298_/C 5.55e-21
C10456 _343_/a_1283_n19# _147_/A 2.59e-19
C10457 _343_/a_193_7# _226_/X 1.14e-19
C10458 _318_/a_1217_7# _248_/A 6.84e-20
C10459 _341_/a_27_7# _244_/B 0.00878f
C10460 _339_/a_27_7# VPWR 0.0783f
C10461 _267_/A _310_/a_448_7# 3.11e-19
C10462 _327_/a_27_7# _232_/X 0.0373f
C10463 _339_/Q _336_/a_1108_7# 1.25e-19
C10464 _271_/A _143_/a_27_7# 0.00778f
C10465 _150_/C _217_/A 8.04e-23
C10466 _252_/a_27_7# _297_/A 0.00441f
C10467 _342_/Q _216_/A 0.0503f
C10468 _255_/B _250_/X 8.18e-19
C10469 _343_/a_1283_n19# _149_/A 0.0055f
C10470 _187_/a_27_7# _144_/A 0.00167f
C10471 _169_/Y _174_/a_27_257# 5.79e-20
C10472 _323_/a_1108_7# _334_/a_27_7# 2.13e-21
C10473 _323_/a_1283_n19# _334_/a_193_7# 9.09e-19
C10474 _329_/a_1270_373# _329_/D 2.49e-19
C10475 _326_/a_27_7# _232_/X 0.00785f
C10476 _336_/a_651_373# _202_/a_93_n19# 7.47e-20
C10477 _216_/A _144_/a_27_7# 0.00152f
C10478 _144_/A _315_/D 0.00584f
C10479 _337_/Q _194_/a_27_7# 0.0371f
C10480 _330_/Q _327_/Q 0.0032f
C10481 _341_/a_27_7# _323_/D 1.83e-22
C10482 input1/X _298_/A 0.00454f
C10483 _312_/a_761_249# _312_/D 2.33e-20
C10484 _254_/A _300_/Y 0.00165f
C10485 cal input3/a_27_7# 0.00367f
C10486 repeater43/X _324_/a_1462_7# -8.59e-19
C10487 _317_/a_193_7# _217_/A 6.04e-21
C10488 input1/X _336_/a_448_7# 0.0139f
C10489 ctlp[3] ctlp[4] 6.04e-20
C10490 _340_/a_27_7# _254_/B 0.00251f
C10491 repeater43/X _318_/a_1283_n19# 0.047f
C10492 _343_/a_1217_7# repeater43/X 5.1e-19
C10493 _316_/a_193_7# _244_/B 0.016f
C10494 _329_/a_193_7# _329_/a_448_7# -0.00779f
C10495 _254_/Y _336_/D 0.0208f
C10496 _329_/a_761_249# _327_/D 5.8e-20
C10497 _346_/Q _242_/A 1.35e-20
C10498 _345_/D VGND 0.119f
C10499 _341_/Q _146_/C 0.407f
C10500 _290_/A _310_/a_27_7# 0.00413f
C10501 _306_/X _194_/A 1.41e-19
C10502 _297_/B _212_/X 0.0751f
C10503 _319_/a_1217_7# VGND -4.3e-19
C10504 _331_/a_1108_7# _304_/X 0.00108f
C10505 _331_/a_1283_n19# _217_/A 0.00192f
C10506 _313_/a_1108_7# VGND 0.0241f
C10507 _271_/A _343_/CLK 0.0569f
C10508 _313_/a_651_373# VPWR -0.00912f
C10509 _181_/X _330_/a_543_7# 1.53e-20
C10510 repeater42/a_27_7# repeater43/X 0.018f
C10511 _323_/a_761_249# _248_/A 6.42e-22
C10512 _292_/Y _290_/Y 0.157f
C10513 _337_/a_1217_7# VPWR 9.35e-20
C10514 _337_/a_639_7# VGND -0.00131f
C10515 _328_/a_1283_n19# output19/a_27_7# 0.00171f
C10516 _335_/a_27_7# _343_/CLK 0.0152f
C10517 ctln[7] _208_/a_78_159# 6.49e-21
C10518 _342_/a_1108_7# _341_/a_1283_n19# 8.54e-21
C10519 _342_/a_1283_n19# _341_/a_1108_7# 1.21e-19
C10520 _342_/a_651_373# _341_/a_761_249# 4.5e-21
C10521 _298_/C _203_/a_209_7# 0.00189f
C10522 result[5] _331_/CLK 0.194f
C10523 _255_/a_30_13# _283_/A 4.06e-22
C10524 clkbuf_1_0_0_clk/a_75_172# _283_/A 7.43e-19
C10525 output31/a_27_7# output33/a_27_7# 5.46e-20
C10526 _298_/C _254_/B 0.109f
C10527 _301_/X _170_/a_76_159# 0.0115f
C10528 _258_/S _306_/X 0.035f
C10529 _286_/B _333_/a_193_7# 5.86e-22
C10530 _320_/a_27_7# _331_/CLK 1.62e-21
C10531 _320_/Q _322_/a_651_373# 0.0268f
C10532 cal _153_/A 0.0134f
C10533 _336_/a_1283_n19# _267_/A 2.28e-22
C10534 _145_/A _315_/D 1.19e-19
C10535 _197_/X _338_/a_1108_7# 1.9e-21
C10536 _298_/A _286_/Y 0.123f
C10537 _345_/a_1296_7# _345_/Q 3.55e-19
C10538 _254_/A VGND 1.4f
C10539 _157_/a_27_7# VPWR 0.12f
C10540 clkbuf_2_3_0_clk/A clkbuf_2_1_0_clk/a_75_172# 0.0419f
C10541 _167_/X _301_/a_245_257# 9.68e-19
C10542 _165_/X _301_/a_51_257# 3.9e-19
C10543 clkbuf_0_clk/X _215_/A 0.02f
C10544 _308_/X _229_/a_489_373# 1.36e-20
C10545 rstn _194_/X 0.151f
C10546 _165_/X clkbuf_1_1_0_clk/a_75_172# 7.88e-21
C10547 _301_/X clkbuf_2_1_0_clk/A 1.39e-19
C10548 _339_/Q _194_/a_27_7# 7.44e-22
C10549 _172_/A _295_/a_676_257# 8.31e-21
C10550 _267_/B _311_/a_27_7# 2.36e-19
C10551 _342_/a_761_249# _229_/a_76_159# 2.51e-19
C10552 _342_/a_193_7# _229_/a_226_7# 3.8e-19
C10553 _277_/Y clkbuf_0_clk/X 0.0113f
C10554 _313_/D _279_/Y 2.97e-20
C10555 _210_/a_307_257# _306_/S 4.83e-19
C10556 _323_/Q VPWR 0.711f
C10557 repeater43/a_27_7# _323_/a_193_7# 2.51e-22
C10558 _319_/Q _321_/a_1108_7# 7.57e-19
C10559 _288_/A _164_/Y 2.53e-19
C10560 _340_/a_651_373# _197_/X 0.00109f
C10561 _218_/a_584_7# _217_/X 0.00205f
C10562 _325_/a_543_7# _315_/D 2.87e-21
C10563 _246_/B _217_/X 1.5e-19
C10564 _226_/X VGND 0.281f
C10565 _164_/Y _162_/X 0.449f
C10566 _302_/a_227_257# _300_/Y 0.00148f
C10567 _279_/Y _197_/X 0.0909f
C10568 _236_/B _232_/a_27_7# 0.0411f
C10569 _292_/A _172_/B 2.77e-19
C10570 _305_/a_76_159# _340_/CLK 0.00155f
C10571 _283_/Y _334_/a_1108_7# 2.26e-21
C10572 _320_/a_543_7# _319_/a_761_249# 2.05e-21
C10573 _320_/a_1283_n19# _319_/a_193_7# 1.97e-20
C10574 _320_/a_1108_7# _319_/a_27_7# 6.18e-19
C10575 _320_/a_761_249# _319_/a_543_7# 2.04e-21
C10576 _320_/a_27_7# _319_/a_1108_7# 7.23e-19
C10577 _333_/a_761_249# _333_/D 0.00216f
C10578 _160_/a_27_7# VPWR 0.126f
C10579 _194_/A _147_/Y 0.00364f
C10580 _290_/A output36/a_27_7# 2.6e-19
C10581 _309_/D VGND 0.087f
C10582 _160_/A _172_/B 1.15e-20
C10583 _343_/a_1462_7# _226_/X 1.19e-19
C10584 _215_/A input1/X 3.34e-20
C10585 _339_/a_1217_7# VPWR 9.01e-20
C10586 _339_/a_639_7# VGND -0.00153f
C10587 _183_/a_471_7# _217_/A 6.48e-22
C10588 _327_/a_1217_7# _232_/X 1.21e-19
C10589 _267_/A _310_/D 0.0174f
C10590 _181_/X _331_/Q 0.0207f
C10591 clkbuf_0_clk/X _304_/X 0.00415f
C10592 _277_/Y input1/X 1.59e-19
C10593 _325_/a_651_373# _217_/A 0.0018f
C10594 _325_/a_1108_7# _324_/D 2.2e-20
C10595 output5/a_27_7# clkc 0.00847f
C10596 _317_/a_1283_n19# VPWR 0.0465f
C10597 _317_/a_761_249# VGND -3.61e-19
C10598 _299_/a_78_159# _299_/a_292_257# -1.09e-21
C10599 _323_/a_27_7# _343_/CLK 0.361f
C10600 _182_/a_215_7# _286_/B 0.00944f
C10601 _182_/a_79_n19# _181_/X 0.00924f
C10602 _258_/S _147_/Y 0.00636f
C10603 _283_/Y _338_/D 0.183f
C10604 _326_/a_1217_7# _232_/X 3.21e-20
C10605 _317_/Q _269_/A 0.0145f
C10606 repeater43/X _335_/a_448_7# -2.34e-19
C10607 _271_/A output29/a_27_7# 7.89e-19
C10608 _258_/S _312_/a_1108_7# 1.48e-21
C10609 _330_/Q _331_/a_1270_373# 1.04e-19
C10610 _172_/A _173_/a_76_159# 0.00308f
C10611 _337_/D _311_/a_193_7# 5.61e-21
C10612 _228_/A _225_/B 3.66e-20
C10613 _292_/A _312_/a_761_249# 6.94e-19
C10614 _248_/A _244_/a_109_257# 0.00285f
C10615 _309_/a_1283_n19# _267_/B 3.39e-20
C10616 _309_/a_761_249# _309_/D 4.29e-21
C10617 _340_/a_543_7# _147_/Y 4.68e-21
C10618 _328_/a_805_7# _232_/X 1.12e-19
C10619 _331_/a_1108_7# VGND 0.0324f
C10620 _331_/a_651_373# VPWR 0.00329f
C10621 result[7] VPWR 0.244f
C10622 _320_/a_1270_373# _346_/SET_B -2.06e-19
C10623 _196_/A _162_/X 0.0046f
C10624 _302_/a_227_257# VGND -5.05e-19
C10625 _302_/a_539_257# VPWR -3.64e-19
C10626 comp clkc 0.0262f
C10627 _214_/a_373_7# _346_/SET_B 2.82e-20
C10628 _344_/a_1032_373# _346_/SET_B -0.0049f
C10629 _316_/a_805_7# _317_/D 4.26e-19
C10630 _343_/a_761_249# cal 0.00455f
C10631 _343_/a_193_7# input1/X 0.00125f
C10632 _290_/A _310_/a_1217_7# 2.56e-19
C10633 _336_/a_761_249# _306_/S 2.67e-20
C10634 _336_/a_543_7# _340_/Q 3.78e-20
C10635 _336_/a_1283_n19# _194_/X 0.00818f
C10636 _336_/a_193_7# _193_/Y 0.00102f
C10637 _206_/A _153_/B 0.806f
C10638 _302_/a_77_159# _314_/Q 0.0149f
C10639 _292_/A _289_/a_121_257# 7.79e-19
C10640 _215_/A _286_/Y 0.866f
C10641 _294_/A output31/a_27_7# 0.0341f
C10642 ctln[7] _190_/A 1.03e-19
C10643 _335_/a_805_7# _334_/D 3.76e-20
C10644 _182_/a_79_n19# _343_/Q 1.62e-20
C10645 _342_/a_543_7# _341_/D 5.07e-22
C10646 _306_/S _260_/a_27_257# 3.06e-20
C10647 _322_/a_27_7# _321_/D 3.39e-19
C10648 _322_/a_1283_n19# _331_/CLK 0.0084f
C10649 _277_/Y _286_/Y 0.0159f
C10650 _325_/a_761_249# _246_/B 4.66e-20
C10651 _270_/a_121_257# _232_/A 8.63e-19
C10652 _342_/D _341_/a_543_7# 1.32e-20
C10653 ctln[1] _335_/a_1283_n19# 4.73e-20
C10654 _179_/a_27_7# _190_/A 3.92e-20
C10655 _169_/Y _216_/A 5.23e-20
C10656 _216_/A _225_/B 0.0233f
C10657 _162_/a_27_7# VGND 0.133f
C10658 clkbuf_0_clk/X _220_/a_93_n19# 7.29e-19
C10659 _177_/a_27_7# _177_/A 0.0152f
C10660 _277_/A _165_/X 7.84e-20
C10661 _271_/A _146_/a_184_13# 1.44e-20
C10662 _250_/a_215_7# _215_/A 0.00122f
C10663 _255_/B _325_/Q 6.89e-20
C10664 _324_/a_761_249# _286_/Y 0.00706f
C10665 _267_/B _311_/a_1217_7# 1.56e-19
C10666 _342_/a_1108_7# _248_/A 0.00541f
C10667 _300_/a_383_7# _284_/A 5.93e-19
C10668 _309_/a_193_7# _337_/Q 8.78e-20
C10669 _327_/a_639_7# _331_/D 8.22e-21
C10670 clkbuf_2_0_0_clk/a_75_172# _194_/X 6.32e-22
C10671 _166_/Y _170_/a_76_159# 1.87e-19
C10672 _285_/A _288_/Y 0.0225f
C10673 repeater43/X _323_/a_448_7# 7.47e-21
C10674 _343_/a_193_7# _286_/Y 9.16e-20
C10675 _187_/a_27_7# _324_/Q 0.00812f
C10676 _281_/Y clkbuf_2_1_0_clk/A 6.44e-20
C10677 result[4] _242_/B 0.00425f
C10678 _192_/a_68_257# _305_/X 0.0165f
C10679 _304_/X _286_/Y 0.0173f
C10680 _307_/X _184_/a_439_7# 1.67e-20
C10681 _324_/Q _315_/D 0.015f
C10682 _330_/D _331_/a_193_7# 4.15e-19
C10683 _320_/a_193_7# _212_/X 1.31e-20
C10684 _320_/a_27_7# _217_/X 4.56e-21
C10685 _162_/X _347_/a_1283_n19# 1.37e-20
C10686 _306_/X _201_/a_27_7# 4.06e-21
C10687 _324_/a_651_373# _324_/Q 3.05e-19
C10688 clkbuf_0_clk/X VGND 1.4f
C10689 clkbuf_2_3_0_clk/A _311_/D 0.0062f
C10690 _211_/a_27_257# _339_/a_27_7# 4.74e-21
C10691 _325_/a_1270_373# VGND 1.86e-19
C10692 _166_/Y clkbuf_2_1_0_clk/A 0.245f
C10693 _339_/a_27_7# _198_/a_93_n19# 4.18e-22
C10694 _283_/Y _343_/CLK 4.37f
C10695 _157_/A _314_/D 1.41e-19
C10696 _344_/a_476_7# _345_/Q 4.67e-20
C10697 _320_/D _319_/a_193_7# 2.25e-20
C10698 _324_/a_27_7# _221_/a_93_n19# 2.47e-20
C10699 repeater43/X _172_/A 1.9e-20
C10700 _340_/D _336_/Q 5.53e-20
C10701 _329_/D clkbuf_2_1_0_clk/A 2.67e-20
C10702 _202_/a_346_7# VPWR -9.07e-19
C10703 _202_/a_250_257# VGND 5.69e-19
C10704 repeater43/X _335_/D 0.158f
C10705 repeater43/X _232_/X 0.0852f
C10706 _297_/A _347_/a_639_7# 0.00466f
C10707 _315_/Q _342_/D 1.72e-21
C10708 _313_/D _313_/a_27_7# 0.0514f
C10709 _219_/a_250_257# _279_/A 0.00527f
C10710 _294_/A _291_/a_39_257# 1.53e-19
C10711 _273_/A _172_/B 0.188f
C10712 _341_/a_27_7# _177_/A 3.3e-20
C10713 _308_/X _207_/C 5.36e-19
C10714 _300_/Y _286_/Y 1.3e-20
C10715 _340_/a_27_7# _196_/A 0.0625f
C10716 input1/X VGND 0.926f
C10717 _308_/S _145_/A 0.106f
C10718 _292_/A trimb[4] 4.11e-20
C10719 trim[1] _292_/A 4.2e-20
C10720 _346_/a_652_n19# _147_/Y 1.04e-20
C10721 _300_/Y _297_/a_27_257# 8.99e-19
C10722 _269_/A _315_/a_193_7# 0.0171f
C10723 _269_/A _298_/A 1.18e-19
C10724 _323_/a_1108_7# _323_/Q 0.0499f
C10725 _323_/a_1283_n19# _192_/B 5.55e-19
C10726 _197_/X _337_/a_1283_n19# 7.4e-19
C10727 _232_/A _243_/a_113_257# 0.0686f
C10728 _342_/a_543_7# _343_/CLK 1.66e-19
C10729 _227_/A _306_/S 0.0444f
C10730 _212_/a_27_7# _327_/Q 0.0655f
C10731 _283_/Y _339_/a_1108_7# 1.48e-19
C10732 _265_/B _297_/Y 0.00721f
C10733 _342_/Q _209_/a_27_257# 1.97e-19
C10734 _277_/Y _240_/B 9.49e-20
C10735 _323_/a_651_373# _226_/X 1.92e-21
C10736 _147_/Y _201_/a_27_7# 6.62e-19
C10737 _275_/A _318_/Q 5.92e-19
C10738 _187_/a_27_7# _228_/A 6.4e-22
C10739 _211_/a_109_257# _334_/Q 1.72e-20
C10740 _335_/D _334_/Q 0.0117f
C10741 _182_/X _343_/Q 8.42e-21
C10742 _305_/a_505_n19# _147_/A 6.61e-21
C10743 _165_/a_215_7# _164_/Y 0.0282f
C10744 _315_/D _228_/A 0.00842f
C10745 _196_/A _298_/C 0.00836f
C10746 output14/a_27_7# ctlp[1] 1.68e-21
C10747 _323_/a_805_7# _149_/A 5.73e-20
C10748 _234_/B _242_/A 0.0154f
C10749 _324_/a_651_373# _228_/A 0.00227f
C10750 _255_/B _326_/Q 1.44e-20
C10751 _297_/B _344_/Q 0.0106f
C10752 _172_/A _191_/B 0.00735f
C10753 _267_/A VPWR 2.13f
C10754 _321_/a_1283_n19# _242_/A 1.2e-21
C10755 repeater43/X _244_/B 0.443f
C10756 _265_/B _310_/a_193_7# 1.18e-19
C10757 _316_/D _330_/a_1108_7# 9.6e-20
C10758 _331_/CLK _330_/a_448_7# 0.00567f
C10759 VGND _286_/Y 3.89f
C10760 VPWR sample 0.268f
C10761 _308_/X _150_/C 0.0562f
C10762 _335_/D _191_/B 0.02f
C10763 _188_/S _192_/B 1.3e-19
C10764 _173_/a_226_7# _147_/Y 0.0402f
C10765 _297_/a_27_257# VGND -0.00253f
C10766 _184_/a_76_159# _146_/C 1.67e-20
C10767 _219_/a_584_7# VGND 5.26e-19
C10768 _239_/a_199_7# _297_/B 2.45e-19
C10769 _309_/a_651_373# _174_/a_27_257# 3.05e-20
C10770 repeater43/X _322_/a_1270_373# -3.58e-20
C10771 _346_/a_193_7# _297_/A 4.11e-20
C10772 _345_/a_381_7# _344_/D 1.53e-19
C10773 _153_/a_109_53# _204_/Y 1.58e-20
C10774 _153_/a_215_257# _335_/Q 0.0199f
C10775 _342_/Q _315_/a_761_249# 5.12e-21
C10776 _343_/Q valid 3.74e-19
C10777 _298_/C _298_/X 0.0875f
C10778 _209_/X _335_/Q 1.57e-20
C10779 _254_/B _207_/C 0.0464f
C10780 _313_/a_1283_n19# _254_/B 4.59e-21
C10781 repeater43/X _323_/D 0.00784f
C10782 _277_/Y _328_/Q 7.2e-21
C10783 _333_/a_761_249# _190_/A 0.00357f
C10784 _333_/a_543_7# _333_/Q 3.11e-20
C10785 _333_/a_1283_n19# _332_/Q 0.00739f
C10786 _254_/Y _336_/a_761_249# 0.0188f
C10787 _345_/a_381_7# _346_/Q 1.82e-21
C10788 _187_/a_27_7# _216_/A 1.31e-19
C10789 _341_/a_193_7# _341_/a_543_7# -0.011f
C10790 _341_/a_27_7# _341_/a_1283_n19# -1.43e-19
C10791 _309_/a_27_7# _267_/A 1.72e-19
C10792 _216_/A _315_/D 0.0191f
C10793 _330_/Q _221_/a_250_257# 2.47e-21
C10794 _255_/B _314_/a_193_7# 4.03e-20
C10795 _250_/a_215_7# VGND 0.0307f
C10796 _234_/B _322_/D 0.00544f
C10797 _324_/a_651_373# _216_/A 3.69e-19
C10798 _324_/a_1108_7# _250_/X 1.06e-20
C10799 _313_/Q clkbuf_2_3_0_clk/A 2.52e-20
C10800 _197_/X _339_/a_1283_n19# 2.62e-20
C10801 _314_/a_27_7# _297_/Y 9.19e-21
C10802 ctlp[4] _346_/SET_B 0.00351f
C10803 _345_/a_27_7# _165_/X 2.07e-19
C10804 _345_/a_193_7# _167_/X 2.35e-20
C10805 _285_/A _337_/Q -1.05e-36
C10806 _167_/a_109_257# clkbuf_2_1_0_clk/A 4.75e-19
C10807 _227_/A _327_/D 2.36e-21
C10808 _338_/a_193_7# _338_/a_543_7# -0.0231f
C10809 _331_/Q _346_/SET_B 4.33e-20
C10810 _221_/a_93_n19# VPWR 0.0224f
C10811 result[4] _318_/a_1283_n19# 4.55e-20
C10812 _347_/Q _306_/S 1.89e-20
C10813 _344_/a_1224_7# _345_/Q 2.97e-19
C10814 _281_/Y _218_/a_93_n19# 0.00887f
C10815 _339_/D _153_/B 0.0019f
C10816 _170_/a_76_159# _297_/Y 2.62e-20
C10817 _189_/a_27_7# _154_/A 1.49e-19
C10818 _231_/a_79_n19# _343_/CLK 1.14e-19
C10819 _250_/X _324_/D 1.19e-21
C10820 _342_/a_639_7# repeater43/X -7.75e-19
C10821 _314_/D _221_/a_250_257# 1.04e-20
C10822 _319_/Q _279_/A 0.00753f
C10823 _209_/a_109_257# _335_/Q 1.51e-20
C10824 _191_/B _203_/a_80_n19# 0.00876f
C10825 _342_/Q _153_/A 6.99e-21
C10826 _255_/B _154_/A 4.24e-21
C10827 _346_/SET_B _312_/a_805_7# 5.66e-19
C10828 _340_/a_1108_7# _194_/A 1.24e-20
C10829 _329_/a_27_7# _217_/A 2.29e-19
C10830 _329_/a_193_7# _304_/X 7.4e-19
C10831 _304_/X _328_/Q 0.00369f
C10832 output32/a_27_7# _338_/Q 2.03e-19
C10833 _332_/a_1283_n19# _332_/a_1108_7# 2.84e-32
C10834 _184_/a_218_7# cal 5.88e-20
C10835 _184_/a_535_334# input1/X 7.48e-19
C10836 _232_/X _331_/a_448_7# 0.00141f
C10837 _240_/B _300_/Y 3.74e-20
C10838 clkbuf_2_1_0_clk/A _297_/Y 0.00595f
C10839 output34/a_27_7# _292_/A 0.035f
C10840 _341_/Q _232_/A 0.0166f
C10841 _323_/a_27_7# output30/a_27_7# 4.04e-20
C10842 _286_/B _295_/a_79_n19# 0.00338f
C10843 _169_/Y _301_/a_240_7# 0.0057f
C10844 _314_/Q _284_/A 1.61e-20
C10845 _317_/D _150_/C 2.98e-19
C10846 _346_/a_27_7# _286_/B 1.52e-20
C10847 _325_/Q _326_/Q 0.289f
C10848 _290_/A _309_/Q 1.61e-20
C10849 _172_/A _337_/Q 0.0016f
C10850 _329_/D _218_/a_93_n19# 1.97e-19
C10851 _164_/A _173_/a_76_159# 9.18e-20
C10852 _267_/A _311_/a_651_373# 0.00269f
C10853 _261_/A _311_/a_448_7# 6.06e-21
C10854 _227_/A _283_/A 0.0252f
C10855 _269_/A _315_/a_1462_7# 4.06e-19
C10856 _343_/CLK _333_/a_27_7# 0.0375f
C10857 _310_/Q _297_/Y 0.031f
C10858 _258_/S _260_/B 0.0732f
C10859 ctlp[0] _320_/Q 0.00734f
C10860 _158_/Y _147_/Y 4.71e-22
C10861 result[2] _315_/a_1108_7# 0.00129f
C10862 _194_/X VPWR 1.06f
C10863 _275_/Y _344_/Q 0.0149f
C10864 output35/a_27_7# _164_/Y 3.06e-19
C10865 _306_/X _157_/a_27_7# 5.02e-19
C10866 _337_/Q _198_/a_250_257# 0.00416f
C10867 _309_/a_543_7# _284_/A 0.0337f
C10868 _227_/A _205_/a_382_257# 4.67e-19
C10869 clkbuf_2_1_0_clk/A _310_/a_193_7# 1.08e-20
C10870 _270_/a_39_257# _242_/B 3.49e-20
C10871 ctln[6] VGND 0.3f
C10872 _343_/a_193_7# _269_/A 0.0146f
C10873 _279_/Y _340_/a_193_7# 0.00235f
C10874 _317_/a_543_7# _244_/B 0.00109f
C10875 _317_/a_193_7# _317_/D 0.0656f
C10876 _177_/a_27_7# _248_/A 0.0513f
C10877 _342_/a_1283_n19# _145_/A 7.77e-19
C10878 _229_/a_76_159# valid 2.85e-19
C10879 _306_/S _297_/B 0.00989f
C10880 _308_/S _324_/Q 0.00271f
C10881 ctln[3] _267_/A 1.21e-19
C10882 _315_/Q _341_/a_193_7# 4.15e-22
C10883 _316_/a_27_7# _316_/a_448_7# -0.00676f
C10884 _310_/a_1108_7# _310_/D 0.0579f
C10885 _310_/a_193_7# _310_/Q 2.21e-19
C10886 _326_/a_1270_373# _181_/X 6.96e-21
C10887 _346_/SET_B _299_/a_292_257# 5.81e-20
C10888 _329_/Q _216_/X 0.0395f
C10889 _233_/a_113_257# _327_/Q 2.77e-20
C10890 _255_/X _215_/A 5.23e-20
C10891 _273_/A trimb[4] 1.23e-19
C10892 trim[1] _273_/A 3.38e-19
C10893 _300_/Y _328_/Q 9.83e-20
C10894 _232_/A _315_/a_639_7# 5.52e-20
C10895 _209_/X _209_/a_373_7# -1.67e-20
C10896 _336_/a_193_7# _336_/a_448_7# -0.00779f
C10897 _327_/a_761_249# _216_/X 2.39e-20
C10898 _227_/A _248_/B 0.0157f
C10899 _240_/B VGND 0.0895f
C10900 _290_/A _311_/a_193_7# 2.68e-19
C10901 _325_/Q _224_/a_256_7# 0.00128f
C10902 _196_/A _332_/D 9.13e-20
C10903 _167_/X VPWR 0.359f
C10904 _343_/a_193_7# _343_/D 0.0584f
C10905 _343_/a_543_7# _185_/A 0.0118f
C10906 _327_/a_761_249# _329_/Q 6.8e-21
C10907 _327_/a_27_7# _238_/B 2.21e-21
C10908 _188_/S _146_/C 0.0113f
C10909 _309_/a_448_7# _344_/D 1.46e-19
C10910 _182_/a_79_n19# _206_/A 4.1e-23
C10911 _153_/A _204_/Y 1.84e-21
C10912 _327_/a_193_7# _327_/a_543_7# -0.0156f
C10913 clkbuf_2_1_0_clk/A _242_/A 0.0182f
C10914 _255_/a_112_257# VPWR 9.73e-21
C10915 result[3] _317_/a_27_7# 6.27e-19
C10916 _318_/Q _317_/a_761_249# 7.38e-22
C10917 _188_/S _157_/A 0.00349f
C10918 _324_/a_1108_7# _255_/B 2.38e-19
C10919 _323_/a_1270_373# cal 5.18e-20
C10920 _306_/a_535_334# _284_/A 7.28e-19
C10921 _328_/a_193_7# _216_/X 5.54e-19
C10922 _315_/Q _316_/a_761_249# 1.06e-19
C10923 _329_/a_1283_n19# _330_/Q 0.00346f
C10924 _268_/a_121_257# _248_/A 1.05e-19
C10925 repeater43/X _330_/a_805_7# 5.66e-19
C10926 trim[1] trim[4] 0.0329f
C10927 _331_/a_193_7# _330_/a_1283_n19# 4.08e-19
C10928 _331_/a_27_7# _330_/a_1108_7# 2.59e-21
C10929 _332_/a_27_7# _207_/X 1.31e-21
C10930 _332_/a_1108_7# _208_/a_215_7# 3.99e-20
C10931 _326_/a_193_7# _326_/a_543_7# -0.0231f
C10932 _162_/X _313_/a_193_7# 1.64e-20
C10933 _255_/B _324_/D 1.61e-20
C10934 _328_/a_761_249# _320_/Q 0.00338f
C10935 _328_/a_193_7# _329_/Q 0.0325f
C10936 _339_/Q _198_/a_250_257# 6.25e-20
C10937 _318_/Q _331_/a_1108_7# 2.2e-20
C10938 _341_/Q _243_/a_199_7# 1.03e-19
C10939 repeater43/X _333_/a_448_7# -2.34e-19
C10940 _329_/a_193_7# VGND 0.0109f
C10941 _329_/a_543_7# VPWR 0.00183f
C10942 _328_/Q VGND 2.92f
C10943 _144_/a_27_7# _217_/A 0.00107f
C10944 _308_/a_218_334# _306_/S 7.74e-19
C10945 _296_/a_295_257# VGND -9.38e-19
C10946 _296_/a_109_7# VPWR -0.00106f
C10947 _259_/a_113_257# _338_/Q 8.99e-19
C10948 _308_/X cal 8.32e-19
C10949 _258_/a_505_n19# _260_/A 7.65e-21
C10950 _251_/X _314_/D 0.0454f
C10951 _341_/a_27_7# _248_/A 0.013f
C10952 _329_/a_1108_7# _297_/B 0.00159f
C10953 _342_/a_27_7# cal 2.72e-19
C10954 _275_/A _286_/B 8.1e-20
C10955 _346_/SET_B _312_/Q 0.394f
C10956 _308_/S _228_/A 3.09e-20
C10957 _281_/Y _328_/D 0.00191f
C10958 _322_/a_1270_373# result[6] 3.25e-20
C10959 _165_/X clkbuf_2_1_0_clk/a_75_172# 3.19e-19
C10960 output22/a_27_7# result[0] 0.00457f
C10961 _290_/A _309_/a_1108_7# 0.014f
C10962 _333_/a_805_7# _206_/A 4.25e-19
C10963 _332_/a_543_7# _332_/D 4.88e-19
C10964 _301_/a_512_257# _347_/Q 1.79e-19
C10965 _301_/a_149_7# _299_/X 0.0168f
C10966 _329_/a_761_249# repeater42/a_27_7# 3.57e-20
C10967 _321_/Q _283_/A 7.39e-19
C10968 _182_/a_79_n19# _147_/A 5.82e-20
C10969 _188_/a_76_159# _182_/X 1.16e-21
C10970 _328_/a_27_7# _328_/a_761_249# -0.0166f
C10971 _223_/a_93_n19# _327_/Q 1.77e-21
C10972 _153_/a_487_257# _153_/A 0.00166f
C10973 _347_/a_1108_7# _347_/D 1.26e-19
C10974 _303_/A _232_/X 0.00286f
C10975 _274_/a_39_257# _216_/X 1.75e-20
C10976 _308_/X _150_/a_193_257# 2.66e-20
C10977 _164_/Y _345_/Q 0.0138f
C10978 _261_/A _311_/D 0.0155f
C10979 _229_/a_76_159# _229_/a_226_7# -2.84e-32
C10980 _237_/a_199_7# _346_/SET_B 3.05e-20
C10981 _275_/Y _306_/S 0.0488f
C10982 _269_/A VGND 0.727f
C10983 _167_/X _306_/a_76_159# 1.05e-20
C10984 _215_/A _336_/a_193_7# 4.56e-22
C10985 _316_/a_193_7# _248_/A 0.0129f
C10986 _329_/D _328_/D 2.74e-19
C10987 clkbuf_2_1_0_clk/A _199_/a_93_n19# 0.0125f
C10988 _346_/a_27_7# _279_/Y 7e-21
C10989 _270_/a_121_257# VPWR 3.17e-19
C10990 _254_/B _202_/a_93_n19# 0.074f
C10991 _317_/Q _318_/a_27_7# 4.17e-21
C10992 output34/a_27_7# _273_/A 0.0121f
C10993 _324_/a_1108_7# _325_/Q 6.5e-21
C10994 _315_/a_193_7# _315_/a_651_373# -0.00701f
C10995 result[0] _341_/a_805_7# 1.5e-19
C10996 _333_/a_448_7# _191_/B 0.0165f
C10997 _331_/Q _331_/a_761_249# 0.0285f
C10998 _326_/Q _224_/a_256_7# 3.08e-19
C10999 _308_/S _216_/A 0.00261f
C11000 _340_/a_761_249# _190_/A 4.08e-21
C11001 _316_/a_193_7# _331_/CLK 0.00171f
C11002 _316_/a_27_7# _316_/D 0.141f
C11003 _344_/Q _171_/a_292_257# 3.89e-19
C11004 _310_/a_1462_7# _310_/Q 7.11e-19
C11005 _343_/D VGND 0.0607f
C11006 clkbuf_0_clk/X _330_/a_27_7# 8.36e-20
C11007 input3/a_27_7# en 0.0188f
C11008 _311_/a_27_7# _297_/Y 1.88e-21
C11009 _225_/B _153_/A 1.89e-21
C11010 _338_/a_651_373# _340_/CLK 0.0268f
C11011 _294_/A _311_/a_1108_7# 1.13e-20
C11012 input1/X _203_/a_209_257# 0.0443f
C11013 output11/a_27_7# _333_/Q 3.49e-20
C11014 _318_/Q clkbuf_0_clk/X 0.00784f
C11015 _301_/a_51_257# VPWR 0.0505f
C11016 _167_/a_373_7# VGND -0.00114f
C11017 cal _254_/B 0.0668f
C11018 _346_/SET_B _347_/a_448_7# 4.73e-21
C11019 _313_/Q _157_/A 1.01e-24
C11020 clkbuf_1_1_0_clk/a_75_172# VPWR 0.071f
C11021 _326_/a_27_7# _248_/A 1.33e-19
C11022 clkbuf_2_1_0_clk/A _336_/Q 1.48e-20
C11023 _334_/a_27_7# _334_/a_761_249# -0.0166f
C11024 input1/a_75_172# _312_/a_193_7# 2.12e-19
C11025 _200_/a_93_n19# _346_/SET_B 8.63e-20
C11026 _181_/X _222_/a_584_7# 6.34e-19
C11027 _290_/A _311_/a_1462_7# 9.05e-19
C11028 _327_/a_27_7# _331_/CLK 0.0816f
C11029 _325_/Q _324_/D 8.92e-19
C11030 _321_/a_193_7# _321_/Q 0.0247f
C11031 _286_/B _345_/D 1.15e-19
C11032 _197_/a_27_7# _254_/B 0.00905f
C11033 _248_/B _297_/B 0.522f
C11034 _338_/a_761_249# _337_/a_193_7# 3.01e-20
C11035 _338_/a_543_7# _337_/a_27_7# 6.11e-21
C11036 _338_/a_27_7# _337_/a_543_7# 1.06e-19
C11037 repeater43/X _304_/a_257_159# 3.1e-19
C11038 _326_/a_27_7# _331_/CLK 0.0412f
C11039 _196_/A _207_/C 1.07e-20
C11040 _311_/a_193_7# _310_/a_27_7# 3.08e-19
C11041 _286_/B _313_/a_1108_7# 0.0019f
C11042 _196_/A _313_/a_1283_n19# 4.6e-20
C11043 _327_/a_27_7# _273_/A 6.96e-21
C11044 _294_/A _275_/Y 0.00945f
C11045 _283_/Y _195_/a_109_257# 2.05e-20
C11046 _255_/X VGND 0.108f
C11047 repeater43/X _177_/A 0.0131f
C11048 _257_/a_448_7# VGND 0.0186f
C11049 _342_/D _149_/a_27_7# 1.32e-19
C11050 output27/a_27_7# _269_/A 0.00937f
C11051 _160_/A _173_/a_76_159# 7.23e-21
C11052 _325_/a_27_7# _223_/a_93_n19# 2.29e-21
C11053 clkc VGND 0.587f
C11054 _341_/a_639_7# _341_/D 0.00445f
C11055 ctln[5] _340_/CLK 1.53e-19
C11056 _326_/a_27_7# _273_/A 1.56e-20
C11057 _311_/Q _284_/A 5.53e-21
C11058 _161_/Y _344_/Q 0.342f
C11059 _258_/a_439_7# _284_/A 3.69e-19
C11060 _321_/a_193_7# _318_/a_193_7# 5.06e-21
C11061 rstn _269_/Y 0.00739f
C11062 _332_/a_639_7# _333_/Q 0.00103f
C11063 _210_/a_27_7# VPWR 0.00104f
C11064 _340_/a_27_7# _337_/a_1108_7# 0.00102f
C11065 _340_/a_193_7# _337_/a_1283_n19# 0.00185f
C11066 _340_/a_1108_7# _337_/a_27_7# 0.00102f
C11067 _340_/a_1283_n19# _337_/a_193_7# 0.00185f
C11068 _210_/a_109_257# VGND 0.00203f
C11069 _307_/a_439_7# _181_/X 6.73e-20
C11070 _254_/A _286_/B 0.0412f
C11071 _317_/Q _246_/B 0.0362f
C11072 repeater43/X _333_/D 0.0133f
C11073 _338_/a_1270_373# _346_/SET_B -2.06e-19
C11074 _338_/a_1108_7# _338_/Q 5.52e-19
C11075 _216_/X _216_/a_27_7# 0.048f
C11076 _181_/X _304_/S 0.0519f
C11077 _329_/Q _319_/a_543_7# 1.7e-20
C11078 _238_/B _319_/a_193_7# 0.0204f
C11079 _326_/a_27_7# _222_/a_93_n19# 0.01f
C11080 _281_/Y _305_/a_76_159# 1.01e-19
C11081 _310_/a_543_7# VGND 0.0212f
C11082 _310_/a_1108_7# VPWR 0.0179f
C11083 _313_/Q _260_/A 5.23e-20
C11084 input4/X _332_/a_543_7# 2.22e-20
C11085 repeater43/X _332_/a_193_7# 0.0018f
C11086 _344_/a_1602_7# _344_/D 1.32e-20
C11087 _344_/a_956_373# _344_/Q 1.59e-19
C11088 _168_/a_109_7# _161_/Y 1.26e-19
C11089 _319_/Q _322_/a_193_7# 1.13e-20
C11090 output21/a_27_7# _331_/a_1283_n19# 2.03e-20
C11091 _294_/A _309_/a_639_7# 0.00429f
C11092 _340_/Q _311_/D 1.64e-21
C11093 _258_/a_76_159# _306_/S 0.0591f
C11094 _334_/a_27_7# _333_/Q 2.29e-21
C11095 repeater43/X _325_/D 0.13f
C11096 _316_/Q _317_/Q 0.0823f
C11097 clkbuf_2_1_0_clk/A _170_/a_489_373# 0.00219f
C11098 _264_/a_199_7# VGND 4.53e-20
C11099 _298_/B _227_/A 7.97e-19
C11100 _340_/a_805_7# _346_/SET_B 8.73e-20
C11101 _181_/X _225_/X 0.0137f
C11102 _182_/X _147_/A 0.0687f
C11103 _196_/A _150_/C 2.51e-19
C11104 _307_/X _181_/X 2.85e-20
C11105 _343_/CLK _298_/C 9.41e-20
C11106 _332_/a_1108_7# _206_/A 8.74e-19
C11107 _339_/a_543_7# _338_/a_27_7# 5.44e-20
C11108 _339_/a_27_7# _338_/a_543_7# 1.2e-19
C11109 _344_/a_27_7# _167_/X 2.91e-21
C11110 _279_/Y _275_/A 3.09e-20
C11111 _256_/a_209_257# _191_/B 0.00131f
C11112 _309_/a_761_249# _310_/a_543_7# 9.16e-21
C11113 _182_/X _149_/A 4.83e-21
C11114 _259_/a_113_257# _309_/D 0.00649f
C11115 _328_/a_1283_n19# _319_/a_27_7# 5.72e-19
C11116 _198_/a_93_n19# _194_/X 1.28e-21
C11117 _229_/a_556_7# _248_/A -0.0013f
C11118 _306_/X _267_/A 9.44e-21
C11119 _334_/Q _333_/D 2.39e-20
C11120 _286_/B _309_/D 0.0055f
C11121 ctln[6] _211_/a_109_7# 1.42e-19
C11122 _318_/Q _286_/Y 0.00658f
C11123 _243_/a_113_257# VPWR 0.0495f
C11124 _175_/Y VPWR 0.812f
C11125 _342_/a_1283_n19# _228_/A 1.13e-21
C11126 _183_/a_553_257# _162_/X 0.00218f
C11127 _327_/a_1270_373# _346_/SET_B -2.06e-19
C11128 _324_/a_1108_7# _326_/Q 0.00247f
C11129 trim[0] trim[2] 0.0574f
C11130 _346_/a_193_7# _346_/a_1032_373# -0.00364f
C11131 _334_/Q _332_/a_193_7# 1.73e-21
C11132 _334_/D _332_/a_1108_7# 2.34e-20
C11133 repeater43/X _341_/a_1283_n19# -0.0119f
C11134 _164_/A _337_/Q 2.28e-20
C11135 _325_/a_1283_n19# _162_/X 3.98e-21
C11136 _169_/Y _346_/D 6.4e-20
C11137 _176_/a_27_7# _323_/Q 1.82e-19
C11138 _165_/a_78_159# _345_/Q 0.00539f
C11139 _203_/a_209_7# _284_/A 1.56e-19
C11140 _340_/a_1108_7# _339_/a_27_7# 4.01e-21
C11141 _340_/a_543_7# _339_/a_761_249# 1.11e-20
C11142 _340_/a_761_249# _339_/a_543_7# 1.11e-20
C11143 _254_/B _284_/A 0.018f
C11144 _333_/D _191_/B 0.0789f
C11145 _320_/a_1108_7# _328_/Q 3.51e-19
C11146 _242_/A _318_/a_651_373# 0.00299f
C11147 _326_/Q _324_/D 0.00314f
C11148 _344_/a_1032_373# _290_/A 0.0113f
C11149 _277_/A VPWR 0.444f
C11150 _343_/Q _225_/X 0.00609f
C11151 _329_/a_27_7# _214_/a_109_257# 1.38e-20
C11152 _324_/a_193_7# _227_/A 0.0404f
C11153 _346_/SET_B _340_/CLK 0.475f
C11154 _294_/A _258_/a_76_159# 9.36e-21
C11155 _336_/a_543_7# VPWR -0.00108f
C11156 _181_/X _331_/a_543_7# 2.2e-19
C11157 _346_/a_193_7# _273_/A 9.3e-20
C11158 _336_/a_193_7# VGND 0.0252f
C11159 _271_/A _234_/B 0.00951f
C11160 _346_/SET_B _347_/D 5.14e-19
C11161 _326_/a_1217_7# _248_/A 5.49e-20
C11162 _313_/D _216_/A 0.0272f
C11163 _320_/Q _282_/a_121_257# 8.96e-19
C11164 _271_/A _321_/a_1283_n19# 0.0161f
C11165 _321_/a_1462_7# _321_/Q 0.00199f
C11166 _292_/A _288_/Y 1.92e-19
C11167 _207_/X _333_/Q 0.00399f
C11168 _189_/a_27_7# _153_/B 0.00608f
C11169 _275_/Y _254_/Y 1.49e-20
C11170 repeater43/X _316_/a_1108_7# -0.0143f
C11171 _300_/a_27_257# _347_/Q 0.00375f
C11172 _300_/a_301_257# _299_/X 0.00249f
C11173 _321_/a_805_7# VPWR 9.28e-19
C11174 _283_/Y _340_/D 5.23e-20
C11175 _216_/X _327_/Q 0.033f
C11176 rstn _335_/a_1283_n19# 0.0285f
C11177 _161_/Y _306_/S 2.37e-19
C11178 _338_/a_639_7# _343_/CLK 7.64e-20
C11179 repeater43/X _208_/a_78_159# 0.0447f
C11180 _329_/a_761_249# _232_/X 2.61e-21
C11181 _329_/Q _327_/Q 1.13e-19
C11182 _320_/Q _212_/X 0.00539f
C11183 _224_/a_584_7# _217_/A 0.00171f
C11184 _267_/A _147_/Y 0.249f
C11185 _188_/S _251_/X 1.14e-20
C11186 _291_/a_121_257# VPWR 7.02e-19
C11187 _327_/a_193_7# _212_/X 0.00669f
C11188 _327_/a_27_7# _217_/X 0.00423f
C11189 _327_/a_761_249# _327_/Q 0.00119f
C11190 _215_/A _299_/X 7.82e-21
C11191 _319_/a_193_7# _331_/CLK 6.73e-20
C11192 _326_/a_1283_n19# repeater43/X 0.0682f
C11193 clkbuf_2_3_0_clk/a_75_172# VGND 0.0574f
C11194 _275_/Y _310_/a_651_373# 0.00178f
C11195 _277_/Y _299_/X 2.8e-19
C11196 _207_/C _204_/a_27_257# 0.00225f
C11197 _326_/a_193_7# _212_/X 9.66e-19
C11198 _326_/a_27_7# _217_/X 0.0286f
C11199 _281_/A _330_/a_1108_7# 1.69e-20
C11200 _341_/a_1108_7# _226_/X 2.8e-21
C11201 _199_/a_256_7# VGND -1.88e-19
C11202 _199_/a_584_7# VPWR -3.19e-19
C11203 repeater43/X _332_/a_1462_7# 5.26e-19
C11204 _281_/Y _330_/a_761_249# 6.87e-20
C11205 ctlp[5] _328_/Q 9.52e-19
C11206 _343_/D _323_/a_651_373# 9.28e-21
C11207 _185_/A _323_/a_639_7# 0.0016f
C11208 _297_/A _303_/A 0.0518f
C11209 _345_/a_27_7# _345_/a_193_7# -0.0541f
C11210 _313_/Q _340_/Q 0.0439f
C11211 _306_/X _194_/X 6.25e-20
C11212 _279_/Y _254_/A 0.00234f
C11213 _145_/A _316_/a_27_7# 5.45e-20
C11214 _334_/Q _208_/a_78_159# 0.0278f
C11215 _328_/a_193_7# _327_/Q 2.66e-21
C11216 ctlp[7] _331_/a_1108_7# 7.34e-21
C11217 _328_/a_27_7# _212_/X 0.0443f
C11218 _260_/B _157_/a_27_7# 7.71e-19
C11219 _183_/a_471_7# _196_/A 5.41e-20
C11220 _344_/a_27_7# _301_/a_51_257# 5.57e-20
C11221 _302_/a_77_159# _347_/a_1283_n19# 5.34e-19
C11222 _302_/a_227_7# _347_/a_27_7# 2.45e-20
C11223 _341_/Q VPWR 1.18f
C11224 _183_/a_27_7# _181_/X 0.00182f
C11225 _346_/a_956_373# _346_/SET_B 4.41e-19
C11226 clk _181_/X 0.138f
C11227 _325_/a_448_7# _181_/X 0.00179f
C11228 _255_/B _181_/a_27_7# 3.93e-19
C11229 _294_/A _161_/Y 4.12e-20
C11230 _300_/a_27_257# _297_/B 1.34e-19
C11231 _340_/CLK _206_/A 3.09e-19
C11232 _340_/CLK _313_/a_761_249# 9.01e-21
C11233 _240_/B _318_/Q 3.34e-20
C11234 input4/X _334_/a_1108_7# 2.73e-21
C11235 repeater43/X _334_/a_543_7# 0.00392f
C11236 _316_/Q _315_/a_193_7# 1.98e-20
C11237 output23/a_27_7# _315_/a_1108_7# 8.68e-19
C11238 _337_/a_448_7# _340_/CLK 0.0253f
C11239 _252_/a_109_257# _228_/A 1.04e-19
C11240 _200_/a_93_n19# _337_/D 6.44e-19
C11241 _342_/a_193_7# _185_/A 3.15e-19
C11242 _325_/a_27_7# _216_/X 0.00124f
C11243 _321_/Q _242_/B 1.18e-20
C11244 _343_/CLK _332_/D 3.72e-20
C11245 _339_/Q _312_/D 0.0592f
C11246 _257_/a_222_53# _305_/a_76_159# 3.22e-21
C11247 _257_/a_79_159# _305_/a_505_n19# 5.21e-20
C11248 clkbuf_2_2_0_clk/a_75_172# _338_/D 2.34e-19
C11249 _344_/a_1182_221# _297_/Y 0.0745f
C11250 _286_/B _202_/a_250_257# 0.00101f
C11251 input4/X _338_/D 6.48e-20
C11252 _334_/a_1108_7# _207_/C 0.0375f
C11253 _163_/a_292_257# _158_/Y 7.38e-20
C11254 ctlp[0] result[7] 0.0502f
C11255 _242_/a_109_257# VGND -0.00114f
C11256 _156_/a_39_257# _347_/D 1.84e-19
C11257 _258_/a_76_159# _254_/Y 2.39e-20
C11258 _315_/a_639_7# VPWR 8.11e-19
C11259 _315_/a_651_373# VGND 7.25e-19
C11260 _183_/a_553_257# _298_/C 3.5e-19
C11261 _227_/A ctln[0] 7.52e-20
C11262 _342_/Q _308_/X 0.0736f
C11263 _196_/A cal 0.00462f
C11264 _286_/B input1/X 0.422f
C11265 _329_/a_27_7# _331_/D 1.87e-19
C11266 clk _343_/Q 9.73e-19
C11267 _274_/a_39_257# _327_/Q 0.0211f
C11268 trimb[2] _162_/A 4.6e-20
C11269 _320_/a_1283_n19# _319_/D 0.00112f
C11270 _339_/a_193_7# _332_/Q 1.41e-20
C11271 _336_/a_1462_7# VGND -7.21e-19
C11272 _271_/A _224_/a_250_257# 2.19e-20
C11273 _342_/a_27_7# _342_/Q 1.34e-19
C11274 _329_/a_193_7# _330_/a_27_7# 7.02e-19
C11275 _329_/a_27_7# _330_/a_193_7# 7.02e-19
C11276 _326_/a_27_7# _325_/a_761_249# 2.29e-20
C11277 _326_/a_193_7# _325_/a_193_7# 6.35e-20
C11278 _334_/a_651_373# _334_/D 8.49e-19
C11279 _334_/a_543_7# _334_/Q 8.84e-21
C11280 repeater43/X _248_/A 1.78f
C11281 _318_/a_193_7# _242_/B 1.16e-19
C11282 _315_/D _314_/a_805_7# 0.00259f
C11283 _196_/A _197_/a_27_7# 0.00188f
C11284 _329_/a_193_7# _318_/Q 2.32e-20
C11285 output31/a_27_7# _285_/A 0.0277f
C11286 _318_/Q _328_/Q 0.158f
C11287 ctln[1] _334_/a_193_7# 9.1e-20
C11288 _314_/a_1283_n19# VGND 0.0279f
C11289 _314_/a_448_7# VPWR 0.0169f
C11290 _346_/SET_B _319_/a_639_7# 0.00103f
C11291 _324_/a_193_7# _297_/B 0.00401f
C11292 _346_/SET_B _313_/a_543_7# 0.0134f
C11293 _315_/D _217_/A 8.11e-20
C11294 _346_/SET_B _337_/a_651_373# 1.78e-33
C11295 _194_/X _147_/Y 2.25e-19
C11296 _157_/A _347_/a_27_7# 0.00953f
C11297 output24/a_27_7# _244_/B 1.14e-19
C11298 _340_/CLK _147_/A 0.111f
C11299 clk _332_/a_1283_n19# 0.0445f
C11300 repeater43/X _331_/CLK 0.307f
C11301 _347_/Q _160_/X 0.0764f
C11302 _299_/X _300_/Y 0.156f
C11303 _147_/A _347_/D 3.46e-20
C11304 _154_/a_27_7# _205_/a_297_7# 1.65e-20
C11305 _324_/a_1108_7# _324_/D 0.0567f
C11306 _311_/D _310_/a_448_7# 1.64e-19
C11307 _311_/a_448_7# _310_/D 2.91e-20
C11308 _311_/a_761_249# _310_/Q 9.29e-22
C11309 _196_/A _150_/a_193_257# 1.14e-20
C11310 repeater42/a_27_7# _227_/A 4.05e-20
C11311 _170_/a_556_7# VGND 5.23e-19
C11312 repeater43/X _190_/A 0.124f
C11313 ctlp[7] clkbuf_0_clk/X 1.5e-19
C11314 _322_/a_639_7# _269_/A 0.00132f
C11315 _270_/a_39_257# _244_/B 2.82e-19
C11316 _279_/Y _302_/a_227_257# 2.18e-19
C11317 _324_/Q _268_/a_39_257# 0.0361f
C11318 _334_/a_193_7# _192_/B 0.00135f
C11319 _334_/a_543_7# _191_/B 9.73e-19
C11320 cal _298_/X 0.0625f
C11321 _345_/a_27_7# VPWR 0.125f
C11322 _319_/Q _331_/Q 0.127f
C11323 _292_/A _337_/Q 0.0088f
C11324 _308_/S _209_/a_27_257# 5.54e-20
C11325 _339_/a_448_7# _340_/CLK 0.0012f
C11326 _273_/A repeater43/X 0.0122f
C11327 _153_/a_297_257# _153_/B 2.64e-20
C11328 _323_/a_1108_7# _175_/Y 8.5e-19
C11329 _304_/S _346_/SET_B 3e-21
C11330 _340_/a_448_7# _337_/Q 6.16e-21
C11331 _345_/a_652_n19# _297_/B 1.08e-19
C11332 _273_/A _288_/Y 0.214f
C11333 _327_/a_1217_7# _217_/X 1.36e-19
C11334 _162_/X _344_/D 0.00949f
C11335 _232_/X _319_/D 1.07e-19
C11336 _286_/B _286_/Y 0.0138f
C11337 _167_/X _147_/Y 0.0121f
C11338 _339_/a_193_7# _337_/a_193_7# 5.08e-20
C11339 _318_/Q _269_/A 0.215f
C11340 _346_/Q _162_/X 0.37f
C11341 repeater43/X _222_/a_93_n19# 0.00136f
C11342 _145_/A _295_/a_79_n19# 0.00139f
C11343 _277_/A _320_/a_543_7# 0.00193f
C11344 _188_/a_76_159# _304_/S 2.11e-20
C11345 _184_/a_505_n19# _341_/Q 4.83e-20
C11346 _342_/Q _254_/B 5.23e-20
C11347 _342_/Q _317_/D 3.58e-20
C11348 _334_/Q _190_/A 0.029f
C11349 _342_/a_805_7# _269_/A 3.43e-19
C11350 _299_/X VGND 1.13f
C11351 _308_/a_439_7# _227_/A 0.00127f
C11352 _301_/X _347_/a_1108_7# 4.92e-19
C11353 _303_/A _347_/a_761_249# 1.66e-19
C11354 _260_/A _347_/a_27_7# 1.98e-19
C11355 _322_/a_27_7# _322_/D 0.0554f
C11356 clkbuf_2_2_0_clk/a_75_172# _343_/CLK 4.73e-19
C11357 _319_/a_193_7# _217_/X 0.00192f
C11358 _346_/SET_B _267_/B 0.303f
C11359 _160_/X _297_/B 0.0853f
C11360 _339_/a_651_373# _346_/SET_B 2.99e-19
C11361 _283_/Y _153_/a_215_257# 2.32e-21
C11362 trim[2] _312_/a_1270_373# 5.7e-21
C11363 _188_/a_505_n19# _147_/A 1.7e-20
C11364 input4/X _343_/CLK 3.47f
C11365 _188_/a_76_159# _307_/X 0.00778f
C11366 _337_/D _340_/CLK 0.0784f
C11367 _192_/a_68_257# _336_/D 3.81e-21
C11368 _246_/B _304_/X 0.0107f
C11369 _258_/a_505_n19# _336_/a_1283_n19# 2.59e-19
C11370 _308_/X _298_/a_181_7# 4.16e-20
C11371 _192_/B _332_/Q 6.42e-20
C11372 _191_/B _190_/A 0.671f
C11373 _157_/A _216_/X 2.74e-20
C11374 _166_/Y _299_/a_78_159# 9.74e-19
C11375 _324_/Q _316_/a_27_7# 6.1e-20
C11376 _292_/A _339_/Q 0.0107f
C11377 _279_/Y clkbuf_0_clk/X 0.157f
C11378 repeater43/X _145_/a_113_7# 1.08e-19
C11379 _341_/a_1108_7# input1/X 1.93e-19
C11380 _196_/A _284_/A 0.534f
C11381 _330_/Q VPWR 0.782f
C11382 _172_/A _260_/a_27_257# 0.0705f
C11383 _145_/A _180_/a_29_13# 0.0486f
C11384 _293_/a_39_257# _336_/Q 1.02e-19
C11385 clk _208_/a_215_7# 5.09e-20
C11386 _343_/CLK _207_/C 0.27f
C11387 _198_/a_250_257# _336_/a_761_249# 2.94e-21
C11388 _198_/a_93_n19# _336_/a_543_7# 2.69e-20
C11389 _317_/a_543_7# _248_/A 0.00215f
C11390 _316_/Q _304_/X 2.51e-21
C11391 _330_/D clkbuf_2_1_0_clk/A 8.1e-20
C11392 _308_/S _153_/A 3.8e-19
C11393 trimb[0] _285_/Y 0.0394f
C11394 _327_/a_1108_7# clkbuf_0_clk/X 0.0531f
C11395 _269_/Y VPWR 0.0938f
C11396 _321_/Q _318_/a_1283_n19# 2.5e-21
C11397 _254_/A _313_/a_27_7# 0.00144f
C11398 _324_/a_805_7# VPWR 2.23e-19
C11399 _324_/a_1270_373# VGND 9.25e-20
C11400 _236_/B _317_/a_193_7# 5.23e-20
C11401 _317_/a_761_249# _316_/D 7.51e-21
C11402 _317_/a_543_7# _331_/CLK 6.54e-19
C11403 ctlp[6] _330_/Q 2.78e-19
C11404 _315_/D _314_/Q 0.0271f
C11405 _306_/S _263_/B 2.32e-20
C11406 _143_/a_181_7# _149_/A 0.00108f
C11407 _314_/D VPWR 0.0946f
C11408 _318_/a_761_249# VPWR 0.0111f
C11409 _318_/a_27_7# VGND 0.0242f
C11410 _343_/a_639_7# VPWR 6.69e-19
C11411 _343_/a_651_373# VGND 9.92e-19
C11412 _218_/a_93_n19# _218_/a_256_7# -3.48e-20
C11413 _272_/a_39_257# _246_/B 0.0104f
C11414 _157_/A _347_/a_1217_7# 3.15e-20
C11415 _281_/Y _181_/X 1.55e-19
C11416 _254_/B _204_/Y 2.22e-20
C11417 _279_/Y input1/X 0.00815f
C11418 _328_/a_1283_n19# clkbuf_0_clk/X 1.29e-20
C11419 _345_/a_652_n19# _275_/Y 4.46e-20
C11420 _311_/D _310_/D 7.12e-19
C11421 _236_/B _331_/a_1283_n19# 1.31e-19
C11422 _316_/D _331_/a_1108_7# 3.7e-21
C11423 _331_/CLK _331_/a_448_7# 0.00108f
C11424 _318_/a_193_7# _318_/a_1283_n19# -5.37e-19
C11425 _273_/A _172_/a_109_257# 0.00231f
C11426 _254_/a_109_257# _254_/A 0.00285f
C11427 cal _204_/a_27_257# 5.42e-20
C11428 _225_/X _206_/A 0.0163f
C11429 _233_/a_113_257# _232_/A 5.94e-21
C11430 _313_/a_543_7# _147_/A 0.0469f
C11431 _341_/a_1108_7# _286_/Y 0.0548f
C11432 _345_/a_586_7# VPWR 0.00166f
C11433 _345_/a_956_373# VGND 1.14e-19
C11434 _319_/Q output14/a_27_7# 6.37e-23
C11435 _339_/D _340_/CLK 0.0427f
C11436 _254_/B _298_/a_181_7# 1.85e-19
C11437 _154_/a_27_7# _298_/A 3.3e-20
C11438 _154_/A _153_/B 0.148f
C11439 _301_/a_51_257# _147_/Y 0.00355f
C11440 _307_/a_505_n19# _191_/B 0.0535f
C11441 _244_/a_109_257# _298_/A 1.32e-19
C11442 _336_/a_27_7# _254_/B 0.00194f
C11443 _283_/A _330_/a_651_373# 3.94e-19
C11444 _343_/CLK _150_/C 1.82e-20
C11445 clk _334_/a_448_7# 0.00212f
C11446 _284_/A _347_/a_1283_n19# 2.64e-21
C11447 _311_/a_27_7# _311_/a_761_249# -6.54e-19
C11448 _307_/a_439_7# _147_/A 0.0017f
C11449 _316_/a_27_7# _228_/A 8.18e-22
C11450 _283_/A _333_/a_543_7# 0.0359f
C11451 repeater43/X _217_/X 0.0196f
C11452 _178_/a_27_7# _191_/B 0.0018f
C11453 _188_/a_535_334# _145_/A 7.27e-19
C11454 clkbuf_2_3_0_clk/A _172_/Y 1.01e-19
C11455 clkbuf_2_1_0_clk/a_75_172# VPWR 0.101f
C11456 _304_/S _147_/A 6.19e-20
C11457 result[3] _242_/A 0.00375f
C11458 _275_/Y _160_/X 0.0157f
C11459 _255_/B _182_/a_79_n19# 2.05e-20
C11460 _260_/B _267_/A 0.0113f
C11461 _294_/A _263_/B 1.46e-19
C11462 _265_/a_109_257# _162_/A 0.00122f
C11463 _181_/a_27_7# _314_/a_193_7# 2.37e-19
C11464 _273_/A _337_/Q 4.78e-19
C11465 _218_/a_584_7# VGND -2.45e-19
C11466 _246_/B VGND 0.161f
C11467 output27/a_27_7# _318_/a_27_7# 1.63e-19
C11468 _239_/a_113_257# _329_/Q 2.58e-20
C11469 _279_/Y _286_/Y 0.03f
C11470 _304_/S _149_/A 0.00193f
C11471 _309_/a_1108_7# _309_/Q 0.00154f
C11472 result[6] _331_/CLK 0.0121f
C11473 _308_/a_535_334# VPWR -1.35e-19
C11474 _308_/a_505_n19# VGND 0.0788f
C11475 _279_/Y _219_/a_584_7# 4.69e-20
C11476 _343_/a_193_7# _323_/a_761_249# 4.61e-21
C11477 _343_/a_27_7# _323_/a_543_7# 6.81e-21
C11478 _343_/a_543_7# _323_/a_27_7# 4.97e-20
C11479 _343_/a_761_249# _323_/a_193_7# 4.99e-21
C11480 output32/a_27_7# clkc 1.6e-21
C11481 _290_/A _312_/Q 0.564f
C11482 _147_/A _225_/X 0.0105f
C11483 _311_/a_448_7# VPWR 0.00229f
C11484 _324_/Q _295_/a_79_n19# 3.74e-21
C11485 _307_/X _147_/A 0.0484f
C11486 _311_/a_1283_n19# VGND 0.0113f
C11487 cal _334_/a_1108_7# 5.52e-19
C11488 _306_/X _336_/a_543_7# 1.47e-20
C11489 _313_/Q _336_/a_1283_n19# 0.00149f
C11490 _313_/D _336_/a_651_373# 2.47e-19
C11491 _283_/Y clkbuf_2_1_0_clk/A 0.0129f
C11492 _316_/Q VGND 1.33f
C11493 result[1] VPWR 0.159f
C11494 _172_/A _227_/A 0.664f
C11495 output22/a_27_7# _228_/A 3.93e-19
C11496 _342_/a_1108_7# _298_/A 1.8e-21
C11497 repeater43/X _296_/Y 1.33e-20
C11498 _307_/X _149_/A 3.41e-20
C11499 result[3] _322_/D 4.6e-20
C11500 _271_/Y VGND 1.45f
C11501 _337_/a_543_7# _337_/Q 0.00294f
C11502 _345_/a_27_7# _344_/a_27_7# 0.00167f
C11503 _216_/X _221_/a_250_257# 0.0051f
C11504 _335_/a_761_249# VGND 0.00158f
C11505 _227_/A _335_/D 0.118f
C11506 _335_/a_1283_n19# VPWR 0.00256f
C11507 _197_/X _336_/a_651_373# 3.66e-19
C11508 comp trimb[4] 0.0899f
C11509 cal _338_/D 0.18f
C11510 input1/a_75_172# _338_/Q 0.0183f
C11511 _184_/a_76_159# VPWR 0.00973f
C11512 _232_/A _223_/a_93_n19# 4.49e-19
C11513 _306_/S _194_/A 0.149f
C11514 _336_/Q _203_/a_303_7# 3.48e-19
C11515 _301_/X _346_/SET_B 0.00907f
C11516 _254_/A _313_/a_1217_7# 1.01e-19
C11517 _225_/B _254_/B 0.332f
C11518 _338_/a_761_249# _340_/Q 3.91e-19
C11519 _338_/a_193_7# _306_/S 0.00477f
C11520 _338_/a_27_7# _193_/Y 0.0141f
C11521 _338_/a_543_7# _194_/X 0.00964f
C11522 _322_/Q _242_/A 1.3e-19
C11523 _333_/a_193_7# _153_/a_109_53# 2.38e-19
C11524 _325_/a_761_249# repeater43/X -0.0024f
C11525 _209_/X _333_/a_27_7# 0.00124f
C11526 _273_/A _339_/Q 4.04e-20
C11527 _318_/a_1217_7# VGND -4.7e-19
C11528 _324_/Q _180_/a_29_13# 0.00661f
C11529 _258_/S _306_/S 0.134f
C11530 _346_/SET_B _174_/a_373_7# 2.37e-19
C11531 _218_/a_93_n19# _330_/D 0.0015f
C11532 _303_/A _248_/A 0.00857f
C11533 _325_/a_27_7# _327_/Q 4.6e-20
C11534 _275_/Y _309_/a_193_7# 0.0159f
C11535 _344_/a_193_7# _347_/Q 1.65e-20
C11536 ctln[4] _283_/Y 0.1f
C11537 _320_/a_27_7# _220_/a_93_n19# 1.38e-21
C11538 clk _206_/A 0.259f
C11539 result[7] _282_/a_121_257# 1.17e-19
C11540 repeater43/X _317_/a_651_373# 1.83e-20
C11541 _251_/X _347_/a_27_7# 6.7e-22
C11542 _309_/a_805_7# VPWR 0.00146f
C11543 _309_/a_1270_373# VGND 6.76e-20
C11544 _340_/a_761_249# _193_/Y 0.00906f
C11545 _340_/a_543_7# _306_/S 0.0117f
C11546 _340_/a_27_7# _340_/D 0.0442f
C11547 _340_/a_1108_7# _194_/X 0.0203f
C11548 _340_/a_1283_n19# _340_/Q 0.0717f
C11549 ctln[1] _192_/B 1.3e-20
C11550 _227_/A _203_/a_80_n19# 1.71e-19
C11551 _315_/a_448_7# _317_/D 0.00791f
C11552 output11/a_27_7# _306_/S 1.03e-19
C11553 _336_/a_543_7# _147_/Y 0.0357f
C11554 _296_/Y _191_/B 0.074f
C11555 _255_/X _192_/a_150_257# 6.99e-19
C11556 _279_/Y ctln[6] 0.0204f
C11557 _228_/A _295_/a_79_n19# 9.04e-22
C11558 _219_/a_256_7# _346_/SET_B 7.48e-19
C11559 _172_/A _347_/Q 3.03e-19
C11560 _164_/A _310_/a_1283_n19# 1.08e-21
C11561 _273_/A _303_/A 1.05e-19
C11562 clk _334_/D 0.143f
C11563 _333_/a_193_7# _209_/a_27_257# 8.8e-19
C11564 _322_/D _322_/Q 1.11e-19
C11565 _220_/a_584_7# _328_/D 4.33e-19
C11566 output7/a_27_7# clk 0.053f
C11567 _339_/a_543_7# _337_/Q 3.1e-21
C11568 _339_/Q _337_/a_543_7# 0.0358f
C11569 repeater43/X _331_/a_805_7# 6.41e-19
C11570 _322_/a_543_7# _318_/D 9.4e-20
C11571 _270_/a_39_257# _177_/A 1.78e-20
C11572 _145_/A _226_/X 1.96e-20
C11573 _146_/a_29_271# _191_/B 4.61e-20
C11574 _183_/a_1241_257# _304_/S 0.0198f
C11575 result[5] VGND 0.0903f
C11576 output15/a_27_7# _283_/A 6.82e-20
C11577 _255_/X _286_/B 0.561f
C11578 _342_/Q _196_/A 0.936f
C11579 _331_/a_448_7# _217_/X 2.05e-21
C11580 _325_/a_1108_7# _304_/S 7.42e-21
C11581 _320_/a_761_249# VPWR 0.00829f
C11582 _320_/a_27_7# VGND 0.0285f
C11583 _257_/a_544_257# _196_/A 0.00396f
C11584 _257_/a_448_7# _286_/B 6.27e-20
C11585 _323_/a_761_249# VGND 0.00165f
C11586 _323_/a_1283_n19# VPWR 0.0319f
C11587 _294_/A _258_/S 0.496f
C11588 _146_/a_184_13# _150_/C 2.02e-19
C11589 clk _191_/a_109_257# 1.26e-19
C11590 clkbuf_0_clk/a_110_7# _191_/B 0.00251f
C11591 _318_/Q _242_/a_109_257# 3.52e-19
C11592 _320_/a_1283_n19# _297_/B 0.0473f
C11593 _185_/A _343_/Q 0.0125f
C11594 _286_/B _210_/a_109_257# 3.12e-20
C11595 _207_/X _207_/a_27_7# 0.00196f
C11596 trim[2] trim[3] 0.0609f
C11597 _344_/a_193_7# _297_/B 0.00537f
C11598 _256_/a_209_7# _255_/X 6.79e-19
C11599 clk _147_/A 0.00685f
C11600 _258_/a_505_n19# VPWR 0.0489f
C11601 _311_/D VPWR 0.371f
C11602 cal _343_/CLK 0.0534f
C11603 _180_/a_29_13# _228_/A 7.51e-20
C11604 _186_/a_297_7# VGND 0.0401f
C11605 result[4] _331_/CLK 0.233f
C11606 _321_/Q _232_/X 0.0892f
C11607 clk _149_/A 2.84e-19
C11608 _312_/Q _310_/a_27_7# 2.51e-19
C11609 _285_/Y VPWR 0.624f
C11610 _329_/a_1283_n19# _216_/X 0.0027f
C11611 _216_/X _251_/X 0.0758f
C11612 _345_/a_1032_373# _344_/a_1602_7# 5.51e-20
C11613 _345_/a_1602_7# _344_/a_1032_373# 7.78e-20
C11614 _172_/A _297_/B 0.933f
C11615 _277_/Y _172_/B 7.95e-21
C11616 _283_/A _194_/A 4.46e-19
C11617 _328_/a_1283_n19# _240_/B 2.42e-20
C11618 _328_/a_651_373# _319_/Q 8.53e-19
C11619 _222_/a_250_257# _286_/Y 1.06e-19
C11620 _279_/Y _328_/Q 0.0018f
C11621 _188_/S VPWR 0.396f
C11622 _343_/a_27_7# _342_/a_448_7# 7.07e-21
C11623 _343_/a_193_7# _342_/a_1108_7# 2.41e-19
C11624 _343_/a_543_7# _342_/a_543_7# 9.97e-20
C11625 _343_/a_761_249# _342_/a_1283_n19# 2.8e-21
C11626 _338_/a_193_7# _283_/A 6.09e-21
C11627 output27/a_27_7# result[5] 0.00252f
C11628 _329_/a_1283_n19# _329_/Q 0.00292f
C11629 _339_/a_543_7# _339_/Q 2.77e-19
C11630 _160_/X _161_/Y 0.0539f
C11631 _328_/a_448_7# _329_/D 4.59e-20
C11632 _232_/X _297_/B 0.00574f
C11633 _320_/a_1270_373# _279_/A 7.08e-21
C11634 _288_/A _265_/B 0.0141f
C11635 _331_/Q _326_/Q 1.07e-20
C11636 _327_/a_193_7# _327_/D 0.0512f
C11637 _329_/a_1108_7# _327_/a_193_7# 9.3e-21
C11638 _327_/a_1108_7# _328_/Q 8.57e-21
C11639 _329_/a_1283_n19# _327_/a_761_249# 9.61e-21
C11640 _171_/a_493_257# VPWR 5.34e-21
C11641 _171_/a_78_159# VGND -0.0119f
C11642 _313_/a_27_7# _297_/a_27_257# 2.69e-20
C11643 _333_/a_193_7# _153_/A 3.05e-19
C11644 _162_/X _265_/B 6.22e-20
C11645 _212_/a_27_7# VPWR 0.0315f
C11646 _210_/a_307_257# _333_/D 6.15e-19
C11647 _287_/a_39_257# _265_/B 1.22e-19
C11648 _281_/Y _346_/SET_B 0.0276f
C11649 _297_/Y _347_/a_1108_7# 1.35e-19
C11650 _181_/X _242_/A 0.00909f
C11651 _216_/A _180_/a_29_13# 1.43e-19
C11652 _301_/X _147_/A 0.112f
C11653 _325_/a_805_7# _212_/X 1.33e-19
C11654 _340_/a_543_7# _283_/A 1.37e-20
C11655 _290_/A _340_/CLK 1.71e-20
C11656 trim[0] _311_/a_543_7# 1.04e-20
C11657 _285_/A _311_/a_1108_7# 4.94e-19
C11658 cal _339_/a_1108_7# 2.66e-21
C11659 input1/X _339_/a_1283_n19# 4.24e-21
C11660 _166_/Y _346_/SET_B 0.0307f
C11661 output13/a_27_7# _271_/Y 1.61e-20
C11662 _329_/a_1108_7# _328_/a_27_7# 1.1e-19
C11663 _329_/a_1283_n19# _328_/a_193_7# 4.84e-20
C11664 _328_/a_1283_n19# _328_/Q 0.0528f
C11665 _182_/X _298_/a_27_7# 2.38e-19
C11666 _330_/D _328_/D 3.15e-20
C11667 _307_/X _150_/a_27_7# 3.03e-20
C11668 _320_/Q _283_/A 0.173f
C11669 _317_/Q _316_/a_193_7# 6.11e-20
C11670 output24/a_27_7# _316_/a_1108_7# 2.41e-19
C11671 _196_/A _336_/a_27_7# 0.0132f
C11672 _286_/B _336_/a_193_7# 0.0143f
C11673 _315_/D _317_/D 0.00828f
C11674 _345_/a_476_7# _172_/B 0.00577f
C11675 _154_/a_27_7# VGND 0.0355f
C11676 _244_/a_109_257# VGND -8.91e-19
C11677 _185_/A _229_/a_76_159# 0.0159f
C11678 _322_/a_1270_373# _321_/Q 1.93e-19
C11679 ctln[7] VGND 0.076f
C11680 _329_/D _346_/SET_B 0.381f
C11681 _254_/Y _194_/A 8.18e-20
C11682 _285_/A _275_/Y 4.09e-20
C11683 _308_/a_76_159# _308_/X 0.00227f
C11684 _342_/D _298_/B 9.02e-21
C11685 _326_/a_193_7# _283_/A 0.00984f
C11686 clkbuf_2_3_0_clk/A _260_/A 0.0112f
C11687 _306_/S _201_/a_27_7# 4.43e-21
C11688 _311_/a_543_7# _311_/Q 1.77e-19
C11689 _176_/a_27_7# _175_/Y 0.00104f
C11690 _179_/a_27_7# VGND 0.0979f
C11691 _318_/a_193_7# _244_/B 6.43e-20
C11692 _145_/A clkbuf_0_clk/X 1.47e-19
C11693 _322_/a_1283_n19# VGND 0.0219f
C11694 _322_/a_448_7# VPWR -0.0035f
C11695 _313_/a_193_7# _284_/A 0.0111f
C11696 _315_/a_193_7# _177_/a_27_7# 3.2e-21
C11697 _177_/a_27_7# _298_/A 0.00495f
C11698 _346_/a_1182_221# _167_/X 0.00809f
C11699 _344_/a_193_7# _275_/Y 0.0103f
C11700 _258_/S _254_/Y 3.03e-19
C11701 _319_/Q _321_/D 0.0114f
C11702 _320_/a_1217_7# VGND 1.19e-19
C11703 input4/X _195_/a_109_257# 8.42e-19
C11704 _298_/a_181_7# _298_/X 4.5e-19
C11705 _157_/A _192_/B 9.79e-21
C11706 _162_/X _314_/a_27_7# 6.06e-20
C11707 result[0] _269_/A 0.0582f
C11708 output12/a_27_7# repeater43/X 1.54e-21
C11709 _305_/a_218_7# VGND 6.45e-20
C11710 _344_/a_1140_373# VPWR 1.26e-20
C11711 _182_/a_79_n19# _154_/A 8.2e-19
C11712 _231_/a_676_257# _217_/A 5.81e-20
C11713 _320_/D _297_/B 0.0295f
C11714 _309_/a_193_7# _161_/Y 1.44e-20
C11715 clkbuf_2_3_0_clk/A _261_/A 3.41e-20
C11716 _332_/a_1283_n19# _335_/Q 9.95e-20
C11717 _332_/a_543_7# _204_/Y 3.4e-21
C11718 _306_/S _173_/a_226_7# 0.0019f
C11719 _342_/a_193_7# _271_/A 1.33e-21
C11720 _162_/X _170_/a_76_159# 0.0404f
C11721 _279_/Y _255_/X 0.0598f
C11722 _275_/Y _172_/A 0.292f
C11723 _291_/a_39_257# _312_/D 1.04e-19
C11724 _227_/A _333_/a_448_7# 1.01e-20
C11725 _313_/Q VPWR 0.308f
C11726 _279_/Y _257_/a_448_7# 0.00353f
C11727 _344_/D _345_/Q 6.44e-20
C11728 _320_/Q _321_/a_193_7# 1.1e-19
C11729 _144_/A _286_/Y 6.44e-20
C11730 _255_/a_30_13# _190_/A 4.36e-21
C11731 _297_/A _227_/A 2.75e-20
C11732 _337_/a_27_7# _306_/S 5.37e-21
C11733 _337_/a_193_7# _340_/Q 6.73e-19
C11734 _337_/a_761_249# _194_/X 0.00741f
C11735 _318_/Q _318_/a_27_7# 0.0475f
C11736 _281_/Y _206_/A 0.00552f
C11737 _145_/A input1/X 1.95e-20
C11738 _342_/a_1108_7# VGND -0.00591f
C11739 _342_/a_651_373# VPWR 7.31e-19
C11740 _292_/A _310_/a_1283_n19# 0.0177f
C11741 repeater43/X _207_/a_109_7# 2.32e-19
C11742 _335_/a_543_7# _335_/D 0.0103f
C11743 _312_/Q _310_/a_1217_7# 7.83e-20
C11744 _184_/a_505_n19# _188_/S 0.0236f
C11745 _239_/a_113_257# _327_/Q 5.62e-20
C11746 _346_/Q _345_/Q 0.0155f
C11747 _199_/a_346_7# _312_/D 1.04e-19
C11748 clkbuf_2_1_0_clk/A _162_/X 0.528f
C11749 _297_/A _314_/a_1108_7# 5.77e-19
C11750 _324_/Q _317_/a_761_249# 1e-19
C11751 _288_/A _310_/Q 0.0233f
C11752 _275_/A _290_/Y 0.00241f
C11753 _329_/a_761_249# _331_/CLK 1.96e-19
C11754 _268_/a_39_257# _315_/a_761_249# 0.00174f
C11755 _252_/a_27_7# _304_/X 2.49e-20
C11756 _343_/a_27_7# _342_/D 4.38e-19
C11757 _165_/X _173_/a_489_373# 7.92e-20
C11758 _169_/Y _196_/A 0.149f
C11759 _189_/a_27_7# _340_/CLK 1.83e-20
C11760 _319_/Q _319_/a_639_7# 7.11e-19
C11761 _240_/B _319_/a_448_7# 7.02e-21
C11762 _181_/X _336_/Q 2.76e-20
C11763 _196_/A _225_/B 0.126f
C11764 _287_/a_39_257# _310_/Q 0.034f
C11765 _209_/X _298_/C 1.4e-19
C11766 _260_/A _192_/B 0.00458f
C11767 _238_/B _319_/D 0.26f
C11768 _333_/a_1462_7# _153_/A 4.34e-19
C11769 _257_/a_79_159# _340_/CLK 0.0136f
C11770 _172_/B VGND 0.461f
C11771 _312_/a_27_7# _311_/a_27_7# 9.35e-20
C11772 _330_/Q _233_/a_199_7# 1.09e-21
C11773 _235_/a_199_7# _331_/Q 3.01e-20
C11774 _157_/A _302_/a_227_7# 0.00918f
C11775 _341_/a_193_7# _315_/a_27_7# 2.08e-20
C11776 _341_/a_27_7# _315_/a_193_7# 8.6e-21
C11777 output12/a_27_7# _191_/B 4.11e-20
C11778 _273_/A input2/a_27_7# 4.62e-20
C11779 _341_/a_27_7# _298_/A 0.00324f
C11780 clkbuf_2_1_0_clk/A _299_/a_493_257# 2.16e-19
C11781 output18/a_27_7# VPWR 0.0883f
C11782 output24/a_27_7# _248_/A 3.73e-20
C11783 _246_/B _330_/a_27_7# -4.86e-37
C11784 _212_/X _221_/a_93_n19# 0.0317f
C11785 _222_/a_250_257# _328_/Q 1.4e-19
C11786 _327_/Q _221_/a_250_257# 0.00596f
C11787 _233_/a_113_257# VPWR 0.0539f
C11788 _254_/A _168_/a_397_257# 0.00102f
C11789 _145_/A _286_/Y 0.352f
C11790 _281_/Y _147_/A 0.0103f
C11791 _318_/Q _246_/B 0.00565f
C11792 _216_/A _313_/a_1108_7# 0.0524f
C11793 _269_/A _316_/D 1.49e-20
C11794 ctln[7] _335_/a_651_373# 0.0264f
C11795 _340_/CLK _310_/a_27_7# 0.0373f
C11796 _263_/B _262_/a_113_257# 0.00506f
C11797 _258_/S _336_/a_1108_7# 4.2e-19
C11798 output24/a_27_7# _331_/CLK 0.0021f
C11799 _309_/a_761_249# _172_/B 8.79e-21
C11800 _283_/A _207_/X 1.44e-20
C11801 _286_/B _336_/a_1462_7# 1.12e-19
C11802 _339_/a_27_7# _306_/S 0.0122f
C11803 _298_/C _209_/a_109_257# 5.55e-20
C11804 _339_/a_193_7# _340_/Q 0.0119f
C11805 _283_/A _201_/a_27_7# 6.57e-21
C11806 _312_/a_761_249# VGND 0.015f
C11807 _312_/a_1283_n19# VPWR 0.0219f
C11808 _297_/A _347_/Q 0.0116f
C11809 _341_/D _342_/Q 0.00805f
C11810 rstn _334_/a_193_7# 1.55e-20
C11811 _166_/Y _147_/A 1.76e-20
C11812 _308_/S _308_/X 0.00163f
C11813 _313_/Q _306_/a_76_159# 0.00257f
C11814 _270_/a_39_257# _331_/CLK 0.00112f
C11815 _196_/A _314_/a_543_7# 2.09e-19
C11816 _251_/X _216_/a_27_7# 1.32e-20
C11817 _335_/Q _204_/a_27_7# 0.00231f
C11818 _204_/Y _204_/a_27_257# 0.00679f
C11819 _208_/a_215_7# _335_/Q 0.0069f
C11820 _208_/a_493_257# _204_/Y 7.08e-19
C11821 input1/a_75_172# input1/X 0.00232f
C11822 _326_/a_1462_7# _283_/A 1.66e-19
C11823 _316_/Q _318_/Q 2.43e-20
C11824 _304_/a_257_159# _227_/A 0.0202f
C11825 _254_/A _216_/A 0.00914f
C11826 _340_/a_193_7# _336_/a_651_373# 1.1e-21
C11827 _316_/a_193_7# _315_/a_193_7# 4.52e-19
C11828 _316_/a_27_7# _315_/a_761_249# 3.93e-20
C11829 repeater43/a_27_7# _269_/A 0.00169f
C11830 _346_/a_1182_221# clkbuf_1_1_0_clk/a_75_172# 2.38e-19
C11831 _231_/a_306_7# VGND 1.35e-19
C11832 _231_/a_512_7# VPWR -5.3e-19
C11833 clkbuf_2_3_0_clk/A _340_/Q 1.26e-20
C11834 _346_/SET_B _297_/Y 0.188f
C11835 _324_/a_1283_n19# _162_/X 1.18e-21
C11836 _325_/a_543_7# _286_/Y 0.0017f
C11837 _294_/Y _338_/Q 7.28e-19
C11838 _279_/Y _336_/a_193_7# 7.4e-21
C11839 _313_/a_1462_7# _284_/A 1.49e-19
C11840 _330_/Q _330_/a_639_7# 4.51e-19
C11841 _169_/Y _347_/a_1283_n19# 7.15e-21
C11842 trimb[0] _162_/A 0.00109f
C11843 _326_/a_651_373# _242_/A 1e-18
C11844 input4/X _340_/D 2.92e-19
C11845 _180_/a_183_257# _283_/A 4.36e-19
C11846 _186_/a_382_257# _308_/X 5.99e-19
C11847 _289_/a_121_257# VGND -4.24e-19
C11848 _281_/A _331_/a_1108_7# 8.39e-21
C11849 _188_/a_505_n19# _255_/B 0.002f
C11850 _342_/a_193_7# _186_/a_79_n19# 9.87e-21
C11851 _258_/a_76_159# _198_/a_250_257# 1.08e-20
C11852 _330_/a_1270_373# VPWR -2.48e-19
C11853 _330_/a_448_7# VGND 0.00311f
C11854 _182_/X _154_/A 2.4e-20
C11855 _329_/a_805_7# _346_/SET_B -0.00125f
C11856 ctlp[4] _279_/A 2.27e-19
C11857 _251_/a_215_7# _191_/B 3.54e-21
C11858 _343_/a_193_7# _177_/a_27_7# 2.23e-19
C11859 _345_/a_1032_373# _288_/A 1.5e-20
C11860 clkbuf_0_clk/X _324_/Q 8.71e-20
C11861 repeater43/a_27_7# _343_/D 4.57e-21
C11862 _337_/a_27_7# _283_/A 1.93e-19
C11863 _291_/a_39_257# _292_/A 0.0182f
C11864 clk _250_/a_78_159# 0.0128f
C11865 _346_/SET_B _310_/a_193_7# 0.0119f
C11866 _307_/X _250_/X 0.00225f
C11867 _333_/a_761_249# VGND 0.011f
C11868 _333_/a_1283_n19# VPWR 0.0199f
C11869 _227_/A _333_/D 8.54e-20
C11870 _275_/A _240_/a_109_257# 0.00378f
C11871 _193_/Y _313_/a_448_7# 1.54e-21
C11872 _345_/a_1032_373# _162_/X 2.94e-19
C11873 output13/a_27_7# ctln[7] 0.00647f
C11874 _165_/X clkbuf_2_3_0_clk/A 0.43f
C11875 _302_/a_227_257# _228_/A 2.95e-20
C11876 _341_/a_543_7# _341_/Q 1.31e-20
C11877 _252_/a_27_7# VGND 0.0307f
C11878 _337_/a_1462_7# _340_/Q 1.92e-19
C11879 _218_/a_250_257# _331_/Q 3.12e-19
C11880 _346_/Q _302_/a_77_159# 3.45e-20
C11881 _216_/A _309_/D 1.05e-19
C11882 output12/a_27_7# _337_/Q 2.41e-20
C11883 _290_/A _267_/B 0.297f
C11884 cal output30/a_27_7# 0.00142f
C11885 _194_/a_27_7# _194_/A 0.0432f
C11886 _254_/Y _201_/a_27_7# 1.42e-20
C11887 rstn _332_/Q 0.391f
C11888 _285_/A _161_/Y 3.66e-19
C11889 _297_/A _297_/B 0.141f
C11890 _185_/A _206_/A 0.0655f
C11891 _286_/B _299_/X 9.51e-19
C11892 _334_/a_1108_7# _204_/Y 4.07e-20
C11893 _227_/A _325_/D 1.46e-20
C11894 _223_/a_93_n19# VPWR 0.00533f
C11895 _258_/S _284_/a_39_257# 0.0113f
C11896 _162_/A _310_/D 0.0255f
C11897 _314_/a_1283_n19# _347_/a_543_7# 1.08e-19
C11898 _308_/S _254_/B 3.51e-20
C11899 _165_/X _172_/Y 0.00552f
C11900 _306_/S _157_/a_27_7# 1.73e-20
C11901 _258_/S _194_/a_27_7# 9.27e-21
C11902 _331_/CLK _319_/D 0.00935f
C11903 _344_/a_193_7# _161_/Y 0.00119f
C11904 _164_/A _297_/B 1.87e-20
C11905 _242_/A _346_/SET_B 0.242f
C11906 _320_/D _320_/a_193_7# -0.0056f
C11907 _271_/A _322_/Q 0.748f
C11908 _323_/a_543_7# _323_/D 0.00206f
C11909 _157_/A _260_/A 0.00571f
C11910 _329_/a_27_7# _331_/a_193_7# 6.62e-19
C11911 _329_/a_193_7# _331_/a_27_7# 6.62e-19
C11912 _172_/A _161_/Y 0.0532f
C11913 _330_/D _330_/a_761_249# 7.46e-21
C11914 _313_/a_761_249# _297_/Y 3.84e-21
C11915 _329_/a_761_249# _217_/X 1.75e-22
C11916 _329_/a_543_7# _212_/X 9.69e-20
C11917 clkbuf_0_clk/X _281_/A 0.165f
C11918 _339_/a_27_7# _283_/A 0.123f
C11919 _200_/a_250_257# clkbuf_2_1_0_clk/A 0.00749f
C11920 output31/a_27_7# _273_/A 0.0129f
C11921 _342_/Q _343_/CLK 0.00449f
C11922 rstn _337_/a_193_7# 2.36e-21
C11923 trimb[1] trimb[4] 0.0645f
C11924 _196_/A _315_/D 2e-20
C11925 _275_/Y _312_/a_448_7# 0.00882f
C11926 comp _288_/Y 4.18e-20
C11927 _182_/a_510_7# VGND 5.54e-20
C11928 _219_/a_93_n19# _219_/a_346_7# -3.48e-20
C11929 _339_/a_805_7# _193_/Y 4.25e-19
C11930 _258_/S _262_/a_113_257# 0.0102f
C11931 _185_/A _147_/A 0.00215f
C11932 clkbuf_0_clk/X _228_/A 0.0128f
C11933 input4/a_27_7# _343_/CLK 1.49e-19
C11934 _255_/B _304_/S 0.0192f
C11935 _281_/Y _339_/D 1.82e-20
C11936 trimb[4] VGND 0.269f
C11937 trim[1] VGND 0.232f
C11938 _315_/Q _341_/Q 4.97e-21
C11939 _185_/A _149_/A 0.00994f
C11940 _316_/a_27_7# _318_/D 6.1e-23
C11941 _258_/a_439_7# _313_/D 2.24e-19
C11942 _258_/a_505_n19# _306_/X 0.0187f
C11943 _324_/Q _286_/Y 0.0858f
C11944 _324_/a_27_7# _216_/X 0.0126f
C11945 _246_/B _223_/a_346_7# 2.46e-19
C11946 _326_/a_1270_373# _326_/Q 4.42e-20
C11947 _189_/a_27_7# _225_/X 8.4e-19
C11948 _317_/Q repeater43/X 0.0178f
C11949 output35/a_27_7# _265_/B 0.00998f
C11950 _177_/a_27_7# VGND 0.0666f
C11951 _304_/a_257_159# _297_/B 1.35e-21
C11952 _227_/A _208_/a_78_159# 1.27e-19
C11953 VPWR output41/a_27_7# 0.114f
C11954 _255_/B _225_/X 0.029f
C11955 _279_/Y _314_/a_1283_n19# 0.00263f
C11956 _307_/X _255_/B 0.032f
C11957 _257_/a_222_53# _147_/A 3.55e-20
C11958 _342_/a_27_7# _342_/a_1283_n19# -1.57e-19
C11959 _342_/a_193_7# _342_/a_543_7# 3.55e-33
C11960 _313_/Q _198_/a_93_n19# 1.35e-21
C11961 _147_/A _297_/Y 9.1e-19
C11962 _258_/S _266_/a_199_7# 1.7e-19
C11963 _344_/a_652_n19# _172_/B 0.00703f
C11964 _288_/A _309_/a_1283_n19# 2.67e-19
C11965 _250_/a_78_159# _250_/a_292_257# -1.09e-21
C11966 _345_/a_193_7# _162_/A 9.3e-21
C11967 clkbuf_0_clk/X _216_/A 0.00153f
C11968 clk _250_/X 0.206f
C11969 _309_/a_1283_n19# _162_/X 3.26e-21
C11970 _157_/A _251_/a_79_n19# 0.0436f
C11971 _309_/a_1283_n19# _287_/a_39_257# 0.0114f
C11972 _242_/A _319_/a_1270_373# 1.79e-19
C11973 _206_/A _335_/Q 0.186f
C11974 _327_/a_27_7# _304_/X 0.00955f
C11975 _211_/a_373_7# _197_/X 2.4e-19
C11976 _337_/Q _193_/Y 0.0258f
C11977 _343_/a_1108_7# _343_/Q 0.00102f
C11978 _197_/X _198_/a_346_7# 0.00172f
C11979 clkbuf_0_clk/X _221_/a_584_7# 0.00118f
C11980 rstn _339_/a_193_7# 3.22e-20
C11981 _232_/A _327_/Q 0.0113f
C11982 _275_/Y _164_/A 5.14e-20
C11983 _347_/a_27_7# VPWR 0.064f
C11984 _326_/a_27_7# _304_/X 0.0117f
C11985 _145_/A _269_/A 1.2e-21
C11986 _277_/A _319_/a_1283_n19# 0.0212f
C11987 _343_/CLK _204_/Y 0.249f
C11988 _334_/Q _205_/a_297_7# 3.78e-19
C11989 _334_/D _335_/Q 0.00648f
C11990 _346_/SET_B _336_/Q 0.00725f
C11991 _308_/a_505_n19# _286_/B 0.0232f
C11992 repeater43/X _321_/a_761_249# 0.00165f
C11993 _319_/Q _280_/a_68_257# 0.0135f
C11994 output28/a_27_7# _269_/A 0.00203f
C11995 _336_/a_193_7# _313_/a_27_7# 2.01e-20
C11996 _268_/a_121_257# VGND -4.23e-19
C11997 _297_/B _347_/a_761_249# 0.0191f
C11998 _314_/a_193_7# _347_/D 0.00138f
C11999 _314_/D _347_/a_193_7# 2.34e-20
C12000 _267_/A _344_/Q 7.17e-20
C12001 _163_/a_78_159# _310_/D 4.32e-21
C12002 _267_/B _310_/a_27_7# 0.0112f
C12003 _237_/a_199_7# _279_/A 1.21e-19
C12004 input4/X _153_/a_215_257# 2.85e-21
C12005 _216_/A input1/X 1.85e-20
C12006 _313_/D _254_/B 2.12e-19
C12007 _325_/Q _304_/S 1.34e-19
C12008 _312_/Q _311_/a_193_7# 0.00479f
C12009 _279_/Y _299_/X 1.72e-20
C12010 _192_/B _205_/a_79_n19# 0.0215f
C12011 _191_/B _205_/a_297_7# 2.28e-19
C12012 _228_/A _286_/Y 0.00591f
C12013 _322_/Q _232_/a_27_7# 6.8e-19
C12014 _175_/Y _226_/a_297_7# 0.0113f
C12015 _254_/A _301_/a_240_7# 0.0257f
C12016 _341_/a_761_249# VPWR 0.00783f
C12017 _341_/a_27_7# VGND -0.0311f
C12018 _340_/CLK _154_/A 1.85e-22
C12019 _238_/B _347_/Q 2.53e-20
C12020 _318_/Q _322_/a_1283_n19# 5.41e-22
C12021 _305_/X VGND 0.527f
C12022 _242_/A _147_/A 1.07e-20
C12023 _338_/a_27_7# VGND -0.0188f
C12024 _338_/a_761_249# VPWR 0.00144f
C12025 _197_/X _254_/B 0.456f
C12026 _207_/C _153_/a_215_257# 2.19e-19
C12027 _281_/Y _250_/a_78_159# 0.00175f
C12028 _339_/a_1217_7# _283_/A 8.24e-19
C12029 _346_/SET_B _336_/a_805_7# -4.85e-19
C12030 _346_/a_193_7# _277_/Y 3.07e-21
C12031 _209_/X _207_/C 0.0268f
C12032 _319_/D _217_/X 1.04e-19
C12033 _275_/Y _312_/D 0.0986f
C12034 _289_/a_39_257# _311_/Q 0.0168f
C12035 _346_/SET_B _314_/a_761_249# -0.00741f
C12036 _250_/a_215_7# _228_/A 1.74e-19
C12037 output34/a_27_7# VGND 0.0684f
C12038 _339_/Q _193_/Y 0.0866f
C12039 _345_/a_1032_373# _165_/a_215_7# 8.34e-19
C12040 _294_/Y _162_/a_27_7# 0.0111f
C12041 _225_/X _298_/a_27_7# 1.37e-19
C12042 _227_/A _248_/A 2.72e-19
C12043 _317_/Q _317_/a_543_7# 8.44e-19
C12044 ctln[1] rstn 0.0467f
C12045 _162_/A VPWR 0.702f
C12046 _340_/a_1283_n19# VPWR 0.0166f
C12047 _340_/a_761_249# VGND -3.55e-19
C12048 _292_/A _297_/B 1.84e-20
C12049 _346_/SET_B _170_/a_489_373# 2.29e-21
C12050 _193_/Y _202_/a_256_7# 7.99e-20
C12051 _316_/a_1217_7# _318_/D 3.42e-21
C12052 _313_/Q _306_/X 0.034f
C12053 _216_/X VPWR 0.923f
C12054 _216_/A _286_/Y 0.144f
C12055 _248_/A _314_/a_1108_7# 6.54e-20
C12056 _325_/Q _317_/a_27_7# 5.09e-19
C12057 result[7] _283_/A 0.0033f
C12058 _327_/a_543_7# _330_/Q 0.00134f
C12059 _316_/a_543_7# VPWR 0.0295f
C12060 _227_/A _331_/CLK 0.0156f
C12061 _316_/a_193_7# VGND 0.00706f
C12062 _344_/D _284_/A 1.44e-20
C12063 _297_/B _160_/A 1.37e-21
C12064 _271_/A _343_/Q 0.4f
C12065 _258_/S _309_/a_193_7# 0.00171f
C12066 _251_/a_510_7# _286_/Y 0.00141f
C12067 _329_/Q VPWR 0.36f
C12068 _221_/a_584_7# _286_/Y 0.00396f
C12069 _227_/A _190_/A 0.00121f
C12070 _255_/B _183_/a_27_7# 0.00131f
C12071 cal _340_/D 1.3e-20
C12072 _326_/Q _222_/a_584_7# 4.55e-19
C12073 _200_/a_93_n19# _311_/a_193_7# 1.72e-20
C12074 _336_/Q _206_/A 9.76e-19
C12075 _313_/a_193_7# _225_/B 4.9e-20
C12076 _255_/B clk 0.0233f
C12077 _309_/a_1108_7# _312_/Q 6.56e-20
C12078 _342_/D _172_/A 0.0131f
C12079 _327_/a_761_249# VPWR 0.016f
C12080 _327_/a_27_7# VGND -0.00885f
C12081 _317_/a_1283_n19# _248_/B 2.89e-21
C12082 _317_/a_1108_7# _232_/A 0.00102f
C12083 _337_/a_448_7# _336_/Q 2.53e-19
C12084 _271_/A ctlp[1] 0.0123f
C12085 _273_/A _227_/A 0.00494f
C12086 _260_/A _340_/Q 7.68e-20
C12087 _197_/a_27_7# _340_/D 0.00204f
C12088 _346_/a_27_7# _346_/D 0.201f
C12089 _238_/B _297_/B 0.153f
C12090 repeater43/X _315_/a_193_7# 0.0194f
C12091 _277_/Y _173_/a_76_159# 2.97e-19
C12092 _250_/a_215_7# _216_/A 0.00516f
C12093 _250_/a_292_257# _250_/X 6.36e-19
C12094 repeater43/X _298_/A 0.0237f
C12095 _326_/a_27_7# VGND -0.0767f
C12096 _326_/a_761_249# VPWR 0.00899f
C12097 _322_/a_761_249# _322_/Q 2.57e-19
C12098 _327_/a_1283_n19# _297_/B 0.00144f
C12099 _285_/A _263_/B 3.67e-20
C12100 _307_/a_76_159# _341_/Q 1.36e-19
C12101 _234_/B _317_/a_193_7# 1e-19
C12102 _345_/a_193_7# _163_/a_78_159# 0.00765f
C12103 _157_/A _251_/X 0.0226f
C12104 _277_/Y _319_/a_193_7# 5.09e-21
C12105 _346_/a_1140_373# clkbuf_2_1_0_clk/A 2.72e-19
C12106 _324_/Q _296_/a_295_257# 0.00194f
C12107 _332_/a_1270_373# VGND 5.8e-20
C12108 _332_/a_805_7# VPWR 3.03e-19
C12109 _327_/a_193_7# repeater42/a_27_7# 0.00618f
C12110 _331_/Q _214_/a_373_7# 3.71e-19
C12111 _167_/a_27_257# _301_/X 3.07e-20
C12112 _328_/a_193_7# VPWR -0.0896f
C12113 _347_/a_639_7# VGND -0.00129f
C12114 _347_/a_1217_7# VPWR 6.49e-20
C12115 _221_/a_93_n19# _221_/a_256_7# -3.48e-20
C12116 _200_/a_346_7# VGND 5.41e-19
C12117 _326_/a_1217_7# _304_/X 1.19e-20
C12118 _306_/S _267_/A 0.025f
C12119 _308_/S _196_/A 0.0274f
C12120 _165_/X _260_/A 1.4e-19
C12121 _192_/B _225_/a_59_35# 2.46e-19
C12122 _328_/a_543_7# _297_/B 4.37e-20
C12123 _321_/a_193_7# result[7] 3.09e-19
C12124 _258_/S _306_/a_505_n19# 0.021f
C12125 _281_/Y _319_/Q 0.00983f
C12126 _304_/S _326_/Q 0.00325f
C12127 _164_/A _171_/a_292_257# 4.85e-19
C12128 _267_/B _310_/a_1217_7# 2.55e-19
C12129 _347_/Q _248_/A 7.95e-21
C12130 _298_/B _226_/a_79_n19# 7.64e-19
C12131 _341_/Q _226_/a_297_7# 3.68e-21
C12132 _212_/a_27_7# _223_/a_250_257# 1.03e-20
C12133 _324_/a_27_7# _216_/a_27_7# 2.02e-19
C12134 _346_/a_652_n19# _160_/X 2.71e-19
C12135 _343_/CLK _315_/a_448_7# 0.0166f
C12136 _334_/Q _298_/A 0.0016f
C12137 clkbuf_2_3_0_clk/A clkbuf_2_0_0_clk/a_75_172# 5.7e-20
C12138 clkbuf_2_2_0_clk/a_75_172# clkbuf_2_1_0_clk/A 5.7e-20
C12139 _167_/X _344_/Q 0.00257f
C12140 _313_/Q _147_/Y 0.391f
C12141 _334_/a_193_7# VPWR -0.279f
C12142 en _343_/CLK 0.00155f
C12143 _147_/A _336_/Q 4.86e-20
C12144 _292_/A _311_/a_1108_7# 0.00329f
C12145 _333_/a_193_7# _254_/B 1.89e-21
C12146 _344_/a_1182_221# _162_/X 0.00299f
C12147 _190_/a_27_7# VPWR 0.161f
C12148 _186_/a_382_257# _196_/A 6.17e-21
C12149 output26/a_27_7# _269_/A 0.0114f
C12150 _324_/Q _269_/A 0.00358f
C12151 _323_/a_193_7# _298_/X 1.38e-19
C12152 _307_/a_505_n19# _227_/A 0.00208f
C12153 clkbuf_2_3_0_clk/A _310_/D 2.02e-36
C12154 _341_/a_1217_7# VGND -4.69e-19
C12155 _342_/D _244_/B 0.00182f
C12156 _251_/X _260_/A 1.44e-20
C12157 _323_/a_27_7# _343_/Q 5.95e-19
C12158 _273_/A _347_/Q 0.0495f
C12159 _338_/a_1217_7# VGND 1.19e-19
C12160 _319_/Q _329_/D 0.448f
C12161 _191_/B _298_/A 0.00209f
C12162 _281_/Y _250_/X 3.9e-20
C12163 _168_/a_109_7# _167_/X 0.0268f
C12164 _149_/a_27_7# _175_/Y 2.92e-19
C12165 _274_/a_39_257# VPWR 0.0574f
C12166 _330_/a_193_7# _330_/a_1108_7# -0.00656f
C12167 _316_/Q _316_/a_448_7# 0.023f
C12168 _227_/A _178_/a_27_7# 3.69e-20
C12169 _275_/Y _292_/A 0.0341f
C12170 _321_/Q _248_/A 0.0166f
C12171 _329_/a_193_7# _281_/A 0.0291f
C12172 _326_/a_1108_7# _246_/B 0.00104f
C12173 _146_/C _232_/A 0.033f
C12174 _325_/a_448_7# _325_/Q 9.74e-21
C12175 _164_/A _161_/Y 0.0462f
C12176 _328_/a_651_373# _279_/A 0.00488f
C12177 _304_/S _224_/a_256_7# 4.82e-20
C12178 _294_/A _267_/A 0.324f
C12179 _275_/Y _160_/A 1.97e-21
C12180 _342_/D _323_/D 3.09e-20
C12181 _321_/Q _331_/CLK 0.316f
C12182 _188_/S _304_/a_79_n19# 2.77e-20
C12183 _229_/a_556_7# VGND -6.44e-19
C12184 _336_/a_805_7# _147_/A 8.03e-20
C12185 _295_/a_676_257# VGND -3.25e-19
C12186 _295_/a_409_7# VPWR -8.63e-19
C12187 _346_/a_193_7# VGND -0.103f
C12188 _346_/a_476_7# VPWR 0.0265f
C12189 _160_/X _173_/a_226_7# 0.0181f
C12190 _337_/D _199_/a_93_n19# 0.00154f
C12191 _193_/Y _336_/D 0.0263f
C12192 _335_/a_27_7# _204_/a_27_7# 9.11e-21
C12193 _335_/a_27_7# _208_/a_215_7# 8.23e-20
C12194 _248_/A _297_/B 0.00585f
C12195 _163_/a_78_159# VPWR 0.0144f
C12196 _343_/a_27_7# _226_/a_79_n19# 1.17e-20
C12197 _236_/a_109_257# VPWR -0.00186f
C12198 _318_/a_193_7# _248_/A 0.00234f
C12199 _345_/a_381_7# _346_/SET_B 0.00297f
C12200 _316_/a_1462_7# VGND -8.48e-19
C12201 _344_/a_956_373# _164_/A 2.32e-19
C12202 _299_/X _313_/a_27_7# 2.68e-19
C12203 _300_/a_735_7# _313_/a_1283_n19# 2.7e-20
C12204 _324_/a_639_7# _331_/CLK 1.61e-19
C12205 _346_/a_1032_373# _297_/B 5.45e-20
C12206 _346_/a_27_7# _314_/Q 1.46e-19
C12207 _340_/CLK _311_/a_193_7# 0.002f
C12208 ctln[4] input4/X 0.0179f
C12209 _332_/Q VPWR 1.86f
C12210 _276_/a_150_257# _242_/A 3.67e-19
C12211 _331_/CLK _297_/B 0.00898f
C12212 _187_/a_27_7# _143_/a_27_7# 9.19e-19
C12213 _315_/Q result[1] 0.194f
C12214 result[0] _316_/Q 8.95e-19
C12215 _318_/a_193_7# _331_/CLK 8.73e-20
C12216 _327_/a_1217_7# VGND -5.03e-19
C12217 _337_/D _336_/Q 1.06e-19
C12218 _143_/a_27_7# _315_/D 5.25e-20
C12219 _342_/a_639_7# _342_/D 0.00445f
C12220 _346_/a_586_7# _346_/D 2.11e-19
C12221 output15/a_27_7# _232_/X 3.2e-21
C12222 _194_/X _306_/S 0.00236f
C12223 _326_/a_1217_7# VGND -4.44e-19
C12224 output14/a_27_7# _322_/a_193_7# 0.0101f
C12225 _254_/A _300_/a_383_7# 6.45e-19
C12226 _215_/A _313_/a_448_7# 0.0162f
C12227 trimb[0] trimb[2] 0.0638f
C12228 _273_/A _297_/B 0.0181f
C12229 _300_/a_27_257# _157_/a_27_7# 9.66e-20
C12230 repeater43/X _324_/a_761_249# -0.0067f
C12231 _286_/B _179_/a_27_7# 0.0489f
C12232 _285_/A _258_/S 0.0135f
C12233 _216_/A _328_/Q 1.43e-20
C12234 _269_/A _228_/A 6.79e-19
C12235 _227_/A _217_/X 4.5e-21
C12236 _180_/a_111_257# VGND -1.94e-19
C12237 _324_/a_27_7# _327_/Q 2.28e-19
C12238 _343_/a_193_7# repeater43/X 0.0196f
C12239 _251_/a_79_n19# _251_/X 9.11e-19
C12240 _331_/Q _330_/a_543_7# 2.45e-19
C12241 _328_/a_1462_7# VPWR 6.83e-20
C12242 _328_/a_805_7# VGND -6.97e-19
C12243 _173_/a_76_159# VGND 0.0185f
C12244 _173_/a_489_373# VPWR 0.0377f
C12245 _251_/X _221_/a_250_257# 5.19e-20
C12246 _298_/B _323_/Q 2.4e-20
C12247 _221_/a_93_n19# _327_/D 0.00253f
C12248 _221_/a_584_7# _328_/Q 2.62e-20
C12249 repeater43/X _304_/X 0.621f
C12250 _305_/a_218_7# _286_/B 9.67e-19
C12251 _206_/A output6/a_27_7# 6.17e-19
C12252 _271_/Y _334_/a_1283_n19# 5.03e-21
C12253 _271_/A _334_/a_448_7# 0.0166f
C12254 _319_/a_543_7# VPWR 0.0201f
C12255 _319_/a_193_7# VGND 0.0383f
C12256 _323_/a_27_7# _229_/a_76_159# 5.24e-22
C12257 _346_/SET_B _220_/a_584_7# 5.68e-20
C12258 _345_/a_193_7# clkbuf_2_3_0_clk/A 5.48e-21
C12259 _346_/SET_B _311_/a_761_249# 0.0111f
C12260 _337_/a_193_7# VPWR -0.262f
C12261 _321_/a_1462_7# result[7] 3.47e-20
C12262 _167_/X _306_/S 2.47e-19
C12263 _216_/a_27_7# VPWR 0.156f
C12264 _258_/S _258_/a_535_334# 0.00181f
C12265 _319_/a_1108_7# _297_/B 1.7e-19
C12266 _343_/CLK _315_/D 0.0617f
C12267 _215_/A _191_/B 1.01e-19
C12268 _313_/D _196_/A 1.46e-19
C12269 _340_/a_27_7# _305_/a_76_159# 1.38e-20
C12270 _334_/a_805_7# VGND -7.97e-19
C12271 _334_/a_1462_7# VPWR 2.22e-19
C12272 clk _209_/a_109_7# 8.26e-19
C12273 _189_/a_27_7# _281_/Y 0.00738f
C12274 _321_/a_1108_7# _280_/a_68_257# 2.62e-20
C12275 _167_/a_27_257# _166_/Y 0.0594f
C12276 _255_/a_112_257# _306_/S 6.78e-20
C12277 _258_/S _172_/A 2.48e-20
C12278 _309_/a_1108_7# _340_/CLK 1.59e-20
C12279 _316_/D _246_/B 0.358f
C12280 _158_/Y _160_/X 0.152f
C12281 _149_/a_27_7# _341_/Q 1.95e-19
C12282 cal _209_/X 0.267f
C12283 _320_/Q _320_/a_1283_n19# 0.00312f
C12284 _238_/B _320_/a_193_7# 6.09e-19
C12285 _200_/a_250_257# _293_/a_39_257# 4.96e-21
C12286 _281_/Y _255_/B 7.93e-20
C12287 _345_/a_1032_373# _345_/Q 0.0581f
C12288 _345_/a_193_7# _172_/Y 1.17e-19
C12289 _345_/a_1182_221# _345_/D 2.73e-19
C12290 _296_/Y _227_/A 0.66f
C12291 _168_/a_109_7# _301_/a_51_257# 0.00126f
C12292 _294_/A _194_/X 0.00114f
C12293 _339_/D _336_/Q 0.0274f
C12294 _325_/a_448_7# _326_/Q 0.00123f
C12295 _196_/A _197_/X 0.0174f
C12296 _258_/S _198_/a_250_257# 4.54e-21
C12297 _324_/a_1108_7# _304_/S 0.0394f
C12298 _283_/Y _332_/a_1283_n19# 6.57e-20
C12299 _327_/a_27_7# _214_/a_27_257# 6.34e-21
C12300 _258_/a_505_n19# _260_/B 5.83e-20
C12301 _188_/a_76_159# _271_/A 0.00338f
C12302 _316_/Q _316_/D 0.149f
C12303 _329_/a_1462_7# _281_/A 3.42e-19
C12304 _254_/Y _267_/A 0.0104f
C12305 _326_/a_27_7# _214_/a_27_257# 0.00953f
C12306 repeater43/X _272_/a_39_257# 0.00232f
C12307 _268_/a_39_257# _317_/D 0.00254f
C12308 _306_/S _296_/a_109_7# 0.00202f
C12309 _304_/S _324_/D 0.0207f
C12310 _340_/a_1283_n19# _198_/a_93_n19# 5.9e-19
C12311 _273_/A _311_/a_1108_7# 3.27e-21
C12312 _254_/A _346_/D 0.116f
C12313 _275_/A _314_/Q 1.44e-20
C12314 _286_/B _172_/B 1.21e-20
C12315 _226_/a_382_257# VPWR -2.33e-19
C12316 _188_/a_218_7# VGND 3.68e-20
C12317 _292_/A _171_/a_292_257# 0.00208f
C12318 _325_/a_27_7# _324_/a_27_7# 0.00102f
C12319 _294_/A _167_/X 3.66e-21
C12320 _346_/a_1224_7# VPWR 2.28e-20
C12321 _346_/a_796_7# VGND -4.28e-19
C12322 _333_/a_27_7# _333_/a_639_7# -0.0015f
C12323 _335_/a_1108_7# _332_/Q 5.62e-20
C12324 _335_/a_1283_n19# _333_/Q 7.66e-19
C12325 _320_/Q _232_/X 0.054f
C12326 _309_/a_448_7# _346_/SET_B 0.00176f
C12327 _335_/a_448_7# _207_/X 1.8e-19
C12328 _342_/a_543_7# _343_/Q 1.73e-19
C12329 _248_/B _221_/a_93_n19# 5.83e-20
C12330 _343_/a_1108_7# _147_/A 4.53e-20
C12331 _343_/a_761_249# _226_/X 5.44e-20
C12332 _339_/a_193_7# VPWR 0.0247f
C12333 _341_/a_193_7# _244_/B 8.07e-19
C12334 _300_/Y _313_/a_448_7# 1.45e-19
C12335 _327_/a_193_7# _232_/X 0.0169f
C12336 _271_/A _143_/a_109_7# 6.22e-20
C12337 _282_/a_39_257# VPWR 0.0417f
C12338 _317_/a_1283_n19# _242_/B 4.65e-19
C12339 _275_/Y _273_/A 0.00811f
C12340 _255_/X _216_/A 6.44e-20
C12341 repeater43/a_27_7# _271_/Y 0.0548f
C12342 _343_/a_1108_7# _149_/A 0.00199f
C12343 _323_/a_1108_7# _334_/a_193_7# 9.49e-21
C12344 _283_/Y _338_/a_651_373# 1.08e-19
C12345 _283_/A _194_/X 0.00709f
C12346 _323_/a_27_7# _334_/a_448_7# 2.62e-20
C12347 _326_/a_193_7# _232_/X 0.00842f
C12348 trimb[2] trimb[3] 0.055f
C12349 output22/a_27_7# _342_/a_27_7# 3.56e-22
C12350 trimb[1] _288_/Y 0.0206f
C12351 _290_/A _297_/Y 0.0244f
C12352 clkbuf_2_3_0_clk/A VPWR 1.11f
C12353 _330_/Q _212_/X 0.118f
C12354 _169_/a_109_257# _267_/A 0.00294f
C12355 clk _154_/A 0.23f
C12356 ctlp[0] _322_/a_448_7# 3.93e-21
C12357 repeater43/X VGND 4.39f
C12358 _312_/a_543_7# _312_/D 2.39e-19
C12359 _292_/A _161_/Y 0.0143f
C12360 _215_/A _337_/Q 1.19e-19
C12361 input1/X _336_/a_651_373# 8.49e-19
C12362 _328_/a_27_7# _232_/X 0.00311f
C12363 _271_/A _206_/A 0.082f
C12364 _340_/a_193_7# _254_/B 1.07e-21
C12365 _288_/Y VGND 0.255f
C12366 _277_/Y _337_/Q 0.0114f
C12367 _327_/Q VPWR 1.94f
C12368 _330_/D _346_/SET_B 0.0101f
C12369 _340_/CLK _153_/B 5.02e-19
C12370 output40/a_27_7# trimb[4] 0.00878f
C12371 _223_/a_93_n19# _223_/a_250_257# -6.97e-22
C12372 _335_/a_27_7# _206_/A 1.12e-21
C12373 output32/a_27_7# trim[1] 0.0074f
C12374 repeater43/X _318_/a_1108_7# 0.0241f
C12375 _161_/Y _160_/A 0.508f
C12376 _267_/B _309_/Q 0.0481f
C12377 _343_/a_1462_7# repeater43/X 4.76e-19
C12378 _316_/a_27_7# _317_/D 0.0119f
C12379 _172_/Y VPWR 0.593f
C12380 _329_/a_193_7# _329_/a_651_373# -0.00701f
C12381 _329_/a_543_7# _327_/D 8.05e-19
C12382 _290_/A _310_/a_193_7# 0.00365f
C12383 ctln[5] _283_/Y 0.0139f
C12384 _297_/B _217_/X 0.44f
C12385 _314_/D _212_/X 1.35e-22
C12386 _319_/Q _242_/A 0.295f
C12387 _271_/A _334_/D 0.167f
C12388 _331_/a_1108_7# _217_/A 1.03e-20
C12389 _319_/a_1462_7# VGND -8.4e-19
C12390 _313_/a_1270_373# VPWR -2.54e-19
C12391 _313_/a_448_7# VGND -0.00529f
C12392 output7/a_27_7# _271_/A 4.11e-19
C12393 _337_/a_1462_7# VPWR 1.18e-19
C12394 _337_/a_805_7# VGND -6.12e-19
C12395 _328_/a_1108_7# output19/a_27_7# 2.13e-19
C12396 _335_/a_27_7# _334_/D 1.05e-19
C12397 _335_/a_193_7# _343_/CLK 0.0051f
C12398 _335_/D _334_/a_27_7# 1.88e-21
C12399 _342_/a_1108_7# _341_/a_1108_7# 5.35e-21
C12400 output7/a_27_7# _335_/a_27_7# 0.0137f
C12401 _301_/X _170_/a_226_7# 2.93e-19
C12402 _250_/a_78_159# _336_/Q 3.73e-20
C12403 input2/a_27_7# comp 0.0152f
C12404 _320_/Q _322_/a_1270_373# 3.72e-19
C12405 _160_/X _160_/a_27_7# 0.00172f
C12406 _334_/Q VGND 0.109f
C12407 input1/X _153_/A 1.61e-20
C12408 ctln[1] VPWR 0.233f
C12409 _344_/a_27_7# _163_/a_78_159# 8.39e-19
C12410 clkbuf_2_1_0_clk/A cal 0.135f
C12411 _254_/Y _194_/X 2.65e-20
C12412 _315_/a_761_249# _286_/Y 9.69e-22
C12413 _271_/A _191_/a_109_257# 1.03e-19
C12414 _320_/D _320_/Q 6.41e-20
C12415 ctln[2] VPWR 0.201f
C12416 output25/a_27_7# _316_/a_1108_7# 1.65e-20
C12417 _147_/Y _347_/a_27_7# 1.41e-19
C12418 result[0] _244_/a_109_257# 0.00131f
C12419 output22/a_27_7# _317_/D 1.62e-19
C12420 rstn _340_/Q 0.0829f
C12421 input4/a_27_7# _340_/D 9.18e-20
C12422 _267_/B _311_/a_193_7# 3.56e-19
C12423 _172_/A _295_/a_306_7# 1.75e-19
C12424 _342_/a_543_7# _229_/a_76_159# 0.00304f
C12425 _296_/Y _297_/B 2.46e-20
C12426 _265_/B _284_/A 0.00647f
C12427 _210_/a_27_7# _306_/S 0.0307f
C12428 _254_/A _314_/Q 4.84e-20
C12429 _271_/A _147_/A 0.352f
C12430 _313_/Q _260_/B 0.00283f
C12431 _144_/A _246_/B 1.6e-20
C12432 _319_/Q _322_/D 0.376f
C12433 _191_/B VGND 0.556f
C12434 _192_/B VPWR 2.02f
C12435 repeater43/a_27_7# _323_/a_761_249# 2.95e-22
C12436 _162_/X _299_/a_78_159# 2.89e-19
C12437 _319_/Q _321_/a_448_7# 4.51e-20
C12438 _258_/a_76_159# _190_/A 1.97e-20
C12439 _327_/a_27_7# _318_/Q 6.11e-19
C12440 _324_/Q _315_/a_651_373# 4.18e-20
C12441 _340_/a_1270_373# _197_/X 3.81e-19
C12442 _271_/A _149_/A 0.231f
C12443 _277_/Y _339_/Q 0.0114f
C12444 _326_/a_27_7# _318_/Q 1.38e-19
C12445 _342_/D _177_/A 0.00335f
C12446 _216_/A _336_/a_193_7# 5.81e-22
C12447 _302_/a_323_257# _300_/Y 0.00637f
C12448 _328_/a_27_7# _320_/D 1.75e-21
C12449 _325_/a_27_7# VPWR 0.0375f
C12450 _283_/Y _334_/a_448_7# 1.84e-19
C12451 ctln[7] _334_/a_1283_n19# 1.25e-21
C12452 _305_/a_505_n19# _340_/CLK 0.00714f
C12453 _157_/A _314_/a_651_373# 2.12e-19
C12454 _211_/a_27_257# _332_/Q 0.0511f
C12455 _323_/a_27_7# _206_/A 6.57e-19
C12456 _333_/a_543_7# _333_/D 0.0102f
C12457 _320_/a_448_7# _319_/a_27_7# 3.28e-20
C12458 clkbuf_0_clk/a_110_7# _297_/B 9.38e-19
C12459 _335_/D _207_/X 0.0223f
C12460 _339_/a_805_7# VGND -6.97e-19
C12461 _339_/a_1462_7# VPWR 6.95e-20
C12462 _341_/a_1462_7# _244_/B 2.71e-19
C12463 _341_/a_805_7# _317_/D 3.41e-19
C12464 _261_/A _310_/D 2.19e-19
C12465 _327_/a_1462_7# _232_/X 1.42e-19
C12466 _333_/a_27_7# _332_/a_1283_n19# 7.4e-21
C12467 _333_/a_1283_n19# _332_/a_27_7# 9.12e-21
C12468 clkbuf_0_clk/X _217_/A 0.00566f
C12469 _325_/a_639_7# _304_/X 0.00432f
C12470 _325_/a_1270_373# _217_/A 2.78e-20
C12471 _317_/a_1108_7# VPWR 0.053f
C12472 _317_/a_543_7# VGND 0.0183f
C12473 _294_/Y clkc 0.0173f
C12474 _323_/a_193_7# _343_/CLK 0.314f
C12475 _323_/a_27_7# _334_/D 4.25e-19
C12476 _169_/Y _344_/D 0.00155f
C12477 _283_/Y _346_/SET_B 0.00158f
C12478 _182_/a_79_n19# _182_/X 7.45e-19
C12479 _182_/a_215_7# _196_/A 0.0114f
C12480 _326_/a_1462_7# _232_/X 7.88e-20
C12481 trimb[2] VPWR 0.211f
C12482 _265_/a_109_257# _310_/D 8.7e-19
C12483 _172_/a_109_257# VGND -6.79e-19
C12484 _336_/a_448_7# _336_/D 0.00232f
C12485 _336_/a_1270_373# _284_/A 1.41e-19
C12486 _330_/Q _331_/a_639_7# 0.00101f
C12487 _172_/A _173_/a_226_7# 0.0036f
C12488 _258_/S _312_/a_448_7# 1.74e-19
C12489 output24/a_27_7# _317_/Q 0.0371f
C12490 _284_/a_39_257# _267_/A 1.66e-21
C12491 _318_/a_193_7# _317_/a_651_373# 6.94e-21
C12492 _169_/B _166_/Y 4.33e-20
C12493 _169_/Y _346_/Q 0.00119f
C12494 _281_/Y _326_/Q 4.18e-20
C12495 _292_/A _312_/a_543_7# 5.3e-19
C12496 _314_/a_27_7# _284_/A 2.83e-19
C12497 _194_/a_27_7# _267_/A 3.72e-19
C12498 _309_/a_1108_7# _267_/B 3.08e-19
C12499 _309_/a_543_7# _309_/D 2.04e-19
C12500 _308_/S _307_/a_535_334# 8.39e-19
C12501 _308_/a_505_n19# _145_/A 1.1e-20
C12502 _317_/Q _270_/a_39_257# 2.38e-19
C12503 _340_/a_1283_n19# _147_/Y 1.67e-21
C12504 _331_/a_448_7# VGND 0.00171f
C12505 _320_/a_639_7# _346_/SET_B 0.00347f
C12506 _310_/a_27_7# _297_/Y 2.31e-21
C12507 _181_/X _162_/X 0.488f
C12508 _294_/A _310_/a_1108_7# 2.04e-21
C12509 _302_/a_227_7# VPWR 0.00524f
C12510 _302_/a_323_257# VGND -5.16e-19
C12511 _169_/Y _168_/a_481_7# 5.38e-20
C12512 _344_/a_1602_7# _346_/SET_B 1.36e-20
C12513 _343_/a_543_7# cal 0.00539f
C12514 _308_/a_218_7# _192_/B 0.00216f
C12515 _290_/A _310_/a_1462_7# 3.59e-19
C12516 _163_/a_493_257# _161_/Y 1.86e-19
C12517 _308_/S _178_/a_193_257# 5.71e-21
C12518 _336_/a_761_249# _193_/Y 1.91e-20
C12519 _336_/a_1283_n19# _340_/Q 5.18e-20
C12520 _336_/a_1108_7# _194_/X 7.1e-19
C12521 _230_/a_27_7# _232_/A 5.39e-19
C12522 _338_/Q _311_/Q 0.344f
C12523 _285_/A _158_/Y 0.00175f
C12524 _337_/Q VGND 1.02f
C12525 _335_/a_1462_7# _343_/CLK 2.64e-19
C12526 _335_/a_651_373# _334_/Q 2.53e-20
C12527 _182_/a_297_257# _343_/Q 1.09e-20
C12528 _322_/a_193_7# _321_/D 2.62e-19
C12529 _303_/A _304_/X 0.0017f
C12530 _325_/a_543_7# _246_/B 1.74e-20
C12531 _315_/a_651_373# _228_/A 8.7e-19
C12532 _342_/D _341_/a_1283_n19# 1.19e-20
C12533 _322_/a_1108_7# _331_/CLK 8.41e-19
C12534 ctln[1] _335_/a_1108_7# 4.83e-20
C12535 _310_/a_27_7# _310_/a_193_7# -0.29f
C12536 clkbuf_2_1_0_clk/A _284_/A 0.00696f
C12537 _321_/a_543_7# _269_/A 3e-21
C12538 _281_/Y _314_/a_193_7# 7.32e-20
C12539 _323_/a_27_7# _149_/A 5.54e-20
C12540 _273_/A _161_/Y 0.207f
C12541 _307_/a_76_159# _188_/S 6.74e-22
C12542 clkbuf_0_clk/X _220_/a_250_257# 5.6e-19
C12543 output13/a_27_7# repeater43/X 1.2e-20
C12544 _310_/Q _284_/A 3.82e-19
C12545 _197_/X _338_/D 0.0733f
C12546 _210_/a_27_7# _283_/A 4.38e-21
C12547 result[6] VGND 0.144f
C12548 _186_/a_79_n19# _147_/A 0.00508f
C12549 _172_/A _226_/a_79_n19# 2.78e-19
C12550 _324_/a_543_7# _286_/Y 0.00337f
C12551 _184_/a_505_n19# _192_/B 1.03e-19
C12552 output25/a_27_7# _331_/CLK 0.0615f
C12553 _318_/Q _316_/a_1462_7# 3.28e-20
C12554 _342_/a_448_7# _248_/A 2.35e-20
C12555 _345_/a_27_7# _344_/Q 1.57e-21
C12556 _309_/a_761_249# _337_/Q 9.17e-20
C12557 _346_/Q _170_/a_226_257# 1.33e-19
C12558 ctln[6] _153_/A 5.33e-20
C12559 _281_/Y _154_/A 9.41e-21
C12560 _186_/a_79_n19# _149_/A 0.00636f
C12561 _146_/C VPWR 0.237f
C12562 _344_/a_27_7# clkbuf_2_3_0_clk/A 3.52e-21
C12563 repeater43/X _323_/a_651_373# 0.00182f
C12564 _172_/A _158_/Y 5.66e-21
C12565 _283_/Y _206_/A 6.63e-20
C12566 _184_/a_439_7# _150_/C 7.82e-19
C12567 _188_/S _226_/a_297_7# 1.49e-19
C12568 _192_/a_68_257# _194_/A 0.00102f
C12569 repeater43/X _214_/a_27_257# 0.00273f
C12570 _217_/A _286_/Y 0.23f
C12571 _330_/D _331_/a_761_249# 8.45e-20
C12572 _320_/a_193_7# _217_/X 3.17e-20
C12573 _162_/X _347_/a_1108_7# 3.16e-20
C12574 _320_/Q _297_/A 1.02e-22
C12575 _157_/A VPWR 0.653f
C12576 _346_/D _286_/Y 6.44e-20
C12577 _225_/X _153_/B 0.00232f
C12578 _324_/a_1270_373# _324_/Q 1.29e-19
C12579 _303_/A _300_/Y 0.00282f
C12580 _325_/a_639_7# VGND -0.00113f
C12581 _339_/a_193_7# _198_/a_93_n19# 3.46e-22
C12582 _283_/Y _334_/D 5.79e-19
C12583 output26/a_27_7# _318_/a_27_7# 9.3e-19
C12584 cal _311_/a_27_7# 8.53e-20
C12585 output7/a_27_7# _283_/Y 3.26e-21
C12586 _286_/B _305_/X 0.174f
C12587 _324_/a_27_7# _221_/a_250_257# 2.08e-20
C12588 _344_/a_1182_221# _345_/Q 0.00917f
C12589 clkbuf_0_clk/X _314_/Q 4.53e-21
C12590 _341_/Q _306_/S 7.1e-20
C12591 _339_/Q VGND 0.844f
C12592 _194_/X _194_/a_27_7# 0.024f
C12593 _338_/Q _254_/B 0.00327f
C12594 _338_/D _312_/a_193_7# 9.32e-21
C12595 _346_/SET_B _312_/a_27_7# 0.00569f
C12596 _292_/A _263_/B 0.00994f
C12597 _342_/Q _209_/X 1.21e-20
C12598 _202_/a_584_7# VPWR -8.09e-19
C12599 _202_/a_256_7# VGND -0.00131f
C12600 _297_/A _347_/a_805_7# 0.00238f
C12601 _160_/X _267_/A 5.23e-20
C12602 output27/a_27_7# result[6] 0.00521f
C12603 _324_/a_1283_n19# _284_/A 1.07e-19
C12604 _258_/S _312_/D 4.29e-19
C12605 _219_/a_256_7# _279_/A 5.31e-19
C12606 _313_/D _313_/a_193_7# -0.00498f
C12607 _347_/a_27_7# _347_/a_193_7# -0.0371f
C12608 _341_/a_193_7# _177_/A 6.62e-20
C12609 _168_/a_397_257# _299_/X 0.00154f
C12610 _340_/a_193_7# _196_/A 0.00888f
C12611 _346_/a_476_7# _147_/Y 4.58e-21
C12612 _269_/A _315_/a_761_249# 0.00748f
C12613 _325_/Q _242_/A 1.04e-20
C12614 input3/a_27_7# _269_/A 0.0117f
C12615 _163_/a_78_159# _147_/Y 1.69e-19
C12616 _323_/a_448_7# _323_/Q 1.22e-19
C12617 _303_/A VGND 0.375f
C12618 _260_/A VPWR 0.987f
C12619 _197_/X _337_/a_1108_7# 0.00102f
C12620 _189_/a_27_7# _336_/Q 0.00156f
C12621 _188_/a_76_159# _231_/a_79_n19# 7.12e-21
C12622 _342_/a_1283_n19# _343_/CLK 1.24e-20
C12623 _212_/a_27_7# _212_/X 0.00213f
C12624 _304_/a_79_n19# _216_/X 0.00204f
C12625 _255_/B _336_/Q 4.84e-20
C12626 _324_/Q _246_/B 2.27e-20
C12627 _172_/A _157_/a_27_7# 0.0221f
C12628 _281_/Y _324_/a_1108_7# 8.39e-20
C12629 _285_/A _160_/a_27_7# 0.00654f
C12630 _197_/X _343_/CLK 9.79e-21
C12631 _216_/A _299_/X 1.79e-20
C12632 _181_/X _298_/C 0.67f
C12633 _343_/D input3/a_27_7# 0.00188f
C12634 _323_/a_1217_7# _149_/A 5.91e-20
C12635 _324_/a_1270_373# _228_/A 2.78e-20
C12636 _261_/A VPWR 0.176f
C12637 _340_/CLK _263_/a_109_257# 5.25e-21
C12638 _239_/a_113_257# VPWR 0.0524f
C12639 _281_/Y _324_/D 0.0105f
C12640 output18/a_27_7# _319_/a_1283_n19# 1.83e-22
C12641 _316_/Q _324_/Q 0.0037f
C12642 _265_/B _310_/a_761_249# 6.87e-19
C12643 _345_/a_27_7# _306_/S 1.37e-20
C12644 _265_/a_109_257# VPWR 6.87e-19
C12645 _335_/D _323_/Q 3.78e-21
C12646 _173_/a_489_373# _147_/Y 3.2e-19
C12647 _342_/a_27_7# _226_/X 0.00141f
C12648 _153_/a_215_257# _204_/Y 1.84e-20
C12649 _153_/a_297_257# _335_/Q 0.00438f
C12650 _342_/D _248_/A 0.00931f
C12651 _342_/Q _315_/a_543_7# 2.36e-20
C12652 _264_/a_113_257# _265_/B 0.00508f
C12653 _314_/Q _286_/Y 5.23e-20
C12654 _167_/a_27_257# _170_/a_489_373# 2.64e-20
C12655 _333_/a_543_7# _190_/A 8.48e-19
C12656 _333_/a_1108_7# _332_/Q 0.0122f
C12657 _333_/a_1283_n19# _333_/Q 0.0654f
C12658 _254_/Y _336_/a_543_7# 0.0298f
C12659 _309_/a_193_7# _267_/A 1.73e-19
C12660 _341_/a_193_7# _341_/a_1283_n19# -4.45e-19
C12661 _283_/Y _337_/D 4.16e-21
C12662 result[4] VGND 0.186f
C12663 _343_/Q _298_/C 0.792f
C12664 repeater43/X _330_/a_27_7# 0.00541f
C12665 _260_/B _347_/a_27_7# 2.11e-20
C12666 clk _153_/B 0.0711f
C12667 repeater43/X _318_/Q 0.17f
C12668 _341_/Q _283_/A 2.03e-19
C12669 _197_/X _339_/a_1108_7# 1.85e-19
C12670 _314_/a_193_7# _297_/Y 0.00158f
C12671 _345_/a_193_7# _165_/X 6.7e-19
C12672 _227_/a_113_7# _327_/Q 4.91e-20
C12673 _251_/a_79_n19# VPWR 0.0502f
C12674 _281_/A _246_/B 9.7e-21
C12675 _338_/a_193_7# _338_/a_1283_n19# -5.93e-19
C12676 _221_/a_250_257# VPWR 0.0363f
C12677 result[4] _318_/a_1108_7# 2.17e-19
C12678 _324_/a_27_7# _251_/X 1.36e-19
C12679 _254_/A _254_/B 0.0788f
C12680 _281_/Y _218_/a_250_257# 0.0083f
C12681 _170_/a_226_7# _297_/Y 5.45e-20
C12682 _342_/a_805_7# repeater43/X -0.00125f
C12683 _191_/B _203_/a_209_257# 0.00254f
C12684 _346_/SET_B _312_/a_1217_7# 4.88e-19
C12685 _329_/a_761_249# _304_/X 5.07e-19
C12686 _326_/a_193_7# _325_/D 4.73e-21
C12687 _336_/D VGND 0.393f
C12688 _217_/A _328_/Q 0.00157f
C12689 _258_/S _292_/A 0.00642f
C12690 _322_/a_1283_n19# output28/a_27_7# 7.51e-19
C12691 _333_/a_27_7# _206_/A 0.615f
C12692 _288_/A _346_/SET_B 0.00365f
C12693 _184_/a_439_7# cal 1.86e-19
C12694 _184_/a_218_7# input1/X 7.76e-19
C12695 _279_/Y _305_/X 0.0108f
C12696 _313_/Q _313_/a_639_7# 2.41e-20
C12697 _329_/D _279_/A 9e-21
C12698 repeater42/a_27_7# _221_/a_93_n19# 0.0117f
C12699 _242_/A _326_/Q 0.0245f
C12700 _340_/a_651_373# _338_/a_27_7# 3.74e-21
C12701 _340_/a_1283_n19# _338_/a_543_7# 3.08e-22
C12702 _341_/Q _248_/B 0.0376f
C12703 _162_/X _346_/SET_B 0.0541f
C12704 _196_/A _295_/a_79_n19# 0.061f
C12705 _306_/a_505_n19# _267_/A 0.00787f
C12706 _167_/X _160_/X 0.0108f
C12707 _317_/D _226_/X 7.97e-20
C12708 _287_/a_39_257# _346_/SET_B 3.07e-19
C12709 _329_/D _218_/a_250_257# 2.92e-19
C12710 _269_/A _318_/D 0.182f
C12711 repeater43/X _241_/a_199_7# 7.51e-20
C12712 _164_/A _173_/a_226_7# 1.05e-19
C12713 _343_/CLK _333_/a_193_7# 7.9e-19
C12714 _316_/Q _228_/A 1.49e-21
C12715 _248_/a_109_257# _327_/Q 9.17e-22
C12716 _323_/D _323_/Q 1.09e-19
C12717 result[4] output27/a_27_7# 2.55e-19
C12718 output26/a_27_7# result[5] 0.00139f
C12719 _309_/D _254_/B 9.65e-21
C12720 clk _181_/a_27_7# 9.98e-19
C12721 _340_/Q VPWR 0.22f
C12722 _309_/a_1283_n19# _284_/A 0.0918f
C12723 _227_/A _205_/a_297_7# 0.0352f
C12724 _273_/A _263_/B 0.00757f
C12725 _317_/a_1283_n19# _244_/B 1.64e-19
C12726 _317_/a_761_249# _317_/D 0.00196f
C12727 _216_/A _246_/B 9.68e-19
C12728 _319_/Q _271_/A 0.0529f
C12729 _229_/a_226_7# valid 1.95e-19
C12730 _315_/Q _341_/a_761_249# 1.93e-21
C12731 result[0] _341_/a_27_7# 0.0128f
C12732 _293_/a_39_257# cal 2.75e-20
C12733 clkbuf_2_3_0_clk/A _147_/Y 0.0194f
C12734 _310_/a_761_249# _310_/Q 3.71e-19
C12735 _310_/a_448_7# _310_/D 0.0145f
C12736 _329_/a_27_7# _218_/a_93_n19# 1.39e-19
C12737 _327_/a_543_7# _216_/X 0.00717f
C12738 _209_/X _225_/B 9.91e-21
C12739 _336_/a_193_7# _336_/a_651_373# -0.00701f
C12740 _196_/A _180_/a_29_13# 3.86e-20
C12741 _325_/Q _224_/a_346_7# 0.00426f
C12742 _270_/a_39_257# _304_/X 1.81e-20
C12743 _264_/a_113_257# _310_/Q 2.9e-20
C12744 _320_/Q _238_/B 0.0206f
C12745 _343_/a_761_249# _343_/D 6.89e-19
C12746 _343_/a_1283_n19# _185_/A 8.3e-20
C12747 _165_/X VPWR 0.485f
C12748 _231_/a_306_7# _144_/A 2.89e-19
C12749 _286_/B _173_/a_76_159# 0.00738f
C12750 _327_/a_193_7# _238_/B 2.55e-19
C12751 _327_/a_543_7# _329_/Q 2e-21
C12752 _172_/Y _147_/Y 0.0947f
C12753 ctln[4] input4/a_27_7# 0.00102f
C12754 _340_/CLK _312_/Q 4.76e-20
C12755 _288_/Y output40/a_27_7# 1.46e-19
C12756 _154_/A _335_/Q 3.19e-19
C12757 _327_/a_193_7# _327_/a_1283_n19# -5.93e-19
C12758 _322_/a_1270_373# result[7] 4.19e-20
C12759 _255_/a_184_257# VPWR -7.16e-19
C12760 _255_/a_30_13# VGND 0.043f
C12761 result[3] _317_/a_193_7# 0.00109f
C12762 _318_/Q _317_/a_543_7# 2.24e-20
C12763 output15/a_27_7# _331_/CLK 1.91e-20
C12764 clkbuf_1_0_0_clk/a_75_172# VGND 0.0557f
C12765 _324_/a_1283_n19# _342_/Q 6.53e-21
C12766 _323_/a_639_7# cal 8.53e-19
C12767 _315_/Q _316_/a_543_7# 3.01e-19
C12768 _329_/a_1108_7# _330_/Q 0.0053f
C12769 _330_/Q _327_/D 0.0012f
C12770 repeater43/X _330_/a_1217_7# 4.9e-19
C12771 _277_/Y _319_/D 2.11e-19
C12772 _332_/a_27_7# _332_/Q 0.0135f
C12773 _331_/a_761_249# _330_/a_1283_n19# 5.29e-20
C12774 _331_/a_27_7# _330_/a_448_7# 1.8e-20
C12775 _331_/a_193_7# _330_/a_1108_7# 7.02e-21
C12776 _332_/a_193_7# _207_/X 9.94e-22
C12777 _326_/a_193_7# _326_/a_1283_n19# -6.53e-19
C12778 _162_/X _313_/a_761_249# 2.93e-19
C12779 _328_/a_761_249# _329_/Q 0.0308f
C12780 _328_/a_543_7# _320_/Q 4.79e-19
C12781 _305_/a_76_159# _197_/a_27_7# 5.76e-19
C12782 trimb[1] input2/a_27_7# 0.00273f
C12783 _298_/B _175_/Y 0.0101f
C12784 _251_/X VPWR 0.564f
C12785 _329_/a_1283_n19# VPWR 0.0335f
C12786 _329_/a_761_249# VGND -0.007f
C12787 _328_/a_27_7# _327_/a_1283_n19# 0.001f
C12788 _308_/a_535_334# _306_/S 2.17e-19
C12789 _296_/a_213_83# VPWR 0.0018f
C12790 _296_/a_493_257# VGND -7.67e-20
C12791 _259_/a_199_7# _338_/Q 4.9e-19
C12792 _308_/X input1/X 0.787f
C12793 _285_/A _267_/A 0.00788f
C12794 _306_/a_76_159# _340_/Q 0.00347f
C12795 input2/a_27_7# VGND 0.0533f
C12796 _341_/a_193_7# _248_/A 0.0149f
C12797 _314_/Q _328_/Q 2.67e-20
C12798 _342_/a_193_7# cal 8.06e-19
C12799 _192_/B _147_/Y 0.0124f
C12800 _162_/X _156_/a_39_257# 0.0414f
C12801 _322_/a_639_7# result[6] 8.64e-19
C12802 _333_/a_639_7# _207_/C 6.89e-19
C12803 _332_/a_1283_n19# _332_/D 4.66e-20
C12804 _301_/a_240_7# _299_/X 0.035f
C12805 _301_/a_51_257# _160_/X 0.0147f
C12806 _319_/Q _330_/D 0.00932f
C12807 _232_/A _245_/a_113_257# 8.93e-20
C12808 _309_/Q _297_/Y 0.00708f
C12809 _330_/Q _283_/A 0.574f
C12810 _329_/a_543_7# repeater42/a_27_7# 1.5e-19
C12811 _182_/a_79_n19# _225_/X 0.07f
C12812 _340_/a_27_7# _346_/SET_B 0.0259f
C12813 _160_/X clkbuf_1_1_0_clk/a_75_172# 0.00959f
C12814 output16/a_27_7# trimb[2] 2.55e-19
C12815 ctlp[2] output38/a_27_7# 3.88e-19
C12816 _200_/a_93_n19# _340_/CLK 6.6e-20
C12817 _328_/a_193_7# _328_/a_761_249# -0.0105f
C12818 _328_/a_27_7# _328_/a_543_7# -0.00936f
C12819 _347_/a_448_7# _347_/D 0.00397f
C12820 _198_/a_93_n19# _260_/A 5.83e-20
C12821 _317_/Q _321_/Q 1.05e-20
C12822 _267_/a_109_257# _263_/B 0.00125f
C12823 _164_/Y _345_/D 2.41e-20
C12824 _167_/X _306_/a_505_n19# 1.05e-21
C12825 _314_/a_27_7# _225_/B 5.23e-20
C12826 _172_/A _267_/A 1.32f
C12827 _258_/S _190_/A 8.9e-20
C12828 output24/a_27_7# VGND 0.113f
C12829 _162_/X _147_/A 0.00857f
C12830 _293_/a_39_257# _284_/A 1.03e-19
C12831 _230_/a_27_7# VPWR 0.0617f
C12832 _316_/a_761_249# _248_/A 0.00936f
C12833 _205_/a_79_n19# VPWR 0.0195f
C12834 _281_/Y _153_/B 0.0566f
C12835 clkbuf_2_1_0_clk/A _199_/a_250_257# 0.00526f
C12836 _269_/A _318_/a_448_7# 2.94e-20
C12837 _169_/Y _170_/a_76_159# 0.00212f
C12838 _297_/A _157_/a_27_7# 0.00154f
C12839 _177_/A _226_/a_79_n19# 3.23e-20
C12840 _258_/S _273_/A 0.0119f
C12841 _308_/X _286_/Y 1.57e-21
C12842 _346_/a_193_7# _279_/Y 6.19e-21
C12843 _343_/a_27_7# _175_/Y 0.0084f
C12844 _270_/a_39_257# VGND 0.0449f
C12845 _254_/B _202_/a_250_257# 3.04e-19
C12846 _320_/Q _248_/A 0.026f
C12847 _330_/Q _248_/B 2.68e-20
C12848 _317_/Q _318_/a_193_7# 9.26e-22
C12849 _342_/a_27_7# _286_/Y 0.00804f
C12850 output22/a_27_7# _341_/D 0.00197f
C12851 result[0] _341_/a_1217_7# 1.07e-20
C12852 _333_/a_651_373# _191_/B 0.0287f
C12853 clkbuf_0_clk/X _331_/D 2.29e-21
C12854 _331_/Q _331_/a_543_7# 0.0313f
C12855 _319_/Q _232_/a_27_7# 1.64e-21
C12856 _326_/Q _224_/a_346_7# 4.01e-19
C12857 _316_/a_193_7# _316_/D 0.0896f
C12858 _236_/B _316_/a_27_7# 1.6e-21
C12859 _316_/a_761_249# _331_/CLK 2.4e-19
C12860 _340_/a_543_7# _190_/A 2.42e-20
C12861 _268_/a_39_257# _343_/CLK 1.11e-20
C12862 _227_/A _298_/A 0.472f
C12863 clkbuf_0_clk/X _330_/a_193_7# 7.74e-20
C12864 _311_/a_193_7# _297_/Y 1.73e-20
C12865 repeater43/X _286_/B 0.00226f
C12866 _338_/a_1270_373# _340_/CLK 6.39e-19
C12867 input1/X _203_/a_209_7# 3.49e-19
C12868 _301_/a_245_257# VPWR -6.18e-20
C12869 _320_/Q _331_/CLK 0.146f
C12870 _306_/X _157_/A 3.21e-21
C12871 input1/X _254_/B 0.163f
C12872 _232_/A VPWR 0.78f
C12873 _169_/Y clkbuf_2_1_0_clk/A 0.0543f
C12874 _326_/a_193_7# _248_/A 5.42e-19
C12875 _334_/a_27_7# _334_/a_543_7# -0.00936f
C12876 _334_/a_193_7# _334_/a_761_249# -0.0157f
C12877 _337_/a_543_7# _194_/A 1.57e-21
C12878 _327_/a_193_7# _331_/CLK 0.582f
C12879 _255_/B _271_/A 1.13e-19
C12880 _321_/a_761_249# _321_/Q 0.022f
C12881 _208_/a_78_159# _207_/X 0.0112f
C12882 _329_/a_27_7# _328_/D 4.4e-21
C12883 repeater43/X _304_/a_306_329# 1.35e-19
C12884 _248_/B _314_/D 0.0377f
C12885 _338_/a_27_7# _337_/a_1283_n19# 1.06e-19
C12886 _338_/a_1283_n19# _337_/a_27_7# 2.16e-20
C12887 _338_/a_543_7# _337_/a_193_7# 1.13e-20
C12888 _338_/a_761_249# _337_/a_761_249# 4.46e-20
C12889 _338_/a_193_7# _337_/a_543_7# 4.67e-20
C12890 _273_/A _320_/Q 1.61e-20
C12891 _234_/a_109_257# VPWR -6.83e-19
C12892 _326_/a_193_7# _331_/CLK 0.0134f
C12893 _326_/a_27_7# _316_/D 3.75e-21
C12894 _292_/A _173_/a_226_7# 2.35e-21
C12895 _181_/X _207_/C 1.26e-19
C12896 _314_/a_27_7# _314_/a_543_7# -0.00482f
C12897 _311_/a_27_7# _310_/a_761_249# 1.1e-21
C12898 _311_/a_193_7# _310_/a_193_7# 2.17e-21
C12899 _311_/a_761_249# _310_/a_27_7# 4.52e-22
C12900 _321_/a_27_7# VPWR 0.0554f
C12901 _327_/a_193_7# _273_/A 1.83e-20
C12902 _258_/S trim[4] 0.00517f
C12903 _341_/Q _298_/B 0.868f
C12904 _165_/a_215_7# _346_/SET_B 3.3e-19
C12905 _325_/a_193_7# _223_/a_93_n19# 6.59e-20
C12906 _341_/a_805_7# _341_/D 0.00213f
C12907 _326_/a_193_7# _273_/A 3.25e-20
C12908 _242_/A _279_/A 0.0106f
C12909 _321_/a_27_7# _318_/a_543_7# 3.23e-21
C12910 rstn VPWR 1.48f
C12911 _232_/X _221_/a_93_n19# 0.0011f
C12912 _164_/A _160_/a_27_7# 1.12e-20
C12913 _281_/Y _181_/a_27_7# 1.21e-19
C12914 _332_/a_805_7# _333_/Q 5.85e-19
C12915 _340_/a_761_249# _337_/a_1283_n19# 0.00151f
C12916 _340_/a_193_7# _337_/a_1108_7# 9.56e-19
C12917 _340_/a_1108_7# _337_/a_193_7# 9.56e-19
C12918 _340_/a_1283_n19# _337_/a_761_249# 0.00151f
C12919 _210_/a_307_257# VGND 2.3e-20
C12920 _254_/A _196_/A 0.0101f
C12921 _338_/a_639_7# _346_/SET_B 0.00231f
C12922 _338_/a_448_7# _338_/Q 8.49e-21
C12923 _238_/B _319_/a_761_249# 0.00145f
C12924 _317_/D _286_/Y 0.0209f
C12925 _244_/B sample 2.81e-19
C12926 _310_/a_1283_n19# VGND 0.0165f
C12927 _310_/a_448_7# VPWR 0.00447f
C12928 _198_/a_584_7# _284_/A 4.53e-19
C12929 _319_/D VGND 0.129f
C12930 input4/X _332_/a_1283_n19# 8.9e-20
C12931 repeater43/X _332_/a_761_249# 8.17e-19
C12932 _306_/X _260_/A 4.3e-21
C12933 _344_/a_1140_373# _344_/Q 5.77e-19
C12934 _344_/a_381_7# _344_/D 0.016f
C12935 _343_/CLK _316_/a_27_7# 2.23e-21
C12936 _286_/B _191_/B 0.224f
C12937 output21/a_27_7# _331_/a_1108_7# 8.79e-20
C12938 _294_/A _309_/a_805_7# 0.0021f
C12939 _343_/Q _207_/C 2.67e-20
C12940 _298_/C _206_/A 0.0702f
C12941 _306_/S _311_/D 1.61e-20
C12942 _258_/a_76_159# _193_/Y 1.86e-19
C12943 _258_/a_505_n19# _306_/S 0.0407f
C12944 _190_/a_27_7# _333_/Q 4.3e-21
C12945 output31/a_27_7# VGND 0.0663f
C12946 _157_/A _147_/Y 2.2e-21
C12947 _340_/a_1217_7# _346_/SET_B -5.4e-19
C12948 _182_/X _225_/X 0.0278f
C12949 _196_/A _226_/X 4.99e-20
C12950 _181_/X _150_/C 0.303f
C12951 _283_/A _335_/a_1283_n19# 3.8e-20
C12952 _307_/X _182_/X 6.6e-20
C12953 output10/a_27_7# _277_/Y 0.0302f
C12954 _323_/D sample 5.52e-19
C12955 _225_/a_59_35# VPWR 0.00688f
C12956 _332_/a_448_7# _206_/A 1.09e-21
C12957 _332_/a_1283_n19# _207_/C 0.00628f
C12958 _339_/a_193_7# _338_/a_543_7# 7.48e-19
C12959 _339_/a_543_7# _338_/a_193_7# 1.16e-19
C12960 _339_/a_1283_n19# _338_/a_27_7# 5.53e-19
C12961 _344_/a_27_7# _165_/X 5.49e-21
C12962 _344_/a_193_7# _167_/X 1.71e-21
C12963 _256_/a_80_n19# _192_/B 0.0161f
C12964 _198_/a_93_n19# _340_/Q 0.0219f
C12965 _198_/a_250_257# _194_/X 0.00127f
C12966 _328_/a_1283_n19# _319_/a_193_7# 1.81e-19
C12967 _328_/a_1108_7# _319_/a_27_7# 0.00118f
C12968 _188_/S _306_/S 0.00545f
C12969 _335_/a_543_7# _205_/a_297_7# 1.89e-20
C12970 ctln[6] _211_/a_373_7# 4.17e-20
C12971 _215_/A _227_/A 0.0121f
C12972 _271_/A _325_/Q 0.0731f
C12973 _342_/a_1108_7# _228_/A 9.26e-22
C12974 _292_/A _158_/Y 0.646f
C12975 _243_/a_199_7# VPWR -2.77e-19
C12976 _183_/a_1241_257# _162_/X 3.74e-19
C12977 _267_/B _312_/Q 0.00386f
C12978 _327_/a_639_7# _346_/SET_B 0.00386f
C12979 result[1] _248_/B 2.84e-20
C12980 _325_/a_27_7# _304_/a_79_n19# 1.92e-20
C12981 _346_/a_193_7# _346_/a_1602_7# -4.26e-19
C12982 output22/a_27_7# _343_/CLK 0.00601f
C12983 repeater43/X _341_/a_1108_7# -0.0113f
C12984 _271_/A _298_/a_27_7# 0.00947f
C12985 _158_/Y _160_/A 0.112f
C12986 _165_/a_292_257# _345_/Q 4.74e-19
C12987 _172_/A _167_/X 4.18e-19
C12988 _340_/a_448_7# _339_/a_27_7# 1.27e-20
C12989 _340_/a_543_7# _339_/a_543_7# 8.59e-19
C12990 _340_/a_27_7# _339_/a_448_7# 5.09e-21
C12991 _226_/X _298_/X 7.63e-21
C12992 _343_/a_1217_7# _175_/Y 6.01e-19
C12993 _242_/a_109_257# _318_/D 8.83e-19
C12994 _342_/a_639_7# sample 3.59e-19
C12995 _163_/a_78_159# _163_/a_292_257# -1.09e-21
C12996 _164_/Y _162_/a_27_7# 4.17e-19
C12997 _190_/A _295_/a_306_7# 4.18e-19
C12998 _242_/A _318_/a_1270_373# 1.12e-19
C12999 _254_/A _347_/a_1283_n19# 0.00218f
C13000 _315_/a_543_7# _315_/D 1.98e-19
C13001 _320_/a_448_7# _328_/Q 8.27e-22
C13002 _318_/Q result[4] 0.031f
C13003 _308_/a_76_159# _209_/X 5.13e-21
C13004 _329_/a_639_7# _330_/D 0.00115f
C13005 _294_/A _311_/D 1.18e-20
C13006 _343_/Q _150_/C 3.81e-20
C13007 _298_/C _147_/A 0.134f
C13008 _294_/A _258_/a_505_n19# 5.65e-21
C13009 _336_/a_1283_n19# VPWR 0.00128f
C13010 _324_/a_761_249# _227_/A 0.0084f
C13011 _336_/a_761_249# VGND 0.00203f
C13012 _328_/a_1270_373# _346_/SET_B -2.06e-19
C13013 _326_/a_1462_7# _248_/A 3.6e-19
C13014 _331_/Q _280_/a_68_257# 3.23e-20
C13015 _271_/A _321_/a_1108_7# 0.00155f
C13016 _315_/D _314_/a_27_7# 0.192f
C13017 _332_/Q _333_/Q 0.324f
C13018 _149_/A _298_/C 0.00954f
C13019 _207_/X _190_/A 5.09e-19
C13020 _260_/A _147_/Y 0.017f
C13021 trimb[0] VPWR 0.249f
C13022 _260_/a_27_257# VGND -3.01e-19
C13023 output21/a_27_7# clkbuf_0_clk/X 1.38e-19
C13024 _227_/A _304_/X 0.00256f
C13025 ctln[5] input4/X 0.022f
C13026 repeater43/X _316_/a_448_7# -1.93e-19
C13027 _300_/a_301_257# _347_/Q 0.0114f
C13028 _279_/Y repeater43/X 1.41e-21
C13029 _300_/a_383_7# _299_/X 0.0144f
C13030 _321_/a_639_7# VGND -0.00169f
C13031 _321_/a_1217_7# VPWR 1.35e-19
C13032 _259_/a_113_257# _337_/Q 9.64e-21
C13033 _216_/X _212_/X 0.248f
C13034 rstn _335_/a_1108_7# 0.0502f
C13035 _286_/B _337_/Q 0.00189f
C13036 _338_/a_805_7# _343_/CLK 4.51e-20
C13037 _341_/a_27_7# _145_/A 3.41e-20
C13038 _329_/a_543_7# _232_/X 1.58e-20
C13039 _329_/Q _212_/X 0.111f
C13040 _320_/Q _217_/X 0.00343f
C13041 _291_/a_39_257# VGND 0.0214f
C13042 _340_/a_27_7# _337_/D 4.29e-21
C13043 _267_/A _312_/a_448_7# 5.68e-19
C13044 _327_/a_543_7# _327_/Q 0.00136f
C13045 _327_/a_761_249# _212_/X 0.00603f
C13046 _327_/a_193_7# _217_/X 0.00609f
C13047 _215_/A _347_/Q 4.35e-21
C13048 clkbuf_2_0_0_clk/a_75_172# VPWR 0.0805f
C13049 _319_/a_761_249# _331_/CLK 2.84e-21
C13050 _326_/a_1108_7# repeater43/X 0.0193f
C13051 _277_/Y _347_/Q 2.82e-20
C13052 _338_/D _338_/Q 0.0301f
C13053 _326_/a_27_7# _331_/a_27_7# 1.73e-19
C13054 _207_/C _204_/a_27_7# 0.0354f
C13055 _208_/a_215_7# _207_/C 3.36e-19
C13056 _281_/A _330_/a_448_7# 2.84e-19
C13057 _326_/a_193_7# _217_/X 0.547f
C13058 _310_/D VPWR 0.966f
C13059 _199_/a_346_7# VGND 3.06e-19
C13060 result[0] repeater43/X 0.00156f
C13061 _281_/Y _330_/a_543_7# 1.4e-19
C13062 _185_/A _323_/a_805_7# 6.97e-19
C13063 _306_/X _340_/Q 1.61e-19
C13064 _313_/Q _306_/S 0.65f
C13065 _342_/a_27_7# _269_/A 0.0149f
C13066 _334_/Q _208_/a_292_257# 3.84e-19
C13067 _300_/Y _227_/A 7.62e-21
C13068 _328_/a_193_7# _212_/X 0.21f
C13069 _328_/a_27_7# _217_/X 0.0176f
C13070 _302_/a_227_7# _347_/a_193_7# 6.03e-20
C13071 _183_/a_471_7# _181_/X 0.0113f
C13072 _344_/a_193_7# _301_/a_51_257# 3.84e-20
C13073 _344_/a_27_7# _301_/a_245_257# 5.17e-21
C13074 _346_/a_1140_373# _346_/SET_B 3.25e-19
C13075 clkbuf_0_clk/X _196_/A 0.00375f
C13076 _325_/a_651_373# _181_/X 0.00436f
C13077 _271_/A _326_/Q 0.00806f
C13078 _188_/S _283_/A 0.226f
C13079 _319_/Q _330_/a_1283_n19# 1.76e-20
C13080 result[5] _321_/a_543_7# 6.66e-22
C13081 _300_/a_301_257# _297_/B 0.00117f
C13082 _300_/Y _314_/a_1108_7# 3.56e-36
C13083 _332_/D _206_/A 0.0165f
C13084 _290_/A _312_/a_27_7# 4.75e-21
C13085 _279_/Y _191_/B 2.32e-19
C13086 _340_/CLK _313_/a_543_7# 4.44e-20
C13087 _197_/X _340_/D 3.79e-19
C13088 input4/X _334_/a_448_7# 0.0012f
C13089 repeater43/X _334_/a_1283_n19# 0.0386f
C13090 _309_/a_27_7# _310_/D 2.82e-20
C13091 trim[0] clkc 0.0891f
C13092 _326_/a_27_7# _217_/a_27_7# 0.00236f
C13093 _252_/a_27_7# _228_/A 5.73e-20
C13094 result[1] _315_/a_27_7# 0.00108f
C13095 _259_/a_113_257# _339_/Q 2.22e-19
C13096 _157_/A _304_/a_79_n19# 7.62e-21
C13097 _299_/X _346_/D 0.0684f
C13098 _342_/a_27_7# _343_/D 5.2e-20
C13099 _342_/a_761_249# _185_/A 3.38e-19
C13100 _172_/A _301_/a_51_257# 1.65e-19
C13101 _149_/A _229_/a_489_373# 5.22e-19
C13102 _325_/a_193_7# _216_/X 1.86e-20
C13103 output10/a_27_7# VGND 0.108f
C13104 _212_/a_27_7# _283_/A 3.7e-21
C13105 _335_/Q _153_/B 0.0255f
C13106 _257_/a_222_53# _305_/a_505_n19# 5.6e-19
C13107 clkbuf_1_0_0_clk/a_75_172# _330_/a_27_7# 3.3e-20
C13108 clkbuf_2_2_0_clk/a_75_172# _346_/SET_B 5.5e-20
C13109 _309_/a_651_373# _265_/B 9.07e-20
C13110 _271_/Y input3/a_27_7# 4.84e-20
C13111 _345_/a_27_7# _160_/X 4.94e-19
C13112 _160_/a_27_7# _160_/A 0.0531f
C13113 _337_/a_27_7# _337_/a_543_7# -0.00482f
C13114 _337_/a_193_7# _337_/a_761_249# -0.0052f
C13115 _344_/a_1032_373# _297_/Y 0.116f
C13116 _286_/B _202_/a_256_7# 8.41e-20
C13117 _215_/A _297_/B 0.00553f
C13118 _161_/Y comp 4.04e-20
C13119 input4/X _346_/SET_B 1.32e-19
C13120 _340_/a_27_7# _339_/D 0.0133f
C13121 _334_/a_448_7# _207_/C 0.0248f
C13122 _164_/A _267_/A 0.101f
C13123 _277_/Y _297_/B 0.0603f
C13124 _308_/a_505_n19# _153_/A 1.27e-19
C13125 _188_/S _248_/B 2.32e-20
C13126 _315_/a_805_7# VPWR 4.17e-19
C13127 _308_/S _209_/X 2.1e-19
C13128 _304_/S _347_/D 2.53e-19
C13129 _311_/Q clkc 1.69e-20
C13130 _324_/a_1283_n19# _315_/D 1.79e-20
C13131 _196_/A input1/X 0.0158f
C13132 trimb[3] VPWR 0.123f
C13133 _227_/A VGND 4f
C13134 _294_/A _313_/Q 0.00411f
C13135 _320_/a_1108_7# _319_/D 2.15e-19
C13136 _274_/a_121_257# _327_/Q 5.18e-20
C13137 _324_/a_27_7# VPWR 0.0665f
C13138 _342_/a_193_7# _342_/Q 0.0022f
C13139 _321_/Q _304_/X 0.013f
C13140 _346_/SET_B _345_/Q 0.0628f
C13141 _346_/a_1182_221# clkbuf_2_3_0_clk/A 0.0124f
C13142 _318_/a_761_249# _242_/B 1.03e-19
C13143 _318_/a_27_7# _318_/D 0.052f
C13144 _326_/a_27_7# _325_/a_543_7# 2.16e-20
C13145 _315_/D _314_/a_1217_7# 4.27e-19
C13146 _334_/a_1270_373# _334_/D 2.49e-19
C13147 _334_/a_1283_n19# _334_/Q 0.00215f
C13148 _273_/A _158_/Y 0.147f
C13149 _314_/a_1108_7# VGND 0.0143f
C13150 _314_/a_651_373# VPWR 0.00303f
C13151 _281_/Y _331_/Q 0.0118f
C13152 _346_/SET_B _319_/a_805_7# 5.85e-19
C13153 _346_/SET_B _313_/a_1283_n19# -0.0135f
C13154 _269_/A _317_/D 0.00769f
C13155 _324_/a_761_249# _297_/B 3.04e-20
C13156 _340_/Q _147_/Y 2.75e-19
C13157 _338_/a_1108_7# _337_/Q 1.73e-21
C13158 _338_/D _337_/a_639_7# 1.98e-20
C13159 _346_/SET_B _337_/a_1270_373# 2.28e-19
C13160 clk _332_/a_1108_7# 0.0538f
C13161 _157_/A _347_/a_193_7# 0.0123f
C13162 repeater43/X _316_/D 0.0108f
C13163 _324_/a_448_7# _324_/D 0.0145f
C13164 _347_/Q _300_/Y 0.0024f
C13165 _314_/a_1283_n19# _314_/Q 0.00451f
C13166 _271_/A _154_/A 9.8e-19
C13167 _311_/D _310_/a_651_373# 1.88e-19
C13168 _338_/Q _343_/CLK 0.0162f
C13169 _322_/a_805_7# _269_/A 5.87e-19
C13170 _293_/a_39_257# _336_/a_27_7# 2.94e-21
C13171 _334_/a_543_7# _323_/Q 9.34e-19
C13172 _279_/Y _302_/a_323_257# 2.23e-20
C13173 _324_/Q _268_/a_121_257# 8.47e-19
C13174 _270_/a_121_257# _244_/B 7.87e-21
C13175 _267_/B _340_/CLK 0.0122f
C13176 input1/X _298_/X 1.07e-21
C13177 _345_/a_193_7# VPWR 0.0467f
C13178 _256_/a_80_n19# _260_/A 7.66e-19
C13179 _339_/a_651_373# _340_/CLK 0.00137f
C13180 _153_/a_403_257# _153_/B 3.09e-19
C13181 _266_/a_113_257# VPWR 0.0725f
C13182 _340_/a_651_373# _337_/Q 3.33e-20
C13183 _267_/A _312_/D 0.00661f
C13184 cal _343_/Q 0.0783f
C13185 _327_/a_1462_7# _217_/X 3.46e-19
C13186 _329_/D _331_/Q 1.01e-19
C13187 _345_/a_476_7# _297_/B 4.08e-19
C13188 repeater43/a_27_7# repeater43/X 0.134f
C13189 _196_/A _286_/Y 2.88e-20
C13190 _165_/X _147_/Y 0.00848f
C13191 _279_/Y _337_/Q 3.88e-20
C13192 _341_/a_27_7# _324_/Q 2.41e-21
C13193 repeater43/X _222_/a_250_257# 0.00141f
C13194 _149_/A _334_/a_1270_373# 5.17e-21
C13195 output24/a_27_7# _318_/Q 2.1e-19
C13196 _317_/Q output25/a_27_7# 5.45e-20
C13197 _277_/A _320_/a_1283_n19# 3.12e-19
C13198 _177_/a_27_7# _228_/A 6.55e-19
C13199 _184_/a_76_159# _298_/B 2.08e-20
C13200 _255_/X _254_/B 8.74e-20
C13201 _306_/S _333_/a_1283_n19# 3.27e-20
C13202 _257_/a_448_7# _254_/B 6.68e-19
C13203 _245_/a_113_257# VPWR 0.0496f
C13204 _298_/C _150_/a_27_7# 0.0122f
C13205 input4/X _206_/A 1.22e-19
C13206 _347_/Q VGND 0.675f
C13207 _303_/A _347_/a_543_7# 6.46e-20
C13208 _196_/A _250_/a_215_7# 7.2e-19
C13209 _260_/A _347_/a_193_7# 5.99e-22
C13210 _322_/a_193_7# _322_/D 0.00526f
C13211 _336_/Q _153_/B 5.48e-21
C13212 _322_/a_1283_n19# _321_/a_543_7# 2.2e-19
C13213 _173_/a_226_257# _172_/Y 1.82e-19
C13214 _298_/X _286_/Y 4e-19
C13215 _318_/a_543_7# _245_/a_113_257# 4.47e-21
C13216 _300_/Y _297_/B 0.0176f
C13217 _232_/a_27_7# _326_/Q 6.5e-20
C13218 _232_/X _243_/a_113_257# 2.04e-21
C13219 _255_/B _231_/a_79_n19# 0.121f
C13220 _339_/a_1270_373# _346_/SET_B 2.19e-19
C13221 _275_/Y _215_/A 0.0131f
C13222 _316_/Q _318_/D 9.93e-20
C13223 _188_/a_76_159# _150_/C 9e-19
C13224 input4/X _334_/D 9.55e-19
C13225 _188_/a_505_n19# _307_/X 0.00209f
C13226 _258_/a_505_n19# _336_/a_1108_7# 4.77e-19
C13227 _246_/B _217_/A 0.652f
C13228 output7/a_27_7# input4/X 1.06e-19
C13229 _277_/Y _275_/Y 0.0526f
C13230 _288_/A _290_/A 1.1e-19
C13231 _192_/B _333_/Q 0.212f
C13232 _206_/A _207_/C 0.0993f
C13233 _297_/B _220_/a_93_n19# 5.9e-21
C13234 _324_/Q _316_/a_193_7# 1.37e-19
C13235 _250_/X _162_/X 0.00609f
C13236 _313_/a_193_7# _313_/a_1108_7# -0.00656f
C13237 _313_/a_27_7# _313_/a_448_7# -0.0068f
C13238 _260_/B _157_/A 0.00115f
C13239 _290_/A _162_/X 0.00612f
C13240 _290_/A _287_/a_39_257# 0.00266f
C13241 _286_/B _336_/D 0.158f
C13242 _321_/Q VGND 1.92f
C13243 _181_/X _284_/A 0.0553f
C13244 _145_/A _180_/a_111_257# 7.69e-19
C13245 input2/a_27_7# output40/a_27_7# 2.3e-22
C13246 repeater43/a_27_7# _191_/B 1.23e-19
C13247 _334_/D _207_/C 0.109f
C13248 _198_/a_250_257# _336_/a_543_7# 3.23e-20
C13249 _317_/a_1283_n19# _248_/A 1.59e-19
C13250 _316_/Q _217_/A 4.94e-20
C13251 output7/a_27_7# _207_/C 4.36e-20
C13252 _327_/a_448_7# clkbuf_0_clk/X 1.1e-19
C13253 _313_/Q _254_/Y 0.0101f
C13254 _279_/Y _339_/Q 4.06e-22
C13255 _339_/a_27_7# _339_/a_543_7# -0.0049f
C13256 _297_/a_27_257# _347_/a_1283_n19# 4.07e-19
C13257 _302_/a_77_159# _346_/SET_B 0.00195f
C13258 _269_/Y ctln[0] 0.0102f
C13259 _254_/A _313_/a_193_7# 0.00189f
C13260 _324_/a_1217_7# VPWR 6.8e-20
C13261 _324_/a_639_7# VGND -0.0012f
C13262 _315_/Q _146_/C 1.86e-20
C13263 _342_/a_1462_7# _342_/Q 1.6e-19
C13264 _317_/a_543_7# _316_/D 3.2e-20
C13265 _317_/a_1283_n19# _331_/CLK 2.74e-21
C13266 _338_/a_27_7# _195_/a_27_257# 0.0105f
C13267 _273_/A _160_/a_27_7# 1.22e-19
C13268 cal _229_/a_76_159# 0.00233f
C13269 _297_/B VGND 1.22f
C13270 repeater42/a_27_7# _330_/Q 4.58e-20
C13271 _183_/a_553_257# _180_/a_29_13# 1.57e-20
C13272 _179_/a_27_7# _209_/a_27_257# 0.00103f
C13273 _318_/a_193_7# VGND 0.00707f
C13274 _318_/a_543_7# VPWR 0.00802f
C13275 _341_/a_27_7# _228_/A 1.09e-19
C13276 _343_/a_805_7# VPWR 3.45e-19
C13277 _343_/a_1270_373# VGND 4.69e-20
C13278 _346_/a_27_7# _276_/a_68_257# 2.72e-22
C13279 _175_/Y _244_/B 0.00256f
C13280 _244_/B _243_/a_113_257# 0.00203f
C13281 output8/a_27_7# ctln[2] 0.0196f
C13282 _272_/a_121_257# _246_/B 8.56e-19
C13283 clk _340_/CLK 7.12e-20
C13284 _273_/A _317_/a_1283_n19# 3.43e-20
C13285 _220_/a_584_7# _279_/A 0.00103f
C13286 ctlp[6] VPWR 0.0877f
C13287 _194_/X _312_/D 7.91e-20
C13288 _345_/a_476_7# _275_/Y 0.00223f
C13289 _147_/A _345_/Q 4.49e-20
C13290 _236_/B _331_/a_1108_7# 1.53e-19
C13291 _331_/CLK _331_/a_651_373# 9.87e-19
C13292 result[7] _331_/CLK 1.79e-19
C13293 _231_/a_512_7# _283_/A 0.00118f
C13294 _318_/a_193_7# _318_/a_1108_7# -0.0069f
C13295 _150_/C _206_/A 9.79e-21
C13296 _309_/a_27_7# VPWR 0.0439f
C13297 cal _204_/a_27_7# 3.26e-19
C13298 _313_/a_1283_n19# _147_/A 0.0984f
C13299 _341_/a_448_7# _286_/Y 0.0148f
C13300 _279_/Y _303_/A 0.085f
C13301 _305_/a_505_n19# _336_/Q 6.6e-20
C13302 _305_/a_76_159# _225_/B 0.0103f
C13303 _345_/a_1140_373# VGND 8.85e-20
C13304 _345_/a_796_7# VPWR 3.95e-19
C13305 _260_/B _260_/A 0.108f
C13306 _339_/D _332_/D 7.3e-21
C13307 _149_/A _207_/C 2.04e-20
C13308 _323_/D _175_/Y 0.00137f
C13309 _162_/A _344_/Q 0.00469f
C13310 _307_/a_218_334# _191_/B 0.00114f
C13311 _292_/A _267_/A 0.00956f
C13312 _336_/a_193_7# _254_/B 2.84e-19
C13313 output27/a_27_7# _321_/Q 2.06e-19
C13314 _283_/A _330_/a_1270_373# 6.3e-20
C13315 _325_/Q _231_/a_79_n19# 1.42e-22
C13316 clk _334_/a_651_373# 0.00152f
C13317 _172_/A _341_/Q 0.00475f
C13318 _194_/a_27_7# _311_/D 3.72e-20
C13319 repeater43/X _331_/a_27_7# 0.0179f
C13320 _327_/a_27_7# _281_/A 3.74e-20
C13321 _160_/A _267_/A 1.39e-19
C13322 _283_/A _333_/a_1283_n19# 0.0595f
C13323 _316_/a_193_7# _228_/A 1.37e-21
C13324 output19/a_27_7# clkbuf_2_1_0_clk/A 0.0517f
C13325 _258_/a_76_159# _215_/A 1.22e-20
C13326 _167_/a_27_257# _162_/X 0.0156f
C13327 _255_/a_30_13# _286_/B 0.0674f
C13328 _277_/A _320_/D 0.0643f
C13329 _307_/X _304_/S 7.53e-20
C13330 _326_/a_27_7# _281_/A 5.81e-20
C13331 _310_/D _171_/a_215_7# 3.85e-20
C13332 _188_/S _298_/B 0.328f
C13333 _327_/Q _212_/X 0.244f
C13334 _309_/a_448_7# _309_/Q 2.82e-21
C13335 _301_/X _347_/D 4.23e-21
C13336 _308_/a_218_334# VGND 9.48e-19
C13337 _308_/a_218_7# VPWR -4.9e-19
C13338 _283_/A _223_/a_93_n19# 1.57e-21
C13339 _154_/a_27_7# _153_/A 2.86e-19
C13340 _343_/a_193_7# _323_/a_543_7# 3.1e-22
C13341 _343_/a_761_249# _323_/a_761_249# 8.24e-21
C13342 _343_/a_1283_n19# _323_/a_27_7# 8.85e-19
C13343 _306_/a_76_159# VPWR 0.0202f
C13344 _294_/Y trimb[4] 0.0206f
C13345 _255_/B _162_/X 0.746f
C13346 _294_/Y trim[1] 0.0015f
C13347 _329_/a_27_7# _181_/X 1.06e-20
C13348 _147_/A _150_/C 0.234f
C13349 _311_/a_651_373# VPWR 0.0127f
C13350 _311_/a_1108_7# VGND 0.00393f
C13351 _263_/a_109_257# _310_/a_193_7# 1.4e-19
C13352 cal _334_/a_448_7# 3.25e-19
C13353 _306_/X _336_/a_1283_n19# 5.03e-21
C13354 _313_/Q _336_/a_1108_7# 9.89e-19
C13355 _285_/A _345_/a_27_7# 1.52e-20
C13356 repeater43/X _217_/a_27_7# 0.00152f
C13357 _179_/a_27_7# _153_/A 4.29e-19
C13358 _149_/A _150_/C 0.388f
C13359 _346_/SET_B _202_/a_93_n19# 0.0174f
C13360 repeater43/X _145_/A 0.00397f
C13361 repeater43/X output28/a_27_7# 0.00142f
C13362 _292_/Y ctlp[3] 6.43e-19
C13363 _345_/a_193_7# _344_/a_27_7# 6.66e-21
C13364 _216_/X _221_/a_256_7# 7.53e-19
C13365 _345_/a_27_7# _344_/a_193_7# 0.00143f
C13366 _337_/a_1283_n19# _337_/Q 0.037f
C13367 _288_/A _310_/a_27_7# 1.04e-20
C13368 _335_/a_543_7# VGND 0.00168f
C13369 _335_/a_1108_7# VPWR -0.0111f
C13370 _184_/a_505_n19# VPWR 0.0549f
C13371 input1/X _338_/D 2.82e-19
C13372 ctln[3] VPWR 0.194f
C13373 cal _346_/SET_B 0.00727f
C13374 _275_/Y VGND 0.663f
C13375 _232_/A _223_/a_250_257# 0.00141f
C13376 _276_/a_68_257# _275_/A 7.47e-20
C13377 _341_/Q _244_/B 6.65e-19
C13378 _193_/Y _194_/A 0.165f
C13379 _225_/B _203_/a_303_7# 0.00208f
C13380 _250_/X _298_/C 9.18e-22
C13381 output31/a_27_7# output32/a_27_7# 0.00185f
C13382 _254_/A _313_/a_1462_7# 2.44e-19
C13383 _340_/a_651_373# _336_/D 2.62e-20
C13384 _326_/a_27_7# _216_/A 9.4e-19
C13385 _212_/a_27_7# _242_/B 1.42e-19
C13386 _338_/a_193_7# _193_/Y 0.00995f
C13387 _338_/a_543_7# _340_/Q 0.00308f
C13388 _338_/a_1283_n19# _194_/X 0.00398f
C13389 _331_/Q _242_/A 7.91e-20
C13390 _345_/a_27_7# _172_/A 3.2e-19
C13391 _279_/Y _336_/D 3.21e-20
C13392 _325_/a_543_7# repeater43/X 0.00182f
C13393 _209_/X _333_/a_193_7# 5.03e-19
C13394 ctlp[7] clkbuf_1_0_0_clk/a_75_172# 2.23e-19
C13395 _324_/Q _180_/a_111_257# 1.5e-19
C13396 _258_/S _193_/Y 9.46e-20
C13397 _318_/a_1462_7# VGND -8.93e-19
C13398 _218_/a_250_257# _330_/D 0.00226f
C13399 _302_/a_77_159# _147_/A 0.0171f
C13400 _325_/a_27_7# _212_/X 3.45e-19
C13401 _325_/a_193_7# _327_/Q 3.06e-20
C13402 _275_/Y _309_/a_761_249# 0.00126f
C13403 _164_/Y clkc 6.6e-20
C13404 _277_/Y _161_/Y 8.73e-20
C13405 _320_/a_193_7# _220_/a_93_n19# 4.59e-20
C13406 _309_/a_1217_7# VPWR 1.06e-19
C13407 _309_/a_639_7# VGND -0.00169f
C13408 _341_/D _286_/Y 0.624f
C13409 _340_/a_193_7# _340_/D 0.0613f
C13410 _340_/a_543_7# _193_/Y 0.00725f
C13411 _340_/a_448_7# _194_/X 2.59e-20
C13412 _340_/a_1108_7# _340_/Q 0.0483f
C13413 clkbuf_2_1_0_clk/A _197_/X 0.0116f
C13414 _185_/A _182_/X 0.00619f
C13415 _258_/a_76_159# _300_/Y 1.55e-20
C13416 _269_/A _298_/X 0.0125f
C13417 _336_/a_1283_n19# _147_/Y 0.0665f
C13418 _145_/A _191_/B 0.0827f
C13419 _219_/a_346_7# _346_/SET_B 0.00103f
C13420 _163_/a_78_159# _344_/Q 1.64e-19
C13421 _322_/D _331_/Q 2.48e-20
C13422 _325_/Q _162_/X 1.93e-20
C13423 _164_/A _310_/a_1108_7# 5.78e-20
C13424 _290_/A _165_/a_215_7# 1.7e-19
C13425 _339_/a_1283_n19# _337_/Q 2.8e-19
C13426 _321_/a_651_373# _322_/Q 5.88e-19
C13427 _346_/a_27_7# _346_/Q 2.16e-19
C13428 _307_/a_76_159# _157_/A 2.58e-21
C13429 repeater43/X _331_/a_1217_7# 2.12e-19
C13430 _331_/a_27_7# _331_/a_448_7# -0.00972f
C13431 _183_/a_27_7# _304_/S 1.31e-19
C13432 clkbuf_0_clk/a_110_7# _157_/a_27_7# 4.24e-21
C13433 _248_/A sample 0.00558f
C13434 _255_/X _196_/A 0.085f
C13435 _342_/Q _181_/X 0.356f
C13436 _320_/a_543_7# VPWR 0.0141f
C13437 _320_/a_193_7# VGND 0.0484f
C13438 _316_/a_27_7# _247_/a_113_257# 7.96e-19
C13439 _257_/a_448_7# _196_/A 2.06e-19
C13440 _185_/A valid 4.65e-19
C13441 _343_/D _298_/X 0.00717f
C13442 _323_/a_1108_7# VPWR 0.00959f
C13443 _323_/a_543_7# VGND 0.0187f
C13444 _344_/a_27_7# VPWR -0.207f
C13445 cal _206_/A 0.0112f
C13446 _312_/Q _297_/Y 0.00285f
C13447 _320_/a_1108_7# _297_/B 0.0653f
C13448 _273_/A _267_/A 0.00869f
C13449 cal _337_/a_448_7# 3.08e-19
C13450 _275_/Y _311_/a_639_7# 3.45e-19
C13451 _318_/Q _227_/A 1.42e-20
C13452 _207_/a_27_7# _332_/Q 0.0223f
C13453 _183_/a_1241_257# _150_/C 0.00746f
C13454 _207_/X _207_/a_109_7# 3.57e-19
C13455 _281_/Y _340_/CLK 2.94e-19
C13456 _344_/a_652_n19# _297_/B 1.04e-20
C13457 clk _225_/X 0.00683f
C13458 _258_/a_218_334# VPWR -0.00162f
C13459 _294_/A _162_/A 1.02e-19
C13460 _258_/a_76_159# VGND 0.00399f
C13461 ctln[4] _197_/X 4.53e-21
C13462 _281_/Y _347_/D 8.9e-21
C13463 clkbuf_2_1_0_clk/A _312_/a_193_7# 1.27e-20
C13464 input1/X _343_/CLK 9.52e-21
C13465 cal _334_/D 0.00133f
C13466 _325_/a_27_7# _325_/a_193_7# -0.294f
C13467 _143_/a_27_7# _286_/Y 1.9e-20
C13468 _183_/a_471_7# _149_/A 1.59e-19
C13469 _330_/Q _232_/X 0.706f
C13470 _342_/D _298_/A 1.07e-19
C13471 _248_/A _221_/a_93_n19# 3.61e-19
C13472 _346_/SET_B _284_/A 0.498f
C13473 _312_/Q _310_/a_193_7# 7.35e-19
C13474 _329_/a_1108_7# _216_/X 7.3e-19
C13475 _216_/X _327_/D 0.00591f
C13476 _172_/A _314_/D 3e-21
C13477 _342_/Q _343_/Q 1.01e-24
C13478 _248_/B _347_/a_27_7# 0.0163f
C13479 _255_/B _298_/C 0.233f
C13480 _211_/a_27_257# VPWR 0.102f
C13481 _328_/a_1270_373# _319_/Q 4.23e-19
C13482 _198_/a_93_n19# VPWR 0.0147f
C13483 _306_/S _190_/a_27_7# 0.0469f
C13484 _341_/a_448_7# _269_/A 0.00883f
C13485 _301_/X _304_/S 3.19e-20
C13486 cal _191_/a_109_257# 1.76e-19
C13487 _343_/a_651_373# _342_/a_27_7# 8.42e-21
C13488 _343_/a_543_7# _342_/a_1283_n19# 7.56e-20
C13489 _147_/A _202_/a_93_n19# 1.89e-19
C13490 _338_/a_761_249# _283_/A 1.01e-20
C13491 trim[4] _267_/A 0.0377f
C13492 _329_/a_1108_7# _329_/Q 7.5e-19
C13493 _339_/a_1283_n19# _339_/Q 0.0437f
C13494 _329_/a_193_7# _327_/a_448_7# 2.89e-20
C13495 _329_/a_1283_n19# _327_/a_543_7# 1.13e-19
C13496 _329_/a_1108_7# _327_/a_761_249# 6.9e-21
C13497 _329_/a_651_373# _327_/a_27_7# 1.75e-20
C13498 _327_/a_761_249# _327_/D 4.93e-19
C13499 repeater43/X _324_/Q 0.0362f
C13500 _273_/A _221_/a_93_n19# 0.0104f
C13501 output16/a_27_7# trimb[3] 0.0077f
C13502 ctlp[2] output39/a_27_7# 3.47e-19
C13503 _171_/a_215_7# VPWR 0.0012f
C13504 _171_/a_292_257# VGND -0.00136f
C13505 _289_/a_39_257# _310_/Q 7.21e-19
C13506 _333_/a_27_7# _154_/A 1.45e-19
C13507 _333_/a_761_249# _153_/A 4.85e-21
C13508 cal _147_/A 0.00325f
C13509 _210_/a_27_7# _333_/D 0.00489f
C13510 rstn _332_/a_27_7# 2.63e-20
C13511 _169_/B _162_/X 0.0457f
C13512 cal _149_/A 0.0446f
C13513 _343_/CLK _286_/Y 0.134f
C13514 _340_/a_1283_n19# _283_/A 6.76e-21
C13515 trim[0] _311_/a_1283_n19# 4.17e-19
C13516 _216_/X _283_/A 0.00113f
C13517 _275_/A _346_/Q 1.44e-20
C13518 _329_/a_27_7# _328_/a_448_7# 1.72e-21
C13519 _329_/a_1108_7# _328_/a_193_7# 5.75e-20
C13520 _328_/a_1108_7# _328_/Q 0.0372f
C13521 output28/a_27_7# result[6] 0.0143f
C13522 _162_/X _326_/Q 3.23e-22
C13523 _150_/C _150_/a_27_7# 0.015f
C13524 _182_/X _298_/a_109_7# 1.07e-19
C13525 result[2] _316_/a_27_7# 3.25e-19
C13526 _313_/Q _160_/X 1.44e-20
C13527 _196_/A _336_/a_193_7# 0.00227f
C13528 _286_/B _336_/a_761_249# 0.00228f
C13529 _177_/A _175_/Y 5.36e-20
C13530 _271_/A _322_/a_193_7# 6.04e-21
C13531 _185_/A _229_/a_226_7# 0.0247f
C13532 _322_/a_639_7# _321_/Q 6.39e-19
C13533 _306_/S _332_/Q 0.00333f
C13534 _161_/Y VGND 1.48f
C13535 output14/a_27_7# _322_/D 0.00495f
C13536 _286_/B _260_/a_27_257# 7.66e-20
C13537 _193_/Y _201_/a_27_7# 0.041f
C13538 _311_/a_1283_n19# _311_/Q 0.0224f
C13539 _326_/a_761_249# _283_/A 0.00183f
C13540 _318_/a_27_7# _317_/D 1.92e-20
C13541 _318_/a_761_249# _244_/B 6.44e-20
C13542 _226_/X output30/a_27_7# 5.29e-20
C13543 _322_/a_651_373# VPWR -0.00876f
C13544 _322_/a_1108_7# VGND 0.00173f
C13545 _216_/X _248_/B 0.456f
C13546 _313_/a_27_7# _336_/D 2.19e-22
C13547 _315_/a_761_249# _177_/a_27_7# 8.97e-20
C13548 _313_/a_761_249# _284_/A 0.0077f
C13549 _344_/a_652_n19# _275_/Y 4.46e-20
C13550 _320_/a_1462_7# VGND 2.24e-19
C13551 _346_/a_1182_221# _165_/X 0.00371f
C13552 _346_/a_1032_373# _167_/X 0.00957f
C13553 rstn _338_/a_543_7# 3.11e-20
C13554 repeater43/X _281_/A 0.0141f
C13555 _318_/Q _321_/Q 9.53e-20
C13556 _324_/Q _191_/B 0.00252f
C13557 _162_/X _314_/a_193_7# 1.63e-19
C13558 trim[2] _346_/SET_B 1.89e-19
C13559 _305_/a_439_7# VGND 2.02e-19
C13560 _344_/a_586_7# VPWR 0.00166f
C13561 trim[3] clkc 0.00318f
C13562 _329_/a_27_7# _346_/SET_B -8.5e-19
C13563 _227_/a_113_7# VPWR -6.72e-20
C13564 _298_/C _298_/a_27_7# 0.134f
C13565 input1/a_75_172# _337_/Q 1.89e-21
C13566 cal _337_/D 0.205f
C13567 _309_/a_761_249# _161_/Y 7.42e-22
C13568 _332_/a_1283_n19# _204_/Y 9.33e-20
C13569 _332_/a_1108_7# _335_/Q 3.19e-19
C13570 output25/a_27_7# VGND 0.101f
C13571 _254_/Y _340_/a_1283_n19# 1.49e-21
C13572 _343_/a_639_7# _323_/D 0.00108f
C13573 _306_/S _173_/a_489_373# 0.00324f
C13574 repeater43/X _228_/A 0.189f
C13575 _149_/a_27_7# _146_/C 1.56e-19
C13576 _243_/a_113_257# _325_/D 2.1e-20
C13577 _162_/X _170_/a_226_7# 0.00496f
C13578 _172_/A _184_/a_76_159# 0.00561f
C13579 _306_/X VPWR 0.102f
C13580 _156_/a_39_257# _284_/A 1.61e-19
C13581 _273_/A _167_/X 0.00913f
C13582 _344_/D _345_/D 2.97e-20
C13583 _168_/a_109_7# clkbuf_2_3_0_clk/A 0.0118f
C13584 _318_/Q _297_/B 2.33e-20
C13585 _337_/a_193_7# _306_/S 4.63e-20
C13586 _337_/a_761_249# _340_/Q 1.21e-20
C13587 _337_/a_27_7# _193_/Y 6.61e-20
C13588 _337_/a_543_7# _194_/X 0.00499f
C13589 _318_/Q _318_/a_193_7# 0.555f
C13590 ctln[5] input4/a_27_7# 9.98e-20
C13591 _335_/a_1283_n19# _335_/D 8.68e-20
C13592 _342_/a_1270_373# VPWR 5.14e-20
C13593 _342_/a_448_7# VGND -0.00503f
C13594 _292_/A _310_/a_1108_7# 0.00297f
C13595 repeater43/X _207_/a_181_7# 3.3e-19
C13596 _239_/a_199_7# _327_/Q 1.13e-20
C13597 _199_/a_584_7# _312_/D 1.25e-19
C13598 _346_/Q _345_/D 3.58e-20
C13599 _315_/Q _232_/A 6.58e-19
C13600 _337_/Q _174_/a_27_257# 7.57e-21
C13601 _297_/A _314_/a_448_7# 7.3e-22
C13602 _324_/Q _317_/a_543_7# 4.4e-21
C13603 _329_/a_543_7# _331_/CLK 0.00512f
C13604 _268_/a_39_257# _315_/a_543_7# 0.00965f
C13605 _341_/D _269_/A 0.0157f
C13606 ctln[6] _343_/CLK 0.0109f
C13607 _246_/B _317_/D 0.00881f
C13608 _343_/a_193_7# _342_/D 2.94e-21
C13609 _308_/a_505_n19# _254_/B 7.07e-21
C13610 _147_/A _284_/A 0.0501f
C13611 _319_/Q _319_/a_805_7# 5.13e-19
C13612 _189_/a_27_7# _332_/D 1.78e-20
C13613 _248_/a_109_257# VPWR -6.14e-19
C13614 _165_/X _319_/a_1283_n19# 1.22e-20
C13615 _254_/A _344_/D 3.64e-20
C13616 output16/a_27_7# VPWR 0.129f
C13617 repeater43/X _216_/A 0.0156f
C13618 _281_/Y _304_/S 0.00729f
C13619 _257_/a_222_53# _340_/CLK 0.00161f
C13620 _320_/a_27_7# _320_/a_448_7# -0.00297f
C13621 _312_/a_27_7# _311_/a_193_7# 1.75e-21
C13622 _312_/a_193_7# _311_/a_27_7# 9.49e-20
C13623 _276_/a_68_257# clkbuf_0_clk/X 0.0509f
C13624 _277_/Y _263_/B 0.202f
C13625 _326_/D _328_/Q 2.47e-21
C13626 _341_/a_193_7# _315_/a_193_7# 9.38e-19
C13627 _341_/a_27_7# _315_/a_761_249# 1.1e-21
C13628 _341_/a_761_249# _315_/a_27_7# 1.02e-21
C13629 result[1] _244_/B 2.06e-20
C13630 _254_/A _346_/Q 0.00719f
C13631 _316_/Q _317_/D 0.186f
C13632 _341_/a_193_7# _298_/A 0.169f
C13633 _332_/a_651_373# _153_/a_215_257# 0.00179f
C13634 _341_/Q _177_/A 0.35f
C13635 clkbuf_2_1_0_clk/A _299_/a_215_7# 0.00901f
C13636 _331_/D _246_/B 1.78e-21
C13637 _345_/a_27_7# _164_/A 0.00133f
C13638 input1/a_75_172# _339_/Q 2.4e-20
C13639 cal _339_/D 0.0237f
C13640 _246_/B _330_/a_193_7# 2.73e-20
C13641 _217_/X _221_/a_93_n19# 0.0106f
C13642 _290_/A _345_/Q 0.731f
C13643 _212_/X _221_/a_250_257# 0.0173f
C13644 _327_/Q _221_/a_256_7# 5.78e-19
C13645 _228_/A _191_/B 1.71e-20
C13646 _233_/a_199_7# VPWR -2.03e-19
C13647 _281_/Y _225_/X 1.43e-20
C13648 _236_/B _269_/A 0.00343f
C13649 _167_/a_109_7# _346_/SET_B 3.41e-21
C13650 _216_/A _313_/a_448_7# 0.0137f
C13651 _339_/D _197_/a_27_7# 4.87e-19
C13652 ctln[7] _335_/a_1270_373# 4.3e-19
C13653 _283_/A _332_/Q 0.0114f
C13654 _274_/a_39_257# _248_/B 1.48e-19
C13655 _286_/B _227_/A 0.231f
C13656 _340_/CLK _310_/a_193_7# 0.00163f
C13657 _147_/Y VPWR 1.05f
C13658 _339_/a_761_249# _340_/Q 0.00976f
C13659 _339_/a_27_7# _193_/Y 0.00719f
C13660 _339_/a_193_7# _306_/S 0.0142f
C13661 _285_/A _285_/Y 0.0967f
C13662 _328_/a_1283_n19# _319_/D 8.96e-19
C13663 _341_/Q _333_/D 1.04e-19
C13664 _312_/a_543_7# VGND 0.00807f
C13665 _312_/a_1108_7# VPWR 0.0135f
C13666 _283_/Y _153_/B 5.23e-20
C13667 _200_/a_93_n19# _199_/a_93_n19# 1.68e-19
C13668 _313_/Q _306_/a_505_n19# 2.53e-20
C13669 _196_/A _314_/a_1283_n19# 1.89e-19
C13670 clkbuf_0_clk/a_110_7# _267_/A 4.6e-19
C13671 _306_/X _306_/a_76_159# 8.81e-19
C13672 _335_/Q _204_/a_277_7# 0.00398f
C13673 _204_/Y _204_/a_27_7# 0.0414f
C13674 _270_/a_39_257# _316_/D 0.0601f
C13675 _208_/a_215_7# _204_/Y 2.18e-19
C13676 output26/a_27_7# result[6] 0.0026f
C13677 _316_/a_543_7# _315_/a_27_7# 1.63e-21
C13678 _316_/a_193_7# _315_/a_761_249# 6.73e-20
C13679 _316_/a_27_7# _315_/a_543_7# 2.89e-19
C13680 _316_/a_761_249# _315_/a_193_7# 1.99e-19
C13681 _346_/a_1032_373# clkbuf_1_1_0_clk/a_75_172# 4.22e-21
C13682 _231_/a_409_7# VGND -0.00137f
C13683 ctln[2] output33/a_27_7# 2.89e-20
C13684 clkbuf_2_3_0_clk/A _306_/S 0.0157f
C13685 _258_/a_505_n19# _172_/A 9.02e-20
C13686 _169_/Y _347_/a_1108_7# 2.33e-21
C13687 _330_/Q _330_/a_805_7# 2.22e-19
C13688 _219_/a_93_n19# clkbuf_0_clk/X 2.12e-20
C13689 _326_/a_1270_373# _242_/A 2.42e-19
C13690 _277_/A _238_/B 0.00478f
C13691 _186_/a_297_7# _308_/X 0.00147f
C13692 output17/a_27_7# VGND 0.091f
C13693 _216_/A _191_/B 2.88e-19
C13694 _342_/a_27_7# _186_/a_297_7# 4.59e-22
C13695 cal _150_/a_27_7# 2.64e-19
C13696 _330_/a_651_373# VGND 0.00105f
C13697 _330_/a_639_7# VPWR 4.53e-19
C13698 _162_/X _324_/D 1.61e-20
C13699 _242_/A _347_/D 1.44e-20
C13700 _273_/A clkbuf_1_1_0_clk/a_75_172# 9.13e-21
C13701 _345_/a_1602_7# _288_/A 3.21e-20
C13702 _306_/S _172_/Y 0.00122f
C13703 _337_/a_193_7# _283_/A 3.01e-19
C13704 _343_/a_27_7# output41/a_27_7# 4.98e-19
C13705 _250_/X _150_/C 2.09e-20
C13706 _172_/A _188_/S 0.578f
C13707 _346_/SET_B _310_/a_761_249# 0.0145f
C13708 _333_/a_543_7# VGND 0.0177f
C13709 _333_/a_1108_7# VPWR 0.0107f
C13710 _288_/A _309_/Q 0.294f
C13711 _302_/a_323_257# _228_/A 4.34e-20
C13712 _341_/a_1283_n19# _341_/Q 0.00102f
C13713 _337_/Q _195_/a_27_257# 1.08e-21
C13714 _218_/a_256_7# _331_/Q 0.00297f
C13715 _319_/Q _331_/a_1283_n19# 7.49e-20
C13716 _309_/a_1283_n19# _289_/a_39_257# 1.92e-21
C13717 _269_/A _343_/CLK 0.253f
C13718 _342_/D VGND 1.36f
C13719 input1/X output30/a_27_7# 2.46e-19
C13720 _276_/a_68_257# _286_/Y 1.17e-21
C13721 _287_/a_39_257# _309_/Q 4.49e-19
C13722 _297_/A _314_/D 0.113f
C13723 rstn _333_/Q 0.0587f
C13724 _286_/B _347_/Q 0.00115f
C13725 _167_/a_27_257# _345_/Q 2.37e-19
C13726 _196_/A _299_/X 0.00235f
C13727 _273_/Y clkc 0.0248f
C13728 _223_/a_250_257# VPWR 0.00842f
C13729 _294_/A clkbuf_2_3_0_clk/A 0.00635f
C13730 _314_/a_1108_7# _347_/a_543_7# 1.18e-19
C13731 _322_/a_193_7# _322_/a_761_249# -0.00517f
C13732 _277_/Y _194_/A 3.64e-20
C13733 _158_/Y comp 1.85e-20
C13734 _306_/a_76_159# _147_/Y 0.00461f
C13735 _232_/X _212_/a_27_7# 0.0036f
C13736 _344_/a_652_n19# _161_/Y 1.13e-20
C13737 _298_/C _154_/A 1.41e-19
C13738 _343_/D _343_/CLK 0.0798f
C13739 _216_/a_27_7# _248_/B 0.0486f
C13740 _294_/Y _288_/Y 0.00483f
C13741 _258_/S _215_/A 2.11e-19
C13742 _306_/S _192_/B 0.0198f
C13743 _216_/A _331_/a_448_7# 2.68e-21
C13744 _339_/D _284_/A -1.01e-24
C13745 _271_/A _331_/Q 0.074f
C13746 _273_/A _310_/a_1108_7# 3.7e-21
C13747 _258_/S _277_/Y 0.119f
C13748 _342_/Q _206_/A 0.00217f
C13749 _293_/a_39_257# _197_/X 8.78e-21
C13750 _271_/A _182_/a_79_n19# 1.7e-19
C13751 _248_/A _175_/Y 0.0748f
C13752 _330_/D _330_/a_543_7# 2.07e-19
C13753 _251_/X _212_/X 6.82e-20
C13754 _327_/Q _327_/D 0.451f
C13755 _329_/a_1283_n19# _212_/X 0.0257f
C13756 _344_/a_1032_373# _344_/a_1602_7# 1.42e-32
C13757 _339_/a_193_7# _283_/A 0.0208f
C13758 _346_/SET_B _336_/a_27_7# 0.0178f
C13759 output30/a_27_7# _286_/Y 0.0288f
C13760 _281_/Y clk 4.57e-20
C13761 _263_/B VGND 0.0766f
C13762 _283_/A _282_/a_39_257# 0.00162f
C13763 _181_/X _315_/D 0.258f
C13764 _188_/S _244_/B 3.36e-22
C13765 _275_/Y _312_/a_651_373# 0.00269f
C13766 _216_/A _337_/Q 5.35e-19
C13767 _199_/a_93_n19# _340_/CLK 3.8e-19
C13768 _321_/D _242_/A 0.0698f
C13769 _258_/S _262_/a_199_7# 0.00181f
C13770 _239_/a_199_7# _157_/A 3.23e-20
C13771 clkbuf_2_3_0_clk/A _283_/A 3.92e-20
C13772 _286_/B _297_/B 0.0107f
C13773 _319_/a_448_7# _319_/D 0.00455f
C13774 _294_/A ctln[2] 1.21e-19
C13775 _160_/X _347_/a_27_7# 2.03e-21
C13776 _299_/X _347_/a_1283_n19# 4.4e-19
C13777 _258_/a_535_334# _313_/Q 4.18e-19
C13778 _286_/a_113_7# VPWR -6.36e-20
C13779 _304_/a_79_n19# VPWR 0.00917f
C13780 _277_/A _331_/CLK 0.044f
C13781 _324_/a_193_7# _216_/X 0.00939f
C13782 _326_/a_639_7# _326_/Q 3.47e-20
C13783 _279_/Y _227_/A 0.00106f
C13784 _340_/CLK _336_/Q 0.00967f
C13785 _313_/Q _172_/A 8.87e-20
C13786 _256_/a_80_n19# VPWR 0.0864f
C13787 _283_/A _327_/Q 0.00618f
C13788 _342_/Q _147_/A 0.0131f
C13789 _279_/Y _314_/a_1108_7# 0.00396f
C13790 _255_/B _150_/C 0.316f
C13791 _277_/A _273_/A 7.73e-20
C13792 _342_/a_1108_7# _308_/X 9.13e-21
C13793 _317_/a_761_249# _247_/a_113_257# 2.25e-20
C13794 _345_/a_27_7# _292_/A 1.84e-19
C13795 _342_/a_193_7# _342_/a_1283_n19# -7.11e-33
C13796 _342_/a_27_7# _342_/a_1108_7# -2.98e-20
C13797 _313_/Q _198_/a_250_257# 5.04e-21
C13798 output26/a_27_7# result[4] 0.00541f
C13799 _346_/a_27_7# _170_/a_76_159# 2.39e-22
C13800 _321_/D _322_/D 0.0102f
C13801 _344_/a_476_7# _172_/B 0.0052f
C13802 _176_/a_27_7# VPWR 0.0839f
C13803 _154_/a_27_7# _254_/B 0.0112f
C13804 _342_/Q _149_/A 0.177f
C13805 _321_/D _321_/a_448_7# 0.00249f
C13806 _244_/a_109_257# _317_/D 8.7e-19
C13807 _333_/a_27_7# _153_/B 1.88e-21
C13808 _260_/A _344_/Q 2.02e-20
C13809 _338_/D _199_/a_256_7# 5.76e-19
C13810 _309_/a_1108_7# _162_/X 1.77e-21
C13811 _267_/B _297_/Y 0.00619f
C13812 _157_/A _251_/a_297_257# 1.14e-19
C13813 _309_/a_1108_7# _287_/a_39_257# 3.07e-19
C13814 _206_/A _204_/Y 0.0856f
C13815 output15/a_27_7# VGND 0.111f
C13816 _303_/A _228_/A 9.76e-20
C13817 _179_/a_27_7# _254_/B 0.031f
C13818 _327_/a_193_7# _304_/X 0.0065f
C13819 _327_/a_27_7# _217_/A 5.01e-19
C13820 _343_/a_448_7# _343_/Q 4.51e-20
C13821 _343_/a_1283_n19# _298_/C 4.68e-20
C13822 _330_/D _331_/Q 0.0472f
C13823 _166_/Y _301_/X 0.036f
C13824 _346_/a_27_7# clkbuf_2_1_0_clk/A 0.00188f
C13825 _338_/Q _265_/B 1.44e-20
C13826 _332_/a_27_7# VPWR 0.093f
C13827 _248_/B _327_/Q 0.0291f
C13828 _347_/a_193_7# VPWR -0.295f
C13829 _326_/a_27_7# _217_/A 0.00105f
C13830 _326_/a_193_7# _304_/X 0.0134f
C13831 _258_/S _300_/Y 2.29e-21
C13832 _277_/A _319_/a_1108_7# 0.00539f
C13833 _292_/Y output38/a_27_7# 3.46e-19
C13834 _169_/Y _346_/SET_B 2.96e-20
C13835 _334_/D _204_/Y 4.68e-19
C13836 _346_/SET_B _225_/B 5.41e-20
C13837 _254_/Y clkbuf_2_3_0_clk/A 0.0143f
C13838 repeater43/X _321_/a_543_7# 0.0101f
C13839 _319_/Q _280_/a_150_257# 8.78e-19
C13840 _308_/a_218_334# _286_/B 6.05e-19
C13841 _308_/a_76_159# _181_/X 6.42e-19
C13842 output7/a_27_7# _204_/Y 1.03e-19
C13843 _305_/a_218_7# _254_/B 3e-21
C13844 _336_/a_193_7# _313_/a_193_7# 8.4e-20
C13845 _250_/a_78_159# _284_/A 0.0227f
C13846 _297_/B _347_/a_543_7# 0.0302f
C13847 _314_/D _347_/a_761_249# 8.15e-21
C13848 _264_/a_113_257# _147_/A 7.42e-21
C13849 _267_/B _310_/a_193_7# 0.0139f
C13850 comp _160_/a_27_7# 6.69e-19
C13851 _283_/A _192_/B 0.755f
C13852 _341_/Q _248_/A 2.6e-20
C13853 _160_/X _162_/A 2.32e-19
C13854 repeater43/X _153_/a_109_53# 0.00246f
C13855 _146_/C _306_/S 8.12e-22
C13856 _312_/Q _311_/a_761_249# 1.41e-19
C13857 _279_/Y _347_/Q 2.07e-20
C13858 _192_/B _205_/a_382_257# 0.00149f
C13859 _331_/Q _232_/a_27_7# 9.52e-21
C13860 _233_/a_113_257# _232_/X 0.0086f
C13861 _276_/a_68_257# _328_/Q 0.00907f
C13862 _346_/Q _286_/Y 4.5e-20
C13863 _332_/D _154_/A 2.28e-19
C13864 _341_/a_193_7# VGND 0.0308f
C13865 _341_/a_543_7# VPWR 0.0163f
C13866 _194_/A VGND 0.181f
C13867 _298_/B _332_/Q 3.29e-21
C13868 _271_/A _182_/X 5.74e-19
C13869 _157_/A _306_/S 1.23e-19
C13870 _342_/a_1108_7# _317_/D 3.95e-19
C13871 _259_/a_113_257# _275_/Y 4.39e-19
C13872 _275_/Y _286_/B 0.0513f
C13873 _225_/X _335_/Q 1.03e-20
C13874 _338_/a_543_7# VPWR 0.0196f
C13875 _338_/a_193_7# VGND 0.00602f
C13876 ctlp[0] VPWR 0.108f
C13877 _281_/Y _250_/a_292_257# 6.81e-21
C13878 _294_/Y _337_/Q 8.23e-22
C13879 _339_/a_1462_7# _283_/A 0.00185f
C13880 _346_/SET_B _336_/a_1217_7# -1.45e-19
C13881 _320_/Q _220_/a_93_n19# 0.0245f
C13882 _325_/Q _150_/C 4.02e-20
C13883 _258_/S VGND 2.01f
C13884 clkbuf_2_1_0_clk/A _319_/a_27_7# 1.56e-21
C13885 _279_/A _347_/a_651_373# 4.72e-20
C13886 _346_/SET_B _314_/a_543_7# -9.91e-19
C13887 _169_/a_109_257# clkbuf_2_3_0_clk/A 1.93e-20
C13888 _150_/C _298_/a_27_7# 8.23e-20
C13889 output25/a_27_7# _318_/Q 0.0137f
C13890 _185_/A clk 0.00226f
C13891 _342_/a_651_373# _323_/D 3.01e-19
C13892 repeater43/X _209_/a_27_257# 1.77e-19
C13893 _334_/Q _153_/a_109_53# 6.95e-19
C13894 _317_/Q _317_/a_1283_n19# 0.0133f
C13895 _336_/a_27_7# _147_/A 3.08e-19
C13896 _242_/A _317_/a_27_7# 2.14e-19
C13897 _325_/a_27_7# _248_/B 2e-20
C13898 _271_/Y _298_/X 4.53e-21
C13899 _340_/a_1108_7# VPWR 0.00265f
C13900 _340_/a_543_7# VGND 0.00287f
C13901 _236_/a_109_257# _242_/B 0.00157f
C13902 _238_/B _330_/Q 9.17e-21
C13903 _184_/a_76_159# _177_/A 1.76e-19
C13904 _325_/Q _317_/a_193_7# 0.00763f
C13905 output11/a_27_7# VGND 0.0606f
C13906 _254_/Y _192_/B 1.1e-20
C13907 _327_/a_1283_n19# _330_/Q 1.65e-19
C13908 _283_/A _331_/a_1270_373# 9.87e-20
C13909 _316_/a_1283_n19# VPWR 0.0404f
C13910 _316_/a_761_249# VGND -0.00151f
C13911 _343_/a_1283_n19# _229_/a_489_373# 8.95e-21
C13912 _343_/a_1108_7# _229_/a_226_7# 3.9e-20
C13913 _260_/B VPWR 0.374f
C13914 _258_/S _309_/a_761_249# 1.29e-19
C13915 _328_/a_27_7# _220_/a_93_n19# 0.00351f
C13916 _320_/Q VGND 0.54f
C13917 _225_/B _206_/A 0.00217f
C13918 _326_/a_1283_n19# _330_/Q 0.00131f
C13919 _200_/a_250_257# _311_/a_193_7# 4.68e-20
C13920 _279_/Y _297_/B 0.0375f
C13921 clkbuf_2_1_0_clk/A _338_/Q 0.315f
C13922 _313_/a_761_249# _225_/B 6.24e-21
C13923 _327_/a_543_7# VPWR 0.024f
C13924 _327_/a_193_7# VGND 0.00102f
C13925 _183_/a_1241_257# _144_/a_27_7# 1.05e-20
C13926 _275_/A clkbuf_2_1_0_clk/A 0.146f
C13927 _346_/a_193_7# _346_/D 0.146f
C13928 _260_/A _306_/S 0.0188f
C13929 repeater42/a_27_7# _216_/X 0.00281f
C13930 repeater43/X _315_/a_761_249# 0.00575f
C13931 _250_/a_493_257# _250_/X 4.03e-20
C13932 _322_/a_543_7# _322_/Q 2.49e-19
C13933 _326_/a_193_7# VGND 0.0341f
C13934 _326_/a_543_7# VPWR 0.0156f
C13935 repeater43/a_27_7# _227_/A 3.62e-21
C13936 _338_/Q _310_/Q 5.37e-20
C13937 _254_/A _265_/B 1.68e-19
C13938 _294_/Y _339_/Q 6.59e-20
C13939 _161_/Y output40/a_27_7# 4.49e-19
C13940 _232_/X _223_/a_93_n19# 2.25e-21
C13941 _315_/Q VPWR 0.584f
C13942 _156_/a_39_257# _225_/B 0.00695f
C13943 _324_/Q _296_/a_493_257# 3.01e-20
C13944 _332_/a_639_7# VGND 3.52e-19
C13945 _332_/a_1217_7# VPWR 6.07e-20
C13946 _251_/a_79_n19# _251_/a_297_257# 3.55e-33
C13947 _328_/a_761_249# VPWR 0.0114f
C13948 _328_/a_27_7# VGND -0.0891f
C13949 _347_/a_805_7# VGND -5.82e-19
C13950 _221_/a_93_n19# _221_/a_346_7# -3.48e-20
C13951 _347_/a_1462_7# VPWR 1.27e-19
C13952 _193_/Y _267_/A 7.21e-19
C13953 repeater43/X _224_/a_93_n19# 2.18e-19
C13954 _341_/Q _178_/a_27_7# 0.0366f
C13955 _200_/a_584_7# VGND -0.00129f
C13956 _189_/a_27_7# cal 1.07e-20
C13957 trim[0] trim[1] 0.0362f
C13958 _345_/a_27_7# _273_/A 6.68e-20
C13959 en _206_/A 0.00784f
C13960 _269_/A output30/a_27_7# 0.0144f
C13961 _191_/B _209_/a_27_257# 0.00513f
C13962 _192_/B _225_/a_145_35# 7.61e-20
C13963 _234_/B _331_/a_1108_7# 6.91e-22
C13964 _308_/S _181_/X 0.352f
C13965 _255_/B cal 3.49e-19
C13966 _328_/a_1283_n19# _297_/B 0.0112f
C13967 _181_/a_27_7# _162_/X 2.02e-19
C13968 _250_/X _284_/A 0.00428f
C13969 _321_/a_761_249# result[7] 3.68e-20
C13970 _314_/Q _347_/a_639_7# 7.55e-19
C13971 _258_/S _306_/a_218_334# 0.00244f
C13972 _164_/Y _171_/a_78_159# 0.00884f
C13973 _290_/A _284_/A 0.00948f
C13974 _298_/B _226_/a_382_257# 2.5e-19
C13975 _146_/C _283_/A 1.77e-20
C13976 _288_/A _344_/a_1032_373# 1.5e-20
C13977 _324_/a_193_7# _216_/a_27_7# 0.00366f
C13978 _343_/CLK _315_/a_651_373# 0.0265f
C13979 _258_/a_76_159# _286_/B 0.0389f
C13980 _346_/a_476_7# _160_/X 5.24e-19
C13981 _169_/Y _147_/A 4.53e-20
C13982 _165_/X _344_/Q 1.68e-19
C13983 input4/X _154_/A 4.53e-21
C13984 _334_/a_761_249# VPWR 0.0208f
C13985 _334_/a_27_7# VGND -0.0985f
C13986 repeater43/X _153_/A 0.0141f
C13987 _225_/X _336_/Q 1.22e-19
C13988 _306_/X _147_/Y 0.0163f
C13989 _320_/Q output27/a_27_7# 0.0132f
C13990 _147_/A _225_/B 0.0297f
C13991 _257_/a_79_159# _197_/a_27_7# 1.08e-21
C13992 ctln[4] _338_/Q 3.73e-20
C13993 _281_/Y _329_/D 0.00913f
C13994 _163_/a_78_159# _160_/X 0.069f
C13995 _301_/X _297_/Y 0.0397f
C13996 _312_/D _311_/D 0.00169f
C13997 clkbuf_1_0_0_clk/a_75_172# _281_/A 6.07e-19
C13998 _344_/a_1032_373# _162_/X 0.00626f
C13999 _309_/D _265_/B 5.07e-19
C14000 _294_/A _260_/A 3.09e-20
C14001 _307_/a_218_334# _227_/A 4.12e-19
C14002 _323_/a_761_249# _298_/X 2.42e-20
C14003 _342_/Q _150_/a_27_7# 0.147f
C14004 _267_/B _336_/Q 5.14e-21
C14005 _326_/Q _150_/C 1.15e-20
C14006 _341_/a_1462_7# VGND -8.91e-19
C14007 _346_/SET_B _315_/D 0.188f
C14008 _338_/a_1462_7# VGND 0.00172f
C14009 _323_/a_193_7# _343_/Q 0.00707f
C14010 clk _335_/Q 0.0125f
C14011 _168_/a_109_7# _165_/X 0.0324f
C14012 _314_/a_543_7# _156_/a_39_257# 4.79e-19
C14013 input3/a_27_7# _191_/B 1.89e-19
C14014 _207_/C _154_/A 0.0123f
C14015 _274_/a_121_257# VPWR 4.98e-19
C14016 _330_/a_193_7# _330_/a_448_7# -0.00482f
C14017 _270_/a_39_257# _324_/Q 2.83e-20
C14018 _330_/Q _248_/A 0.284f
C14019 _329_/a_761_249# _281_/A 0.0234f
C14020 _146_/C _248_/B 8.29e-20
C14021 output35/a_27_7# _309_/Q 2.38e-19
C14022 _304_/S _224_/a_346_7# 6.18e-20
C14023 _254_/A _170_/a_76_159# 0.00271f
C14024 _342_/a_27_7# _177_/a_27_7# 7.66e-20
C14025 _334_/Q _153_/A 4.12e-19
C14026 _321_/Q _316_/D 0.184f
C14027 _330_/Q _331_/CLK 0.139f
C14028 _157_/A _248_/B 3.32e-20
C14029 _295_/a_306_7# VGND -5.05e-19
C14030 _295_/a_512_7# VPWR 0.00219f
C14031 _346_/a_652_n19# VGND 0.0193f
C14032 _346_/a_1182_221# VPWR 0.0034f
C14033 _337_/Q _310_/a_639_7# 4.62e-19
C14034 _337_/D _199_/a_250_257# 8.8e-20
C14035 _160_/X _173_/a_489_373# 0.0387f
C14036 _335_/a_27_7# _204_/a_277_7# 7.9e-21
C14037 _188_/S _177_/A 0.0102f
C14038 _163_/a_292_257# VPWR -5.64e-19
C14039 _248_/A _314_/D 3e-21
C14040 _335_/a_193_7# _208_/a_215_7# 7.06e-20
C14041 _335_/a_1283_n19# _208_/a_78_159# 2.99e-19
C14042 _329_/a_27_7# _319_/Q 0.0505f
C14043 _343_/a_193_7# _226_/a_79_n19# 6.88e-20
C14044 _345_/a_562_373# _346_/SET_B 6.46e-19
C14045 _254_/A clkbuf_2_1_0_clk/A 0.00987f
C14046 _347_/Q _313_/a_27_7# 1.7e-21
C14047 _299_/X _313_/a_193_7# 4.4e-19
C14048 _273_/A _330_/Q 4.75e-21
C14049 _324_/a_805_7# _331_/CLK 3.6e-19
C14050 _346_/a_193_7# _314_/Q 0.00128f
C14051 _340_/CLK _311_/a_761_249# 3.02e-19
C14052 _283_/A _260_/A 9.26e-21
C14053 _333_/Q VPWR 0.381f
C14054 _207_/X VGND 1.03f
C14055 _342_/Q _250_/a_78_159# 0.00633f
C14056 _191_/B _153_/A 0.247f
C14057 _254_/Y _157_/A 2.32e-21
C14058 _318_/a_761_249# _331_/CLK 1.66e-20
C14059 _236_/B _318_/a_27_7# 3.82e-20
C14060 _254_/A _310_/Q 3.47e-20
C14061 _201_/a_27_7# VGND 0.0871f
C14062 _327_/a_1462_7# VGND -9.09e-19
C14063 _301_/X _242_/A 0.00167f
C14064 _342_/a_805_7# _342_/D 0.00213f
C14065 _346_/a_796_7# _346_/D 3.69e-19
C14066 _162_/a_27_7# _265_/B 1.04e-19
C14067 _298_/C _153_/B 7.18e-20
C14068 _227_/A _144_/A 1.94e-20
C14069 repeater43/X _318_/D 0.00213f
C14070 _194_/X _193_/Y 0.117f
C14071 _340_/Q _306_/S 0.0367f
C14072 _326_/a_1462_7# VGND -8.11e-19
C14073 _211_/a_27_257# _332_/a_27_7# 5.13e-19
C14074 cal _298_/a_27_7# 0.017f
C14075 _286_/B _161_/Y 3.51e-19
C14076 _215_/A _313_/a_651_373# 0.0263f
C14077 _300_/a_301_257# _157_/a_27_7# 6.09e-20
C14078 _254_/A _300_/a_735_7# 0.00202f
C14079 _273_/A _314_/D 3.56e-19
C14080 _290_/A trim[2] 0.00504f
C14081 repeater43/X _324_/a_543_7# -9.96e-19
C14082 _296_/Y _341_/Q 7.2e-20
C14083 ctln[6] _340_/D 7.01e-21
C14084 _242_/B _327_/Q 0.00421f
C14085 _180_/a_183_257# VGND -2.84e-19
C14086 _332_/a_448_7# _153_/B 0.00783f
C14087 _324_/a_193_7# _327_/Q 1.53e-19
C14088 _324_/a_27_7# _212_/X 0.00118f
C14089 _255_/B _284_/A 0.202f
C14090 _343_/a_761_249# repeater43/X 0.0138f
C14091 _251_/a_297_257# _251_/X 1.69e-19
C14092 _328_/a_1217_7# VGND -4.95e-19
C14093 _298_/B _192_/B 1.83e-19
C14094 _331_/Q _330_/a_1283_n19# 1.66e-20
C14095 _173_/a_226_7# VGND 0.00671f
C14096 _173_/a_226_257# VPWR -7.25e-19
C14097 _341_/Q _146_/a_29_271# 0.0221f
C14098 clkbuf_2_1_0_clk/A _309_/D 1.69e-19
C14099 repeater43/X _217_/A 0.0283f
C14100 _177_/a_27_7# _317_/D 0.0317f
C14101 _285_/A _162_/A 0.0854f
C14102 _271_/Y _334_/a_1108_7# 8.39e-21
C14103 _271_/A _334_/a_651_373# 0.0267f
C14104 _319_/a_761_249# VGND 0.0209f
C14105 _319_/a_1283_n19# VPWR 0.0302f
C14106 _215_/A _157_/a_27_7# 6.12e-20
C14107 _346_/SET_B _311_/a_543_7# 0.00803f
C14108 _338_/Q _311_/a_27_7# 9.44e-20
C14109 _337_/a_27_7# VGND -0.0566f
C14110 _337_/a_761_249# VPWR 0.00848f
C14111 _165_/X _306_/S 0.00642f
C14112 _164_/Y _172_/B 1.96e-19
C14113 _342_/a_27_7# _341_/a_27_7# 1.22e-20
C14114 _309_/D _310_/Q 0.00185f
C14115 clkbuf_2_1_0_clk/a_75_172# _331_/CLK 0.00197f
C14116 _319_/a_448_7# _297_/B 2.28e-19
C14117 _340_/a_27_7# _305_/a_505_n19# 7.53e-21
C14118 _344_/a_193_7# _162_/A 9.3e-21
C14119 _334_/a_1217_7# VGND -5.03e-19
C14120 output8/a_27_7# VPWR 0.125f
C14121 clk _209_/a_373_7# 2.05e-19
C14122 clk _336_/Q 6.78e-20
C14123 _254_/Y _260_/A 0.203f
C14124 _167_/a_109_257# _166_/Y -5.55e-35
C14125 _167_/a_373_7# _346_/Q 7.65e-19
C14126 _236_/B _246_/B 2.04e-19
C14127 _301_/a_149_7# _267_/A 2.13e-20
C14128 _341_/a_1283_n19# _188_/S 2.1e-20
C14129 _309_/a_448_7# _340_/CLK 5.27e-20
C14130 _255_/a_184_257# _306_/S 4.99e-20
C14131 input1/X _209_/X 2.44e-20
C14132 _329_/Q _320_/a_1283_n19# 3.78e-19
C14133 _320_/Q _320_/a_1108_7# 0.00173f
C14134 _238_/B _320_/a_761_249# 6.14e-21
C14135 _315_/D _156_/a_39_257# 5.52e-19
C14136 _307_/a_76_159# VPWR 0.0347f
C14137 _145_/A _227_/A 0.165f
C14138 _323_/D output41/a_27_7# 1.21e-19
C14139 _345_/a_1602_7# _345_/Q 0.0364f
C14140 _345_/a_1032_373# _345_/D 1.3e-19
C14141 _294_/A _340_/Q 0.00426f
C14142 result[1] _248_/A 8.01e-20
C14143 _343_/a_651_373# _343_/CLK 5.9e-20
C14144 _325_/a_651_373# _326_/Q 0.00219f
C14145 _339_/D _225_/B 3.1e-20
C14146 _324_/a_448_7# _304_/S 0.0219f
C14147 _292_/A _285_/Y 0.00674f
C14148 _172_/A _162_/A 0.00163f
C14149 clkbuf_2_3_0_clk/A _160_/X 0.0131f
C14150 _172_/A _216_/X 7.61e-21
C14151 _316_/Q _236_/B 1e-20
C14152 _251_/X _306_/S 2.72e-21
C14153 result[1] _331_/CLK 1.73e-19
C14154 _326_/D _246_/B 9.06e-21
C14155 _326_/a_193_7# _214_/a_27_257# 2.85e-19
C14156 _166_/Y _297_/Y 1.3e-20
C14157 _268_/a_121_257# _317_/D 2.33e-20
C14158 _184_/a_76_159# _248_/A 7.45e-20
C14159 _306_/S _296_/a_213_83# 0.0207f
C14160 _315_/D _147_/A 1.25e-20
C14161 _340_/a_1283_n19# _198_/a_250_257# 2.03e-19
C14162 _342_/a_651_373# _177_/A 4.9e-20
C14163 _226_/a_297_7# VPWR -1.59e-19
C14164 _226_/a_79_n19# VGND 0.00575f
C14165 _216_/X _232_/X 0.0367f
C14166 _188_/a_439_7# VGND -5.95e-19
C14167 _325_/a_193_7# _324_/a_27_7# 1.23e-20
C14168 _325_/a_27_7# _324_/a_193_7# 0.00182f
C14169 _294_/A _165_/X 1.07e-20
C14170 _149_/A _315_/D 5.23e-20
C14171 _346_/a_1296_7# VPWR 1.34e-19
C14172 _346_/a_1056_7# VGND -5.94e-19
C14173 _160_/X _172_/Y 0.0234f
C14174 rstn _207_/a_27_7# 0.096f
C14175 _335_/a_1108_7# _333_/Q 1.19e-20
C14176 _335_/a_1283_n19# _190_/A 7.41e-20
C14177 _329_/Q _232_/X 0.0229f
C14178 _169_/a_109_257# _260_/A 5.38e-19
C14179 _158_/Y VGND 0.187f
C14180 _248_/B _221_/a_250_257# 4.68e-19
C14181 clkbuf_0_clk/X _314_/a_27_7# 0.0176f
C14182 clkbuf_0_clk/a_110_7# _314_/a_448_7# 9.3e-20
C14183 _309_/a_651_373# _346_/SET_B 0.00383f
C14184 _305_/X _254_/B 0.00347f
C14185 _343_/a_1108_7# _225_/X 2.43e-20
C14186 _343_/a_1283_n19# _150_/C 1.21e-20
C14187 _343_/a_543_7# _226_/X 0.00168f
C14188 _341_/a_27_7# _317_/D 0.012f
C14189 _341_/a_761_249# _244_/B 1.69e-20
C14190 _339_/a_761_249# VPWR 0.0105f
C14191 _339_/a_27_7# VGND -0.0902f
C14192 _327_/a_761_249# _232_/X 0.00613f
C14193 _308_/a_76_159# _206_/A 1.06e-20
C14194 _282_/a_121_257# VPWR -3.8e-19
C14195 _271_/A _143_/a_181_7# 4.57e-20
C14196 _150_/C _324_/D 1.64e-22
C14197 _342_/Q _250_/X 0.0247f
C14198 _169_/Y _174_/a_109_7# 5.74e-20
C14199 _323_/a_1283_n19# _334_/a_543_7# 1.52e-20
C14200 _283_/Y _338_/a_1270_373# 4.43e-20
C14201 _283_/A _340_/Q 0.00455f
C14202 _326_/a_761_249# _232_/X 0.00307f
C14203 _321_/D _318_/a_639_7# 0.00103f
C14204 _235_/a_113_257# _331_/a_1108_7# 2.49e-19
C14205 _292_/Y _290_/A 1.83e-19
C14206 _320_/Q ctlp[5] 0.00126f
C14207 _330_/Q _217_/X 0.0877f
C14208 _312_/a_1283_n19# _312_/D 3.82e-21
C14209 _312_/a_27_7# _312_/Q 0.0038f
C14210 _300_/Y _157_/a_27_7# 0.00159f
C14211 _281_/Y _242_/A 0.0045f
C14212 input1/X _336_/a_1270_373# 2.49e-19
C14213 _328_/a_193_7# _232_/X 0.00214f
C14214 clkbuf_0_clk/X clkbuf_2_1_0_clk/A 0.966f
C14215 _212_/X VPWR 1.28f
C14216 _223_/a_93_n19# _223_/a_256_7# -3.48e-20
C14217 _332_/D _153_/B 0.034f
C14218 _256_/a_80_n19# _147_/Y 0.00119f
C14219 _316_/Q _343_/CLK 0.0045f
C14220 repeater43/X _318_/a_448_7# 0.00395f
C14221 _269_/A _247_/a_113_257# 2.42e-19
C14222 _316_/a_193_7# _317_/D 0.0144f
C14223 _316_/a_543_7# _244_/B 0.00391f
C14224 _329_/a_27_7# _329_/a_639_7# -0.0015f
C14225 _329_/a_1283_n19# _329_/a_1108_7# 5.68e-32
C14226 _166_/Y _242_/A 1.84e-19
C14227 _298_/B _146_/C 4.81e-20
C14228 _318_/a_1283_n19# _327_/Q 2.14e-19
C14229 _309_/a_193_7# clkbuf_2_3_0_clk/A 4.46e-21
C14230 _271_/Y _343_/CLK 0.0949f
C14231 _313_/a_651_373# VGND 0.0024f
C14232 _313_/a_639_7# VPWR 1.06e-19
C14233 _157_/A _300_/a_27_257# 0.00525f
C14234 ctln[7] _204_/a_27_257# 1.85e-19
C14235 _337_/a_1217_7# VGND -4.52e-19
C14236 _328_/a_27_7# ctlp[5] 7.04e-20
C14237 _335_/a_193_7# _334_/D 4.34e-19
C14238 _335_/a_761_249# _343_/CLK 0.00109f
C14239 repeater42/a_27_7# _327_/Q 0.0118f
C14240 _181_/X _333_/a_193_7# 4.58e-22
C14241 _321_/Q output28/a_27_7# 0.0311f
C14242 _271_/A _304_/S 0.00636f
C14243 _250_/a_78_159# _225_/B 7.06e-20
C14244 cal _154_/A 0.00197f
C14245 _344_/a_193_7# _163_/a_78_159# 0.0103f
C14246 _254_/Y _340_/Q 0.00273f
C14247 result[6] _318_/D 1.65e-20
C14248 clkbuf_2_1_0_clk/A input1/X 0.32f
C14249 _165_/a_78_159# _172_/B 0.0033f
C14250 _157_/a_27_7# VGND 0.0592f
C14251 _167_/X _301_/a_149_7# 0.00324f
C14252 _147_/Y _347_/a_193_7# 3.37e-22
C14253 _274_/a_39_257# _232_/X 0.00505f
C14254 rstn _306_/S 0.136f
C14255 _320_/Q _330_/a_27_7# 0.0312f
C14256 _172_/A _295_/a_409_7# 1.4e-19
C14257 _283_/Y _340_/CLK 0.00802f
C14258 _309_/D _311_/a_27_7# 1.16e-19
C14259 _267_/B _311_/a_761_249# 4.11e-21
C14260 _342_/a_1283_n19# _229_/a_76_159# 0.00126f
C14261 _327_/a_27_7# _331_/D 1.55e-19
C14262 _306_/X _260_/B 1.74e-19
C14263 _318_/Q _320_/Q 0.00196f
C14264 _271_/A _225_/X 0.00376f
C14265 _307_/X _271_/A 8.83e-20
C14266 _323_/Q VGND 0.244f
C14267 _169_/B _284_/A 1.61e-20
C14268 _258_/a_505_n19# _190_/A 1.21e-21
C14269 _319_/Q _321_/a_651_373# 1.63e-19
C14270 _327_/a_193_7# _318_/Q 1.35e-19
C14271 _326_/a_27_7# _331_/D 7.1e-19
C14272 _188_/S _248_/A 1.55e-20
C14273 _164_/Y trimb[4] 1.16e-19
C14274 _276_/a_68_257# _299_/X 2.53e-20
C14275 _340_/a_639_7# _197_/X 5.71e-19
C14276 _331_/a_193_7# _246_/B 1.73e-20
C14277 output19/a_27_7# _346_/SET_B 1.38e-20
C14278 _306_/a_505_n19# clkbuf_2_3_0_clk/A 0.00226f
C14279 _324_/Q _227_/A 0.128f
C14280 _326_/a_193_7# _318_/Q 4.8e-20
C14281 clk output6/a_27_7# 0.00714f
C14282 ctln[5] _197_/X 1.61e-20
C14283 _325_/a_193_7# VPWR -0.0971f
C14284 _302_/a_539_257# _300_/Y 0.00175f
C14285 _325_/a_651_373# _324_/a_1108_7# 4.58e-21
C14286 _344_/Q _310_/D 6.12e-20
C14287 ctln[7] _334_/a_1108_7# 2.6e-21
C14288 _271_/A _317_/a_27_7# 0.00105f
C14289 _157_/A _314_/a_1270_373# 5.17e-20
C14290 _211_/a_109_257# _332_/Q 0.0292f
C14291 _323_/a_193_7# _206_/A 1.47e-19
C14292 _160_/a_27_7# VGND 0.134f
C14293 _255_/B _342_/Q 0.0546f
C14294 _149_/a_27_7# VPWR 0.142f
C14295 _335_/D _332_/Q 0.00117f
C14296 _212_/a_27_7# _248_/A 8.74e-20
C14297 _251_/X _248_/B 0.0532f
C14298 _273_/A _285_/Y 0.376f
C14299 clkbuf_0_clk/a_110_7# _314_/D 0.00284f
C14300 _341_/a_1217_7# _317_/D 1.59e-19
C14301 _339_/a_1217_7# VGND -4.51e-19
C14302 _255_/B _144_/a_27_7# 9.65e-19
C14303 clkbuf_2_1_0_clk/A _286_/Y 0.0106f
C14304 _328_/a_27_7# _318_/Q 5.18e-21
C14305 _308_/S _206_/A 2.51e-19
C14306 _333_/a_27_7# _332_/a_1108_7# 3.51e-21
C14307 _333_/a_193_7# _332_/a_1283_n19# 9e-20
C14308 _333_/a_1283_n19# _332_/a_193_7# 6.46e-20
C14309 _333_/a_1108_7# _332_/a_27_7# 1.36e-19
C14310 _306_/S _225_/a_59_35# 1.45e-19
C14311 _259_/a_113_257# _263_/B 0.0495f
C14312 _325_/a_805_7# _304_/X 0.0021f
C14313 _317_/a_1283_n19# VGND 0.0254f
C14314 _317_/a_448_7# VPWR 0.00193f
C14315 _281_/Y _336_/Q 0.455f
C14316 _323_/a_193_7# _334_/D 7.39e-21
C14317 _323_/a_761_249# _343_/CLK 0.00777f
C14318 _182_/a_510_7# _196_/A 0.00742f
C14319 repeater42/a_27_7# _325_/a_27_7# 1.81e-20
C14320 result[2] _269_/A 0.0792f
C14321 repeater43/X _335_/a_1270_373# -2.06e-19
C14322 _297_/A _347_/a_27_7# 0.226f
C14323 _258_/a_76_159# _313_/a_27_7# 0.00103f
C14324 _330_/Q _331_/a_805_7# 4.96e-19
C14325 clkbuf_0_clk/X _278_/a_68_257# 1.49e-19
C14326 _318_/a_543_7# _317_/a_448_7# 6.21e-20
C14327 _258_/S output32/a_27_7# 0.0218f
C14328 input4/X _153_/B 8.1e-20
C14329 _292_/A _312_/a_1283_n19# 0.0118f
C14330 _314_/a_193_7# _284_/A 0.00228f
C14331 _312_/a_1217_7# _312_/Q 1.74e-20
C14332 _340_/a_1108_7# _147_/Y 2.01e-21
C14333 _331_/a_651_373# VGND 0.00418f
C14334 result[7] VGND 0.31f
C14335 _331_/a_639_7# VPWR 5.21e-19
C14336 _320_/a_805_7# _346_/SET_B 5.87e-19
C14337 _310_/a_193_7# _297_/Y 2.12e-20
C14338 _172_/A _216_/a_27_7# 1.61e-20
C14339 _302_/a_539_257# VGND -9.17e-19
C14340 _223_/a_93_n19# _325_/D 0.00541f
C14341 _283_/A _232_/A 1.33e-20
C14342 _344_/a_381_7# _346_/SET_B 0.00243f
C14343 _215_/A _267_/A 0.132f
C14344 _343_/a_1283_n19# cal 0.00527f
C14345 _308_/a_439_7# _192_/B 7.35e-19
C14346 _336_/a_543_7# _193_/Y 7.16e-19
C14347 _336_/a_1108_7# _340_/Q 2.99e-21
C14348 _336_/a_1283_n19# _306_/S 9.96e-21
C14349 _163_/a_215_7# _161_/Y 0.00494f
C14350 _277_/Y _267_/A 0.0192f
C14351 _207_/C _153_/B 1.32e-19
C14352 _255_/a_30_13# _209_/a_27_257# 4.93e-21
C14353 _294_/Y output31/a_27_7# 0.00815f
C14354 _313_/D _346_/SET_B 0.0395f
C14355 _234_/B _269_/A 2.26e-21
C14356 _303_/A _217_/A 7.64e-20
C14357 _342_/a_1108_7# _341_/D 1.95e-22
C14358 _182_/a_79_n19# _298_/C 1.94e-19
C14359 _322_/a_448_7# _331_/CLK 3.38e-20
C14360 _322_/a_761_249# _321_/D 0.00127f
C14361 _325_/a_1283_n19# _246_/B 1.13e-19
C14362 _342_/D _341_/a_1108_7# 1.15e-20
C14363 _310_/a_27_7# _310_/a_761_249# -0.0166f
C14364 ctln[1] _335_/a_448_7# 7.79e-19
C14365 _308_/S _147_/A 0.0126f
C14366 _240_/a_109_257# _319_/D 0.00121f
C14367 _227_/A _228_/A 0.179f
C14368 _323_/a_193_7# _149_/A 1.13e-19
C14369 _297_/B _174_/a_27_257# 2.28e-19
C14370 rstn _283_/A 2.87e-20
C14371 _264_/a_113_257# _310_/a_27_7# 8.51e-20
C14372 _232_/A _248_/B 0.176f
C14373 _197_/X _346_/SET_B 0.404f
C14374 _186_/a_382_257# _147_/A 0.00112f
C14375 _184_/a_76_159# _146_/a_29_271# 8.98e-21
C14376 _324_/a_1283_n19# _286_/Y 0.00129f
C14377 _340_/CLK _312_/a_27_7# 0.0383f
C14378 _188_/S _178_/a_27_7# 0.0205f
C14379 _342_/a_651_373# _248_/A 0.00504f
C14380 _325_/Q _144_/a_27_7# 1.07e-19
C14381 output27/a_27_7# result[7] 1.4e-20
C14382 _297_/A _216_/X 0.00594f
C14383 _271_/A clk 0.0322f
C14384 repeater43/X _323_/a_1270_373# 3.23e-20
C14385 result[6] _318_/a_448_7# 3.73e-20
C14386 _344_/a_193_7# clkbuf_2_3_0_clk/A 1.81e-20
C14387 _313_/Q _190_/A 9.04e-21
C14388 clk _335_/a_27_7# 0.00351f
C14389 _257_/a_79_159# _336_/a_27_7# 0.0102f
C14390 result[4] _318_/D 0.00585f
C14391 _192_/a_150_257# _194_/A 3.83e-19
C14392 repeater43/X _214_/a_109_257# 1.97e-19
C14393 _330_/D _331_/a_543_7# 1.53e-19
C14394 _320_/a_761_249# _217_/X 1.65e-21
C14395 _164_/A _162_/A 8.07e-20
C14396 _216_/A _227_/A 0.581f
C14397 _293_/a_39_257# _254_/A 0.0493f
C14398 _328_/a_1462_7# _320_/D 3.31e-21
C14399 _325_/a_805_7# VGND -4.63e-19
C14400 _160_/X _260_/A 6.44e-20
C14401 _343_/CLK _244_/a_109_257# 0.0012f
C14402 _339_/a_761_249# _198_/a_93_n19# 7.02e-22
C14403 _321_/a_27_7# _321_/a_193_7# -0.327f
C14404 ctln[7] _343_/CLK 0.516f
C14405 _172_/A clkbuf_2_3_0_clk/A 0.00893f
C14406 _271_/A _317_/a_1217_7# 1.16e-19
C14407 _324_/Q _297_/B 2.13e-21
C14408 _196_/A _305_/X 4.44e-20
C14409 cal _311_/a_193_7# 6.21e-20
C14410 input1/X _311_/a_27_7# 7.95e-21
C14411 _344_/a_1032_373# _345_/Q 0.00107f
C14412 _324_/a_193_7# _251_/a_79_n19# 1.15e-20
C14413 _286_/B _194_/A 0.637f
C14414 _165_/a_78_159# trimb[4] 1.52e-19
C14415 repeater43/X _308_/X 1.62e-21
C14416 _299_/X _344_/D 2.21e-20
C14417 _342_/a_27_7# repeater43/X 0.00374f
C14418 _340_/Q _194_/a_27_7# 0.0107f
C14419 _259_/a_113_257# _258_/S 0.0139f
C14420 _255_/a_30_13# _153_/A 4.56e-21
C14421 _346_/SET_B _312_/a_193_7# 0.00291f
C14422 _258_/S _286_/B 0.351f
C14423 _326_/a_1283_n19# _223_/a_93_n19# 1.3e-19
C14424 _304_/X _221_/a_93_n19# 0.00319f
C14425 _202_/a_346_7# VGND -0.00162f
C14426 _346_/Q _299_/X 0.00982f
C14427 output13/a_27_7# _323_/Q 1.22e-19
C14428 _317_/Q _243_/a_113_257# 5.49e-19
C14429 _297_/A _347_/a_1217_7# 3.71e-19
C14430 _300_/Y _267_/A 5.23e-20
C14431 _215_/A _194_/X 1.9e-22
C14432 ctlp[7] output15/a_27_7# 8.28e-20
C14433 _172_/A _172_/Y 0.647f
C14434 _219_/a_346_7# _279_/A 9.56e-19
C14435 _294_/Y _291_/a_39_257# 5.44e-20
C14436 _277_/Y _194_/X 2.27e-19
C14437 _341_/a_761_249# _177_/A 0.00106f
C14438 _232_/X _327_/Q 0.25f
C14439 _168_/a_481_7# _299_/X 1.66e-19
C14440 _340_/a_761_249# _196_/A 5.42e-19
C14441 _210_/a_109_257# _209_/X 9.42e-19
C14442 _321_/Q _281_/A 0.00686f
C14443 _269_/A _315_/a_543_7# 0.00354f
C14444 _324_/D _284_/A 1.96e-20
C14445 _197_/X _206_/A 7.01e-19
C14446 _289_/a_39_257# _346_/SET_B 0.00768f
C14447 _323_/a_651_373# _323_/Q 6.5e-19
C14448 _294_/A _310_/D 0.00667f
C14449 clkbuf_2_1_0_clk/A _328_/Q 5.7e-19
C14450 _197_/X _337_/a_448_7# 8.81e-19
C14451 _275_/Y _174_/a_27_257# 0.0108f
C14452 _189_/a_27_7# _225_/B 4.57e-20
C14453 _342_/a_1108_7# _343_/CLK 8.02e-20
C14454 _212_/a_27_7# _217_/X 2.6e-19
C14455 _303_/A _314_/Q 0.228f
C14456 _265_/B clkc 0.00113f
C14457 _167_/X _215_/A 9.98e-21
C14458 _304_/a_257_159# _216_/X 0.0288f
C14459 _255_/B _225_/B 2.82e-20
C14460 _323_/a_27_7# clk 0.00185f
C14461 _281_/Y _324_/a_448_7# 0.006f
C14462 _344_/Q VPWR 0.78f
C14463 _257_/a_79_159# _225_/B 7.73e-19
C14464 _216_/A _347_/Q 3.17e-21
C14465 _281_/A _297_/B 2.89e-21
C14466 _277_/Y _167_/X 0.00205f
C14467 _309_/Q _284_/A 0.635f
C14468 _182_/X _298_/C 5.46e-20
C14469 ctln[1] _335_/D 0.0216f
C14470 _323_/a_1462_7# _149_/A 2.91e-19
C14471 _256_/a_80_n19# _260_/B -9.39e-21
C14472 _322_/D _242_/A 0.0105f
C14473 _172_/A _192_/B 1.15e-19
C14474 _232_/A _315_/a_27_7# 6.15e-19
C14475 _267_/A VGND 2.36f
C14476 _296_/Y _188_/S 0.00839f
C14477 repeater43/X _317_/D 0.881f
C14478 _239_/a_199_7# VPWR -3.26e-19
C14479 clkbuf_0_clk/X _328_/D 9.33e-19
C14480 _144_/a_27_7# _326_/Q 4.57e-22
C14481 _297_/B _228_/A 0.0445f
C14482 _313_/D _147_/A 0.156f
C14483 output18/a_27_7# _319_/a_1108_7# 1.15e-19
C14484 _265_/B _310_/a_543_7# 2.14e-19
C14485 _345_/a_193_7# _306_/S 5.65e-20
C14486 _168_/a_109_7# VPWR 0.0214f
C14487 _207_/a_27_7# VPWR 0.0295f
C14488 VGND sample 0.172f
C14489 _335_/D _192_/B 0.0185f
C14490 _188_/S _146_/a_29_271# 0.00125f
C14491 _342_/a_193_7# _226_/X 0.0012f
C14492 _309_/a_27_7# _344_/Q 1.7e-21
C14493 _153_/a_403_257# _335_/Q 6.88e-19
C14494 _346_/a_27_7# _299_/a_78_159# 3.97e-19
C14495 _342_/Q _315_/a_1283_n19# 2.43e-21
C14496 _298_/C valid 2.77e-19
C14497 _276_/a_68_257# _320_/a_27_7# 2.1e-20
C14498 _342_/a_1283_n19# _149_/A 0.00645f
C14499 _333_/a_1283_n19# _190_/A 3.89e-19
C14500 _333_/a_1108_7# _333_/Q 0.00287f
C14501 _248_/A _223_/a_93_n19# 7.92e-19
C14502 _162_/X _340_/CLK 1.61e-20
C14503 _254_/Y _336_/a_1283_n19# 0.0479f
C14504 _325_/a_27_7# _232_/X 3.16e-19
C14505 _345_/a_381_7# _166_/Y 1.33e-19
C14506 _341_/a_193_7# _341_/a_1108_7# -0.00656f
C14507 _341_/a_27_7# _341_/a_448_7# -0.00642f
C14508 _309_/a_761_249# _267_/A 1.16e-19
C14509 _200_/a_93_n19# _340_/a_27_7# 3.54e-21
C14510 _292_/Y output39/a_27_7# 0.025f
C14511 repeater43/X _331_/D 0.0614f
C14512 _162_/X _347_/D 2.32e-20
C14513 _250_/X _315_/D 1.98e-20
C14514 repeater43/X _330_/a_193_7# 0.00223f
C14515 _216_/X _325_/D 2.82e-20
C14516 _260_/B _347_/a_193_7# 9.55e-20
C14517 _210_/a_27_7# _298_/A 8.84e-20
C14518 _334_/Q _254_/B 2.28e-20
C14519 output33/a_27_7# VPWR 0.0681f
C14520 _164_/A _163_/a_78_159# 0.00175f
C14521 _197_/X _339_/a_448_7# 3.41e-21
C14522 _345_/a_652_n19# _165_/X 3.46e-20
C14523 _251_/a_297_257# VPWR -0.00242f
C14524 ctlp[7] _320_/Q 4.56e-22
C14525 _338_/a_27_7# _338_/a_448_7# -0.00297f
C14526 _338_/a_193_7# _338_/a_1108_7# -0.00817f
C14527 _221_/a_256_7# VPWR -4.57e-19
C14528 _221_/a_93_n19# VGND -0.00346f
C14529 result[4] _318_/a_448_7# 2.81e-19
C14530 _324_/a_193_7# _251_/X 0.00134f
C14531 _216_/A _297_/B 6.35e-20
C14532 _341_/Q _205_/a_297_7# 1.05e-20
C14533 _273_/A _223_/a_93_n19# 7.01e-19
C14534 _342_/a_1217_7# repeater43/X -1.57e-19
C14535 _191_/B _203_/a_209_7# 1.34e-19
C14536 _192_/B _203_/a_80_n19# 0.0117f
C14537 _342_/Q _154_/A 1.61e-20
C14538 _346_/SET_B _312_/a_1462_7# 6.45e-19
C14539 _191_/B _254_/B 0.384f
C14540 _326_/a_761_249# _325_/D 4.86e-21
C14541 _329_/a_543_7# _304_/X 0.0111f
C14542 _322_/a_1108_7# output28/a_27_7# 0.00173f
C14543 _333_/a_193_7# _206_/A 0.596f
C14544 _184_/a_439_7# input1/X 5.09e-19
C14545 _279_/Y _194_/A 0.0113f
C14546 _313_/Q _313_/a_805_7# 2.13e-20
C14547 _231_/a_79_n19# _304_/S 0.00632f
C14548 _294_/A _266_/a_113_257# 0.00502f
C14549 output34/a_27_7# trim[3] 0.00949f
C14550 _258_/a_439_7# _337_/Q 1.07e-22
C14551 _337_/Q _311_/Q 1.5e-20
C14552 _341_/D _177_/a_27_7# 4.53e-20
C14553 _181_/X _295_/a_79_n19# 0.0401f
C14554 _196_/A _295_/a_676_257# 6.39e-19
C14555 cal _153_/B 1.16e-19
C14556 _328_/Q _278_/a_68_257# 2.67e-19
C14557 _165_/X _160_/X 0.155f
C14558 _167_/X _300_/Y 1.1e-19
C14559 _200_/a_93_n19# _200_/a_250_257# -6.97e-22
C14560 _283_/Y clk 0.00332f
C14561 _267_/A _311_/a_639_7# 0.00152f
C14562 _297_/A _216_/a_27_7# 1.47e-20
C14563 _292_/A _162_/A 2.13e-19
C14564 _310_/Q clkc 3.69e-20
C14565 _343_/CLK _333_/a_761_249# 9.01e-21
C14566 _258_/S _279_/Y 2.25e-20
C14567 _175_/Y _298_/A 0.01f
C14568 _230_/a_27_7# _242_/B 0.0472f
C14569 _275_/A ctlp[3] 0.0121f
C14570 _197_/X _337_/D 0.258f
C14571 _241_/a_113_257# _327_/Q 0.00116f
C14572 _306_/S VPWR 1.9f
C14573 _307_/X _231_/a_79_n19# 5.29e-19
C14574 _194_/X VGND 0.828f
C14575 _162_/A _160_/A 0.0195f
C14576 _309_/a_1108_7# _284_/A 0.0603f
C14577 _158_/Y output40/a_27_7# 3.44e-19
C14578 _277_/Y _301_/a_51_257# 6.24e-20
C14579 _286_/B _201_/a_27_7# 1.83e-19
C14580 _346_/a_956_373# _162_/X 2.41e-19
C14581 _277_/Y clkbuf_1_1_0_clk/a_75_172# 0.0255f
C14582 _317_/a_543_7# _317_/D 0.00306f
C14583 _315_/Q _341_/a_543_7# 1.17e-21
C14584 result[0] _341_/a_193_7# 8.59e-19
C14585 _293_/a_39_257# input1/X 0.0399f
C14586 _308_/S _250_/a_78_159# 5.1e-19
C14587 output11/a_27_7# _279_/Y 0.0344f
C14588 _310_/a_651_373# _310_/D 8.49e-19
C14589 _310_/a_543_7# _310_/Q 2.05e-19
C14590 _329_/a_27_7# _218_/a_250_257# 2.62e-19
C14591 _329_/a_193_7# _218_/a_93_n19# 3.18e-19
C14592 _346_/SET_B _299_/a_215_7# 9.69e-19
C14593 _218_/a_93_n19# _328_/Q 1.13e-20
C14594 _232_/A _242_/B 0.00103f
C14595 _172_/A _146_/C 4.35e-19
C14596 _335_/a_1108_7# _207_/a_27_7# 4.86e-20
C14597 _336_/a_27_7# _336_/a_639_7# -0.0015f
C14598 _327_/a_1283_n19# _216_/X 5.09e-19
C14599 _324_/a_27_7# _248_/B 6.49e-20
C14600 _196_/A _180_/a_111_257# 6.42e-20
C14601 _181_/X _180_/a_29_13# 9.13e-19
C14602 _270_/a_39_257# _217_/A 1.09e-19
C14603 _325_/Q _224_/a_584_7# 0.00353f
C14604 _309_/a_27_7# _306_/S 0.00447f
C14605 _329_/Q _238_/B 0.00474f
C14606 _172_/A _157_/A 0.123f
C14607 _343_/a_543_7# _343_/D 4.36e-19
C14608 _343_/a_1108_7# _185_/A 2.14e-19
C14609 _167_/X VGND 0.27f
C14610 _231_/a_409_7# _144_/A 7.67e-19
C14611 _286_/B _173_/a_226_7# 0.00781f
C14612 _327_/a_1283_n19# _329_/Q 1.62e-19
C14613 _327_/a_1108_7# _320_/Q 5.65e-21
C14614 _187_/a_27_7# _255_/B 0.00262f
C14615 _154_/A _204_/Y 0.0109f
C14616 _327_/a_193_7# _327_/a_1108_7# -0.00817f
C14617 _255_/B _315_/D 0.135f
C14618 _248_/A _347_/a_27_7# 1.61e-20
C14619 _255_/a_112_257# VGND -1.96e-19
C14620 _157_/A _232_/X 9.54e-25
C14621 _318_/Q _317_/a_1283_n19# 8.4e-19
C14622 result[3] _317_/a_761_249# 2.01e-19
C14623 _340_/a_27_7# _340_/CLK 0.26f
C14624 _323_/a_805_7# cal 4.57e-19
C14625 _275_/Y _216_/A 0.00704f
C14626 _333_/D _332_/Q 7.95e-20
C14627 _337_/Q _254_/B 1.07f
C14628 _341_/a_27_7# _341_/D 0.149f
C14629 _315_/Q _316_/a_1283_n19# 1.08e-20
C14630 _294_/A VPWR 0.475f
C14631 _305_/a_505_n19# cal 1.88e-20
C14632 _329_/a_448_7# _330_/Q 0.00171f
C14633 _161_/Y _174_/a_27_257# 0.0115f
C14634 repeater43/X _330_/a_1462_7# 7.65e-19
C14635 _331_/D _331_/a_448_7# 0.0214f
C14636 _169_/B _169_/Y 0.00398f
C14637 _332_/a_193_7# _332_/Q 7.29e-19
C14638 _332_/a_27_7# _333_/Q 0.0134f
C14639 _343_/a_1283_n19# _342_/Q 9.83e-20
C14640 _331_/a_543_7# _330_/a_1283_n19# 0.00122f
C14641 _197_/X _339_/D 0.233f
C14642 _326_/a_27_7# _326_/a_448_7# -0.00656f
C14643 _326_/a_193_7# _326_/a_1108_7# -0.0069f
C14644 _162_/X _313_/a_543_7# 2.08e-20
C14645 _305_/a_505_n19# _197_/a_27_7# 0.00143f
C14646 _328_/a_1283_n19# _320_/Q 0.00141f
C14647 _328_/a_193_7# _238_/B 7.43e-20
C14648 _328_/a_543_7# _329_/Q 0.0406f
C14649 _330_/a_639_7# _212_/X 7.16e-20
C14650 clkbuf_2_1_0_clk/A _336_/a_193_7# 1.18e-21
C14651 repeater43/X _333_/a_1270_373# -2.06e-19
C14652 _329_/a_1108_7# VPWR 0.0125f
C14653 _329_/a_543_7# VGND -0.00247f
C14654 _338_/a_27_7# _338_/D 0.485f
C14655 _327_/D VPWR 0.0943f
C14656 _308_/a_218_7# _306_/S 5.54e-19
C14657 _281_/Y _330_/D 0.0709f
C14658 _296_/a_109_7# VGND -9.03e-19
C14659 _344_/a_27_7# _344_/Q 0.00224f
C14660 _341_/a_761_249# _248_/A 0.00886f
C14661 _306_/a_76_159# _306_/S 0.0511f
C14662 _342_/a_761_249# cal 4.92e-19
C14663 output23/a_27_7# _269_/A 0.0045f
C14664 _294_/A _309_/a_27_7# 0.151f
C14665 _343_/CLK _177_/a_27_7# 3.56e-21
C14666 _146_/C _244_/B 0.00668f
C14667 _172_/A _260_/A 0.447f
C14668 _162_/X _156_/a_121_257# 0.00131f
C14669 _341_/Q _298_/A 1.1f
C14670 _322_/a_805_7# result[6] 4.25e-19
C14671 _332_/a_448_7# _340_/CLK 1.82e-21
C14672 _333_/a_805_7# _207_/C 2.96e-19
C14673 _332_/a_1108_7# _332_/D 1.31e-19
C14674 _301_/a_240_7# _347_/Q 0.00113f
C14675 _344_/a_652_n19# _267_/A 1.33e-21
C14676 _162_/X _304_/S 0.00495f
C14677 _340_/a_193_7# _346_/SET_B 0.0206f
C14678 _182_/a_297_257# _225_/X 0.00562f
C14679 _182_/a_79_n19# _150_/C 0.00364f
C14680 _200_/a_250_257# _340_/CLK 7.75e-21
C14681 _328_/a_193_7# _328_/a_543_7# -0.0102f
C14682 _347_/a_651_373# _347_/D 0.00135f
C14683 _317_/Q _330_/Q 4.61e-19
C14684 _329_/D _330_/D 0.0131f
C14685 _164_/A _172_/Y 3.74e-20
C14686 _283_/A VPWR 1.33f
C14687 clkbuf_2_3_0_clk/a_75_172# clkbuf_2_1_0_clk/A 0.00167f
C14688 _314_/a_193_7# _225_/B 1.91e-19
C14689 _292_/A _163_/a_78_159# 0.00946f
C14690 _277_/A _277_/Y 0.0208f
C14691 _216_/X _248_/A 0.00778f
C14692 _339_/Q _254_/B 5.58e-20
C14693 _327_/a_1283_n19# _274_/a_39_257# 2.15e-19
C14694 _205_/a_382_257# VPWR -1.79e-19
C14695 _271_/A _185_/A 0.017f
C14696 _316_/a_543_7# _248_/A 0.00309f
C14697 _288_/A _267_/B 0.319f
C14698 clkbuf_2_1_0_clk/A _199_/a_256_7# 0.00126f
C14699 _216_/a_27_7# _325_/D 2.42e-21
C14700 _169_/Y _170_/a_226_7# 0.0184f
C14701 _254_/A _299_/a_78_159# 3.65e-21
C14702 _325_/Q _315_/D 4.28e-20
C14703 _163_/a_78_159# _160_/A 0.00587f
C14704 _343_/a_193_7# _175_/Y 0.0148f
C14705 _342_/D _145_/A 3.63e-20
C14706 _270_/a_121_257# VGND -4.17e-19
C14707 _254_/B _202_/a_256_7# 0.00429f
C14708 _216_/X _331_/CLK 0.0171f
C14709 _342_/a_193_7# _286_/Y 0.00744f
C14710 output34/a_27_7# _273_/Y 0.0019f
C14711 _333_/a_448_7# _192_/B 9.1e-20
C14712 _333_/a_1270_373# _191_/B 1.45e-19
C14713 _230_/a_27_7# _318_/a_1283_n19# 0.00465f
C14714 result[0] _341_/a_1462_7# 2.78e-20
C14715 _239_/a_113_257# _232_/X 0.00328f
C14716 _331_/Q _331_/a_1283_n19# 0.0469f
C14717 _308_/S _250_/X 0.00124f
C14718 _287_/a_39_257# _267_/B 0.0441f
C14719 _316_/a_543_7# _331_/CLK 3.51e-20
C14720 _316_/a_761_249# _316_/D 5.8e-19
C14721 _344_/Q _171_/a_215_7# 0.0026f
C14722 _294_/A _306_/a_76_159# 0.0472f
C14723 output36/a_27_7# output37/a_27_7# 6.12e-19
C14724 clkbuf_0_clk/X _330_/a_761_249# 5.43e-19
C14725 clkbuf_2_3_0_clk/A _312_/D 6.85e-20
C14726 _311_/a_27_7# clkc 6.57e-22
C14727 input3/a_27_7# _227_/A 0.0131f
C14728 _294_/Y _311_/a_1108_7# 1.3e-20
C14729 _301_/a_51_257# VGND 0.0509f
C14730 _301_/a_512_257# VPWR 2.15e-20
C14731 _273_/A _162_/A 0.129f
C14732 _320_/Q _316_/D 0.031f
C14733 _329_/Q _331_/CLK 0.00215f
C14734 _194_/A _313_/a_27_7# 1.48e-22
C14735 _248_/B VPWR 3.09f
C14736 _346_/SET_B _347_/a_1270_373# -3.58e-20
C14737 _181_/a_27_7# _284_/A 0.00303f
C14738 _258_/a_76_159# _216_/A 4.57e-20
C14739 clkbuf_1_1_0_clk/a_75_172# VGND 0.0706f
C14740 _326_/a_761_249# _248_/A 1.11e-19
C14741 _273_/A _216_/X 0.0332f
C14742 _334_/a_193_7# _334_/a_543_7# -0.0231f
C14743 clk _333_/a_27_7# 7.86e-21
C14744 _321_/a_543_7# _321_/Q 0.0363f
C14745 _327_/a_761_249# _331_/CLK 0.0194f
C14746 _260_/A _203_/a_80_n19# 1.16e-19
C14747 _208_/a_78_159# _332_/Q 0.00803f
C14748 _208_/a_292_257# _207_/X 3.24e-19
C14749 _328_/Q _328_/D 2.48e-19
C14750 _301_/a_240_7# _297_/B 2.97e-20
C14751 _338_/a_27_7# _337_/a_1108_7# 2.42e-22
C14752 _338_/a_193_7# _337_/a_1283_n19# 7.59e-20
C14753 _338_/a_1108_7# _337_/a_27_7# 3.41e-22
C14754 _338_/a_761_249# _337_/a_543_7# 4.05e-19
C14755 _338_/a_543_7# _337_/a_761_249# 6.57e-19
C14756 _319_/Q output19/a_27_7# 2.21e-19
C14757 _273_/A _329_/Q 1.3e-20
C14758 _326_/a_761_249# _331_/CLK 3.26e-20
C14759 _326_/a_27_7# _236_/B 1.61e-19
C14760 _258_/S _313_/a_27_7# 1.26e-19
C14761 _341_/a_27_7# _343_/CLK 0.0294f
C14762 _286_/B _313_/a_651_373# 0.00112f
C14763 _314_/a_193_7# _314_/a_543_7# 3.55e-33
C14764 _172_/A _251_/a_79_n19# 0.0173f
C14765 _311_/a_193_7# _310_/a_761_249# 8.57e-22
C14766 _311_/a_761_249# _310_/a_193_7# 1.64e-21
C14767 _321_/a_193_7# VPWR 0.0334f
C14768 _338_/a_27_7# _343_/CLK 6.76e-20
C14769 _254_/Y VPWR 1.61f
C14770 repeater43/X _298_/X 0.00976f
C14771 _325_/a_193_7# _223_/a_250_257# 1.32e-19
C14772 _341_/a_1217_7# _341_/D 8.48e-19
C14773 _234_/B _318_/a_27_7# 8.66e-19
C14774 _326_/a_761_249# _273_/A 6.54e-20
C14775 _321_/a_193_7# _318_/a_543_7# 6.89e-20
C14776 _321_/a_27_7# _318_/a_1283_n19# 7.61e-21
C14777 rstn ctln[0] 0.0526f
C14778 _227_/A _153_/A 3.43e-19
C14779 _332_/a_1217_7# _333_/Q 2.37e-19
C14780 trim[4] _162_/A 0.00457f
C14781 _340_/a_761_249# _337_/a_1108_7# 1.64e-19
C14782 _340_/a_543_7# _337_/a_1283_n19# 4.09e-19
C14783 _340_/a_1283_n19# _337_/a_543_7# 4.09e-19
C14784 _340_/a_1108_7# _337_/a_761_249# 1.64e-19
C14785 _210_/a_27_7# VGND 0.0613f
C14786 _326_/a_27_7# _326_/D 0.0456f
C14787 _192_/a_68_257# _192_/B 0.00553f
C14788 result[2] _246_/B 5.9e-20
C14789 _286_/B _157_/a_27_7# 0.00113f
C14790 _279_/Y _337_/a_27_7# 1.12e-21
C14791 _338_/a_651_373# _338_/Q 3.34e-20
C14792 _344_/a_27_7# _306_/S 5.27e-20
C14793 _238_/B _319_/a_543_7# 0.00299f
C14794 _310_/a_1108_7# VGND 0.00399f
C14795 _310_/a_651_373# VPWR 0.0114f
C14796 repeater43/X _332_/a_543_7# 2.05e-19
C14797 _344_/a_562_373# _344_/D 3.6e-19
C14798 _343_/CLK _316_/a_193_7# 1.22e-19
C14799 _196_/A _191_/B 0.194f
C14800 _185_/A _323_/a_27_7# 0.0187f
C14801 _297_/A _302_/a_227_7# 0.00833f
C14802 _294_/A _309_/a_1217_7# 8.93e-19
C14803 _193_/Y _311_/D 1.29e-20
C14804 _316_/Q result[2] 0.187f
C14805 clkbuf_2_1_0_clk/A _170_/a_556_7# 0.00149f
C14806 _172_/A _340_/Q 9.79e-21
C14807 _340_/CLK _332_/D 0.0159f
C14808 _190_/a_27_7# _190_/A 0.0471f
C14809 _274_/a_39_257# _248_/A 6.56e-20
C14810 _346_/a_27_7# _346_/SET_B 0.0954f
C14811 _340_/a_1462_7# _346_/SET_B -9.14e-19
C14812 _182_/X _150_/C 0.0707f
C14813 _325_/D _327_/Q 4.3e-20
C14814 _169_/a_109_257# VPWR -0.00183f
C14815 _225_/a_145_35# VPWR -1.45e-19
C14816 _332_/a_1108_7# _207_/C 9.68e-19
C14817 _339_/a_1108_7# _338_/a_27_7# 9.17e-19
C14818 _339_/a_1283_n19# _338_/a_193_7# 0.00184f
C14819 _271_/A _242_/A 0.0152f
C14820 _344_/a_193_7# _165_/X 2.65e-20
C14821 _271_/A _335_/Q 0.00288f
C14822 _256_/a_209_257# _192_/B 0.00288f
C14823 repeater43/a_27_7# _334_/a_27_7# 0.00579f
C14824 _234_/B _246_/B 2.58e-21
C14825 _198_/a_93_n19# _306_/S 0.00137f
C14826 _315_/D _326_/Q 1.07e-20
C14827 _335_/a_27_7# _335_/Q 0.00397f
C14828 _341_/Q _304_/X 4.59e-21
C14829 _191_/B _298_/X 4.56e-21
C14830 _243_/a_113_257# VGND 0.00287f
C14831 _175_/Y VGND 0.405f
C14832 _299_/X _170_/a_76_159# 0.00672f
C14833 _327_/a_805_7# _346_/SET_B 0.00126f
C14834 _325_/a_27_7# _304_/a_257_159# 1.71e-20
C14835 clk _162_/X 1.01e-19
C14836 _346_/a_193_7# _346_/a_381_7# -0.00419f
C14837 _308_/S _255_/B 0.277f
C14838 repeater43/X _341_/a_448_7# 2.63e-21
C14839 _271_/A _298_/a_109_7# 2.71e-19
C14840 _236_/a_109_257# _248_/A 1.03e-19
C14841 output15/a_27_7# output28/a_27_7# 4.36e-21
C14842 _172_/A _165_/X 0.00559f
C14843 _343_/a_1462_7# _175_/Y 4.63e-19
C14844 _340_/a_193_7# _339_/a_448_7# 9.08e-22
C14845 _254_/Y _306_/a_76_159# 5.65e-20
C14846 _254_/B _336_/D 0.247f
C14847 _342_/a_805_7# sample 1.67e-19
C14848 _190_/A _295_/a_409_7# 0.00172f
C14849 _333_/D _192_/B 5.8e-19
C14850 _242_/A _318_/a_639_7# 0.00111f
C14851 _254_/A _347_/a_1108_7# 0.00194f
C14852 _344_/D _172_/B 9.62e-20
C14853 _279_/Y _339_/a_27_7# 0.00675f
C14854 clkbuf_2_1_0_clk/A _299_/X 0.00701f
C14855 _315_/a_27_7# VPWR 0.0901f
C14856 _284_/a_39_257# _266_/a_113_257# 7.86e-19
C14857 _292_/A clkbuf_2_3_0_clk/A 1.18e-20
C14858 _277_/A VGND 0.667f
C14859 _308_/a_505_n19# _209_/X 2.87e-21
C14860 _329_/a_805_7# _330_/D 4.89e-19
C14861 _182_/a_79_n19# cal 1.26e-19
C14862 _343_/Q _226_/X 0.026f
C14863 _298_/C _225_/X 0.0109f
C14864 _324_/a_543_7# _227_/A 0.0191f
C14865 _336_/a_1108_7# VPWR 0.00566f
C14866 _346_/a_476_7# _273_/A 1e-19
C14867 _336_/a_543_7# VGND -9.95e-19
C14868 _307_/X _298_/C 0.0969f
C14869 _271_/A _322_/D 1.79e-21
C14870 _324_/a_27_7# _324_/a_193_7# -0.299f
C14871 _328_/a_639_7# _346_/SET_B -7.75e-19
C14872 _346_/Q _172_/B 7.47e-21
C14873 input1/X _312_/a_639_7# 9.82e-20
C14874 _315_/D _314_/a_193_7# 0.0226f
C14875 _332_/Q _190_/A 0.954f
C14876 _297_/A _157_/A 0.498f
C14877 _345_/a_27_7# _277_/Y 1.14e-20
C14878 _343_/a_639_7# _298_/A 3.64e-20
C14879 _346_/SET_B _319_/a_27_7# 0.0637f
C14880 clkbuf_0_clk/X _299_/a_78_159# 7.68e-19
C14881 _227_/A _217_/A 2.18e-19
C14882 _292_/A _172_/Y 1.9e-20
C14883 repeater43/X _316_/a_651_373# 0.00383f
C14884 _300_/a_735_7# _299_/X 0.0256f
C14885 _300_/a_383_7# _347_/Q 7.31e-19
C14886 _147_/A _347_/a_1270_373# 1.76e-19
C14887 _172_/A _251_/X 1.91e-19
C14888 _342_/Q _153_/B 4.74e-20
C14889 _321_/a_805_7# VGND -7.97e-19
C14890 _321_/a_1462_7# VPWR 1.53e-19
C14891 _216_/X _217_/X 0.707f
C14892 _344_/Q _147_/Y 4.82e-19
C14893 _196_/A _337_/Q 4.74e-21
C14894 rstn _335_/a_448_7# 0.0154f
C14895 repeater43/X _204_/a_27_257# 7.43e-20
C14896 _338_/a_1217_7# _343_/CLK 4.22e-20
C14897 _322_/a_27_7# _269_/A 0.0264f
C14898 _301_/X _162_/X 0.0965f
C14899 _341_/a_193_7# _145_/A 0.00452f
C14900 repeater43/X _208_/a_493_257# 1.41e-19
C14901 _160_/A _172_/Y 3.14e-21
C14902 _325_/a_27_7# _325_/D 0.484f
C14903 _329_/a_1283_n19# _232_/X 6.54e-19
C14904 _238_/B _327_/Q 2.68e-20
C14905 _329_/Q _217_/X 0.0841f
C14906 _291_/a_121_257# VGND -4.61e-19
C14907 comp _285_/Y 0.0198f
C14908 _327_/a_761_249# _217_/X 0.00164f
C14909 _327_/a_1283_n19# _327_/Q 0.0257f
C14910 _327_/a_543_7# _212_/X 0.00348f
C14911 _326_/a_448_7# repeater43/X 0.0337f
C14912 _275_/Y _310_/a_639_7# 9.32e-19
C14913 _326_/a_27_7# _331_/a_193_7# 0.00113f
C14914 _326_/a_193_7# _331_/a_27_7# 1.71e-20
C14915 _346_/SET_B _338_/Q 0.01f
C14916 _207_/C _204_/a_277_7# 0.0382f
C14917 ctln[2] _292_/A 7.06e-20
C14918 clkbuf_2_2_0_clk/a_75_172# _340_/CLK 0.0378f
C14919 _275_/A _346_/SET_B 0.0106f
C14920 _326_/a_761_249# _217_/X 0.0191f
C14921 _326_/a_1283_n19# _327_/Q 6.04e-20
C14922 _281_/A _330_/a_651_373# 3.42e-19
C14923 _199_/a_584_7# VGND 6.01e-19
C14924 input4/X _340_/CLK 1.28e-19
C14925 _188_/a_218_7# _341_/D 5.9e-19
C14926 _345_/a_193_7# _345_/a_652_n19# -5.22e-20
C14927 _296_/Y _216_/X 3.57e-19
C14928 _255_/a_30_13# _254_/B 4.85e-20
C14929 _313_/Q _193_/Y 7.97e-20
C14930 _297_/A _260_/A 5.87e-21
C14931 _306_/X _306_/S 0.666f
C14932 _334_/Q _204_/a_27_257# 0.114f
C14933 _300_/a_27_257# VPWR 0.019f
C14934 _342_/a_193_7# _269_/A 0.0138f
C14935 output12/a_27_7# _333_/a_1283_n19# 1.49e-20
C14936 _281_/Y _333_/a_27_7# 1.14e-20
C14937 _328_/a_761_249# _212_/X 7.46e-19
C14938 _328_/a_193_7# _217_/X 0.0169f
C14939 ctlp[7] result[7] 0.0274f
C14940 _341_/Q VGND 0.329f
C14941 _344_/a_27_7# _301_/a_512_257# 1.6e-21
C14942 _284_/a_39_257# VPWR 0.0411f
C14943 _298_/B VPWR 0.855f
C14944 _346_/a_586_7# _346_/SET_B 0.00237f
C14945 _211_/a_27_257# _283_/A 0.062f
C14946 _198_/a_93_n19# _283_/A 2.69e-22
C14947 clkbuf_0_clk/X _181_/X 4.21e-20
C14948 result[5] _234_/B 9.44e-20
C14949 _325_/a_1270_373# _181_/X 6.96e-20
C14950 _342_/Q _181_/a_27_7# 0.00256f
C14951 _294_/Y _161_/Y 3.07e-19
C14952 _300_/a_383_7# _297_/B 2.96e-21
C14953 _194_/a_27_7# VPWR 0.0677f
C14954 _340_/CLK _313_/a_1283_n19# 5.21e-21
C14955 output33/a_27_7# _312_/a_1108_7# 6.32e-20
C14956 input4/X _334_/a_651_373# 2.57e-19
C14957 repeater43/X _334_/a_1108_7# -0.0181f
C14958 _229_/a_76_159# _226_/X 0.0146f
C14959 _309_/a_193_7# _310_/D 1.68e-19
C14960 _326_/a_193_7# _217_/a_27_7# 0.00473f
C14961 _232_/a_27_7# _242_/A 0.023f
C14962 _232_/X _230_/a_27_7# 6.91e-21
C14963 result[1] _315_/a_193_7# 3.49e-19
C14964 _147_/A _295_/a_79_n19# 1.46e-19
C14965 _146_/C _177_/A 0.167f
C14966 _335_/D _205_/a_79_n19# 0.00206f
C14967 _259_/a_199_7# _339_/Q 0.00146f
C14968 _157_/A _304_/a_257_159# 1.97e-21
C14969 _342_/a_193_7# _343_/D 3.21e-19
C14970 _347_/Q _346_/D 0.0137f
C14971 clkbuf_0_clk/a_110_7# _216_/X 2.02e-19
C14972 _255_/X _305_/a_76_159# 5.28e-19
C14973 _331_/D clkbuf_1_0_0_clk/a_75_172# 1.43e-19
C14974 _239_/a_113_257# _297_/A 1.56e-19
C14975 repeater43/X _341_/D 0.416f
C14976 _333_/a_1108_7# _207_/a_27_7# 1.45e-20
C14977 clkbuf_1_0_0_clk/a_75_172# _330_/a_193_7# 5.93e-20
C14978 _309_/a_1270_373# _265_/B 1.25e-19
C14979 _345_/a_193_7# _160_/X 2.37e-19
C14980 _337_/a_193_7# _337_/a_543_7# -0.0132f
C14981 _344_/a_1602_7# _297_/Y 0.0513f
C14982 _309_/a_27_7# _284_/a_39_257# 2.94e-21
C14983 _215_/A _314_/D 1.24e-19
C14984 _184_/a_76_159# _298_/A 3.79e-21
C14985 _317_/Q _212_/a_27_7# 2.13e-20
C14986 _299_/a_78_159# _286_/Y 0.0507f
C14987 _237_/a_113_257# clkbuf_0_clk/X 0.0477f
C14988 _340_/a_193_7# _339_/D 0.0165f
C14989 _290_/A _289_/a_39_257# 0.00687f
C14990 _163_/a_215_7# _158_/Y 0.0172f
C14991 _232_/X _232_/A 0.0448f
C14992 _242_/B VPWR 0.84f
C14993 _313_/D _257_/a_79_159# 3.01e-19
C14994 _315_/a_639_7# VGND 2.71e-19
C14995 _315_/a_1217_7# VPWR 1.42e-19
C14996 _183_/a_27_7# _298_/C 4.48e-19
C14997 _181_/X input1/X 0.00572f
C14998 _182_/X cal 0.00704f
C14999 clk _298_/C 0.00831f
C15000 _274_/a_39_257# _217_/X 0.00177f
C15001 _324_/a_193_7# VPWR -0.0762f
C15002 _294_/A _306_/X 0.0134f
C15003 _339_/a_543_7# _332_/Q 7.26e-21
C15004 _342_/a_761_249# _342_/Q 2.48e-19
C15005 _321_/Q _217_/A 1.61e-20
C15006 _330_/Q _304_/X 0.043f
C15007 _346_/SET_B _345_/D 0.0303f
C15008 _262_/a_113_257# VPWR 0.0744f
C15009 _346_/a_1032_373# clkbuf_2_3_0_clk/A 0.00688f
C15010 _326_/a_27_7# _325_/a_1283_n19# 7.57e-21
C15011 _334_/a_1108_7# _334_/Q 7.95e-19
C15012 _318_/a_543_7# _242_/B 1.95e-19
C15013 _318_/a_193_7# _318_/D 0.0515f
C15014 _315_/D _314_/a_1462_7# 4.32e-19
C15015 output31/a_27_7# trim[0] 0.00764f
C15016 _314_/a_1270_373# VPWR 1.09e-19
C15017 _314_/a_448_7# VGND -0.00611f
C15018 _346_/SET_B _319_/a_1217_7# -3.08e-19
C15019 _324_/a_543_7# _297_/B 1.58e-20
C15020 _346_/SET_B _313_/a_1108_7# -0.0236f
C15021 clkbuf_2_3_0_clk/A _331_/CLK 0.0449f
C15022 _343_/a_27_7# VPWR 0.064f
C15023 _346_/SET_B _337_/a_639_7# -7.75e-19
C15024 _338_/D _337_/a_805_7# 1.33e-20
C15025 _248_/A _327_/Q 0.0137f
C15026 _306_/S _147_/Y 0.0295f
C15027 _157_/A _347_/a_761_249# 0.00327f
C15028 clk _332_/a_448_7# 5.25e-19
C15029 repeater43/X _236_/B 0.221f
C15030 _230_/a_27_7# _244_/B 5.56e-19
C15031 _324_/a_651_373# _324_/D 8.49e-19
C15032 _258_/S _174_/a_27_257# 1.02e-19
C15033 _311_/D _310_/a_1270_373# 7.93e-21
C15034 _311_/Q _310_/a_1283_n19# 0.00114f
C15035 _314_/a_1108_7# _314_/Q 0.00126f
C15036 _314_/a_639_7# _314_/D 5.51e-19
C15037 _311_/a_1283_n19# _310_/Q 1.57e-20
C15038 repeater42/a_27_7# _324_/a_27_7# 7.8e-21
C15039 _283_/Y _335_/Q 1.54e-19
C15040 rstn _335_/D 0.0311f
C15041 _341_/a_1462_7# _145_/A 2.44e-19
C15042 _322_/a_1217_7# _269_/A 1.14e-19
C15043 _273_/A clkbuf_2_3_0_clk/A 0.00568f
C15044 _293_/a_39_257# _336_/a_193_7# 1.74e-20
C15045 _331_/CLK _327_/Q 0.526f
C15046 _279_/Y _302_/a_539_257# 5.07e-21
C15047 cal valid 0.081f
C15048 _345_/a_652_n19# VPWR 0.0209f
C15049 _345_/a_27_7# VGND 0.0378f
C15050 _314_/D _304_/X 1.17e-19
C15051 _256_/a_209_257# _260_/A 1.48e-19
C15052 _339_/a_1270_373# _340_/CLK 1.74e-20
C15053 _153_/a_487_257# _153_/B 0.00136f
C15054 _254_/A _346_/SET_B 0.232f
C15055 _297_/B _346_/D 0.013f
C15056 _286_/B _267_/A 0.22f
C15057 output31/a_27_7# _311_/Q 3.21e-19
C15058 _323_/a_651_373# _175_/Y 5.12e-22
C15059 repeater43/X _143_/a_27_7# 5.25e-21
C15060 _266_/a_199_7# VPWR -3.89e-19
C15061 _281_/Y _162_/X 0.00817f
C15062 _306_/a_76_159# _194_/a_27_7# 8.91e-21
C15063 _340_/a_1270_373# _337_/Q 3e-20
C15064 input1/X _343_/Q 1.43e-21
C15065 _345_/a_1182_221# _297_/B 7.49e-20
C15066 _341_/a_1283_n19# _146_/C 0.001f
C15067 _261_/A _312_/D 0.0555f
C15068 _238_/a_109_257# _242_/A 0.00282f
C15069 _326_/D repeater43/X 0.175f
C15070 _232_/A _244_/B 0.376f
C15071 _273_/A _327_/Q 0.598f
C15072 _181_/X _286_/Y 0.419f
C15073 _339_/a_27_7# _337_/a_1283_n19# 0.00733f
C15074 _339_/a_1283_n19# _337_/a_27_7# 0.00733f
C15075 _315_/D _279_/A 9e-19
C15076 result[3] _269_/A 0.0168f
C15077 _273_/A _172_/Y 0.342f
C15078 _235_/a_113_257# _246_/B 0.00444f
C15079 _272_/a_39_257# _330_/Q 2.94e-19
C15080 _341_/a_193_7# _324_/Q 1.45e-21
C15081 _166_/Y _162_/X 0.00685f
C15082 _277_/A _320_/a_1108_7# 7.56e-19
C15083 _184_/a_505_n19# _298_/B 6.07e-19
C15084 _222_/a_93_n19# _327_/Q 0.0394f
C15085 _306_/S _333_/a_1108_7# 2.74e-20
C15086 _200_/a_93_n19# cal 0.00987f
C15087 _245_/a_199_7# VPWR -3.55e-19
C15088 _216_/A _263_/B 4.53e-21
C15089 _330_/Q _220_/a_93_n19# 6.99e-22
C15090 _160_/X VPWR 3.15f
C15091 _294_/A _147_/Y 0.16f
C15092 _305_/a_505_n19# _336_/a_27_7# 0.00189f
C15093 _302_/a_77_159# _347_/D 8.67e-20
C15094 _312_/a_27_7# _297_/Y 1.56e-21
C15095 _329_/a_27_7# _331_/Q 0.00827f
C15096 _322_/a_761_249# _322_/D 2.33e-20
C15097 _322_/a_1283_n19# _234_/B 4.17e-20
C15098 _248_/B _227_/a_113_7# 1.37e-19
C15099 _319_/a_543_7# _217_/X 1.48e-21
C15100 _346_/SET_B _309_/D 0.00546f
C15101 _347_/Q _314_/Q 1.2e-19
C15102 _255_/B _231_/a_676_257# 9.16e-19
C15103 _339_/a_639_7# _346_/SET_B -7.75e-19
C15104 _209_/X _154_/a_27_7# 2.37e-21
C15105 _290_/A _312_/a_1462_7# 6.07e-19
C15106 _188_/a_505_n19# _150_/C 0.0119f
C15107 repeater43/X _343_/CLK 0.304f
C15108 _309_/a_1462_7# _310_/D 4.08e-19
C15109 _188_/a_218_334# _307_/X 1.17e-19
C15110 _258_/a_76_159# _336_/a_651_373# 8.53e-19
C15111 _325_/a_27_7# _248_/A 0.0194f
C15112 _192_/B _190_/A 0.239f
C15113 _166_/Y _299_/a_493_257# 2.2e-19
C15114 _209_/X _179_/a_27_7# 0.00141f
C15115 _172_/A _336_/a_1283_n19# 1.37e-21
C15116 _324_/Q _316_/a_761_249# 1.31e-19
C15117 _313_/a_193_7# _313_/a_448_7# -0.00779f
C15118 _290_/A _287_/a_121_257# 1.45e-20
C15119 _320_/Q output26/a_27_7# 1.38e-19
C15120 _325_/a_27_7# _331_/CLK 0.04f
C15121 _196_/A _336_/D 7.8e-19
C15122 _330_/Q VGND 1.57f
C15123 _145_/A _180_/a_183_257# 0.00107f
C15124 _188_/S _298_/A 0.712f
C15125 _320_/a_27_7# clkbuf_2_1_0_clk/A 4.13e-19
C15126 _163_/a_215_7# _160_/a_27_7# 1.35e-19
C15127 _332_/a_27_7# _207_/a_27_7# 7.82e-19
C15128 repeater43/a_27_7# _323_/Q 7.83e-20
C15129 _317_/a_1108_7# _248_/A 2.67e-20
C15130 _285_/A _310_/D 0.00769f
C15131 _327_/a_651_373# clkbuf_0_clk/X 0.00177f
C15132 _306_/X _254_/Y 6.37e-20
C15133 _297_/a_27_257# _347_/a_1108_7# 1.39e-19
C15134 _343_/a_1108_7# _271_/A 1.83e-20
C15135 _322_/Q _269_/A 1.56e-20
C15136 _273_/A _325_/a_27_7# 1.09e-19
C15137 VPWR ctln[0] 0.202f
C15138 _269_/Y VGND 0.442f
C15139 _326_/a_193_7# _324_/Q 1.48e-22
C15140 _165_/X _164_/A 8.39e-19
C15141 output21/a_27_7# clkbuf_1_0_0_clk/a_75_172# 2.45e-20
C15142 _324_/a_1462_7# VPWR 7.79e-20
C15143 _324_/a_805_7# VGND -5.41e-19
C15144 _254_/A _313_/a_761_249# 0.00142f
C15145 _313_/a_27_7# _157_/a_27_7# 0.00644f
C15146 _248_/a_109_257# _248_/B 7.13e-19
C15147 _317_/a_1283_n19# _316_/D 5.19e-21
C15148 _317_/a_1108_7# _331_/CLK 2.11e-21
C15149 _338_/a_27_7# _195_/a_109_257# 4.99e-20
C15150 _338_/a_193_7# _195_/a_27_257# 4.22e-19
C15151 _343_/CLK _334_/Q 0.00644f
C15152 cal _229_/a_226_7# 0.00126f
C15153 input1/X _229_/a_76_159# 0.00322f
C15154 _232_/A _241_/a_113_257# 1.93e-19
C15155 _314_/D VGND 0.45f
C15156 _179_/a_27_7# _209_/a_109_257# 6.34e-20
C15157 clkbuf_2_3_0_clk/A _267_/a_109_257# 9.31e-19
C15158 _318_/a_1283_n19# VPWR 0.0469f
C15159 _318_/a_761_249# VGND 0.00894f
C15160 _341_/a_193_7# _228_/A 5.56e-19
C15161 _343_/a_639_7# VGND 4.97e-19
C15162 _343_/a_1217_7# VPWR 7.83e-20
C15163 _286_/B _194_/X 0.00437f
C15164 _338_/D _337_/Q 1.61e-20
C15165 _338_/Q _337_/D 2.67e-20
C15166 _325_/a_27_7# _222_/a_93_n19# 2.19e-19
C15167 clk _332_/D 4.43e-19
C15168 _273_/A _317_/a_1108_7# 1.48e-20
C15169 _297_/A _251_/X 0.0293f
C15170 _297_/B _314_/Q 0.0228f
C15171 repeater42/a_27_7# VPWR 0.143f
C15172 _273_/A trimb[2] 0.0252f
C15173 _318_/a_193_7# _318_/a_448_7# -0.00482f
C15174 _225_/X _207_/C 4.39e-19
C15175 _309_/a_193_7# VPWR 0.0331f
C15176 _306_/a_76_159# _160_/X 6.95e-22
C15177 _313_/a_1108_7# _147_/A 0.0417f
C15178 _341_/a_651_373# _286_/Y 8.49e-19
C15179 _343_/CLK _191_/B 0.00695f
C15180 _345_/a_1056_7# VPWR 4.32e-19
C15181 _172_/A _310_/D 0.00116f
C15182 _286_/a_113_7# _306_/S 3.09e-20
C15183 _304_/a_79_n19# _306_/S 1.35e-19
C15184 output11/a_27_7# _195_/a_27_257# 3.91e-21
C15185 _256_/a_80_n19# _306_/S 2.06e-20
C15186 _292_/A _261_/A 4.08e-20
C15187 _336_/a_761_249# _254_/B 4.87e-20
C15188 clk _334_/a_1270_373# 9.84e-20
C15189 _320_/Q _281_/A 0.0469f
C15190 _167_/X _286_/B 9.24e-19
C15191 repeater43/X _331_/a_193_7# 0.0131f
C15192 _254_/A _147_/A 0.0142f
C15193 _316_/a_761_249# _228_/A 2.35e-21
C15194 _283_/A _333_/a_1108_7# 0.0395f
C15195 _178_/a_27_7# _192_/B 1.92e-19
C15196 _216_/A _194_/A 3.29e-21
C15197 _229_/a_76_159# _286_/Y 1.78e-19
C15198 clkbuf_2_1_0_clk/a_75_172# VGND 0.0649f
C15199 _309_/a_27_7# _309_/a_193_7# -0.332f
C15200 _279_/Y _267_/A 2.23e-20
C15201 _255_/a_112_257# _286_/B 9.86e-19
C15202 _255_/a_30_13# _196_/A 2.96e-20
C15203 _258_/a_505_n19# _215_/A 4.31e-20
C15204 _304_/S _150_/C 0.0781f
C15205 cal _340_/CLK 0.00847f
C15206 _326_/a_193_7# _281_/A 7.55e-21
C15207 _294_/Y _263_/B 3.06e-19
C15208 output23/a_27_7# _316_/Q 0.0309f
C15209 _281_/Y _298_/C 6.98e-22
C15210 _254_/Y _147_/Y 0.43f
C15211 _327_/Q _217_/X 0.949f
C15212 _277_/Y _311_/D 0.376f
C15213 clkbuf_0_clk/X _346_/SET_B 0.24f
C15214 _333_/a_27_7# _335_/Q 0.002f
C15215 _197_/a_27_7# _340_/CLK 0.0132f
C15216 _258_/S _216_/A 2.78e-20
C15217 _308_/a_535_334# VGND 4.33e-19
C15218 _308_/a_439_7# VPWR -4.69e-19
C15219 _265_/B _172_/B 8.1e-20
C15220 _306_/S _332_/a_27_7# 4.17e-21
C15221 _343_/a_1283_n19# _323_/a_193_7# 5.86e-19
C15222 _343_/a_761_249# _323_/a_543_7# 8.5e-20
C15223 _343_/a_543_7# _323_/a_761_249# 7.14e-21
C15224 _343_/a_1108_7# _323_/a_27_7# 1.05e-19
C15225 _306_/a_505_n19# VPWR 0.0639f
C15226 _288_/A _297_/Y 1.3f
C15227 _328_/a_27_7# _281_/A 9.17e-21
C15228 _339_/Q _338_/D 0.0317f
C15229 _180_/a_29_13# _150_/a_27_7# 5.79e-20
C15230 _188_/S _215_/A 4.33e-19
C15231 _181_/X _328_/Q 7.22e-21
C15232 trim[2] _312_/Q 0.00254f
C15233 _147_/A _226_/X 0.00233f
C15234 _225_/X _150_/C 0.134f
C15235 _317_/Q _223_/a_93_n19# 1.07e-19
C15236 _146_/C _331_/CLK 5.37e-22
C15237 _311_/a_1270_373# VPWR 1.32e-19
C15238 _307_/X _150_/C 0.0875f
C15239 _311_/a_448_7# VGND -0.00652f
C15240 _285_/A _345_/a_193_7# 1.81e-20
C15241 _162_/X _297_/Y 0.0701f
C15242 _313_/D _336_/a_639_7# 5.63e-20
C15243 _306_/X _336_/a_1108_7# 1.25e-20
C15244 _181_/X _296_/a_295_257# 3.47e-19
C15245 _287_/a_39_257# _297_/Y 8.35e-20
C15246 result[1] VGND 0.131f
C15247 _308_/X _227_/A 0.0227f
C15248 _149_/A _226_/X 0.111f
C15249 _346_/SET_B _202_/a_250_257# 0.00287f
C15250 _309_/D _147_/A 7.79e-20
C15251 _337_/Q _313_/a_193_7# 2.58e-21
C15252 _304_/a_257_159# _251_/X 1.57e-21
C15253 _337_/a_1108_7# _337_/Q 0.0565f
C15254 _345_/a_193_7# _344_/a_193_7# 7.32e-19
C15255 _216_/X _221_/a_346_7# 1.68e-19
C15256 _157_/A _190_/A 9.42e-22
C15257 _288_/A _310_/a_193_7# 3.49e-20
C15258 output32/a_27_7# _310_/a_1108_7# 9.48e-20
C15259 _279_/Y _221_/a_93_n19# 5.71e-20
C15260 _335_/a_1283_n19# VGND -8.38e-19
C15261 _335_/a_448_7# VPWR -0.00208f
C15262 _197_/X _336_/a_639_7# 2.93e-19
C15263 result[0] sample 0.0571f
C15264 _184_/a_218_334# VPWR -7.6e-20
C15265 _184_/a_76_159# VGND 0.00795f
C15266 input1/X _346_/SET_B 0.154f
C15267 _309_/a_27_7# _306_/a_505_n19# 3.16e-21
C15268 _309_/a_193_7# _306_/a_76_159# 3.5e-20
C15269 _302_/a_77_159# _304_/S 1.85e-19
C15270 _273_/A _157_/A 2.67e-20
C15271 _237_/a_113_257# _328_/Q 0.0057f
C15272 _326_/a_193_7# _216_/A 7.42e-20
C15273 _338_/a_27_7# _340_/D 0.0012f
C15274 _338_/a_1108_7# _194_/X 0.00563f
C15275 _345_/a_193_7# _172_/A 1.86e-19
C15276 input4/X clk 0.0208f
C15277 _219_/a_93_n19# _319_/a_193_7# 6.71e-20
C15278 _325_/a_1283_n19# repeater43/X 0.00575f
C15279 _188_/a_76_159# input1/X 1.38e-22
C15280 _209_/X _333_/a_761_249# 3.39e-19
C15281 _317_/a_27_7# _317_/a_193_7# -0.031f
C15282 _324_/Q _180_/a_183_257# 2.13e-19
C15283 _302_/a_227_257# _147_/A 3.88e-19
C15284 _182_/a_79_n19# _204_/Y 5.91e-22
C15285 _325_/a_193_7# _212_/X 5.95e-19
C15286 _325_/a_27_7# _217_/X 0.0101f
C15287 _325_/a_761_249# _327_/Q 7.82e-20
C15288 _275_/Y _309_/a_543_7# 0.0049f
C15289 _344_/a_27_7# _160_/X 7.85e-20
C15290 _304_/a_79_n19# _283_/A 0.00275f
C15291 _320_/a_193_7# _220_/a_250_257# 1.8e-19
C15292 clk _207_/C 0.0184f
C15293 _212_/a_27_7# _304_/X 0.0418f
C15294 repeater43/X _317_/a_639_7# 0.0048f
C15295 _309_/a_1462_7# VPWR 1.16e-19
C15296 _309_/a_805_7# VGND -7.97e-19
C15297 _340_/a_761_249# _340_/D 6.55e-19
C15298 _340_/a_1283_n19# _193_/Y 1.75e-19
C15299 _227_/A _203_/a_209_7# 2.49e-20
C15300 _258_/a_505_n19# _300_/Y 1.51e-21
C15301 _286_/B _301_/a_51_257# 8.38e-20
C15302 _296_/Y _192_/B 1.18e-20
C15303 _227_/A _254_/B 0.0774f
C15304 _260_/B _306_/S 0.158f
C15305 _336_/a_1108_7# _147_/Y 0.0422f
C15306 _346_/SET_B _286_/Y 0.0125f
C15307 _260_/A _190_/A 0.0108f
C15308 _346_/SET_B _297_/a_27_257# 0.013f
C15309 ctln[5] ctln[6] 0.00244f
C15310 _219_/a_584_7# _346_/SET_B 6.32e-19
C15311 output13/a_27_7# _269_/Y 1.57e-19
C15312 _283_/Y output6/a_27_7# 8.91e-19
C15313 _146_/C _145_/a_113_7# 1.39e-19
C15314 _340_/CLK _284_/A 0.0867f
C15315 _271_/A _323_/a_27_7# 7.54e-21
C15316 _321_/a_1270_373# _322_/Q 1.29e-19
C15317 _346_/a_193_7# _346_/Q 8.01e-20
C15318 _284_/A _347_/D 9.79e-21
C15319 output12/a_27_7# _332_/Q 8.3e-19
C15320 _339_/a_1108_7# _337_/Q 1.07e-19
C15321 _269_/A _343_/Q 1.63e-19
C15322 repeater43/X _331_/a_1462_7# 2.97e-19
C15323 _181_/a_27_7# _315_/D 0.0344f
C15324 _307_/a_505_n19# _157_/A 9.69e-21
C15325 _292_/A _165_/X 1.33e-19
C15326 _231_/a_512_7# _298_/A 1.81e-19
C15327 _346_/a_27_7# _319_/Q 2.07e-20
C15328 _285_/A VPWR 0.714f
C15329 _331_/a_193_7# _331_/a_448_7# -0.00297f
C15330 _146_/C _178_/a_27_7# 5.27e-19
C15331 _330_/Q _214_/a_27_257# 0.00425f
C15332 _325_/a_27_7# _296_/Y 1.1e-21
C15333 _183_/a_471_7# _304_/S 1.43e-19
C15334 _304_/a_79_n19# _248_/B 0.0491f
C15335 _188_/a_76_159# _286_/Y 0.0604f
C15336 _342_/Q _182_/X 2.54e-19
C15337 _255_/X _181_/X 3.51e-19
C15338 _313_/Q _215_/A 0.0168f
C15339 _339_/Q _343_/CLK 1.07e-20
C15340 _320_/a_1283_n19# VPWR 0.0187f
C15341 _320_/a_761_249# VGND 0.0236f
C15342 _283_/A _332_/a_27_7# 0.00101f
C15343 _323_/a_448_7# VPWR 0.00417f
C15344 _323_/a_1283_n19# VGND 0.0323f
C15345 _277_/Y _313_/Q 1.5e-20
C15346 output19/a_27_7# _279_/A 0.0375f
C15347 _232_/A _177_/A 0.00644f
C15348 _294_/Y _258_/S 0.489f
C15349 _333_/D _205_/a_79_n19# 2.6e-20
C15350 _189_/a_27_7# _340_/a_193_7# 4.57e-20
C15351 _322_/a_27_7# _318_/a_27_7# 8.76e-19
C15352 clkbuf_0_clk/a_110_7# _192_/B 0.00125f
C15353 input1/X _206_/A 0.0293f
C15354 _344_/a_193_7# VPWR 0.0413f
C15355 result[3] _242_/a_109_257# 2.04e-19
C15356 _320_/a_448_7# _297_/B 0.0138f
C15357 _275_/Y _311_/a_805_7# 1.19e-19
C15358 _343_/D _343_/Q 2.83e-19
C15359 _185_/A _298_/C 0.0173f
C15360 _186_/a_79_n19# _271_/A 0.0148f
C15361 _286_/B _210_/a_27_7# 6.38e-20
C15362 _207_/a_27_7# _333_/Q 0.0129f
C15363 _345_/a_1182_221# _161_/Y 0.0136f
C15364 _183_/a_27_7# _150_/C 0.00212f
C15365 _207_/X _207_/a_181_7# 4.43e-19
C15366 _281_/Y _332_/D 0.00176f
C15367 _344_/a_476_7# _297_/B 1.5e-19
C15368 clkbuf_0_clk/X _147_/A 3.09e-20
C15369 _258_/a_535_334# VPWR -8.41e-19
C15370 _258_/a_505_n19# VGND 0.0583f
C15371 _285_/A _309_/a_27_7# 1.99e-20
C15372 _311_/D VGND 0.0723f
C15373 trimb[1] _285_/Y 0.00356f
C15374 _254_/Y _256_/a_80_n19# 5.34e-21
C15375 _325_/a_27_7# _325_/a_761_249# -0.0166f
C15376 _271_/A _232_/a_27_7# 0.00905f
C15377 _172_/A VPWR 5.53f
C15378 _248_/A _221_/a_250_257# 2.32e-19
C15379 repeater43/X output30/a_27_7# 2.61e-21
C15380 _312_/Q _310_/a_761_249# 5.74e-20
C15381 _346_/Q _173_/a_76_159# 3.66e-20
C15382 _285_/Y VGND 0.138f
C15383 output28/a_27_7# result[7] 0.00704f
C15384 _223_/a_93_n19# _298_/A 5.9e-21
C15385 _211_/a_109_257# VPWR 0.00216f
C15386 _198_/a_250_257# VPWR 0.0215f
C15387 _232_/X VPWR 1.12f
C15388 _222_/a_346_7# _286_/Y 4.05e-20
C15389 _335_/D VPWR 0.138f
C15390 _341_/a_651_373# _269_/A 0.00128f
C15391 _245_/a_113_257# _244_/B 0.0446f
C15392 _188_/S VGND 0.377f
C15393 comp _162_/A 0.227f
C15394 _232_/A _325_/D 3.75e-19
C15395 _267_/A _313_/a_27_7# 5.7e-20
C15396 _343_/a_543_7# _342_/a_1108_7# 3.37e-20
C15397 _343_/a_1283_n19# _342_/a_1283_n19# 5.11e-20
C15398 _343_/a_193_7# _342_/a_651_373# 4.57e-20
C15399 _251_/a_79_n19# _190_/A 2.55e-19
C15400 _338_/a_543_7# _283_/A 3.73e-20
C15401 _319_/Q _319_/a_27_7# 0.00851f
C15402 _339_/a_639_7# _339_/D 1.57e-19
C15403 _339_/a_1108_7# _339_/Q 0.00699f
C15404 _194_/a_27_7# _147_/Y 3.95e-19
C15405 _327_/a_543_7# _327_/D 2.8e-19
C15406 _327_/a_651_373# _328_/Q 1.87e-19
C15407 _273_/A _221_/a_250_257# 0.00854f
C15408 _309_/a_27_7# _172_/A 2.37e-19
C15409 _171_/a_493_257# VGND -3.15e-19
C15410 _313_/a_761_249# _297_/a_27_257# 3.35e-20
C15411 trim[4] _265_/a_109_257# 0.00115f
C15412 _333_/a_543_7# _153_/A 1.54e-21
C15413 _333_/a_193_7# _154_/A 1.61e-19
C15414 cal _225_/X 0.554f
C15415 input1/X _147_/A 0.0109f
C15416 _286_/B _175_/Y 0.0271f
C15417 _212_/a_27_7# VGND 0.0334f
C15418 _216_/A _180_/a_183_257# 2.39e-20
C15419 rstn _332_/a_193_7# 1.6e-19
C15420 _254_/a_109_257# _267_/A 3.99e-19
C15421 _269_/A _229_/a_76_159# 1.5e-20
C15422 input1/X _149_/A 0.0133f
C15423 _340_/a_1108_7# _283_/A 1.86e-21
C15424 cal _267_/B 9.25e-20
C15425 _341_/a_1283_n19# _232_/A 2.86e-21
C15426 trim[0] _311_/a_1108_7# 4.74e-19
C15427 _212_/a_27_7# _318_/a_1108_7# 1.92e-20
C15428 _320_/a_27_7# _328_/D 8.73e-21
C15429 _283_/Y _271_/A 3.09e-20
C15430 _269_/A _316_/a_1270_373# 1.79e-19
C15431 _150_/C _150_/a_109_257# 6.95e-19
C15432 _240_/B _346_/SET_B 0.0013f
C15433 _283_/Y _335_/a_27_7# 0.00213f
C15434 _275_/A _319_/Q 0.0171f
C15435 result[2] _316_/a_193_7# 0.00255f
C15436 _203_/a_80_n19# VPWR 0.0656f
C15437 _286_/B _336_/a_543_7# 0.00525f
C15438 _345_/a_1032_373# _172_/B 0.00363f
C15439 _339_/a_27_7# _195_/a_27_257# 3.22e-21
C15440 _244_/B VPWR 0.803f
C15441 _185_/A _229_/a_489_373# 6.62e-20
C15442 _322_/a_805_7# _321_/Q 3.79e-19
C15443 _306_/S _333_/Q 0.0165f
C15444 _164_/A _310_/D 0.0023f
C15445 _325_/Q _316_/a_27_7# 1.09e-19
C15446 output8/a_27_7# output33/a_27_7# 6.6e-19
C15447 _308_/a_218_334# _308_/X 8.5e-19
C15448 _196_/A _260_/a_27_257# 0.00657f
C15449 _346_/a_796_7# _346_/Q 2.52e-20
C15450 _326_/a_543_7# _283_/A 3.07e-19
C15451 _296_/Y _157_/A 0.0134f
C15452 _311_/a_1108_7# _311_/Q 9.16e-19
C15453 _146_/a_29_271# _146_/C 0.0232f
C15454 _172_/A _306_/a_76_159# 1.09e-19
C15455 _318_/a_193_7# _317_/D 5.61e-20
C15456 _147_/A _286_/Y 5.24e-20
C15457 _322_/a_1270_373# VPWR -1.7e-19
C15458 _330_/Q _330_/a_27_7# 0.00452f
C15459 _147_/A _297_/a_27_257# 0.00905f
C15460 _313_/a_543_7# _284_/A 0.00523f
C15461 _315_/a_543_7# _177_/a_27_7# 3.96e-21
C15462 _298_/C _335_/Q 1.61e-20
C15463 _344_/a_476_7# _275_/Y 0.00223f
C15464 _337_/a_651_373# _284_/A 1.57e-19
C15465 _346_/a_1032_373# _165_/X 0.00674f
C15466 rstn _338_/a_1283_n19# 0.00974f
C15467 _320_/D VPWR 0.0882f
C15468 _323_/D VPWR 0.249f
C15469 _318_/Q _330_/Q 0.00156f
C15470 _302_/a_77_159# _301_/X 0.0279f
C15471 _290_/A _338_/Q 0.0915f
C15472 _149_/A _286_/Y 0.00793f
C15473 _280_/a_68_257# _331_/a_1283_n19# 0.00316f
C15474 _165_/X _331_/CLK 2.27e-20
C15475 _290_/A _275_/A 0.0476f
C15476 _344_/a_796_7# VPWR 4.85e-19
C15477 _255_/B _295_/a_79_n19# 0.0322f
C15478 _329_/a_193_7# _346_/SET_B -0.00409f
C15479 _346_/SET_B _328_/Q 0.386f
C15480 _231_/a_512_7# _304_/X 1.5e-20
C15481 _298_/C _298_/a_109_7# 6.43e-19
C15482 input1/X _337_/D 3.81e-21
C15483 _332_/a_1108_7# _204_/Y 5.56e-20
C15484 _343_/a_805_7# _323_/D 4.47e-19
C15485 _162_/X _170_/a_489_373# 0.0318f
C15486 clkbuf_0_clk/a_110_7# _157_/A 0.00126f
C15487 _250_/a_215_7# _147_/A 0.0722f
C15488 _273_/A _165_/X 0.356f
C15489 _313_/Q VGND 0.459f
C15490 _285_/A _309_/a_1217_7# 2.55e-21
C15491 _326_/a_1283_n19# _232_/A 3.52e-20
C15492 _254_/Y _260_/B 0.0754f
C15493 _194_/X _313_/a_27_7# 2.51e-22
C15494 _304_/S _284_/A 1.29e-20
C15495 _320_/Q _321_/a_543_7# 2.91e-20
C15496 _168_/a_109_257# clkbuf_2_3_0_clk/A 0.00117f
C15497 _337_/a_543_7# _340_/Q 3.02e-20
C15498 _337_/a_1283_n19# _194_/X 6.97e-20
C15499 _337_/a_193_7# _193_/Y 2.67e-19
C15500 _251_/X _248_/A 1.61e-20
C15501 ctln[6] _206_/A 0.00874f
C15502 _318_/Q _318_/a_761_249# 0.0197f
C15503 _324_/a_27_7# _297_/A 0.00888f
C15504 _342_/a_651_373# VGND 0.00286f
C15505 _342_/a_639_7# VPWR 3.84e-19
C15506 _335_/a_1108_7# _335_/D 0.00115f
C15507 _239_/a_113_257# _217_/X 1.47e-19
C15508 _166_/Y _345_/Q 3.52e-20
C15509 _315_/Q _248_/B 0.00883f
C15510 rstn _208_/a_78_159# 2.54e-21
C15511 trim[1] _310_/Q 3.7e-19
C15512 _286_/B _341_/Q 3.81e-19
C15513 _329_/a_1283_n19# _331_/CLK 4.42e-20
C15514 _160_/X _147_/Y 0.315f
C15515 _307_/a_76_159# _306_/S 0.00163f
C15516 _322_/a_27_7# result[5] 0.00303f
C15517 _251_/X _190_/A 2.78e-20
C15518 _319_/Q _319_/a_1217_7# 0.00115f
C15519 _306_/X _309_/a_193_7# 1.3e-21
C15520 _255_/B _180_/a_29_13# 2.54e-19
C15521 _273_/A _251_/X 6.76e-19
C15522 _241_/a_113_257# VPWR 0.0744f
C15523 _257_/a_544_257# _340_/CLK 4.95e-19
C15524 _320_/a_193_7# _320_/a_448_7# -0.00297f
C15525 _304_/X _223_/a_93_n19# 0.0322f
C15526 _267_/B _284_/A 0.0158f
C15527 clk cal 0.00753f
C15528 _312_/a_27_7# _311_/a_761_249# 1.1e-21
C15529 _276_/a_150_257# clkbuf_0_clk/X 0.0013f
C15530 _340_/a_27_7# _336_/Q 1.72e-20
C15531 _341_/a_193_7# _315_/a_761_249# 8.57e-22
C15532 _341_/a_761_249# _315_/a_193_7# 1.3e-21
C15533 _341_/a_761_249# _298_/A 0.0198f
C15534 clkbuf_0_clk/a_110_7# _260_/A 0.00617f
C15535 _319_/Q _254_/A 6.19e-21
C15536 output18/a_27_7# VGND 0.107f
C15537 _345_/a_193_7# _164_/A 4.38e-19
C15538 _344_/a_27_7# _344_/a_193_7# -0.035f
C15539 _290_/A _345_/D 5.11e-20
C15540 _217_/X _221_/a_250_257# 0.00241f
C15541 _230_/a_27_7# _248_/A 0.0541f
C15542 _212_/X _221_/a_256_7# 7.63e-19
C15543 _327_/Q _221_/a_346_7# 3.76e-19
C15544 output35/a_27_7# _297_/Y 5.97e-20
C15545 _233_/a_113_257# VGND -0.00247f
C15546 _320_/a_1217_7# _328_/D 1.74e-20
C15547 _216_/A _313_/a_651_373# 8.49e-19
C15548 _283_/A _333_/Q 0.371f
C15549 _340_/CLK _310_/a_761_249# 5.61e-20
C15550 _196_/A _227_/A 0.103f
C15551 _258_/S _336_/a_651_373# 1.55e-19
C15552 result[2] _316_/a_1462_7# 2.44e-19
C15553 _230_/a_27_7# _331_/CLK 1.44e-20
C15554 _339_/a_193_7# _193_/Y 0.00795f
C15555 _339_/a_761_249# _306_/S 0.00394f
C15556 _294_/A output8/a_27_7# 1.3e-19
C15557 _339_/a_543_7# _340_/Q 0.00328f
C15558 _339_/a_1283_n19# _194_/X 0.0116f
C15559 _298_/C _336_/Q 0.0129f
C15560 _200_/a_250_257# _199_/a_93_n19# 0.00113f
C15561 _312_/a_448_7# VPWR 0.00322f
C15562 _312_/a_1283_n19# VGND 0.0232f
C15563 _299_/X _299_/a_78_159# 0.00758f
C15564 _344_/a_27_7# _172_/A 0.00312f
C15565 _270_/a_121_257# _316_/D 9.54e-19
C15566 _196_/A _314_/a_1108_7# 7.06e-19
C15567 _204_/Y _204_/a_277_7# 0.00269f
C15568 _205_/a_297_7# _332_/Q 5.96e-19
C15569 _240_/B _147_/A 3.48e-21
C15570 _232_/A _248_/A 0.0362f
C15571 _264_/a_113_257# _340_/CLK 0.0144f
C15572 _300_/a_27_257# _347_/a_193_7# 6.64e-22
C15573 _292_/A trimb[0] 4.11e-20
C15574 _316_/Q result[3] 9.87e-19
C15575 _340_/a_1108_7# _336_/a_1108_7# 9.66e-21
C15576 _316_/a_193_7# _315_/a_543_7# 6.61e-19
C15577 _316_/a_761_249# _315_/a_761_249# 1.55e-20
C15578 _316_/a_543_7# _315_/a_193_7# 6.54e-21
C15579 _216_/A _157_/a_27_7# 1.25e-19
C15580 _231_/a_512_7# VGND 0.0491f
C15581 _272_/a_39_257# _223_/a_93_n19# 3.47e-19
C15582 clkbuf_2_3_0_clk/A _193_/Y 4.43e-20
C15583 _346_/SET_B clkc 3.26e-20
C15584 _330_/Q _330_/a_1217_7# 8.51e-21
C15585 _331_/CLK _232_/A 0.293f
C15586 en valid 0.00291f
C15587 _227_/A _298_/X 2.26e-20
C15588 _345_/a_27_7# _286_/B 2.06e-20
C15589 _321_/a_27_7# _248_/A 1.04e-20
C15590 clkbuf_2_1_0_clk/A _338_/a_27_7# 1.88e-19
C15591 clkbuf_2_0_0_clk/a_75_172# _338_/a_1283_n19# 1.67e-20
C15592 cal _150_/a_109_257# 2.07e-19
C15593 _330_/a_805_7# VPWR 2.22e-19
C15594 _330_/a_1270_373# VGND 3.3e-19
C15595 _273_/A _232_/A 1.25e-20
C15596 _343_/a_543_7# _177_/a_27_7# 1.95e-20
C15597 _344_/a_1182_221# _171_/a_78_159# 3.22e-19
C15598 _269_/A _206_/A 0.117f
C15599 _337_/a_761_249# _283_/A 5.66e-20
C15600 _321_/a_27_7# _331_/CLK 0.633f
C15601 _338_/Q _310_/a_27_7# 4.67e-20
C15602 _346_/SET_B _310_/a_543_7# 0.00975f
C15603 _333_/a_448_7# VPWR -0.00164f
C15604 _333_/a_1283_n19# VGND 0.0161f
C15605 _341_/a_1108_7# _341_/Q 1.84e-19
C15606 _294_/Y _158_/Y 2.83e-19
C15607 _297_/A VPWR 0.372f
C15608 _337_/a_1462_7# _193_/Y 3.96e-19
C15609 _315_/Q _315_/a_27_7# 0.0126f
C15610 output22/a_27_7# _315_/a_1283_n19# 0.00124f
C15611 clkbuf_0_clk/a_110_7# _251_/a_79_n19# 3.42e-19
C15612 _343_/a_27_7# _176_/a_27_7# 2.46e-20
C15613 _218_/a_346_7# _331_/Q 0.00328f
C15614 _166_/Y _302_/a_77_159# 6.24e-20
C15615 _322_/Q _246_/B 0.00561f
C15616 _319_/Q _331_/a_1108_7# 8.29e-20
C15617 _198_/a_93_n19# _198_/a_250_257# -6.97e-22
C15618 _309_/a_1108_7# _289_/a_39_257# 3.05e-21
C15619 _292_/A _310_/D 0.879f
C15620 _336_/a_27_7# _340_/CLK 0.00796f
C15621 _258_/S _300_/a_383_7# 2.16e-21
C15622 rstn _190_/A 3.39e-20
C15623 _197_/X _153_/B 0.00912f
C15624 _167_/a_109_257# _345_/Q 8.3e-20
C15625 _185_/A _207_/C 2.09e-19
C15626 _343_/D _206_/A 0.0897f
C15627 _196_/A _347_/Q 1.27e-19
C15628 _223_/a_93_n19# VGND 0.00317f
C15629 _216_/A _317_/a_1283_n19# 2.29e-20
C15630 _223_/a_256_7# VPWR -9.17e-19
C15631 _164_/A VPWR 0.336f
C15632 _160_/A _310_/D 0.0186f
C15633 _324_/a_27_7# _325_/D 0.00271f
C15634 _267_/A _174_/a_27_257# 7.62e-20
C15635 _322_/a_193_7# _322_/a_543_7# -0.0129f
C15636 clk _284_/A 0.0354f
C15637 _164_/Y _297_/B 6.14e-21
C15638 _344_/a_476_7# _161_/Y 3.35e-21
C15639 _258_/a_76_159# _254_/B 8.84e-21
C15640 _320_/D _320_/a_543_7# 5.55e-19
C15641 _255_/X _206_/A 0.00654f
C15642 _345_/Q _297_/Y 1.11e-19
C15643 _332_/a_651_373# _154_/A 3.01e-19
C15644 _192_/a_68_257# VPWR 0.0339f
C15645 _309_/a_27_7# _164_/A 0.00148f
C15646 _330_/D _330_/a_1283_n19# 1.81e-21
C15647 _313_/a_1283_n19# _297_/Y 2.37e-21
C15648 _329_/a_1283_n19# _217_/X 0.00207f
C15649 _329_/a_1108_7# _212_/X 0.00892f
C15650 _212_/X _327_/D 0.00572f
C15651 _343_/D _191_/a_109_257# 1.74e-19
C15652 _225_/a_59_35# _190_/A 0.0135f
C15653 _339_/a_761_249# _283_/A 0.0219f
C15654 _346_/SET_B _336_/a_193_7# 0.0115f
C15655 _216_/X _215_/A 1.48e-19
C15656 _200_/a_346_7# clkbuf_2_1_0_clk/A 7.79e-20
C15657 _283_/A _282_/a_121_257# 7.34e-20
C15658 _275_/Y _312_/a_1270_373# 5.04e-20
C15659 _316_/D _243_/a_113_257# 8.5e-20
C15660 _199_/a_250_257# _340_/CLK 6.41e-21
C15661 _324_/a_1270_373# _181_/X 1.89e-19
C15662 _271_/A _162_/X 1.49e-20
C15663 _292_/A trimb[3] 4.71e-19
C15664 _185_/A _150_/C 1.43e-19
C15665 _312_/D VPWR 0.0967f
C15666 _342_/Q _304_/S 0.0127f
C15667 _196_/A _297_/B 7.5e-20
C15668 ctln[2] output5/a_27_7# 1.42e-19
C15669 _290_/A _162_/a_27_7# 4.25e-21
C15670 _319_/Q clkbuf_0_clk/X 0.923f
C15671 result[0] _341_/Q 3.66e-20
C15672 _300_/Y _347_/a_27_7# 0.0103f
C15673 _160_/X _347_/a_193_7# 0.0013f
C15674 _347_/Q _347_/a_1283_n19# 0.0197f
C15675 _299_/X _347_/a_1108_7# 5.19e-20
C15676 _304_/S _144_/a_27_7# 0.0147f
C15677 _304_/a_257_159# VPWR 0.0714f
C15678 _316_/a_1283_n19# _242_/B 8.46e-21
C15679 _326_/a_805_7# _326_/Q 3.15e-20
C15680 _332_/D _336_/Q 4.14e-21
C15681 _305_/a_505_n19# _197_/X 2.1e-21
C15682 _340_/CLK _225_/B 0.0074f
C15683 _256_/a_209_257# VPWR -0.00511f
C15684 _306_/X _172_/A 2.93e-20
C15685 _296_/Y _251_/X 2.08e-21
C15686 result[2] repeater43/X 0.00574f
C15687 _283_/A _212_/X 0.00908f
C15688 _298_/A _332_/Q 1.22e-19
C15689 _177_/A VPWR 0.448f
C15690 _227_/A _204_/a_27_257# 4.49e-19
C15691 input4/X _335_/Q 3.02e-19
C15692 input1/a_75_172# _194_/X 1.53e-19
C15693 VGND output41/a_27_7# 0.104f
C15694 _255_/X _147_/A 1.4e-19
C15695 _342_/Q _225_/X 1.46e-19
C15696 _145_/A _296_/a_109_7# 6.88e-20
C15697 _279_/Y _314_/a_448_7# 0.00325f
C15698 _317_/Q _327_/Q 4.67e-21
C15699 _307_/X _342_/Q 8.34e-20
C15700 _281_/Y cal 0.00833f
C15701 _345_/a_193_7# _292_/A 2e-19
C15702 _216_/X _304_/X 0.081f
C15703 _342_/a_27_7# _342_/a_448_7# -0.00346f
C15704 _342_/a_193_7# _342_/a_1108_7# 1.42e-32
C15705 _306_/X _198_/a_250_257# 8.57e-21
C15706 _346_/a_193_7# _170_/a_76_159# 1.49e-21
C15707 _321_/D _321_/a_651_373# 2.65e-19
C15708 _333_/a_193_7# _153_/B 1.73e-20
C15709 _338_/D _199_/a_346_7# 6.13e-19
C15710 _273_/A trimb[0] 0.0121f
C15711 _283_/Y _312_/a_27_7# 7.16e-20
C15712 _333_/D VPWR 0.347f
C15713 _294_/Y _160_/a_27_7# 0.00936f
C15714 _157_/A _251_/a_215_7# 0.0364f
C15715 _318_/Q _212_/a_27_7# 0.0326f
C15716 _207_/C _335_/Q 0.0213f
C15717 _327_/a_193_7# _217_/A 6.45e-20
C15718 ctlp[7] _330_/Q 2.54e-19
C15719 _337_/Q _340_/D 2.05e-19
C15720 _315_/Q _315_/a_1217_7# 1.61e-19
C15721 clkbuf_0_clk/a_110_7# _251_/X 0.00213f
C15722 _343_/a_1108_7# _298_/C 5.02e-20
C15723 _343_/a_651_373# _343_/Q 0.00104f
C15724 _346_/a_193_7# clkbuf_2_1_0_clk/A 8.08e-20
C15725 _332_/a_193_7# VPWR -0.0978f
C15726 _315_/D _347_/a_448_7# 0.00163f
C15727 rstn _339_/a_543_7# 9.92e-21
C15728 _275_/Y _164_/Y 1.59e-20
C15729 _232_/A _217_/X 5e-21
C15730 _248_/B _212_/X 6.79e-20
C15731 _347_/a_27_7# VGND -0.082f
C15732 _347_/a_761_249# VPWR 0.00546f
C15733 _325_/a_543_7# _296_/a_109_7# 3.54e-21
C15734 _326_/a_761_249# _304_/X 0.0103f
C15735 _326_/a_193_7# _217_/A 7.13e-19
C15736 repeater43/X _234_/B 0.0162f
C15737 _325_/D VPWR 0.465f
C15738 _308_/a_535_334# _286_/B 4.9e-19
C15739 _308_/a_505_n19# _181_/X 0.00194f
C15740 repeater43/X _321_/a_1283_n19# -0.0071f
C15741 output23/a_27_7# _341_/a_27_7# 1.83e-20
C15742 _336_/a_543_7# _313_/a_27_7# 8.2e-21
C15743 _336_/a_761_249# _313_/a_193_7# 8.05e-21
C15744 _297_/B _347_/a_1283_n19# 0.0133f
C15745 _314_/D _347_/a_543_7# 2.97e-20
C15746 _336_/a_193_7# _313_/a_761_249# 1.72e-20
C15747 _305_/a_439_7# _254_/B 0.00171f
C15748 _250_/a_292_257# _284_/A 2.94e-19
C15749 _267_/B _310_/a_761_249# 0.00725f
C15750 _309_/D _310_/a_27_7# 0.00251f
C15751 output25/a_27_7# _317_/D 3.46e-19
C15752 repeater43/X _153_/a_215_257# 0.00481f
C15753 repeater43/X _209_/X 4.05e-20
C15754 _267_/B _264_/a_113_257# 2.49e-19
C15755 _192_/B _205_/a_297_7# 1.29e-19
C15756 _341_/Q _316_/D 8.1e-20
C15757 _273_/A _310_/D 0.00644f
C15758 _172_/A _147_/Y 0.0563f
C15759 trimb[2] comp 2.27e-20
C15760 _233_/a_199_7# _232_/X 1.41e-19
C15761 _325_/a_193_7# _283_/A 1.73e-20
C15762 _341_/a_1283_n19# VPWR 0.0635f
C15763 _168_/a_397_257# _267_/A 4.46e-21
C15764 _341_/a_761_249# VGND -0.00176f
C15765 _309_/a_1217_7# _164_/A 1.07e-19
C15766 _216_/X _220_/a_93_n19# 0.0394f
C15767 _327_/a_27_7# _218_/a_93_n19# 0.00351f
C15768 _319_/Q _286_/Y 2.41e-19
C15769 _259_/a_199_7# _275_/Y 6.75e-20
C15770 _275_/Y _196_/A 3.29e-20
C15771 _225_/X _204_/Y 6.01e-22
C15772 _338_/a_761_249# VGND 0.00751f
C15773 _338_/a_1283_n19# VPWR 0.00573f
C15774 _150_/C _335_/Q 3.44e-20
C15775 _281_/Y _250_/a_493_257# 2.47e-19
C15776 _346_/SET_B _336_/a_1462_7# -9.14e-19
C15777 _320_/Q _220_/a_250_257# 0.0921f
C15778 _329_/Q _220_/a_93_n19# 0.0568f
C15779 _275_/A output39/a_27_7# 3.76e-19
C15780 ctlp[4] output19/a_27_7# 5.3e-19
C15781 clkbuf_2_1_0_clk/A _319_/a_193_7# 1.43e-20
C15782 trimb[1] _162_/A 0.0941f
C15783 _346_/SET_B _314_/a_1283_n19# 0.0556f
C15784 _339_/Q _340_/D 1.04e-20
C15785 _292_/A VPWR 1.27f
C15786 _315_/a_805_7# _248_/A 9.55e-19
C15787 _216_/A _267_/A 0.0897f
C15788 repeater43/X _209_/a_109_257# 3.13e-19
C15789 _334_/Q _153_/a_215_257# -4.44e-34
C15790 _317_/Q _317_/a_1108_7# 0.00576f
C15791 _336_/a_193_7# _147_/A 5.3e-19
C15792 _230_/a_27_7# _317_/a_651_373# 1.54e-19
C15793 _242_/A _317_/a_193_7# 8.58e-20
C15794 _324_/a_27_7# _248_/A 3.67e-20
C15795 _209_/X _334_/Q 1.63e-19
C15796 _325_/a_193_7# _248_/B 3.12e-21
C15797 _340_/a_448_7# VPWR 0.00267f
C15798 _340_/a_1283_n19# VGND -0.00144f
C15799 _162_/A VGND 0.783f
C15800 _160_/A VPWR 0.236f
C15801 _300_/Y _347_/a_1217_7# 5.17e-19
C15802 trim[4] _310_/D 8.19e-19
C15803 _216_/X VGND 0.686f
C15804 _250_/X _286_/Y 0.0943f
C15805 _290_/A _286_/Y 1.4e-20
C15806 _316_/a_1108_7# VPWR 0.0129f
C15807 _316_/a_543_7# VGND -6.2e-19
C15808 _281_/Y _284_/A 0.019f
C15809 _343_/a_651_373# _229_/a_76_159# 1.34e-19
C15810 _344_/a_27_7# _164_/A 0.011f
C15811 _324_/a_27_7# _331_/CLK 6.01e-20
C15812 _271_/A _298_/C 0.0146f
C15813 _258_/S _309_/a_543_7# 2.7e-19
C15814 _328_/a_193_7# _220_/a_93_n19# 0.00158f
C15815 _328_/a_27_7# _220_/a_250_257# 6.8e-20
C15816 _329_/Q VGND 1.38f
C15817 _238_/B VPWR 0.871f
C15818 _208_/a_78_159# VPWR 0.00422f
C15819 _242_/A _331_/a_1283_n19# 1.58e-21
C15820 _326_/a_1108_7# _330_/Q 1.52e-20
C15821 _309_/a_27_7# _292_/A 5.13e-22
C15822 _255_/B clkbuf_0_clk/X 9.93e-21
C15823 _219_/a_250_257# _328_/Q 7.8e-21
C15824 _279_/Y _314_/D 0.038f
C15825 _342_/Q clk 0.757f
C15826 _313_/a_1283_n19# _336_/Q 1.14e-20
C15827 _313_/a_543_7# _225_/B 1.86e-20
C15828 _209_/X _191_/B 0.27f
C15829 _342_/D _308_/X 3.81e-19
C15830 _317_/a_651_373# _232_/A 8.99e-22
C15831 _327_/a_761_249# VGND -5.27e-19
C15832 _327_/a_1283_n19# VPWR 0.0169f
C15833 _203_/a_80_n19# _147_/Y 0.0131f
C15834 _273_/A trimb[3] 0.00719f
C15835 _342_/a_27_7# _342_/D 0.158f
C15836 _260_/A _193_/Y 9.04e-20
C15837 _346_/a_652_n19# _346_/D 0.013f
C15838 _273_/A _324_/a_27_7# 0.00326f
C15839 repeater43/X _315_/a_543_7# 0.0166f
C15840 _195_/a_27_257# _194_/X 0.0111f
C15841 _277_/Y _173_/a_489_373# 0.00297f
C15842 _326_/a_1283_n19# VPWR 0.0142f
C15843 _326_/a_761_249# VGND 0.00468f
C15844 _185_/A cal 0.0467f
C15845 _322_/a_1283_n19# _322_/Q 0.00965f
C15846 _307_/a_218_334# _341_/Q 1.04e-20
C15847 _234_/B _317_/a_543_7# 1.39e-21
C15848 _306_/S _344_/Q 8.72e-20
C15849 _169_/B _254_/A 1.41e-20
C15850 _324_/Q _296_/a_109_7# 0.00412f
C15851 _332_/a_805_7# VGND 1.88e-19
C15852 _332_/a_1462_7# VPWR 1.26e-19
C15853 _299_/X _346_/SET_B 0.0595f
C15854 _315_/D _347_/D 0.234f
C15855 _327_/a_543_7# repeater42/a_27_7# 7.41e-19
C15856 _328_/a_543_7# VPWR 0.0211f
C15857 _328_/a_193_7# VGND 0.0112f
C15858 _347_/a_1217_7# VGND 7.36e-20
C15859 _341_/Q _178_/a_109_257# 4.36e-19
C15860 _193_/Y _261_/A 9.92e-20
C15861 output10/a_27_7# _343_/CLK 0.0124f
C15862 _345_/a_193_7# _273_/A 3.42e-20
C15863 _191_/B _209_/a_109_257# 1.53e-19
C15864 _255_/B input1/X 0.00651f
C15865 _328_/a_1108_7# _297_/B 0.0122f
C15866 _321_/a_543_7# result[7] 2.6e-19
C15867 _314_/Q _347_/a_805_7# 4.25e-19
C15868 _248_/A _245_/a_113_257# 3.8e-19
C15869 _164_/Y _171_/a_292_257# 3.04e-21
C15870 _164_/A _171_/a_215_7# 4.79e-20
C15871 _258_/S _306_/a_535_334# 0.00106f
C15872 _257_/a_79_159# input1/X 1.14e-20
C15873 _257_/a_222_53# cal 6.01e-22
C15874 _298_/B _226_/a_297_7# 2.59e-20
C15875 _263_/B _311_/Q 0.00797f
C15876 _273_/A _266_/a_113_257# 1.9e-20
C15877 _259_/a_113_257# _311_/D 3.36e-20
C15878 _288_/A _344_/a_1602_7# 3.21e-20
C15879 _324_/a_761_249# _216_/a_27_7# 9.03e-19
C15880 _346_/a_1182_221# _160_/X 0.00169f
C15881 _346_/a_562_373# _299_/X 4.36e-19
C15882 _346_/a_381_7# _347_/Q 0.00197f
C15883 _343_/CLK _315_/a_1270_373# 5.21e-19
C15884 _258_/a_76_159# _196_/A 9.36e-21
C15885 _258_/a_505_n19# _286_/B 0.00817f
C15886 _334_/a_543_7# VPWR 0.0302f
C15887 _227_/A _343_/CLK 0.0132f
C15888 _334_/a_193_7# VGND -0.00466f
C15889 _225_/X _225_/B 0.00313f
C15890 _257_/a_222_53# _197_/a_27_7# 7e-20
C15891 _331_/CLK _245_/a_113_257# 0.0348f
C15892 _163_/a_292_257# _160_/X 0.00386f
C15893 _345_/Q _170_/a_489_373# 6.46e-20
C15894 _190_/a_27_7# VGND 0.0818f
C15895 _319_/Q _240_/B 0.151f
C15896 _342_/Q _150_/a_109_257# 0.00214f
C15897 _216_/a_27_7# _304_/X 1.83e-20
C15898 _342_/D _317_/D 1.15e-19
C15899 _216_/A _194_/X 2.28e-22
C15900 _323_/a_27_7# _298_/C 6.19e-20
C15901 _323_/a_761_249# _343_/Q 1.36e-20
C15902 _188_/S _286_/B 0.0102f
C15903 _294_/A _344_/Q 2.74e-20
C15904 clk _204_/Y 0.0993f
C15905 _192_/B _298_/A 3.09e-19
C15906 _331_/D _330_/a_651_373# 4.57e-20
C15907 _314_/a_1283_n19# _156_/a_39_257# 6.45e-19
C15908 _168_/a_109_257# _165_/X 0.00295f
C15909 _168_/a_397_257# _167_/X 0.00514f
C15910 _172_/A _304_/a_79_n19# 1.78e-20
C15911 _270_/a_121_257# _324_/Q 1.51e-20
C15912 _274_/a_39_257# VGND 0.0342f
C15913 _330_/a_193_7# _330_/a_651_373# -0.00701f
C15914 _275_/Y trim[3] 1.12e-19
C15915 ctln[3] _292_/A 3.65e-19
C15916 _341_/Q _144_/A 0.0272f
C15917 _329_/a_543_7# _281_/A 0.0395f
C15918 trim[4] _266_/a_113_257# 0.00294f
C15919 _164_/Y _161_/Y 1.09f
C15920 _329_/a_27_7# _281_/Y 0.0119f
C15921 _328_/a_639_7# _279_/A 0.00102f
C15922 _304_/S _224_/a_584_7# 3.63e-20
C15923 _294_/Y _267_/A 0.154f
C15924 _254_/A _170_/a_226_7# 7.23e-19
C15925 _342_/a_193_7# _177_/a_27_7# 3.28e-20
C15926 _255_/B _286_/Y 0.0958f
C15927 _236_/B _321_/Q 0.0163f
C15928 _330_/Q _316_/D 0.0995f
C15929 _248_/A VPWR 3.92f
C15930 _319_/a_27_7# _279_/A 2.62e-21
C15931 _295_/a_409_7# VGND -0.00119f
C15932 _346_/a_1032_373# VPWR 0.0088f
C15933 _346_/a_476_7# VGND 0.00961f
C15934 _149_/a_27_7# _315_/a_27_7# 2.75e-20
C15935 clkbuf_2_3_0_clk/A _215_/A 0.00807f
C15936 _271_/Y _208_/a_215_7# 2.37e-19
C15937 _160_/X _173_/a_226_257# 0.0011f
C15938 _337_/Q _310_/a_805_7# 1.78e-19
C15939 _167_/X _216_/A 7.14e-21
C15940 _335_/a_543_7# _204_/a_27_257# 6.78e-20
C15941 _335_/a_1108_7# _208_/a_78_159# 3.94e-19
C15942 _163_/a_78_159# VGND 0.00274f
C15943 _163_/a_493_257# VPWR -8.36e-20
C15944 _343_/a_193_7# _226_/a_382_257# 1.51e-20
C15945 _343_/a_27_7# _226_/a_297_7# 3.16e-21
C15946 _277_/Y clkbuf_2_3_0_clk/A 0.908f
C15947 _319_/Q _328_/Q 1.3f
C15948 _329_/a_193_7# _319_/Q 0.562f
C15949 _236_/a_109_257# VGND -0.00108f
C15950 _331_/CLK VPWR 6.98f
C15951 _318_/a_543_7# _248_/A 7.75e-20
C15952 _347_/Q _313_/a_193_7# 2.23e-21
C15953 _299_/X _313_/a_761_249# 2.31e-21
C15954 _346_/a_381_7# _297_/B 4.49e-19
C15955 _340_/CLK _311_/a_543_7# 1.77e-19
C15956 _337_/Q _265_/B 0.182f
C15957 _332_/Q VGND 0.375f
C15958 _190_/A VPWR 1.49f
C15959 _318_/Q _223_/a_93_n19# 8.33e-22
C15960 cal _335_/Q 0.00122f
C15961 _338_/Q _309_/Q 0.00112f
C15962 _329_/a_27_7# _329_/D 0.478f
C15963 result[0] result[1] 0.0416f
C15964 _263_/B _254_/B 4.63e-19
C15965 _236_/B _318_/a_193_7# 2.08e-19
C15966 _318_/a_543_7# _331_/CLK 3.78e-20
C15967 _273_/A VPWR 5.3f
C15968 _342_/a_1217_7# _342_/D 8.5e-19
C15969 _219_/a_93_n19# _319_/D 3.78e-20
C15970 _294_/A output33/a_27_7# 0.0253f
C15971 _277_/Y _172_/Y 1.36e-19
C15972 _340_/Q _193_/Y 1.22f
C15973 _196_/A _161_/Y 0.00244f
C15974 repeater43/a_27_7# _269_/Y 2.23e-19
C15975 clk _153_/a_487_257# 3.52e-19
C15976 cal _298_/a_109_7# 2.83e-19
C15977 output14/a_27_7# _322_/a_543_7# 2.3e-19
C15978 _215_/A _313_/a_1270_373# 3.5e-19
C15979 _299_/X _156_/a_39_257# 1.25e-19
C15980 _275_/A _279_/A 0.0151f
C15981 repeater43/X _324_/a_1283_n19# 0.0424f
C15982 _145_/A _341_/Q 0.473f
C15983 _242_/B _212_/X 1.31e-19
C15984 _345_/a_1182_221# _158_/Y 0.00433f
C15985 trim[0] _258_/S 3.46e-19
C15986 _305_/a_76_159# _305_/X 0.00308f
C15987 _218_/a_584_7# _346_/SET_B 6.4e-19
C15988 _222_/a_93_n19# VPWR 0.0105f
C15989 _332_/a_651_373# _153_/B 0.00209f
C15990 _324_/a_193_7# _212_/X 4.15e-19
C15991 _324_/a_27_7# _217_/X 1.22e-20
C15992 _343_/a_543_7# repeater43/X 0.00412f
C15993 _319_/Q _269_/A 0.0145f
C15994 _331_/Q _330_/a_1108_7# 5.37e-19
C15995 _328_/a_1462_7# VGND -8.76e-19
C15996 _173_/a_489_373# VGND -0.00129f
C15997 _173_/a_556_7# VPWR -1.5e-19
C15998 _341_/Q _146_/a_112_13# 7.47e-21
C15999 _221_/a_256_7# _327_/D 4.89e-19
C16000 _284_/A _297_/Y 0.00538f
C16001 _283_/A _207_/a_27_7# 1.06e-22
C16002 _271_/A _334_/a_1270_373# 4.61e-19
C16003 _319_/a_543_7# VGND 0.0427f
C16004 _319_/a_1108_7# VPWR 0.0215f
C16005 _346_/SET_B _311_/a_1283_n19# 4.89e-19
C16006 _338_/Q _311_/a_193_7# 1.49e-20
C16007 _344_/a_27_7# _292_/A 0.00116f
C16008 _337_/a_543_7# VPWR 0.0035f
C16009 _337_/a_193_7# VGND 0.0305f
C16010 _231_/a_79_n19# _162_/X 0.00545f
C16011 trim[4] VPWR 0.17f
C16012 _304_/X _327_/Q 0.147f
C16013 _299_/X _147_/A 0.0138f
C16014 _342_/a_27_7# _341_/a_193_7# 1.2e-22
C16015 _342_/a_193_7# _341_/a_27_7# 7.41e-20
C16016 _216_/a_27_7# VGND 0.0596f
C16017 _343_/Q _154_/a_27_7# 3.59e-21
C16018 _258_/S _311_/Q 0.329f
C16019 _297_/B _313_/a_193_7# 9.97e-21
C16020 _215_/A _192_/B 7.68e-20
C16021 _344_/a_27_7# _160_/A 2.33e-22
C16022 _313_/Q _286_/B 0.164f
C16023 _325_/Q _286_/Y 1.56e-21
C16024 _334_/a_1462_7# VGND -9.48e-19
C16025 clk _225_/B 1.28e-19
C16026 _189_/a_27_7# ctln[6] 1.29e-20
C16027 _167_/a_109_7# _166_/Y 0.00187f
C16028 _341_/a_1108_7# _188_/S 9.63e-19
C16029 _297_/A _147_/Y 7.04e-21
C16030 _320_/Q _320_/a_448_7# 9.75e-20
C16031 _329_/Q _320_/a_1108_7# 4.44e-20
C16032 _339_/Q _265_/B 5.43e-21
C16033 _315_/D _156_/a_121_257# 1.04e-19
C16034 _187_/a_27_7# _304_/S 0.00117f
C16035 _345_/a_1602_7# _345_/D 5.75e-20
C16036 _345_/a_381_7# _345_/Q 1.44e-19
C16037 _307_/a_505_n19# VPWR 0.0704f
C16038 _281_/Y _342_/Q 3.38e-20
C16039 _324_/Q _243_/a_113_257# 1.12e-19
C16040 _304_/S _315_/D 0.0102f
C16041 _275_/Y _338_/D 7.04e-21
C16042 _294_/A _306_/S 0.495f
C16043 _145_/a_113_7# VPWR -3.62e-20
C16044 _325_/a_1270_373# _326_/Q 9.84e-20
C16045 _309_/a_27_7# trim[4] 1.96e-19
C16046 cal _199_/a_93_n19# 0.00221f
C16047 _323_/D _176_/a_27_7# 0.00558f
C16048 _164_/A _147_/Y 1.65e-19
C16049 _146_/C _298_/A 0.00616f
C16050 output12/a_27_7# rstn 1.22e-21
C16051 _178_/a_27_7# VPWR 0.089f
C16052 _336_/Q _202_/a_93_n19# 2.26e-20
C16053 _260_/B _172_/A 0.0141f
C16054 _329_/a_1217_7# _281_/Y 2.55e-19
C16055 _157_/A _298_/A 2.12e-19
C16056 clkbuf_2_1_0_clk/A _337_/Q 0.0246f
C16057 _340_/a_1108_7# _198_/a_250_257# 6.51e-20
C16058 _307_/X _315_/D 1.8e-20
C16059 _226_/a_382_257# VGND -6.04e-19
C16060 _272_/a_39_257# _327_/Q 1.03e-20
C16061 clk en 0.0697f
C16062 _292_/A _171_/a_215_7# 0.00516f
C16063 cal _336_/Q 0.109f
C16064 _325_/a_27_7# _324_/a_761_249# 8.8e-19
C16065 _346_/a_1224_7# VGND 8.27e-20
C16066 _337_/Q _310_/Q 0.722f
C16067 _165_/a_78_159# _161_/Y 0.0407f
C16068 _169_/Y _301_/X 3.78e-19
C16069 rstn _207_/a_109_7# 5.27e-19
C16070 _335_/a_1108_7# _190_/A 2.18e-19
C16071 clkbuf_0_clk/X _314_/a_193_7# 0.0186f
C16072 _309_/a_1270_373# _346_/SET_B -2.06e-19
C16073 _335_/a_1270_373# _207_/X 2.86e-20
C16074 _197_/a_27_7# _336_/Q 0.0621f
C16075 _267_/a_109_257# VPWR -2.18e-19
C16076 _160_/A _171_/a_215_7# 0.00197f
C16077 _343_/a_1108_7# _150_/C 2.02e-20
C16078 _343_/a_1283_n19# _226_/X 4.18e-19
C16079 _194_/A _254_/B 0.0407f
C16080 _339_/a_193_7# VGND -0.00466f
C16081 _339_/a_543_7# VPWR 0.0104f
C16082 result[4] _234_/B 2.96e-20
C16083 _341_/a_193_7# _317_/D 0.0138f
C16084 _341_/a_543_7# _244_/B 3.94e-20
C16085 _308_/a_505_n19# _206_/A 6.71e-20
C16086 _327_/a_543_7# _232_/X 0.00784f
C16087 _282_/a_39_257# VGND 0.0474f
C16088 _275_/Y _273_/Y 6.2e-21
C16089 _325_/a_27_7# _304_/X 0.225f
C16090 input4/X _271_/A 2.12e-19
C16091 _343_/a_27_7# _149_/a_27_7# 4.33e-21
C16092 _283_/A _306_/S 0.00713f
C16093 _326_/a_543_7# _232_/X 0.00379f
C16094 _321_/D _318_/a_805_7# 2.96e-19
C16095 _254_/A _279_/A 1.02e-19
C16096 input4/X _335_/a_27_7# 7.37e-19
C16097 _258_/S _254_/B 8.96e-19
C16098 _321_/Q _331_/a_193_7# 2.66e-20
C16099 _330_/Q _331_/a_27_7# 0.0406f
C16100 trim[2] _297_/Y 2.3e-19
C16101 _290_/A clkc 0.00291f
C16102 clkbuf_2_3_0_clk/A VGND 0.916f
C16103 _329_/Q ctlp[5] 0.0474f
C16104 _341_/a_543_7# _323_/D 4.33e-20
C16105 _255_/B _296_/a_295_257# 0.00583f
C16106 _312_/a_193_7# _312_/Q 0.0147f
C16107 _312_/a_1108_7# _312_/D 1.91e-21
C16108 _328_/a_761_249# _232_/X 5.02e-19
C16109 _200_/a_93_n19# _197_/X 0.0423f
C16110 _320_/a_27_7# _346_/SET_B 0.101f
C16111 _271_/Y _206_/A 0.00871f
C16112 _271_/A _207_/C 0.112f
C16113 _340_/a_543_7# _254_/B 1.03e-20
C16114 _327_/Q VGND 1.56f
C16115 _217_/X VPWR 3.16f
C16116 _223_/a_93_n19# _223_/a_346_7# -5.12e-20
C16117 _324_/a_1462_7# _212_/X 2.7e-20
C16118 _335_/a_27_7# _207_/C 1.57e-20
C16119 _335_/a_761_249# _206_/A 3.36e-20
C16120 repeater43/X _318_/a_651_373# 0.00247f
C16121 _309_/D _309_/Q 1.3e-20
C16122 _316_/a_761_249# _317_/D 0.00394f
C16123 _172_/Y VGND 0.0703f
C16124 clkbuf_2_1_0_clk/A _339_/Q 0.0157f
C16125 _288_/A _162_/X 0.0083f
C16126 _154_/a_27_7# _204_/a_27_7# 5.6e-21
C16127 _306_/S _248_/B 6.44e-20
C16128 _318_/a_1283_n19# _212_/X 1.76e-20
C16129 _318_/a_1108_7# _327_/Q 1.03e-19
C16130 _288_/A _287_/a_39_257# 0.00296f
C16131 _271_/Y _334_/D 3.67e-19
C16132 _326_/Q _286_/Y 0.0829f
C16133 _313_/a_805_7# VPWR 1.05e-19
C16134 _313_/a_1270_373# VGND 4.01e-19
C16135 _289_/a_39_257# _312_/Q 0.00116f
C16136 _281_/Y _336_/a_27_7# 1.21e-21
C16137 output7/a_27_7# _271_/Y 0.0164f
C16138 _337_/a_1462_7# VGND -8.98e-19
C16139 _330_/Q _217_/a_27_7# 0.00179f
C16140 _328_/a_193_7# ctlp[5] 6.7e-20
C16141 _324_/Q _341_/Q 0.0943f
C16142 _335_/a_761_249# _334_/D 9.68e-19
C16143 _335_/a_543_7# _343_/CLK 0.00148f
C16144 _275_/Y _343_/CLK 2.24e-19
C16145 repeater42/a_27_7# _212_/X 0.0674f
C16146 _286_/B _333_/a_1283_n19# 1.03e-19
C16147 _250_/a_292_257# _225_/B 4.06e-20
C16148 ctln[1] VGND 0.151f
C16149 _254_/Y _306_/S 0.00573f
C16150 _315_/a_1283_n19# _286_/Y 1.21e-19
C16151 _342_/D _196_/A 1.66e-20
C16152 _318_/Q _216_/X 0.00469f
C16153 _296_/Y VPWR 0.223f
C16154 _157_/A _215_/A 0.00723f
C16155 ctln[2] VGND 0.0737f
C16156 _320_/Q _331_/D 2.15e-20
C16157 _272_/a_39_257# _317_/a_1108_7# 2.63e-20
C16158 _165_/X _301_/a_149_7# 3.26e-20
C16159 _167_/X _301_/a_240_7# 0.00192f
C16160 _274_/a_121_257# _232_/X 2.15e-19
C16161 _315_/Q _244_/B 0.0114f
C16162 _188_/a_76_159# _186_/a_297_7# 5.6e-21
C16163 rstn _193_/Y 0.0697f
C16164 _320_/Q _330_/a_193_7# 0.545f
C16165 _172_/A _295_/a_512_7# 4.17e-19
C16166 _283_/Y _332_/D 3.27e-20
C16167 _342_/a_1283_n19# _229_/a_226_7# 0.00389f
C16168 _327_/a_193_7# _331_/D 7.24e-20
C16169 _342_/Q _185_/A 3.63e-20
C16170 _344_/a_27_7# _273_/A 3.39e-22
C16171 _271_/A _150_/C 0.016f
C16172 _192_/B VGND 2.51f
C16173 _146_/a_29_271# VPWR 0.0572f
C16174 input4/X _323_/a_27_7# 2.43e-19
C16175 _162_/X _299_/a_493_257# 2.76e-20
C16176 _314_/a_193_7# _297_/a_27_257# 1.02e-19
C16177 _319_/Q _321_/a_1270_373# 4.59e-20
C16178 _346_/SET_B _171_/a_78_159# 9.26e-19
C16179 _336_/Q _284_/A 0.266f
C16180 _340_/a_805_7# _197_/X 5.24e-19
C16181 clk _315_/D 1.24e-20
C16182 clkbuf_0_clk/a_110_7# VPWR 0.2f
C16183 _302_/a_227_7# _300_/Y 0.00108f
C16184 _333_/a_27_7# _298_/C 4.16e-21
C16185 _325_/a_761_249# VPWR 0.0063f
C16186 _325_/a_27_7# VGND -0.0677f
C16187 _305_/a_535_334# _340_/CLK 3.23e-19
C16188 _211_/a_27_257# _190_/A 4.73e-21
C16189 _271_/A _317_/a_193_7# 4.3e-19
C16190 _323_/a_27_7# _207_/C 9.18e-21
C16191 _323_/a_761_249# _206_/A 8.15e-21
C16192 _255_/B _255_/X 0.00226f
C16193 _319_/Q clkbuf_2_3_0_clk/a_75_172# 2.04e-20
C16194 _335_/D _333_/Q 5.39e-19
C16195 _257_/a_79_159# _255_/X 8.99e-21
C16196 _248_/B _327_/D 7.08e-21
C16197 _339_/a_1462_7# VGND -8.76e-19
C16198 _333_/a_761_249# _332_/a_1283_n19# 4.37e-22
C16199 _333_/a_1108_7# _332_/a_193_7# 5.13e-19
C16200 _333_/a_193_7# _332_/a_1108_7# 7.59e-19
C16201 _333_/a_1283_n19# _332_/a_761_249# 2.05e-20
C16202 clkbuf_0_clk/X _324_/D 4.09e-19
C16203 _313_/D _340_/CLK 0.0539f
C16204 output20/a_27_7# clkbuf_0_clk/X 0.0541f
C16205 _325_/a_1217_7# _304_/X 9.18e-19
C16206 _294_/A _254_/Y 0.0859f
C16207 _317_/a_1108_7# VGND 0.0132f
C16208 _317_/a_651_373# VPWR 0.00155f
C16209 _281_/Y _225_/B 0.0143f
C16210 _212_/a_27_7# _316_/D 0.00823f
C16211 _215_/A _260_/A 0.0127f
C16212 _323_/a_543_7# _343_/CLK 0.0217f
C16213 _182_/a_215_7# _182_/X 0.00213f
C16214 repeater42/a_27_7# _325_/a_193_7# 1.59e-20
C16215 trimb[2] VGND 0.198f
C16216 _297_/A _347_/a_193_7# 0.0307f
C16217 _341_/Q _228_/A 0.00749f
C16218 _330_/Q _331_/a_1217_7# 1.93e-19
C16219 _172_/A _173_/a_226_257# 4.91e-19
C16220 _258_/a_76_159# _313_/a_193_7# 2e-20
C16221 _258_/a_505_n19# _313_/a_27_7# 4.78e-20
C16222 _277_/Y _260_/A 0.0204f
C16223 clkbuf_0_clk/X _278_/a_150_257# 1.47e-21
C16224 output24/a_27_7# result[2] 0.00541f
C16225 _292_/A _147_/Y 3.76e-21
C16226 _317_/Q _230_/a_27_7# 9.27e-21
C16227 _337_/Q _311_/a_27_7# 0.00298f
C16228 _169_/Y _166_/Y 2.16e-20
C16229 _292_/A _312_/a_1108_7# 0.00418f
C16230 _325_/Q _269_/A 1.8e-20
C16231 _314_/a_761_249# _284_/A 2.56e-21
C16232 _197_/X _340_/CLK 0.0292f
C16233 _312_/a_1462_7# _312_/Q 5.4e-19
C16234 _308_/S _307_/a_439_7# 3.65e-19
C16235 _160_/A _147_/Y 7.7e-21
C16236 _331_/a_1270_373# VGND 3.79e-19
C16237 _320_/a_1217_7# _346_/SET_B 1.14e-19
C16238 _331_/a_805_7# VPWR 2.56e-19
C16239 _301_/X _315_/D 3.12e-21
C16240 _310_/a_27_7# clkc 7.41e-22
C16241 _294_/Y _310_/a_1108_7# 1.52e-20
C16242 _302_/a_227_7# VGND 0.0459f
C16243 _283_/A _248_/B 0.00879f
C16244 _223_/a_250_257# _325_/D 6.81e-20
C16245 _276_/a_68_257# _297_/B 2.03e-21
C16246 _344_/a_562_373# _346_/SET_B 4.13e-19
C16247 _162_/A output40/a_27_7# 0.0146f
C16248 _337_/a_543_7# _198_/a_93_n19# 1.85e-20
C16249 _343_/a_1108_7# cal 0.00508f
C16250 _343_/a_1283_n19# input1/X 0.0042f
C16251 clkbuf_0_clk/X _279_/A 0.011f
C16252 _277_/Y _261_/A 1.36e-19
C16253 _317_/Q _232_/A 0.632f
C16254 _336_/a_1283_n19# _193_/Y 3.7e-21
C16255 _172_/A _307_/a_76_159# 0.00924f
C16256 _255_/a_30_13# _209_/a_109_257# 3.77e-21
C16257 _274_/a_39_257# _318_/Q 0.00463f
C16258 _157_/A _300_/Y 0.662f
C16259 _254_/B _201_/a_27_7# 1.08e-19
C16260 clkbuf_0_clk/X _218_/a_250_257# 1.32e-19
C16261 _322_/a_543_7# _321_/D 1.69e-19
C16262 _325_/a_1108_7# _246_/B 1.27e-19
C16263 _341_/Q _216_/A 5.41e-20
C16264 _308_/S _225_/X 2.67e-20
C16265 _310_/a_193_7# _310_/a_761_249# -0.0105f
C16266 _310_/a_27_7# _310_/a_543_7# -0.00469f
C16267 _307_/X _308_/S 0.00189f
C16268 _323_/a_761_249# _149_/A 1.13e-19
C16269 _283_/Y clkbuf_2_2_0_clk/a_75_172# 3.95e-19
C16270 _301_/a_51_257# _301_/a_240_7# -6e-19
C16271 _283_/Y input4/X 0.383f
C16272 _162_/X _298_/C 3.09e-20
C16273 _186_/a_297_7# _147_/A 0.0047f
C16274 _186_/a_79_n19# _150_/C 9.87e-21
C16275 _324_/a_1108_7# _286_/Y 0.0107f
C16276 _340_/CLK _312_/a_193_7# 0.00969f
C16277 _188_/S _178_/a_109_257# 5.04e-20
C16278 repeater43/X _322_/a_27_7# -1.89e-19
C16279 _342_/a_1270_373# _248_/A 9.62e-20
C16280 _309_/a_1283_n19# _337_/Q 2.98e-19
C16281 _251_/a_79_n19# _215_/A 0.0026f
C16282 _339_/Q _311_/a_27_7# 0.0176f
C16283 _326_/Q _328_/Q 0.00299f
C16284 clkbuf_2_0_0_clk/a_75_172# _193_/Y 1.35e-19
C16285 ctln[6] _154_/A 3.2e-19
C16286 _154_/a_27_7# _206_/A 0.0115f
C16287 _146_/C VGND 0.872f
C16288 _186_/a_297_7# _149_/A 4.57e-21
C16289 _273_/A _227_/a_113_7# 6.23e-20
C16290 _260_/B _297_/A 1.18e-20
C16291 _219_/a_93_n19# _297_/B 0.0469f
C16292 _346_/SET_B _172_/B 0.553f
C16293 ctln[7] _206_/A 9.7e-20
C16294 clk _335_/a_193_7# 8.07e-21
C16295 _283_/Y _207_/C 1.69e-19
C16296 _337_/a_27_7# _254_/B 3.49e-21
C16297 _306_/X _190_/A 2.11e-20
C16298 _257_/a_79_159# _336_/a_193_7# 2.53e-20
C16299 repeater43/X _214_/a_109_7# 8.94e-22
C16300 _324_/D _286_/Y 0.00809f
C16301 _320_/a_543_7# _217_/X 1.03e-21
C16302 _294_/A _336_/a_1108_7# 7.8e-20
C16303 _179_/a_27_7# _206_/A 8.2e-21
C16304 _157_/A VGND 1.35f
C16305 _293_/a_121_257# _254_/A 5.59e-19
C16306 _304_/a_79_n19# _325_/D 2.84e-20
C16307 output21/a_27_7# _320_/Q 1.53e-19
C16308 _214_/a_27_257# _327_/Q 0.0422f
C16309 _300_/Y _260_/A 6.44e-20
C16310 _325_/a_1217_7# VGND -3.66e-19
C16311 _339_/a_543_7# _198_/a_93_n19# 7.73e-22
C16312 ctln[7] _334_/D 5.23e-20
C16313 _321_/a_27_7# _321_/a_761_249# -0.0166f
C16314 input1/X _311_/a_193_7# 2.97e-21
C16315 _271_/A _317_/a_1462_7# 3.73e-19
C16316 _196_/A _194_/A 0.00515f
C16317 _181_/X _305_/X 4.63e-22
C16318 _320_/D _319_/a_1283_n19# 7.86e-19
C16319 _298_/B _306_/S 1.18e-21
C16320 _347_/Q _344_/D 0.00131f
C16321 _160_/X _344_/Q 1.46e-21
C16322 _342_/a_193_7# repeater43/X 0.00402f
C16323 _165_/a_215_7# _162_/X 3.3e-21
C16324 _306_/S _194_/a_27_7# 4.98e-21
C16325 _259_/a_199_7# _258_/S 1.85e-19
C16326 _188_/S _144_/A 9.48e-19
C16327 _346_/SET_B _312_/a_761_249# 0.0036f
C16328 _258_/S _196_/A 0.0311f
C16329 _271_/A cal 0.0533f
C16330 _326_/a_1283_n19# _223_/a_250_257# 6.05e-21
C16331 _326_/a_1108_7# _223_/a_93_n19# 1.26e-20
C16332 _202_/a_584_7# VGND -7.74e-19
C16333 _279_/A _286_/Y 0.0764f
C16334 _304_/X _221_/a_250_257# 0.00152f
C16335 _346_/Q _347_/Q 4.51e-20
C16336 _297_/A _347_/a_1462_7# 3.42e-19
C16337 _332_/a_27_7# _332_/a_193_7# -0.0297f
C16338 clkbuf_2_1_0_clk/A clkbuf_1_0_0_clk/a_75_172# 0.00207f
C16339 _273_/A _248_/a_109_257# 0.00362f
C16340 trimb[0] comp 0.0055f
C16341 _215_/A _340_/Q 1.3e-20
C16342 _219_/a_584_7# _279_/A 0.00103f
C16343 _313_/Q _313_/a_27_7# 0.00107f
C16344 _273_/A output16/a_27_7# 0.0366f
C16345 _319_/Q _299_/X 8.44e-20
C16346 _347_/a_193_7# _347_/a_761_249# -0.00517f
C16347 _347_/a_27_7# _347_/a_543_7# -0.00482f
C16348 _341_/a_651_373# _177_/a_27_7# 0.00111f
C16349 _341_/a_543_7# _177_/A 1.53e-19
C16350 _277_/Y _340_/Q -1.05e-36
C16351 _232_/X _212_/X 0.113f
C16352 _167_/X _300_/a_383_7# 1.17e-19
C16353 _168_/a_109_7# _160_/X 2.8e-20
C16354 _335_/Q _204_/Y 0.247f
C16355 _340_/a_543_7# _196_/A 0.0067f
C16356 _330_/Q _281_/A 0.014f
C16357 _210_/a_307_257# _209_/X 1.27e-21
C16358 _216_/X _286_/B 8.24e-20
C16359 _269_/A _315_/a_1283_n19# 0.00655f
C16360 _323_/a_1270_373# _323_/Q 3.69e-19
C16361 _149_/A _154_/a_27_7# 1.14e-19
C16362 _260_/A VGND 0.541f
C16363 _197_/X _337_/a_651_373# 3.67e-19
C16364 _275_/Y _174_/a_109_257# 0.0086f
C16365 _342_/a_448_7# _343_/CLK 2.28e-19
C16366 _190_/A _147_/Y 0.00209f
C16367 _281_/Y _315_/D 0.00755f
C16368 _283_/Y _339_/a_1270_373# 8.07e-21
C16369 output12/a_27_7# VPWR 0.104f
C16370 _342_/Q _336_/Q 7.62e-20
C16371 _165_/X _215_/A 3.15e-20
C16372 _323_/a_193_7# clk 0.00154f
C16373 _281_/Y _324_/a_651_373# 4.47e-19
C16374 _273_/A _147_/Y 1.87e-21
C16375 _294_/A _284_/a_39_257# 0.00391f
C16376 _257_/a_222_53# _225_/B 0.00197f
C16377 _169_/Y _297_/Y 0.00531f
C16378 _342_/D _341_/D 5.92e-20
C16379 _277_/Y _165_/X 1.11f
C16380 _273_/A _312_/a_1108_7# 2.69e-21
C16381 _325_/a_27_7# _214_/a_27_257# 7.38e-22
C16382 _308_/S clk 1.61e-19
C16383 _326_/a_27_7# _181_/X 0.00376f
C16384 _294_/A _194_/a_27_7# 9.76e-21
C16385 _185_/A en 8.7e-19
C16386 _256_/a_209_257# _260_/B 1.89e-20
C16387 _297_/B _344_/D 0.00185f
C16388 _232_/A _315_/a_193_7# 1.02e-19
C16389 _248_/B _315_/a_27_7# 4.61e-19
C16390 _232_/A _298_/A 1.35e-22
C16391 _145_/A _188_/S 0.315f
C16392 _261_/A VGND 0.0313f
C16393 _239_/a_113_257# VGND -0.00101f
C16394 _314_/D _228_/A 0.0123f
C16395 result[1] _324_/Q 1.3e-19
C16396 _331_/CLK _330_/a_639_7# 9.32e-19
C16397 _346_/Q _297_/B 0.0789f
C16398 _168_/a_109_257# VPWR 6.37e-19
C16399 _314_/Q _267_/A 1.3e-20
C16400 _265_/a_109_257# VGND -9.42e-19
C16401 _207_/a_109_7# VPWR -2.51e-19
C16402 _217_/a_27_7# _212_/a_27_7# 7.59e-20
C16403 _173_/a_556_7# _147_/Y 3.04e-19
C16404 _309_/a_193_7# _344_/Q 3.43e-20
C16405 _342_/a_1108_7# _147_/A 2.38e-21
C16406 _319_/Q _318_/a_27_7# 3.34e-19
C16407 _293_/a_39_257# _337_/Q 1.62e-19
C16408 _346_/a_193_7# _299_/a_78_159# 1.88e-19
C16409 _342_/Q _315_/a_1108_7# 1.86e-21
C16410 _251_/X _215_/A 0.0177f
C16411 _330_/Q _216_/A 3.22e-21
C16412 _197_/X _225_/X 1.57e-19
C16413 _333_/a_651_373# _332_/Q 1.15e-19
C16414 _333_/a_1108_7# _190_/A 0.0107f
C16415 _323_/a_27_7# cal 0.0138f
C16416 _248_/A _223_/a_250_257# 2.26e-19
C16417 _342_/a_1108_7# _149_/A 0.00199f
C16418 _254_/Y _336_/a_1108_7# 0.0546f
C16419 _325_/a_193_7# _232_/X 1.87e-19
C16420 _341_/a_193_7# _341_/a_448_7# -0.00297f
C16421 repeater43/X _330_/a_761_249# 0.00351f
C16422 _279_/Y _347_/a_27_7# 0.00227f
C16423 _167_/X _346_/D 3.71e-20
C16424 _288_/A output35/a_27_7# 7.49e-20
C16425 _294_/A _262_/a_113_257# 2.16e-20
C16426 repeater43/X result[3] 3.13e-19
C16427 _298_/B _283_/A 0.00247f
C16428 _332_/a_27_7# _208_/a_78_159# 3.13e-22
C16429 _316_/D _223_/a_93_n19# 0.00382f
C16430 _345_/a_476_7# _165_/X 0.00153f
C16431 _251_/a_79_n19# VGND 0.0288f
C16432 _251_/a_215_7# VPWR -0.00126f
C16433 _338_/a_193_7# _338_/a_448_7# -0.00779f
C16434 _275_/A ctlp[4] 2.69e-20
C16435 _221_/a_346_7# VPWR -8.08e-19
C16436 _221_/a_250_257# VGND -0.00147f
C16437 result[4] _318_/a_651_373# 3.52e-19
C16438 _160_/X _306_/S 0.613f
C16439 _318_/Q _327_/Q 1.75f
C16440 _216_/A _314_/D 6.01e-20
C16441 _281_/Y _218_/a_346_7# 0.00147f
C16442 _298_/B _205_/a_382_257# 7.88e-20
C16443 _186_/a_79_n19# cal 4.95e-19
C16444 _342_/a_1462_7# repeater43/X -6.42e-19
C16445 _240_/B _279_/A 1.81e-19
C16446 _191_/B _203_/a_303_7# 9.72e-21
C16447 _192_/B _203_/a_209_257# 0.00274f
C16448 _323_/Q _254_/B 2.38e-20
C16449 _294_/Y _345_/a_27_7# 1.08e-20
C16450 _251_/X _304_/X 0.00132f
C16451 _322_/a_27_7# result[6] 0.0251f
C16452 _333_/a_761_249# _206_/A 0.0523f
C16453 _333_/a_27_7# _207_/C 0.0108f
C16454 trim[1] _346_/SET_B 7.38e-20
C16455 _319_/Q _246_/B 0.00764f
C16456 _167_/a_27_257# _299_/X 0.0011f
C16457 _232_/X _331_/a_639_7# 9.29e-19
C16458 _345_/a_956_373# _290_/A 3.3e-19
C16459 _286_/B _295_/a_409_7# 8.4e-21
C16460 _306_/a_535_334# _267_/A 1.94e-19
C16461 _210_/a_27_7# _153_/A 0.0116f
C16462 _336_/a_27_7# _336_/Q 3.02e-20
C16463 _200_/a_93_n19# _200_/a_256_7# -6.6e-20
C16464 _267_/A _311_/a_805_7# 5.78e-19
C16465 _343_/CLK _333_/a_543_7# 4.44e-20
C16466 _149_/a_27_7# _244_/B 0.0259f
C16467 _241_/a_199_7# _327_/Q 0.00132f
C16468 _304_/a_79_n19# _248_/A 1.16e-20
C16469 _231_/a_79_n19# _150_/C 0.00943f
C16470 _286_/B _332_/Q 0.00119f
C16471 _337_/Q _198_/a_584_7# 0.00188f
C16472 _193_/Y VPWR 0.548f
C16473 _275_/Y _344_/D 0.163f
C16474 _340_/Q VGND 1.54f
C16475 _309_/a_448_7# _284_/A 0.0139f
C16476 _342_/D _343_/CLK 0.00305f
C16477 clkbuf_2_1_0_clk/A _319_/D 1.34e-20
C16478 _294_/A _160_/X 0.00174f
C16479 _328_/Q _279_/A 0.0392f
C16480 _317_/a_1283_n19# _317_/D 4.6e-19
C16481 repeater43/X _322_/Q 0.242f
C16482 _252_/a_109_257# _304_/S 7.61e-21
C16483 _275_/Y _346_/Q 5.18e-20
C16484 _279_/Y _216_/X 2.37e-21
C16485 _254_/Y _194_/a_27_7# 1.6e-20
C16486 _315_/Q _341_/a_1283_n19# 1.55e-22
C16487 result[0] _341_/a_761_249# 2.66e-19
C16488 _308_/S _250_/a_292_257# 1.56e-21
C16489 _316_/a_27_7# _316_/a_639_7# -0.0015f
C16490 _310_/a_1270_373# _310_/D 3.05e-19
C16491 _310_/a_1283_n19# _310_/Q 0.0178f
C16492 _329_/a_761_249# _218_/a_93_n19# 1.26e-19
C16493 _329_/a_193_7# _218_/a_250_257# 0.00139f
C16494 _199_/a_93_n19# _199_/a_250_257# -6.97e-22
C16495 _218_/a_250_257# _328_/Q 3.24e-21
C16496 _248_/A _176_/a_27_7# 1.35e-20
C16497 _289_/a_39_257# _267_/B 0.00168f
C16498 _256_/a_80_n19# _190_/A 0.0921f
C16499 _325_/a_27_7# _318_/Q 3.46e-21
C16500 _327_/a_1108_7# _216_/X 1.21e-19
C16501 _273_/A _286_/a_113_7# 2.73e-19
C16502 _324_/a_193_7# _248_/B 2.17e-19
C16503 _273_/A _304_/a_79_n19# 1.04e-20
C16504 _333_/a_193_7# _225_/X 2.58e-21
C16505 _290_/A _311_/a_1283_n19# 0.0158f
C16506 _283_/Y cal 0.053f
C16507 _309_/a_193_7# _306_/S 5.64e-19
C16508 _343_/a_448_7# _185_/A 0.00225f
C16509 _165_/X VGND 1.02f
C16510 _231_/a_512_7# _144_/A 0.0015f
C16511 _286_/B _173_/a_489_373# 1.25e-19
C16512 _327_/a_1108_7# _329_/Q 5.32e-20
C16513 _277_/Y rstn 0.00156f
C16514 _327_/a_193_7# _327_/a_448_7# -0.00482f
C16515 _232_/A _304_/X 6.84e-20
C16516 _248_/A _347_/a_193_7# 3.56e-19
C16517 _255_/a_184_257# VGND -3.87e-19
C16518 result[3] _317_/a_543_7# 6.24e-20
C16519 _340_/a_193_7# _340_/CLK 0.0267f
C16520 output15/a_27_7# _236_/B 7.16e-21
C16521 _288_/A _345_/Q 0.00962f
C16522 _188_/S _324_/Q 0.105f
C16523 clk _197_/X 1.04e-20
C16524 _323_/a_1217_7# cal 1.75e-19
C16525 _333_/D _333_/Q 3.33e-19
C16526 output5/a_27_7# VPWR 0.0794f
C16527 _341_/a_193_7# _341_/D 0.00908f
C16528 _329_/a_651_373# _330_/Q 0.00147f
C16529 _305_/a_505_n19# input1/X 8.21e-20
C16530 _162_/X _345_/Q 0.0305f
C16531 _161_/Y _174_/a_109_257# 5.14e-19
C16532 _332_/a_761_249# _332_/Q 2.57e-19
C16533 _332_/a_27_7# _190_/A 6.1e-21
C16534 _332_/a_193_7# _333_/Q 0.0263f
C16535 _338_/D _194_/A 8.74e-21
C16536 _336_/Q _225_/B 0.793f
C16537 _164_/Y _158_/Y 0.581f
C16538 _227_/A _209_/X 2.47e-19
C16539 _326_/a_193_7# _326_/a_448_7# -0.00779f
C16540 _328_/a_1108_7# _320_/Q 0.00542f
C16541 _285_/A _344_/Q 3.38e-19
C16542 _339_/Q _198_/a_584_7# 0.00311f
C16543 _317_/Q _245_/a_113_257# 0.00107f
C16544 _251_/X VGND 0.122f
C16545 repeater43/X _333_/a_639_7# -7.75e-19
C16546 _338_/a_27_7# _346_/SET_B 0.111f
C16547 _338_/a_193_7# _338_/D 0.513f
C16548 _329_/a_1283_n19# VGND 0.025f
C16549 _329_/a_448_7# VPWR -0.0026f
C16550 _308_/a_439_7# _306_/S 4.26e-19
C16551 _296_/a_213_83# VGND 0.0283f
C16552 _281_/Y _308_/S 1.8e-21
C16553 _306_/a_76_159# _193_/Y 3.39e-21
C16554 comp VPWR 0.647f
C16555 _344_/a_193_7# _344_/Q 5.22e-20
C16556 _341_/a_543_7# _248_/A 0.0126f
C16557 _306_/a_505_n19# _306_/S 0.0696f
C16558 _342_/a_543_7# cal 5.36e-19
C16559 _319_/Q result[5] 3.52e-19
C16560 _297_/A _212_/X 1.14e-19
C16561 _294_/A _309_/a_193_7# 0.0222f
C16562 _279_/Y _190_/a_27_7# 5.96e-19
C16563 _338_/Q _312_/Q 0.524f
C16564 _319_/Q _320_/a_27_7# 2.23e-19
C16565 _181_/a_27_7# _286_/Y 3.06e-19
C16566 _322_/a_1217_7# result[6] 3.42e-19
C16567 _332_/a_448_7# _332_/D 0.00345f
C16568 _301_/a_512_257# _160_/X 6.75e-19
C16569 _290_/A _309_/a_1270_373# 1.55e-19
C16570 _309_/Q clkc 1.06e-19
C16571 repeater42/a_27_7# _327_/D 0.0172f
C16572 _182_/a_297_257# _150_/C 2.58e-20
C16573 _182_/a_215_7# _225_/X 2.49e-19
C16574 _340_/a_761_249# _346_/SET_B 0.00704f
C16575 _196_/A _226_/a_79_n19# 1.32e-19
C16576 _172_/A _344_/Q 0.123f
C16577 _267_/A _311_/Q 0.00183f
C16578 output12/a_27_7# _211_/a_27_257# 0.0127f
C16579 _196_/A _339_/a_27_7# 1.54e-19
C16580 _314_/a_761_249# _225_/B 3.67e-19
C16581 result[4] _322_/a_27_7# 9.94e-21
C16582 _292_/A _163_/a_292_257# 0.00209f
C16583 _255_/B _246_/B 1.18e-20
C16584 _242_/A _315_/D 6.44e-20
C16585 _215_/A _336_/a_1283_n19# 8.48e-22
C16586 _327_/a_27_7# _346_/SET_B 0.0401f
C16587 _317_/Q VPWR 0.887f
C16588 _162_/X _150_/C 0.00264f
C16589 _230_/a_27_7# VGND 0.0315f
C16590 _316_/a_1283_n19# _248_/A 1.22e-19
C16591 _205_/a_79_n19# VGND -0.00251f
C16592 _205_/a_297_7# VPWR -2.93e-19
C16593 ctln[6] _153_/B 0.603f
C16594 clkbuf_2_1_0_clk/A _199_/a_346_7# 8.1e-19
C16595 _163_/a_292_257# _160_/A 3.35e-20
C16596 _326_/a_27_7# _346_/SET_B 4.29e-21
C16597 _188_/S _228_/A 0.0495f
C16598 _226_/a_79_n19# _298_/X 6.92e-20
C16599 _343_/a_761_249# _175_/Y 0.00151f
C16600 _254_/B _202_/a_346_7# 0.0039f
C16601 clkbuf_2_3_0_clk/A _286_/B 0.303f
C16602 _342_/a_27_7# sample 0.0268f
C16603 _342_/a_761_249# _286_/Y 1.43e-20
C16604 _217_/a_27_7# _223_/a_93_n19# 2.37e-20
C16605 _333_/a_651_373# _192_/B 8.03e-20
C16606 _341_/Q _153_/A 0.00249f
C16607 _331_/Q _331_/a_1108_7# 0.0335f
C16608 _230_/a_27_7# _318_/a_1108_7# 0.00127f
C16609 _287_/a_121_257# _267_/B 0.00141f
C16610 _316_/a_543_7# _316_/D 3.87e-19
C16611 _316_/a_1283_n19# _331_/CLK 2.4e-20
C16612 _294_/A _306_/a_505_n19# 0.0186f
C16613 _149_/A _177_/a_27_7# 7.89e-19
C16614 _329_/a_27_7# _330_/D 0.0124f
C16615 clkbuf_0_clk/X _330_/a_543_7# 8.72e-20
C16616 repeater43/X _181_/X 0.135f
C16617 _279_/Y _332_/Q 0.00466f
C16618 _301_/a_149_7# VPWR -9.74e-19
C16619 _301_/a_245_257# VGND -6.83e-19
C16620 _320_/Q _236_/B 9.19e-21
C16621 _260_/B _190_/A 0.274f
C16622 _232_/A VGND 1.15f
C16623 _346_/SET_B _347_/a_639_7# -7.75e-19
C16624 cal _312_/a_27_7# 0.00373f
C16625 _258_/a_505_n19# _216_/A 1.1e-19
C16626 _321_/Q _234_/B 8.26e-20
C16627 _326_/a_543_7# _248_/A 9.84e-20
C16628 _200_/a_93_n19# _338_/Q 0.00787f
C16629 clk _333_/a_193_7# 7.42e-20
C16630 _327_/a_543_7# _331_/CLK 0.0302f
C16631 _321_/a_1283_n19# _321_/Q 0.0664f
C16632 _342_/Q _271_/A 0.0293f
C16633 _208_/a_292_257# _332_/Q 6.43e-21
C16634 _207_/X _204_/a_27_257# 2.15e-19
C16635 _208_/a_78_159# _333_/Q 0.0017f
C16636 _227_/A _314_/a_27_7# 1.17e-20
C16637 _286_/B _172_/Y 0.638f
C16638 repeater43/X _304_/a_288_7# 1.02e-19
C16639 _338_/a_543_7# _337_/a_543_7# 1.95e-20
C16640 _338_/a_1108_7# _337_/a_193_7# 3.35e-20
C16641 _318_/a_1108_7# _232_/A 8.18e-22
C16642 _326_/a_193_7# _236_/B 9.56e-22
C16643 _326_/a_543_7# _331_/CLK 5.68e-20
C16644 _234_/a_109_257# VGND -0.00128f
C16645 _315_/Q _248_/A 0.00803f
C16646 _341_/a_193_7# _343_/CLK 0.00432f
C16647 _258_/S _313_/a_193_7# 1.23e-20
C16648 _305_/a_76_159# _336_/D 6.63e-19
C16649 _277_/A _346_/D 0.00258f
C16650 _311_/a_1283_n19# _310_/a_27_7# 6.54e-19
C16651 _311_/a_761_249# _310_/a_761_249# 1.8e-21
C16652 _286_/B _313_/a_1270_373# 8.5e-21
C16653 _321_/a_761_249# VPWR 0.0314f
C16654 _321_/a_27_7# VGND -0.103f
C16655 _327_/a_543_7# _273_/A 1.12e-21
C16656 _277_/Y clkbuf_2_0_0_clk/a_75_172# 7.71e-19
C16657 output10/a_27_7# clkbuf_2_1_0_clk/A 0.0101f
C16658 _304_/a_257_159# _212_/X 1.5e-20
C16659 _338_/a_193_7# _343_/CLK 1.21e-19
C16660 _169_/B _299_/X 6.64e-19
C16661 _188_/S _216_/A 1.07e-19
C16662 _160_/A _173_/a_226_257# 5.09e-21
C16663 _215_/A _310_/D 1.93e-20
C16664 _315_/Q _331_/CLK 1.44e-20
C16665 _234_/B _318_/a_193_7# 0.0102f
C16666 _341_/a_1462_7# _341_/D 0.00186f
C16667 _328_/a_761_249# _331_/CLK 1.16e-21
C16668 _321_/a_193_7# _318_/a_1283_n19# 1.06e-20
C16669 _161_/Y _344_/D 0.123f
C16670 rstn VGND 1.94f
C16671 _232_/X _221_/a_256_7# 2.44e-19
C16672 output31/a_27_7# _311_/a_27_7# 1.11e-20
C16673 result[6] _322_/Q 2.35e-19
C16674 _164_/Y _160_/a_27_7# 5.6e-21
C16675 _332_/a_1462_7# _333_/Q 3.49e-19
C16676 _267_/A _254_/B 0.0249f
C16677 output8/a_27_7# _292_/A 3.84e-19
C16678 _340_/a_543_7# _337_/a_1108_7# 0.002f
C16679 _340_/a_1108_7# _337_/a_543_7# 0.002f
C16680 repeater43/X _343_/Q 0.0142f
C16681 _326_/a_193_7# _326_/D -0.0114f
C16682 _196_/A _157_/a_27_7# 0.0276f
C16683 _290_/A _171_/a_78_159# 0.00772f
C16684 _279_/Y _337_/a_193_7# 1.03e-20
C16685 _344_/a_193_7# _306_/S 5.65e-20
C16686 _329_/Q _319_/a_448_7# 5.12e-21
C16687 _238_/B _319_/a_1283_n19# 0.00111f
C16688 repeater43/X ctlp[1] 1.88e-20
C16689 _317_/D sample 0.00544f
C16690 _310_/a_1270_373# VPWR 1e-19
C16691 _310_/a_448_7# VGND 0.00326f
C16692 output15/a_27_7# output29/a_27_7# 3.1e-20
C16693 _325_/Q _246_/B 0.0099f
C16694 repeater43/X _332_/a_1283_n19# 0.0526f
C16695 _290_/Y _285_/Y 9.56e-19
C16696 output11/a_27_7# _343_/CLK 3.06e-19
C16697 _181_/X _191_/B 0.00811f
C16698 _286_/B _192_/B 0.238f
C16699 _165_/a_78_159# _158_/Y 0.0117f
C16700 _319_/Q _322_/a_1283_n19# 1.74e-21
C16701 output21/a_27_7# result[7] 7.2e-19
C16702 _185_/A _323_/a_193_7# 0.00993f
C16703 _294_/A _309_/a_1462_7# 0.00206f
C16704 _298_/C _207_/C 0.0615f
C16705 clkbuf_0_clk/X _331_/Q 4.53e-21
C16706 _172_/A _306_/S 0.019f
C16707 _346_/a_193_7# _346_/SET_B 0.325f
C16708 _182_/X _226_/X 0.00543f
C16709 _325_/a_27_7# _286_/B 9.4e-22
C16710 output10/a_27_7# ctln[4] 0.00177f
C16711 _325_/D _212_/X 4.69e-19
C16712 _225_/a_59_35# VGND 0.0419f
C16713 output27/a_27_7# _321_/a_27_7# 2.43e-21
C16714 _316_/Q _325_/Q 0.0172f
C16715 _347_/Q _314_/a_27_7# 1.13e-20
C16716 _339_/a_1283_n19# _338_/a_761_249# 8.55e-19
C16717 _339_/a_1108_7# _338_/a_193_7# 5.12e-19
C16718 _271_/A _204_/Y 0.0087f
C16719 repeater43/a_27_7# _334_/a_193_7# 0.00341f
C16720 _309_/a_1283_n19# _310_/a_1283_n19# 0.00161f
C16721 _198_/a_256_7# _340_/Q 0.00124f
C16722 _198_/a_93_n19# _193_/Y 0.0577f
C16723 _294_/A _285_/A 0.0489f
C16724 _335_/a_193_7# _335_/Q 0.0138f
C16725 _335_/a_27_7# _204_/Y 2.52e-20
C16726 _281_/Y _197_/X 0.0956f
C16727 _321_/a_1108_7# _246_/B 3.41e-20
C16728 _323_/Q _298_/X 0.103f
C16729 _324_/Q _231_/a_512_7# 1.66e-19
C16730 _243_/a_199_7# VGND 1.21e-19
C16731 _299_/X _170_/a_226_7# 0.00857f
C16732 _347_/Q _170_/a_76_159# 1.01e-19
C16733 _324_/a_27_7# _215_/A 2.04e-20
C16734 _327_/a_1217_7# _346_/SET_B 7.36e-19
C16735 _324_/a_1270_373# _326_/Q 3.8e-20
C16736 _309_/D _312_/Q 3.27e-20
C16737 _325_/a_193_7# _304_/a_257_159# 1.2e-20
C16738 _334_/Q _332_/a_1283_n19# 5.27e-19
C16739 repeater43/X _341_/a_651_373# 7.07e-21
C16740 clkbuf_2_3_0_clk/A _338_/a_1108_7# 9.92e-22
C16741 _271_/A _298_/a_181_7# 3.8e-19
C16742 _256_/a_80_n19# clkbuf_0_clk/a_110_7# 9.1e-20
C16743 _343_/Q _191_/B 1.05e-19
C16744 _165_/a_215_7# _345_/Q 0.00196f
C16745 _340_/a_1283_n19# _339_/a_1283_n19# 0.00114f
C16746 _226_/X valid 1.36e-19
C16747 _342_/a_1217_7# sample 1.2e-20
C16748 _342_/D output30/a_27_7# 0.00437f
C16749 _190_/A _295_/a_512_7# 0.0438f
C16750 _242_/A _318_/a_805_7# 4.25e-19
C16751 _157_/a_27_7# _347_/a_1283_n19# 4.92e-21
C16752 output22/a_27_7# _304_/S 1.37e-19
C16753 clkbuf_2_1_0_clk/A _347_/Q 3.06e-19
C16754 _279_/Y _339_/a_193_7# 2.28e-19
C16755 _315_/a_193_7# VPWR -0.295f
C16756 trimb[0] trimb[1] 0.0574f
C16757 result[3] result[4] 0.0661f
C16758 _298_/A VPWR 2.67f
C16759 _149_/a_27_7# _177_/A 0.0303f
C16760 _342_/Q _186_/a_79_n19# 0.059f
C16761 _298_/C _150_/C 7.27e-19
C16762 _338_/Q _340_/CLK 0.518f
C16763 _336_/a_448_7# VPWR -0.00265f
C16764 _181_/X _331_/a_448_7# 7.28e-19
C16765 _324_/a_1283_n19# _227_/A 3.53e-20
C16766 _336_/a_1283_n19# VGND 0.024f
C16767 _346_/a_1182_221# _273_/A 5.64e-20
C16768 _332_/a_1283_n19# _191_/B 1.05e-20
C16769 _328_/a_805_7# _346_/SET_B -0.00125f
C16770 _324_/a_27_7# _324_/a_761_249# -0.0166f
C16771 _317_/a_27_7# _316_/a_27_7# 3e-19
C16772 input1/X _312_/a_805_7# 4.33e-20
C16773 _313_/Q _216_/A 0.0219f
C16774 _334_/a_27_7# _343_/CLK 0.0214f
C16775 repeater43/X _229_/a_76_159# 0.0128f
C16776 _315_/D _314_/a_761_249# 0.0231f
C16777 _333_/Q _190_/A 0.597f
C16778 _275_/A _347_/D 3.62e-19
C16779 _294_/A _172_/A 5.74e-19
C16780 _216_/X _144_/A 0.00133f
C16781 trimb[0] VGND 0.205f
C16782 _343_/a_805_7# _298_/A 5.75e-21
C16783 _345_/a_193_7# _277_/Y 3.31e-20
C16784 _346_/SET_B _319_/a_193_7# 0.0245f
C16785 _338_/D _337_/a_27_7# 1.93e-19
C16786 _194_/X _254_/B 0.0171f
C16787 _216_/X _331_/a_27_7# 6.49e-19
C16788 _324_/a_27_7# _304_/X 0.00881f
C16789 _314_/a_27_7# _297_/B 0.0389f
C16790 _255_/X _153_/B 3.06e-20
C16791 _321_/a_1217_7# VGND -5.03e-19
C16792 _324_/Q _223_/a_93_n19# 2.29e-19
C16793 rstn _335_/a_651_373# 8.98e-19
C16794 _338_/a_1462_7# _343_/CLK 1.47e-19
C16795 repeater43/X _204_/a_27_7# 1.74e-19
C16796 _341_/a_761_249# _145_/A 4.5e-20
C16797 _322_/a_193_7# _269_/A 0.0193f
C16798 repeater43/X _208_/a_215_7# 0.0537f
C16799 _279_/Y _327_/Q 5.94e-19
C16800 _325_/a_193_7# _325_/D 0.513f
C16801 _320_/Q _331_/a_193_7# 2.1e-21
C16802 _297_/B _170_/a_76_159# 1.17e-20
C16803 _238_/B _212_/X 1.21e-20
C16804 _232_/X _327_/D 0.0192f
C16805 _329_/a_1108_7# _232_/X 5.23e-20
C16806 _265_/B _311_/a_1108_7# 4.35e-20
C16807 _327_/a_1108_7# _327_/Q 0.00914f
C16808 _327_/a_543_7# _217_/X 0.00155f
C16809 _246_/B _326_/Q 0.59f
C16810 clkbuf_2_0_0_clk/a_75_172# VGND 0.0547f
C16811 _326_/a_651_373# repeater43/X 0.00205f
C16812 _275_/Y _310_/a_805_7# 3.81e-19
C16813 _290_/A _172_/B 0.429f
C16814 _326_/a_761_249# _331_/a_27_7# 9.17e-22
C16815 _326_/a_193_7# _331_/a_193_7# 1.65e-20
C16816 _326_/a_543_7# _217_/X 0.0299f
C16817 _326_/a_1283_n19# _212_/X 7.49e-21
C16818 clkbuf_2_1_0_clk/A _297_/B 0.00767f
C16819 _310_/D VGND 0.0996f
C16820 input4/X _332_/D 4.27e-20
C16821 _188_/a_439_7# _341_/D 6.45e-20
C16822 _281_/Y _330_/a_1108_7# 2.03e-20
C16823 _286_/B _146_/C 5.82e-23
C16824 _275_/Y _265_/B 0.0156f
C16825 _172_/A _283_/A 0.00746f
C16826 _345_/a_193_7# _345_/a_476_7# -2.46e-20
C16827 _306_/X _193_/Y 4.89e-22
C16828 _334_/Q _204_/a_27_7# 0.0018f
C16829 _342_/a_761_249# _269_/A 0.00206f
C16830 _341_/a_1283_n19# _149_/a_27_7# 9.5e-19
C16831 _343_/CLK _207_/X 0.00844f
C16832 _300_/a_301_257# VPWR 0.0385f
C16833 _281_/Y _333_/a_193_7# 3.05e-20
C16834 output12/a_27_7# _333_/a_1108_7# 4.49e-19
C16835 _328_/a_761_249# _217_/X 2.3e-19
C16836 _328_/a_543_7# _212_/X 0.0111f
C16837 _302_/a_77_159# _347_/a_651_373# 1.39e-19
C16838 _302_/a_227_7# _347_/a_543_7# 2.68e-20
C16839 _157_/A _286_/B 0.0113f
C16840 _284_/a_121_257# VPWR 2.67e-19
C16841 _211_/a_109_257# _283_/A 0.00202f
C16842 _346_/a_796_7# _346_/SET_B 0.00126f
C16843 output8/a_27_7# _273_/A 0.00233f
C16844 _232_/X _283_/A 0.0362f
C16845 _255_/B _179_/a_27_7# 0.00763f
C16846 _325_/a_639_7# _181_/X 0.00105f
C16847 output13/a_27_7# rstn 0.0135f
C16848 _283_/Y input4/a_27_7# 0.00125f
C16849 _339_/a_27_7# _338_/D 2.44e-20
C16850 trim[2] _312_/a_27_7# 2.83e-20
C16851 _279_/Y _192_/B 6.73e-19
C16852 _340_/CLK _313_/a_1108_7# 3.88e-21
C16853 _229_/a_226_7# _226_/X 0.0178f
C16854 repeater43/X _334_/a_448_7# 0.00442f
C16855 _337_/a_639_7# _340_/CLK 0.00434f
C16856 result[1] _315_/a_761_249# 1.27e-19
C16857 _316_/Q _315_/a_1283_n19# 0.0034f
C16858 _335_/a_1462_7# _335_/Q 2.71e-19
C16859 _235_/a_113_257# _321_/Q 0.00403f
C16860 _215_/A VPWR 3.9f
C16861 _342_/a_1283_n19# _185_/A 1.68e-21
C16862 _164_/A _344_/Q 0.182f
C16863 _172_/A _248_/B 1.77e-21
C16864 _255_/X _305_/a_505_n19# 5.46e-21
C16865 _277_/Y VPWR 1.45f
C16866 clkbuf_1_0_0_clk/a_75_172# _330_/a_761_249# 0.00105f
C16867 _260_/B clkbuf_0_clk/a_110_7# 5.48e-20
C16868 _345_/a_652_n19# _160_/X 5.9e-20
C16869 _271_/A en 0.00643f
C16870 _344_/a_381_7# _297_/Y 0.0146f
C16871 _309_/a_193_7# _284_/a_39_257# 7.16e-20
C16872 _286_/B _202_/a_584_7# 2.11e-19
C16873 ctlp[1] result[6] 3e-19
C16874 _184_/a_505_n19# _298_/A 3.73e-20
C16875 _254_/A _340_/CLK 5.73e-20
C16876 _340_/a_761_249# _339_/D 8.19e-21
C16877 repeater43/X _346_/SET_B 0.00367f
C16878 _237_/a_199_7# clkbuf_0_clk/X 2.41e-19
C16879 _290_/A _289_/a_121_257# 4.18e-19
C16880 _164_/Y _267_/A 0.169f
C16881 _232_/X _248_/B 0.00109f
C16882 _313_/D _257_/a_222_53# 1.91e-19
C16883 _315_/a_805_7# VGND 1.45e-19
C16884 _315_/a_1462_7# VPWR 1.96e-19
C16885 _183_/a_471_7# _298_/C 9.95e-19
C16886 _282_/a_39_257# _316_/D 0.00101f
C16887 _288_/A _284_/A 0.0365f
C16888 _182_/X input1/X 0.0258f
C16889 trimb[3] VGND 0.229f
C16890 _340_/a_27_7# _202_/a_93_n19# 2.29e-20
C16891 _324_/a_27_7# VGND -0.0862f
C16892 _274_/a_121_257# _217_/X 4.18e-19
C16893 _324_/a_761_249# VPWR 0.00181f
C16894 _342_/a_543_7# _342_/Q 1.59e-19
C16895 _254_/Y _172_/A 1.9e-20
C16896 _309_/a_27_7# _215_/A 0.0132f
C16897 _262_/a_199_7# VPWR -2.88e-19
C16898 _330_/Q _217_/A 0.00486f
C16899 _326_/a_193_7# _325_/a_1283_n19# 3.09e-20
C16900 _346_/a_1602_7# clkbuf_2_3_0_clk/A 0.00601f
C16901 _162_/X _284_/A 0.00726f
C16902 _188_/a_76_159# repeater43/X 2.54e-20
C16903 _318_/a_1283_n19# _242_/B 4.8e-19
C16904 _318_/a_761_249# _318_/D 6.55e-19
C16905 _329_/a_1283_n19# _318_/Q 4.85e-21
C16906 _286_/B _260_/A 0.0179f
C16907 _287_/a_39_257# _284_/A 6.79e-20
C16908 _277_/Y _309_/a_27_7# 1.09e-19
C16909 ctln[1] _334_/a_1283_n19# 3.76e-19
C16910 _314_/a_651_373# VGND 0.00142f
C16911 _314_/a_639_7# VPWR 6.67e-19
C16912 _346_/SET_B _319_/a_1462_7# -9.14e-19
C16913 _324_/a_1283_n19# _297_/B 1.43e-21
C16914 _346_/SET_B _313_/a_448_7# 0.00153f
C16915 _343_/a_193_7# VPWR 0.0227f
C16916 _340_/a_27_7# cal 4.31e-20
C16917 _346_/SET_B _337_/a_805_7# -0.00125f
C16918 _338_/a_651_373# _337_/Q 4.11e-20
C16919 _193_/Y _147_/Y 3.48e-19
C16920 _248_/A _212_/X 0.0108f
C16921 _307_/X _180_/a_29_13# 1.02e-20
C16922 clk _332_/a_651_373# 0.0174f
C16923 _304_/X VPWR 0.598f
C16924 _157_/A _347_/a_543_7# 0.00408f
C16925 _324_/a_1270_373# _324_/D 3.05e-19
C16926 _340_/a_27_7# _197_/a_27_7# 0.00852f
C16927 _283_/Y _204_/Y 2.54e-20
C16928 _216_/A _223_/a_93_n19# 0.0311f
C16929 _293_/a_121_257# _336_/a_193_7# 1.19e-20
C16930 _331_/CLK _212_/X 0.0783f
C16931 _316_/D _327_/Q 0.00956f
C16932 input1/X valid 7.35e-20
C16933 _345_/a_476_7# VPWR 0.0598f
C16934 _345_/a_193_7# VGND 0.0172f
C16935 _309_/D _340_/CLK 0.72f
C16936 _259_/a_113_257# _261_/A 0.0424f
C16937 _308_/S _209_/a_373_7# 2.38e-20
C16938 _308_/S _336_/Q 1.35e-20
C16939 _196_/A _267_/A 0.0561f
C16940 _162_/A _174_/a_27_257# 7.92e-20
C16941 _266_/a_113_257# VGND 0.00209f
C16942 _341_/a_1108_7# _146_/C 4.02e-21
C16943 cal _298_/C 0.512f
C16944 _297_/B _278_/a_68_257# 9.35e-22
C16945 _345_/a_1032_373# _297_/B 1.09e-19
C16946 _248_/B _244_/B 0.018f
C16947 _273_/A _212_/X 0.244f
C16948 _275_/Y _310_/Q 0.0122f
C16949 _339_/a_27_7# _337_/a_1108_7# 8.22e-19
C16950 _339_/a_193_7# _337_/a_1283_n19# 0.00304f
C16951 _339_/a_1108_7# _337_/a_27_7# 8.22e-19
C16952 _339_/a_1283_n19# _337_/a_193_7# 0.00304f
C16953 _172_/A _169_/a_109_257# 0.00306f
C16954 _272_/a_121_257# _330_/Q 2.89e-21
C16955 _235_/a_199_7# _246_/B 1.42e-19
C16956 _341_/a_761_249# _324_/Q 7.52e-20
C16957 output24/a_27_7# result[3] 2.55e-19
C16958 result[2] output25/a_27_7# 2.55e-19
C16959 _277_/A _320_/a_448_7# 0.00162f
C16960 _318_/Q _230_/a_27_7# 1.5e-19
C16961 _339_/a_27_7# _343_/CLK 1.49e-20
C16962 _254_/Y _203_/a_80_n19# 3.92e-20
C16963 _222_/a_93_n19# _212_/X 0.0736f
C16964 _222_/a_250_257# _327_/Q 6.75e-20
C16965 _308_/X _175_/Y 1.1e-19
C16966 _200_/a_250_257# cal 0.0301f
C16967 _200_/a_93_n19# input1/X 0.00391f
C16968 _245_/a_113_257# VGND 2.98e-19
C16969 _272_/a_39_257# VPWR 0.0326f
C16970 input4/X _207_/C 3.46e-19
C16971 repeater43/X _206_/A 1.04f
C16972 _342_/a_27_7# _175_/Y 2.5e-19
C16973 _300_/Y VPWR 0.159f
C16974 _329_/a_193_7# _331_/Q 2.53e-19
C16975 _322_/a_543_7# _322_/D 2.39e-19
C16976 _322_/a_1108_7# _234_/B 3.52e-19
C16977 _338_/Q _267_/B 0.72f
C16978 valid _286_/Y 8.35e-19
C16979 output12/a_27_7# _332_/a_27_7# 6.84e-20
C16980 _255_/B _231_/a_306_7# 8.57e-19
C16981 _210_/a_27_7# _254_/B 0.0669f
C16982 _339_/a_805_7# _346_/SET_B -0.00123f
C16983 _220_/a_93_n19# VPWR 0.0118f
C16984 _318_/Q _232_/A 2.97e-20
C16985 _320_/Q _219_/a_93_n19# 5.25e-20
C16986 _183_/a_27_7# _295_/a_79_n19# 2.57e-21
C16987 repeater43/X _334_/D 0.448f
C16988 _188_/a_535_334# _307_/X 1.86e-19
C16989 _164_/A _306_/S 1.2e-20
C16990 _325_/a_193_7# _248_/A 0.0127f
C16991 _231_/a_79_n19# _144_/a_27_7# 2.22e-20
C16992 _290_/A trimb[4] 3e-20
C16993 clk _295_/a_79_n19# 0.00109f
C16994 _254_/a_109_257# clkbuf_2_3_0_clk/A 0.00244f
C16995 ctln[1] repeater43/a_27_7# 1.44e-19
C16996 ctln[4] _275_/Y 1.83e-20
C16997 _277_/Y ctln[3] 4.28e-20
C16998 output7/a_27_7# repeater43/X 0.0708f
C16999 _324_/Q _216_/X 0.0147f
C17000 _166_/Y _299_/a_215_7# 0.00202f
C17001 _324_/Q _316_/a_543_7# 0.00232f
C17002 _279_/Y _157_/A 0.0408f
C17003 _187_/a_27_7# _271_/A 8.87e-20
C17004 _228_/A _347_/a_27_7# 2.48e-22
C17005 _313_/a_193_7# _313_/a_651_373# -0.00701f
C17006 _149_/a_27_7# _248_/A 4.47e-19
C17007 _271_/A _315_/D 0.0104f
C17008 _289_/a_39_257# _297_/Y 0.00114f
C17009 _325_/a_193_7# _331_/CLK 0.00589f
C17010 _325_/a_27_7# _316_/D 1.58e-21
C17011 trimb[1] VPWR 0.178f
C17012 _320_/a_193_7# clkbuf_2_1_0_clk/A 2.39e-20
C17013 _334_/Q _206_/A 0.0147f
C17014 _332_/a_193_7# _207_/a_27_7# 3.43e-19
C17015 _327_/a_1270_373# clkbuf_0_clk/X 3.61e-19
C17016 _306_/S _192_/a_68_257# 7.09e-20
C17017 _273_/A _325_/a_193_7# 6.91e-20
C17018 _328_/a_27_7# _219_/a_93_n19# 0.00285f
C17019 _161_/Y _265_/B 3e-19
C17020 VPWR VGND 4.77f
C17021 _254_/A _313_/a_543_7# 5.81e-19
C17022 _324_/a_1217_7# VGND -3.95e-19
C17023 _313_/a_193_7# _157_/a_27_7# 8.95e-19
C17024 result[0] _146_/C 1.24e-20
C17025 _236_/B _317_/a_1283_n19# 2.84e-19
C17026 _317_/a_1108_7# _316_/D 2.97e-20
C17027 _317_/a_448_7# _331_/CLK 1.16e-20
C17028 _338_/a_193_7# _195_/a_109_257# 6.68e-20
C17029 repeater43/X _147_/A 0.00194f
C17030 _334_/D _334_/Q 0.454f
C17031 cal _229_/a_489_373# 4.36e-19
C17032 input1/X _229_/a_226_7# 0.00124f
C17033 _188_/S _224_/a_93_n19# 3.1e-20
C17034 _285_/A _284_/a_39_257# 0.0332f
C17035 _183_/a_27_7# _180_/a_29_13# 3.3e-19
C17036 _175_/Y _254_/B 1.26e-20
C17037 _318_/a_1108_7# VPWR 0.0146f
C17038 _318_/a_543_7# VGND 0.00482f
C17039 _343_/a_1462_7# VPWR 3.62e-19
C17040 _343_/a_805_7# VGND 2.44e-19
C17041 _191_/B _206_/A 1.75f
C17042 _346_/a_652_n19# _276_/a_68_257# 1.47e-21
C17043 _341_/a_761_249# _228_/A 0.00111f
C17044 _175_/Y _317_/D 1.61e-20
C17045 _286_/B _340_/Q 0.00216f
C17046 repeater43/X _149_/A 0.0343f
C17047 _325_/a_193_7# _222_/a_93_n19# 9.34e-19
C17048 _325_/a_27_7# _222_/a_250_257# 2.53e-19
C17049 _346_/SET_B _337_/Q 0.173f
C17050 ctlp[6] VGND 0.125f
C17051 clkbuf_0_clk/X _347_/D 2e-20
C17052 _346_/a_27_7# _301_/X 1.07e-19
C17053 _314_/D _314_/Q 3.43e-21
C17054 _294_/A _164_/A 7.75e-19
C17055 _307_/a_76_159# _296_/Y 0.0095f
C17056 _318_/a_193_7# _318_/a_651_373# -0.00701f
C17057 _292_/A _344_/Q 0.371f
C17058 _309_/a_761_249# VPWR 0.0232f
C17059 _309_/a_27_7# VGND -0.0942f
C17060 _313_/a_448_7# _147_/A 0.0282f
C17061 _298_/C _284_/A 2.09e-19
C17062 _334_/D _191_/B 8.6e-20
C17063 _343_/CLK _323_/Q 1.66e-19
C17064 _254_/A _304_/S 2.27e-20
C17065 _341_/a_1270_373# _286_/Y 2.49e-19
C17066 _279_/Y _260_/A 0.00995f
C17067 _305_/a_218_334# _225_/B 0.0013f
C17068 _345_/a_796_7# VGND 2.15e-19
C17069 _345_/a_1224_7# VPWR 7.19e-20
C17070 _216_/X _281_/A 0.00249f
C17071 _281_/Y _340_/a_193_7# 9.32e-21
C17072 _258_/a_505_n19# _300_/a_383_7# 2.1e-21
C17073 _292_/Y ctlp[2] 8.52e-20
C17074 _315_/a_27_7# _244_/B 0.0171f
C17075 _307_/a_218_7# _191_/B 2.46e-19
C17076 _160_/A _344_/Q 0.00642f
C17077 _301_/a_149_7# _147_/Y 3.58e-19
C17078 _336_/a_543_7# _254_/B 1.68e-19
C17079 _197_/X _199_/a_93_n19# 0.0415f
C17080 clk _334_/a_639_7# 4.17e-19
C17081 _329_/Q _281_/A 0.00288f
C17082 _172_/A _298_/B 0.00793f
C17083 _308_/X _341_/Q 0.0116f
C17084 _165_/X _286_/B 0.00643f
C17085 _167_/X _196_/A 2.22e-19
C17086 _326_/D _331_/a_651_373# 3.38e-20
C17087 _216_/X _228_/A 0.07f
C17088 _311_/a_193_7# _311_/a_1283_n19# -7.11e-33
C17089 repeater43/X _331_/a_761_249# 0.0133f
C17090 _277_/Y _344_/a_27_7# 7.15e-21
C17091 _191_/a_109_257# _191_/B 0.00102f
C17092 _283_/A _333_/a_448_7# 0.0227f
C17093 _316_/a_543_7# _228_/A 1.61e-21
C17094 output27/a_27_7# VPWR 0.0997f
C17095 _229_/a_226_7# _286_/Y 2.84e-20
C17096 _309_/a_27_7# _309_/a_761_249# -0.0166f
C17097 _255_/a_184_257# _286_/B 0.00154f
C17098 _255_/a_30_13# _181_/X 0.0058f
C17099 input1/X _340_/CLK 0.085f
C17100 _331_/a_27_7# _327_/Q 7.33e-20
C17101 _298_/B _335_/D 1.18e-20
C17102 _285_/A _262_/a_113_257# 1.36e-20
C17103 _212_/X _217_/X 0.727f
C17104 _306_/S _333_/D 0.128f
C17105 _197_/X _336_/Q 0.268f
C17106 _333_/a_27_7# _204_/Y 0.00132f
C17107 _333_/a_193_7# _335_/Q 3.67e-19
C17108 _191_/B _147_/A 0.955f
C17109 _308_/a_218_7# VGND 2.27e-20
C17110 _306_/S _332_/a_193_7# 2.71e-21
C17111 _275_/Y _311_/a_27_7# 0.0081f
C17112 _327_/a_27_7# _319_/Q 3.58e-20
C17113 _149_/A _191_/B 6.44e-20
C17114 _343_/a_1108_7# _323_/a_193_7# 3.74e-21
C17115 _343_/a_193_7# _323_/a_1108_7# 1.02e-20
C17116 _154_/a_27_7# _154_/A 0.0569f
C17117 _328_/a_193_7# _281_/A 4.24e-21
C17118 _306_/a_76_159# VGND -0.00714f
C17119 _306_/a_218_334# VPWR -0.0017f
C17120 _342_/Q _162_/X 0.00641f
C17121 _251_/X _286_/B 1.37e-21
C17122 _146_/C _316_/D 2.32e-20
C17123 _339_/Q _346_/SET_B 0.0296f
C17124 _225_/X _226_/X 4.27e-19
C17125 _317_/Q _223_/a_250_257# 3.84e-19
C17126 _311_/a_651_373# VGND 9.28e-19
C17127 _311_/a_639_7# VPWR 0.00344f
C17128 _162_/X _144_/a_27_7# 0.0101f
C17129 _181_/X _296_/a_493_257# 2.86e-19
C17130 clkbuf_2_1_0_clk/A _161_/Y 2.09e-21
C17131 _179_/a_27_7# _154_/A 3.03e-20
C17132 _216_/X _216_/A 0.624f
C17133 _346_/SET_B _202_/a_256_7# 0.00162f
C17134 _297_/B _328_/D 9.33e-19
C17135 _297_/A _248_/B 0.21f
C17136 _324_/a_193_7# _172_/A 1.1e-21
C17137 _335_/a_27_7# _335_/a_193_7# -0.296f
C17138 _217_/a_27_7# _327_/Q 0.0337f
C17139 _232_/X _242_/B 0.00167f
C17140 _345_/a_476_7# _344_/a_27_7# 1.68e-22
C17141 _345_/a_27_7# _344_/a_476_7# 0.00128f
C17142 _328_/a_1283_n19# _239_/a_113_257# 3.06e-20
C17143 _288_/A _310_/a_761_249# 2.92e-21
C17144 trim[1] _310_/a_27_7# 5.45e-21
C17145 _335_/a_651_373# VPWR -0.00901f
C17146 _335_/a_1108_7# VGND 0.00185f
C17147 _279_/Y _221_/a_250_257# 6.22e-20
C17148 _197_/X _336_/a_805_7# 1.48e-19
C17149 _184_/a_535_334# VPWR -7.81e-19
C17150 _184_/a_505_n19# VGND 0.0833f
C17151 _309_/a_193_7# _306_/a_505_n19# 2.41e-20
C17152 ctln[3] VGND 0.0752f
C17153 _267_/B _309_/D 0.163f
C17154 _341_/Q _254_/B 0.0245f
C17155 _347_/D _286_/Y 3.63e-20
C17156 _341_/Q _317_/D 0.00141f
C17157 _237_/a_199_7# _328_/Q 2.26e-19
C17158 _340_/D _194_/A 1.47e-20
C17159 output14/a_27_7# _269_/A 0.0318f
C17160 _303_/A _346_/SET_B 0.00263f
C17161 _320_/a_27_7# _279_/A 1.96e-20
C17162 _340_/a_639_7# _336_/D 7.09e-21
C17163 _326_/a_761_249# _216_/A 1.47e-19
C17164 _338_/a_448_7# _194_/X 8.94e-19
C17165 _333_/a_1283_n19# _153_/a_109_53# 0.00488f
C17166 _285_/A _160_/X 0.0173f
C17167 _219_/a_250_257# _319_/a_193_7# 8.34e-20
C17168 _325_/a_1108_7# repeater43/X -0.00933f
C17169 _209_/X _333_/a_543_7# 2.92e-20
C17170 _188_/S _217_/A 5.08e-20
C17171 _283_/A _312_/D 0.00155f
C17172 _302_/a_323_257# _147_/A 8.77e-19
C17173 _325_/a_761_249# _212_/X 0.00323f
C17174 _325_/a_193_7# _217_/X 8.75e-20
C17175 _325_/a_543_7# _327_/Q 4.35e-20
C17176 _344_/a_193_7# _160_/X 4.1e-20
C17177 _304_/a_257_159# _283_/A 9.12e-19
C17178 _157_/A _313_/a_27_7# 8.02e-19
C17179 _212_/a_27_7# _217_/A 0.00257f
C17180 _309_/a_1217_7# VGND -4.44e-19
C17181 repeater43/X _317_/a_805_7# 0.00163f
C17182 _340_/a_448_7# _306_/S 7.93e-20
C17183 _340_/a_651_373# _340_/Q 9.07e-20
C17184 _340_/a_543_7# _340_/D 0.00108f
C17185 _340_/a_1108_7# _193_/Y 2.43e-19
C17186 _337_/Q _147_/A 1.24e-20
C17187 _244_/B _242_/B 4.64e-20
C17188 _227_/A _203_/a_303_7# 2.19e-20
C17189 _324_/Q _216_/a_27_7# 0.00243f
C17190 _315_/a_639_7# _317_/D 0.00112f
C17191 _279_/Y _340_/Q 1.44e-20
C17192 output11/a_27_7# _340_/D 1.32e-19
C17193 _269_/A valid 0.19f
C17194 _145_/A _192_/B 2.63e-21
C17195 _336_/a_448_7# _147_/Y 0.0251f
C17196 clkbuf_2_2_0_clk/a_75_172# cal 2.6e-19
C17197 clkbuf_2_3_0_clk/A input1/a_75_172# 0.0147f
C17198 _322_/a_27_7# _321_/Q 0.0061f
C17199 _172_/A _160_/X 0.0113f
C17200 output13/a_27_7# VPWR 0.123f
C17201 _333_/a_1283_n19# _209_/a_27_257# 0.00129f
C17202 _271_/A _323_/a_193_7# 1.21e-20
C17203 _339_/Q _337_/a_448_7# 0.0185f
C17204 _346_/a_652_n19# _346_/Q 3.87e-19
C17205 _346_/a_27_7# _166_/Y 1.11e-19
C17206 output12/a_27_7# _333_/Q 1.19e-19
C17207 _283_/A _333_/D 0.193f
C17208 output29/a_27_7# result[7] 0.00541f
C17209 _325_/a_193_7# _296_/Y 9.31e-21
C17210 _304_/a_257_159# _248_/B 0.0943f
C17211 _188_/a_505_n19# _286_/Y 0.052f
C17212 _306_/X _215_/A 3.52e-21
C17213 clkbuf_0_clk/X _304_/S 0.011f
C17214 _320_/a_1108_7# VPWR 0.015f
C17215 _320_/a_543_7# VGND 0.0348f
C17216 _273_/A _344_/Q 0.0162f
C17217 output35/a_27_7# _284_/A 0.00246f
C17218 _343_/D valid 2.22e-19
C17219 _323_/a_651_373# VPWR 0.00257f
C17220 _323_/a_1108_7# VGND 0.00923f
C17221 _283_/A _332_/a_193_7# 2.88e-20
C17222 _248_/B _177_/A 3.63e-20
C17223 _322_/a_193_7# _318_/a_27_7# 4.51e-21
C17224 _322_/a_27_7# _318_/a_193_7# 1.14e-20
C17225 _214_/a_27_257# VPWR 0.081f
C17226 _344_/a_27_7# VGND 0.0178f
C17227 _344_/a_652_n19# VPWR 0.0095f
C17228 cal _207_/C 0.193f
C17229 input1/X _313_/a_543_7# 1.6e-20
C17230 _294_/A _292_/A 0.147f
C17231 _320_/a_651_373# _297_/B 8.49e-19
C17232 _283_/A _325_/D 0.00946f
C17233 _186_/a_382_257# _271_/A 2.25e-19
C17234 _207_/a_109_7# _333_/Q 5.36e-19
C17235 _345_/a_1032_373# _161_/Y 0.00386f
C17236 _343_/a_27_7# _323_/D 0.0144f
C17237 _149_/a_27_7# _146_/a_29_271# 1.94e-21
C17238 _183_/a_471_7# _150_/C 0.137f
C17239 _324_/a_27_7# _318_/Q 1.07e-21
C17240 ctln[6] _340_/CLK 0.00708f
C17241 _344_/a_1182_221# _297_/B 8.68e-22
C17242 _260_/A _313_/a_27_7# 6.45e-20
C17243 _294_/A _160_/A 3.63e-20
C17244 _294_/Y _162_/A 1.07f
C17245 _285_/A _309_/a_193_7# 9.05e-20
C17246 _258_/a_218_334# VGND -4.43e-19
C17247 _258_/a_218_7# VPWR -2.54e-19
C17248 _325_/a_27_7# _325_/a_543_7# -0.00936f
C17249 _325_/a_193_7# _325_/a_761_249# -0.0105f
C17250 _346_/SET_B _336_/D 0.0196f
C17251 _184_/a_76_159# _184_/a_218_7# -8.88e-34
C17252 _265_/B _263_/B 2.04e-20
C17253 _346_/Q _173_/a_226_7# 5.42e-20
C17254 _146_/C _144_/A 0.00965f
C17255 _337_/D _337_/Q 0.075f
C17256 _211_/a_109_7# VPWR 1.5e-19
C17257 _211_/a_27_257# VGND -0.00794f
C17258 output32/a_27_7# _310_/D 2.39e-19
C17259 _342_/Q _298_/C 0.0547f
C17260 _254_/A _301_/X 0.682f
C17261 _279_/Y _251_/X 2.68e-20
C17262 _222_/a_584_7# _286_/Y 2.09e-19
C17263 _198_/a_256_7# VPWR -6.42e-19
C17264 _198_/a_93_n19# VGND 0.00256f
C17265 output15/a_27_7# _234_/B 3.12e-21
C17266 _245_/a_199_7# _244_/B 7.84e-19
C17267 _267_/A _313_/a_193_7# 4.65e-20
C17268 _343_/a_1108_7# _342_/a_1283_n19# 8.59e-22
C17269 _248_/B _325_/D 1.16e-21
C17270 output17/a_27_7# clkbuf_2_1_0_clk/A 7.55e-19
C17271 output15/a_27_7# _321_/a_1283_n19# 1.75e-19
C17272 _216_/a_27_7# _228_/A 6.73e-19
C17273 _319_/Q _319_/a_193_7# 0.004f
C17274 _157_/A _144_/A 4.06e-20
C17275 _339_/a_448_7# _339_/Q 2.2e-20
C17276 output33/a_27_7# _273_/A 0.02f
C17277 _286_/B _225_/a_59_35# 1.55e-19
C17278 _242_/B _241_/a_113_257# 0.00671f
C17279 _232_/X _318_/a_1283_n19# 1.24e-20
C17280 _309_/a_193_7# _172_/A 6.93e-19
C17281 _171_/a_215_7# VGND 0.0301f
C17282 _338_/D _194_/X 0.0121f
C17283 _333_/a_1283_n19# _153_/A 0.0101f
C17284 _224_/a_93_n19# _223_/a_93_n19# 5.13e-19
C17285 cal _150_/C 0.00653f
C17286 _196_/A _175_/Y 9.43e-19
C17287 _307_/X input1/X 1.9e-20
C17288 _323_/a_27_7# _323_/a_193_7# -0.163f
C17289 ctlp[5] VPWR 0.0908f
C17290 _215_/A _147_/Y 0.0272f
C17291 repeater42/a_27_7# _232_/X 0.0105f
C17292 _275_/A _281_/Y 7.01e-21
C17293 _303_/A _147_/A 6.09e-19
C17294 _169_/Y _162_/X 0.0202f
C17295 _269_/A _229_/a_226_7# 4.98e-20
C17296 _277_/Y _147_/Y 0.017f
C17297 _162_/X _225_/B 0.00355f
C17298 _343_/CLK sample 0.229f
C17299 input1/X _267_/B 1.47e-20
C17300 _341_/a_1283_n19# _248_/B 8.11e-22
C17301 _275_/A _166_/Y 1.72e-19
C17302 _328_/Q _347_/D 2.04e-20
C17303 _328_/a_651_373# _328_/Q 1.4e-19
C17304 _346_/a_1032_373# _306_/S 3.24e-36
C17305 _150_/C _150_/a_193_257# 1.89e-19
C17306 _304_/S _286_/Y 0.00933f
C17307 _283_/Y _335_/a_193_7# 3.53e-19
C17308 _317_/Q _316_/a_1283_n19# 5.76e-19
C17309 result[2] _316_/a_761_249# 9.25e-19
C17310 _309_/a_1108_7# _171_/a_78_159# 1.18e-20
C17311 _203_/a_209_257# VPWR -0.00479f
C17312 _286_/B _336_/a_1283_n19# 0.00413f
C17313 _242_/A _316_/a_27_7# 1.22e-21
C17314 _216_/A _216_/a_27_7# 0.026f
C17315 _306_/X _300_/Y 2.69e-20
C17316 _339_/a_193_7# _195_/a_27_257# 2.26e-20
C17317 _145_/A _146_/C 0.025f
C17318 _175_/Y _298_/X 0.0229f
C17319 _185_/A _229_/a_226_257# 1.66e-19
C17320 _322_/a_1217_7# _321_/Q 2.56e-19
C17321 _297_/A _300_/a_27_257# 2.68e-19
C17322 _306_/S _190_/A 0.506f
C17323 _308_/a_535_334# _308_/X 1.23e-19
C17324 _325_/Q _316_/a_193_7# 8.51e-20
C17325 _339_/Q _337_/D 0.162f
C17326 _339_/D _337_/Q 0.00404f
C17327 _346_/a_1056_7# _346_/Q 6.07e-20
C17328 _145_/A _157_/A 3.78e-19
C17329 _326_/a_1283_n19# _283_/A 0.0028f
C17330 _231_/a_79_n19# _315_/D 0.0443f
C17331 _340_/a_27_7# _336_/a_27_7# 1.42e-21
C17332 _273_/A _306_/S 0.0434f
C17333 _318_/a_761_249# _317_/D 8.13e-20
C17334 _322_/a_639_7# VPWR 7.56e-19
C17335 _330_/Q _331_/D 0.0322f
C17336 _322_/a_651_373# VGND 0.0014f
C17337 _307_/X _286_/Y 0.078f
C17338 _315_/a_27_7# _177_/A 5.32e-20
C17339 _313_/a_1283_n19# _284_/A 0.00331f
C17340 _330_/Q _330_/a_193_7# 0.00348f
C17341 _298_/C _204_/Y 1.9e-20
C17342 _346_/a_1602_7# _165_/X 0.0307f
C17343 rstn _338_/a_1108_7# 5.75e-19
C17344 input3/a_27_7# output41/a_27_7# 5.19e-19
C17345 _162_/X _314_/a_543_7# 2.04e-19
C17346 _250_/a_78_159# _191_/B 0.029f
C17347 _344_/a_1056_7# VPWR 3.31e-19
C17348 _255_/B _295_/a_676_257# 6.49e-19
C17349 clkbuf_2_1_0_clk/A _263_/B 5.66e-20
C17350 _281_/A _327_/Q 1.8e-20
C17351 _329_/a_761_249# _346_/SET_B -0.00742f
C17352 _330_/a_27_7# VPWR 0.0574f
C17353 _227_/a_113_7# VGND -1.06e-19
C17354 _298_/C _298_/a_181_7# 7.87e-19
C17355 _231_/a_512_7# _217_/A 3.35e-19
C17356 _327_/a_1283_n19# _248_/B 5.43e-19
C17357 _318_/Q VPWR 2.23f
C17358 _306_/S _173_/a_556_7# 8.54e-19
C17359 _308_/X _184_/a_76_159# 0.0269f
C17360 _325_/a_27_7# _324_/Q 1.08e-19
C17361 _227_/A _333_/a_639_7# 4.47e-21
C17362 _306_/X VGND 0.894f
C17363 _285_/A _309_/a_1462_7# 1.69e-21
C17364 _326_/a_1108_7# _232_/A 1.16e-20
C17365 clk clkbuf_0_clk/X 3.27e-20
C17366 _263_/B _310_/Q 9.05e-20
C17367 _194_/X _313_/a_193_7# 2.08e-22
C17368 output32/a_27_7# _266_/a_113_257# 3.66e-20
C17369 _320_/Q _321_/a_1283_n19# 5.86e-20
C17370 _319_/Q repeater43/X 0.0237f
C17371 _228_/A _327_/Q 6.16e-19
C17372 _168_/a_397_257# clkbuf_2_3_0_clk/A 3.44e-19
C17373 _286_/B _310_/D 7.04e-21
C17374 _337_/a_27_7# _340_/D 1.88e-21
C17375 _337_/a_1108_7# _194_/X 0.00274f
C17376 _337_/a_761_249# _193_/Y 8.36e-22
C17377 _337_/a_1283_n19# _340_/Q 0.00444f
C17378 _318_/Q _318_/a_543_7# 0.0304f
C17379 _324_/a_193_7# _297_/A 5.06e-20
C17380 _248_/A _327_/D 0.00102f
C17381 _279_/Y rstn 0.521f
C17382 _335_/a_448_7# _335_/D 0.0214f
C17383 _342_/a_1270_373# VGND 6.94e-20
C17384 _342_/a_805_7# VPWR 2.03e-19
C17385 _166_/Y _345_/D 4.6e-20
C17386 _343_/CLK _194_/X 2.62e-19
C17387 _258_/S _265_/B 0.0172f
C17388 _329_/a_1108_7# _331_/CLK 3.83e-20
C17389 _300_/Y _147_/Y 1.22e-22
C17390 _294_/A _273_/A 0.117f
C17391 _196_/A _341_/Q 7.78e-19
C17392 _331_/CLK _327_/D 0.0381f
C17393 _252_/a_27_7# _324_/D 3.71e-20
C17394 _147_/A _336_/D 8.42e-20
C17395 _319_/Q _319_/a_1462_7# 0.00212f
C17396 _322_/a_193_7# result[5] 0.00245f
C17397 clkbuf_2_3_0_clk/A _216_/A 0.00617f
C17398 _339_/D _339_/Q 1.04e-19
C17399 _248_/a_109_257# VGND -9.98e-19
C17400 _255_/X _340_/CLK 3.74e-20
C17401 output16/a_27_7# VGND 0.0626f
C17402 _273_/A _327_/D 0.0233f
C17403 _241_/a_199_7# VPWR -1.99e-19
C17404 _217_/A _223_/a_93_n19# 0.0101f
C17405 _304_/X _223_/a_250_257# 0.00144f
C17406 _312_/a_543_7# _311_/a_27_7# 9.1e-21
C17407 _312_/a_193_7# _311_/a_761_249# 8.57e-22
C17408 _285_/A _344_/a_193_7# 1.81e-20
C17409 clk input1/X 0.00773f
C17410 _306_/S _178_/a_27_7# 8.18e-19
C17411 _340_/a_27_7# _225_/B 2.43e-19
C17412 _340_/a_193_7# _336_/Q 1.58e-20
C17413 _321_/Q _322_/Q 0.0145f
C17414 _341_/a_1283_n19# _315_/a_27_7# 2.95e-20
C17415 _341_/a_761_249# _315_/a_761_249# 4.11e-21
C17416 _341_/a_193_7# _315_/a_543_7# 2.73e-20
C17417 _341_/a_27_7# _315_/a_1283_n19# 3.39e-20
C17418 result[1] _317_/D 3.06e-20
C17419 _255_/a_30_13# _206_/A 6.99e-22
C17420 _283_/A _248_/A 0.282f
C17421 _254_/A _166_/Y 7.19e-19
C17422 _216_/A _327_/Q 0.0509f
C17423 _341_/a_543_7# _298_/A 0.00516f
C17424 _290_/A _288_/Y 3.45e-20
C17425 _345_/a_27_7# _164_/Y 7.4e-20
C17426 _341_/Q _298_/X 7.28e-20
C17427 _212_/X _221_/a_346_7# 0.00286f
C17428 _327_/Q _221_/a_584_7# 1.59e-19
C17429 _344_/a_27_7# _344_/a_652_n19# -0.00438f
C17430 _228_/A _192_/B 1.07e-20
C17431 _233_/a_199_7# VGND -9.65e-20
C17432 _283_/A _331_/CLK 0.00967f
C17433 _320_/a_1462_7# _328_/D 4.94e-20
C17434 _294_/A trim[4] 0.276f
C17435 _346_/a_27_7# _242_/A 3.09e-20
C17436 _321_/D _269_/A 0.29f
C17437 _216_/A _313_/a_1270_373# 2.49e-19
C17438 _256_/a_80_n19# _215_/A 2.9e-19
C17439 _283_/A _190_/A 0.00724f
C17440 _340_/CLK _310_/a_543_7# 1.57e-19
C17441 _277_/Y _286_/a_113_7# 1.81e-19
C17442 _181_/X _227_/A 0.195f
C17443 _309_/a_1108_7# _172_/B 5.13e-20
C17444 output8/a_27_7# output5/a_27_7# 0.0128f
C17445 cal _202_/a_93_n19# 1.53e-20
C17446 _147_/Y VGND 3.03f
C17447 _230_/a_27_7# _316_/D 1.51e-20
C17448 _339_/a_761_249# _193_/Y 0.00834f
C17449 _339_/a_543_7# _306_/S 0.012f
C17450 _339_/a_27_7# _340_/D 0.0145f
C17451 _339_/a_1108_7# _194_/X 0.0119f
C17452 _298_/B _333_/D 0.00279f
C17453 _298_/C _225_/B 0.00815f
C17454 _312_/a_651_373# VPWR 0.00825f
C17455 _312_/a_1108_7# VGND 0.015f
C17456 rstn _334_/a_1283_n19# 8.16e-19
C17457 _273_/A _283_/A 0.00744f
C17458 _297_/A _160_/X 3.08e-21
C17459 _299_/X _299_/a_292_257# 0.00119f
C17460 _347_/Q _299_/a_78_159# 7.7e-20
C17461 _344_/a_193_7# _172_/A 2.28e-19
C17462 output40/a_27_7# VPWR 0.0949f
C17463 output32/a_27_7# VPWR 0.0743f
C17464 _264_/a_199_7# _340_/CLK 1.5e-19
C17465 _179_/a_27_7# _153_/B 3.43e-21
C17466 _248_/B _248_/A 0.0656f
C17467 _346_/a_476_7# _301_/a_240_7# 3.53e-21
C17468 _162_/X _315_/D 0.0152f
C17469 _316_/a_543_7# _315_/a_761_249# 7.57e-19
C17470 _316_/a_1283_n19# _315_/a_193_7# 4.2e-19
C17471 _304_/a_288_7# _227_/A 5.69e-19
C17472 _340_/a_1283_n19# _336_/a_651_373# 2.2e-21
C17473 _272_/a_39_257# _223_/a_250_257# 0.00117f
C17474 _326_/a_27_7# _326_/Q 0.00778f
C17475 clk _286_/Y 0.0956f
C17476 _338_/Q _297_/Y 0.012f
C17477 _164_/A _160_/X 0.0241f
C17478 cal _197_/a_27_7# 0.0208f
C17479 _325_/a_448_7# _286_/Y 0.00675f
C17480 _330_/Q _330_/a_1462_7# 5.05e-19
C17481 clkbuf_2_1_0_clk/A _194_/A 4.44e-19
C17482 _316_/D _232_/A 0.0973f
C17483 _331_/CLK _248_/B 3.74e-19
C17484 _324_/Q _146_/C 0.00252f
C17485 _345_/a_193_7# _286_/B 7.88e-20
C17486 _216_/A _192_/B 0.00109f
C17487 _250_/X _191_/B 0.0802f
C17488 _304_/S _328_/Q 4.32e-20
C17489 _321_/a_193_7# _248_/A 1.78e-20
C17490 _271_/A _333_/a_193_7# 1.23e-21
C17491 _188_/a_218_7# _255_/B 6.3e-19
C17492 clkbuf_2_1_0_clk/A _338_/a_193_7# 9.91e-21
C17493 clkbuf_2_0_0_clk/a_75_172# _338_/a_1108_7# 5.46e-19
C17494 _304_/a_79_n19# _304_/X 0.00747f
C17495 _330_/a_1217_7# VPWR 8.33e-21
C17496 _330_/a_639_7# VGND 5.32e-19
C17497 _344_/a_1032_373# _171_/a_78_159# 4.96e-19
C17498 _157_/A _324_/Q 0.0551f
C17499 _258_/S clkbuf_2_1_0_clk/A 0.00631f
C17500 _227_/A _343_/Q 3.44e-19
C17501 _273_/A _248_/B 0.0956f
C17502 output21/a_27_7# _330_/Q 0.0023f
C17503 _337_/a_543_7# _283_/A 1.88e-19
C17504 _321_/a_27_7# _316_/D 1.12e-21
C17505 _321_/a_193_7# _331_/CLK 0.587f
C17506 _338_/Q _310_/a_193_7# 9.31e-20
C17507 clk _250_/a_215_7# 2.44e-20
C17508 _308_/X _188_/S 0.115f
C17509 _346_/SET_B _310_/a_1283_n19# -7.41e-19
C17510 _346_/SET_B _319_/D 0.0627f
C17511 _325_/a_27_7# _216_/A 3.17e-19
C17512 _333_/a_1108_7# VGND -0.00654f
C17513 _333_/a_651_373# VPWR -0.0085f
C17514 _242_/A _319_/a_27_7# 0.00671f
C17515 _341_/a_448_7# _341_/Q 1.16e-22
C17516 _258_/S _310_/Q 0.0278f
C17517 _315_/Q _315_/a_193_7# 0.00298f
C17518 output22/a_27_7# _315_/a_1108_7# 2.72e-19
C17519 _343_/a_193_7# _176_/a_27_7# 6.56e-20
C17520 _254_/Y _190_/A 0.0211f
C17521 _331_/Q _246_/B 0.0135f
C17522 _198_/a_93_n19# _198_/a_256_7# -6.6e-20
C17523 _336_/a_193_7# _340_/CLK 8.38e-19
C17524 output31/a_27_7# _346_/SET_B 1.94e-19
C17525 _153_/a_109_53# _332_/Q 0.0323f
C17526 _223_/a_250_257# VGND 0.00251f
C17527 _223_/a_346_7# VPWR -9.64e-19
C17528 _301_/X _286_/Y 1.61e-20
C17529 _324_/a_193_7# _325_/D 0.00389f
C17530 repeater43/X _255_/B 1.25e-19
C17531 _304_/S _269_/A 1.56e-20
C17532 _320_/Q clkbuf_2_1_0_clk/A 0.0474f
C17533 _314_/a_1283_n19# _347_/a_448_7# 2.28e-19
C17534 _296_/Y _306_/S 0.0527f
C17535 _325_/a_651_373# _284_/A 1.1e-20
C17536 _283_/A _178_/a_27_7# 0.0131f
C17537 _344_/a_1182_221# _161_/Y 0.00439f
C17538 repeater43/a_27_7# rstn 0.00706f
C17539 input4/X input4/a_27_7# 0.00293f
C17540 _346_/D _347_/a_27_7# 4.25e-21
C17541 _311_/D _254_/B 0.00186f
C17542 _275_/A _242_/A 0.565f
C17543 _339_/D _336_/D 7.14e-21
C17544 _323_/a_448_7# _323_/D 0.00455f
C17545 _345_/D _297_/Y 3.09e-20
C17546 _342_/Q _207_/C 4.53e-21
C17547 _192_/a_150_257# VPWR 3.79e-19
C17548 _309_/a_193_7# _164_/A 0.00164f
C17549 _345_/a_1056_7# _164_/A 1.33e-19
C17550 _202_/a_93_n19# _284_/A 0.0113f
C17551 _319_/Q result[6] 0.0017f
C17552 _330_/D _330_/a_1108_7# 8.65e-22
C17553 _329_/a_448_7# _212_/X 2.2e-20
C17554 _329_/a_1108_7# _217_/X 0.00204f
C17555 _329_/a_651_373# _327_/Q 9.23e-20
C17556 _217_/X _327_/D 0.00674f
C17557 _146_/C _228_/A 0.326f
C17558 _209_/a_27_257# _332_/Q 0.0131f
C17559 _328_/a_27_7# clkbuf_2_1_0_clk/A 2.11e-20
C17560 _225_/a_145_35# _190_/A 6.69e-19
C17561 _339_/a_543_7# _283_/A 0.0355f
C17562 _200_/a_584_7# clkbuf_2_1_0_clk/A 3.41e-19
C17563 output30/a_27_7# sample 0.00317f
C17564 _346_/SET_B _336_/a_761_249# 0.0068f
C17565 ctln[6] clk 8.04e-20
C17566 _281_/Y clkbuf_0_clk/X 0.144f
C17567 _290_/Y trimb[2] 0.0193f
C17568 _283_/Y _197_/X 4.53e-21
C17569 _236_/B _243_/a_113_257# 1.23e-19
C17570 _275_/Y _312_/a_639_7# 0.00121f
C17571 _259_/a_113_257# VPWR 0.0513f
C17572 _316_/D _243_/a_199_7# 1.91e-19
C17573 _260_/B _215_/A 0.00971f
C17574 _286_/B VPWR 2.62f
C17575 _290_/A _337_/Q 0.00759f
C17576 _199_/a_256_7# _340_/CLK 6.26e-20
C17577 cal _284_/A 0.0259f
C17578 _157_/A _228_/A 0.69f
C17579 _345_/a_27_7# _165_/a_78_159# 8.39e-19
C17580 _185_/A _226_/X 0.323f
C17581 _315_/a_27_7# _248_/A 0.00737f
C17582 _254_/A _297_/Y 0.0486f
C17583 _181_/X _297_/B 1.62e-19
C17584 _300_/Y _347_/a_193_7# 0.00991f
C17585 _347_/Q _347_/a_1108_7# 0.00191f
C17586 _258_/a_218_7# _306_/X 4.61e-19
C17587 _258_/a_439_7# _313_/Q -4.44e-34
C17588 _255_/B _191_/B 0.00971f
C17589 _286_/a_113_7# VGND 1.93e-19
C17590 _304_/a_79_n19# VGND 0.0252f
C17591 _331_/CLK _315_/a_27_7# 4.53e-21
C17592 _304_/a_306_329# VPWR -0.00273f
C17593 _324_/a_543_7# _216_/X 0.00135f
C17594 _326_/a_1217_7# _326_/Q 4.66e-20
C17595 _332_/D _225_/B 2.61e-20
C17596 _256_/a_80_n19# VGND 0.036f
C17597 _279_/Y _324_/a_27_7# 3.03e-19
C17598 _256_/a_209_7# VPWR -3.74e-19
C17599 _329_/D clkbuf_0_clk/X 0.0102f
C17600 _283_/A _217_/X 0.131f
C17601 _309_/a_27_7# _286_/B 7.48e-19
C17602 _227_/A _204_/a_27_7# 3.1e-19
C17603 input4/X _204_/Y 4.3e-20
C17604 _227_/A _208_/a_215_7# 1.57e-19
C17605 _291_/a_39_257# _346_/SET_B 1.43e-19
C17606 _279_/Y _314_/a_651_373# 0.00488f
C17607 _342_/Q _150_/C 0.063f
C17608 _317_/Q _212_/X 3e-21
C17609 _281_/Y input1/X 0.00636f
C17610 repeater43/X _325_/Q 0.00628f
C17611 _216_/X _217_/A 0.0133f
C17612 _315_/D _298_/C 1.8e-20
C17613 _346_/a_652_n19# _170_/a_76_159# 2.42e-21
C17614 _144_/a_27_7# _150_/C 7.8e-19
C17615 ctlp[1] _321_/Q 6.98e-19
C17616 _326_/a_1283_n19# _242_/B 1.35e-20
C17617 _344_/a_1032_373# _172_/B 5.45e-19
C17618 _176_/a_27_7# VGND 0.0536f
C17619 _157_/A _216_/A 0.00594f
C17620 repeater43/X _298_/a_27_7# 5.62e-20
C17621 _144_/A _232_/A 6.36e-20
C17622 _338_/D _199_/a_584_7# 2.44e-19
C17623 _338_/Q _199_/a_93_n19# 0.0118f
C17624 _320_/a_27_7# ctlp[4] 4.07e-19
C17625 _210_/a_109_257# _225_/X 5.43e-19
C17626 _283_/Y _312_/a_193_7# 6.46e-20
C17627 _242_/A _319_/a_1217_7# 1.61e-19
C17628 _157_/A _251_/a_510_7# 0.00245f
C17629 _324_/Q _251_/a_79_n19# 0.0581f
C17630 _267_/B clkc 1.38e-19
C17631 _207_/C _204_/Y 0.383f
C17632 _341_/D _341_/Q 0.0753f
C17633 _327_/a_761_249# _217_/A 2.17e-20
C17634 _327_/a_543_7# _304_/X 3.38e-20
C17635 _315_/Q _315_/a_1462_7# 4.85e-19
C17636 _260_/A _228_/A 7.34e-20
C17637 _343_/a_1270_373# _343_/Q 4.51e-20
C17638 _346_/a_652_n19# clkbuf_2_1_0_clk/A 8.1e-20
C17639 _332_/a_761_249# VPWR 0.0168f
C17640 _332_/a_27_7# VGND 0.0459f
C17641 rstn _339_/a_1283_n19# 1.95e-20
C17642 _343_/CLK _175_/Y 1.34e-20
C17643 _248_/B _217_/X 0.00655f
C17644 _320_/Q _278_/a_68_257# 0.00651f
C17645 _347_/a_193_7# VGND 0.0148f
C17646 _347_/a_543_7# VPWR 0.00821f
C17647 _290_/A _339_/Q 0.0186f
C17648 _326_/a_543_7# _304_/X 0.00692f
C17649 _326_/a_761_249# _217_/A 4.81e-19
C17650 _325_/a_543_7# _296_/a_213_83# 3.39e-21
C17651 _153_/A _332_/Q 0.492f
C17652 ctlp[7] VPWR 0.0464f
C17653 _338_/Q _336_/Q 6.79e-20
C17654 _323_/D _244_/B 1.61e-20
C17655 repeater43/X _321_/a_1108_7# -0.0198f
C17656 _292_/A _160_/X 0.0117f
C17657 _336_/a_193_7# _313_/a_543_7# 2.54e-20
C17658 _336_/a_1283_n19# _313_/a_27_7# 4.16e-21
C17659 _250_/a_493_257# _284_/A 1.19e-20
C17660 _267_/A _344_/D 3.63e-20
C17661 _314_/Q _347_/a_27_7# 0.0106f
C17662 _297_/B _347_/a_1108_7# 0.0576f
C17663 _314_/a_1283_n19# _347_/D 0.00609f
C17664 _254_/A _242_/A 8.1e-20
C17665 _309_/D _310_/a_193_7# 4.59e-19
C17666 _232_/X _241_/a_113_257# 7.45e-19
C17667 _163_/a_215_7# _310_/D 6.51e-21
C17668 _267_/B _310_/a_543_7# 0.0018f
C17669 _306_/a_76_159# _286_/B 0.0116f
C17670 _258_/S _311_/a_27_7# 0.0113f
C17671 _281_/Y _286_/Y 0.0288f
C17672 _160_/X _160_/A 0.374f
C17673 _346_/Q _267_/A 2.48e-20
C17674 repeater43/X _153_/a_297_257# 5.63e-19
C17675 _313_/Q _254_/B 0.0011f
C17676 _312_/Q _311_/a_1283_n19# 0.00684f
C17677 _327_/a_27_7# _279_/A 1.31e-21
C17678 repeater42/a_27_7# _325_/D 2.06e-20
C17679 _328_/a_27_7# _278_/a_68_257# 2.81e-21
C17680 _166_/Y _286_/Y 0.0606f
C17681 _168_/a_481_7# _267_/A 8.28e-20
C17682 _216_/A _260_/A 0.729f
C17683 clk _269_/A 0.0532f
C17684 _341_/a_1108_7# VPWR -0.00292f
C17685 _341_/a_543_7# VGND -0.00279f
C17686 _296_/Y _248_/B 3.63e-20
C17687 _216_/X _220_/a_250_257# 4.6e-19
C17688 _145_/A _232_/A 0.00175f
C17689 _327_/a_193_7# _218_/a_93_n19# 0.00158f
C17690 _327_/a_27_7# _218_/a_250_257# 6.8e-20
C17691 _338_/a_543_7# VGND 0.00153f
C17692 _338_/a_1108_7# VPWR 0.0106f
C17693 _184_/a_505_n19# _286_/B 2e-21
C17694 _227_/A _346_/SET_B 1.11e-19
C17695 ctlp[0] VGND 0.12f
C17696 _281_/Y _250_/a_215_7# 0.00464f
C17697 output9/a_27_7# output34/a_27_7# 5.88e-21
C17698 _346_/a_1182_221# _277_/Y 4.22e-21
C17699 _329_/a_193_7# _280_/a_68_257# 1.64e-20
C17700 _320_/Q _220_/a_256_7# 9.29e-19
C17701 _329_/Q _220_/a_250_257# 0.0256f
C17702 _341_/Q _143_/a_27_7# 0.00272f
C17703 _308_/a_76_159# _298_/C 0.00293f
C17704 clkbuf_2_1_0_clk/A _319_/a_761_249# 7.74e-22
C17705 _346_/SET_B _314_/a_1108_7# 0.00587f
C17706 clkbuf_2_1_0_clk/A _337_/a_27_7# 3.61e-22
C17707 _248_/A _242_/B 0.577f
C17708 output25/a_27_7# result[3] 0.0104f
C17709 _343_/D clk 0.00132f
C17710 _271_/A _316_/a_27_7# 2.07e-19
C17711 _342_/a_639_7# _323_/D 5.63e-20
C17712 _285_/A _164_/A 9.41e-21
C17713 _319_/Q result[4] 0.00665f
C17714 _317_/Q _317_/a_448_7# 2.15e-19
C17715 _336_/a_761_249# _147_/A 3.98e-19
C17716 _242_/A _317_/a_761_249# 9.61e-19
C17717 _251_/a_79_n19# _228_/A 0.0324f
C17718 clkbuf_0_clk/a_110_7# _248_/B 3.1e-21
C17719 _337_/Q _310_/a_27_7# 0.0625f
C17720 _340_/a_651_373# VPWR 0.00255f
C17721 _340_/a_1108_7# VGND -0.00735f
C17722 _236_/a_109_257# _318_/D 0.0032f
C17723 _331_/CLK _242_/B 0.00782f
C17724 _260_/a_27_257# _147_/A 0.00101f
C17725 _325_/Q _317_/a_543_7# 4.5e-19
C17726 _184_/a_76_159# _298_/X 8.95e-20
C17727 _279_/Y VPWR 1.88f
C17728 _316_/a_1283_n19# VGND -0.00529f
C17729 _316_/a_448_7# VPWR 0.0022f
C17730 _327_/a_448_7# _330_/Q 8.97e-19
C17731 repeater43/X _326_/Q 0.258f
C17732 _343_/a_27_7# _248_/A 0.00813f
C17733 _324_/a_193_7# _331_/CLK 2.36e-20
C17734 _344_/a_193_7# _164_/A 0.00945f
C17735 _169_/Y _345_/Q 1.49e-19
C17736 _260_/B VGND 0.31f
C17737 _258_/S _309_/a_1283_n19# 1.58e-20
C17738 _328_/a_193_7# _220_/a_250_257# 1.26e-19
C17739 _172_/A _297_/A 3.97e-20
C17740 _208_/a_292_257# VPWR -7.48e-19
C17741 trim[4] _284_/a_39_257# 0.00777f
C17742 _242_/A _331_/a_1108_7# 3.82e-21
C17743 _255_/X clk 0.0114f
C17744 _309_/a_193_7# _292_/A 9.64e-20
C17745 _313_/a_1108_7# _336_/Q 1.12e-19
C17746 _327_/a_1108_7# VPWR 0.018f
C17747 _327_/a_543_7# VGND -0.00132f
C17748 _325_/a_639_7# _255_/B 1.66e-20
C17749 _182_/a_79_n19# _154_/a_27_7# 2.07e-21
C17750 _342_/a_193_7# _342_/D 0.0196f
C17751 _346_/a_476_7# _346_/D 0.0336f
C17752 _273_/A _324_/a_193_7# 0.00176f
C17753 _341_/Q _343_/CLK 3.03e-20
C17754 _297_/A _232_/X 8.3e-19
C17755 repeater43/X _315_/a_1283_n19# -8.73e-19
C17756 _273_/A _262_/a_113_257# 0.0101f
C17757 _172_/A _164_/A 1.19e-19
C17758 _195_/a_27_257# _340_/Q 0.0144f
C17759 _322_/a_1108_7# _322_/Q 0.00224f
C17760 _326_/a_1108_7# VPWR -4.48e-19
C17761 _326_/a_543_7# VGND 0.0209f
C17762 _185_/A input1/X 0.0526f
C17763 _234_/B _317_/a_1283_n19# 1.85e-20
C17764 _277_/Y _319_/a_1283_n19# 1.01e-20
C17765 _345_/a_1182_221# _163_/a_78_159# 3.22e-19
C17766 _324_/Q _251_/X 0.00205f
C17767 _251_/a_79_n19# _216_/A 0.00615f
C17768 _281_/Y ctln[6] 0.0375f
C17769 _254_/A _336_/Q 0.00143f
C17770 _347_/Q _346_/SET_B 0.485f
C17771 _315_/Q VGND 1.22f
C17772 _324_/Q _296_/a_213_83# 0.00672f
C17773 result[0] VPWR 0.222f
C17774 _332_/a_1217_7# VGND 9.98e-20
C17775 _328_/a_1283_n19# VPWR 0.0236f
C17776 _328_/a_761_249# VGND -0.00137f
C17777 _347_/a_1462_7# VGND 2.42e-19
C17778 repeater43/X _224_/a_256_7# 5.78e-20
C17779 _298_/B _178_/a_27_7# 5.76e-19
C17780 _341_/Q _178_/a_193_257# 2.85e-19
C17781 _227_/A _206_/A 0.96f
C17782 _344_/a_27_7# _286_/B 1.56e-19
C17783 _191_/B _209_/a_109_7# 1.96e-19
C17784 _342_/Q cal 0.00122f
C17785 _328_/a_448_7# _297_/B 5.27e-20
C17786 _321_/a_1283_n19# result[7] 5.9e-19
C17787 _164_/Y _171_/a_493_257# 6.82e-19
C17788 _257_/a_222_53# input1/X 1.18e-19
C17789 _273_/A _266_/a_199_7# 3.99e-19
C17790 _339_/Q _310_/a_27_7# 0.00883f
C17791 _324_/a_543_7# _216_/a_27_7# 0.00527f
C17792 _258_/a_218_334# _286_/B 8.46e-19
C17793 _258_/a_505_n19# _196_/A 1.16e-21
C17794 _346_/a_1032_373# _160_/X 0.00133f
C17795 _346_/a_956_373# _299_/X 7.27e-19
C17796 _167_/X _344_/D 2.27e-20
C17797 _334_/a_761_249# VGND 0.00201f
C17798 _334_/a_1283_n19# VPWR 0.0372f
C17799 _227_/A _334_/D 1.85e-19
C17800 repeater43/X _154_/A 0.00156f
C17801 _333_/a_1283_n19# _254_/B 1.34e-20
C17802 _163_/a_493_257# _160_/X 7.5e-19
C17803 _331_/CLK _245_/a_199_7# 6.79e-20
C17804 _316_/D _245_/a_113_257# 1.27e-19
C17805 _186_/a_297_7# _182_/X 1.73e-20
C17806 _307_/a_218_7# _227_/A 1.22e-19
C17807 _323_/a_1283_n19# _298_/X 4.95e-21
C17808 _167_/X _346_/Q 0.0208f
C17809 _342_/Q _150_/a_193_257# 9.42e-19
C17810 _309_/D _336_/Q 0.00105f
C17811 _216_/a_27_7# _217_/A 4.02e-19
C17812 _216_/A _340_/Q 1.71e-20
C17813 input1/X _310_/a_193_7# 1.52e-20
C17814 clkbuf_0_clk/X _242_/A 0.0918f
C17815 _273_/A _160_/X 0.336f
C17816 _323_/a_651_373# _176_/a_27_7# 1.34e-19
C17817 _323_/a_193_7# _298_/C 6.33e-21
C17818 _323_/a_543_7# _343_/Q 5.46e-19
C17819 _188_/S _196_/A 0.149f
C17820 _314_/a_1108_7# _156_/a_39_257# 0.00178f
C17821 _168_/a_481_7# _167_/X 0.00176f
C17822 _168_/a_397_257# _165_/X 0.00584f
C17823 input3/a_27_7# _192_/B 9.56e-21
C17824 _172_/A _304_/a_257_159# 4.41e-21
C17825 _274_/a_121_257# VGND -3.46e-19
C17826 _316_/Q _316_/a_639_7# 0.00497f
C17827 _329_/a_1283_n19# _281_/A 8.8e-19
C17828 _320_/Q _328_/D 0.0278f
C17829 _308_/S _298_/C 0.00144f
C17830 _325_/a_639_7# _325_/Q 2.06e-20
C17831 _281_/Y _328_/Q 0.00118f
C17832 _329_/a_193_7# _281_/Y 0.0143f
C17833 _328_/a_805_7# _279_/A 4.57e-19
C17834 _346_/SET_B _297_/B 1.75f
C17835 _172_/A _177_/A 0.00101f
C17836 _254_/A _170_/a_489_373# 7.53e-20
C17837 _342_/a_761_249# _177_/a_27_7# 0.00223f
C17838 _227_/A _147_/A 0.00637f
C17839 _236_/B _330_/Q 0.014f
C17840 _334_/Q _154_/A 8.28e-19
C17841 _293_/a_39_257# _194_/A 0.00142f
C17842 _342_/a_27_7# output41/a_27_7# 7.48e-21
C17843 _324_/Q _232_/A 0.505f
C17844 _319_/a_193_7# _279_/A 1.84e-20
C17845 _251_/X _228_/A 0.0299f
C17846 _295_/a_512_7# VGND 0.0502f
C17847 _294_/Y _265_/a_109_257# 0.00131f
C17848 _346_/a_1182_221# VGND 0.0058f
C17849 _346_/a_1602_7# VPWR 0.00609f
C17850 _297_/a_27_257# _297_/Y 0.0256f
C17851 _337_/Q _310_/a_1217_7# 3.64e-20
C17852 comp _344_/Q 8.78e-20
C17853 _160_/X _173_/a_556_7# 5.06e-19
C17854 _149_/a_27_7# _298_/A 8.35e-19
C17855 _333_/a_27_7# _333_/a_193_7# -0.333f
C17856 _335_/a_543_7# _204_/a_27_7# 8.04e-21
C17857 _335_/a_1283_n19# _204_/a_27_257# 1.62e-20
C17858 _227_/A _149_/A 2.2e-19
C17859 _165_/X _216_/A 2.4e-20
C17860 _163_/a_292_257# VGND -0.00122f
C17861 _163_/a_215_7# VPWR -5.14e-20
C17862 _329_/a_761_249# _319_/Q 0.0192f
C17863 _316_/D VPWR 0.834f
C17864 _318_/a_1283_n19# _248_/A 5.81e-20
C17865 _172_/A _333_/D 1.05e-21
C17866 _347_/Q _313_/a_761_249# 7e-20
C17867 _293_/a_39_257# _258_/S 2.96e-19
C17868 _346_/a_476_7# _314_/Q 5e-21
C17869 _340_/CLK _311_/a_1283_n19# 1.27e-20
C17870 _333_/Q VGND 0.875f
C17871 _328_/a_27_7# _328_/D 0.0475f
C17872 _326_/D _330_/Q 4.26e-20
C17873 cal _204_/Y 1.23e-19
C17874 _191_/B _154_/A 0.0151f
C17875 _192_/B _153_/A 0.00305f
C17876 _329_/a_193_7# _329_/D 0.513f
C17877 _329_/D _328_/Q 3.92e-21
C17878 repeater42/a_27_7# _248_/A 2.21e-20
C17879 repeater43/X _235_/a_199_7# 7.04e-21
C17880 _321_/D _318_/a_27_7# 0.0135f
C17881 _318_/a_1283_n19# _331_/CLK 1.08e-19
C17882 _336_/a_27_7# _202_/a_93_n19# 1.88e-19
C17883 _335_/D _333_/D 1.39e-20
C17884 _342_/a_1462_7# _342_/D 0.00187f
C17885 output12/a_27_7# _283_/A 0.0224f
C17886 output33/a_27_7# output5/a_27_7# 0.0123f
C17887 _219_/a_250_257# _319_/D 5.46e-20
C17888 _306_/S _193_/Y 0.584f
C17889 _194_/X _340_/D 0.00204f
C17890 cal _298_/a_181_7# 3.53e-19
C17891 _277_/A _276_/a_68_257# 0.0239f
C17892 repeater42/a_27_7# _331_/CLK 0.0664f
C17893 repeater43/a_27_7# VPWR 0.225f
C17894 repeater43/X _324_/a_1108_7# -0.0197f
C17895 _242_/B _217_/X 0.00148f
C17896 _305_/a_505_n19# _305_/X 1.87e-19
C17897 _305_/a_76_159# _194_/A 0.0401f
C17898 cal _336_/a_27_7# 5.07e-21
C17899 _345_/a_1032_373# _158_/Y 0.0128f
C17900 _251_/X _216_/A 0.00259f
C17901 _222_/a_250_257# VPWR 0.0202f
C17902 _285_/A _292_/A 0.0361f
C17903 _232_/X _325_/D 4.51e-20
C17904 _324_/a_543_7# _327_/Q 7.59e-19
C17905 _342_/Q _284_/A 0.638f
C17906 _343_/a_1283_n19# repeater43/X 4.72e-19
C17907 repeater42/a_27_7# _273_/A 4.16e-19
C17908 _331_/Q _330_/a_448_7# 6.16e-20
C17909 _173_/a_226_257# VGND -5.12e-19
C17910 clkbuf_2_3_0_clk/A _346_/D 5.85e-21
C17911 repeater43/X _324_/D 0.299f
C17912 _309_/a_193_7# _273_/A 2.67e-20
C17913 _177_/A _244_/B 0.375f
C17914 _285_/A _160_/A 0.00806f
C17915 _271_/A _334_/a_639_7# 2.23e-19
C17916 _175_/Y output30/a_27_7# 4.04e-19
C17917 _313_/a_27_7# VPWR 0.025f
C17918 _319_/a_448_7# VPWR 0.00443f
C17919 _319_/a_1283_n19# VGND 0.0131f
C17920 _323_/a_761_249# _229_/a_226_7# 3.06e-21
C17921 _323_/a_543_7# _229_/a_76_159# 3.34e-21
C17922 _338_/Q _311_/a_761_249# 5.07e-21
C17923 _346_/SET_B _311_/a_1108_7# 0.0102f
C17924 _344_/a_193_7# _292_/A 2e-19
C17925 _337_/a_1283_n19# VPWR 0.0126f
C17926 _337_/a_761_249# VGND -0.00214f
C17927 _217_/A _327_/Q 0.851f
C17928 _304_/X _212_/X 0.472f
C17929 _301_/a_51_257# _344_/D 1.03e-19
C17930 _347_/Q _147_/A 0.00535f
C17931 _231_/a_676_257# _162_/X 6.33e-19
C17932 _183_/a_553_257# _341_/Q 2.76e-20
C17933 _242_/A _286_/Y 1.95e-19
C17934 _342_/a_761_249# _341_/a_27_7# 2.14e-21
C17935 _342_/a_27_7# _341_/a_761_249# 1.1e-21
C17936 _342_/a_193_7# _341_/a_193_7# 1.91e-20
C17937 _297_/B _313_/a_761_249# 3.21e-20
C17938 _313_/Q _196_/A 4.12e-20
C17939 _306_/X _286_/B 0.0654f
C17940 _320_/Q _322_/a_27_7# 0.0211f
C17941 _344_/a_193_7# _160_/A 4.62e-20
C17942 _232_/A _228_/A 2.68e-20
C17943 _343_/CLK _269_/Y 0.025f
C17944 _346_/Q _301_/a_51_257# 8.6e-19
C17945 output8/a_27_7# VGND 0.0721f
C17946 _167_/a_373_7# _166_/Y 0.00212f
C17947 _289_/a_39_257# _287_/a_39_257# 3.42e-20
C17948 _341_/D _184_/a_76_159# 2.04e-21
C17949 _320_/Q _320_/a_651_373# 3.49e-19
C17950 _238_/B _320_/a_1283_n19# 6.05e-19
C17951 _307_/a_76_159# VGND 0.00845f
C17952 _307_/a_218_334# VPWR 1.19e-19
C17953 _292_/A _172_/A 4.7e-20
C17954 _281_/Y _255_/X 0.507f
C17955 _345_/a_381_7# _345_/D 0.021f
C17956 _345_/a_562_373# _345_/Q 1.94e-19
C17957 _254_/a_109_257# VPWR 2.54e-19
C17958 _294_/A _193_/Y 0.00273f
C17959 output17/a_27_7# ctlp[3] 0.0152f
C17960 _275_/Y _346_/SET_B 0.338f
C17961 rstn _195_/a_27_257# 0.0576f
C17962 _343_/a_639_7# _343_/CLK 4.94e-20
C17963 _325_/a_639_7# _326_/Q 3.7e-19
C17964 _309_/a_193_7# trim[4] 7.44e-20
C17965 _172_/A _160_/A 6.14e-20
C17966 cal _199_/a_250_257# 6.01e-20
C17967 input1/X _199_/a_93_n19# 0.00759f
C17968 _178_/a_109_257# VPWR -0.00125f
C17969 _340_/a_27_7# _197_/X 0.00982f
C17970 _329_/a_1462_7# _281_/Y 4.06e-19
C17971 _315_/D _150_/C 0.111f
C17972 _340_/a_651_373# _198_/a_93_n19# 4.61e-20
C17973 _226_/a_297_7# VGND 0.047f
C17974 _272_/a_39_257# _212_/X 9.42e-20
C17975 _279_/Y _211_/a_27_257# 0.00103f
C17976 _325_/a_1108_7# _227_/A 1.4e-19
C17977 _216_/A _232_/A 0.00157f
C17978 cal _225_/B 0.237f
C17979 _325_/a_27_7# _324_/a_543_7# 1.97e-19
C17980 input1/X _336_/Q 0.0727f
C17981 _174_/a_27_257# _310_/D 1.9e-19
C17982 _294_/Y _165_/X 1.01e-20
C17983 _346_/a_1296_7# VGND 4.49e-19
C17984 _255_/a_30_13# _255_/B 0.0137f
C17985 rstn _207_/a_181_7# 7.76e-19
C17986 _238_/B _232_/X 0.00191f
C17987 _297_/B _147_/A 0.459f
C17988 clkbuf_0_clk/X _314_/a_761_249# 1.37e-19
C17989 _309_/a_639_7# _346_/SET_B -2.04e-20
C17990 _335_/D _208_/a_78_159# 8.16e-19
C17991 _335_/a_639_7# _207_/X 6.67e-19
C17992 _197_/a_27_7# _225_/B 0.00306f
C17993 _343_/a_1108_7# _226_/X 2.19e-19
C17994 _212_/X _220_/a_93_n19# 0.0096f
C17995 _341_/a_1283_n19# _244_/B 0.0103f
C17996 _341_/a_761_249# _317_/D 0.00684f
C17997 _339_/a_761_249# VGND -0.00335f
C17998 _339_/a_1283_n19# VPWR 0.0152f
C17999 _327_/a_1283_n19# _232_/X 0.0143f
C18000 _308_/a_76_159# _207_/C 3.27e-20
C18001 _282_/a_121_257# VGND 2.61e-20
C18002 _319_/Q _319_/D 0.0741f
C18003 _325_/a_27_7# _217_/A 0.0462f
C18004 _325_/a_193_7# _304_/X 0.0257f
C18005 _294_/A output5/a_27_7# 3.1e-19
C18006 _343_/a_1270_373# _149_/A 4.43e-20
C18007 _283_/A _193_/Y 0.0063f
C18008 _326_/a_1283_n19# _232_/X 0.00424f
C18009 _286_/B _147_/Y 0.0852f
C18010 input4/X _335_/a_193_7# 5.66e-19
C18011 _336_/a_27_7# _284_/A 0.0132f
C18012 _330_/Q _331_/a_193_7# 0.02f
C18013 _330_/Q output29/a_27_7# 6.46e-19
C18014 _265_/B _267_/A 0.0271f
C18015 _144_/A VPWR 0.578f
C18016 _318_/a_27_7# _317_/a_27_7# 4.08e-21
C18017 _255_/B _296_/a_493_257# 2.89e-19
C18018 _312_/a_761_249# _312_/Q 0.00238f
C18019 _312_/a_448_7# _312_/D 0.00422f
C18020 cal en 0.0615f
C18021 _317_/a_1108_7# _217_/A 1.5e-20
C18022 _331_/a_27_7# VPWR 0.0769f
C18023 _200_/a_250_257# _197_/X 0.00116f
C18024 _328_/a_543_7# _232_/X 0.00192f
C18025 _320_/a_193_7# _346_/SET_B 0.0135f
C18026 _185_/A _269_/A 6e-19
C18027 _340_/a_1283_n19# _254_/B 6.54e-21
C18028 _212_/X VGND 2.41f
C18029 _335_/a_193_7# _207_/C 8.46e-21
C18030 _335_/a_543_7# _206_/A 4.33e-19
C18031 repeater43/X _318_/a_1270_373# -3.58e-20
C18032 _316_/a_543_7# _317_/D 0.012f
C18033 _290_/A _310_/a_1283_n19# 0.00788f
C18034 _240_/B _242_/A 0.157f
C18035 _313_/a_639_7# VGND -0.00137f
C18036 _313_/a_1217_7# VPWR 3.82e-20
C18037 _323_/a_448_7# _248_/A 6.79e-20
C18038 _258_/a_76_159# _346_/SET_B 0.0187f
C18039 _328_/a_761_249# ctlp[5] 2.49e-21
C18040 _335_/a_543_7# _334_/D 8.71e-19
C18041 _335_/a_1283_n19# _343_/CLK 0.0139f
C18042 _321_/D result[5] 2.63e-19
C18043 _185_/A _343_/D 0.0239f
C18044 _308_/a_76_159# _150_/C 7.6e-20
C18045 output15/a_27_7# _322_/Q 0.024f
C18046 output31/a_27_7# _290_/A 7.71e-21
C18047 repeater42/a_27_7# _217_/X 0.0712f
C18048 _286_/B _333_/a_1108_7# 2.81e-21
C18049 _250_/a_215_7# _336_/Q 2.37e-19
C18050 _250_/a_493_257# _225_/B 6.94e-21
C18051 _216_/X _331_/D 1.69e-19
C18052 _217_/a_27_7# VPWR 0.127f
C18053 _341_/D _188_/S 6.92e-19
C18054 _344_/a_27_7# _163_/a_215_7# 7.36e-20
C18055 _254_/Y _193_/Y 8.25e-20
C18056 _285_/A _273_/A 0.292f
C18057 _320_/D _238_/B 0.0334f
C18058 _315_/a_1108_7# _286_/Y 2.86e-19
C18059 _145_/A VPWR 0.951f
C18060 output28/a_27_7# VPWR 0.104f
C18061 _317_/a_27_7# _246_/B 1.49e-19
C18062 _165_/X _301_/a_240_7# 6.92e-20
C18063 _318_/Q _316_/a_1283_n19# 1.43e-19
C18064 _320_/Q _330_/a_761_249# 0.0184f
C18065 _342_/a_1108_7# _229_/a_226_7# 4.3e-19
C18066 _344_/a_193_7# _273_/A 3.42e-20
C18067 _271_/A _226_/X 0.176f
C18068 _146_/a_112_13# VPWR -9.59e-20
C18069 input4/X _323_/a_193_7# 1.05e-20
C18070 _162_/X _299_/a_215_7# 1.37e-20
C18071 _242_/A _328_/Q 0.231f
C18072 _169_/Y _284_/A 1.3e-20
C18073 _232_/X _248_/A 0.351f
C18074 _275_/Y _147_/A 0.00507f
C18075 _225_/B _284_/A 0.0103f
C18076 _337_/Q _309_/Q 0.00337f
C18077 _340_/a_1217_7# _197_/X 4.17e-20
C18078 _316_/Q _317_/a_27_7# 1.29e-19
C18079 _172_/A _190_/A 4.31e-19
C18080 _324_/a_27_7# _324_/Q 5.63e-19
C18081 _326_/a_543_7# _318_/Q 7.26e-20
C18082 _216_/A _336_/a_1283_n19# 3.71e-21
C18083 _325_/a_193_7# VGND 0.0202f
C18084 _325_/a_543_7# VPWR 0.00635f
C18085 _301_/X _299_/X 0.00158f
C18086 _333_/a_193_7# _298_/C 1.08e-20
C18087 _232_/X _331_/CLK 0.0823f
C18088 _273_/A _172_/A 0.109f
C18089 clkbuf_2_1_0_clk/A _267_/A 1.26f
C18090 _285_/A trim[4] 0.0586f
C18091 _271_/A _317_/a_761_249# 1.98e-19
C18092 _320_/a_761_249# _319_/a_651_373# 2.64e-21
C18093 _320_/a_651_373# _319_/a_761_249# 1.59e-21
C18094 _333_/a_448_7# _333_/D 0.0158f
C18095 _149_/a_27_7# VGND 0.065f
C18096 _257_/a_222_53# _255_/X 6.93e-21
C18097 _279_/Y _248_/a_109_257# 2e-19
C18098 _273_/A _232_/X 0.013f
C18099 _267_/A _310_/Q 3.88e-20
C18100 _333_/a_543_7# _332_/a_1283_n19# 1.29e-19
C18101 _333_/a_1283_n19# _332_/a_543_7# 5.68e-19
C18102 _333_/a_1108_7# _332_/a_761_249# 3.2e-20
C18103 _325_/a_1462_7# _304_/X 0.00223f
C18104 _297_/Y clkc 0.0116f
C18105 _317_/a_1270_373# VPWR 4.98e-19
C18106 _317_/a_448_7# VGND -0.00454f
C18107 _317_/Q _283_/A 9.62e-21
C18108 _236_/B _212_/a_27_7# 1.88e-19
C18109 _188_/S _143_/a_27_7# 2.01e-19
C18110 ctln[6] _336_/Q 3.56e-20
C18111 _323_/a_1283_n19# _343_/CLK 7.75e-20
C18112 _182_/a_510_7# _182_/X 3.62e-19
C18113 _283_/Y _338_/Q 0.0101f
C18114 _297_/A _347_/a_761_249# 0.0291f
C18115 _242_/A _269_/A 0.0156f
C18116 _161_/Y _346_/SET_B 0.0223f
C18117 _258_/a_505_n19# _313_/a_193_7# 6.6e-20
C18118 _336_/a_1217_7# _284_/A 1.51e-19
C18119 output36/a_27_7# input2/a_27_7# 0.0114f
C18120 _330_/Q _331_/a_1462_7# 4.02e-19
C18121 _337_/Q _311_/a_193_7# 0.00205f
C18122 repeater43/X _153_/B 0.00295f
C18123 _292_/A _312_/a_448_7# 5.99e-21
C18124 _232_/X _222_/a_93_n19# 7.88e-19
C18125 _197_/X _332_/D 4.82e-19
C18126 _314_/a_543_7# _284_/A 1.92e-21
C18127 _215_/A _344_/Q 6.33e-19
C18128 input1/a_75_172# VPWR 0.0898f
C18129 _248_/A _244_/B 0.34f
C18130 _309_/a_448_7# _309_/D 0.00198f
C18131 _290_/A _291_/a_39_257# 0.00999f
C18132 _331_/a_639_7# VGND 6.12e-19
C18133 output24/a_27_7# _325_/Q 1.25e-19
C18134 _304_/a_79_n19# _286_/B 8.25e-19
C18135 _320_/a_1462_7# _346_/SET_B 3.86e-19
C18136 _277_/Y _344_/Q 4.41e-20
C18137 _290_/Y trimb[0] 3.84e-19
C18138 _310_/a_193_7# clkc 6.82e-21
C18139 _320_/Q _322_/Q 0.246f
C18140 _256_/a_80_n19# _286_/B 9.73e-22
C18141 _279_/Y _147_/Y 0.00882f
C18142 _327_/a_27_7# _331_/Q 0.00878f
C18143 _331_/CLK _244_/B 0.34f
C18144 _306_/S _298_/A 0.569f
C18145 _343_/a_448_7# cal 0.00177f
C18146 _343_/a_1108_7# input1/X 9.59e-19
C18147 _270_/a_39_257# _325_/Q 0.0168f
C18148 _337_/a_543_7# _198_/a_250_257# 3.96e-21
C18149 _337_/a_1283_n19# _198_/a_93_n19# 1.09e-20
C18150 _190_/A _203_/a_80_n19# 0.00721f
C18151 _336_/a_651_373# _340_/Q 7.03e-21
C18152 _336_/a_448_7# _306_/S 6.06e-21
C18153 _254_/B _332_/Q 8.18e-19
C18154 _302_/a_227_7# _314_/Q 1.44e-19
C18155 _172_/A _307_/a_505_n19# 0.00177f
C18156 _323_/a_27_7# _226_/X 2.03e-21
C18157 _326_/a_27_7# _331_/Q 4.52e-21
C18158 _324_/Q _245_/a_113_257# 3.18e-21
C18159 _174_/a_27_257# VPWR 0.119f
C18160 _323_/D _248_/A 0.115f
C18161 _322_/D _269_/A 0.087f
C18162 _277_/Y _168_/a_109_7# 0.00201f
C18163 _182_/a_215_7# _298_/C 2.83e-21
C18164 _322_/a_1283_n19# _321_/D 0.00155f
C18165 _310_/a_193_7# _310_/a_543_7# -0.0102f
C18166 _308_/S _150_/C 5.9e-20
C18167 _321_/a_448_7# _269_/A 4.68e-21
C18168 _323_/a_543_7# _149_/A 1.05e-19
C18169 _324_/a_27_7# _228_/A 0.0483f
C18170 _334_/Q _153_/B 1.08e-20
C18171 _172_/A _178_/a_27_7# 3.48e-19
C18172 _219_/a_93_n19# _330_/Q 0.0387f
C18173 _344_/a_1182_221# _158_/Y 8.2e-19
C18174 _258_/a_76_159# _147_/A 0.00238f
C18175 output41/a_27_7# _298_/X 0.0295f
C18176 _186_/a_297_7# _225_/X 1.01e-21
C18177 _186_/a_79_n19# _226_/X 8.21e-19
C18178 _308_/X _226_/a_382_257# 1.31e-19
C18179 _196_/A _347_/a_27_7# 2.98e-20
C18180 _324_/a_448_7# _286_/Y 3.16e-19
C18181 _340_/CLK _312_/a_761_249# 2.86e-19
C18182 _309_/a_27_7# _174_/a_27_257# 9.74e-21
C18183 _188_/S _178_/a_193_257# 2.84e-19
C18184 repeater43/X _322_/a_193_7# -0.00112f
C18185 _342_/a_639_7# _248_/A 8.3e-19
C18186 _345_/a_27_7# _344_/D 2.32e-20
C18187 _309_/a_1108_7# _337_/Q 9.75e-19
C18188 _276_/a_68_257# clkbuf_2_1_0_clk/a_75_172# 7.29e-20
C18189 _191_/B _153_/B 3.34e-19
C18190 _339_/Q _311_/a_193_7# 0.00296f
C18191 clkbuf_2_1_0_clk/A _194_/X 0.0131f
C18192 _271_/Y clk 0.0709f
C18193 _292_/A _164_/A 0.0118f
C18194 repeater43/X _323_/a_805_7# 5.85e-19
C18195 _303_/A _279_/A 6.44e-20
C18196 _219_/a_250_257# _297_/B 9.84e-19
C18197 _345_/a_27_7# _346_/Q 2.7e-20
C18198 repeater43/X _214_/a_373_7# 4.17e-20
C18199 _330_/D _331_/a_1108_7# 2.32e-20
C18200 _320_/a_1283_n19# _217_/X 1.64e-19
C18201 _320_/a_1108_7# _212_/X 1.11e-20
C18202 output26/a_27_7# VPWR 0.1f
C18203 _324_/Q VPWR 2.35f
C18204 _164_/A _160_/A 2.57e-19
C18205 _167_/X _170_/a_76_159# 0.00748f
C18206 _164_/Y _162_/A 0.00442f
C18207 _250_/X _227_/A 3.67e-19
C18208 _324_/a_27_7# _216_/A 0.00541f
C18209 _214_/a_27_257# _212_/X 0.0524f
C18210 _214_/a_109_257# _327_/Q 0.0469f
C18211 _325_/a_1462_7# VGND -2.54e-19
C18212 _321_/a_193_7# _321_/a_761_249# -0.0105f
C18213 _321_/a_27_7# _321_/a_543_7# -0.00936f
C18214 _280_/a_68_257# _246_/B 3.19e-19
C18215 _157_/A _314_/Q 0.00581f
C18216 cal _311_/a_543_7# 1.11e-20
C18217 _320_/D _319_/a_1108_7# 2.63e-20
C18218 _167_/X clkbuf_2_1_0_clk/A 1.26f
C18219 _145_/a_113_7# _244_/B 1.61e-19
C18220 output15/a_27_7# ctlp[1] 0.00402f
C18221 _342_/a_761_249# repeater43/X -0.00312f
C18222 _193_/Y _194_/a_27_7# 2.23e-19
C18223 _338_/Q _312_/a_27_7# 2.23e-21
C18224 _255_/a_30_13# _154_/A 2.64e-21
C18225 _346_/SET_B _312_/a_543_7# 0.00248f
C18226 _315_/D _284_/A 0.0399f
C18227 _271_/A input1/X 0.00974f
C18228 input4/X _197_/X 1.07e-20
C18229 _166_/Y _299_/X 0.00845f
C18230 _313_/Q _313_/a_193_7# 0.00952f
C18231 _215_/A _306_/S 0.0164f
C18232 _306_/X _313_/a_27_7# 0.0047f
C18233 _290_/Y trimb[3] 0.00303f
C18234 _341_/Q _247_/a_113_257# 1.69e-20
C18235 ctln[4] _194_/X 5.08e-20
C18236 _277_/Y _306_/S 0.577f
C18237 _347_/a_193_7# _347_/a_543_7# -0.0129f
C18238 _341_/a_1283_n19# _177_/A 5.77e-20
C18239 _292_/A _312_/D 9.68e-20
C18240 _232_/X _217_/X 0.0761f
C18241 _236_/B _233_/a_113_257# 0.0486f
C18242 _168_/a_109_257# _160_/X 8.64e-21
C18243 _167_/X _300_/a_735_7# 1.84e-19
C18244 _341_/a_27_7# valid 2.12e-20
C18245 _210_/a_27_7# _209_/X 1.56e-19
C18246 _283_/A _298_/A 0.261f
C18247 _267_/A _311_/a_27_7# 0.102f
C18248 _269_/A _315_/a_1108_7# 0.015f
C18249 _161_/Y _147_/A 0.00388f
C18250 _163_/a_215_7# _147_/Y 1.5e-20
C18251 _260_/B _286_/B 0.00586f
C18252 output24/a_27_7# _315_/a_1283_n19# 6.01e-21
C18253 _317_/Q _315_/a_27_7# 3.22e-21
C18254 _294_/Y _310_/D 0.0148f
C18255 _179_/a_27_7# _225_/X 0.0222f
C18256 _329_/a_543_7# clkbuf_2_1_0_clk/A 3.51e-21
C18257 _197_/X _337_/a_1270_373# 3.4e-20
C18258 _275_/Y _174_/a_109_7# 0.00206f
C18259 _195_/a_27_257# VPWR 0.0854f
C18260 _281_/A VPWR 0.32f
C18261 _340_/a_27_7# _340_/a_193_7# -0.0343f
C18262 ctlp[5] _212_/X 2.5e-22
C18263 _346_/a_27_7# _162_/X 2.89e-19
C18264 _172_/A _296_/Y 0.0378f
C18265 _260_/A _314_/Q 1.44e-20
C18266 _255_/X _336_/Q 0.00775f
C18267 _342_/Q _225_/B 4.96e-20
C18268 _323_/a_761_249# clk 7.2e-19
C18269 _344_/Q VGND 0.646f
C18270 clkbuf_0_clk/X _330_/D 1.15e-19
C18271 _257_/a_544_257# _225_/B 0.00237f
C18272 _319_/Q _321_/Q 0.0153f
C18273 _325_/a_193_7# _214_/a_27_257# 5.18e-20
C18274 _279_/Y _256_/a_80_n19# 0.00104f
C18275 clkbuf_2_3_0_clk/A _254_/B 0.172f
C18276 _326_/a_193_7# _181_/X 5.88e-19
C18277 _271_/A _286_/Y 0.00703f
C18278 _228_/A VPWR 1.38f
C18279 _306_/S _304_/X 6.2e-20
C18280 _172_/A _146_/a_29_271# 3.82e-20
C18281 _308_/X _192_/B 0.0181f
C18282 ctlp[6] _281_/A 0.00818f
C18283 _248_/B _298_/A 1.84e-19
C18284 _239_/a_199_7# VGND -3.15e-19
C18285 _294_/A _215_/A 2.31e-19
C18286 _237_/a_113_257# _320_/Q 0.00256f
C18287 _331_/CLK _330_/a_805_7# 3.81e-19
C18288 _168_/a_397_257# VPWR 0.0234f
C18289 _168_/a_109_7# VGND 0.00228f
C18290 _207_/a_27_7# VGND 0.0473f
C18291 _207_/a_181_7# VPWR -2.98e-19
C18292 _294_/A _277_/Y 0.00865f
C18293 _297_/A _248_/A 1.63e-19
C18294 _172_/A clkbuf_0_clk/a_110_7# 0.143f
C18295 _319_/Q _297_/B 0.668f
C18296 _327_/a_193_7# _237_/a_113_257# 2.41e-20
C18297 _342_/a_1283_n19# _150_/C 0.00156f
C18298 _319_/Q _318_/a_193_7# 1.2e-20
C18299 _309_/a_761_249# _344_/Q 7.6e-21
C18300 repeater43/X _322_/a_1462_7# 3.18e-19
C18301 _346_/a_652_n19# _299_/a_78_159# 2.85e-19
C18302 _342_/Q _315_/a_448_7# 8.53e-21
C18303 _322_/a_27_7# result[7] 4.28e-20
C18304 _313_/a_27_7# _147_/Y 2e-19
C18305 _255_/B _227_/A 0.0211f
C18306 _297_/A _331_/CLK 4.53e-21
C18307 _301_/a_51_257# _170_/a_76_159# 0.00111f
C18308 _188_/S _183_/a_553_257# 5.52e-19
C18309 _323_/a_193_7# cal 0.00918f
C18310 _333_/a_1270_373# _332_/Q 1.85e-19
C18311 _323_/a_27_7# input1/X 4.25e-20
C18312 _254_/Y _336_/a_448_7# 0.0162f
C18313 _341_/a_193_7# _341_/a_651_373# -2.09e-19
C18314 _309_/a_1283_n19# _267_/A 7.49e-21
C18315 _279_/Y _332_/a_27_7# 4.76e-19
C18316 _320_/Q ctlp[1] 9.72e-20
C18317 _165_/X _346_/D 3.91e-21
C18318 _308_/S cal 2.32e-20
C18319 repeater43/X _330_/a_543_7# 0.00149f
C18320 _279_/Y _347_/a_193_7# 0.00126f
C18321 _216_/A VPWR 1.28f
C18322 _260_/B _347_/a_543_7# 4.42e-20
C18323 _332_/a_193_7# _208_/a_78_159# 1.14e-20
C18324 output33/a_27_7# VGND 0.0363f
C18325 _196_/A _190_/a_27_7# 0.0214f
C18326 _331_/D _327_/Q 0.0155f
C18327 _164_/Y _163_/a_78_159# 0.00144f
C18328 _273_/A _297_/A 6.56e-19
C18329 _316_/D _223_/a_250_257# 0.00325f
C18330 _314_/a_1283_n19# _297_/Y 1.24e-19
C18331 _330_/a_27_7# _212_/X 5.33e-20
C18332 output20/a_27_7# clkbuf_1_0_0_clk/a_75_172# 1.5e-19
C18333 clkbuf_2_1_0_clk/A _301_/a_51_257# 0.00453f
C18334 _251_/a_510_7# VPWR -9.97e-19
C18335 _251_/a_297_257# VGND -0.00181f
C18336 _338_/a_193_7# _338_/a_651_373# -0.00701f
C18337 _221_/a_584_7# VPWR -7.98e-19
C18338 result[4] _318_/a_1270_373# 6.15e-21
C18339 _221_/a_256_7# VGND -2.72e-19
C18340 _300_/Y _306_/S 2.26e-21
C18341 clkbuf_2_1_0_clk/A clkbuf_1_1_0_clk/a_75_172# 0.0109f
C18342 _318_/Q _212_/X 0.518f
C18343 _346_/SET_B _263_/B 0.00923f
C18344 _290_/A _297_/B 0.00619f
C18345 _186_/a_382_257# cal 8.66e-20
C18346 _324_/a_1283_n19# _296_/a_109_7# 1.43e-20
C18347 _273_/A _164_/A 2.3e-20
C18348 _344_/a_27_7# _174_/a_27_257# 0.00127f
C18349 _305_/a_505_n19# _337_/Q 7.21e-20
C18350 _215_/A _283_/A 0.00459f
C18351 _194_/X _311_/a_27_7# 1.92e-20
C18352 _192_/B _254_/B 0.00777f
C18353 _294_/Y _345_/a_193_7# 1.08e-20
C18354 _326_/a_1283_n19# _325_/D 2.42e-19
C18355 _251_/X _217_/A 6.56e-19
C18356 _277_/Y _283_/A 1.9e-20
C18357 _304_/X _327_/D 0.422f
C18358 _309_/a_27_7# _216_/A 5.32e-19
C18359 _334_/a_193_7# _298_/X 2.03e-20
C18360 _288_/A _338_/Q 1.14e-19
C18361 _322_/a_193_7# result[6] 0.025f
C18362 _333_/a_543_7# _206_/A 0.0401f
C18363 _333_/a_193_7# _207_/C 0.00964f
C18364 _232_/X _331_/a_805_7# 4.57e-19
C18365 _345_/a_1140_373# _290_/A 7.68e-19
C18366 _294_/Y _266_/a_113_257# 0.0104f
C18367 _290_/Y VPWR 0.393f
C18368 rstn _153_/A 2.04e-20
C18369 _323_/a_27_7# _286_/Y 1.17e-19
C18370 _182_/X _229_/a_556_7# 5.33e-21
C18371 clkbuf_0_clk/a_110_7# _203_/a_80_n19# 4.01e-21
C18372 _181_/X _295_/a_306_7# 0.00397f
C18373 _336_/a_27_7# _225_/B 5.27e-20
C18374 _336_/a_193_7# _336_/Q -1.36e-19
C18375 _275_/A _162_/X 4.53e-21
C18376 _200_/a_93_n19# _200_/a_346_7# -3.48e-20
C18377 ctln[7] clk 0.00237f
C18378 _164_/A _173_/a_556_7# 5.57e-20
C18379 _267_/A _311_/a_1217_7# 7.12e-20
C18380 _343_/CLK _333_/a_1283_n19# 4.29e-21
C18381 _292_/A _160_/A 9.11e-19
C18382 _269_/A output6/a_27_7# 9.93e-19
C18383 _317_/Q _242_/B 2.78e-19
C18384 clk _179_/a_27_7# 0.00437f
C18385 _242_/A _242_/a_109_257# 0.002f
C18386 _215_/A _248_/B 6.44e-20
C18387 _241_/a_113_257# _217_/X 6.31e-20
C18388 _241_/a_199_7# _212_/X 3.32e-20
C18389 _286_/B _333_/Q 0.00468f
C18390 trim[4] _164_/A 6.14e-20
C18391 _306_/S VGND 2.66f
C18392 _309_/a_651_373# _284_/A 8.49e-19
C18393 _299_/X _297_/Y 0.0406f
C18394 _317_/a_1108_7# _317_/D 9.98e-19
C18395 _177_/A _248_/A 0.0182f
C18396 repeater43/X _331_/Q 0.13f
C18397 _283_/A _304_/X 0.611f
C18398 _229_/a_556_7# valid 5.7e-20
C18399 _315_/a_27_7# _315_/a_193_7# -0.00693f
C18400 result[0] _341_/a_543_7# 8.92e-19
C18401 _340_/CLK _305_/X 5.69e-20
C18402 output11/a_27_7# ctln[5] 0.00197f
C18403 _325_/a_27_7# _331_/D 5.01e-20
C18404 _310_/a_1108_7# _310_/Q 0.00134f
C18405 _279_/Y _260_/B 0.00852f
C18406 _341_/Q _209_/X 6.2e-21
C18407 _227_/A _298_/a_27_7# 1.11e-20
C18408 _329_/a_543_7# _218_/a_93_n19# 2.29e-19
C18409 _199_/a_93_n19# _199_/a_256_7# -6.6e-20
C18410 _306_/a_76_159# _216_/A 2.02e-21
C18411 _308_/X _146_/C 0.00846f
C18412 _338_/a_27_7# _340_/CLK 0.0938f
C18413 _289_/a_121_257# _267_/B 7.52e-21
C18414 _256_/a_209_257# _190_/A 3.39e-19
C18415 _254_/Y _215_/A 4.87e-20
C18416 _327_/a_448_7# _216_/X 3.45e-19
C18417 _298_/C _295_/a_79_n19# 0.00106f
C18418 _283_/Y input1/X 5.13e-19
C18419 _290_/A _311_/a_1108_7# 0.00868f
C18420 _309_/a_761_249# _306_/S 1.08e-20
C18421 _277_/Y _254_/Y 7.39e-19
C18422 _160_/X comp 3.03e-20
C18423 _343_/a_1108_7# _343_/D 9.3e-21
C18424 _343_/a_651_373# _185_/A 0.00496f
C18425 _167_/a_27_257# _297_/B 0.0873f
C18426 _327_/a_1283_n19# _238_/B 1.13e-20
C18427 _342_/D _147_/A 2.07e-20
C18428 _327_/a_193_7# _327_/a_651_373# -0.00701f
C18429 _342_/Q _315_/D 0.398f
C18430 _248_/B _304_/X 0.258f
C18431 _232_/A _217_/A 3.76e-19
C18432 _308_/S _284_/A 1.93e-19
C18433 _322_/a_1217_7# result[7] 9.64e-22
C18434 _187_/a_27_7# _144_/a_27_7# 3.2e-20
C18435 _318_/Q _317_/a_448_7# 3.59e-20
C18436 _288_/A _345_/D 6.2e-21
C18437 _340_/a_761_249# _340_/CLK 6.15e-20
C18438 _144_/a_27_7# _315_/D 1.99e-20
C18439 _323_/a_1462_7# cal 3.67e-19
C18440 _342_/D _149_/A 0.0173f
C18441 _333_/D _190_/A 0.0054f
C18442 _248_/A _325_/D 3.2e-19
C18443 _341_/a_761_249# _341_/D 0.0221f
C18444 _290_/A _275_/Y 0.0164f
C18445 _315_/Q _316_/a_448_7# 6.05e-20
C18446 _294_/Y VPWR 0.414f
C18447 _294_/A VGND 2.48f
C18448 _329_/a_1270_373# _330_/Q 8.78e-20
C18449 _162_/X _345_/D 0.00217f
C18450 _161_/Y _174_/a_109_7# 7.38e-19
C18451 _313_/D _202_/a_93_n19# 3.03e-21
C18452 _272_/a_39_257# _283_/A 4.08e-19
C18453 _255_/B _297_/B 4.31e-20
C18454 _332_/a_193_7# _190_/A 1.23e-20
C18455 _332_/a_761_249# _333_/Q 0.014f
C18456 _332_/a_543_7# _332_/Q 4.32e-19
C18457 _346_/SET_B _194_/A 0.0103f
C18458 _277_/A clkbuf_2_1_0_clk/A 0.196f
C18459 _332_/a_1283_n19# _207_/X 2.26e-19
C18460 _331_/CLK _325_/D 0.00633f
C18461 _326_/a_193_7# _326_/a_651_373# -0.00701f
C18462 _328_/a_1108_7# _329_/Q 0.0056f
C18463 _328_/a_448_7# _320_/Q 5.91e-19
C18464 _317_/Q _245_/a_199_7# 4.76e-19
C18465 _307_/a_76_159# _286_/B 0.00571f
C18466 repeater43/X _333_/a_805_7# -0.00125f
C18467 _329_/a_1108_7# VGND 0.00207f
C18468 _329_/a_651_373# VPWR -0.00782f
C18469 _338_/a_761_249# _338_/D 0.043f
C18470 _338_/a_193_7# _346_/SET_B 0.0251f
C18471 _327_/D VGND 0.127f
C18472 _313_/D cal 1.05e-21
C18473 _180_/a_29_13# _298_/C 0.0311f
C18474 _197_/X _202_/a_93_n19# 0.0161f
C18475 _240_/a_109_257# VPWR 5.3e-19
C18476 _258_/S _346_/SET_B 0.044f
C18477 _273_/A _325_/D 6.54e-20
C18478 _341_/a_1283_n19# _248_/A 1.54e-21
C18479 _165_/a_78_159# _163_/a_78_159# 5.04e-19
C18480 _344_/a_652_n19# _344_/Q 1.4e-19
C18481 _342_/a_1283_n19# cal 0.00151f
C18482 _182_/a_79_n19# _191_/B 4.1e-22
C18483 _144_/A _223_/a_250_257# 2.02e-19
C18484 _294_/A _309_/a_761_249# 0.022f
C18485 _294_/Y _309_/a_27_7# 2.82e-21
C18486 _254_/A _162_/X 0.0583f
C18487 _319_/Q _320_/a_193_7# 6.54e-20
C18488 _343_/CLK output41/a_27_7# 0.0178f
C18489 cal _197_/X 0.087f
C18490 _298_/B _298_/A 0.126f
C18491 _263_/B _147_/A 9.79e-21
C18492 _315_/Q result[0] 0.104f
C18493 _300_/Y _248_/B 1.57e-20
C18494 _271_/A _269_/A 0.0139f
C18495 _340_/a_543_7# _346_/SET_B 0.00812f
C18496 _328_/a_27_7# _328_/a_448_7# -0.00642f
C18497 _325_/D _222_/a_93_n19# 2.27e-20
C18498 _197_/X _197_/a_27_7# 0.0307f
C18499 _145_/a_113_7# _177_/A 4.53e-21
C18500 _336_/a_1462_7# _336_/Q 1.15e-19
C18501 _283_/A VGND 4.74f
C18502 _320_/Q _346_/SET_B 0.0119f
C18503 _314_/a_543_7# _225_/B 0.00358f
C18504 _196_/A _339_/a_193_7# 6.65e-20
C18505 _227_/A _326_/Q 1.64e-19
C18506 _327_/a_193_7# _346_/SET_B 0.0101f
C18507 _271_/A _343_/D 4.32e-20
C18508 _205_/a_382_257# VGND -6.65e-19
C18509 _316_/a_1108_7# _248_/A 0.00608f
C18510 _163_/a_493_257# _160_/A 2.54e-19
C18511 _343_/a_543_7# _175_/Y 8.71e-19
C18512 _254_/B _202_/a_584_7# 0.00275f
C18513 _342_/a_193_7# sample 0.0198f
C18514 _342_/a_543_7# _286_/Y 5.9e-21
C18515 clkbuf_2_3_0_clk/A _196_/A 0.0123f
C18516 _292_/A _273_/A 0.214f
C18517 _242_/A _318_/a_27_7# 0.0129f
C18518 _331_/Q _331_/a_448_7# 0.0144f
C18519 result[7] _322_/Q 0.105f
C18520 _340_/a_448_7# _190_/A 8.77e-21
C18521 _319_/D _279_/A 2.31e-20
C18522 _316_/a_1283_n19# _316_/D 3.61e-20
C18523 _316_/a_1108_7# _331_/CLK 3.7e-19
C18524 _294_/A _306_/a_218_334# 7.09e-19
C18525 _327_/a_1283_n19# _248_/A 2.96e-20
C18526 _329_/a_193_7# _330_/D 0.0154f
C18527 _311_/a_1283_n19# _297_/Y 0.00143f
C18528 _343_/Q _226_/a_79_n19# 0.00382f
C18529 _279_/Y _333_/Q 3.81e-19
C18530 _325_/Q _318_/a_193_7# 1.35e-22
C18531 _301_/a_240_7# VPWR -0.00129f
C18532 _301_/a_512_257# VGND -5.06e-19
C18533 _238_/B _331_/CLK 0.282f
C18534 _273_/A _160_/A 0.649f
C18535 _328_/a_27_7# _346_/SET_B 0.0354f
C18536 _248_/B VGND 0.44f
C18537 _346_/SET_B _347_/a_805_7# -0.00125f
C18538 _330_/Q _234_/B 2.34e-19
C18539 _326_/a_1283_n19# _248_/A 0.0577f
C18540 _334_/a_27_7# _334_/a_448_7# -0.00642f
C18541 _334_/a_193_7# _334_/a_1108_7# -0.00656f
C18542 cal _312_/a_193_7# 9.22e-20
C18543 input1/X _312_/a_27_7# 2.78e-19
C18544 _200_/a_250_257# _338_/Q 4.36e-19
C18545 _293_/a_39_257# _194_/X 0.0011f
C18546 _204_/a_27_257# _332_/Q 0.0123f
C18547 _327_/a_1283_n19# _331_/CLK 0.0332f
C18548 _321_/a_1108_7# _321_/Q 0.0402f
C18549 _321_/a_1283_n19# _330_/Q 1.12e-19
C18550 _304_/a_79_n19# _144_/A 9.32e-20
C18551 _208_/a_493_257# _332_/Q 2.44e-20
C18552 _208_/a_215_7# _207_/X 0.00435f
C18553 _260_/A _254_/B 1.03f
C18554 clkbuf_0_clk/a_110_7# _297_/A 4.94e-21
C18555 _273_/A _238_/B 2.04e-20
C18556 _326_/a_1283_n19# _331_/CLK 5.87e-21
C18557 _326_/a_761_249# _236_/B 7e-22
C18558 _258_/S _313_/a_761_249# 1.19e-20
C18559 _341_/a_761_249# _343_/CLK 1.48e-21
C18560 _337_/Q _263_/a_109_257# 0.00161f
C18561 _305_/a_505_n19# _336_/D 0.00245f
C18562 _286_/B _313_/a_639_7# 3.37e-19
C18563 _314_/a_27_7# _314_/a_448_7# -0.00346f
C18564 _255_/a_30_13# _153_/B 9.22e-19
C18565 _311_/a_1108_7# _310_/a_27_7# 3.45e-20
C18566 _311_/a_1283_n19# _310_/a_193_7# 0.00117f
C18567 _311_/a_543_7# _310_/a_761_249# 2.05e-21
C18568 _311_/a_761_249# _310_/a_543_7# 6.99e-21
C18569 _321_/a_543_7# VPWR 0.032f
C18570 _321_/a_193_7# VGND 0.0233f
C18571 _327_/a_1283_n19# _273_/A 5.67e-19
C18572 _338_/a_761_249# _343_/CLK 8.57e-20
C18573 _254_/Y VGND 0.109f
C18574 repeater43/X valid 1.07e-19
C18575 ctln[6] _283_/Y 0.0139f
C18576 _292_/A trim[4] 8.11e-20
C18577 _322_/D _318_/a_27_7# 5.87e-20
C18578 _315_/Q _316_/D 0.00427f
C18579 _326_/a_1283_n19# _273_/A 2.16e-20
C18580 _321_/a_761_249# _318_/a_1283_n19# 1.84e-20
C18581 _321_/a_448_7# _318_/a_27_7# 3.02e-21
C18582 _313_/D _284_/A 3.97e-20
C18583 _323_/a_27_7# _269_/A 0.019f
C18584 _232_/X _221_/a_346_7# 1.39e-19
C18585 _153_/a_109_53# VPWR 0.0017f
C18586 _227_/A _154_/A 0.0128f
C18587 output31/a_27_7# _311_/a_193_7# 6.78e-20
C18588 _340_/a_1108_7# _337_/a_1283_n19# 6.64e-20
C18589 _340_/a_1283_n19# _337_/a_1108_7# 6.64e-20
C18590 output11/a_27_7# _206_/A 8.31e-20
C18591 _326_/a_761_249# _326_/D 2.33e-20
C18592 _260_/B _313_/a_27_7# 0.00395f
C18593 _298_/B _215_/A 3.15e-19
C18594 _275_/Y _310_/a_27_7# 0.0117f
C18595 _242_/A _246_/B 0.00709f
C18596 cal _333_/a_193_7# 1.09e-21
C18597 _288_/A _162_/a_27_7# 2.88e-20
C18598 _238_/B _319_/a_1108_7# 1.77e-19
C18599 _197_/X _284_/A 0.0132f
C18600 _310_/a_651_373# VGND 9.39e-19
C18601 _310_/a_639_7# VPWR 0.0045f
C18602 _162_/X _162_/a_27_7# 0.00177f
C18603 repeater43/X _332_/a_1108_7# 0.0132f
C18604 _165_/a_292_257# _158_/Y 8.87e-20
C18605 _196_/A _192_/B 0.25f
C18606 _319_/Q _322_/a_1108_7# 1.74e-21
C18607 _343_/D _323_/a_27_7# 0.0134f
C18608 _185_/A _323_/a_761_249# 0.0114f
C18609 _296_/Y _304_/a_257_159# 3.45e-20
C18610 _258_/a_218_7# _306_/S 0.00134f
C18611 _334_/a_1108_7# _332_/Q 3.49e-21
C18612 _334_/a_1283_n19# _333_/Q 1.41e-19
C18613 _231_/a_79_n19# _286_/Y 1.31e-20
C18614 result[1] result[2] 0.0461f
C18615 _316_/Q _242_/A 0.00248f
C18616 _228_/A _227_/a_113_7# 1.07e-19
C18617 _346_/a_652_n19# _346_/SET_B 0.0209f
C18618 _258_/S _147_/A 0.00271f
C18619 _315_/D _225_/B 7.44e-20
C18620 _325_/D _217_/X 4.23e-20
C18621 _325_/a_193_7# _286_/B 3.39e-19
C18622 _169_/a_109_257# VGND -0.0011f
C18623 _209_/a_27_257# VPWR 0.0983f
C18624 _225_/a_145_35# VGND 2.93e-19
C18625 output27/a_27_7# _321_/a_193_7# 1.22e-19
C18626 _347_/Q _314_/a_193_7# 5.77e-20
C18627 _339_/a_193_7# _338_/a_448_7# 1.94e-19
C18628 _339_/a_651_373# _338_/a_27_7# 2.22e-19
C18629 _339_/a_1108_7# _338_/a_761_249# 1.97e-19
C18630 _339_/a_1283_n19# _338_/a_543_7# 0.0027f
C18631 _271_/Y _335_/Q 1.26e-20
C18632 _342_/D _150_/a_27_7# 3.52e-20
C18633 _309_/a_1283_n19# _310_/a_1108_7# 4.62e-21
C18634 _309_/a_1108_7# _310_/a_1283_n19# 6.49e-20
C18635 _309_/a_651_373# _310_/a_761_249# 1.09e-20
C18636 _198_/a_346_7# _340_/Q 0.00406f
C18637 _198_/a_584_7# _194_/X 2.89e-19
C18638 _198_/a_250_257# _193_/Y 0.0507f
C18639 _290_/A _161_/Y 0.00778f
C18640 _146_/a_29_271# _177_/A 0.00759f
C18641 _335_/a_761_249# _335_/Q 0.00177f
C18642 _335_/a_193_7# _204_/Y 1.44e-20
C18643 _299_/X _170_/a_489_373# 1.13e-19
C18644 _347_/Q _170_/a_226_7# 0.00166f
C18645 _324_/a_193_7# _215_/A 2.67e-20
C18646 _327_/a_1462_7# _346_/SET_B 0.00117f
C18647 clkbuf_0_clk/X _162_/X 0.0114f
C18648 _308_/S _342_/Q 0.0476f
C18649 repeater43/X _341_/a_1270_373# -1.63e-20
C18650 _334_/Q _332_/a_1108_7# 0.00142f
C18651 _331_/CLK _248_/A 0.477f
C18652 _256_/a_209_257# clkbuf_0_clk/a_110_7# 8.66e-21
C18653 _343_/Q _323_/Q 0.103f
C18654 _346_/a_1032_373# _331_/CLK 6.18e-22
C18655 _340_/a_651_373# _339_/a_761_249# 1.09e-20
C18656 _340_/a_1283_n19# _339_/a_1108_7# 5.4e-21
C18657 _340_/a_1108_7# _339_/a_1283_n19# 2.22e-21
C18658 _334_/a_27_7# _206_/A 0.00406f
C18659 _342_/a_1462_7# sample 3.07e-20
C18660 _315_/a_448_7# _315_/D 0.00196f
C18661 _242_/A _318_/a_1217_7# 1.32e-19
C18662 _315_/a_27_7# VGND -0.00378f
C18663 _315_/a_761_249# VPWR 0.00631f
C18664 ctln[5] _339_/a_27_7# 1.22e-19
C18665 _285_/A comp 9.92e-20
C18666 _273_/A _248_/A 1.25f
C18667 input3/a_27_7# VPWR 0.156f
C18668 _342_/Q _186_/a_382_257# 0.00212f
C18669 _298_/C _226_/X 1.17e-20
C18670 _214_/a_27_257# _327_/D 3.02e-20
C18671 _324_/a_1108_7# _227_/A 1.04e-20
C18672 _336_/a_651_373# VPWR -0.00933f
C18673 _346_/a_1032_373# _273_/A 1.04e-19
C18674 _336_/a_1108_7# VGND 0.00324f
C18675 _324_/a_27_7# _324_/a_543_7# -0.00944f
C18676 _317_/a_193_7# _316_/a_27_7# 3.22e-19
C18677 _324_/a_193_7# _324_/a_761_249# -0.0105f
C18678 _328_/a_1217_7# _346_/SET_B -5.48e-19
C18679 _166_/Y _172_/B 7.4e-21
C18680 _306_/X _216_/A 5.18e-20
C18681 _334_/a_27_7# _334_/D 0.484f
C18682 _334_/a_193_7# _343_/CLK 0.00539f
C18683 repeater43/X _229_/a_226_7# 0.00624f
C18684 _315_/D _314_/a_543_7# 0.0373f
C18685 _337_/D _194_/A 0.00662f
C18686 _273_/A _331_/CLK 0.0269f
C18687 _346_/SET_B _319_/a_761_249# 0.0124f
C18688 _242_/B _304_/X 1.06e-19
C18689 _346_/SET_B _337_/a_27_7# 0.00773f
C18690 _338_/D _337_/a_193_7# 2.41e-19
C18691 _248_/A _222_/a_93_n19# 0.00976f
C18692 _289_/a_39_257# _284_/A 2.28e-21
C18693 _227_/A _324_/D 0.0388f
C18694 _224_/a_93_n19# VPWR 0.00221f
C18695 _216_/X _331_/a_193_7# 0.00237f
C18696 repeater43/X _316_/a_639_7# -2.15e-19
C18697 _300_/a_27_257# _300_/Y 0.00766f
C18698 _300_/a_301_257# _160_/X 0.0139f
C18699 _340_/Q _254_/B 0.0097f
C18700 _324_/a_193_7# _304_/X 0.00114f
C18701 _324_/a_27_7# _217_/A 1.61e-19
C18702 _314_/a_193_7# _297_/B 9.07e-19
C18703 _314_/a_27_7# _314_/D 0.0543f
C18704 _321_/a_1462_7# VGND -9.48e-19
C18705 _324_/Q _223_/a_250_257# 7.77e-20
C18706 rstn _335_/a_1270_373# 2.49e-19
C18707 _343_/a_27_7# _343_/a_193_7# -0.0287f
C18708 _322_/a_761_249# _269_/A 0.00583f
C18709 _341_/a_543_7# _145_/A 1.06e-20
C18710 _331_/CLK _222_/a_93_n19# 9.61e-19
C18711 _279_/Y _212_/X 6.29e-21
C18712 _330_/Q clkbuf_2_1_0_clk/A 0.0011f
C18713 _325_/a_761_249# _325_/D 0.043f
C18714 _337_/Q _312_/Q 1.8e-20
C18715 _308_/a_505_n19# _336_/Q 3.67e-20
C18716 result[5] _242_/A 1.23e-19
C18717 _238_/B _217_/X 3.43e-21
C18718 _171_/a_78_159# _297_/Y 1.02e-19
C18719 _153_/A VPWR 0.22f
C18720 ctlp[0] output28/a_27_7# 7.69e-19
C18721 output14/a_27_7# result[6] 0.0108f
C18722 _320_/a_27_7# _242_/A 4.98e-20
C18723 _215_/A _160_/X 2.67e-20
C18724 _327_/a_1283_n19# _217_/X 0.0154f
C18725 _327_/a_448_7# _327_/Q 0.00128f
C18726 _319_/a_1108_7# _331_/CLK 1.11e-21
C18727 _326_/a_1270_373# repeater43/X -2.06e-19
C18728 _273_/A _222_/a_93_n19# 0.0378f
C18729 _326_/a_27_7# _331_/a_543_7# 1.04e-20
C18730 _326_/a_543_7# _331_/a_27_7# 4.74e-20
C18731 _168_/a_397_257# _147_/Y 3.31e-21
C18732 _277_/Y _160_/X 0.6f
C18733 ctln[2] trim[3] 0.0563f
C18734 _207_/X _206_/A 0.0102f
C18735 _326_/a_1283_n19# _217_/X 0.00168f
C18736 ctlp[1] result[7] 0.0812f
C18737 _281_/Y _330_/a_448_7# 1.52e-19
C18738 _273_/A trim[4] 2.3e-19
C18739 _345_/a_193_7# _345_/a_1182_221# -2.22e-21
C18740 _343_/CLK _332_/Q 0.0209f
C18741 _334_/Q _204_/a_277_7# 5e-19
C18742 _162_/X _286_/Y 0.00996f
C18743 _275_/Y _169_/B 1.64e-21
C18744 _300_/a_383_7# VPWR 2.16e-19
C18745 _300_/a_27_257# VGND -0.00299f
C18746 _341_/a_1108_7# _149_/a_27_7# 4.2e-19
C18747 _342_/a_543_7# _269_/A 0.00804f
C18748 _334_/D _207_/X 0.00156f
C18749 ctln[6] _333_/a_27_7# 5.48e-21
C18750 _328_/a_1283_n19# _212_/X 1.04e-19
C18751 _328_/a_543_7# _217_/X 0.0119f
C18752 _162_/X _297_/a_27_257# 1.75e-19
C18753 _302_/a_227_7# _347_/a_1283_n19# 9.97e-20
C18754 _157_/A _196_/A 0.314f
C18755 _298_/B VGND 0.147f
C18756 _284_/a_39_257# VGND 0.0111f
C18757 _346_/a_1056_7# _346_/SET_B 0.0013f
C18758 _344_/a_193_7# _301_/a_149_7# 1.4e-20
C18759 _344_/a_27_7# _301_/a_240_7# 5.46e-22
C18760 _211_/a_109_7# _283_/A 0.00364f
C18761 _307_/a_505_n19# _190_/A 0.00133f
C18762 _216_/A _147_/Y 0.0281f
C18763 result[5] _322_/D 0.156f
C18764 _281_/Y _252_/a_27_7# 0.00124f
C18765 _325_/a_805_7# _181_/X 4.26e-19
C18766 output41/a_27_7# output30/a_27_7# 9.03e-19
C18767 _158_/Y _346_/SET_B 0.0107f
C18768 _194_/a_27_7# VGND 0.0458f
C18769 result[5] _321_/a_448_7# 2.96e-21
C18770 _290_/Y output16/a_27_7# 5.45e-20
C18771 _339_/a_193_7# _338_/D 0.00112f
C18772 _339_/a_27_7# _346_/SET_B 0.0142f
C18773 trim[2] _312_/a_193_7# 6.11e-21
C18774 _317_/Q _232_/X 6.96e-21
C18775 _340_/CLK _313_/a_448_7# 5.89e-20
C18776 _229_/a_489_373# _226_/X 0.00139f
C18777 input4/X _334_/a_639_7# 7.07e-20
C18778 repeater43/X _334_/a_651_373# 0.00149f
C18779 result[1] _315_/a_543_7# 2.48e-19
C18780 _316_/Q _315_/a_1108_7# 0.00146f
C18781 _337_/a_805_7# _340_/CLK 0.0021f
C18782 _335_/D _205_/a_297_7# 6.33e-19
C18783 _335_/a_1462_7# _204_/Y 7.37e-20
C18784 _235_/a_113_257# _330_/Q 0.0093f
C18785 _324_/Q _304_/a_79_n19# 0.00333f
C18786 _342_/a_543_7# _343_/D 2.36e-19
C18787 _200_/a_93_n19# _337_/Q 0.0385f
C18788 _342_/a_1108_7# _185_/A 1.28e-19
C18789 _172_/A _301_/a_149_7# 7.15e-21
C18790 _255_/X _305_/a_218_334# 3.91e-21
C18791 _339_/Q _312_/Q 0.086f
C18792 clkbuf_1_0_0_clk/a_75_172# _330_/a_543_7# 9.47e-20
C18793 clkbuf_2_3_0_clk/A _338_/D 1.43e-19
C18794 clkbuf_2_2_0_clk/a_75_172# _338_/Q 0.0016f
C18795 _345_/a_476_7# _160_/X 5.37e-20
C18796 _309_/a_193_7# _284_/a_121_257# 3.97e-20
C18797 _337_/a_193_7# _337_/a_1108_7# -0.00656f
C18798 _337_/a_27_7# _337_/a_448_7# -0.00346f
C18799 clkbuf_2_1_0_clk/a_75_172# clkbuf_2_1_0_clk/A 0.0353f
C18800 _344_/a_562_373# _297_/Y 0.0023f
C18801 _187_/a_27_7# _315_/D 1.36e-19
C18802 _340_/a_543_7# _339_/D 0.0089f
C18803 _334_/a_639_7# _207_/C 0.00425f
C18804 _242_/B VGND 0.169f
C18805 _318_/D VPWR 0.598f
C18806 _315_/a_1217_7# VGND 5.56e-20
C18807 _340_/a_193_7# _202_/a_93_n19# 8.43e-19
C18808 _320_/a_1270_373# _319_/D 5.63e-21
C18809 _324_/a_193_7# VGND -2.68e-19
C18810 _324_/a_543_7# VPWR 0.0139f
C18811 _342_/a_1283_n19# _342_/Q 0.0213f
C18812 _340_/CLK _191_/B 2.55e-20
C18813 _309_/a_193_7# _215_/A 5.31e-21
C18814 _326_/a_761_249# _325_/a_1283_n19# 6.36e-19
C18815 _326_/a_193_7# _325_/a_1108_7# 3.42e-19
C18816 _262_/a_113_257# VGND -0.00248f
C18817 _318_/a_1108_7# _242_/B 5.17e-19
C18818 _318_/a_543_7# _318_/D 4.36e-19
C18819 _347_/Q _279_/A 0.00244f
C18820 _196_/A _260_/A 0.617f
C18821 _318_/Q _327_/D 0.00539f
C18822 _277_/Y _309_/a_193_7# 1e-20
C18823 ctln[1] _334_/a_1108_7# 8.63e-19
C18824 _314_/a_805_7# VPWR 3.64e-19
C18825 _324_/a_1108_7# _297_/B 1.05e-20
C18826 _346_/SET_B _313_/a_651_373# 0.00472f
C18827 _343_/a_27_7# VGND 0.0385f
C18828 _343_/a_761_249# VPWR 0.012f
C18829 _340_/a_193_7# cal 7.67e-21
C18830 _340_/a_27_7# input1/X 1.29e-21
C18831 _180_/a_29_13# _150_/C 0.00779f
C18832 _346_/SET_B _337_/a_1217_7# -1.33e-20
C18833 _248_/A _217_/X 0.0797f
C18834 _317_/Q _244_/B 0.0356f
C18835 _157_/A _347_/a_1283_n19# 3.82e-19
C18836 clk _332_/a_1270_373# 4.42e-19
C18837 _217_/A VPWR 1.97f
C18838 repeater43/X _321_/D 0.168f
C18839 _160_/X _300_/Y 1.94e-21
C18840 _154_/a_27_7# _335_/Q 1.76e-21
C18841 _324_/a_1217_7# _217_/A 7.57e-20
C18842 _286_/B _344_/Q 1.45e-19
C18843 _340_/a_193_7# _197_/a_27_7# 8.64e-19
C18844 _346_/D VPWR 0.256f
C18845 _216_/A _223_/a_250_257# 0.00272f
C18846 ctln[7] _335_/Q 0.182f
C18847 _316_/D _212_/X 0.013f
C18848 _331_/CLK _217_/X 0.785f
C18849 _236_/B _327_/Q 0.00611f
C18850 _334_/a_448_7# _323_/Q 1.1e-19
C18851 _345_/a_1182_221# VPWR -0.00291f
C18852 _345_/a_652_n19# VGND 0.0105f
C18853 _297_/B _324_/D 0.00981f
C18854 _318_/a_1283_n19# _304_/X 3.31e-20
C18855 _179_/a_27_7# _335_/Q 3.26e-21
C18856 _259_/a_199_7# _261_/A 7.87e-19
C18857 _308_/S _225_/B 0.00227f
C18858 _322_/a_1283_n19# _242_/A 1.08e-19
C18859 _265_/B _311_/D 9.22e-21
C18860 _172_/B _297_/Y 0.00623f
C18861 _346_/SET_B _157_/a_27_7# 0.00692f
C18862 _200_/a_93_n19# _339_/Q 9.24e-20
C18863 _266_/a_199_7# VGND 1.94e-19
C18864 input1/X _298_/C 0.242f
C18865 _283_/A _330_/a_27_7# 0.001f
C18866 _345_/a_1602_7# _297_/B 1.3e-20
C18867 repeater42/a_27_7# _304_/X 0.0058f
C18868 _273_/A _217_/X 0.123f
C18869 _232_/A _317_/D 3.01e-19
C18870 _168_/a_109_7# _286_/B 3.83e-19
C18871 _318_/Q _283_/A 0.00628f
C18872 _339_/a_193_7# _337_/a_1108_7# 1.39e-19
C18873 _339_/a_761_249# _337_/a_1283_n19# 0.00117f
C18874 _339_/a_1283_n19# _337_/a_761_249# 0.00117f
C18875 _339_/a_1108_7# _337_/a_193_7# 1.39e-19
C18876 _330_/Q _218_/a_93_n19# 0.0124f
C18877 _326_/D _327_/Q 0.00759f
C18878 _341_/a_543_7# _324_/Q 4.46e-21
C18879 _256_/a_80_n19# _228_/A 1.2e-19
C18880 _277_/A _320_/a_651_373# 9.87e-19
C18881 _339_/a_193_7# _343_/CLK 1.43e-20
C18882 _337_/D _201_/a_27_7# 1.07e-19
C18883 _222_/a_250_257# _212_/X 0.00368f
C18884 _222_/a_256_7# _327_/Q 0.00273f
C18885 _222_/a_93_n19# _217_/X 0.00413f
C18886 _254_/Y _203_/a_209_257# 5.11e-20
C18887 _200_/a_250_257# input1/X 0.00407f
C18888 _200_/a_256_7# cal 0.00108f
C18889 _297_/B _279_/A 0.0309f
C18890 _272_/a_121_257# VPWR 1.18e-19
C18891 _245_/a_199_7# VGND -3.11e-19
C18892 _160_/X VGND 0.358f
C18893 _342_/a_193_7# _175_/Y 0.00196f
C18894 _290_/A _263_/B 0.0911f
C18895 _219_/a_93_n19# _216_/X 0.0221f
C18896 _260_/A _347_/a_1283_n19# 1.43e-21
C18897 input4/X _337_/a_639_7# 1.5e-20
C18898 _329_/a_761_249# _331_/Q 9.96e-21
C18899 _322_/a_1283_n19# _322_/D 1.42e-20
C18900 clkbuf_2_3_0_clk/A _343_/CLK 1.56e-19
C18901 _322_/a_1283_n19# _321_/a_448_7# 6.58e-21
C18902 _345_/Q _345_/D 0.0232f
C18903 _255_/B _231_/a_409_7# 2.74e-19
C18904 _294_/A output32/a_27_7# 0.00285f
C18905 _339_/a_1217_7# _346_/SET_B 1.3e-20
C18906 _226_/a_79_n19# _147_/A 0.0244f
C18907 _220_/a_250_257# VPWR 0.0225f
C18908 _329_/Q _219_/a_93_n19# 2.08e-20
C18909 _320_/Q _219_/a_250_257# 1e-19
C18910 _318_/Q _248_/B 4.68e-19
C18911 _188_/a_535_334# _150_/C 1.85e-19
C18912 ctln[2] _273_/Y 0.0293f
C18913 _325_/a_761_249# _248_/A 1.63e-19
C18914 _313_/D _336_/a_27_7# 7.85e-20
C18915 _337_/Q _340_/CLK 0.317f
C18916 _172_/A _298_/A 0.0093f
C18917 clk _295_/a_676_257# 4.19e-19
C18918 _304_/a_79_n19# _216_/A 0.0508f
C18919 _298_/C _286_/Y 0.15f
C18920 _149_/A _226_/a_79_n19# 0.00166f
C18921 _313_/a_27_7# _313_/a_639_7# -0.0015f
C18922 _256_/a_80_n19# _216_/A 6.68e-19
C18923 _289_/a_121_257# _297_/Y 1.75e-20
C18924 repeater43/X _304_/S 0.581f
C18925 _325_/a_761_249# _331_/CLK 3.29e-20
C18926 _325_/a_193_7# _316_/D 6.04e-21
C18927 _317_/Q _241_/a_113_257# 3.85e-19
C18928 _337_/a_27_7# _337_/D 0.146f
C18929 _335_/D _298_/A 1.8e-20
C18930 _167_/X _299_/a_78_159# 0.0109f
C18931 _197_/X _336_/a_27_7# 0.00132f
C18932 _320_/a_761_249# clkbuf_2_1_0_clk/A 1.62e-19
C18933 clkbuf_0_clk/a_110_7# _190_/A 6.26e-20
C18934 _317_/a_651_373# _248_/A 2.55e-19
C18935 output35/a_27_7# _162_/a_27_7# 9.56e-20
C18936 _339_/a_27_7# _339_/a_448_7# -0.00676f
C18937 _271_/A _318_/a_27_7# 2.74e-19
C18938 _328_/a_193_7# _219_/a_93_n19# 0.00121f
C18939 _328_/a_27_7# _219_/a_250_257# 6.49e-19
C18940 _273_/A _325_/a_761_249# 8.43e-20
C18941 _302_/a_539_257# _346_/SET_B 1.36e-19
C18942 ctln[0] VGND 0.0398f
C18943 _225_/a_59_35# _254_/B 0.0552f
C18944 _324_/a_1462_7# VGND -7.51e-19
C18945 _254_/A _313_/a_1283_n19# 0.0138f
C18946 _281_/Y _305_/X 2.58e-19
C18947 repeater43/X _225_/X 3.33e-20
C18948 _326_/D _325_/a_27_7# 0.00157f
C18949 _169_/B _161_/Y 0.00233f
C18950 _307_/X repeater43/X 3.34e-21
C18951 cal _229_/a_226_257# 7.95e-20
C18952 input1/X _229_/a_489_373# 0.0235f
C18953 _188_/S _224_/a_250_257# 1.57e-19
C18954 clkbuf_2_1_0_clk/A _311_/D 8.54e-20
C18955 ctln[1] _343_/CLK 0.0928f
C18956 _314_/Q VPWR 0.181f
C18957 _318_/a_1283_n19# VGND 0.0149f
C18958 _318_/a_448_7# VPWR -0.00144f
C18959 _183_/a_471_7# _180_/a_29_13# 1.9e-19
C18960 _341_/a_543_7# _228_/A 0.0112f
C18961 _196_/A _340_/Q 0.00426f
C18962 _323_/Q _206_/A 0.0912f
C18963 _343_/a_1217_7# VGND 4.56e-20
C18964 _286_/B _306_/S 2.93f
C18965 _315_/Q _324_/Q 0.375f
C18966 _325_/a_761_249# _222_/a_93_n19# 4.85e-19
C18967 _325_/a_193_7# _222_/a_250_257# 6.57e-19
C18968 _193_/Y _312_/D 2.29e-21
C18969 _346_/a_193_7# _301_/X 8.1e-20
C18970 repeater42/a_27_7# VGND 0.0176f
C18971 _307_/a_76_159# _145_/A 0.00254f
C18972 _211_/a_27_257# _153_/A 1.49e-19
C18973 _318_/a_27_7# _318_/a_639_7# -0.00188f
C18974 _309_/a_543_7# VPWR 0.0384f
C18975 _309_/a_193_7# VGND 0.0305f
C18976 repeater43/X _317_/a_27_7# 0.238f
C18977 _313_/a_651_373# _147_/A 0.00127f
C18978 _275_/Y _309_/Q 1.37e-21
C18979 _334_/D _323_/Q 9.09e-20
C18980 _343_/CLK _192_/B 0.0148f
C18981 _345_/a_1056_7# VGND 2.47e-19
C18982 _345_/a_1296_7# VPWR 2.11e-19
C18983 _339_/Q _340_/CLK 0.366f
C18984 _315_/a_193_7# _244_/B 0.0144f
C18985 _301_/a_240_7# _147_/Y 2.9e-19
C18986 _162_/A _344_/D 4.28e-20
C18987 _244_/B _298_/A 0.0668f
C18988 _307_/a_439_7# _191_/B 2.32e-19
C18989 _336_/a_1283_n19# _254_/B 2.41e-19
C18990 _283_/A _330_/a_1217_7# 7.3e-21
C18991 _341_/D _146_/C 0.00652f
C18992 _197_/X _199_/a_250_257# 0.00157f
C18993 _234_/B _233_/a_113_257# 0.0044f
C18994 clk _334_/a_805_7# 2.11e-19
C18995 _274_/a_39_257# _219_/a_93_n19# 5.13e-20
C18996 _165_/X _196_/A 0.00133f
C18997 _313_/D _225_/B 1.8e-19
C18998 _321_/a_1283_n19# _233_/a_113_257# 1.5e-19
C18999 _339_/D _337_/a_27_7# 1.09e-20
C19000 repeater43/X _331_/a_543_7# 0.00887f
C19001 _311_/a_193_7# _311_/a_1108_7# 1.42e-32
C19002 _311_/a_27_7# _311_/a_448_7# -0.0036f
C19003 _277_/Y _344_/a_193_7# 3.31e-20
C19004 _271_/A _246_/B 0.00581f
C19005 _191_/a_109_257# _323_/Q 0.00332f
C19006 _181_/a_27_7# _227_/A 0.00107f
C19007 _147_/A _157_/a_27_7# 0.0103f
C19008 _229_/a_76_159# sample 2.44e-19
C19009 _327_/a_27_7# _281_/Y 0.0128f
C19010 _309_/a_193_7# _309_/a_761_249# -0.0105f
C19011 _309_/a_27_7# _309_/a_543_7# -0.00951f
C19012 _331_/a_27_7# _212_/X 7.79e-19
C19013 _331_/a_193_7# _327_/Q 5.62e-20
C19014 output23/a_27_7# result[1] 0.00382f
C19015 _197_/X _225_/B 0.00587f
C19016 _172_/A _215_/A 0.0338f
C19017 _333_/a_761_249# _335_/Q 4.08e-21
C19018 _333_/a_193_7# _204_/Y 2.77e-20
C19019 _191_/B _225_/X 0.0106f
C19020 _330_/Q _328_/D 0.0058f
C19021 _294_/A _286_/B 0.0788f
C19022 _342_/a_1462_7# _175_/Y 5.5e-20
C19023 _307_/X _191_/B 0.151f
C19024 _321_/D result[6] 0.00239f
C19025 _319_/Q _320_/Q 0.0473f
C19026 _277_/Y _172_/A 0.00739f
C19027 _308_/a_439_7# VGND 0.0019f
C19028 _303_/A _347_/D 0.0335f
C19029 _275_/Y _311_/a_193_7# 0.00745f
C19030 _258_/S _290_/A 0.0324f
C19031 _316_/Q _271_/A 4.61e-19
C19032 _327_/a_193_7# _319_/Q -1.23e-36
C19033 trim[1] _297_/Y 1.12e-19
C19034 _288_/A clkc 4.05e-19
C19035 _306_/a_505_n19# VGND 0.065f
C19036 _306_/a_535_334# VPWR -8.05e-19
C19037 _149_/A _323_/Q 0.0291f
C19038 ctln[6] _332_/a_448_7# 0.00857f
C19039 _150_/C _226_/X 0.00475f
C19040 _311_/a_805_7# VPWR 0.00221f
C19041 _324_/Q _295_/a_512_7# 2.06e-19
C19042 _263_/B _310_/a_27_7# 1.65e-19
C19043 _271_/A _271_/Y 0.423f
C19044 _326_/a_193_7# _319_/Q 4.18e-21
C19045 cal _334_/a_639_7# 1.85e-19
C19046 _306_/X _336_/a_651_373# 1.75e-20
C19047 _327_/a_27_7# _329_/D 2.69e-20
C19048 _181_/X _296_/a_109_7# 0.00106f
C19049 _271_/Y _335_/a_27_7# 1.11e-19
C19050 _315_/Q _228_/A 0.005f
C19051 _346_/SET_B _202_/a_346_7# 7.7e-19
C19052 _335_/a_27_7# _335_/a_761_249# -0.0166f
C19053 clkbuf_1_1_0_clk/a_75_172# _299_/a_78_159# 1.31e-20
C19054 _217_/a_27_7# _212_/X 0.0189f
C19055 _260_/B _216_/A 0.0106f
C19056 _337_/Q _313_/a_543_7# 6.91e-21
C19057 output9/a_27_7# _275_/Y 0.0128f
C19058 _337_/a_651_373# _337_/Q 0.00164f
C19059 _345_/a_193_7# _344_/a_476_7# 9.08e-21
C19060 _345_/a_652_n19# _344_/a_652_n19# 3.55e-19
C19061 _345_/a_1182_221# _344_/a_27_7# 9.11e-19
C19062 _345_/a_476_7# _344_/a_193_7# 4.15e-20
C19063 _146_/C _143_/a_27_7# 0.0436f
C19064 trim[1] _310_/a_193_7# 7.46e-20
C19065 _288_/A _310_/a_543_7# 3.76e-22
C19066 _328_/a_27_7# _319_/Q 0.616f
C19067 _254_/A _302_/a_77_159# 0.00172f
C19068 _335_/a_1270_373# VPWR -2.59e-19
C19069 _335_/a_448_7# VGND -7.77e-19
C19070 cal _338_/Q 0.211f
C19071 _184_/a_218_7# VPWR -4.21e-19
C19072 _184_/a_218_334# VGND -4.29e-19
C19073 _309_/a_193_7# _306_/a_218_334# 6.02e-21
C19074 _235_/a_113_257# _212_/a_27_7# 4.12e-20
C19075 _339_/a_27_7# _339_/D 0.189f
C19076 _320_/a_193_7# _279_/A 1.55e-20
C19077 _286_/B _283_/A 0.0106f
C19078 _338_/a_448_7# _340_/Q 0.00981f
C19079 _338_/a_651_373# _194_/X 0.00387f
C19080 _333_/a_1108_7# _153_/a_109_53# 3.41e-20
C19081 _333_/a_1283_n19# _153_/a_215_257# 0.0161f
C19082 repeater43/X clk 0.423f
C19083 _326_/D _325_/a_1217_7# 4.27e-20
C19084 _232_/X _304_/X 0.0879f
C19085 _325_/a_448_7# repeater43/X 8.79e-20
C19086 _215_/A _203_/a_80_n19# 1.12e-19
C19087 _313_/Q clkbuf_2_1_0_clk/A 0.0182f
C19088 _317_/a_27_7# _317_/a_543_7# -0.00482f
C19089 _302_/a_539_257# _147_/A 0.00135f
C19090 _325_/a_543_7# _212_/X 0.00138f
C19091 _165_/X _165_/a_78_159# 0.00626f
C19092 _344_/a_652_n19# _160_/X 1.45e-20
C19093 _346_/a_796_7# _301_/X 4.56e-20
C19094 _308_/a_76_159# _308_/S 2.83e-19
C19095 _157_/A _313_/a_193_7# 0.00707f
C19096 _346_/SET_B _267_/A 0.0751f
C19097 _309_/a_1462_7# VGND -8.78e-19
C19098 repeater43/X _317_/a_1217_7# 5.29e-19
C19099 _146_/C _343_/CLK 8.11e-19
C19100 _340_/a_651_373# _306_/S 0.00432f
C19101 ctln[5] _194_/X 3.25e-19
C19102 _279_/Y _306_/S 0.0792f
C19103 _336_/a_651_373# _147_/Y 6.7e-20
C19104 _286_/B _248_/B 7.2e-20
C19105 _285_/A trimb[1] 0.0013f
C19106 _276_/a_68_257# clkbuf_2_3_0_clk/A 2e-20
C19107 _322_/a_193_7# _321_/Q 0.0083f
C19108 _172_/A _300_/Y 4.32e-20
C19109 _255_/B _194_/A 7.65e-20
C19110 output13/a_27_7# ctln[0] 3e-19
C19111 ctln[7] output6/a_27_7# 1.2e-19
C19112 _163_/a_215_7# _344_/Q 4.46e-19
C19113 _333_/a_1283_n19# _209_/a_109_257# 0.00123f
C19114 _333_/a_1108_7# _209_/a_27_257# 0.00111f
C19115 clk _334_/Q 0.0605f
C19116 _340_/CLK _336_/D 0.00115f
C19117 _337_/Q _267_/B 0.159f
C19118 _271_/Y _323_/a_27_7# 2.03e-20
C19119 _321_/a_805_7# _322_/Q 1.81e-19
C19120 _346_/a_476_7# _346_/Q 0.00474f
C19121 _346_/a_193_7# _166_/Y 5.16e-21
C19122 _269_/A _298_/C 3.67e-20
C19123 _339_/Q _337_/a_651_373# 0.0282f
C19124 _307_/a_76_159# _324_/Q 5.47e-19
C19125 _311_/a_27_7# _311_/D 0.15f
C19126 trim[0] VPWR 0.284f
C19127 _343_/a_193_7# _244_/B 1.78e-21
C19128 _285_/A VGND 1.28f
C19129 _330_/Q _214_/a_109_7# 2.92e-19
C19130 _272_/a_39_257# _232_/X 0.00112f
C19131 _232_/a_27_7# _246_/B 1.04e-20
C19132 _304_/a_306_329# _248_/B 0.0022f
C19133 _258_/S _257_/a_79_159# 0.00102f
C19134 _320_/a_448_7# VPWR 0.00147f
C19135 _320_/a_1283_n19# VGND 0.0235f
C19136 repeater43/X _280_/a_68_257# 1.17e-19
C19137 _277_/A ctlp[3] 5.12e-20
C19138 _254_/Y _286_/B 0.0188f
C19139 _323_/a_1270_373# VPWR 5.95e-21
C19140 _323_/a_448_7# VGND 0.00122f
C19141 _145_/A _149_/a_27_7# 8.21e-19
C19142 output18/a_27_7# clkbuf_2_1_0_clk/A 0.0561f
C19143 _181_/a_27_7# _297_/B 3.37e-19
C19144 output39/a_27_7# output17/a_27_7# 5.88e-21
C19145 _214_/a_109_257# VPWR -0.018f
C19146 _322_/a_193_7# _318_/a_193_7# 2.64e-20
C19147 _322_/a_27_7# _318_/a_761_249# 8.42e-22
C19148 clk _191_/B 0.368f
C19149 input1/X _207_/C 1.8e-20
C19150 _292_/A output5/a_27_7# 3.25e-20
C19151 _344_/a_193_7# VGND 0.0132f
C19152 _344_/a_476_7# VPWR 0.0512f
C19153 _232_/X _220_/a_93_n19# 0.00128f
C19154 ctlp[7] _283_/A 0.0712f
C19155 _318_/Q _242_/B 0.0898f
C19156 input1/X _313_/a_1283_n19# 7.1e-21
C19157 _194_/A _310_/a_27_7# 7.14e-20
C19158 _346_/SET_B _221_/a_93_n19# 6.71e-19
C19159 _320_/a_1270_373# _297_/B 3.05e-19
C19160 _343_/D _298_/C 4.96e-20
C19161 cal _337_/a_639_7# 2.01e-19
C19162 _186_/a_297_7# _271_/A 0.00208f
C19163 _207_/a_181_7# _333_/Q 4.47e-19
C19164 _343_/a_193_7# _323_/D 0.013f
C19165 _345_/a_1602_7# _161_/Y 0.0166f
C19166 ctln[6] _332_/D 0.18f
C19167 _344_/a_1032_373# _297_/B 1.6e-20
C19168 _260_/A _313_/a_193_7# 2.15e-20
C19169 _311_/Q VPWR 0.202f
C19170 _258_/a_535_334# VGND -1.68e-19
C19171 _258_/a_439_7# VPWR -3.68e-19
C19172 _285_/A _309_/a_761_249# 7.1e-21
C19173 _277_/A _299_/a_78_159# 4.98e-20
C19174 _325_/a_193_7# _325_/a_543_7# -0.0102f
C19175 _325_/a_27_7# _325_/a_1283_n19# -9.15e-20
C19176 _161_/Y _309_/Q 1.63e-19
C19177 _258_/S _310_/a_27_7# 0.0299f
C19178 _172_/A VGND 2.19f
C19179 _308_/X VPWR 1.09f
C19180 result[4] _321_/D 2.25e-19
C19181 _338_/Q _284_/A 1.64e-19
C19182 _342_/a_27_7# VPWR 0.0753f
C19183 _254_/A cal 2.67e-20
C19184 _292_/A comp 3.35e-20
C19185 _312_/Q _310_/a_1283_n19# 2.44e-19
C19186 _346_/Q _173_/a_489_373# 6.46e-20
C19187 _255_/X _298_/C 9.37e-20
C19188 _211_/a_373_7# VPWR -4.76e-19
C19189 _211_/a_109_257# VGND -0.00224f
C19190 _198_/a_346_7# VPWR -7.08e-19
C19191 _198_/a_250_257# VGND -0.00277f
C19192 _232_/X VGND 1.39f
C19193 _335_/D VGND 0.292f
C19194 _341_/a_639_7# _269_/A 6.35e-19
C19195 _340_/D _190_/a_27_7# 1.77e-19
C19196 _245_/a_113_257# _317_/D 0.00334f
C19197 _303_/A _304_/S 0.00193f
C19198 _267_/A _313_/a_761_249# 2.04e-20
C19199 comp _160_/A 1.19e-19
C19200 _343_/a_651_373# _342_/a_543_7# 1.8e-21
C19201 _343_/a_1108_7# _342_/a_1108_7# 2.44e-20
C19202 _219_/a_93_n19# _327_/Q 0.00109f
C19203 _339_/Q _267_/B 0.0122f
C19204 _338_/a_1108_7# _283_/A 8.39e-21
C19205 _169_/a_109_257# _286_/B 1.15e-19
C19206 _319_/Q _319_/a_761_249# 0.00571f
C19207 _196_/A _225_/a_59_35# 4.51e-19
C19208 _242_/B _241_/a_199_7# 2.22e-34
C19209 _232_/X _318_/a_1108_7# 2.08e-21
C19210 output32/a_27_7# _284_/a_39_257# 9.03e-19
C19211 _338_/D _340_/Q 0.0103f
C19212 _346_/SET_B _194_/X 0.28f
C19213 _333_/a_1108_7# _153_/A 0.00814f
C19214 cal _226_/X 0.00426f
C19215 input1/X _150_/C 0.0947f
C19216 _224_/a_250_257# _223_/a_93_n19# 1.47e-19
C19217 _307_/a_76_159# _228_/A 8.19e-22
C19218 _323_/a_27_7# _323_/a_761_249# -6.54e-19
C19219 _324_/Q _212_/X 0.00198f
C19220 rstn _332_/a_543_7# 5.16e-20
C19221 cal _309_/D 9.82e-20
C19222 _271_/A _154_/a_27_7# 0.00165f
C19223 _290_/A _173_/a_226_7# 3.48e-21
C19224 _241_/a_113_257# _304_/X 5.76e-20
C19225 _279_/Y _283_/A 0.00838f
C19226 _283_/Y _271_/Y 2.55e-19
C19227 _328_/a_1270_373# _328_/Q 1.44e-19
C19228 _346_/a_1602_7# _306_/S 2.48e-20
C19229 _283_/Y _335_/a_761_249# 1.21e-19
C19230 ctln[7] _335_/a_27_7# 0.0504f
C19231 _182_/a_79_n19# _227_/A 0.0112f
C19232 _317_/Q _316_/a_1108_7# 6.56e-19
C19233 result[2] _316_/a_543_7# 1.84e-19
C19234 _203_/a_80_n19# VGND 0.0544f
C19235 _203_/a_209_7# VPWR -6.62e-19
C19236 _286_/B _336_/a_1108_7# 0.0046f
C19237 _345_/a_381_7# _172_/B 5.7e-20
C19238 _167_/X _346_/SET_B 0.0331f
C19239 _339_/a_761_249# _195_/a_27_257# 7.65e-21
C19240 _339_/a_193_7# _195_/a_109_257# 6.22e-21
C19241 _254_/B VPWR 0.403f
C19242 _271_/A _322_/a_1283_n19# 8.83e-19
C19243 _244_/B VGND 0.449f
C19244 _317_/D VPWR 1.07f
C19245 _297_/A _300_/a_301_257# 2.33e-19
C19246 _185_/A _229_/a_556_7# 0.00294f
C19247 _322_/a_1462_7# _321_/Q 5.11e-19
C19248 _340_/D _332_/Q 4.29e-21
C19249 _164_/Y _310_/D 0.0157f
C19250 _267_/A _147_/A 0.387f
C19251 _346_/a_1224_7# _346_/Q 2.7e-19
C19252 _327_/a_27_7# _242_/A 1.63e-19
C19253 _326_/a_1108_7# _283_/A 0.0101f
C19254 _343_/Q _175_/Y 0.223f
C19255 _231_/a_676_257# _315_/D 2.58e-19
C19256 _307_/a_76_159# _216_/A 1.89e-19
C19257 _340_/a_193_7# _336_/a_27_7# 2.51e-22
C19258 _340_/a_27_7# _336_/a_193_7# 2.81e-21
C19259 _146_/a_184_13# _146_/C 3.7e-19
C19260 _318_/a_543_7# _317_/D 0.00121f
C19261 _322_/a_805_7# VPWR 3.85e-19
C19262 _150_/C _286_/Y 0.0112f
C19263 _326_/a_1283_n19# _317_/Q 0.0119f
C19264 _315_/a_193_7# _177_/A 2.16e-20
C19265 _313_/a_1108_7# _284_/A 0.00635f
C19266 _330_/Q _330_/a_761_249# 0.00199f
C19267 _177_/A _298_/A 0.0392f
C19268 _326_/a_27_7# _242_/A 0.604f
C19269 _279_/Y _248_/B 0.114f
C19270 _346_/D _147_/Y 0.0413f
C19271 _337_/a_639_7# _284_/A 4.11e-20
C19272 _320_/D VGND 0.171f
C19273 clkbuf_2_3_0_clk/A _344_/D 2.84e-20
C19274 _323_/D VGND 0.44f
C19275 _302_/a_323_257# _301_/X 3.63e-19
C19276 _162_/X _314_/a_1283_n19# 2.56e-20
C19277 ctln[6] input4/X 0.0108f
C19278 _281_/Y repeater43/X 3.15e-19
C19279 _331_/D VPWR 0.134f
C19280 _344_/a_796_7# VGND 1.26e-19
C19281 _344_/a_1224_7# VPWR 2.92e-19
C19282 _281_/A _212_/X 3.07e-20
C19283 _342_/Q _295_/a_79_n19# 0.0758f
C19284 _255_/B _295_/a_306_7# 8.46e-19
C19285 _330_/a_193_7# VPWR -0.289f
C19286 _329_/a_543_7# _346_/SET_B -9.96e-19
C19287 _309_/a_1108_7# _161_/Y 6e-21
C19288 clkbuf_2_3_0_clk/A _346_/Q 0.407f
C19289 _342_/a_1108_7# _271_/A 5.67e-21
C19290 _164_/A _215_/A 0.0024f
C19291 _254_/A _284_/A 0.0994f
C19292 _333_/D _298_/A 6.43e-20
C19293 _308_/X _184_/a_505_n19# 0.0213f
C19294 _325_/a_193_7# _324_/Q 8.79e-20
C19295 _291_/a_39_257# _312_/Q 0.0105f
C19296 _227_/A _333_/a_805_7# 1.27e-21
C19297 _277_/Y _164_/A 8.86e-21
C19298 _279_/Y _254_/Y 4.01e-19
C19299 _194_/X _313_/a_761_249# 4.21e-22
C19300 _306_/S _313_/a_27_7# 2.28e-19
C19301 _168_/a_481_7# clkbuf_2_3_0_clk/A 4.91e-20
C19302 _228_/A _212_/X 3.96e-20
C19303 ctln[6] _207_/C 2.69e-19
C19304 _337_/a_1283_n19# _306_/S 0.00956f
C19305 _337_/a_193_7# _340_/D 1.73e-20
C19306 _337_/a_543_7# _193_/Y 1.3e-20
C19307 _337_/a_1108_7# _340_/Q 0.00384f
C19308 _318_/Q _318_/a_1283_n19# 0.0772f
C19309 _342_/a_639_7# VGND -0.00138f
C19310 _342_/a_1217_7# VPWR 8.96e-20
C19311 _305_/X _336_/Q 2.92e-21
C19312 _290_/A _158_/Y 3.05e-19
C19313 _346_/Q _172_/Y 3.58e-19
C19314 repeater43/X _329_/D 2.97e-19
C19315 _343_/CLK _340_/Q 4.08e-19
C19316 _286_/B _300_/a_27_257# 2.04e-20
C19317 repeater42/a_27_7# _318_/Q 0.104f
C19318 _273_/A output5/a_27_7# 0.00523f
C19319 _329_/a_448_7# _331_/CLK 0.0063f
C19320 _286_/B _298_/B 2.05e-19
C19321 _297_/A _304_/X 2.18e-19
C19322 _314_/a_27_7# _347_/a_27_7# 1.1e-19
C19323 _258_/S _169_/B 1.44e-20
C19324 _343_/a_1283_n19# _342_/D 8.24e-21
C19325 _286_/B _194_/a_27_7# 0.00144f
C19326 _160_/X output40/a_27_7# 3.35e-19
C19327 _306_/a_76_159# _254_/B 1.5e-21
C19328 _265_/B _162_/A 0.246f
C19329 _241_/a_113_257# VGND -0.003f
C19330 _170_/a_76_159# _347_/a_27_7# 2.86e-21
C19331 _320_/a_27_7# _320_/a_639_7# -0.00188f
C19332 _217_/A _223_/a_250_257# 0.00732f
C19333 _304_/X _223_/a_256_7# 0.00219f
C19334 _162_/X _299_/X 0.573f
C19335 _309_/D _284_/A 0.0545f
C19336 _312_/a_543_7# _311_/a_193_7# 1.37e-20
C19337 _312_/a_761_249# _311_/a_761_249# 1.8e-21
C19338 _321_/Q _331_/Q 0.213f
C19339 _330_/Q _322_/Q 6.49e-19
C19340 _340_/a_761_249# _336_/Q 4.11e-21
C19341 _216_/A _212_/X 0.0811f
C19342 _341_/a_543_7# _315_/a_761_249# 2.05e-21
C19343 _341_/a_1108_7# _315_/a_27_7# 4.2e-21
C19344 _341_/a_27_7# _315_/a_1108_7# 7.13e-19
C19345 _341_/a_761_249# _315_/a_543_7# 2.04e-21
C19346 _281_/Y _191_/B 0.0123f
C19347 _341_/a_1283_n19# _298_/A 0.0347f
C19348 _273_/A comp 2.5e-19
C19349 _332_/a_27_7# _153_/A 6.68e-19
C19350 _229_/a_76_159# _175_/Y 0.0332f
C19351 _318_/a_1108_7# _241_/a_113_257# 1.87e-19
C19352 _345_/a_193_7# _164_/Y 8.08e-20
C19353 _345_/a_476_7# _164_/A 1.32e-19
C19354 _202_/a_93_n19# _202_/a_250_257# -6.97e-22
C19355 _341_/D _232_/A 2.19e-22
C19356 _277_/Y _312_/D 3e-19
C19357 _194_/X _147_/A 6.57e-22
C19358 _317_/Q _248_/A 0.0077f
C19359 _344_/a_193_7# _344_/a_652_n19# -5.22e-20
C19360 _344_/a_27_7# _344_/a_476_7# -0.0112f
C19361 output35/a_27_7# clkc 0.00168f
C19362 _283_/A _316_/D 0.197f
C19363 _301_/a_51_257# _346_/SET_B 8.42e-21
C19364 _346_/a_193_7# _242_/A 2.32e-20
C19365 ctlp[4] _297_/B 6.51e-20
C19366 _341_/Q _343_/Q 1.64e-21
C19367 _346_/SET_B clkbuf_1_1_0_clk/a_75_172# 4.01e-19
C19368 output13/a_27_7# _335_/D 9.42e-20
C19369 _340_/CLK _310_/a_1283_n19# 9.11e-21
C19370 _182_/X _227_/A 2.98e-19
C19371 _267_/a_109_257# _193_/Y 3.46e-20
C19372 input1/X _202_/a_93_n19# 4.42e-20
C19373 _317_/Q _331_/CLK 0.416f
C19374 _236_/B _230_/a_27_7# 0.0358f
C19375 _339_/a_1108_7# _340_/Q 0.00153f
C19376 _339_/a_193_7# _340_/D 0.016f
C19377 _339_/a_543_7# _193_/Y 0.00562f
C19378 _312_/a_1270_373# VPWR 1.14e-19
C19379 _312_/a_448_7# VGND 0.00179f
C19380 _297_/A _300_/Y 0.0102f
C19381 rstn _334_/a_1108_7# 6.12e-21
C19382 _299_/X _299_/a_493_257# 9.1e-21
C19383 _294_/A _254_/a_109_257# 1.97e-19
C19384 cal input1/X 0.0724f
C19385 _273_/A _317_/Q 4.27e-19
C19386 _149_/a_27_7# _228_/A 3.35e-21
C19387 _304_/a_578_7# _227_/A 0.00206f
C19388 _316_/a_543_7# _315_/a_543_7# 3.02e-21
C19389 _316_/a_1108_7# _315_/a_193_7# 7.76e-20
C19390 _167_/X _147_/A 6.15e-21
C19391 input4/X _269_/A 0.00198f
C19392 _326_/a_193_7# _326_/Q 0.00475f
C19393 _144_/A _306_/S 1.69e-20
C19394 _232_/X _214_/a_27_257# 0.0124f
C19395 input1/X _197_/a_27_7# 2.14e-21
C19396 _339_/Q _261_/a_109_257# 0.00481f
C19397 _292_/Y _275_/A 0.0345f
C19398 _236_/B _232_/A 0.106f
C19399 _316_/D _248_/B 0.0012f
C19400 rstn _338_/D 1.18e-19
C19401 _301_/X _303_/A 3.46e-19
C19402 _255_/a_30_13# _225_/X 1.5e-19
C19403 clkbuf_2_1_0_clk/A _338_/a_761_249# 9e-22
C19404 _342_/a_1108_7# _186_/a_79_n19# 6.65e-20
C19405 _188_/a_439_7# _255_/B 0.00222f
C19406 _309_/Q _263_/B 3.11e-19
C19407 _319_/Q _317_/a_1283_n19# 2.97e-21
C19408 _304_/a_257_159# _304_/X 9.21e-19
C19409 _330_/a_805_7# VGND 2.78e-19
C19410 _162_/a_27_7# _284_/A 1.59e-19
C19411 _343_/a_193_7# _177_/A 3.13e-21
C19412 _269_/A _207_/C 0.00942f
C19413 _337_/a_1283_n19# _283_/A 3.02e-19
C19414 repeater43/X _185_/A 0.376f
C19415 _321_/a_193_7# _316_/D 1.03e-20
C19416 _321_/a_761_249# _331_/CLK 0.0428f
C19417 _143_/a_27_7# _232_/A 4.01e-20
C19418 _338_/Q _310_/a_761_249# 9.17e-20
C19419 _346_/SET_B _310_/a_1108_7# -0.00865f
C19420 _325_/a_193_7# _216_/A 4.88e-19
C19421 _333_/a_1270_373# VPWR 1.16e-19
C19422 _333_/a_448_7# VGND -0.00251f
C19423 _342_/a_193_7# _188_/S 1.73e-21
C19424 _242_/A _319_/a_193_7# 0.00966f
C19425 _283_/Y ctln[7] 0.0222f
C19426 _297_/A VGND 1.38f
C19427 _337_/D _194_/X 0.0273f
C19428 _315_/Q _315_/a_761_249# 1.41e-19
C19429 _343_/a_761_249# _176_/a_27_7# 0.00165f
C19430 _346_/Q _302_/a_227_7# 5.45e-20
C19431 output21/a_27_7# VPWR 0.136f
C19432 _290_/A _160_/a_27_7# 4.25e-21
C19433 _198_/a_93_n19# _198_/a_346_7# -3.48e-20
C19434 _281_/Y _337_/Q 1.79e-20
C19435 _334_/a_448_7# _175_/Y 1.27e-20
C19436 _216_/X clkbuf_2_1_0_clk/A 1.35e-19
C19437 _174_/a_27_257# _344_/Q 0.0403f
C19438 cal _286_/Y 0.0015f
C19439 _336_/a_761_249# _340_/CLK 3.33e-20
C19440 _343_/D _207_/C 0.00131f
C19441 _153_/a_109_53# _333_/Q 0.0352f
C19442 _153_/a_215_257# _332_/Q 0.0672f
C19443 _286_/B _160_/X 0.0136f
C19444 _343_/CLK _205_/a_79_n19# 1.25e-19
C19445 _223_/a_256_7# VGND -0.00141f
C19446 _223_/a_584_7# VPWR -8.86e-19
C19447 _164_/Y VPWR 0.461f
C19448 _164_/A VGND 0.223f
C19449 _209_/X _332_/Q 0.00269f
C19450 _324_/a_761_249# _325_/D 1.43e-20
C19451 _340_/CLK _260_/a_27_257# 0.00102f
C19452 _329_/Q clkbuf_2_1_0_clk/A 0.0417f
C19453 _314_/a_1283_n19# _347_/a_651_373# 4.01e-20
C19454 _145_/A _306_/S 0.00891f
C19455 _293_/a_39_257# _313_/Q 0.0151f
C19456 _322_/a_193_7# _322_/a_1108_7# -0.00656f
C19457 clkbuf_0_clk/X _284_/A 0.408f
C19458 _263_/B _311_/a_193_7# 4.8e-21
C19459 _344_/a_1032_373# _161_/Y 0.00614f
C19460 _346_/D _347_/a_193_7# 3.03e-20
C19461 _304_/X _325_/D 0.251f
C19462 _279_/Y _300_/a_27_257# 4.07e-20
C19463 _343_/CLK _232_/A 1.83e-19
C19464 _292_/A _215_/A 1.68e-20
C19465 output14/a_27_7# _321_/Q 8.34e-19
C19466 _332_/a_639_7# _154_/A 8.34e-20
C19467 _192_/a_68_257# VGND 0.0267f
C19468 _341_/Q _204_/a_27_7# 4.61e-21
C19469 _330_/Q _181_/X 9.16e-19
C19470 _202_/a_250_257# _284_/A 0.00545f
C19471 _330_/D _330_/a_448_7# 0.00197f
C19472 _329_/a_651_373# _212_/X 1.11e-19
C19473 _277_/A _346_/SET_B 0.164f
C19474 _287_/a_39_257# _311_/a_1283_n19# 7.94e-22
C19475 _209_/a_27_257# _333_/Q 0.0465f
C19476 _209_/a_109_257# _332_/Q 0.00502f
C19477 _328_/a_193_7# clkbuf_2_1_0_clk/A 5.9e-21
C19478 _325_/a_543_7# _306_/S 2.36e-21
C19479 _185_/A _191_/B 4.63e-19
C19480 _339_/a_1283_n19# _283_/A 0.0649f
C19481 _346_/SET_B _336_/a_543_7# 0.00906f
C19482 _346_/a_796_7# _242_/A 1.3e-20
C19483 rstn _337_/a_1108_7# 1.14e-21
C19484 _210_/a_109_257# _207_/C 9.63e-21
C19485 _275_/Y _312_/a_805_7# 5.18e-19
C19486 _259_/a_199_7# VPWR -2.74e-19
C19487 _236_/B _243_/a_199_7# 6.36e-20
C19488 _196_/A VPWR 2.56f
C19489 _199_/a_346_7# _340_/CLK 5.03e-20
C19490 input1/X _284_/A 0.0103f
C19491 _345_/a_193_7# _165_/a_78_159# 0.0103f
C19492 _339_/D _194_/X 2.05e-20
C19493 _226_/a_79_n19# _298_/a_27_7# 7.06e-19
C19494 _269_/A _317_/a_193_7# 5.13e-20
C19495 _315_/a_193_7# _248_/A 0.0116f
C19496 _312_/D VGND 0.188f
C19497 _248_/A _298_/A 0.095f
C19498 _254_/Y _254_/a_109_257# 8.6e-19
C19499 rstn _343_/CLK 0.103f
C19500 _144_/A _283_/A 6.42e-20
C19501 _319_/a_639_7# _319_/D 9.32e-19
C19502 _181_/X _314_/D 0.00236f
C19503 _300_/Y _347_/a_761_249# 6.89e-19
C19504 _258_/a_439_7# _306_/X 0.00109f
C19505 _304_/a_257_159# VGND 0.102f
C19506 _316_/a_1283_n19# _318_/D 4.06e-21
C19507 _304_/a_591_329# VPWR -8.57e-19
C19508 _316_/D _315_/a_27_7# 3.86e-19
C19509 _324_/a_1283_n19# _216_/X 1.52e-20
C19510 _326_/a_1462_7# _326_/Q 1.17e-19
C19511 _283_/A _331_/a_27_7# 0.00155f
C19512 _256_/a_209_257# VGND -0.00111f
C19513 _256_/a_303_7# VPWR -6.83e-19
C19514 _279_/Y _324_/a_193_7# 0.00252f
C19515 repeater43/X _242_/A 0.404f
C19516 _177_/A VGND 1.01f
C19517 _227_/A _204_/a_277_7# 4.19e-19
C19518 _309_/a_193_7# _286_/B 2.14e-19
C19519 repeater43/X _335_/Q 0.057f
C19520 VPWR _298_/X 0.279f
C19521 _342_/Q _226_/X 1.57e-19
C19522 _318_/Q _232_/X 0.156f
C19523 _255_/a_30_13# clk 0.00301f
C19524 _279_/Y _314_/a_1270_373# 8.2e-20
C19525 clkbuf_2_0_0_clk/a_75_172# _338_/D 0.00927f
C19526 _313_/D _197_/X 2.28e-19
C19527 _258_/S _309_/Q 1.81e-20
C19528 _346_/a_476_7# _170_/a_76_159# 2.12e-20
C19529 output10/a_27_7# _340_/CLK 2.26e-20
C19530 _326_/a_1108_7# _242_/B 8.53e-22
C19531 _175_/Y _206_/A 1.45e-20
C19532 _144_/A _248_/B 0.0378f
C19533 _320_/a_193_7# ctlp[4] 4.21e-19
C19534 _260_/A _344_/D 8.89e-20
C19535 _284_/A _286_/Y 0.018f
C19536 _338_/Q _199_/a_250_257# 0.00484f
C19537 _254_/A _264_/a_113_257# 2.21e-19
C19538 _210_/a_307_257# _225_/X 3.29e-21
C19539 _333_/D VGND 0.25f
C19540 output20/a_27_7# _320_/Q 1.8e-21
C19541 _183_/a_553_257# _251_/X 1.22e-21
C19542 _324_/Q _251_/a_297_257# 0.00517f
C19543 _242_/A _319_/a_1462_7# 2.57e-19
C19544 _327_/a_543_7# _217_/A 3.71e-20
C19545 _329_/a_27_7# clkbuf_0_clk/X 0.0013f
C19546 _332_/a_193_7# VGND 0.00647f
C19547 _332_/a_543_7# VPWR 0.0103f
C19548 _217_/a_27_7# _283_/A 0.00926f
C19549 _334_/D _175_/Y 5.78e-21
C19550 _329_/Q _278_/a_68_257# 0.0238f
C19551 _320_/Q _278_/a_150_257# 2.2e-19
C19552 _347_/a_1283_n19# VPWR 0.0107f
C19553 _347_/a_761_249# VGND -0.00224f
C19554 _145_/A _283_/A 0.00738f
C19555 _326_/a_1283_n19# _304_/X 2.87e-19
C19556 _326_/a_193_7# _324_/D 1.93e-21
C19557 _285_/A output40/a_27_7# 0.0116f
C19558 _285_/A output32/a_27_7# 2.51e-20
C19559 repeater43/X _322_/D 0.00772f
C19560 _153_/A _333_/Q 0.705f
C19561 _334_/Q _335_/Q 0.794f
C19562 _325_/D VGND 0.158f
C19563 repeater43/X _321_/a_448_7# 0.00283f
C19564 _336_/a_1283_n19# _313_/a_193_7# 3.32e-21
C19565 _314_/Q _347_/a_193_7# 0.0109f
C19566 _297_/B _347_/a_448_7# 0.0167f
C19567 _314_/a_1108_7# _347_/D 9.04e-19
C19568 _250_/a_215_7# _284_/A 7.64e-19
C19569 _232_/X _241_/a_199_7# 6.35e-22
C19570 _234_/B _327_/Q 1.17e-19
C19571 _267_/B _310_/a_1283_n19# 1.94e-19
C19572 _306_/a_505_n19# _286_/B 0.0482f
C19573 _321_/a_1283_n19# _327_/Q 2.54e-20
C19574 _188_/a_76_159# _341_/Q 0.0174f
C19575 _258_/S _311_/a_193_7# 2.49e-19
C19576 _216_/X _218_/a_93_n19# 0.102f
C19577 _318_/Q _244_/B 1.65e-20
C19578 _320_/Q _279_/A 0.0306f
C19579 repeater43/X _153_/a_403_257# 2.69e-19
C19580 _306_/X _254_/B 4.8e-21
C19581 _165_/a_78_159# VPWR 0.0206f
C19582 _309_/D _264_/a_113_257# 0.00155f
C19583 _312_/Q _311_/a_1108_7# 0.0162f
C19584 _327_/a_193_7# _279_/A 2.36e-21
C19585 _191_/B _335_/Q 0.00248f
C19586 _328_/a_193_7# _278_/a_68_257# 2.05e-20
C19587 _175_/Y _147_/A 0.107f
C19588 _254_/A _336_/a_27_7# 4.88e-21
C19589 _145_/A _248_/B 1.44e-20
C19590 _341_/a_1283_n19# VGND 0.0156f
C19591 _341_/a_448_7# VPWR 0.00151f
C19592 _216_/X _220_/a_256_7# 2.97e-19
C19593 _327_/a_193_7# _218_/a_250_257# 1.26e-19
C19594 _324_/Q _306_/S 0.056f
C19595 _292_/A trimb[1] 4.11e-20
C19596 _294_/A _174_/a_27_257# 2.83e-20
C19597 _337_/Q _297_/Y 7.03e-20
C19598 _338_/a_448_7# VPWR -0.00338f
C19599 _338_/a_1283_n19# VGND 0.0836f
C19600 _323_/Q _298_/a_27_7# 5.11e-20
C19601 _178_/a_27_7# _298_/A 0.0248f
C19602 _149_/A _175_/Y 0.0613f
C19603 clkbuf_2_3_0_clk/A _265_/B 1.8e-20
C19604 _320_/Q _220_/a_346_7# 1.5e-20
C19605 _329_/Q _220_/a_256_7# 7.19e-19
C19606 _346_/a_1032_373# _277_/Y 8.04e-20
C19607 _326_/a_1283_n19# _272_/a_39_257# 0.00175f
C19608 _275_/Y _312_/Q 0.0251f
C19609 _308_/a_505_n19# _298_/C 6.85e-19
C19610 _328_/a_27_7# _279_/A 0.00816f
C19611 clkbuf_2_1_0_clk/A _337_/a_193_7# 2.28e-20
C19612 trim[3] VPWR 0.297f
C19613 _292_/A VGND 0.76f
C19614 _215_/A _190_/A 4.6e-19
C19615 _271_/A _316_/a_193_7# 0.00219f
C19616 _317_/Q _317_/a_651_373# 6.48e-19
C19617 _336_/a_543_7# _147_/A 5.76e-19
C19618 _290_/A _267_/A 0.0149f
C19619 clkbuf_2_0_0_clk/a_75_172# _343_/CLK 0.00348f
C19620 _340_/a_1270_373# VPWR -1.81e-20
C19621 _340_/a_448_7# VGND -0.00664f
C19622 _160_/A VGND 0.327f
C19623 _347_/Q _347_/D 3.63e-20
C19624 _337_/Q _310_/a_193_7# 0.00464f
C19625 _277_/Y _273_/A 0.00687f
C19626 _316_/D _242_/B 2.09e-20
C19627 input1/a_75_172# _283_/A 3.51e-19
C19628 _325_/Q _317_/a_1283_n19# 6.04e-20
C19629 cal _269_/A 0.0362f
C19630 _327_/a_651_373# _330_/Q 3.12e-19
C19631 _283_/A _331_/a_1217_7# 1.61e-19
C19632 _316_/a_651_373# VPWR 0.00185f
C19633 _345_/a_27_7# _346_/SET_B 0.0141f
C19634 _316_/a_1108_7# VGND 0.00814f
C19635 _343_/a_193_7# _248_/A 0.00153f
C19636 _344_/a_27_7# _164_/Y 1.02e-21
C19637 _344_/a_652_n19# _164_/A 2.32e-19
C19638 _300_/a_27_257# _313_/a_27_7# 3.92e-20
C19639 _341_/Q _206_/A 9.11e-19
C19640 _324_/a_761_249# _331_/CLK 0.00402f
C19641 _258_/S _309_/a_1108_7# 7.95e-20
C19642 _162_/X _171_/a_78_159# 0.0578f
C19643 _328_/a_761_249# _220_/a_250_257# 1.06e-19
C19644 _248_/A _304_/X 0.187f
C19645 _204_/a_27_257# VPWR 0.0653f
C19646 _238_/B VGND 0.242f
C19647 _326_/a_27_7# _271_/A 1.97e-21
C19648 _208_/a_493_257# VPWR -3.65e-19
C19649 _208_/a_78_159# VGND -0.0052f
C19650 _184_/a_76_159# _343_/Q 3.77e-19
C19651 _325_/a_805_7# _255_/B 2.63e-21
C19652 _209_/X _192_/B 6.75e-19
C19653 _327_/a_448_7# VPWR -0.00295f
C19654 _327_/a_1283_n19# VGND 0.00954f
C19655 _345_/a_1224_7# _292_/A 7.98e-20
C19656 _342_/a_761_249# _342_/D 0.0221f
C19657 _260_/A _340_/D 0.0105f
C19658 _346_/a_1182_221# _346_/D 1.96e-19
C19659 _331_/CLK _304_/X 0.132f
C19660 _254_/B _147_/Y 0.00868f
C19661 repeater43/X _315_/a_1108_7# -0.00152f
C19662 _273_/A _262_/a_199_7# 7.31e-19
C19663 _277_/Y _173_/a_556_7# 8.42e-19
C19664 _195_/a_27_257# _306_/S 0.0532f
C19665 _195_/a_109_257# _340_/Q 0.00294f
C19666 _195_/a_109_7# _194_/X 7.93e-19
C19667 _326_/a_448_7# VPWR -0.00257f
C19668 _326_/a_1283_n19# VGND 0.00519f
C19669 _322_/a_448_7# _322_/Q 2.11e-20
C19670 _343_/D cal 0.0345f
C19671 _328_/a_448_7# _330_/Q 2.77e-19
C19672 _318_/Q _241_/a_113_257# 0.053f
C19673 _345_/a_1032_373# _163_/a_78_159# 4.96e-19
C19674 _251_/a_297_257# _216_/A 1.4e-19
C19675 _339_/Q _297_/Y 8.16e-20
C19676 _273_/A _304_/X 0.0863f
C19677 _169_/Y _254_/A 0.00868f
C19678 _329_/a_1217_7# clkbuf_0_clk/X 1.88e-19
C19679 _346_/a_1224_7# clkbuf_2_1_0_clk/A 7.32e-19
C19680 _332_/a_1462_7# VGND 2.38e-19
C19681 _306_/S _228_/A 0.00692f
C19682 _328_/a_543_7# VGND 0.0115f
C19683 _328_/a_1108_7# VPWR 0.0133f
C19684 _344_/a_193_7# _286_/B 7.88e-20
C19685 _307_/a_505_n19# _215_/A 2.98e-20
C19686 _191_/B _209_/a_373_7# 5.66e-20
C19687 _191_/B _336_/Q 7.86e-19
C19688 _255_/X cal 2.83e-19
C19689 _342_/Q input1/X 0.00648f
C19690 _321_/a_1108_7# result[7] 3.22e-19
C19691 _297_/B _347_/D 0.0453f
C19692 _164_/Y _171_/a_215_7# 0.0081f
C19693 _272_/a_39_257# _248_/A 0.013f
C19694 result[6] _242_/A 1.12e-20
C19695 _341_/Q _147_/A 0.0908f
C19696 _339_/Q _310_/a_193_7# 8.78e-20
C19697 _346_/a_1602_7# _160_/X 0.00147f
C19698 _258_/a_535_334# _286_/B 2.57e-19
C19699 _165_/X _344_/D 3.51e-20
C19700 clkbuf_2_3_0_clk/A clkbuf_2_1_0_clk/A 0.472f
C19701 _334_/a_543_7# VGND -0.00248f
C19702 _334_/a_1108_7# VPWR 0.0206f
C19703 _215_/A _178_/a_27_7# 0.00205f
C19704 _163_/a_215_7# _160_/X 3.42e-19
C19705 _172_/Y _170_/a_76_159# 2.9e-20
C19706 _296_/a_295_257# _284_/A 8.11e-19
C19707 _341_/Q _149_/A 0.0232f
C19708 cal _210_/a_109_257# 0.00223f
C19709 _172_/A _286_/B 1.07f
C19710 _324_/Q _283_/A 0.0743f
C19711 _296_/Y _298_/A 1.46e-21
C19712 _330_/Q _346_/SET_B 0.0248f
C19713 _307_/a_439_7# _227_/A 3.59e-19
C19714 _165_/X _346_/Q 0.521f
C19715 _341_/D VPWR 0.136f
C19716 _216_/X _328_/D 0.14f
C19717 _304_/S _227_/A 0.574f
C19718 _327_/a_27_7# _330_/D 0.00177f
C19719 _216_/A _306_/S 0.0102f
C19720 _286_/B _198_/a_250_257# 2.77e-19
C19721 _273_/A _272_/a_39_257# 0.00108f
C19722 _273_/A _300_/Y 1.8e-20
C19723 _323_/a_761_249# _298_/C 0.00205f
C19724 _323_/a_1283_n19# _343_/Q 0.00157f
C19725 _294_/Y _344_/Q 1.52e-19
C19726 _188_/S _181_/X 0.156f
C19727 _146_/a_29_271# _298_/A 4.43e-19
C19728 clkbuf_2_1_0_clk/A _172_/Y 2.15e-20
C19729 _338_/D VPWR 0.295f
C19730 _168_/a_481_7# _165_/X 2.54e-19
C19731 _172_/A _304_/a_306_329# 4.7e-21
C19732 ctln[3] trim[3] 0.0032f
C19733 _329_/Q _328_/D 0.0864f
C19734 _316_/Q _316_/a_805_7# 0.00228f
C19735 _298_/B _144_/A 7.96e-22
C19736 _281_/A _327_/D 1.48e-20
C19737 _329_/a_1108_7# _281_/A 0.00808f
C19738 _325_/a_805_7# _325_/Q 1.81e-20
C19739 _277_/Y _267_/a_109_257# 2.38e-19
C19740 result[6] _322_/D 0.0109f
C19741 _329_/a_761_249# _281_/Y 0.00555f
C19742 _346_/SET_B _314_/D 0.00444f
C19743 _342_/a_543_7# _177_/a_27_7# 0.00943f
C19744 _317_/a_1283_n19# _326_/Q 2.32e-19
C19745 _342_/Q _286_/Y 0.306f
C19746 _227_/A _225_/X 0.00712f
C19747 _321_/D _321_/Q 0.141f
C19748 _324_/Q _248_/B 0.139f
C19749 _307_/X _227_/A 1.73e-19
C19750 _293_/a_121_257# _194_/A 8.71e-20
C19751 _342_/a_193_7# output41/a_27_7# 4.39e-20
C19752 _248_/A VGND 1.73f
C19753 _346_/a_381_7# VPWR 0.00144f
C19754 _346_/a_1032_373# VGND 0.0321f
C19755 _337_/Q _310_/a_1462_7# 4.75e-20
C19756 _337_/Q _199_/a_93_n19# 2.39e-19
C19757 _233_/a_113_257# _322_/Q 0.00101f
C19758 _333_/a_27_7# _333_/a_761_249# -0.0173f
C19759 _335_/a_1108_7# _204_/a_27_257# 4.39e-20
C19760 output11/a_27_7# _153_/B 4.18e-19
C19761 _163_/a_493_257# VGND -2.6e-19
C19762 _335_/a_1283_n19# _208_/a_215_7# 2.82e-19
C19763 _236_/B VPWR 0.548f
C19764 _329_/a_543_7# _319_/Q 0.0299f
C19765 _273_/A trimb[1] 8.63e-19
C19766 _331_/CLK VGND 2.13f
C19767 _318_/a_1108_7# _248_/A 0.00159f
C19768 _345_/a_586_7# _346_/SET_B 4.73e-19
C19769 _344_/a_1056_7# _164_/A 0.00127f
C19770 _299_/X _313_/a_1283_n19# 4.36e-21
C19771 _347_/Q _313_/a_543_7# 3.46e-21
C19772 _267_/A _310_/a_27_7# 2.93e-20
C19773 _340_/CLK _311_/a_1108_7# 8.25e-20
C19774 _162_/X _172_/B 0.0333f
C19775 _328_/a_193_7# _328_/D -0.01f
C19776 _190_/A VGND 1.23f
C19777 _323_/Q _154_/A 9.71e-20
C19778 _329_/a_761_249# _329_/D 0.043f
C19779 _283_/A _195_/a_27_257# 2.95e-21
C19780 _283_/Y _338_/a_27_7# 5.97e-19
C19781 _321_/D _318_/a_193_7# 0.00921f
C19782 _326_/a_27_7# _232_/a_27_7# 2.01e-21
C19783 _236_/B _318_/a_543_7# 1.23e-19
C19784 _286_/B _203_/a_80_n19# 3.17e-19
C19785 _283_/A _281_/A 0.0204f
C19786 _318_/a_1108_7# _331_/CLK 1.37e-21
C19787 _273_/Y VPWR 0.0458f
C19788 _337_/Q _336_/Q 0.0175f
C19789 _336_/a_193_7# _202_/a_93_n19# 3.02e-19
C19790 _336_/a_27_7# _202_/a_250_257# 5.06e-20
C19791 _273_/A VGND 1.52f
C19792 _294_/A _216_/A 1.46e-19
C19793 _219_/a_256_7# _319_/D 3.04e-21
C19794 _143_/a_27_7# VPWR 0.0596f
C19795 _294_/Y output33/a_27_7# 9.71e-19
C19796 _340_/Q _340_/D 3.85e-19
C19797 _326_/D VPWR 0.128f
C19798 repeater43/X _324_/a_448_7# -2.34e-19
C19799 _145_/A _298_/B 0.0373f
C19800 _283_/A _228_/A 0.00779f
C19801 _275_/Y _340_/CLK 0.169f
C19802 cal _336_/a_193_7# 5.46e-21
C19803 input1/X _336_/a_27_7# 0.618f
C19804 _345_/a_1602_7# _158_/Y 1.82e-19
C19805 _305_/a_505_n19# _194_/A 0.0313f
C19806 output17/a_27_7# ctlp[4] 2.93e-20
C19807 ctlp[3] output18/a_27_7# 1.62e-19
C19808 _222_/a_256_7# VPWR -7.99e-19
C19809 _222_/a_93_n19# VGND -0.0042f
C19810 _332_/a_639_7# _153_/B 0.00121f
C19811 _324_/a_1283_n19# _327_/Q 3.96e-20
C19812 _255_/X _284_/A 1.61e-20
C19813 _343_/a_1108_7# repeater43/X 0.00781f
C19814 _329_/a_27_7# _329_/a_193_7# -0.296f
C19815 _173_/a_556_7# VGND 6.39e-19
C19816 _221_/a_584_7# _327_/D 5.27e-20
C19817 _284_/A clkc 1.13e-20
C19818 _296_/Y _215_/A 0.0067f
C19819 _206_/A _269_/Y 4.61e-20
C19820 _271_/A _334_/a_805_7# 1.32e-19
C19821 _319_/a_651_373# VPWR 1.79e-19
C19822 _319_/a_1108_7# VGND -0.00595f
C19823 _313_/a_193_7# VPWR -0.308f
C19824 _337_/a_1108_7# VPWR -0.00194f
C19825 _337_/a_543_7# VGND -0.00365f
C19826 _346_/SET_B _311_/a_448_7# 1.7e-19
C19827 trim[4] VGND 0.274f
C19828 _301_/a_245_257# _344_/D 1.55e-20
C19829 _183_/a_1241_257# _341_/Q 2.36e-19
C19830 _304_/X _217_/X 0.0514f
C19831 _217_/A _212_/X 0.0811f
C19832 _342_/a_761_249# _341_/a_193_7# 1.69e-20
C19833 _342_/a_27_7# _341_/a_543_7# 6.7e-21
C19834 _342_/a_193_7# _341_/a_761_249# 2.39e-20
C19835 _342_/a_543_7# _341_/a_27_7# 2.76e-20
C19836 output27/a_27_7# _331_/CLK 0.0604f
C19837 _339_/Q _199_/a_93_n19# 0.0586f
C19838 _297_/B _313_/a_543_7# 3.69e-20
C19839 _306_/X _196_/A 1.62e-20
C19840 _217_/a_27_7# _242_/B 3.09e-20
C19841 _308_/S _295_/a_79_n19# 0.0358f
C19842 _320_/Q _322_/a_193_7# 0.457f
C19843 _248_/B _228_/A 0.101f
C19844 _343_/CLK VPWR 3.75f
C19845 clkbuf_0_clk/X _225_/B 0.00486f
C19846 _320_/Q _320_/a_1270_373# 6.38e-20
C19847 _238_/B _320_/a_1108_7# 1.21e-19
C19848 _254_/A _315_/D 2.53e-20
C19849 _216_/A _283_/A 0.792f
C19850 _179_/a_27_7# _298_/C 0.00349f
C19851 _345_/a_956_373# _345_/Q 6.89e-19
C19852 _345_/a_562_373# _345_/D 4.93e-19
C19853 _307_/a_535_334# VPWR 1.11e-19
C19854 _307_/a_505_n19# VGND 0.0645f
C19855 result[4] _242_/A 0.00508f
C19856 _167_/X _167_/a_27_257# 0.00107f
C19857 clkbuf_0_clk/a_110_7# _215_/A 0.0638f
C19858 _343_/a_805_7# _343_/CLK 7.8e-21
C19859 _145_/a_113_7# VGND 3.99e-20
C19860 rstn _195_/a_109_257# 0.00297f
C19861 _339_/Q _336_/Q 0.0689f
C19862 _325_/a_805_7# _326_/Q 2.11e-19
C19863 _324_/a_639_7# _304_/S 0.00431f
C19864 _309_/a_761_249# trim[4] 2.67e-20
C19865 input1/X _199_/a_250_257# 0.00574f
C19866 _164_/Y _147_/Y 1.26e-21
C19867 _178_/a_27_7# VGND 0.0389f
C19868 _178_/a_193_257# VPWR -3.12e-19
C19869 _304_/S _297_/B 0.00244f
C19870 _296_/Y _304_/X 4.53e-21
C19871 _279_/Y _172_/A 0.0101f
C19872 _188_/S _229_/a_76_159# 8.31e-21
C19873 _324_/Q _315_/a_27_7# 1.76e-19
C19874 _340_/a_193_7# _197_/X 0.00685f
C19875 _320_/Q _246_/a_109_257# 0.00355f
C19876 _183_/a_27_7# _227_/A 0.00298f
C19877 _218_/a_93_n19# _327_/Q 0.00121f
C19878 _343_/a_1283_n19# _323_/Q 0.00149f
C19879 _272_/a_121_257# _212_/X 8.18e-22
C19880 _279_/Y _211_/a_109_257# 1.04e-19
C19881 clkbuf_2_3_0_clk/A _311_/a_27_7# 3.66e-20
C19882 _328_/a_1283_n19# _320_/a_1283_n19# 0.00378f
C19883 _302_/a_77_159# _299_/X 2.14e-21
C19884 clk _227_/A 0.0132f
C19885 _216_/A _248_/B 0.262f
C19886 _279_/Y _232_/X 0.00117f
C19887 input1/X _225_/B 0.77f
C19888 _325_/a_193_7# _324_/a_543_7# 5.95e-19
C19889 _325_/a_27_7# _324_/a_1283_n19# 0.00228f
C19890 _174_/a_109_257# _310_/D 1.63e-19
C19891 _157_/A _314_/a_27_7# 3.56e-19
C19892 _255_/a_112_257# _255_/B 2.75e-19
C19893 clkbuf_0_clk/X _314_/a_543_7# 0.00246f
C19894 _309_/a_805_7# _346_/SET_B -8.28e-19
C19895 _207_/a_27_7# _153_/a_109_53# 7.76e-21
C19896 _267_/a_109_257# VGND -7.81e-19
C19897 _335_/a_805_7# _207_/X 4.25e-19
C19898 _339_/a_1108_7# VPWR 0.0126f
C19899 _339_/a_543_7# VGND -0.00654f
C19900 result[4] _322_/D 0.013f
C19901 _217_/X _220_/a_93_n19# 0.0078f
C19902 _212_/X _220_/a_250_257# 5.12e-19
C19903 _341_/a_1108_7# _244_/B 0.0051f
C19904 _341_/a_543_7# _317_/D 0.00276f
C19905 _263_/a_109_257# _263_/B 0.00178f
C19906 _327_/a_1108_7# _232_/X 0.00848f
C19907 _258_/a_76_159# _340_/CLK 0.00368f
C19908 _341_/Q _150_/a_27_7# 0.0051f
C19909 _325_/a_193_7# _217_/A 0.192f
C19910 _325_/a_761_249# _304_/X 0.0221f
C19911 _207_/X _153_/B 0.00231f
C19912 input4/X _271_/Y 0.0168f
C19913 repeater43/X _271_/A 0.183f
C19914 _283_/Y _338_/a_1217_7# 7.28e-20
C19915 _254_/Y _216_/A 7.5e-20
C19916 _326_/a_1108_7# _232_/X 0.00356f
C19917 _196_/A _147_/Y 0.0159f
C19918 _294_/A _294_/Y 0.572f
C19919 input4/X _335_/a_761_249# 2.15e-19
C19920 repeater43/X _335_/a_27_7# -0.00131f
C19921 _336_/a_193_7# _284_/A 0.00465f
C19922 _330_/Q _331_/a_761_249# 0.00808f
C19923 trim[2] clkc 0.128f
C19924 _329_/D _319_/D 1.08e-21
C19925 _318_/a_27_7# _317_/a_193_7# 4.89e-19
C19926 _318_/a_193_7# _317_/a_27_7# 8.46e-19
C19927 _169_/B _267_/A 0.00403f
C19928 _312_/a_543_7# _312_/Q 0.0018f
C19929 _265_/a_109_257# _265_/B 4.68e-19
C19930 _331_/a_193_7# VPWR 0.0251f
C19931 output29/a_27_7# VPWR 0.0986f
C19932 _200_/a_256_7# _197_/X 0.00215f
C19933 _320_/a_761_249# _346_/SET_B 0.00195f
C19934 _271_/Y _207_/C 0.0271f
C19935 _340_/a_1108_7# _254_/B 6.06e-21
C19936 _217_/X VGND 0.428f
C19937 _288_/A trimb[4] 2.44e-19
C19938 _288_/A trim[1] 0.00431f
C19939 _335_/a_1283_n19# _206_/A 0.00139f
C19940 _335_/a_761_249# _207_/C 7.65e-21
C19941 repeater43/X _318_/a_639_7# 0.00386f
C19942 _260_/B _254_/B 0.0119f
C19943 _316_/a_448_7# _244_/B 0.00899f
C19944 _290_/A _310_/a_1108_7# 0.0158f
C19945 _260_/A _314_/a_27_7# 1.8e-20
C19946 _271_/A _334_/Q 0.0105f
C19947 _313_/a_805_7# VGND -4.6e-19
C19948 _246_/B _150_/C 5.21e-21
C19949 _346_/SET_B _311_/D 0.00458f
C19950 _258_/a_505_n19# _346_/SET_B 0.00399f
C19951 _324_/Q _298_/B 0.00287f
C19952 _335_/D _334_/a_1283_n19# 2.18e-19
C19953 _335_/a_1108_7# _343_/CLK 0.0047f
C19954 _335_/a_27_7# _334_/Q 0.00159f
C19955 _315_/a_27_7# _228_/A 0.009f
C19956 ctln[3] _343_/CLK 8.64e-21
C19957 _308_/a_505_n19# _150_/C 2.7e-20
C19958 output15/a_27_7# _331_/Q 4.11e-19
C19959 _342_/Q _269_/A 1.3e-20
C19960 _277_/A _319_/Q 0.198f
C19961 _167_/a_27_257# _301_/a_51_257# 8.04e-20
C19962 _344_/a_1182_221# _163_/a_78_159# 1.58e-19
C19963 _214_/a_27_257# _331_/CLK 5.4e-19
C19964 _247_/a_113_257# _232_/A 0.0089f
C19965 _271_/A _191_/B 0.0116f
C19966 _296_/Y VGND 0.0939f
C19967 _317_/a_193_7# _246_/B 1.14e-19
C19968 _318_/Q _316_/a_1108_7# 3.16e-19
C19969 _147_/Y _347_/a_1283_n19# 2.74e-19
C19970 _315_/Q _317_/D 0.0121f
C19971 result[0] _244_/B 2.41e-19
C19972 rstn _340_/D 0.281f
C19973 clkbuf_2_1_0_clk/A _260_/A 0.00794f
C19974 _320_/Q _330_/a_543_7# 0.0296f
C19975 _286_/B _164_/A 1.53e-20
C19976 _267_/B _311_/a_1108_7# 7.04e-19
C19977 _342_/a_1108_7# _229_/a_489_373# 2.28e-19
C19978 _327_/a_543_7# _331_/D 4.95e-20
C19979 _273_/A _214_/a_27_257# 3.02e-21
C19980 _326_/Q _221_/a_93_n19# 3.47e-19
C19981 _146_/a_29_271# VGND 0.0134f
C19982 _146_/a_184_13# VPWR -2.14e-19
C19983 repeater43/X _323_/a_27_7# 0.0171f
C19984 _184_/a_76_159# _147_/A 0.0151f
C19985 _327_/a_1283_n19# _318_/Q 0.00315f
C19986 repeater43/X _330_/D 0.00459f
C19987 _336_/Q _336_/D 1.55e-20
C19988 _192_/a_68_257# _192_/a_150_257# 8.88e-34
C19989 _188_/a_76_159# _188_/S 3.99e-19
C19990 clkbuf_0_clk/X _315_/D 0.00619f
C19991 _183_/a_553_257# VPWR 0.00369f
C19992 _316_/Q _317_/a_193_7# 1.27e-19
C19993 _326_/a_1283_n19# _318_/Q 2.76e-20
C19994 _324_/a_193_7# _324_/Q 0.00337f
C19995 _324_/a_1283_n19# _157_/A 8.86e-22
C19996 clkbuf_0_clk/a_110_7# VGND 0.0925f
C19997 _301_/X _347_/Q 0.0324f
C19998 _342_/D valid 0.00306f
C19999 _328_/a_1283_n19# _320_/D 1.62e-20
C20000 _325_/a_761_249# VGND 0.00265f
C20001 _325_/a_1283_n19# VPWR 0.0475f
C20002 _275_/Y _267_/B 0.00714f
C20003 _263_/a_109_257# _194_/A 1.29e-19
C20004 _232_/X _316_/D 0.0763f
C20005 _344_/D _310_/D 1.24e-19
C20006 clkbuf_2_1_0_clk/A _261_/A 6.98e-22
C20007 _271_/A _317_/a_543_7# 4.45e-19
C20008 _333_/a_651_373# _333_/D 0.00247f
C20009 _323_/a_1283_n19# _206_/A 1.95e-21
C20010 _323_/a_761_249# _207_/C 3.56e-21
C20011 _286_/B _192_/a_68_257# 0.0586f
C20012 _340_/Q _265_/B 2.45e-21
C20013 _342_/Q _255_/X 0.0174f
C20014 _207_/a_27_7# _153_/A 1.75e-19
C20015 _339_/a_27_7# _153_/B 1.22e-19
C20016 _257_/a_544_257# _255_/X 4.62e-21
C20017 _327_/Q _328_/D 2.92e-20
C20018 _261_/A _310_/Q 8.23e-20
C20019 _306_/S _209_/a_27_257# 0.0616f
C20020 _333_/a_1283_n19# _332_/a_1283_n19# 3.64e-19
C20021 _317_/a_639_7# VPWR 5.61e-19
C20022 _317_/a_651_373# VGND 0.00264f
C20023 _323_/a_1108_7# _343_/CLK 2.92e-19
C20024 _263_/B _312_/Q 0.00249f
C20025 _297_/A _347_/a_543_7# 0.0395f
C20026 _298_/B _228_/A 2.3e-19
C20027 repeater43/X _232_/a_27_7# 0.0221f
C20028 _336_/a_1462_7# _284_/A 2.71e-19
C20029 _259_/a_113_257# _312_/D 2.14e-21
C20030 _258_/a_505_n19# _313_/a_761_249# 0.00337f
C20031 _337_/Q _311_/a_761_249# 3e-20
C20032 _292_/A _312_/a_651_373# 5.85e-19
C20033 _232_/X _222_/a_250_257# 3.32e-21
C20034 _314_/a_1283_n19# _284_/A 7.74e-21
C20035 _172_/A _313_/a_27_7# 2.04e-20
C20036 _276_/a_68_257# VPWR 0.029f
C20037 _290_/A _291_/a_121_257# 7.04e-19
C20038 _321_/Q _280_/a_68_257# 0.00631f
C20039 _331_/a_805_7# VGND 3.11e-19
C20040 _331_/a_1462_7# VPWR 2.07e-19
C20041 _304_/a_257_159# _286_/B 4.05e-19
C20042 _310_/a_1283_n19# _297_/Y 0.00305f
C20043 _320_/Q _331_/Q 0.0208f
C20044 _169_/B _167_/X 0.0865f
C20045 _256_/a_80_n19# _196_/A 0.0376f
C20046 _344_/a_1140_373# _346_/SET_B -6.31e-19
C20047 _316_/D _244_/B 0.0129f
C20048 _343_/a_651_373# cal 0.00195f
C20049 _337_/a_1108_7# _198_/a_93_n19# 3.97e-19
C20050 _190_/A _203_/a_209_257# 0.00593f
C20051 _254_/B _333_/Q 8.37e-19
C20052 _301_/X _297_/B 0.692f
C20053 _281_/Y _227_/A 0.0447f
C20054 _345_/Q _171_/a_78_159# 2.82e-21
C20055 _172_/A _307_/a_218_334# 0.00171f
C20056 output31/a_27_7# _297_/Y 0.00154f
C20057 _323_/a_193_7# _226_/X 1.04e-21
C20058 _326_/a_193_7# _331_/Q 9.15e-21
C20059 _174_/a_109_257# VPWR 0.00721f
C20060 _313_/Q _346_/SET_B 0.0123f
C20061 _322_/a_1108_7# _321_/D 0.00253f
C20062 _271_/A result[6] 2.02e-20
C20063 _323_/a_1283_n19# _149_/A 0.00149f
C20064 _248_/A _330_/a_27_7# 2.21e-19
C20065 _324_/a_193_7# _228_/A 0.192f
C20066 _234_/B _230_/a_27_7# 3.33e-20
C20067 _286_/B _333_/D 3.71e-19
C20068 _318_/Q _248_/A 0.0103f
C20069 _344_/a_1032_373# _158_/Y 0.00357f
C20070 ctln[7] input4/X 0.0322f
C20071 _283_/Y repeater43/X 4.65e-19
C20072 _258_/a_505_n19# _147_/A 1.75e-19
C20073 _283_/A _153_/a_109_53# 2.21e-19
C20074 _315_/D _286_/Y 0.0393f
C20075 _196_/A _332_/a_27_7# 3.49e-21
C20076 _197_/X _338_/Q 0.0231f
C20077 _331_/CLK _330_/a_27_7# 0.18f
C20078 VPWR output30/a_27_7# 0.107f
C20079 _196_/A _347_/a_193_7# 3.71e-19
C20080 _186_/a_297_7# _150_/C 7.06e-19
C20081 _308_/X _226_/a_297_7# 1.8e-19
C20082 _324_/a_651_373# _286_/Y 0.00109f
C20083 _184_/a_439_7# _192_/B 6.44e-20
C20084 _318_/Q _331_/CLK 0.313f
C20085 _340_/CLK _312_/a_543_7# 1.66e-19
C20086 _219_/a_93_n19# VPWR 0.0233f
C20087 _309_/a_193_7# _174_/a_27_257# 1.24e-20
C20088 _306_/S _153_/A 0.472f
C20089 repeater43/X _322_/a_761_249# 3.39e-20
C20090 _342_/a_805_7# _248_/A 4.44e-19
C20091 _342_/D _229_/a_226_7# 3.02e-20
C20092 _345_/a_193_7# _344_/D 1.61e-20
C20093 _286_/B _325_/D 6.5e-23
C20094 _299_/X _284_/A 2.53e-19
C20095 _339_/Q _311_/a_761_249# 7.15e-21
C20096 _343_/Q output41/a_27_7# 0.00114f
C20097 _176_/a_27_7# _298_/X 0.038f
C20098 _234_/B _232_/A 2.17e-20
C20099 clkbuf_2_1_0_clk/A _340_/Q 0.103f
C20100 _154_/a_27_7# _207_/C 5.54e-21
C20101 result[6] _318_/a_639_7# 6.41e-20
C20102 repeater43/X _323_/a_1217_7# 2.37e-19
C20103 _255_/X _336_/a_27_7# 1.37e-21
C20104 _321_/a_1283_n19# _232_/A 3.26e-21
C20105 _279_/Y _297_/A 0.0211f
C20106 ctln[7] _207_/C 1.18e-20
C20107 clk _335_/a_543_7# 9.36e-20
C20108 _188_/S _147_/A 0.0466f
C20109 _273_/A _318_/Q 6.58e-19
C20110 _345_/a_193_7# _346_/Q 1.3e-19
C20111 _330_/D _331_/a_448_7# 1.1e-19
C20112 _320_/a_1108_7# _217_/X 6.88e-20
C20113 _308_/a_505_n19# cal 8.22e-22
C20114 _308_/a_76_159# input1/X 0.0484f
C20115 _242_/A _319_/D 0.0346f
C20116 _167_/X _170_/a_226_7# 0.00191f
C20117 _324_/a_193_7# _216_/A 6.64e-19
C20118 _214_/a_109_7# _327_/Q 2.27e-19
C20119 _214_/a_27_257# _217_/X 3.07e-20
C20120 _214_/a_109_257# _212_/X 0.00559f
C20121 _188_/S _149_/A 0.00168f
C20122 _321_/a_27_7# _234_/B 5.09e-20
C20123 _309_/Q _267_/A 1.23e-19
C20124 output18/a_27_7# _346_/SET_B 5.4e-20
C20125 _283_/Y _334_/Q 3.15e-20
C20126 _321_/a_193_7# _321_/a_543_7# -0.0102f
C20127 _268_/a_39_257# _316_/a_27_7# 0.00547f
C20128 _172_/A _144_/A 4.53e-21
C20129 _324_/a_1283_n19# _251_/a_79_n19# 1.01e-20
C20130 _165_/a_215_7# trimb[4] 3.56e-19
C20131 output38/a_27_7# _285_/Y 4.43e-20
C20132 _165_/X clkbuf_2_1_0_clk/A 0.0207f
C20133 _342_/a_543_7# repeater43/X 4.36e-19
C20134 _251_/X _314_/a_27_7# 0.00727f
C20135 _338_/Q _312_/a_193_7# 2.28e-20
C20136 _346_/SET_B _312_/a_1283_n19# -8.97e-19
C20137 _324_/D _221_/a_93_n19# 3.06e-20
C20138 _166_/Y _347_/Q 1.49e-20
C20139 _332_/a_193_7# _332_/a_761_249# -0.00395f
C20140 _279_/Y _192_/a_68_257# 0.00193f
C20141 _306_/X _313_/a_193_7# 2.3e-20
C20142 _313_/Q _313_/a_761_249# 4.37e-20
C20143 _258_/S _312_/Q 0.503f
C20144 _340_/a_27_7# _338_/a_27_7# 1.55e-21
C20145 _291_/a_39_257# _297_/Y 7.76e-19
C20146 _232_/X _331_/a_27_7# 0.00342f
C20147 _345_/a_27_7# _290_/A 0.00805f
C20148 rstn _153_/a_215_257# 1.5e-20
C20149 _337_/D _311_/D 5.87e-21
C20150 _341_/a_1108_7# _177_/A 2.29e-20
C20151 _277_/Y _193_/Y 5.71e-21
C20152 ctln[4] _340_/Q 2.15e-20
C20153 _169_/B _301_/a_51_257# 1.58e-20
C20154 _341_/a_193_7# valid 3.89e-20
C20155 _236_/B _233_/a_199_7# 9.95e-19
C20156 _168_/a_397_257# _160_/X 6.72e-20
C20157 _325_/Q _243_/a_113_257# 0.00189f
C20158 _216_/X _181_/X 0.00938f
C20159 _261_/A _311_/a_27_7# 0.00997f
C20160 _267_/A _311_/a_193_7# 0.0244f
C20161 _175_/Y _298_/a_27_7# 4.23e-20
C20162 en _269_/A 0.0304f
C20163 _289_/a_39_257# _338_/Q 0.0504f
C20164 output14/a_27_7# _320_/Q 5.61e-19
C20165 output24/a_27_7# _315_/a_1108_7# 5.54e-22
C20166 _260_/B _196_/A 0.923f
C20167 _313_/D _254_/A 9.18e-22
C20168 _305_/a_76_159# _192_/B 7.06e-21
C20169 _195_/a_109_257# VPWR 0.00116f
C20170 _255_/B _341_/Q 0.0496f
C20171 ctlp[5] _217_/X 1.61e-20
C20172 output12/a_27_7# VGND 0.128f
C20173 _345_/Q _172_/B 0.019f
C20174 _346_/a_193_7# _162_/X 1.05e-19
C20175 _172_/A _145_/A 0.304f
C20176 _255_/X _225_/B 0.00763f
C20177 _323_/a_543_7# clk 7.98e-19
C20178 _281_/Y _324_/a_639_7# 6.89e-19
C20179 _344_/D VPWR 0.273f
C20180 _283_/A _224_/a_93_n19# 0.00697f
C20181 _294_/Y _284_/a_39_257# 0.00799f
C20182 _216_/A _160_/X 2.04e-20
C20183 _257_/a_448_7# _225_/B 0.0102f
C20184 _319_/Q _330_/Q 0.0246f
C20185 _275_/Y _261_/a_109_257# 0.0013f
C20186 output9/a_27_7# _267_/A 1.3e-19
C20187 _217_/a_27_7# _232_/X 0.00928f
C20188 _325_/a_761_249# _214_/a_27_257# 1.06e-20
C20189 _279_/Y _256_/a_209_257# 5.04e-20
C20190 _326_/a_761_249# _181_/X 3.56e-19
C20191 _343_/D en 4.29e-19
C20192 _185_/A _227_/A 0.00533f
C20193 _281_/Y _297_/B 3.8e-19
C20194 _200_/a_93_n19# _194_/A 0.00972f
C20195 _254_/A _197_/X 3.87e-22
C20196 _346_/Q VPWR 0.217f
C20197 _273_/A output40/a_27_7# 0.00294f
C20198 _232_/A _315_/a_543_7# 6.56e-20
C20199 output32/a_27_7# _273_/A 0.0135f
C20200 _336_/a_27_7# _336_/a_193_7# -0.33f
C20201 _340_/CLK _263_/B 0.0109f
C20202 _313_/Q _147_/A 0.0617f
C20203 _283_/A _153_/A 0.0276f
C20204 _237_/a_113_257# _329_/Q 0.00125f
C20205 _237_/a_199_7# _320_/Q 1.89e-19
C20206 _331_/CLK _330_/a_1217_7# 1.82e-21
C20207 _166_/Y _297_/B 0.0644f
C20208 _168_/a_481_7# VPWR -4.36e-19
C20209 _168_/a_109_257# VGND -0.00137f
C20210 _207_/a_109_7# VGND 0.00104f
C20211 _309_/a_27_7# _344_/D 1.95e-19
C20212 _342_/a_1283_n19# _226_/X 3.45e-21
C20213 _346_/a_476_7# _299_/a_78_159# 0.00875f
C20214 _322_/a_193_7# result[7] 7.86e-20
C20215 output25/a_27_7# _317_/a_27_7# 4.09e-21
C20216 _313_/a_193_7# _147_/Y 1.58e-19
C20217 _301_/a_51_257# _170_/a_226_7# 2.83e-19
C20218 _188_/S _183_/a_1241_257# 0.0168f
C20219 _333_/a_651_373# _190_/A 6.05e-19
C20220 _323_/a_761_249# cal 0.00365f
C20221 _329_/D _297_/B 0.216f
C20222 _254_/Y _336_/a_651_373# 0.0265f
C20223 _309_/a_1108_7# _267_/A 4.62e-20
C20224 _341_/a_27_7# _341_/a_639_7# -0.0015f
C20225 _279_/Y _332_/a_193_7# 1.86e-19
C20226 _345_/a_27_7# _167_/a_27_257# 5.01e-20
C20227 _162_/X _173_/a_76_159# 3.69e-19
C20228 repeater43/X _330_/a_1283_n19# 0.00442f
C20229 _308_/S input1/X 0.283f
C20230 output32/a_27_7# trim[4] 0.00124f
C20231 _294_/Y _262_/a_113_257# 0.00788f
C20232 _164_/A _163_/a_215_7# 0.00176f
C20233 _332_/a_193_7# _208_/a_292_257# 6.84e-21
C20234 _331_/D _212_/X 0.119f
C20235 _314_/a_1108_7# _297_/Y 2.18e-19
C20236 _197_/X _339_/a_639_7# 9.22e-20
C20237 _315_/D _328_/Q 3.88e-19
C20238 _330_/a_193_7# _212_/X 5.87e-20
C20239 clkbuf_2_1_0_clk/A _301_/a_245_257# 0.00134f
C20240 _251_/a_215_7# VGND -0.0174f
C20241 repeater43/X _333_/a_27_7# 0.00601f
C20242 _221_/a_346_7# VGND -0.00195f
C20243 _338_/a_27_7# _338_/a_639_7# -0.00188f
C20244 _338_/a_1283_n19# _338_/a_1108_7# -2.84e-32
C20245 _318_/Q _217_/X 0.0441f
C20246 _145_/A _244_/B 0.112f
C20247 _324_/a_1283_n19# _296_/a_213_83# 1.29e-20
C20248 _344_/a_193_7# _174_/a_27_257# 4.49e-20
C20249 _325_/Q _341_/Q 7.55e-20
C20250 _192_/B _203_/a_303_7# 5.7e-19
C20251 _319_/Q clkbuf_2_1_0_clk/a_75_172# 2.49e-19
C20252 _194_/X _311_/a_193_7# 1.34e-20
C20253 _243_/a_113_257# _326_/Q 0.0224f
C20254 _217_/A _327_/D 6.2e-20
C20255 _341_/Q _298_/a_27_7# 3.6e-19
C20256 _322_/a_761_249# result[6] 0.00812f
C20257 _329_/a_543_7# output20/a_27_7# 3.66e-21
C20258 _333_/a_761_249# _207_/C 2.69e-19
C20259 _333_/a_1283_n19# _206_/A 0.0839f
C20260 _294_/Y _266_/a_199_7# 7.55e-19
C20261 _313_/Q _337_/D 7.38e-21
C20262 _297_/A _313_/a_27_7# 2.57e-21
C20263 clkbuf_0_clk/a_110_7# _203_/a_209_257# 7.27e-21
C20264 _334_/a_193_7# _343_/Q 5.23e-21
C20265 _196_/A _295_/a_512_7# 2.02e-19
C20266 _181_/X _295_/a_409_7# 0.00427f
C20267 _172_/A _174_/a_27_257# 0.0726f
C20268 _336_/a_193_7# _225_/B 1e-20
C20269 _336_/a_761_249# _336_/Q 6.81e-22
C20270 _322_/Q _282_/a_39_257# 0.0146f
C20271 _308_/S _286_/Y 6.44e-20
C20272 _267_/A _311_/a_1462_7# 8.56e-20
C20273 _343_/CLK _333_/a_1108_7# 3.88e-21
C20274 _334_/Q _333_/a_27_7# 0.00642f
C20275 _149_/a_27_7# _317_/D 0.00126f
C20276 _267_/B _312_/a_543_7# 2.29e-21
C20277 _231_/a_306_7# _150_/C 0.00103f
C20278 _188_/S _150_/a_27_7# 0.0765f
C20279 _242_/A _227_/A 1.3e-20
C20280 _196_/A _333_/Q 0.00219f
C20281 _340_/D VPWR 0.242f
C20282 _286_/B _190_/A 0.0907f
C20283 _193_/Y VGND 0.263f
C20284 _309_/a_1270_373# _284_/A 3.05e-19
C20285 _227_/A _335_/Q 0.339f
C20286 _283_/Y _339_/Q 3.04e-19
C20287 _347_/Q _297_/Y 0.712f
C20288 _294_/Y _160_/X 0.00721f
C20289 _343_/a_448_7# _269_/A 2.94e-20
C20290 _273_/A _286_/B 0.0435f
C20291 _317_/a_448_7# _317_/D 0.00445f
C20292 _283_/A _217_/A 0.123f
C20293 _275_/Y _166_/Y 6.68e-20
C20294 result[0] _341_/a_1283_n19# 2.84e-19
C20295 _333_/a_27_7# _191_/B 0.0322f
C20296 _308_/S _250_/a_215_7# 4.52e-20
C20297 _340_/CLK _194_/A 0.0095f
C20298 _325_/a_193_7# _331_/D 7.99e-21
C20299 _310_/a_448_7# _310_/Q 9.03e-20
C20300 _317_/Q _304_/X 0.00299f
C20301 _329_/a_543_7# _218_/a_250_257# 4.99e-19
C20302 _329_/a_1283_n19# _218_/a_93_n19# 6.16e-19
C20303 _199_/a_93_n19# _199_/a_346_7# -3.48e-20
C20304 _322_/Q _327_/Q 0.0103f
C20305 _316_/D _177_/A 1.61e-20
C20306 _338_/a_193_7# _340_/CLK 0.575f
C20307 cal _154_/a_27_7# 0.00319f
C20308 _256_/a_209_7# _190_/A 0.00297f
C20309 _247_/a_113_257# VPWR 0.0532f
C20310 _327_/a_651_373# _216_/X 1.44e-20
C20311 _346_/SET_B _347_/a_27_7# 0.0126f
C20312 _324_/a_543_7# _248_/B 7.32e-20
C20313 _258_/S _340_/CLK 0.368f
C20314 _309_/a_543_7# _306_/S 7.17e-20
C20315 _265_/B _310_/D 0.413f
C20316 _343_/a_448_7# _343_/D 0.0023f
C20317 _172_/A _324_/Q 0.441f
C20318 _208_/a_78_159# _208_/a_292_257# -1.09e-21
C20319 _175_/Y _154_/A 4.56e-21
C20320 _326_/D _304_/a_79_n19# 3.56e-20
C20321 _167_/a_109_257# _297_/B 0.0268f
C20322 cal _179_/a_27_7# 0.0267f
C20323 _327_/a_1108_7# _238_/B 6.24e-20
C20324 ctln[4] rstn 5.44e-19
C20325 _321_/a_543_7# _242_/B 4.61e-21
C20326 _288_/A _288_/Y 0.0112f
C20327 repeater43/X _162_/X 1.3e-20
C20328 _327_/a_27_7# _327_/a_639_7# -0.0014f
C20329 _322_/a_1462_7# result[7] 1.19e-19
C20330 _248_/B _217_/A 4.28e-19
C20331 _345_/Q trimb[4] 3.49e-20
C20332 _340_/a_543_7# _340_/CLK 5.06e-19
C20333 _181_/X _216_/a_27_7# 0.00707f
C20334 output5/a_27_7# VGND 0.0532f
C20335 _315_/Q _316_/a_651_373# 2.8e-19
C20336 _341_/a_543_7# _341_/D 0.036f
C20337 _329_/a_639_7# _330_/Q 3.26e-19
C20338 _161_/Y _174_/a_373_7# 1.12e-19
C20339 _255_/B _314_/D 2.35e-20
C20340 _331_/D _331_/a_639_7# 0.00132f
C20341 _332_/a_1283_n19# _332_/Q 0.0246f
C20342 _332_/a_543_7# _333_/Q 0.00925f
C20343 _316_/D _325_/D 9.7e-21
C20344 _332_/a_1108_7# _207_/X 5.5e-36
C20345 _326_/a_27_7# _326_/a_639_7# -0.0015f
C20346 _297_/B _297_/Y 0.0449f
C20347 _328_/a_448_7# _329_/Q 0.0254f
C20348 _328_/a_1283_n19# _238_/B 0.0163f
C20349 trimb[1] comp 0.0654f
C20350 _305_/a_76_159# _260_/A 0.00761f
C20351 _317_/Q _272_/a_39_257# 0.00775f
C20352 _341_/Q _326_/Q 2.6e-19
C20353 repeater43/X _333_/a_1217_7# -2.96e-19
C20354 _338_/a_761_249# _346_/SET_B 0.0053f
C20355 _338_/a_543_7# _338_/D 0.0336f
C20356 _329_/a_448_7# VGND -0.00369f
C20357 _329_/a_1270_373# VPWR -1.4e-19
C20358 _347_/Q _242_/A 1.95e-19
C20359 _313_/D input1/X 5.81e-20
C20360 _197_/X _202_/a_250_257# 0.00641f
C20361 _344_/a_476_7# _344_/Q 2.15e-19
C20362 _344_/a_27_7# _344_/D 0.0892f
C20363 _341_/a_1108_7# _248_/A 1.96e-19
C20364 _342_/a_1108_7# cal 6.65e-19
C20365 _342_/a_1283_n19# input1/X 6.96e-19
C20366 comp VGND 0.545f
C20367 _286_/B _178_/a_27_7# 1.04e-20
C20368 _294_/A _309_/a_543_7# 0.0355f
C20369 _294_/Y _309_/a_193_7# 1.03e-20
C20370 input1/X _197_/X 0.00504f
C20371 _301_/a_240_7# _160_/X 0.00212f
C20372 _329_/a_651_373# repeater42/a_27_7# 1.47e-20
C20373 _346_/SET_B _162_/A 5.96e-20
C20374 _340_/a_1283_n19# _346_/SET_B -0.00538f
C20375 _182_/X _226_/a_79_n19# 0.00116f
C20376 _196_/A _226_/a_297_7# 1.74e-19
C20377 _216_/X _346_/SET_B 0.408f
C20378 _328_/a_193_7# _328_/a_448_7# -0.00831f
C20379 _324_/Q _244_/B 0.0154f
C20380 _227_/A _336_/Q 0.00175f
C20381 _343_/CLK _176_/a_27_7# 0.00104f
C20382 _334_/a_1462_7# _343_/Q 3.65e-20
C20383 _162_/X _191_/B 3e-21
C20384 _267_/B _263_/B 0.289f
C20385 _321_/Q _242_/A 0.00371f
C20386 clkbuf_2_0_0_clk/a_75_172# clkbuf_2_1_0_clk/A 0.0191f
C20387 _329_/Q _346_/SET_B 0.494f
C20388 _172_/A _228_/A 0.0198f
C20389 _215_/A _298_/A 0.0271f
C20390 _271_/A _270_/a_39_257# 0.00816f
C20391 _167_/X _306_/a_439_7# 1.31e-20
C20392 _292_/A _163_/a_215_7# 0.00429f
C20393 _327_/a_761_249# _346_/SET_B 0.0176f
C20394 _317_/Q VGND 1.11f
C20395 result[2] VPWR 0.241f
C20396 _343_/CLK _332_/a_27_7# 1.32e-20
C20397 _339_/Q _312_/a_27_7# 1.35e-19
C20398 _279_/Y _248_/A 0.0449f
C20399 _144_/a_27_7# _246_/B 1.44e-21
C20400 _205_/a_297_7# VGND 0.0396f
C20401 _163_/a_215_7# _160_/A 7.42e-19
C20402 _177_/a_27_7# _150_/C 1.29e-19
C20403 _172_/A _168_/a_397_257# 4.82e-20
C20404 input4/X _338_/a_27_7# 5.7e-19
C20405 _343_/a_1283_n19# _175_/Y 0.0705f
C20406 _342_/a_761_249# sample 4.8e-19
C20407 _342_/a_1283_n19# _286_/Y 1.4e-21
C20408 _242_/A _297_/B 0.01f
C20409 _315_/Q _341_/D 0.00381f
C20410 _341_/Q _154_/A 6.88e-20
C20411 _298_/B _153_/A 1.08e-21
C20412 _331_/Q _331_/a_651_373# 8.49e-19
C20413 result[7] _331_/Q 0.00105f
C20414 _242_/A _318_/a_193_7# 0.0148f
C20415 _266_/a_113_257# _265_/B 1.09e-20
C20416 _316_/a_448_7# _331_/CLK 1.68e-20
C20417 _316_/a_1108_7# _316_/D 1.09e-19
C20418 _279_/Y _331_/CLK 2.04e-20
C20419 _310_/D _310_/Q 0.012f
C20420 _329_/a_761_249# _330_/D 0.0101f
C20421 _311_/a_1108_7# _297_/Y 3.56e-36
C20422 _316_/Q _342_/Q 1.53e-20
C20423 _343_/Q _226_/a_382_257# 5.25e-20
C20424 _301_/a_149_7# VGND 0.00105f
C20425 ctln[5] _332_/Q 0.00346f
C20426 _279_/Y _190_/A 0.0135f
C20427 _320_/Q _321_/D 0.00688f
C20428 _328_/a_193_7# _346_/SET_B 0.0127f
C20429 input1/X _312_/a_193_7# 2.08e-19
C20430 _321_/Q _322_/D 9.99e-20
C20431 _326_/a_1108_7# _248_/A 0.0202f
C20432 _334_/a_193_7# _334_/a_448_7# -0.00779f
C20433 _293_/a_39_257# _340_/Q 0.00845f
C20434 _181_/X _327_/Q 0.0251f
C20435 _290_/A _311_/D 7.04e-21
C20436 _204_/a_27_7# _332_/Q 2.3e-19
C20437 _204_/a_27_257# _333_/Q 0.00152f
C20438 _327_/a_1108_7# _331_/CLK 0.0642f
C20439 _321_/a_448_7# _321_/Q 0.0257f
C20440 _321_/a_1108_7# _330_/Q 2.84e-20
C20441 _279_/Y _273_/A 0.0811f
C20442 _304_/a_257_159# _144_/A 3.24e-20
C20443 _343_/a_27_7# input3/a_27_7# 2.13e-21
C20444 _329_/a_1283_n19# _328_/D 2.52e-20
C20445 _285_/A _290_/Y 1.73e-20
C20446 _324_/a_27_7# _314_/a_27_7# 9.14e-21
C20447 _172_/A _216_/A 0.00875f
C20448 _338_/a_193_7# _337_/a_651_373# 3.04e-21
C20449 _338_/a_651_373# _337_/a_193_7# 2.36e-20
C20450 _304_/X _298_/A 0.00423f
C20451 _326_/a_543_7# _236_/B 7.33e-22
C20452 _234_/B VPWR 0.43f
C20453 _326_/a_1108_7# _331_/CLK 6.56e-21
C20454 _326_/a_1283_n19# _316_/D 1.73e-19
C20455 _144_/A _177_/A 2.99e-20
C20456 result[0] _248_/A 0.0033f
C20457 _258_/S _313_/a_543_7# 4.3e-20
C20458 _147_/A _347_/a_27_7# 5.08e-19
C20459 _172_/A _251_/a_510_7# 2.72e-19
C20460 _311_/a_193_7# _310_/a_1108_7# 2.56e-21
C20461 _286_/B _313_/a_805_7# 3.04e-19
C20462 _321_/a_1283_n19# VPWR 0.0295f
C20463 _321_/a_761_249# VGND 0.00728f
C20464 _275_/Y _297_/Y 0.00672f
C20465 _327_/a_1108_7# _273_/A 2.56e-19
C20466 ctln[4] clkbuf_2_0_0_clk/a_75_172# 1.31e-19
C20467 _290_/A _285_/Y 5.22e-19
C20468 _216_/A _232_/X 0.00112f
C20469 _338_/a_543_7# _343_/CLK 5.91e-20
C20470 _169_/Y _299_/X 0.512f
C20471 _188_/S _250_/X 3.26e-21
C20472 _325_/a_1108_7# _223_/a_93_n19# 8.81e-20
C20473 _299_/X _225_/B 2.82e-20
C20474 _322_/D _318_/a_193_7# 3.83e-19
C20475 _346_/SET_B _190_/a_27_7# 1.28e-19
C20476 _326_/a_1108_7# _273_/A 3.96e-19
C20477 _328_/a_1283_n19# _331_/CLK 7.23e-22
C20478 _321_/a_543_7# _318_/a_1283_n19# 1.57e-20
C20479 _321_/a_448_7# _318_/a_193_7# 9.94e-21
C20480 _323_/a_193_7# _269_/A 0.00304f
C20481 _228_/A _244_/B 0.0107f
C20482 _237_/a_113_257# _327_/Q 3.64e-20
C20483 _232_/X _221_/a_584_7# 7.11e-20
C20484 _288_/A _337_/Q 0.00253f
C20485 _153_/a_215_257# VPWR 0.00345f
C20486 output8/a_27_7# trim[3] 0.0137f
C20487 repeater43/X _298_/C 0.0134f
C20488 _209_/X VPWR 0.194f
C20489 _326_/a_543_7# _326_/D 2.69e-19
C20490 _296_/Y _286_/B 0.00623f
C20491 _340_/CLK _201_/a_27_7# 1.04e-20
C20492 _260_/B _313_/a_193_7# 0.00217f
C20493 _275_/Y _310_/a_193_7# 0.0113f
C20494 _287_/a_39_257# _337_/Q 0.0319f
C20495 _277_/A _279_/A 0.00133f
C20496 _274_/a_39_257# _346_/SET_B 4.63e-19
C20497 _238_/B _319_/a_448_7# 0.00264f
C20498 _310_/a_1270_373# VGND 4.61e-20
C20499 _310_/a_805_7# VPWR 0.00221f
C20500 repeater43/X _332_/a_448_7# 1.27e-21
C20501 _344_/a_1224_7# _344_/Q 2.92e-19
C20502 _181_/X _192_/B 0.644f
C20503 output19/a_27_7# _328_/Q 1.53e-20
C20504 _165_/a_493_257# _158_/Y 2.89e-19
C20505 _343_/D _323_/a_193_7# 0.0185f
C20506 _185_/A _323_/a_543_7# 0.00913f
C20507 _258_/a_439_7# _306_/S 9.15e-19
C20508 _334_/a_1108_7# _333_/Q 2.16e-20
C20509 _265_/B VPWR 1.48f
C20510 _267_/B _194_/A 2.69e-20
C20511 _277_/Y _215_/A 0.00634f
C20512 _308_/X _306_/S 0.0079f
C20513 _346_/a_476_7# _346_/SET_B 0.055f
C20514 _145_/A _177_/A 0.00587f
C20515 _172_/B _284_/A 9.79e-21
C20516 _216_/A _203_/a_80_n19# 1.99e-20
C20517 _325_/a_27_7# _181_/X 0.0146f
C20518 _209_/a_109_257# VPWR -0.0178f
C20519 _330_/Q _326_/Q 0.00102f
C20520 _163_/a_78_159# _346_/SET_B 0.00118f
C20521 _347_/Q _314_/a_761_249# 1.81e-20
C20522 _339_/a_1108_7# _338_/a_543_7# 5.26e-20
C20523 _271_/Y _204_/Y 5.52e-20
C20524 _309_/a_1108_7# _310_/a_1108_7# 8.64e-19
C20525 _337_/a_27_7# _340_/CLK 0.257f
C20526 _198_/a_256_7# _193_/Y 1.43e-19
C20527 _198_/a_584_7# _340_/Q 0.00105f
C20528 _258_/S _267_/B 0.089f
C20529 _294_/A trim[0] 0.0727f
C20530 _275_/Y _242_/A 2.2e-20
C20531 _294_/Y _285_/A 0.864f
C20532 _335_/a_543_7# _335_/Q 0.00154f
C20533 _335_/a_761_249# _204_/Y 2.43e-20
C20534 ctln[6] _197_/X 0.01f
C20535 _183_/a_553_257# _304_/a_79_n19# 1.04e-19
C20536 _323_/Q valid 1.65e-21
C20537 _299_/X _170_/a_226_257# 2.03e-19
C20538 _325_/a_543_7# _304_/a_257_159# 8.66e-20
C20539 _325_/a_1283_n19# _304_/a_79_n19# 2.28e-19
C20540 _308_/S _255_/X 1.05e-21
C20541 _315_/Q _343_/CLK 0.246f
C20542 repeater43/X _341_/a_639_7# -7.75e-19
C20543 _316_/D _248_/A 0.0186f
C20544 _309_/a_27_7# _265_/B 0.00892f
C20545 _343_/Q _192_/B 1.41e-19
C20546 _294_/Y _344_/a_193_7# 1.08e-20
C20547 _298_/C _191_/B 0.0698f
C20548 _184_/a_76_159# _298_/a_27_7# 9.09e-22
C20549 _242_/B _318_/D 0.196f
C20550 _340_/a_1108_7# _339_/a_1108_7# 3.65e-19
C20551 _334_/a_193_7# _206_/A 1.03e-19
C20552 _242_/A _318_/a_1462_7# 1.49e-19
C20553 result[0] _145_/a_113_7# 1.63e-21
C20554 output14/a_27_7# result[7] 0.00724f
C20555 _331_/CLK _316_/D 0.114f
C20556 _344_/a_1140_373# _290_/A 5.59e-19
C20557 ctln[5] _339_/a_193_7# 1.71e-19
C20558 _315_/a_543_7# VPWR -0.0042f
C20559 _315_/a_193_7# VGND 0.00787f
C20560 _298_/A VGND 0.691f
C20561 input3/a_27_7# ctln[0] 7.38e-21
C20562 _342_/Q _186_/a_297_7# 0.00191f
C20563 _294_/A _311_/Q 2.54e-20
C20564 _214_/a_109_257# _327_/D 9.29e-20
C20565 _336_/a_448_7# VGND -0.00194f
C20566 _336_/a_1270_373# VPWR -2.59e-19
C20567 output38/a_27_7# _162_/A 1.07e-21
C20568 _324_/a_448_7# _227_/A 0.0126f
C20569 _294_/A _258_/a_439_7# 4.16e-21
C20570 _328_/a_1462_7# _346_/SET_B -9.14e-19
C20571 _317_/a_761_249# _316_/a_27_7# 8.7e-21
C20572 _317_/a_193_7# _316_/a_193_7# 1.56e-20
C20573 _324_/a_193_7# _324_/a_543_7# -0.0102f
C20574 input1/a_75_172# _312_/D 1.92e-19
C20575 _334_/a_761_249# _343_/CLK 3.04e-20
C20576 _334_/a_193_7# _334_/D 0.513f
C20577 repeater43/X _229_/a_489_373# 0.00694f
C20578 _315_/D _314_/a_1283_n19# 0.00159f
C20579 _273_/A _316_/D 7.03e-20
C20580 _314_/a_27_7# VPWR 0.115f
C20581 _346_/SET_B _319_/a_543_7# 0.00999f
C20582 _242_/B _217_/A 4.21e-20
C20583 clkbuf_0_clk/X _299_/a_215_7# 5.95e-19
C20584 _255_/B _188_/S 0.00379f
C20585 cal.t0 0 0.0245f
C20586 cal.t1 0 0.0387f
C20587 cal.n0 0 0.0814f
C20588 cal.n1 0 1.48f
C20589 clk.t5 0 0.0112f
C20590 clk.t1 0 0.0238f
C20591 clk.t4 0 0.0112f
C20592 clk.t0 0 0.0238f
C20593 clk.t7 0 0.0112f
C20594 clk.t3 0 0.0238f
C20595 clk.t2 0 0.0112f
C20596 clk.t6 0 0.0238f
C20597 clk.n0 0 0.0544f
C20598 clk.n1 0 0.0717f
C20599 clk.n2 0 0.0717f
C20600 clk.n3 0 0.067f
C20601 clk.n4 0 0.0339f
C20602 clk.n5 0 0.779f
C20603 VGND.t374 0 0.0792f
C20604 VGND.n0 0 0.0243f
C20605 VGND.n1 0 0.0547f
C20606 VGND.t288 0 0.0409f
C20607 VGND.n2 0 0.062f
C20608 VGND.n3 0 0.0285f
C20609 VGND.n4 0 0.015f
C20610 VGND.n5 0 0.037f
C20611 VGND.n6 0 0.0166f
C20612 VGND.n7 0 0.0375f
C20613 VGND.n8 0 0.0166f
C20614 VGND.n9 0 0.0331f
C20615 VGND.n10 0 0.0166f
C20616 VGND.n11 0 0.0166f
C20617 VGND.n12 0 0.00981f
C20618 VGND.n13 0 0.028f
C20619 VGND.n14 0 0.0261f
C20620 VGND.n15 0 0.015f
C20621 VGND.n16 0 0.00373f
C20622 VGND.n17 0 0.0166f
C20623 VGND.n18 0 0.0278f
C20624 VGND.n19 0 0.0166f
C20625 VGND.n20 0 0.0331f
C20626 VGND.n21 0 0.0278f
C20627 VGND.n22 0 0.0331f
C20628 VGND.t24 0 0.128f
C20629 VGND.n23 0 0.154f
C20630 VGND.n24 0 0.0263f
C20631 VGND.n25 0 0.0331f
C20632 VGND.n26 0 0.0367f
C20633 VGND.n27 0 0.026f
C20634 VGND.n28 0 0.0253f
C20635 VGND.n29 0 0.0259f
C20636 VGND.n30 0 0.0279f
C20637 VGND.n31 0 0.0291f
C20638 VGND.n32 0 0.0291f
C20639 VGND.n33 0 0.0278f
C20640 VGND.n34 0 0.00234f
C20641 VGND.n35 0 0.00369f
C20642 VGND.n36 0 0.00234f
C20643 VGND.n37 0 7.2e-19
C20644 VGND.n38 0 0.00207f
C20645 VGND.n39 0 0.00207f
C20646 VGND.n40 0 0.00207f
C20647 VGND.n41 0 0.00297f
C20648 VGND.n42 0 0.00234f
C20649 VGND.n43 0 0.00274f
C20650 VGND.n44 0 0.00173f
C20651 VGND.n45 0 0.0039f
C20652 VGND.n46 0 0.00269f
C20653 VGND.n47 0 0.00207f
C20654 VGND.n48 0 0.00287f
C20655 VGND.n49 0 0.00173f
C20656 VGND.n51 0 0.00274f
C20657 VGND.n52 0 0.00173f
C20658 VGND.n53 0 0.00261f
C20659 VGND.n54 0 0.00207f
C20660 VGND.n55 0 0.00135f
C20661 VGND.n56 0 7.2e-19
C20662 VGND.n57 0 9.9e-19
C20663 VGND.n58 0 0.00207f
C20664 VGND.n59 0 0.00315f
C20665 VGND.n60 0 0.00297f
C20666 VGND.n61 0 0.00234f
C20667 VGND.n62 0 0.0271f
C20668 VGND.t270 0 0.0946f
C20669 VGND.n63 0 0.0183f
C20670 VGND.n64 0 0.0961f
C20671 VGND.n65 0 0.0252f
C20672 VGND.n66 0 0.0271f
C20673 VGND.n67 0 0.0321f
C20674 VGND.n68 0 0.0271f
C20675 VGND.t281 0 0.0946f
C20676 VGND.n69 0 0.0183f
C20677 VGND.n70 0 0.0961f
C20678 VGND.n71 0 0.0252f
C20679 VGND.n72 0 0.0271f
C20680 VGND.n73 0 0.0321f
C20681 VGND.n74 0 0.0452f
C20682 VGND.t269 0 0.128f
C20683 VGND.n75 0 0.154f
C20684 VGND.n76 0 0.0263f
C20685 VGND.n77 0 0.0452f
C20686 VGND.n78 0 0.00234f
C20687 VGND.n79 0 0.00287f
C20688 VGND.n80 0 0.00207f
C20689 VGND.n81 0 0.00274f
C20690 VGND.n82 0 0.00403f
C20691 VGND.n83 0 0.00493f
C20692 VGND.n84 0 0.00126f
C20693 VGND.n85 0 0.00173f
C20694 VGND.n87 0 0.00274f
C20695 VGND.n88 0 0.00173f
C20696 VGND.n89 0 0.00207f
C20697 VGND.n90 0 0.00603f
C20698 VGND.n91 0 0.00234f
C20699 VGND.n92 0 0.00135f
C20700 VGND.n93 0 0.00189f
C20701 VGND.n94 0 0.00369f
C20702 VGND.n95 0 0.00252f
C20703 VGND.n96 0 7.2e-19
C20704 VGND.n97 0 7.2e-19
C20705 VGND.n98 0 0.00162f
C20706 VGND.n99 0 0.0331f
C20707 VGND.n100 0 0.0343f
C20708 VGND.n101 0 0.0343f
C20709 VGND.n102 0 0.0331f
C20710 VGND.n103 0 0.0319f
C20711 VGND.n104 0 0.0416f
C20712 VGND.n105 0 0.0243f
C20713 VGND.t130 0 0.0812f
C20714 VGND.t388 0 0.0813f
C20715 VGND.n106 0 0.139f
C20716 VGND.n107 0 0.03f
C20717 VGND.t60 0 0.128f
C20718 VGND.n108 0 0.154f
C20719 VGND.n109 0 0.0517f
C20720 VGND.n110 0 0.0319f
C20721 VGND.n111 0 0.0339f
C20722 VGND.t97 0 0.0792f
C20723 VGND.n112 0 0.0243f
C20724 VGND.n113 0 0.0547f
C20725 VGND.n114 0 0.0259f
C20726 VGND.n115 0 0.0259f
C20727 VGND.n116 0 0.00126f
C20728 VGND.n117 0 0.00274f
C20729 VGND.n118 0 0.00173f
C20730 VGND.n119 0 0.00413f
C20731 VGND.n120 0 0.00261f
C20732 VGND.n121 0 0.00207f
C20733 VGND.n122 0 0.00135f
C20734 VGND.n123 0 0.00423f
C20735 VGND.n124 0 0.00414f
C20736 VGND.n125 0 0.00148f
C20737 VGND.n126 0 0.026f
C20738 VGND.n127 0 0.178f
C20739 VGND.n128 0 0.0636f
C20740 VGND.n129 0 0.0314f
C20741 VGND.t111 0 0.226f
C20742 VGND.n130 0 0.344f
C20743 VGND.t238 0 0.171f
C20744 VGND.n131 0 0.059f
C20745 VGND.n132 0 0.0503f
C20746 VGND.n133 0 0.304f
C20747 VGND.n134 0 0.037f
C20748 VGND.t123 0 0.0813f
C20749 VGND.t237 0 0.157f
C20750 VGND.n135 0 0.199f
C20751 VGND.t90 0 0.0799f
C20752 VGND.n136 0 0.0723f
C20753 VGND.t260 0 0.0445f
C20754 VGND.t233 0 0.0445f
C20755 VGND.n137 0 0.244f
C20756 VGND.n138 0 0.0159f
C20757 VGND.n139 0 0.0367f
C20758 VGND.n140 0 0.0266f
C20759 VGND.n141 0 0.0166f
C20760 VGND.t212 0 0.0429f
C20761 VGND.n142 0 0.148f
C20762 VGND.n143 0 0.0241f
C20763 VGND.n144 0 0.00981f
C20764 VGND.n145 0 0.00828f
C20765 VGND.n146 0 0.0192f
C20766 VGND.n147 0 0.0733f
C20767 VGND.n148 0 0.015f
C20768 VGND.n149 0 0.0166f
C20769 VGND.n150 0 0.0166f
C20770 VGND.n151 0 0.0336f
C20771 VGND.n152 0 0.0482f
C20772 VGND.n153 0 0.0251f
C20773 VGND.n154 0 0.0172f
C20774 VGND.n155 0 0.0496f
C20775 VGND.n156 0 0.139f
C20776 VGND.n157 0 0.037f
C20777 VGND.n158 0 0.00828f
C20778 VGND.n159 0 0.015f
C20779 VGND.n160 0 0.00981f
C20780 VGND.n161 0 0.0584f
C20781 VGND.n162 0 0.0651f
C20782 VGND.n163 0 0.015f
C20783 VGND.n164 0 0.0597f
C20784 VGND.n165 0 0.0166f
C20785 VGND.n166 0 0.0166f
C20786 VGND.n167 0 0.0328f
C20787 VGND.n168 0 0.0249f
C20788 VGND.n169 0 0.0119f
C20789 VGND.t147 0 0.132f
C20790 VGND.n170 0 0.0976f
C20791 VGND.n171 0 0.0503f
C20792 VGND.n172 0 0.0888f
C20793 VGND.t132 0 0.232f
C20794 VGND.n173 0 0.389f
C20795 VGND.n174 0 0.0563f
C20796 VGND.t219 0 0.226f
C20797 VGND.n175 0 0.355f
C20798 VGND.n176 0 0.0332f
C20799 VGND.n177 0 0.0318f
C20800 VGND.n178 0 0.0348f
C20801 VGND.t267 0 0.0792f
C20802 VGND.n179 0 0.054f
C20803 VGND.n180 0 0.0243f
C20804 VGND.n181 0 0.014f
C20805 VGND.n182 0 0.0331f
C20806 VGND.n183 0 0.0166f
C20807 VGND.n184 0 0.0368f
C20808 VGND.n185 0 0.0166f
C20809 VGND.n186 0 0.0166f
C20810 VGND.n187 0 0.0149f
C20811 VGND.n188 0 0.00837f
C20812 VGND.n189 0 0.00828f
C20813 VGND.n190 0 0.0501f
C20814 VGND.n191 0 0.00828f
C20815 VGND.n192 0 0.0303f
C20816 VGND.n193 0 0.0384f
C20817 VGND.n194 0 0.0221f
C20818 VGND.n195 0 0.059f
C20819 VGND.n196 0 0.0166f
C20820 VGND.n197 0 0.0597f
C20821 VGND.n198 0 0.0166f
C20822 VGND.n199 0 0.015f
C20823 VGND.n200 0 0.0119f
C20824 VGND.n201 0 0.0604f
C20825 VGND.t226 0 0.226f
C20826 VGND.n202 0 0.344f
C20827 VGND.n203 0 0.0651f
C20828 VGND.n204 0 0.051f
C20829 VGND.n205 0 0.254f
C20830 VGND.n206 0 0.0249f
C20831 VGND.n207 0 0.0328f
C20832 VGND.n208 0 0.0144f
C20833 VGND.n209 0 0.00819f
C20834 VGND.n210 0 0.009f
C20835 VGND.n211 0 0.0816f
C20836 VGND.n212 0 0.00189f
C20837 VGND.n213 0 8.1e-19
C20838 VGND.n214 0 5.1e-19
C20839 VGND.n215 0 0.00135f
C20840 VGND.n216 0 9e-19
C20841 VGND.n217 0 0.00872f
C20842 VGND.n218 0 0.00198f
C20843 VGND.n219 0 7.2e-19
C20844 VGND.n220 0 0.0191f
C20845 VGND.n221 0 0.049f
C20846 VGND.n222 0 0.229f
C20847 VGND.n223 0 0.0944f
C20848 VGND.n224 0 0.168f
C20849 VGND.n225 0 0.219f
C20850 VGND.n226 0 0.19f
C20851 VGND.n227 0 0.213f
C20852 VGND.n228 0 0.19f
C20853 VGND.n229 0 0.19f
C20854 VGND.n230 0 0.19f
C20855 VGND.n231 0 0.19f
C20856 VGND.n232 0 0.19f
C20857 VGND.n233 0 0.19f
C20858 VGND.n234 0 0.19f
C20859 VGND.n235 0 0.19f
C20860 VGND.n236 0 0.19f
C20861 VGND.n237 0 0.19f
C20862 VGND.n238 0 0.19f
C20863 VGND.n239 0 0.19f
C20864 VGND.n240 0 0.19f
C20865 VGND.n241 0 0.19f
C20866 VGND.n242 0 0.19f
C20867 VGND.n243 0 0.19f
C20868 VGND.n244 0 0.19f
C20869 VGND.n245 0 0.19f
C20870 VGND.n246 0 0.19f
C20871 VGND.n247 0 0.19f
C20872 VGND.n248 0 0.0316f
C20873 VGND.n249 0 0.0317f
C20874 VGND.n250 0 0.0252f
C20875 VGND.n251 0 0.03f
C20876 VGND.n252 0 0.0553f
C20877 VGND.n253 0 0.0191f
C20878 VGND.t138 0 0.0837f
C20879 VGND.t17 0 0.0837f
C20880 VGND.n254 0 0.324f
C20881 VGND.t79 0 0.0837f
C20882 VGND.t333 0 0.0837f
C20883 VGND.n255 0 0.324f
C20884 VGND.t168 0 0.128f
C20885 VGND.n256 0 0.154f
C20886 VGND.n257 0 0.0255f
C20887 VGND.n258 0 0.00627f
C20888 VGND.t78 0 0.0816f
C20889 VGND.n259 0 0.139f
C20890 VGND.n260 0 0.00234f
C20891 VGND.n261 0 0.00369f
C20892 VGND.n262 0 0.00234f
C20893 VGND.n263 0 7.2e-19
C20894 VGND.n264 0 0.00207f
C20895 VGND.n265 0 0.00207f
C20896 VGND.n266 0 0.00207f
C20897 VGND.n267 0 0.00297f
C20898 VGND.n268 0 0.00234f
C20899 VGND.n269 0 0.178f
C20900 VGND.n271 0 0.00274f
C20901 VGND.n272 0 0.00173f
C20902 VGND.n273 0 0.00413f
C20903 VGND.n274 0 0.00207f
C20904 VGND.n275 0 0.00287f
C20905 VGND.n276 0 0.0039f
C20906 VGND.n277 0 0.00269f
C20907 VGND.n278 0 0.00173f
C20908 VGND.n280 0 0.00274f
C20909 VGND.n281 0 0.00173f
C20910 VGND.n282 0 0.00369f
C20911 VGND.n283 0 0.00234f
C20912 VGND.n284 0 7.2e-19
C20913 VGND.n285 0 0.00207f
C20914 VGND.n286 0 0.00207f
C20915 VGND.n287 0 0.00207f
C20916 VGND.n288 0 0.00297f
C20917 VGND.n289 0 0.00234f
C20918 VGND.n290 0 0.00234f
C20919 VGND.n291 0 0.0331f
C20920 VGND.n292 0 0.0496f
C20921 VGND.n293 0 0.0513f
C20922 VGND.n294 0 0.0265f
C20923 VGND.n295 0 0.0492f
C20924 VGND.n296 0 0.057f
C20925 VGND.n297 0 0.0468f
C20926 VGND.n298 0 0.0367f
C20927 VGND.n299 0 0.00414f
C20928 VGND.t329 0 0.0837f
C20929 VGND.n300 0 0.0291f
C20930 VGND.n301 0 0.0774f
C20931 VGND.n302 0 0.0944f
C20932 VGND.n303 0 0.0566f
C20933 VGND.n304 0 9.9e-19
C20934 VGND.n305 0 0.00162f
C20935 VGND.n306 0 8.1e-19
C20936 VGND.n307 0 0.213f
C20937 VGND.t272 0 0.0792f
C20938 VGND.n308 0 0.0243f
C20939 VGND.n309 0 0.0547f
C20940 VGND.n310 0 0.0291f
C20941 VGND.n311 0 0.0513f
C20942 VGND.t384 0 0.121f
C20943 VGND.t240 0 0.155f
C20944 VGND.n312 0 0.0449f
C20945 VGND.n313 0 0.163f
C20946 VGND.n314 0 0.123f
C20947 VGND.n315 0 0.0368f
C20948 VGND.t241 0 0.0837f
C20949 VGND.t131 0 0.0445f
C20950 VGND.t108 0 0.0445f
C20951 VGND.n316 0 0.243f
C20952 VGND.n317 0 0.032f
C20953 VGND.n318 0 0.0351f
C20954 VGND.t385 0 0.0837f
C20955 VGND.n319 0 0.324f
C20956 VGND.n320 0 0.0509f
C20957 VGND.n321 0 0.015f
C20958 VGND.n322 0 0.00373f
C20959 VGND.n323 0 0.0166f
C20960 VGND.n324 0 0.0544f
C20961 VGND.n325 0 0.00981f
C20962 VGND.n326 0 0.00891f
C20963 VGND.n327 0 0.0321f
C20964 VGND.n328 0 0.0651f
C20965 VGND.n329 0 0.0144f
C20966 VGND.n330 0 0.0597f
C20967 VGND.n331 0 0.0166f
C20968 VGND.n332 0 0.059f
C20969 VGND.n333 0 0.0166f
C20970 VGND.n334 0 0.0166f
C20971 VGND.n335 0 0.0166f
C20972 VGND.n336 0 0.00981f
C20973 VGND.n337 0 0.0687f
C20974 VGND.n338 0 0.0292f
C20975 VGND.n339 0 0.015f
C20976 VGND.n340 0 0.0227f
C20977 VGND.n341 0 0.0166f
C20978 VGND.n342 0 0.0254f
C20979 VGND.n343 0 0.0166f
C20980 VGND.n344 0 0.0044f
C20981 VGND.n345 0 0.0166f
C20982 VGND.n346 0 0.00972f
C20983 VGND.n347 0 0.0283f
C20984 VGND.n348 0 0.0583f
C20985 VGND.n349 0 0.0151f
C20986 VGND.n350 0 0.0331f
C20987 VGND.n351 0 0.0166f
C20988 VGND.n352 0 0.0166f
C20989 VGND.n353 0 0.00981f
C20990 VGND.t346 0 0.0792f
C20991 VGND.n354 0 0.0243f
C20992 VGND.n355 0 0.0547f
C20993 VGND.n356 0 0.00837f
C20994 VGND.t361 0 0.126f
C20995 VGND.n357 0 0.178f
C20996 VGND.n358 0 0.0144f
C20997 VGND.t85 0 0.0837f
C20998 VGND.n359 0 0.00828f
C20999 VGND.t16 0 0.0792f
C21000 VGND.n360 0 0.0243f
C21001 VGND.n361 0 0.0654f
C21002 VGND.n362 0 0.00819f
C21003 VGND.t345 0 0.082f
C21004 VGND.n363 0 0.0934f
C21005 VGND.n364 0 0.0151f
C21006 VGND.n365 0 0.0217f
C21007 VGND.t52 0 0.0816f
C21008 VGND.n366 0 0.139f
C21009 VGND.n367 0 0.00151f
C21010 VGND.n368 0 0.0045f
C21011 VGND.n369 0 0.00207f
C21012 VGND.n370 0 0.00287f
C21013 VGND.n371 0 0.00173f
C21014 VGND.n372 0 0.00269f
C21015 VGND.n373 0 0.0039f
C21016 VGND.n374 0 0.00269f
C21017 VGND.n375 0 0.00173f
C21018 VGND.n377 0 0.00274f
C21019 VGND.n378 0 0.00173f
C21020 VGND.n379 0 0.00207f
C21021 VGND.n380 0 0.0175f
C21022 VGND.n381 0 0.00234f
C21023 VGND.n382 0 0.00135f
C21024 VGND.n383 0 0.00189f
C21025 VGND.n384 0 0.00369f
C21026 VGND.n385 0 0.00252f
C21027 VGND.n386 0 7.2e-19
C21028 VGND.n387 0 7.2e-19
C21029 VGND.n388 0 0.00162f
C21030 VGND.n389 0 0.0533f
C21031 VGND.t114 0 0.0792f
C21032 VGND.n390 0 0.0547f
C21033 VGND.n391 0 0.0411f
C21034 VGND.n392 0 0.057f
C21035 VGND.n393 0 0.0331f
C21036 VGND.n394 0 0.0457f
C21037 VGND.t223 0 0.082f
C21038 VGND.n395 0 0.0934f
C21039 VGND.n396 0 0.0217f
C21040 VGND.n397 0 0.213f
C21041 VGND.t45 0 0.0792f
C21042 VGND.n398 0 0.0243f
C21043 VGND.n399 0 0.0547f
C21044 VGND.n400 0 0.047f
C21045 VGND.n401 0 0.0379f
C21046 VGND.t35 0 0.0837f
C21047 VGND.n402 0 0.186f
C21048 VGND.n403 0 0.015f
C21049 VGND.n404 0 0.0535f
C21050 VGND.t137 0 0.0837f
C21051 VGND.t279 0 0.0445f
C21052 VGND.t163 0 0.0445f
C21053 VGND.n405 0 0.243f
C21054 VGND.n406 0 0.0321f
C21055 VGND.n407 0 0.0349f
C21056 VGND.n408 0 0.186f
C21057 VGND.t3 0 0.126f
C21058 VGND.n409 0 0.223f
C21059 VGND.n410 0 0.0394f
C21060 VGND.n411 0 0.012f
C21061 VGND.n412 0 0.015f
C21062 VGND.n413 0 0.00644f
C21063 VGND.n414 0 0.0401f
C21064 VGND.t154 0 0.126f
C21065 VGND.n415 0 0.178f
C21066 VGND.n416 0 0.0484f
C21067 VGND.n417 0 0.00981f
C21068 VGND.n418 0 0.023f
C21069 VGND.n419 0 0.00837f
C21070 VGND.n420 0 0.0227f
C21071 VGND.n421 0 0.0239f
C21072 VGND.n422 0 0.0149f
C21073 VGND.n423 0 0.0254f
C21074 VGND.n424 0 0.0166f
C21075 VGND.n425 0 0.00325f
C21076 VGND.n426 0 0.0166f
C21077 VGND.n427 0 0.0357f
C21078 VGND.n428 0 0.0166f
C21079 VGND.n429 0 0.0104f
C21080 VGND.n430 0 0.0245f
C21081 VGND.n431 0 0.0379f
C21082 VGND.n432 0 0.0144f
C21083 VGND.n433 0 0.0331f
C21084 VGND.n434 0 0.0166f
C21085 VGND.n435 0 0.0166f
C21086 VGND.n436 0 0.00981f
C21087 VGND.t100 0 0.0792f
C21088 VGND.n437 0 0.0243f
C21089 VGND.n438 0 0.0547f
C21090 VGND.n439 0 0.028f
C21091 VGND.t28 0 0.082f
C21092 VGND.n440 0 0.0934f
C21093 VGND.n441 0 0.0452f
C21094 VGND.t44 0 0.128f
C21095 VGND.n442 0 0.154f
C21096 VGND.n443 0 0.0266f
C21097 VGND.n444 0 0.0304f
C21098 VGND.n445 0 0.0414f
C21099 VGND.n446 0 0.0326f
C21100 VGND.t83 0 0.0837f
C21101 VGND.t194 0 0.0837f
C21102 VGND.n447 0 0.325f
C21103 VGND.n448 0 0.023f
C21104 VGND.n449 0 0.00972f
C21105 VGND.n450 0 0.0166f
C21106 VGND.n451 0 0.015f
C21107 VGND.n452 0 0.0191f
C21108 VGND.n453 0 0.0293f
C21109 VGND.n454 0 0.0275f
C21110 VGND.n455 0 0.015f
C21111 VGND.n456 0 0.085f
C21112 VGND.n457 0 0.0213f
C21113 VGND.n458 0 0.0153f
C21114 VGND.n459 0 0.054f
C21115 VGND.t205 0 0.125f
C21116 VGND.n460 0 0.118f
C21117 VGND.n461 0 0.0478f
C21118 VGND.n462 0 0.085f
C21119 VGND.n463 0 0.00837f
C21120 VGND.n464 0 0.0112f
C21121 VGND.n465 0 0.00891f
C21122 VGND.n466 0 0.028f
C21123 VGND.n467 0 0.0384f
C21124 VGND.n468 0 0.00981f
C21125 VGND.n469 0 0.0513f
C21126 VGND.n470 0 0.0166f
C21127 VGND.n471 0 0.00682f
C21128 VGND.n472 0 0.0166f
C21129 VGND.n473 0 0.015f
C21130 VGND.n474 0 0.00828f
C21131 VGND.n475 0 0.0314f
C21132 VGND.n476 0 0.0291f
C21133 VGND.n477 0 0.00981f
C21134 VGND.n478 0 0.0166f
C21135 VGND.n479 0 0.0331f
C21136 VGND.n480 0 0.0166f
C21137 VGND.n481 0 0.0143f
C21138 VGND.n482 0 0.009f
C21139 VGND.n483 0 0.0291f
C21140 VGND.n484 0 0.229f
C21141 VGND.n485 0 0.00169f
C21142 VGND.n486 0 8.1e-19
C21143 VGND.n487 0 5.1e-19
C21144 VGND.n488 0 0.00135f
C21145 VGND.n489 0 9e-19
C21146 VGND.n490 0 0.0182f
C21147 VGND.n491 0 0.00198f
C21148 VGND.n492 0 7.2e-19
C21149 VGND.n493 0 0.0217f
C21150 VGND.n494 0 0.184f
C21151 VGND.n495 0 0.0252f
C21152 VGND.n496 0 0.0375f
C21153 VGND.t185 0 0.0813f
C21154 VGND.n497 0 0.139f
C21155 VGND.n498 0 0.0349f
C21156 VGND.t207 0 0.0812f
C21157 VGND.n499 0 0.139f
C21158 VGND.n500 0 0.0317f
C21159 VGND.n501 0 0.0481f
C21160 VGND.t198 0 0.082f
C21161 VGND.n502 0 0.0934f
C21162 VGND.n503 0 0.0555f
C21163 VGND.t136 0 0.0813f
C21164 VGND.n504 0 0.139f
C21165 VGND.n505 0 0.0496f
C21166 VGND.n506 0 0.00234f
C21167 VGND.n507 0 0.00369f
C21168 VGND.n508 0 0.00234f
C21169 VGND.n509 0 7.2e-19
C21170 VGND.n510 0 0.00207f
C21171 VGND.n511 0 0.00207f
C21172 VGND.n512 0 0.00207f
C21173 VGND.n513 0 0.00297f
C21174 VGND.n514 0 0.00234f
C21175 VGND.n515 0 0.00274f
C21176 VGND.n516 0 0.00173f
C21177 VGND.n517 0 0.00234f
C21178 VGND.t152 0 0.0792f
C21179 VGND.t180 0 0.082f
C21180 VGND.n518 0 0.0934f
C21181 VGND.n519 0 0.045f
C21182 VGND.n520 0 0.0514f
C21183 VGND.t259 0 0.0813f
C21184 VGND.n521 0 0.139f
C21185 VGND.n522 0 0.0349f
C21186 VGND.n523 0 0.0116f
C21187 VGND.t115 0 0.0813f
C21188 VGND.n524 0 0.139f
C21189 VGND.n525 0 0.0496f
C21190 VGND.n526 0 0.00756f
C21191 VGND.n527 0 0.0157f
C21192 VGND.n528 0 0.0733f
C21193 VGND.n529 0 0.015f
C21194 VGND.n530 0 0.0166f
C21195 VGND.n531 0 0.0166f
C21196 VGND.t244 0 0.157f
C21197 VGND.n532 0 0.199f
C21198 VGND.n533 0 0.0336f
C21199 VGND.n534 0 0.0482f
C21200 VGND.n535 0 0.0251f
C21201 VGND.n536 0 0.0172f
C21202 VGND.n537 0 0.00828f
C21203 VGND.n538 0 0.00494f
C21204 VGND.n539 0 0.0347f
C21205 VGND.n540 0 0.015f
C21206 VGND.n541 0 0.0123f
C21207 VGND.n542 0 0.0166f
C21208 VGND.n543 0 0.0253f
C21209 VGND.n544 0 0.0166f
C21210 VGND.t155 0 0.0812f
C21211 VGND.n545 0 0.139f
C21212 VGND.n546 0 0.0107f
C21213 VGND.n547 0 0.0104f
C21214 VGND.n548 0 0.0165f
C21215 VGND.n549 0 0.00828f
C21216 VGND.n550 0 0.003f
C21217 VGND.n551 0 0.0278f
C21218 VGND.n552 0 0.015f
C21219 VGND.n553 0 0.00373f
C21220 VGND.n554 0 0.0166f
C21221 VGND.n555 0 0.0262f
C21222 VGND.n556 0 0.0166f
C21223 VGND.n557 0 0.06f
C21224 VGND.n558 0 0.0166f
C21225 VGND.n559 0 0.0288f
C21226 VGND.n560 0 0.0221f
C21227 VGND.n561 0 0.0137f
C21228 VGND.n562 0 0.00828f
C21229 VGND.n563 0 0.055f
C21230 VGND.n564 0 0.0509f
C21231 VGND.n565 0 0.0127f
C21232 VGND.n566 0 0.00675f
C21233 VGND.n567 0 0.00153f
C21234 VGND.n568 0 0.0308f
C21235 VGND.n569 0 0.00198f
C21236 VGND.n570 0 0.0179f
C21237 VGND.n571 0 0.00153f
C21238 VGND.n572 0 0.00282f
C21239 VGND.n573 0 0.00144f
C21240 VGND.n574 0 0.00651f
C21241 VGND.n575 0 0.00261f
C21242 VGND.n576 0 0.00234f
C21243 VGND.n577 0 0.00234f
C21244 VGND.n578 0 0.00225f
C21245 VGND.n579 0 0.00144f
C21246 VGND.n580 0 0.00148f
C21247 VGND.n581 0 8.57e-19
C21248 VGND.n582 0 0.00126f
C21249 VGND.n583 0 0.00135f
C21250 VGND.n584 0 0.00297f
C21251 VGND.n585 0 0.00315f
C21252 VGND.n586 0 0.00207f
C21253 VGND.n587 0 9.9e-19
C21254 VGND.n588 0 0.00261f
C21255 VGND.n589 0 0.00207f
C21256 VGND.n590 0 0.00135f
C21257 VGND.n591 0 7.2e-19
C21258 VGND.n592 0 0.00126f
C21259 VGND.n593 0 0.00414f
C21260 VGND.n594 0 0.00423f
C21261 VGND.n595 0 0.00126f
C21262 VGND.n596 0 0.00912f
C21263 VGND.n597 0 0.0101f
C21264 VGND.n598 0 0.00126f
C21265 VGND.n599 0 0.00824f
C21266 VGND.n600 0 0.00413f
C21267 VGND.n601 0 0.317f
C21268 VGND.n602 0 0.317f
C21269 VGND.n603 0 0.00269f
C21270 VGND.n604 0 0.00207f
C21271 VGND.n605 0 0.00287f
C21272 VGND.n606 0 0.00173f
C21273 VGND.n608 0 0.00274f
C21274 VGND.n609 0 0.00173f
C21275 VGND.n610 0 0.00413f
C21276 VGND.n611 0 0.00207f
C21277 VGND.n612 0 0.00287f
C21278 VGND.n613 0 0.0039f
C21279 VGND.n614 0 0.00269f
C21280 VGND.n615 0 0.00173f
C21281 VGND.n617 0 0.00274f
C21282 VGND.n618 0 0.00173f
C21283 VGND.n619 0 0.00369f
C21284 VGND.n620 0 0.00234f
C21285 VGND.n621 0 7.2e-19
C21286 VGND.n622 0 0.00207f
C21287 VGND.n623 0 0.00207f
C21288 VGND.n624 0 0.00207f
C21289 VGND.n625 0 0.00297f
C21290 VGND.n626 0 0.00234f
C21291 VGND.n627 0 0.00234f
C21292 VGND.n628 0 0.0331f
C21293 VGND.n629 0 0.0367f
C21294 VGND.t337 0 0.128f
C21295 VGND.n630 0 0.154f
C21296 VGND.n631 0 0.0396f
C21297 VGND.n632 0 0.0258f
C21298 VGND.n633 0 0.028f
C21299 VGND.t89 0 0.082f
C21300 VGND.n634 0 0.0934f
C21301 VGND.n635 0 0.0217f
C21302 VGND.n636 0 0.00414f
C21303 VGND.n637 0 0.00423f
C21304 VGND.n638 0 0.00126f
C21305 VGND.t31 0 0.128f
C21306 VGND.n639 0 0.154f
C21307 VGND.n640 0 0.0685f
C21308 VGND.t82 0 0.157f
C21309 VGND.n641 0 0.192f
C21310 VGND.n642 0 0.0321f
C21311 VGND.n643 0 0.0321f
C21312 VGND.t338 0 0.082f
C21313 VGND.n644 0 0.0934f
C21314 VGND.n645 0 0.0157f
C21315 VGND.n646 0 8.1e-19
C21316 VGND.n647 0 7.2e-19
C21317 VGND.t214 0 0.0813f
C21318 VGND.n648 0 0.139f
C21319 VGND.n649 0 0.0166f
C21320 VGND.n650 0 0.0346f
C21321 VGND.t193 0 0.0837f
C21322 VGND.n651 0 0.185f
C21323 VGND.n652 0 0.0166f
C21324 VGND.t308 0 0.124f
C21325 VGND.n653 0 0.225f
C21326 VGND.n654 0 0.038f
C21327 VGND.t165 0 0.0813f
C21328 VGND.n655 0 0.139f
C21329 VGND.n656 0 0.0349f
C21330 VGND.t283 0 0.0812f
C21331 VGND.n657 0 0.139f
C21332 VGND.n658 0 0.00981f
C21333 VGND.n659 0 0.0166f
C21334 VGND.n660 0 0.0438f
C21335 VGND.n661 0 0.0166f
C21336 VGND.t239 0 0.0792f
C21337 VGND.n662 0 0.0367f
C21338 VGND.t181 0 0.128f
C21339 VGND.n663 0 0.154f
C21340 VGND.n664 0 0.0166f
C21341 VGND.n665 0 0.0283f
C21342 VGND.n666 0 0.0166f
C21343 VGND.n667 0 0.0166f
C21344 VGND.n668 0 0.015f
C21345 VGND.t182 0 0.0837f
C21346 VGND.n669 0 0.0222f
C21347 VGND.t309 0 0.0837f
C21348 VGND.n670 0 0.00828f
C21349 VGND.n671 0 0.0267f
C21350 VGND.t166 0 0.0813f
C21351 VGND.n672 0 0.139f
C21352 VGND.n673 0 0.0349f
C21353 VGND.n674 0 0.0159f
C21354 VGND.t284 0 0.0812f
C21355 VGND.n675 0 0.139f
C21356 VGND.t327 0 0.0445f
C21357 VGND.t304 0 0.0445f
C21358 VGND.n676 0 0.243f
C21359 VGND.n677 0 0.0107f
C21360 VGND.n678 0 0.0205f
C21361 VGND.n679 0 0.0165f
C21362 VGND.n680 0 0.00828f
C21363 VGND.n681 0 0.0293f
C21364 VGND.n682 0 0.035f
C21365 VGND.n683 0 0.015f
C21366 VGND.n684 0 0.0166f
C21367 VGND.n685 0 0.00367f
C21368 VGND.n686 0 0.0296f
C21369 VGND.n687 0 0.325f
C21370 VGND.n688 0 0.0285f
C21371 VGND.n689 0 0.0227f
C21372 VGND.n690 0 0.0254f
C21373 VGND.n691 0 0.0044f
C21374 VGND.n692 0 0.0166f
C21375 VGND.n693 0 0.00972f
C21376 VGND.n694 0 0.0151f
C21377 VGND.n695 0 0.0583f
C21378 VGND.n696 0 0.0331f
C21379 VGND.n697 0 0.0273f
C21380 VGND.n698 0 0.0275f
C21381 VGND.n699 0 0.019f
C21382 VGND.n700 0 0.0496f
C21383 VGND.n701 0 0.213f
C21384 VGND.n702 0 0.229f
C21385 VGND.n703 0 0.0252f
C21386 VGND.n704 0 0.009f
C21387 VGND.n705 0 0.0143f
C21388 VGND.n706 0 0.0166f
C21389 VGND.n707 0 0.0331f
C21390 VGND.n708 0 0.0243f
C21391 VGND.n709 0 0.0547f
C21392 VGND.n710 0 0.0366f
C21393 VGND.n711 0 0.00981f
C21394 VGND.n712 0 0.00828f
C21395 VGND.n713 0 0.015f
C21396 VGND.n714 0 0.00708f
C21397 VGND.n715 0 0.0248f
C21398 VGND.n716 0 0.0351f
C21399 VGND.n717 0 0.0107f
C21400 VGND.n718 0 0.00891f
C21401 VGND.n719 0 0.0165f
C21402 VGND.n720 0 0.00828f
C21403 VGND.n721 0 0.0149f
C21404 VGND.n722 0 0.0349f
C21405 VGND.n723 0 0.0349f
C21406 VGND.n724 0 0.038f
C21407 VGND.n725 0 0.00972f
C21408 VGND.n726 0 0.023f
C21409 VGND.n727 0 0.00828f
C21410 VGND.n728 0 0.015f
C21411 VGND.n729 0 0.00613f
C21412 VGND.n730 0 0.0434f
C21413 VGND.n731 0 0.00341f
C21414 VGND.n732 0 0.00963f
C21415 VGND.n733 0 0.00837f
C21416 VGND.n734 0 0.0285f
C21417 VGND.t357 0 0.0812f
C21418 VGND.n735 0 0.139f
C21419 VGND.n736 0 0.0349f
C21420 VGND.n737 0 0.0176f
C21421 VGND.n738 0 0.0119f
C21422 VGND.n739 0 0.00207f
C21423 VGND.n740 0 0.00287f
C21424 VGND.n741 0 0.00173f
C21425 VGND.n742 0 0.00269f
C21426 VGND.n743 0 0.0039f
C21427 VGND.n744 0 0.00269f
C21428 VGND.n745 0 0.00173f
C21429 VGND.n747 0 0.00274f
C21430 VGND.n748 0 0.00173f
C21431 VGND.n749 0 0.00207f
C21432 VGND.n750 0 0.00603f
C21433 VGND.n751 0 0.00234f
C21434 VGND.n752 0 0.00135f
C21435 VGND.n753 0 0.00189f
C21436 VGND.n754 0 0.00369f
C21437 VGND.n755 0 0.00252f
C21438 VGND.n756 0 7.2e-19
C21439 VGND.n757 0 7.2e-19
C21440 VGND.n758 0 0.00162f
C21441 VGND.n759 0 0.0331f
C21442 VGND.n760 0 0.0151f
C21443 VGND.t222 0 0.0799f
C21444 VGND.n761 0 0.0723f
C21445 VGND.n762 0 0.00981f
C21446 VGND.n763 0 0.0327f
C21447 VGND.t334 0 0.0792f
C21448 VGND.n764 0 0.0618f
C21449 VGND.n765 0 0.0283f
C21450 VGND.n766 0 0.0339f
C21451 VGND.n767 0 0.009f
C21452 VGND.n768 0 0.0651f
C21453 VGND.n769 0 0.213f
C21454 VGND.n770 0 0.00456f
C21455 VGND.t12 0 0.0792f
C21456 VGND.n771 0 0.0243f
C21457 VGND.n772 0 0.0658f
C21458 VGND.n773 0 0.0243f
C21459 VGND.n774 0 0.0321f
C21460 VGND.t320 0 0.0812f
C21461 VGND.t135 0 0.128f
C21462 VGND.n775 0 0.198f
C21463 VGND.n776 0 0.0796f
C21464 VGND.n777 0 0.0271f
C21465 VGND.t40 0 0.0946f
C21466 VGND.n778 0 0.0183f
C21467 VGND.n779 0 0.0961f
C21468 VGND.n780 0 0.0252f
C21469 VGND.n781 0 0.0436f
C21470 VGND.n782 0 0.0335f
C21471 VGND.t113 0 0.0792f
C21472 VGND.n783 0 0.054f
C21473 VGND.n784 0 0.0243f
C21474 VGND.n785 0 0.014f
C21475 VGND.n786 0 0.0499f
C21476 VGND.n787 0 0.0166f
C21477 VGND.n788 0 0.015f
C21478 VGND.n789 0 0.0383f
C21479 VGND.n790 0 0.0448f
C21480 VGND.n791 0 0.00972f
C21481 VGND.n792 0 0.0166f
C21482 VGND.n793 0 0.0166f
C21483 VGND.n794 0 0.0345f
C21484 VGND.n795 0 0.0252f
C21485 VGND.n796 0 0.0166f
C21486 VGND.n797 0 0.0316f
C21487 VGND.n798 0 0.0166f
C21488 VGND.n799 0 0.0324f
C21489 VGND.n800 0 0.0166f
C21490 VGND.n801 0 0.0689f
C21491 VGND.n802 0 0.0166f
C21492 VGND.n803 0 0.0144f
C21493 VGND.n804 0 0.0443f
C21494 VGND.n805 0 0.00456f
C21495 VGND.n806 0 0.00891f
C21496 VGND.n807 0 0.0173f
C21497 VGND.n808 0 0.0165f
C21498 VGND.n809 0 0.0628f
C21499 VGND.n810 0 0.139f
C21500 VGND.n811 0 0.0109f
C21501 VGND.n812 0 0.00891f
C21502 VGND.n813 0 0.00981f
C21503 VGND.n814 0 0.0166f
C21504 VGND.n815 0 0.015f
C21505 VGND.n816 0 0.0316f
C21506 VGND.n817 0 0.0428f
C21507 VGND.n818 0 0.00981f
C21508 VGND.n819 0 0.0166f
C21509 VGND.n820 0 0.0331f
C21510 VGND.n821 0 0.0166f
C21511 VGND.n822 0 0.0379f
C21512 VGND.n823 0 0.0144f
C21513 VGND.n824 0 0.00819f
C21514 VGND.n825 0 0.009f
C21515 VGND.t344 0 0.0792f
C21516 VGND.n826 0 0.0284f
C21517 VGND.n827 0 0.074f
C21518 VGND.n828 0 0.0438f
C21519 VGND.t294 0 0.0946f
C21520 VGND.n829 0 0.0183f
C21521 VGND.n830 0 0.0961f
C21522 VGND.n831 0 0.0252f
C21523 VGND.n832 0 0.0271f
C21524 VGND.n833 0 0.0321f
C21525 VGND.t76 0 0.0792f
C21526 VGND.n834 0 0.0604f
C21527 VGND.n835 0 0.0442f
C21528 VGND.n836 0 0.068f
C21529 VGND.n837 0 0.00819f
C21530 VGND.n838 0 0.0428f
C21531 VGND.t321 0 0.0837f
C21532 VGND.t379 0 0.0445f
C21533 VGND.t351 0 0.0445f
C21534 VGND.n839 0 0.243f
C21535 VGND.n840 0 0.032f
C21536 VGND.n841 0 0.0351f
C21537 VGND.t50 0 0.0837f
C21538 VGND.n842 0 0.325f
C21539 VGND.n843 0 0.0424f
C21540 VGND.n844 0 0.015f
C21541 VGND.n845 0 0.0109f
C21542 VGND.n846 0 0.0166f
C21543 VGND.n847 0 0.0166f
C21544 VGND.n848 0 0.00513f
C21545 VGND.n849 0 0.0246f
C21546 VGND.n850 0 0.0686f
C21547 VGND.n851 0 0.0144f
C21548 VGND.n852 0 0.0166f
C21549 VGND.n853 0 0.0166f
C21550 VGND.n854 0 0.00981f
C21551 VGND.n855 0 0.0488f
C21552 VGND.n856 0 0.0353f
C21553 VGND.n857 0 0.0242f
C21554 VGND.n858 0 0.015f
C21555 VGND.n859 0 0.0166f
C21556 VGND.n860 0 0.0166f
C21557 VGND.n861 0 0.00981f
C21558 VGND.n862 0 0.0445f
C21559 VGND.n863 0 0.0379f
C21560 VGND.n864 0 0.015f
C21561 VGND.n865 0 0.0239f
C21562 VGND.n866 0 0.0166f
C21563 VGND.n867 0 0.00981f
C21564 VGND.n868 0 0.0339f
C21565 VGND.n869 0 0.0371f
C21566 VGND.n870 0 0.015f
C21567 VGND.n871 0 0.0331f
C21568 VGND.n872 0 0.0166f
C21569 VGND.n873 0 0.0166f
C21570 VGND.n874 0 0.00981f
C21571 VGND.n875 0 0.0279f
C21572 VGND.n876 0 0.0261f
C21573 VGND.n877 0 0.0945f
C21574 VGND.n878 0 8.1e-19
C21575 VGND.n879 0 0.00198f
C21576 VGND.n880 0 1.46e-19
C21577 VGND.n881 0 0.00185f
C21578 VGND.n882 0 9.77e-19
C21579 VGND.n883 0 0.0298f
C21580 VGND.n884 0 0.229f
C21581 VGND.n885 0 0.0299f
C21582 VGND.t323 0 0.0818f
C21583 VGND.n886 0 0.139f
C21584 VGND.t363 0 0.082f
C21585 VGND.n887 0 0.00549f
C21586 VGND.t364 0 0.0799f
C21587 VGND.n888 0 0.0723f
C21588 VGND.t204 0 0.128f
C21589 VGND.n889 0 0.198f
C21590 VGND.n890 0 0.00234f
C21591 VGND.n891 0 0.00369f
C21592 VGND.n892 0 0.00234f
C21593 VGND.n893 0 7.2e-19
C21594 VGND.n894 0 0.00207f
C21595 VGND.n895 0 0.00207f
C21596 VGND.n896 0 0.00207f
C21597 VGND.n897 0 0.00297f
C21598 VGND.n898 0 0.00234f
C21599 VGND.n899 0 0.00274f
C21600 VGND.n900 0 0.00173f
C21601 VGND.n901 0 0.00234f
C21602 VGND.t18 0 0.0792f
C21603 VGND.n902 0 0.0243f
C21604 VGND.n903 0 0.0547f
C21605 VGND.t183 0 0.0792f
C21606 VGND.n904 0 0.0421f
C21607 VGND.n905 0 0.0555f
C21608 VGND.n906 0 0.0321f
C21609 VGND.t184 0 0.121f
C21610 VGND.n907 0 0.0597f
C21611 VGND.n908 0 0.138f
C21612 VGND.n909 0 0.0143f
C21613 VGND.n910 0 0.0166f
C21614 VGND.n911 0 0.0166f
C21615 VGND.n912 0 0.00981f
C21616 VGND.n913 0 0.0643f
C21617 VGND.n914 0 0.0271f
C21618 VGND.t19 0 0.0946f
C21619 VGND.n915 0 0.0183f
C21620 VGND.n916 0 0.0961f
C21621 VGND.n917 0 0.0449f
C21622 VGND.n918 0 0.0341f
C21623 VGND.n919 0 0.0345f
C21624 VGND.n920 0 0.0242f
C21625 VGND.n921 0 0.00837f
C21626 VGND.n922 0 0.0149f
C21627 VGND.n923 0 0.0166f
C21628 VGND.n924 0 0.00981f
C21629 VGND.n925 0 0.0452f
C21630 VGND.n926 0 0.00585f
C21631 VGND.n927 0 0.015f
C21632 VGND.n928 0 0.0436f
C21633 VGND.n929 0 0.0166f
C21634 VGND.n930 0 0.0116f
C21635 VGND.n931 0 0.0166f
C21636 VGND.n932 0 0.0379f
C21637 VGND.n933 0 0.0166f
C21638 VGND.n934 0 0.0331f
C21639 VGND.n935 0 0.0166f
C21640 VGND.n936 0 0.0166f
C21641 VGND.n937 0 0.00981f
C21642 VGND.n938 0 0.0287f
C21643 VGND.n939 0 0.0388f
C21644 VGND.n940 0 0.015f
C21645 VGND.n941 0 0.0548f
C21646 VGND.n942 0 0.0166f
C21647 VGND.n943 0 0.0166f
C21648 VGND.n944 0 0.00981f
C21649 VGND.n945 0 0.0291f
C21650 VGND.n946 0 0.00549f
C21651 VGND.n947 0 0.015f
C21652 VGND.n948 0 0.01f
C21653 VGND.n949 0 0.0166f
C21654 VGND.n950 0 0.0409f
C21655 VGND.n951 0 0.0166f
C21656 VGND.n952 0 0.0336f
C21657 VGND.n953 0 0.0166f
C21658 VGND.n954 0 0.00981f
C21659 VGND.n955 0 0.0045f
C21660 VGND.n956 0 0.0379f
C21661 VGND.n957 0 0.015f
C21662 VGND.n958 0 0.0331f
C21663 VGND.n959 0 0.0166f
C21664 VGND.t285 0 0.0792f
C21665 VGND.n960 0 0.0516f
C21666 VGND.n961 0 0.0414f
C21667 VGND.n962 0 0.0153f
C21668 VGND.n963 0 0.0127f
C21669 VGND.n964 0 0.00828f
C21670 VGND.n965 0 0.00153f
C21671 VGND.n966 0 0.00304f
C21672 VGND.t386 0 0.0812f
C21673 VGND.n967 0 0.139f
C21674 VGND.n968 0 0.0628f
C21675 VGND.n969 0 7.62e-19
C21676 VGND.n970 0 0.00376f
C21677 VGND.n971 0 0.00234f
C21678 VGND.n972 0 0.00234f
C21679 VGND.n973 0 0.00225f
C21680 VGND.n974 0 0.00144f
C21681 VGND.n975 0 0.00148f
C21682 VGND.n976 0 8.57e-19
C21683 VGND.n977 0 0.00126f
C21684 VGND.n978 0 0.00135f
C21685 VGND.n979 0 0.00297f
C21686 VGND.n980 0 0.00315f
C21687 VGND.n981 0 0.00207f
C21688 VGND.n982 0 9.9e-19
C21689 VGND.n983 0 0.00261f
C21690 VGND.n984 0 0.00207f
C21691 VGND.n985 0 0.00135f
C21692 VGND.n986 0 7.2e-19
C21693 VGND.n987 0 0.00126f
C21694 VGND.n988 0 0.00414f
C21695 VGND.n989 0 0.00423f
C21696 VGND.n990 0 0.00117f
C21697 VGND.n991 0 0.00912f
C21698 VGND.n992 0 0.0101f
C21699 VGND.n993 0 0.00126f
C21700 VGND.n994 0 0.00824f
C21701 VGND.n995 0 0.00413f
C21702 VGND.n996 0 0.192f
C21703 VGND.n997 0 0.00269f
C21704 VGND.n998 0 0.00207f
C21705 VGND.n999 0 0.00287f
C21706 VGND.n1000 0 0.00173f
C21707 VGND.n1002 0 0.00274f
C21708 VGND.n1003 0 0.00173f
C21709 VGND.n1004 0 0.00413f
C21710 VGND.n1005 0 0.00207f
C21711 VGND.n1006 0 0.00287f
C21712 VGND.n1007 0 0.0039f
C21713 VGND.n1008 0 0.00269f
C21714 VGND.n1009 0 0.00173f
C21715 VGND.n1011 0 0.00274f
C21716 VGND.n1012 0 0.00173f
C21717 VGND.n1013 0 0.00369f
C21718 VGND.n1014 0 0.00234f
C21719 VGND.n1015 0 7.2e-19
C21720 VGND.n1016 0 0.00207f
C21721 VGND.n1017 0 0.00207f
C21722 VGND.n1018 0 0.00207f
C21723 VGND.n1019 0 0.00297f
C21724 VGND.n1020 0 0.00234f
C21725 VGND.n1021 0 0.00234f
C21726 VGND.n1022 0 0.0258f
C21727 VGND.n1023 0 0.0348f
C21728 VGND.n1024 0 0.051f
C21729 VGND.n1025 0 0.0277f
C21730 VGND.n1026 0 0.0253f
C21731 VGND.n1027 0 0.00837f
C21732 VGND.n1028 0 0.00414f
C21733 VGND.n1029 0 0.00423f
C21734 VGND.n1030 0 0.00126f
C21735 VGND.t170 0 0.128f
C21736 VGND.n1031 0 0.154f
C21737 VGND.n1032 0 0.0263f
C21738 VGND.n1033 0 0.0521f
C21739 VGND.n1034 0 0.0339f
C21740 VGND.t236 0 0.0946f
C21741 VGND.n1035 0 0.0183f
C21742 VGND.n1036 0 0.0961f
C21743 VGND.n1037 0 0.0252f
C21744 VGND.n1038 0 0.0271f
C21745 VGND.n1039 0 0.0492f
C21746 VGND.n1040 0 0.046f
C21747 VGND.n1041 0 0.138f
C21748 VGND.n1042 0 0.0463f
C21749 VGND.t358 0 0.082f
C21750 VGND.n1043 0 0.0934f
C21751 VGND.n1044 0 0.00463f
C21752 VGND.t51 0 0.128f
C21753 VGND.n1045 0 0.154f
C21754 VGND.n1046 0 0.0516f
C21755 VGND.n1047 0 9.9e-19
C21756 VGND.n1048 0 0.00162f
C21757 VGND.n1049 0 9e-19
C21758 VGND.n1050 0 0.213f
C21759 VGND.t221 0 0.0837f
C21760 VGND.n1051 0 0.186f
C21761 VGND.t220 0 0.0816f
C21762 VGND.n1052 0 0.139f
C21763 VGND.n1053 0 0.00828f
C21764 VGND.n1054 0 0.00408f
C21765 VGND.t331 0 0.0812f
C21766 VGND.n1055 0 0.139f
C21767 VGND.t291 0 0.0445f
C21768 VGND.t263 0 0.0445f
C21769 VGND.n1056 0 0.243f
C21770 VGND.n1057 0 0.0159f
C21771 VGND.n1058 0 0.0107f
C21772 VGND.n1059 0 0.0205f
C21773 VGND.n1060 0 0.0165f
C21774 VGND.n1061 0 0.0349f
C21775 VGND.t192 0 0.0813f
C21776 VGND.n1062 0 0.139f
C21777 VGND.n1063 0 0.0407f
C21778 VGND.n1064 0 0.00828f
C21779 VGND.n1065 0 0.00819f
C21780 VGND.n1066 0 0.0549f
C21781 VGND.n1067 0 0.0378f
C21782 VGND.n1068 0 0.0151f
C21783 VGND.n1069 0 0.0453f
C21784 VGND.n1070 0 0.0221f
C21785 VGND.t382 0 0.082f
C21786 VGND.n1071 0 0.0934f
C21787 VGND.n1072 0 0.0217f
C21788 VGND.n1073 0 0.0137f
C21789 VGND.n1074 0 0.00828f
C21790 VGND.n1075 0 0.0472f
C21791 VGND.n1076 0 0.0324f
C21792 VGND.n1077 0 0.015f
C21793 VGND.n1078 0 0.0236f
C21794 VGND.n1079 0 0.0166f
C21795 VGND.n1080 0 0.0106f
C21796 VGND.n1081 0 0.00549f
C21797 VGND.n1082 0 0.0379f
C21798 VGND.n1083 0 0.0142f
C21799 VGND.n1084 0 0.0331f
C21800 VGND.n1085 0 0.0166f
C21801 VGND.n1086 0 0.0166f
C21802 VGND.n1087 0 0.0506f
C21803 VGND.t360 0 0.163f
C21804 VGND.n1088 0 0.231f
C21805 VGND.n1089 0 0.0277f
C21806 VGND.n1090 0 0.00981f
C21807 VGND.n1091 0 0.023f
C21808 VGND.n1092 0 0.009f
C21809 VGND.t297 0 0.0792f
C21810 VGND.n1093 0 0.0243f
C21811 VGND.n1094 0 0.0547f
C21812 VGND.n1095 0 0.00828f
C21813 VGND.n1096 0 0.00828f
C21814 VGND.t359 0 0.082f
C21815 VGND.n1097 0 0.0934f
C21816 VGND.n1098 0 0.015f
C21817 VGND.n1099 0 0.0217f
C21818 VGND.t203 0 0.0816f
C21819 VGND.n1100 0 0.139f
C21820 VGND.n1101 0 0.00828f
C21821 VGND.t15 0 0.0792f
C21822 VGND.n1102 0 0.0407f
C21823 VGND.n1103 0 0.0547f
C21824 VGND.n1104 0 0.00837f
C21825 VGND.n1105 0 0.0357f
C21826 VGND.n1106 0 0.00207f
C21827 VGND.n1107 0 0.00207f
C21828 VGND.n1108 0 0.00287f
C21829 VGND.n1109 0 0.00173f
C21830 VGND.n1110 0 0.00269f
C21831 VGND.n1111 0 0.0039f
C21832 VGND.n1112 0 0.00269f
C21833 VGND.n1113 0 0.00173f
C21834 VGND.n1115 0 0.00274f
C21835 VGND.n1116 0 0.00173f
C21836 VGND.n1117 0 0.00207f
C21837 VGND.n1118 0 0.00603f
C21838 VGND.n1119 0 0.00234f
C21839 VGND.n1120 0 0.00135f
C21840 VGND.n1121 0 0.00189f
C21841 VGND.n1122 0 0.00369f
C21842 VGND.n1123 0 0.00252f
C21843 VGND.n1124 0 7.2e-19
C21844 VGND.n1125 0 7.2e-19
C21845 VGND.n1126 0 0.00162f
C21846 VGND.n1127 0 0.0245f
C21847 VGND.n1128 0 0.00545f
C21848 VGND.n1129 0 0.0093f
C21849 VGND.t2 0 0.161f
C21850 VGND.n1130 0 0.234f
C21851 VGND.n1131 0 0.0418f
C21852 VGND.n1132 0 0.0331f
C21853 VGND.n1133 0 0.0254f
C21854 VGND.n1134 0 0.0334f
C21855 VGND.n1135 0 0.0259f
C21856 VGND.n1136 0 0.0331f
C21857 VGND.n1137 0 0.053f
C21858 VGND.n1138 0 0.0423f
C21859 VGND.n1139 0 0.213f
C21860 VGND.n1140 0 0.0279f
C21861 VGND.n1141 0 0.0166f
C21862 VGND.n1142 0 0.00645f
C21863 VGND.n1143 0 0.0166f
C21864 VGND.n1144 0 0.035f
C21865 VGND.n1145 0 0.015f
C21866 VGND.t0 0 0.0792f
C21867 VGND.n1146 0 0.0623f
C21868 VGND.n1147 0 0.015f
C21869 VGND.t150 0 0.158f
C21870 VGND.n1148 0 0.185f
C21871 VGND.n1149 0 0.0649f
C21872 VGND.t356 0 0.0812f
C21873 VGND.n1150 0 0.139f
C21874 VGND.t336 0 0.0445f
C21875 VGND.t317 0 0.0445f
C21876 VGND.n1151 0 0.244f
C21877 VGND.n1152 0 0.0159f
C21878 VGND.n1153 0 0.0205f
C21879 VGND.n1154 0 0.00402f
C21880 VGND.n1155 0 0.0116f
C21881 VGND.n1156 0 0.00846f
C21882 VGND.n1157 0 0.0162f
C21883 VGND.n1158 0 0.077f
C21884 VGND.n1159 0 0.0628f
C21885 VGND.n1160 0 0.0723f
C21886 VGND.n1161 0 0.0208f
C21887 VGND.n1162 0 0.0213f
C21888 VGND.n1163 0 0.0563f
C21889 VGND.n1164 0 0.0243f
C21890 VGND.n1165 0 0.0166f
C21891 VGND.n1166 0 0.00981f
C21892 VGND.n1167 0 0.0373f
C21893 VGND.n1168 0 0.0059f
C21894 VGND.n1169 0 0.0242f
C21895 VGND.n1170 0 0.0166f
C21896 VGND.n1171 0 0.0166f
C21897 VGND.n1172 0 0.0166f
C21898 VGND.n1173 0 0.0132f
C21899 VGND.n1174 0 0.00586f
C21900 VGND.n1175 0 0.024f
C21901 VGND.n1176 0 0.0166f
C21902 VGND.n1177 0 0.00981f
C21903 VGND.n1178 0 0.015f
C21904 VGND.n1179 0 0.0566f
C21905 VGND.n1180 0 0.0331f
C21906 VGND.t1 0 0.0792f
C21907 VGND.n1181 0 0.0658f
C21908 VGND.n1182 0 0.04f
C21909 VGND.n1183 0 0.0166f
C21910 VGND.n1184 0 0.00981f
C21911 VGND.n1185 0 0.009f
C21912 VGND.n1186 0 0.0336f
C21913 VGND.n1187 0 0.00981f
C21914 VGND.t63 0 0.0792f
C21915 VGND.n1188 0 0.00837f
C21916 VGND.n1189 0 0.00819f
C21917 VGND.n1190 0 0.0554f
C21918 VGND.n1191 0 0.0166f
C21919 VGND.n1192 0 0.0391f
C21920 VGND.t178 0 0.157f
C21921 VGND.n1193 0 0.2f
C21922 VGND.n1194 0 0.0496f
C21923 VGND.t49 0 0.0813f
C21924 VGND.n1195 0 0.139f
C21925 VGND.n1196 0 0.0109f
C21926 VGND.n1197 0 0.031f
C21927 VGND.n1198 0 0.0166f
C21928 VGND.n1199 0 0.0326f
C21929 VGND.n1200 0 0.0166f
C21930 VGND.t164 0 0.0792f
C21931 VGND.n1201 0 0.067f
C21932 VGND.n1202 0 0.0442f
C21933 VGND.n1203 0 0.014f
C21934 VGND.n1204 0 0.0604f
C21935 VGND.n1205 0 0.0166f
C21936 VGND.n1206 0 0.069f
C21937 VGND.n1207 0 0.0151f
C21938 VGND.n1208 0 0.00972f
C21939 VGND.n1209 0 0.00344f
C21940 VGND.n1210 0 0.034f
C21941 VGND.n1211 0 0.0248f
C21942 VGND.n1212 0 0.0166f
C21943 VGND.n1213 0 0.0166f
C21944 VGND.n1214 0 0.0166f
C21945 VGND.n1215 0 0.0406f
C21946 VGND.n1216 0 0.00564f
C21947 VGND.n1217 0 0.00398f
C21948 VGND.n1218 0 0.0166f
C21949 VGND.n1219 0 0.015f
C21950 VGND.n1220 0 0.00828f
C21951 VGND.n1221 0 0.019f
C21952 VGND.n1222 0 0.0414f
C21953 VGND.n1223 0 0.0166f
C21954 VGND.n1224 0 0.0296f
C21955 VGND.n1225 0 0.0324f
C21956 VGND.n1226 0 0.058f
C21957 VGND.n1227 0 0.0166f
C21958 VGND.n1228 0 0.0144f
C21959 VGND.n1229 0 0.00891f
C21960 VGND.n1230 0 0.00386f
C21961 VGND.n1231 0 0.0299f
C21962 VGND.n1232 0 0.00574f
C21963 VGND.n1233 0 0.0278f
C21964 VGND.n1234 0 0.0547f
C21965 VGND.n1235 0 0.0457f
C21966 VGND.n1236 0 0.0166f
C21967 VGND.n1237 0 0.0166f
C21968 VGND.n1238 0 0.0143f
C21969 VGND.n1239 0 0.0367f
C21970 VGND.n1240 0 0.026f
C21971 VGND.n1241 0 0.229f
C21972 VGND.n1242 0 8.1e-19
C21973 VGND.n1243 0 0.00198f
C21974 VGND.n1244 0 1.46e-19
C21975 VGND.n1245 0 0.00185f
C21976 VGND.n1246 0 9.77e-19
C21977 VGND.n1247 0 0.0316f
C21978 VGND.n1248 0 0.184f
C21979 VGND.n1249 0 0.229f
C21980 VGND.t13 0 0.0792f
C21981 VGND.n1250 0 0.0243f
C21982 VGND.n1251 0 0.0547f
C21983 VGND.n1252 0 0.053f
C21984 VGND.t93 0 0.0792f
C21985 VGND.n1253 0 0.0245f
C21986 VGND.n1254 0 0.0567f
C21987 VGND.n1255 0 0.0343f
C21988 VGND.t42 0 0.0792f
C21989 VGND.t126 0 0.0792f
C21990 VGND.n1256 0 0.0243f
C21991 VGND.n1257 0 0.0547f
C21992 VGND.n1258 0 0.0231f
C21993 VGND.n1259 0 0.00126f
C21994 VGND.n1260 0 0.00274f
C21995 VGND.n1261 0 0.00173f
C21996 VGND.n1262 0 0.00413f
C21997 VGND.n1263 0 0.00261f
C21998 VGND.n1264 0 0.00207f
C21999 VGND.n1265 0 0.00135f
C22000 VGND.n1266 0 0.00423f
C22001 VGND.n1267 0 0.00414f
C22002 VGND.n1268 0 0.00148f
C22003 VGND.n1269 0 0.0519f
C22004 VGND.t34 0 0.124f
C22005 VGND.n1270 0 0.225f
C22006 VGND.t26 0 0.082f
C22007 VGND.n1271 0 0.0907f
C22008 VGND.n1272 0 0.015f
C22009 VGND.n1273 0 0.0524f
C22010 VGND.n1274 0 0.0166f
C22011 VGND.n1275 0 0.0508f
C22012 VGND.n1276 0 0.00828f
C22013 VGND.n1277 0 0.00153f
C22014 VGND.n1278 0 0.00369f
C22015 VGND.n1279 0 0.00144f
C22016 VGND.n1280 0 0.00225f
C22017 VGND.n1281 0 0.00247f
C22018 VGND.n1282 0 0.0345f
C22019 VGND.n1283 0 8.41e-19
C22020 VGND.n1284 0 0.00371f
C22021 VGND.n1285 0 0.00234f
C22022 VGND.n1286 0 0.00234f
C22023 VGND.n1287 0 0.00234f
C22024 VGND.n1288 0 7.2e-19
C22025 VGND.n1289 0 0.00207f
C22026 VGND.n1290 0 0.00207f
C22027 VGND.n1291 0 0.00207f
C22028 VGND.n1292 0 0.00297f
C22029 VGND.n1293 0 0.00234f
C22030 VGND.n1294 0 0.317f
C22031 VGND.n1295 0 0.317f
C22032 VGND.n1296 0 0.00269f
C22033 VGND.n1297 0 0.00207f
C22034 VGND.n1298 0 0.00287f
C22035 VGND.n1299 0 0.00173f
C22036 VGND.n1301 0 0.00274f
C22037 VGND.n1302 0 0.00173f
C22038 VGND.n1303 0 0.00413f
C22039 VGND.n1304 0 0.00207f
C22040 VGND.n1305 0 0.00287f
C22041 VGND.n1306 0 0.0039f
C22042 VGND.n1307 0 0.00269f
C22043 VGND.n1308 0 0.00173f
C22044 VGND.n1310 0 0.00274f
C22045 VGND.n1311 0 0.00173f
C22046 VGND.n1312 0 0.00369f
C22047 VGND.n1313 0 0.00234f
C22048 VGND.n1314 0 7.2e-19
C22049 VGND.n1315 0 0.00207f
C22050 VGND.n1316 0 0.00207f
C22051 VGND.n1317 0 0.00207f
C22052 VGND.n1318 0 0.00297f
C22053 VGND.n1319 0 0.00234f
C22054 VGND.n1320 0 0.00234f
C22055 VGND.n1321 0 0.0217f
C22056 VGND.n1322 0 0.00376f
C22057 VGND.t372 0 0.0816f
C22058 VGND.n1323 0 0.139f
C22059 VGND.n1324 0 0.043f
C22060 VGND.n1325 0 0.0387f
C22061 VGND.n1326 0 0.0378f
C22062 VGND.n1327 0 0.0107f
C22063 VGND.t70 0 0.0837f
C22064 VGND.n1328 0 0.185f
C22065 VGND.n1329 0 0.0166f
C22066 VGND.n1330 0 0.153f
C22067 VGND.n1331 0 0.0499f
C22068 VGND.n1332 0 0.0425f
C22069 VGND.n1333 0 0.00981f
C22070 VGND.n1334 0 0.00414f
C22071 VGND.t391 0 0.0792f
C22072 VGND.n1335 0 0.0243f
C22073 VGND.n1336 0 0.0547f
C22074 VGND.n1337 0 0.0291f
C22075 VGND.t340 0 0.0813f
C22076 VGND.n1338 0 0.139f
C22077 VGND.n1339 0 0.0349f
C22078 VGND.n1340 0 0.0279f
C22079 VGND.n1341 0 8.1e-19
C22080 VGND.n1342 0 0.00387f
C22081 VGND.n1343 0 7.2e-19
C22082 VGND.t252 0 0.0792f
C22083 VGND.n1344 0 0.0243f
C22084 VGND.n1345 0 0.0623f
C22085 VGND.n1346 0 0.04f
C22086 VGND.t251 0 0.0837f
C22087 VGND.n1347 0 0.186f
C22088 VGND.n1348 0 0.0166f
C22089 VGND.n1349 0 0.0596f
C22090 VGND.n1350 0 0.0143f
C22091 VGND.n1351 0 0.0279f
C22092 VGND.n1352 0 0.213f
C22093 VGND.n1353 0 0.138f
C22094 VGND.n1354 0 0.0166f
C22095 VGND.n1355 0 0.00645f
C22096 VGND.n1356 0 0.0166f
C22097 VGND.n1357 0 0.035f
C22098 VGND.n1358 0 0.015f
C22099 VGND.t143 0 0.0792f
C22100 VGND.n1359 0 0.0623f
C22101 VGND.n1360 0 0.015f
C22102 VGND.t292 0 0.158f
C22103 VGND.n1361 0 0.185f
C22104 VGND.n1362 0 0.0458f
C22105 VGND.n1363 0 0.015f
C22106 VGND.t120 0 0.082f
C22107 VGND.n1364 0 0.0934f
C22108 VGND.n1365 0 0.0266f
C22109 VGND.t246 0 0.0445f
C22110 VGND.n1366 0 0.0159f
C22111 VGND.t368 0 0.0445f
C22112 VGND.n1367 0 0.244f
C22113 VGND.n1368 0 0.0367f
C22114 VGND.n1369 0 0.028f
C22115 VGND.n1370 0 0.0106f
C22116 VGND.n1371 0 0.011f
C22117 VGND.n1372 0 0.045f
C22118 VGND.n1373 0 0.0801f
C22119 VGND.n1374 0 0.0292f
C22120 VGND.n1375 0 0.0221f
C22121 VGND.n1376 0 0.011f
C22122 VGND.n1377 0 0.0473f
C22123 VGND.n1378 0 0.00891f
C22124 VGND.n1379 0 0.00765f
C22125 VGND.n1380 0 0.0213f
C22126 VGND.n1381 0 0.0563f
C22127 VGND.n1382 0 0.0243f
C22128 VGND.n1383 0 0.0166f
C22129 VGND.n1384 0 0.00981f
C22130 VGND.n1385 0 0.0373f
C22131 VGND.n1386 0 0.0059f
C22132 VGND.n1387 0 0.0242f
C22133 VGND.n1388 0 0.0166f
C22134 VGND.n1389 0 0.0166f
C22135 VGND.n1390 0 0.0166f
C22136 VGND.n1391 0 0.0132f
C22137 VGND.n1392 0 0.00586f
C22138 VGND.n1393 0 0.024f
C22139 VGND.n1394 0 0.0166f
C22140 VGND.n1395 0 0.00981f
C22141 VGND.n1396 0 0.015f
C22142 VGND.n1397 0 0.0566f
C22143 VGND.n1398 0 0.0331f
C22144 VGND.t144 0 0.0792f
C22145 VGND.n1399 0 0.0658f
C22146 VGND.n1400 0 0.04f
C22147 VGND.n1401 0 0.0166f
C22148 VGND.n1402 0 0.00981f
C22149 VGND.n1403 0 0.009f
C22150 VGND.n1404 0 0.0261f
C22151 VGND.n1405 0 0.00494f
C22152 VGND.n1406 0 0.00547f
C22153 VGND.n1407 0 0.0106f
C22154 VGND.n1408 0 0.0142f
C22155 VGND.n1409 0 0.0166f
C22156 VGND.n1410 0 0.0333f
C22157 VGND.n1411 0 0.0499f
C22158 VGND.t145 0 0.163f
C22159 VGND.n1412 0 0.228f
C22160 VGND.n1413 0 0.0196f
C22161 VGND.n1414 0 0.00981f
C22162 VGND.n1415 0 0.023f
C22163 VGND.n1416 0 0.00828f
C22164 VGND.n1417 0 0.0466f
C22165 VGND.n1418 0 0.00223f
C22166 VGND.n1419 0 0.015f
C22167 VGND.n1420 0 0.0234f
C22168 VGND.n1421 0 0.0166f
C22169 VGND.n1422 0 0.00567f
C22170 VGND.n1423 0 0.0166f
C22171 VGND.n1424 0 0.0058f
C22172 VGND.n1425 0 0.0166f
C22173 VGND.n1426 0 0.0585f
C22174 VGND.n1427 0 0.0166f
C22175 VGND.n1428 0 0.0132f
C22176 VGND.n1429 0 0.0166f
C22177 VGND.n1430 0 0.0379f
C22178 VGND.n1431 0 0.0166f
C22179 VGND.n1432 0 0.0331f
C22180 VGND.n1433 0 0.0166f
C22181 VGND.n1434 0 0.0166f
C22182 VGND.n1435 0 0.00981f
C22183 VGND.n1436 0 0.00828f
C22184 VGND.n1437 0 0.0337f
C22185 VGND.n1438 0 0.0215f
C22186 VGND.n1439 0 0.015f
C22187 VGND.n1440 0 0.0423f
C22188 VGND.n1441 0 0.0166f
C22189 VGND.n1442 0 0.0373f
C22190 VGND.n1443 0 0.0166f
C22191 VGND.n1444 0 0.0331f
C22192 VGND.n1445 0 0.0166f
C22193 VGND.t307 0 0.0792f
C22194 VGND.n1446 0 0.0536f
C22195 VGND.n1447 0 0.0243f
C22196 VGND.n1448 0 0.014f
C22197 VGND.n1449 0 0.00603f
C22198 VGND.n1450 0 0.206f
C22199 VGND.n1451 0 0.00274f
C22200 VGND.n1452 0 0.00173f
C22201 VGND.n1453 0 0.00413f
C22202 VGND.n1454 0 0.00207f
C22203 VGND.n1455 0 0.00287f
C22204 VGND.n1456 0 0.00269f
C22205 VGND.n1457 0 0.00173f
C22206 VGND.n1459 0 0.00274f
C22207 VGND.n1460 0 0.00173f
C22208 VGND.n1461 0 0.00234f
C22209 VGND.t91 0 0.128f
C22210 VGND.n1462 0 0.154f
C22211 VGND.n1463 0 0.0519f
C22212 VGND.n1464 0 0.0291f
C22213 VGND.n1465 0 0.0254f
C22214 VGND.n1466 0 0.0239f
C22215 VGND.n1467 0 0.0236f
C22216 VGND.n1468 0 0.059f
C22217 VGND.n1469 0 0.0597f
C22218 VGND.n1470 0 0.0878f
C22219 VGND.t172 0 0.0946f
C22220 VGND.n1471 0 0.0192f
C22221 VGND.n1472 0 0.0961f
C22222 VGND.n1473 0 0.0309f
C22223 VGND.n1474 0 0.0271f
C22224 VGND.n1475 0 0.0321f
C22225 VGND.n1476 0 0.0653f
C22226 VGND.n1477 0 0.0331f
C22227 VGND.n1478 0 0.00414f
C22228 VGND.t257 0 0.0792f
C22229 VGND.n1479 0 0.0243f
C22230 VGND.n1480 0 0.0547f
C22231 VGND.n1481 0 0.0291f
C22232 VGND.t75 0 0.128f
C22233 VGND.n1482 0 0.154f
C22234 VGND.n1483 0 0.0766f
C22235 VGND.n1484 0 0.0404f
C22236 VGND.n1485 0 0.0324f
C22237 VGND.n1486 0 0.094f
C22238 VGND.n1487 0 0.009f
C22239 VGND.t256 0 0.082f
C22240 VGND.n1488 0 0.0938f
C22241 VGND.n1489 0 0.028f
C22242 VGND.t228 0 0.128f
C22243 VGND.n1490 0 0.198f
C22244 VGND.n1491 0 0.0119f
C22245 VGND.t148 0 0.156f
C22246 VGND.n1492 0 0.198f
C22247 VGND.n1493 0 0.0788f
C22248 VGND.n1494 0 0.0192f
C22249 VGND.n1495 0 0.0559f
C22250 VGND.n1496 0 0.00287f
C22251 VGND.n1497 0 0.00207f
C22252 VGND.n1498 0 0.00274f
C22253 VGND.n1499 0 0.317f
C22254 VGND.n1500 0 0.317f
C22255 VGND.n1501 0 0.00207f
C22256 VGND.n1502 0 0.00287f
C22257 VGND.n1503 0 0.00173f
C22258 VGND.n1504 0 0.00269f
C22259 VGND.n1505 0 0.0039f
C22260 VGND.n1506 0 0.00269f
C22261 VGND.n1507 0 0.00173f
C22262 VGND.n1509 0 0.00274f
C22263 VGND.n1510 0 0.00173f
C22264 VGND.n1511 0 0.00207f
C22265 VGND.n1512 0 0.00603f
C22266 VGND.n1513 0 0.00234f
C22267 VGND.n1514 0 0.00135f
C22268 VGND.n1515 0 0.00189f
C22269 VGND.n1516 0 0.00369f
C22270 VGND.n1517 0 0.00252f
C22271 VGND.n1518 0 7.2e-19
C22272 VGND.n1519 0 7.2e-19
C22273 VGND.n1520 0 0.00162f
C22274 VGND.n1521 0 0.00549f
C22275 VGND.n1522 0 0.0444f
C22276 VGND.t158 0 0.128f
C22277 VGND.n1523 0 0.154f
C22278 VGND.n1524 0 0.0295f
C22279 VGND.n1525 0 0.0564f
C22280 VGND.n1526 0 0.0351f
C22281 VGND.n1527 0 0.0655f
C22282 VGND.t348 0 0.128f
C22283 VGND.n1528 0 0.154f
C22284 VGND.n1529 0 0.0257f
C22285 VGND.n1530 0 0.0409f
C22286 VGND.n1531 0 0.0246f
C22287 VGND.n1532 0 0.0367f
C22288 VGND.n1533 0 0.213f
C22289 VGND.n1534 0 0.0223f
C22290 VGND.t56 0 0.155f
C22291 VGND.n1535 0 0.0449f
C22292 VGND.n1536 0 0.163f
C22293 VGND.n1537 0 0.0443f
C22294 VGND.n1538 0 0.0488f
C22295 VGND.n1539 0 0.0365f
C22296 VGND.t104 0 0.0837f
C22297 VGND.n1540 0 0.0538f
C22298 VGND.n1541 0 0.0417f
C22299 VGND.n1542 0 0.037f
C22300 VGND.n1543 0 0.015f
C22301 VGND.n1544 0 0.0166f
C22302 VGND.n1545 0 0.0166f
C22303 VGND.n1546 0 0.0318f
C22304 VGND.t188 0 0.0816f
C22305 VGND.n1547 0 0.139f
C22306 VGND.n1548 0 0.0387f
C22307 VGND.n1549 0 0.022f
C22308 VGND.t209 0 0.0792f
C22309 VGND.n1550 0 0.0732f
C22310 VGND.n1551 0 0.0284f
C22311 VGND.n1552 0 0.014f
C22312 VGND.n1553 0 0.0331f
C22313 VGND.n1554 0 0.0166f
C22314 VGND.n1555 0 0.0379f
C22315 VGND.n1556 0 0.0166f
C22316 VGND.n1557 0 0.00549f
C22317 VGND.n1558 0 0.0166f
C22318 VGND.n1559 0 0.0282f
C22319 VGND.n1560 0 0.0166f
C22320 VGND.n1561 0 0.0229f
C22321 VGND.n1562 0 0.0166f
C22322 VGND.n1563 0 0.00619f
C22323 VGND.n1564 0 0.015f
C22324 VGND.n1565 0 0.00828f
C22325 VGND.n1566 0 0.0119f
C22326 VGND.n1567 0 0.0137f
C22327 VGND.t96 0 0.151f
C22328 VGND.n1568 0 0.126f
C22329 VGND.n1569 0 0.0297f
C22330 VGND.n1570 0 0.0252f
C22331 VGND.n1571 0 0.0901f
C22332 VGND.n1572 0 0.02f
C22333 VGND.n1573 0 0.0221f
C22334 VGND.n1574 0 0.015f
C22335 VGND.n1575 0 0.0558f
C22336 VGND.n1576 0 0.0176f
C22337 VGND.n1577 0 0.0252f
C22338 VGND.n1578 0 0.0298f
C22339 VGND.n1579 0 0.00828f
C22340 VGND.n1580 0 0.00981f
C22341 VGND.n1581 0 0.0394f
C22342 VGND.t162 0 0.0803f
C22343 VGND.n1582 0 0.062f
C22344 VGND.n1583 0 0.0413f
C22345 VGND.n1584 0 0.0597f
C22346 VGND.n1585 0 0.0651f
C22347 VGND.n1586 0 0.0314f
C22348 VGND.n1587 0 0.00981f
C22349 VGND.n1588 0 0.0166f
C22350 VGND.n1589 0 0.015f
C22351 VGND.t118 0 0.157f
C22352 VGND.n1590 0 0.192f
C22353 VGND.n1591 0 0.0875f
C22354 VGND.t202 0 0.0427f
C22355 VGND.n1592 0 0.106f
C22356 VGND.n1593 0 0.00846f
C22357 VGND.t38 0 0.0837f
C22358 VGND.t352 0 0.0445f
C22359 VGND.t325 0 0.0445f
C22360 VGND.n1594 0 0.243f
C22361 VGND.n1595 0 0.032f
C22362 VGND.n1596 0 0.0351f
C22363 VGND.t161 0 0.0837f
C22364 VGND.n1597 0 0.324f
C22365 VGND.n1598 0 0.0232f
C22366 VGND.n1599 0 0.0265f
C22367 VGND.n1600 0 0.0148f
C22368 VGND.n1601 0 0.0166f
C22369 VGND.n1602 0 0.0258f
C22370 VGND.n1603 0 0.0105f
C22371 VGND.n1604 0 0.0119f
C22372 VGND.n1605 0 0.0354f
C22373 VGND.t69 0 0.082f
C22374 VGND.n1606 0 0.128f
C22375 VGND.n1607 0 0.045f
C22376 VGND.n1608 0 0.0119f
C22377 VGND.n1609 0 0.015f
C22378 VGND.n1610 0 0.00981f
C22379 VGND.n1611 0 0.0166f
C22380 VGND.n1612 0 0.0291f
C22381 VGND.n1613 0 0.0336f
C22382 VGND.n1614 0 0.0456f
C22383 VGND.n1615 0 0.00891f
C22384 VGND.n1616 0 0.0112f
C22385 VGND.n1617 0 0.052f
C22386 VGND.n1618 0 0.0976f
C22387 VGND.n1619 0 0.015f
C22388 VGND.n1620 0 0.0597f
C22389 VGND.n1621 0 0.0166f
C22390 VGND.n1622 0 0.059f
C22391 VGND.n1623 0 0.0166f
C22392 VGND.n1624 0 0.0166f
C22393 VGND.n1625 0 0.0166f
C22394 VGND.n1626 0 0.00981f
C22395 VGND.n1627 0 0.009f
C22396 VGND.n1628 0 0.00819f
C22397 VGND.n1629 0 0.0221f
C22398 VGND.n1630 0 0.206f
C22399 VGND.t216 0 0.226f
C22400 VGND.n1631 0 0.342f
C22401 VGND.n1632 0 0.0439f
C22402 VGND.n1633 0 0.0153f
C22403 VGND.n1634 0 0.0944f
C22404 VGND.n1635 0 8.1e-19
C22405 VGND.n1636 0 0.00198f
C22406 VGND.n1637 0 1.46e-19
C22407 VGND.n1638 0 0.00185f
C22408 VGND.n1639 0 9.77e-19
C22409 VGND.n1640 0 0.0255f
C22410 VGND.n1641 0 0.138f
C22411 VGND.n1642 0 0.00126f
C22412 VGND.n1643 0 0.0232f
C22413 VGND.n1644 0 0.0257f
C22414 VGND.n1645 0 0.0107f
C22415 VGND.t175 0 0.0812f
C22416 VGND.n1646 0 0.139f
C22417 VGND.n1647 0 0.0349f
C22418 VGND.n1648 0 0.0273f
C22419 VGND.n1649 0 0.0275f
C22420 VGND.n1650 0 0.0108f
C22421 VGND.t200 0 0.0812f
C22422 VGND.n1651 0 0.139f
C22423 VGND.n1652 0 0.0349f
C22424 VGND.n1653 0 0.0292f
C22425 VGND.t117 0 0.0812f
C22426 VGND.t94 0 0.0813f
C22427 VGND.n1654 0 0.139f
C22428 VGND.n1655 0 0.0331f
C22429 VGND.n1656 0 0.0554f
C22430 VGND.t159 0 0.128f
C22431 VGND.n1657 0 0.154f
C22432 VGND.n1658 0 0.0514f
C22433 VGND.n1659 0 0.0337f
C22434 VGND.n1660 0 0.0265f
C22435 VGND.t282 0 0.0837f
C22436 VGND.t106 0 0.126f
C22437 VGND.n1661 0 0.178f
C22438 VGND.n1662 0 0.186f
C22439 VGND.t335 0 0.0445f
C22440 VGND.t316 0 0.0445f
C22441 VGND.n1663 0 0.243f
C22442 VGND.n1664 0 0.0173f
C22443 VGND.n1665 0 0.0247f
C22444 VGND.n1666 0 0.0329f
C22445 VGND.n1667 0 0.0453f
C22446 VGND.n1668 0 0.0378f
C22447 VGND.n1669 0 0.015f
C22448 VGND.n1670 0 0.00828f
C22449 VGND.n1671 0 0.0249f
C22450 VGND.n1672 0 0.0439f
C22451 VGND.n1673 0 0.00981f
C22452 VGND.n1674 0 0.0321f
C22453 VGND.n1675 0 0.0456f
C22454 VGND.n1676 0 0.0166f
C22455 VGND.t160 0 0.0946f
C22456 VGND.n1677 0 0.0183f
C22457 VGND.n1678 0 0.0961f
C22458 VGND.n1679 0 0.0322f
C22459 VGND.n1680 0 0.0271f
C22460 VGND.n1681 0 0.0166f
C22461 VGND.n1682 0 0.0345f
C22462 VGND.n1683 0 0.0252f
C22463 VGND.n1684 0 0.0166f
C22464 VGND.n1685 0 0.0316f
C22465 VGND.n1686 0 0.0166f
C22466 VGND.n1687 0 0.0324f
C22467 VGND.n1688 0 0.0166f
C22468 VGND.n1689 0 0.0331f
C22469 VGND.n1690 0 0.0166f
C22470 VGND.n1691 0 0.0513f
C22471 VGND.n1692 0 0.0166f
C22472 VGND.n1693 0 0.0445f
C22473 VGND.n1694 0 0.0166f
C22474 VGND.n1695 0 0.00513f
C22475 VGND.n1696 0 0.0149f
C22476 VGND.n1697 0 0.00837f
C22477 VGND.n1698 0 0.019f
C22478 VGND.n1699 0 0.0273f
C22479 VGND.n1700 0 0.0275f
C22480 VGND.n1701 0 0.0166f
C22481 VGND.n1702 0 0.0144f
C22482 VGND.n1703 0 0.00819f
C22483 VGND.n1704 0 0.00459f
C22484 VGND.n1705 0 0.049f
C22485 VGND.n1706 0 0.0301f
C22486 VGND.n1707 0 0.00828f
C22487 VGND.n1708 0 0.0172f
C22488 VGND.n1709 0 0.0349f
C22489 VGND.n1710 0 0.139f
C22490 VGND.n1711 0 0.0338f
C22491 VGND.n1712 0 0.00828f
C22492 VGND.n1713 0 0.00981f
C22493 VGND.n1714 0 0.00347f
C22494 VGND.n1715 0 0.0166f
C22495 VGND.n1716 0 0.015f
C22496 VGND.n1717 0 0.0361f
C22497 VGND.t67 0 0.0813f
C22498 VGND.n1718 0 0.139f
C22499 VGND.n1719 0 0.0402f
C22500 VGND.n1720 0 0.00828f
C22501 VGND.n1721 0 0.0165f
C22502 VGND.n1722 0 0.00891f
C22503 VGND.n1723 0 0.00963f
C22504 VGND.n1724 0 0.0166f
C22505 VGND.n1725 0 0.015f
C22506 VGND.n1726 0 0.00376f
C22507 VGND.t37 0 0.0813f
C22508 VGND.n1727 0 0.139f
C22509 VGND.n1728 0 0.0411f
C22510 VGND.n1729 0 0.00828f
C22511 VGND.n1730 0 0.0172f
C22512 VGND.n1731 0 0.0166f
C22513 VGND.n1732 0 0.0166f
C22514 VGND.n1733 0 0.015f
C22515 VGND.n1734 0 0.0253f
C22516 VGND.n1735 0 0.028f
C22517 VGND.n1736 0 0.00981f
C22518 VGND.t7 0 0.0792f
C22519 VGND.n1737 0 0.0547f
C22520 VGND.n1738 0 0.0314f
C22521 VGND.n1739 0 0.0166f
C22522 VGND.n1740 0 0.0491f
C22523 VGND.n1741 0 0.0136f
C22524 VGND.n1742 0 0.00369f
C22525 VGND.n1743 0 0.00234f
C22526 VGND.n1744 0 7.2e-19
C22527 VGND.n1745 0 0.00207f
C22528 VGND.n1746 0 0.00207f
C22529 VGND.n1747 0 0.00207f
C22530 VGND.n1748 0 0.00297f
C22531 VGND.n1749 0 0.00234f
C22532 VGND.n1750 0 0.00274f
C22533 VGND.n1751 0 0.00173f
C22534 VGND.n1752 0 0.00234f
C22535 VGND.n1753 0 0.0122f
C22536 VGND.t53 0 0.0813f
C22537 VGND.n1754 0 0.139f
C22538 VGND.n1755 0 0.0349f
C22539 VGND.t86 0 0.0792f
C22540 VGND.n1756 0 0.0284f
C22541 VGND.n1757 0 0.074f
C22542 VGND.n1758 0 0.0143f
C22543 VGND.n1759 0 0.0331f
C22544 VGND.n1760 0 0.0166f
C22545 VGND.n1761 0 0.0166f
C22546 VGND.n1762 0 0.00981f
C22547 VGND.n1763 0 0.028f
C22548 VGND.n1764 0 0.0386f
C22549 VGND.n1765 0 0.015f
C22550 VGND.n1766 0 0.00462f
C22551 VGND.n1767 0 0.0166f
C22552 VGND.n1768 0 0.00586f
C22553 VGND.n1769 0 0.0166f
C22554 VGND.n1770 0 0.00586f
C22555 VGND.n1771 0 0.0166f
C22556 VGND.n1772 0 0.00418f
C22557 VGND.n1773 0 0.0166f
C22558 VGND.n1774 0 0.0319f
C22559 VGND.n1775 0 0.0166f
C22560 VGND.n1776 0 0.0416f
C22561 VGND.n1777 0 0.0166f
C22562 VGND.n1778 0 0.00972f
C22563 VGND.n1779 0 0.0243f
C22564 VGND.t80 0 0.0812f
C22565 VGND.n1780 0 0.139f
C22566 VGND.n1781 0 0.0105f
C22567 VGND.n1782 0 0.00837f
C22568 VGND.n1783 0 0.0172f
C22569 VGND.n1784 0 0.00828f
C22570 VGND.n1785 0 0.00828f
C22571 VGND.n1786 0 0.0535f
C22572 VGND.n1787 0 0.013f
C22573 VGND.n1788 0 0.015f
C22574 VGND.n1789 0 0.0334f
C22575 VGND.n1790 0 0.0166f
C22576 VGND.n1791 0 0.00418f
C22577 VGND.n1792 0 0.0166f
C22578 VGND.n1793 0 0.00488f
C22579 VGND.n1794 0 0.0166f
C22580 VGND.n1795 0 0.032f
C22581 VGND.n1796 0 0.0166f
C22582 VGND.n1797 0 0.00437f
C22583 VGND.n1798 0 0.0166f
C22584 VGND.n1799 0 0.0379f
C22585 VGND.n1800 0 0.0166f
C22586 VGND.n1801 0 0.0428f
C22587 VGND.n1802 0 0.0166f
C22588 VGND.t54 0 0.0792f
C22589 VGND.n1803 0 0.0509f
C22590 VGND.n1804 0 0.038f
C22591 VGND.n1805 0 0.0153f
C22592 VGND.n1806 0 0.0127f
C22593 VGND.n1807 0 0.00828f
C22594 VGND.n1808 0 0.00153f
C22595 VGND.n1809 0 0.00135f
C22596 VGND.n1810 0 0.00297f
C22597 VGND.n1811 0 0.00315f
C22598 VGND.n1812 0 0.00207f
C22599 VGND.n1813 0 9.9e-19
C22600 VGND.n1814 0 0.00261f
C22601 VGND.n1815 0 0.00207f
C22602 VGND.n1816 0 0.00135f
C22603 VGND.n1817 0 7.2e-19
C22604 VGND.n1818 0 0.00126f
C22605 VGND.n1819 0 0.00414f
C22606 VGND.n1820 0 0.00423f
C22607 VGND.n1821 0 0.00126f
C22608 VGND.n1822 0 0.00912f
C22609 VGND.n1823 0 0.0101f
C22610 VGND.n1824 0 0.00126f
C22611 VGND.n1825 0 0.00824f
C22612 VGND.n1826 0 0.00413f
C22613 VGND.n1827 0 0.317f
C22614 VGND.n1828 0 0.317f
C22615 VGND.n1829 0 0.0039f
C22616 VGND.n1830 0 0.00269f
C22617 VGND.n1831 0 0.00207f
C22618 VGND.n1832 0 0.00287f
C22619 VGND.n1833 0 0.00173f
C22620 VGND.n1835 0 0.317f
C22621 VGND.n1836 0 0.317f
C22622 VGND.n1837 0 0.00207f
C22623 VGND.n1838 0 0.00287f
C22624 VGND.n1839 0 0.00269f
C22625 VGND.n1840 0 0.00173f
C22626 VGND.n1842 0 0.00274f
C22627 VGND.n1843 0 0.00173f
C22628 VGND.n1844 0 0.00369f
C22629 VGND.n1845 0 0.00234f
C22630 VGND.n1846 0 7.2e-19
C22631 VGND.n1847 0 0.00207f
C22632 VGND.n1848 0 0.00207f
C22633 VGND.n1849 0 0.00207f
C22634 VGND.n1850 0 0.00297f
C22635 VGND.n1851 0 0.00234f
C22636 VGND.n1852 0 0.00144f
C22637 VGND.n1853 0 0.00225f
C22638 VGND.n1854 0 0.00234f
C22639 VGND.n1855 0 0.00234f
C22640 VGND.n1856 0 0.00651f
C22641 VGND.n1857 0 0.00261f
C22642 VGND.n1858 0 0.00282f
C22643 VGND.n1859 0 0.00144f
C22644 VGND.n1860 0 0.00453f
C22645 VGND.n1861 0 0.00153f
C22646 VGND.n1862 0 0.0254f
C22647 VGND.n1863 0 0.00198f
C22648 VGND.n1864 0 0.00234f
C22649 VGND.n1865 0 0.0373f
C22650 VGND.n1866 0 0.00513f
C22651 VGND.n1867 0 0.0345f
C22652 VGND.n1868 0 0.0321f
C22653 VGND.n1869 0 0.0435f
C22654 VGND.t68 0 0.0946f
C22655 VGND.n1870 0 0.0183f
C22656 VGND.n1871 0 0.0961f
C22657 VGND.n1872 0 0.0272f
C22658 VGND.n1873 0 0.0271f
C22659 VGND.n1874 0 0.0514f
C22660 VGND.n1875 0 0.0244f
C22661 VGND.n1876 0 0.0254f
C22662 VGND.n1877 0 0.0334f
C22663 VGND.n1878 0 0.0468f
C22664 VGND.n1879 0 0.0379f
C22665 VGND.t20 0 0.128f
C22666 VGND.n1880 0 0.154f
C22667 VGND.n1881 0 0.0272f
C22668 VGND.n1882 0 0.00408f
C22669 VGND.n1883 0 0.0313f
C22670 VGND.n1884 0 0.0261f
C22671 VGND.n1885 0 0.0257f
C22672 VGND.t390 0 0.0792f
C22673 VGND.n1886 0 0.0547f
C22674 VGND.t245 0 0.0445f
C22675 VGND.t224 0 0.0445f
C22676 VGND.n1887 0 0.0279f
C22677 VGND.n1888 0 0.244f
C22678 VGND.n1889 0 0.0163f
C22679 VGND.n1890 0 0.00981f
C22680 VGND.n1891 0 0.015f
C22681 VGND.n1892 0 0.0243f
C22682 VGND.n1893 0 0.0337f
C22683 VGND.n1894 0 0.00981f
C22684 VGND.n1895 0 0.0541f
C22685 VGND.n1896 0 0.0166f
C22686 VGND.n1897 0 0.0166f
C22687 VGND.n1898 0 0.0166f
C22688 VGND.n1899 0 0.015f
C22689 VGND.n1900 0 0.019f
C22690 VGND.n1901 0 0.037f
C22691 VGND.n1902 0 0.0275f
C22692 VGND.n1903 0 0.0166f
C22693 VGND.n1904 0 0.0144f
C22694 VGND.n1905 0 0.00891f
C22695 VGND.n1906 0 0.00549f
C22696 VGND.n1907 0 0.00625f
C22697 VGND.n1908 0 0.00981f
C22698 VGND.n1909 0 0.0413f
C22699 VGND.n1910 0 0.0166f
C22700 VGND.n1911 0 0.0125f
C22701 VGND.n1912 0 0.0166f
C22702 VGND.n1913 0 0.0166f
C22703 VGND.n1914 0 0.00335f
C22704 VGND.n1915 0 0.0166f
C22705 VGND.n1916 0 0.0166f
C22706 VGND.n1917 0 0.015f
C22707 VGND.n1918 0 0.00437f
C22708 VGND.n1919 0 0.0291f
C22709 VGND.n1920 0 0.00981f
C22710 VGND.t176 0 0.0792f
C22711 VGND.n1921 0 0.0547f
C22712 VGND.n1922 0 0.0243f
C22713 VGND.n1923 0 0.0166f
C22714 VGND.n1924 0 0.0166f
C22715 VGND.n1925 0 0.0428f
C22716 VGND.n1926 0 0.0504f
C22717 VGND.n1927 0 0.0143f
C22718 VGND.n1928 0 0.009f
C22719 VGND.n1929 0 0.0367f
C22720 VGND.n1930 0 0.00981f
C22721 VGND.t107 0 0.121f
C22722 VGND.n1931 0 0.112f
C22723 VGND.n1932 0 0.0166f
C22724 VGND.n1933 0 0.0504f
C22725 VGND.n1934 0 0.0166f
C22726 VGND.n1935 0 0.0395f
C22727 VGND.n1936 0 0.0166f
C22728 VGND.n1937 0 0.0166f
C22729 VGND.n1938 0 0.0331f
C22730 VGND.n1939 0 0.0369f
C22731 VGND.n1940 0 0.0144f
C22732 VGND.n1941 0 0.009f
C22733 VGND.n1942 0 0.00819f
C22734 VGND.n1943 0 0.0234f
C22735 VGND.n1944 0 0.0443f
C22736 VGND.n1945 0 0.00981f
C22737 VGND.n1946 0 0.0166f
C22738 VGND.n1947 0 0.0166f
C22739 VGND.n1948 0 0.015f
C22740 VGND.n1949 0 0.0298f
C22741 VGND.n1950 0 0.0488f
C22742 VGND.n1951 0 0.00981f
C22743 VGND.n1952 0 0.0166f
C22744 VGND.n1953 0 0.0166f
C22745 VGND.t119 0 0.0792f
C22746 VGND.n1954 0 0.068f
C22747 VGND.n1955 0 0.0442f
C22748 VGND.n1956 0 0.0604f
C22749 VGND.n1957 0 0.0686f
C22750 VGND.n1958 0 0.0142f
C22751 VGND.n1959 0 0.00972f
C22752 VGND.n1960 0 0.015f
C22753 VGND.n1961 0 0.00828f
C22754 VGND.n1962 0 0.0448f
C22755 VGND.n1963 0 0.0362f
C22756 VGND.n1964 0 0.00981f
C22757 VGND.t191 0 0.0792f
C22758 VGND.n1965 0 0.0547f
C22759 VGND.n1966 0 0.0344f
C22760 VGND.n1967 0 0.0166f
C22761 VGND.n1968 0 0.0166f
C22762 VGND.n1969 0 0.015f
C22763 VGND.n1970 0 0.0375f
C22764 VGND.n1971 0 0.0287f
C22765 VGND.n1972 0 0.00981f
C22766 VGND.t389 0 0.0792f
C22767 VGND.n1973 0 0.0566f
C22768 VGND.n1974 0 0.04f
C22769 VGND.n1975 0 0.0166f
C22770 VGND.n1976 0 0.0312f
C22771 VGND.n1977 0 0.0136f
C22772 VGND.n1978 0 0.0063f
C22773 VGND.n1979 0 0.00824f
C22774 VGND.n1980 0 0.00413f
C22775 VGND.n1981 0 0.018f
C22776 VGND.n1982 0 0.0039f
C22777 VGND.n1983 0 0.00269f
C22778 VGND.n1984 0 0.00207f
C22779 VGND.n1985 0 0.00287f
C22780 VGND.n1986 0 0.00173f
C22781 VGND.n1988 0 0.317f
C22782 VGND.n1989 0 0.317f
C22783 VGND.n1990 0 0.00207f
C22784 VGND.n1991 0 0.00287f
C22785 VGND.n1992 0 0.00269f
C22786 VGND.n1993 0 0.00173f
C22787 VGND.n1995 0 0.018f
C22788 VGND.n1996 0 0.00274f
C22789 VGND.n1997 0 0.00173f
C22790 VGND.n1998 0 0.00413f
C22791 VGND.n1999 0 0.00824f
C22792 VGND.n2000 0 0.0063f
C22793 VGND.n2001 0 0.00234f
C22794 VGND.n2002 0 0.0254f
C22795 VGND.n2003 0 0.00198f
C22796 VGND.n2004 0 0.00453f
C22797 VGND.n2005 0 0.00153f
C22798 VGND.n2006 0 0.00282f
C22799 VGND.n2007 0 0.00144f
C22800 VGND.n2008 0 0.00651f
C22801 VGND.n2009 0 0.00261f
C22802 VGND.n2010 0 0.00234f
C22803 VGND.n2011 0 0.00234f
C22804 VGND.n2012 0 0.00225f
C22805 VGND.n2013 0 0.00144f
C22806 VGND.n2014 0 0.00148f
C22807 VGND.n2015 0 8.57e-19
C22808 VGND.n2016 0 0.0252f
C22809 VGND.n2017 0 0.229f
C22810 VGND.n2018 0 0.229f
C22811 VGND.n2019 0 0.026f
C22812 VGND.n2020 0 0.009f
C22813 VGND.n2021 0 0.0388f
C22814 VGND.n2022 0 0.00981f
C22815 VGND.t140 0 0.0792f
C22816 VGND.n2023 0 0.0689f
C22817 VGND.n2024 0 0.0243f
C22818 VGND.n2025 0 0.0166f
C22819 VGND.n2026 0 0.0166f
C22820 VGND.n2027 0 0.0331f
C22821 VGND.n2028 0 0.0369f
C22822 VGND.n2029 0 0.0151f
C22823 VGND.n2030 0 0.00972f
C22824 VGND.n2031 0 0.015f
C22825 VGND.n2032 0 0.019f
C22826 VGND.n2033 0 0.0273f
C22827 VGND.n2034 0 0.0275f
C22828 VGND.n2035 0 0.0166f
C22829 VGND.n2036 0 0.0144f
C22830 VGND.n2037 0 0.019f
C22831 VGND.n2038 0 0.026f
C22832 VGND.n2039 0 0.00828f
C22833 VGND.n2040 0 0.0766f
C22834 VGND.n2041 0 0.0463f
C22835 VGND.t210 0 0.158f
C22836 VGND.n2042 0 0.185f
C22837 VGND.n2043 0 0.0213f
C22838 VGND.n2044 0 0.00765f
C22839 VGND.n2045 0 0.00891f
C22840 VGND.n2046 0 0.0137f
C22841 VGND.n2047 0 0.0281f
C22842 VGND.n2048 0 0.0221f
C22843 VGND.n2049 0 0.0523f
C22844 VGND.n2050 0 0.0166f
C22845 VGND.n2051 0 0.0166f
C22846 VGND.n2052 0 0.0387f
C22847 VGND.n2053 0 0.0379f
C22848 VGND.n2054 0 0.0142f
C22849 VGND.n2055 0 0.00891f
C22850 VGND.n2056 0 0.00783f
C22851 VGND.n2057 0 0.00207f
C22852 VGND.n2058 0 0.00315f
C22853 VGND.n2059 0 0.00162f
C22854 VGND.n2060 0 0.00162f
C22855 VGND.n2061 0 0.00189f
C22856 VGND.n2062 0 9.9e-19
C22857 VGND.n2063 0 0.00162f
C22858 VGND.n2064 0 0.00171f
C22859 VGND.n2065 0 0.00494f
C22860 VGND.n2066 0 9.9e-19
C22861 VGND.n2067 0 0.00189f
C22862 VGND.n2068 0 0.00162f
C22863 VGND.n2069 0 0.00342f
C22864 VGND.n2070 0 0.00387f
C22865 VGND.n2071 0 7.2e-19
C22866 VGND.n2072 0 0.00162f
C22867 VGND.n2073 0 0.00207f
C22868 VGND.n2074 0 0.00207f
C22869 VGND.n2075 0 0.00162f
C22870 VGND.n2076 0 0.00234f
C22871 VGND.n2077 0 0.00234f
C22872 VGND.n2078 0 0.00234f
C22873 VGND.n2079 0 0.00297f
C22874 VGND.n2080 0 0.00842f
C22875 VGND.n2081 0 0.00144f
C22876 VGND.n2082 0 0.00135f
C22877 VGND.n2083 0 2.7e-19
C22878 VGND.n2084 0 0.003f
C22879 VGND.n2085 0 0.0179f
C22880 VGND.n2086 0 0.00126f
C22881 VGND.n2087 0 0.00207f
C22882 VGND.n2088 0 0.00126f
C22883 VGND.n2089 0 0.00126f
C22884 VGND.n2090 0 0.00701f
C22885 VGND.n2091 0 0.0041f
C22886 VGND.n2092 0 0.018f
C22887 VGND.n2093 0 0.00287f
C22888 VGND.n2094 0 0.00207f
C22889 VGND.n2095 0 0.00274f
C22890 VGND.n2096 0 0.00403f
C22891 VGND.n2097 0 0.00493f
C22892 VGND.n2098 0 0.00126f
C22893 VGND.n2099 0 0.00173f
C22894 VGND.n2101 0 0.317f
C22895 VGND.n2102 0 0.317f
C22896 VGND.n2103 0 0.00207f
C22897 VGND.n2104 0 0.00287f
C22898 VGND.n2105 0 0.00173f
C22899 VGND.n2106 0 0.00269f
C22900 VGND.n2107 0 0.0039f
C22901 VGND.n2108 0 0.00269f
C22902 VGND.n2109 0 0.00173f
C22903 VGND.n2111 0 0.00274f
C22904 VGND.n2112 0 0.00173f
C22905 VGND.n2113 0 0.00207f
C22906 VGND.n2114 0 0.00603f
C22907 VGND.n2115 0 0.00234f
C22908 VGND.n2116 0 0.00135f
C22909 VGND.n2117 0 0.00189f
C22910 VGND.n2118 0 0.00369f
C22911 VGND.n2119 0 0.00252f
C22912 VGND.n2120 0 7.2e-19
C22913 VGND.n2121 0 7.2e-19
C22914 VGND.n2122 0 8.1e-19
C22915 VGND.n2123 0 0.213f
C22916 VGND.n2124 0 0.0245f
C22917 VGND.n2125 0 0.0646f
C22918 VGND.n2126 0 0.00828f
C22919 VGND.n2127 0 0.00828f
C22920 VGND.t306 0 0.082f
C22921 VGND.n2128 0 0.0934f
C22922 VGND.n2129 0 0.015f
C22923 VGND.n2130 0 0.065f
C22924 VGND.t373 0 0.128f
C22925 VGND.n2131 0 0.198f
C22926 VGND.n2132 0 0.0628f
C22927 VGND.t302 0 0.0445f
C22928 VGND.t277 0 0.0445f
C22929 VGND.n2133 0 0.243f
C22930 VGND.n2134 0 0.0159f
C22931 VGND.t264 0 0.0812f
C22932 VGND.n2135 0 0.139f
C22933 VGND.n2136 0 0.0107f
C22934 VGND.n2137 0 0.0205f
C22935 VGND.n2138 0 0.0165f
C22936 VGND.n2139 0 0.0173f
C22937 VGND.n2140 0 0.0317f
C22938 VGND.n2141 0 0.0375f
C22939 VGND.n2142 0 0.0543f
C22940 VGND.n2143 0 0.00981f
C22941 VGND.n2144 0 0.0119f
C22942 VGND.n2145 0 0.0217f
C22943 VGND.t22 0 0.0816f
C22944 VGND.n2146 0 0.139f
C22945 VGND.n2147 0 0.0496f
C22946 VGND.n2148 0 0.0534f
C22947 VGND.n2149 0 0.015f
C22948 VGND.n2150 0 0.00674f
C22949 VGND.n2151 0 0.0104f
C22950 VGND.n2152 0 0.00765f
C22951 VGND.n2153 0 0.00891f
C22952 VGND.n2154 0 0.0321f
C22953 VGND.n2155 0 0.0651f
C22954 VGND.n2156 0 0.0144f
C22955 VGND.n2157 0 0.0597f
C22956 VGND.n2158 0 0.0166f
C22957 VGND.n2159 0 0.059f
C22958 VGND.n2160 0 0.0166f
C22959 VGND.n2161 0 0.0166f
C22960 VGND.n2162 0 0.0166f
C22961 VGND.t289 0 0.155f
C22962 VGND.n2163 0 0.0449f
C22963 VGND.n2164 0 0.163f
C22964 VGND.n2165 0 0.0295f
C22965 VGND.n2166 0 0.0603f
C22966 VGND.n2167 0 0.0327f
C22967 VGND.n2168 0 0.00981f
C22968 VGND.n2169 0 0.0243f
C22969 VGND.t370 0 0.0792f
C22970 VGND.n2170 0 0.0547f
C22971 VGND.n2171 0 0.0348f
C22972 VGND.t48 0 0.0792f
C22973 VGND.n2172 0 0.0681f
C22974 VGND.t87 0 0.0837f
C22975 VGND.n2173 0 0.185f
C22976 VGND.n2174 0 0.0273f
C22977 VGND.t353 0 0.158f
C22978 VGND.n2175 0 0.258f
C22979 VGND.n2176 0 0.0122f
C22980 VGND.n2177 0 0.0287f
C22981 VGND.n2178 0 0.0513f
C22982 VGND.n2179 0 0.0825f
C22983 VGND.n2180 0 0.014f
C22984 VGND.n2181 0 0.0411f
C22985 VGND.n2182 0 0.0329f
C22986 VGND.n2183 0 0.0279f
C22987 VGND.n2184 0 0.015f
C22988 VGND.n2185 0 0.00828f
C22989 VGND.n2186 0 0.00828f
C22990 VGND.n2187 0 0.0192f
C22991 VGND.t265 0 0.0799f
C22992 VGND.n2188 0 0.0723f
C22993 VGND.n2189 0 0.0245f
C22994 VGND.n2190 0 0.00981f
C22995 VGND.n2191 0 0.0166f
C22996 VGND.n2192 0 0.015f
C22997 VGND.n2193 0 0.0379f
C22998 VGND.n2194 0 0.00444f
C22999 VGND.n2195 0 0.00981f
C23000 VGND.n2196 0 0.0166f
C23001 VGND.n2197 0 0.0221f
C23002 VGND.n2198 0 0.015f
C23003 VGND.n2199 0 0.00828f
C23004 VGND.n2200 0 0.0247f
C23005 VGND.n2201 0 0.0329f
C23006 VGND.n2202 0 0.0338f
C23007 VGND.n2203 0 0.0151f
C23008 VGND.n2204 0 0.00756f
C23009 VGND.n2205 0 0.00828f
C23010 VGND.n2206 0 0.0287f
C23011 VGND.n2207 0 0.0547f
C23012 VGND.n2208 0 0.0506f
C23013 VGND.n2209 0 0.00981f
C23014 VGND.n2210 0 0.0166f
C23015 VGND.n2211 0 0.015f
C23016 VGND.n2212 0 0.062f
C23017 VGND.n2213 0 0.0578f
C23018 VGND.n2214 0 0.00981f
C23019 VGND.n2215 0 0.0149f
C23020 VGND.n2216 0 0.00837f
C23021 VGND.n2217 0 0.0834f
C23022 VGND.t9 0 0.148f
C23023 VGND.n2218 0 0.0882f
C23024 VGND.n2219 0 0.0584f
C23025 VGND.n2220 0 0.0214f
C23026 VGND.n2221 0 0.00756f
C23027 VGND.n2222 0 0.009f
C23028 VGND.n2223 0 0.0316f
C23029 VGND.n2224 0 0.094f
C23030 VGND.n2225 0 0.094f
C23031 VGND.n2226 0 0.0316f
C23032 VGND.n2227 0 9.77e-19
C23033 VGND.n2228 0 0.00185f
C23034 VGND.n2229 0 1.46e-19
C23035 VGND.n2230 0 0.00198f
C23036 VGND.n2231 0 0.00162f
C23037 VGND.n2232 0 0.00207f
C23038 VGND.n2233 0 0.00315f
C23039 VGND.n2234 0 0.00162f
C23040 VGND.n2235 0 0.00162f
C23041 VGND.n2236 0 0.00189f
C23042 VGND.n2237 0 9.9e-19
C23043 VGND.n2238 0 0.00162f
C23044 VGND.n2239 0 0.00153f
C23045 VGND.n2240 0 0.0157f
C23046 VGND.n2241 0 9.9e-19
C23047 VGND.n2242 0 0.00189f
C23048 VGND.n2243 0 0.00162f
C23049 VGND.n2244 0 0.00342f
C23050 VGND.n2245 0 0.00387f
C23051 VGND.n2246 0 7.2e-19
C23052 VGND.n2247 0 0.00162f
C23053 VGND.n2248 0 0.00207f
C23054 VGND.n2249 0 0.00207f
C23055 VGND.n2250 0 0.00162f
C23056 VGND.n2251 0 0.00234f
C23057 VGND.n2252 0 0.00234f
C23058 VGND.n2253 0 0.00234f
C23059 VGND.n2254 0 0.00297f
C23060 VGND.n2255 0 0.00144f
C23061 VGND.n2256 0 0.00151f
C23062 VGND.t319 0 0.0818f
C23063 VGND.n2257 0 0.139f
C23064 VGND.t71 0 0.124f
C23065 VGND.n2258 0 0.125f
C23066 VGND.n2259 0 0.0318f
C23067 VGND.n2260 0 1.12e-19
C23068 VGND.n2261 0 0.00126f
C23069 VGND.n2262 0 0.00207f
C23070 VGND.n2263 0 0.00126f
C23071 VGND.n2264 0 0.00126f
C23072 VGND.n2265 0 0.00701f
C23073 VGND.n2266 0 0.0041f
C23074 VGND.n2267 0 0.018f
C23075 VGND.n2269 0 0.00403f
C23076 VGND.n2270 0 0.00173f
C23077 VGND.n2271 0 0.00126f
C23078 VGND.n2272 0 0.00493f
C23079 VGND.n2273 0 0.00675f
C23080 VGND.n2274 0 0.0853f
C23081 VGND.n2275 0 0.0148f
C23082 VGND.t23 0 0.0792f
C23083 VGND.n2276 0 0.0547f
C23084 VGND.n2277 0 0.0243f
C23085 VGND.n2278 0 0.0166f
C23086 VGND.n2279 0 0.00972f
C23087 VGND.n2280 0 0.00828f
C23088 VGND.n2281 0 0.0639f
C23089 VGND.t367 0 0.0799f
C23090 VGND.n2282 0 0.0723f
C23091 VGND.n2283 0 0.0486f
C23092 VGND.n2284 0 0.0348f
C23093 VGND.n2285 0 0.015f
C23094 VGND.n2286 0 0.0166f
C23095 VGND.n2287 0 0.00981f
C23096 VGND.n2288 0 0.00828f
C23097 VGND.n2289 0 0.0766f
C23098 VGND.n2290 0 0.0334f
C23099 VGND.n2291 0 0.0346f
C23100 VGND.n2292 0 0.015f
C23101 VGND.n2293 0 0.0166f
C23102 VGND.n2294 0 0.0555f
C23103 VGND.n2295 0 0.0275f
C23104 VGND.n2296 0 0.019f
C23105 VGND.n2297 0 0.00828f
C23106 VGND.n2298 0 0.0795f
C23107 VGND.n2299 0 0.0369f
C23108 VGND.n2300 0 0.0571f
C23109 VGND.n2301 0 0.015f
C23110 VGND.n2302 0 0.0166f
C23111 VGND.t74 0 0.0792f
C23112 VGND.n2303 0 0.0547f
C23113 VGND.n2304 0 0.0411f
C23114 VGND.n2305 0 0.0166f
C23115 VGND.n2306 0 0.00981f
C23116 VGND.n2307 0 0.00819f
C23117 VGND.n2308 0 0.0538f
C23118 VGND.n2309 0 0.0548f
C23119 VGND.n2310 0 0.0368f
C23120 VGND.n2311 0 0.0151f
C23121 VGND.n2312 0 0.00972f
C23122 VGND.n2313 0 0.012f
C23123 VGND.n2314 0 0.0217f
C23124 VGND.t112 0 0.0816f
C23125 VGND.n2315 0 0.139f
C23126 VGND.n2316 0 0.00756f
C23127 VGND.n2317 0 0.0396f
C23128 VGND.n2318 0 0.0351f
C23129 VGND.n2319 0 0.0655f
C23130 VGND.n2320 0 0.0144f
C23131 VGND.n2321 0 0.0166f
C23132 VGND.t195 0 0.0792f
C23133 VGND.n2322 0 0.0547f
C23134 VGND.n2323 0 0.0243f
C23135 VGND.n2324 0 0.0166f
C23136 VGND.n2325 0 0.0291f
C23137 VGND.n2326 0 0.00981f
C23138 VGND.n2327 0 0.00412f
C23139 VGND.n2328 0 0.015f
C23140 VGND.n2329 0 0.0389f
C23141 VGND.n2330 0 0.0166f
C23142 VGND.n2331 0 0.0166f
C23143 VGND.n2332 0 0.00972f
C23144 VGND.n2333 0 0.009f
C23145 VGND.n2334 0 0.0104f
C23146 VGND.n2335 0 0.0578f
C23147 VGND.n2336 0 0.0144f
C23148 VGND.n2337 0 0.0489f
C23149 VGND.n2338 0 0.0166f
C23150 VGND.n2339 0 0.0366f
C23151 VGND.n2340 0 0.0275f
C23152 VGND.n2341 0 0.019f
C23153 VGND.n2342 0 0.00819f
C23154 VGND.n2343 0 0.00593f
C23155 VGND.n2344 0 0.0362f
C23156 VGND.n2345 0 0.0151f
C23157 VGND.n2346 0 0.0331f
C23158 VGND.n2347 0 0.0166f
C23159 VGND.n2348 0 0.0166f
C23160 VGND.n2349 0 0.00981f
C23161 VGND.n2350 0 0.00828f
C23162 VGND.n2351 0 0.0112f
C23163 VGND.n2352 0 0.0531f
C23164 VGND.n2353 0 0.015f
C23165 VGND.n2354 0 0.00972f
C23166 VGND.n2355 0 0.00549f
C23167 VGND.n2356 0 0.0578f
C23168 VGND.n2357 0 0.0151f
C23169 VGND.n2358 0 0.0387f
C23170 VGND.n2359 0 0.0166f
C23171 VGND.t177 0 0.0792f
C23172 VGND.n2360 0 0.0509f
C23173 VGND.n2361 0 0.0243f
C23174 VGND.n2362 0 0.0153f
C23175 VGND.n2363 0 0.0127f
C23176 VGND.n2364 0 0.00828f
C23177 VGND.n2365 0 0.00153f
C23178 VGND.n2366 0 0.00423f
C23179 VGND.n2367 0 0.00126f
C23180 VGND.n2368 0 0.00912f
C23181 VGND.n2369 0 0.0101f
C23182 VGND.n2370 0 0.00126f
C23183 VGND.n2371 0 0.00824f
C23184 VGND.n2372 0 0.00234f
C23185 VGND.n2373 0 0.00297f
C23186 VGND.n2374 0 0.00315f
C23187 VGND.n2375 0 0.00207f
C23188 VGND.n2376 0 9.9e-19
C23189 VGND.n2377 0 0.00261f
C23190 VGND.n2378 0 0.00207f
C23191 VGND.n2379 0 0.00135f
C23192 VGND.n2380 0 7.2e-19
C23193 VGND.n2381 0 0.00126f
C23194 VGND.n2382 0 0.00135f
C23195 VGND.n2383 0 0.00126f
C23196 VGND.n2384 0 0.00153f
C23197 VGND.n2385 0 0.0026f
C23198 VGND.n2386 0 0.00198f
C23199 VGND.n2387 0 5.42e-19
C23200 VGND.n2388 0 0.00153f
C23201 VGND.n2389 0 5.1e-19
C23202 VGND.n2390 0 0.00144f
C23203 VGND.n2391 0 0.00169f
C23204 VGND.n2392 0 0.00261f
C23205 VGND.n2393 0 0.00234f
C23206 VGND.n2394 0 0.00369f
C23207 VGND.n2395 0 0.00297f
C23208 VGND.n2396 0 0.00207f
C23209 VGND.n2397 0 0.00207f
C23210 VGND.n2398 0 0.00207f
C23211 VGND.n2399 0 7.2e-19
C23212 VGND.n2400 0 0.00234f
C23213 VGND.n2401 0 0.00234f
C23214 VGND.n2402 0 0.00225f
C23215 VGND.n2403 0 0.00144f
C23216 VGND.n2404 0 0.00148f
C23217 VGND.n2405 0 8.57e-19
C23218 VGND.n2406 0 0.0254f
C23219 VGND.n2407 0 0.0945f
C23220 VGND.n2408 0 0.229f
C23221 VGND.n2409 0 0.0331f
C23222 VGND.n2410 0 0.0379f
C23223 VGND.n2411 0 0.0278f
C23224 VGND.n2412 0 0.053f
C23225 VGND.n2413 0 0.0435f
C23226 VGND.t312 0 0.119f
C23227 VGND.n2414 0 0.053f
C23228 VGND.n2415 0 0.0433f
C23229 VGND.n2416 0 0.0834f
C23230 VGND.n2417 0 0.00981f
C23231 VGND.t149 0 0.0792f
C23232 VGND.t376 0 0.0792f
C23233 VGND.n2418 0 0.0567f
C23234 VGND.n2419 0 0.0245f
C23235 VGND.n2420 0 0.053f
C23236 VGND.t142 0 0.0792f
C23237 VGND.n2421 0 0.0547f
C23238 VGND.n2422 0 0.0534f
C23239 VGND.n2423 0 0.0331f
C23240 VGND.t290 0 0.0445f
C23241 VGND.n2424 0 0.0166f
C23242 VGND.t261 0 0.0445f
C23243 VGND.n2425 0 0.244f
C23244 VGND.n2426 0 0.0279f
C23245 VGND.n2427 0 0.00981f
C23246 VGND.n2428 0 0.0166f
C23247 VGND.n2429 0 0.0149f
C23248 VGND.n2430 0 0.00837f
C23249 VGND.n2431 0 0.0647f
C23250 VGND.n2432 0 0.0451f
C23251 VGND.n2433 0 0.00981f
C23252 VGND.n2434 0 0.0166f
C23253 VGND.n2435 0 0.015f
C23254 VGND.n2436 0 0.0375f
C23255 VGND.n2437 0 0.0578f
C23256 VGND.n2438 0 0.0547f
C23257 VGND.n2439 0 0.0243f
C23258 VGND.n2440 0 0.0149f
C23259 VGND.n2441 0 0.00837f
C23260 VGND.n2442 0 0.00828f
C23261 VGND.n2443 0 0.0158f
C23262 VGND.n2444 0 0.0374f
C23263 VGND.n2445 0 0.0162f
C23264 VGND.n2446 0 0.00981f
C23265 VGND.n2447 0 0.0447f
C23266 VGND.n2448 0 0.0166f
C23267 VGND.n2449 0 0.0324f
C23268 VGND.n2450 0 0.0166f
C23269 VGND.n2451 0 0.0166f
C23270 VGND.n2452 0 0.0144f
C23271 VGND.n2453 0 0.00891f
C23272 VGND.n2454 0 0.00549f
C23273 VGND.n2455 0 0.005f
C23274 VGND.n2456 0 0.0166f
C23275 VGND.n2457 0 0.00616f
C23276 VGND.n2458 0 0.0166f
C23277 VGND.n2459 0 0.015f
C23278 VGND.n2460 0 0.028f
C23279 VGND.n2461 0 0.047f
C23280 VGND.n2462 0 0.00981f
C23281 VGND.t311 0 0.0792f
C23282 VGND.n2463 0 0.0547f
C23283 VGND.n2464 0 0.0243f
C23284 VGND.n2465 0 0.0166f
C23285 VGND.n2466 0 0.0166f
C23286 VGND.n2467 0 0.0143f
C23287 VGND.n2468 0 0.009f
C23288 VGND.n2469 0 0.0392f
C23289 VGND.n2470 0 0.0386f
C23290 VGND.n2471 0 0.00981f
C23291 VGND.t229 0 0.0792f
C23292 VGND.n2472 0 0.0547f
C23293 VGND.n2473 0 0.0243f
C23294 VGND.n2474 0 0.0166f
C23295 VGND.n2475 0 0.0166f
C23296 VGND.n2476 0 0.015f
C23297 VGND.n2477 0 0.0554f
C23298 VGND.n2478 0 0.00509f
C23299 VGND.n2479 0 0.00981f
C23300 VGND.n2480 0 0.0166f
C23301 VGND.n2481 0 0.015f
C23302 VGND.n2482 0 0.0349f
C23303 VGND.n2483 0 0.0431f
C23304 VGND.n2484 0 0.0512f
C23305 VGND.n2485 0 0.00981f
C23306 VGND.t332 0 0.121f
C23307 VGND.n2486 0 0.138f
C23308 VGND.n2487 0 0.0166f
C23309 VGND.n2488 0 0.0166f
C23310 VGND.n2489 0 0.0166f
C23311 VGND.n2490 0 0.0142f
C23312 VGND.n2491 0 0.00846f
C23313 VGND.n2492 0 0.0155f
C23314 VGND.n2493 0 0.00414f
C23315 VGND.n2494 0 0.009f
C23316 VGND.n2495 0 0.00972f
C23317 VGND.n2496 0 0.0166f
C23318 VGND.n2497 0 0.0166f
C23319 VGND.n2498 0 0.00325f
C23320 VGND.n2499 0 0.0166f
C23321 VGND.n2500 0 0.015f
C23322 VGND.n2501 0 0.019f
C23323 VGND.n2502 0 0.0273f
C23324 VGND.n2503 0 0.0275f
C23325 VGND.n2504 0 0.0468f
C23326 VGND.n2505 0 0.0166f
C23327 VGND.n2506 0 0.0473f
C23328 VGND.n2507 0 0.0136f
C23329 VGND.n2508 0 0.00612f
C23330 VGND.n2509 0 0.00824f
C23331 VGND.n2510 0 0.00413f
C23332 VGND.n2511 0 0.018f
C23333 VGND.n2512 0 0.0039f
C23334 VGND.n2513 0 0.00269f
C23335 VGND.n2514 0 0.00207f
C23336 VGND.n2515 0 0.00287f
C23337 VGND.n2516 0 0.00173f
C23338 VGND.n2518 0 0.206f
C23339 VGND.n2519 0 0.12f
C23340 VGND.n2520 0 0.308f
C23341 VGND.n2521 0 4.5f
C23342 VGND.n2522 0 3.67f
C23343 VGND.n2523 0 0.12f
C23344 VGND.n2524 0 0.00207f
C23345 VGND.n2525 0 0.00287f
C23346 VGND.n2526 0 0.00173f
C23347 VGND.n2527 0 0.00269f
C23348 VGND.n2528 0 0.0039f
C23349 VGND.n2529 0 0.00269f
C23350 VGND.n2530 0 0.00173f
C23351 VGND.n2532 0 0.317f
C23352 VGND.n2533 0 0.317f
C23353 VGND.n2534 0 0.00287f
C23354 VGND.n2535 0 0.00207f
C23355 VGND.n2536 0 0.00274f
C23356 VGND.n2537 0 0.00403f
C23357 VGND.n2538 0 0.00493f
C23358 VGND.n2539 0 0.00126f
C23359 VGND.n2540 0 0.00173f
C23360 VGND.n2542 0 0.018f
C23361 VGND.n2543 0 0.00274f
C23362 VGND.n2544 0 0.00173f
C23363 VGND.n2545 0 0.0041f
C23364 VGND.n2546 0 0.00701f
C23365 VGND.n2547 0 0.00252f
C23366 VGND.n2548 0 0.00369f
C23367 VGND.n2549 0 0.00189f
C23368 VGND.n2550 0 0.00135f
C23369 VGND.n2551 0 0.00207f
C23370 VGND.n2552 0 0.00126f
C23371 VGND.n2553 0 0.00126f
C23372 VGND.n2554 0 0.00207f
C23373 VGND.n2555 0 0.0392f
C23374 VGND.n2556 0 0.003f
C23375 VGND.n2557 0 5.29e-19
C23376 VGND.n2558 0 0.00126f
C23377 VGND.n2559 0 2.7e-19
C23378 VGND.n2560 0 0.00135f
C23379 VGND.n2561 0 0.00407f
C23380 VGND.n2562 0 0.00511f
C23381 VGND.n2563 0 0.00144f
C23382 VGND.n2564 0 0.00297f
C23383 VGND.n2565 0 0.00234f
C23384 VGND.n2566 0 0.00234f
C23385 VGND.n2567 0 0.00234f
C23386 VGND.n2568 0 0.00234f
C23387 VGND.n2569 0 0.00162f
C23388 VGND.n2570 0 0.00207f
C23389 VGND.n2571 0 0.00207f
C23390 VGND.n2572 0 0.00162f
C23391 VGND.n2573 0 0.00342f
C23392 VGND.n2574 0 0.00162f
C23393 VGND.n2575 0 0.00189f
C23394 VGND.n2576 0 0.054f
C23395 VGND.n2577 0 9.92e-19
C23396 VGND.n2578 0 0.0205f
C23397 VGND.n2579 0 0.0173f
C23398 VGND.n2580 0 0.0631f
C23399 VGND.n2581 0 0.0271f
C23400 VGND.t171 0 0.0946f
C23401 VGND.n2582 0 0.0183f
C23402 VGND.n2583 0 0.0961f
C23403 VGND.n2584 0 0.041f
C23404 VGND.n2585 0 0.0402f
C23405 VGND.n2586 0 0.0321f
C23406 VGND.n2587 0 0.00565f
C23407 VGND.n2588 0 0.0319f
C23408 VGND.n2589 0 0.011f
C23409 VGND.t371 0 0.0812f
C23410 VGND.n2590 0 0.139f
C23411 VGND.n2591 0 0.077f
C23412 VGND.n2592 0 0.0563f
C23413 VGND.t8 0 0.0792f
C23414 VGND.n2593 0 0.0547f
C23415 VGND.n2594 0 0.025f
C23416 VGND.n2595 0 0.0868f
C23417 VGND.n2596 0 0.00981f
C23418 VGND.n2597 0 0.0151f
C23419 VGND.n2598 0 0.00819f
C23420 VGND.n2599 0 0.00765f
C23421 VGND.n2600 0 0.0213f
C23422 VGND.t174 0 0.158f
C23423 VGND.n2601 0 0.185f
C23424 VGND.n2602 0 0.0613f
C23425 VGND.n2603 0 0.0888f
C23426 VGND.n2604 0 0.00828f
C23427 VGND.n2605 0 0.0162f
C23428 VGND.n2606 0 0.0106f
C23429 VGND.n2607 0 0.0149f
C23430 VGND.n2608 0 0.00837f
C23431 VGND.n2609 0 0.00828f
C23432 VGND.n2610 0 0.0422f
C23433 VGND.n2611 0 0.055f
C23434 VGND.n2612 0 0.00981f
C23435 VGND.n2613 0 0.0166f
C23436 VGND.n2614 0 0.0166f
C23437 VGND.n2615 0 0.0345f
C23438 VGND.n2616 0 0.0252f
C23439 VGND.n2617 0 0.0166f
C23440 VGND.n2618 0 0.0316f
C23441 VGND.n2619 0 0.0166f
C23442 VGND.n2620 0 0.015f
C23443 VGND.n2621 0 0.011f
C23444 VGND.n2622 0 0.0551f
C23445 VGND.t355 0 0.124f
C23446 VGND.n2623 0 0.125f
C23447 VGND.n2624 0 0.0251f
C23448 VGND.n2625 0 0.0243f
C23449 VGND.n2626 0 0.015f
C23450 VGND.n2627 0 0.0081f
C23451 VGND.n2628 0 0.00783f
C23452 VGND.n2629 0 0.00171f
C23453 VGND.n2630 0 0.00162f
C23454 VGND.n2631 0 9.9e-19
C23455 VGND.n2632 0 0.00189f
C23456 VGND.n2633 0 0.00162f
C23457 VGND.n2634 0 0.00162f
C23458 VGND.n2635 0 0.00315f
C23459 VGND.n2636 0 0.00207f
C23460 VGND.n2637 0 7.2e-19
C23461 VGND.n2638 0 7.2e-19
C23462 VGND.n2639 0 0.00162f
C23463 VGND.n2640 0 0.00198f
C23464 VGND.n2641 0 1.46e-19
C23465 VGND.n2642 0 0.00185f
C23466 VGND.n2643 0 9.77e-19
C23467 VGND.n2644 0 0.0251f
C23468 VGND.n2645 0 0.131f
C23469 VGND.n2646 0 0.184f
C23470 VGND.t208 0 0.0812f
C23471 VGND.n2647 0 0.139f
C23472 VGND.n2648 0 0.03f
C23473 VGND.n2649 0 0.009f
C23474 VGND.n2650 0 0.0163f
C23475 VGND.n2651 0 0.00828f
C23476 VGND.n2652 0 0.0105f
C23477 VGND.n2653 0 0.0505f
C23478 VGND.n2654 0 0.015f
C23479 VGND.n2655 0 0.00546f
C23480 VGND.n2656 0 0.0166f
C23481 VGND.n2657 0 0.00981f
C23482 VGND.n2658 0 0.0497f
C23483 VGND.n2659 0 0.0454f
C23484 VGND.n2660 0 0.015f
C23485 VGND.n2661 0 0.0331f
C23486 VGND.n2662 0 0.0166f
C23487 VGND.n2663 0 0.0166f
C23488 VGND.n2664 0 0.00981f
C23489 VGND.n2665 0 0.00828f
C23490 VGND.n2666 0 0.00588f
C23491 VGND.n2667 0 0.033f
C23492 VGND.n2668 0 0.015f
C23493 VGND.n2669 0 0.0191f
C23494 VGND.n2670 0 0.0166f
C23495 VGND.n2671 0 0.0334f
C23496 VGND.n2672 0 0.0166f
C23497 VGND.n2673 0 0.00418f
C23498 VGND.n2674 0 0.0166f
C23499 VGND.n2675 0 0.00586f
C23500 VGND.n2676 0 0.0166f
C23501 VGND.n2677 0 0.0285f
C23502 VGND.n2678 0 0.0166f
C23503 VGND.n2679 0 0.00821f
C23504 VGND.n2680 0 0.0166f
C23505 VGND.n2681 0 0.00586f
C23506 VGND.n2682 0 0.0166f
C23507 VGND.n2683 0 0.0155f
C23508 VGND.n2684 0 0.0166f
C23509 VGND.n2685 0 0.0361f
C23510 VGND.n2686 0 0.0166f
C23511 VGND.n2687 0 0.00583f
C23512 VGND.n2688 0 0.0166f
C23513 VGND.n2689 0 0.0341f
C23514 VGND.n2690 0 0.0166f
C23515 VGND.n2691 0 0.0372f
C23516 VGND.n2692 0 0.0166f
C23517 VGND.n2693 0 0.0511f
C23518 VGND.n2694 0 0.0166f
C23519 VGND.t300 0 0.0792f
C23520 VGND.n2695 0 0.0509f
C23521 VGND.n2696 0 0.0314f
C23522 VGND.n2697 0 0.0153f
C23523 VGND.n2698 0 0.0127f
C23524 VGND.n2699 0 0.00828f
C23525 VGND.n2700 0 0.00153f
C23526 VGND.n2701 0 0.00423f
C23527 VGND.n2702 0 0.00126f
C23528 VGND.n2703 0 0.00912f
C23529 VGND.n2704 0 0.0101f
C23530 VGND.n2705 0 0.00126f
C23531 VGND.n2706 0 0.00824f
C23532 VGND.n2707 0 0.00234f
C23533 VGND.n2708 0 0.00297f
C23534 VGND.n2709 0 0.00315f
C23535 VGND.n2710 0 0.00207f
C23536 VGND.n2711 0 9.9e-19
C23537 VGND.n2712 0 0.00261f
C23538 VGND.n2713 0 0.00207f
C23539 VGND.n2714 0 0.00135f
C23540 VGND.n2715 0 7.2e-19
C23541 VGND.n2716 0 0.00126f
C23542 VGND.n2717 0 0.00135f
C23543 VGND.n2718 0 0.00126f
C23544 VGND.n2719 0 0.0379f
C23545 VGND.n2720 0 0.00198f
C23546 VGND.n2721 0 0.00954f
C23547 VGND.n2722 0 0.00153f
C23548 VGND.n2723 0 0.00282f
C23549 VGND.n2724 0 0.00144f
C23550 VGND.n2725 0 0.00651f
C23551 VGND.n2726 0 0.00261f
C23552 VGND.n2727 0 0.00234f
C23553 VGND.n2728 0 0.00234f
C23554 VGND.n2729 0 0.00225f
C23555 VGND.n2730 0 0.00144f
C23556 VGND.n2731 0 0.00148f
C23557 VGND.n2732 0 8.57e-19
C23558 VGND.n2733 0 0.0252f
C23559 VGND.n2734 0 0.229f
C23560 VGND.n2735 0 0.184f
C23561 VGND.n2736 0 0.009f
C23562 VGND.t32 0 0.128f
C23563 VGND.n2737 0 0.198f
C23564 VGND.n2738 0 0.0532f
C23565 VGND.n2739 0 0.0304f
C23566 VGND.n2740 0 0.0278f
C23567 VGND.n2741 0 0.013f
C23568 VGND.t365 0 0.0812f
C23569 VGND.n2742 0 0.139f
C23570 VGND.t179 0 0.0445f
C23571 VGND.n2743 0 0.14f
C23572 VGND.t234 0 0.0445f
C23573 VGND.t350 0 0.0445f
C23574 VGND.n2744 0 0.243f
C23575 VGND.n2745 0 0.0173f
C23576 VGND.n2746 0 0.019f
C23577 VGND.n2747 0 0.0275f
C23578 VGND.n2748 0 0.0383f
C23579 VGND.n2749 0 0.0166f
C23580 VGND.n2750 0 0.00596f
C23581 VGND.n2751 0 0.0166f
C23582 VGND.n2752 0 0.015f
C23583 VGND.n2753 0 0.00553f
C23584 VGND.n2754 0 0.0693f
C23585 VGND.n2755 0 0.00981f
C23586 VGND.n2756 0 0.0321f
C23587 VGND.n2757 0 0.0271f
C23588 VGND.n2758 0 0.0166f
C23589 VGND.t21 0 0.0946f
C23590 VGND.n2759 0 0.0183f
C23591 VGND.n2760 0 0.0961f
C23592 VGND.n2761 0 0.0252f
C23593 VGND.n2762 0 0.0271f
C23594 VGND.n2763 0 0.0166f
C23595 VGND.n2764 0 0.0345f
C23596 VGND.n2765 0 0.0252f
C23597 VGND.n2766 0 0.0166f
C23598 VGND.n2767 0 0.0453f
C23599 VGND.n2768 0 0.0166f
C23600 VGND.n2769 0 0.0421f
C23601 VGND.n2770 0 0.0166f
C23602 VGND.n2771 0 0.0166f
C23603 VGND.n2772 0 0.0331f
C23604 VGND.n2773 0 0.037f
C23605 VGND.n2774 0 0.015f
C23606 VGND.n2775 0 0.00981f
C23607 VGND.n2776 0 0.00453f
C23608 VGND.n2777 0 0.0166f
C23609 VGND.n2778 0 0.0124f
C23610 VGND.n2779 0 0.0166f
C23611 VGND.n2780 0 0.015f
C23612 VGND.n2781 0 0.0119f
C23613 VGND.n2782 0 0.0451f
C23614 VGND.n2783 0 0.00828f
C23615 VGND.n2784 0 0.0163f
C23616 VGND.n2785 0 0.0628f
C23617 VGND.t315 0 0.0812f
C23618 VGND.n2786 0 0.139f
C23619 VGND.n2787 0 0.0301f
C23620 VGND.n2788 0 0.0452f
C23621 VGND.n2789 0 0.00972f
C23622 VGND.t380 0 0.0792f
C23623 VGND.n2790 0 0.0547f
C23624 VGND.n2791 0 0.0243f
C23625 VGND.n2792 0 0.0166f
C23626 VGND.n2793 0 0.0166f
C23627 VGND.n2794 0 0.015f
C23628 VGND.n2795 0 0.00828f
C23629 VGND.n2796 0 0.0442f
C23630 VGND.n2797 0 0.0483f
C23631 VGND.n2798 0 0.0321f
C23632 VGND.n2799 0 0.0271f
C23633 VGND.t286 0 0.0946f
C23634 VGND.n2800 0 0.0192f
C23635 VGND.n2801 0 0.0961f
C23636 VGND.n2802 0 0.0298f
C23637 VGND.n2803 0 0.0472f
C23638 VGND.n2804 0 0.015f
C23639 VGND.n2805 0 0.0221f
C23640 VGND.n2806 0 0.0081f
C23641 VGND.n2807 0 0.0106f
C23642 VGND.n2808 0 0.00376f
C23643 VGND.n2809 0 0.0166f
C23644 VGND.n2810 0 0.0166f
C23645 VGND.n2811 0 0.00462f
C23646 VGND.n2812 0 0.0166f
C23647 VGND.n2813 0 0.00586f
C23648 VGND.n2814 0 0.0166f
C23649 VGND.n2815 0 0.00437f
C23650 VGND.n2816 0 0.0166f
C23651 VGND.n2817 0 0.0149f
C23652 VGND.n2818 0 0.00837f
C23653 VGND.n2819 0 0.00819f
C23654 VGND.n2820 0 0.0567f
C23655 VGND.n2821 0 0.00837f
C23656 VGND.n2822 0 0.0137f
C23657 VGND.t232 0 0.082f
C23658 VGND.n2823 0 0.0934f
C23659 VGND.n2824 0 0.0261f
C23660 VGND.n2825 0 0.0191f
C23661 VGND.n2826 0 0.0063f
C23662 VGND.n2827 0 0.00824f
C23663 VGND.n2828 0 0.00413f
C23664 VGND.n2829 0 0.018f
C23665 VGND.n2830 0 0.00269f
C23666 VGND.n2831 0 0.00207f
C23667 VGND.n2832 0 0.00287f
C23668 VGND.n2833 0 0.00173f
C23669 VGND.n2835 0 0.317f
C23670 VGND.n2836 0 0.317f
C23671 VGND.n2837 0 0.00207f
C23672 VGND.n2838 0 0.00287f
C23673 VGND.n2839 0 0.0039f
C23674 VGND.n2840 0 0.00269f
C23675 VGND.n2841 0 0.00173f
C23676 VGND.n2843 0 0.018f
C23677 VGND.n2844 0 0.00274f
C23678 VGND.n2845 0 0.00173f
C23679 VGND.n2846 0 0.00413f
C23680 VGND.n2847 0 0.00824f
C23681 VGND.n2848 0 0.0063f
C23682 VGND.n2849 0 0.00765f
C23683 VGND.n2850 0 0.00405f
C23684 VGND.n2851 0 0.0155f
C23685 VGND.n2852 0 0.059f
C23686 VGND.n2853 0 0.0597f
C23687 VGND.n2854 0 0.0878f
C23688 VGND.n2855 0 0.0142f
C23689 VGND.n2856 0 0.0166f
C23690 VGND.n2857 0 0.0166f
C23691 VGND.n2858 0 0.059f
C23692 VGND.n2859 0 0.0166f
C23693 VGND.n2860 0 0.0449f
C23694 VGND.n2861 0 0.0166f
C23695 VGND.t43 0 0.155f
C23696 VGND.n2862 0 0.163f
C23697 VGND.t167 0 0.148f
C23698 VGND.n2863 0 0.093f
C23699 VGND.n2864 0 0.07f
C23700 VGND.n2865 0 0.0147f
C23701 VGND.n2866 0 0.0166f
C23702 VGND.n2867 0 0.0482f
C23703 VGND.n2868 0 0.00981f
C23704 VGND.n2869 0 0.00828f
C23705 VGND.n2870 0 0.0105f
C23706 VGND.n2871 0 0.0287f
C23707 VGND.n2872 0 0.015f
C23708 VGND.n2873 0 0.0279f
C23709 VGND.n2874 0 0.0166f
C23710 VGND.n2875 0 0.00236f
C23711 VGND.n2876 0 0.00963f
C23712 VGND.n2877 0 0.0152f
C23713 VGND.n2878 0 0.0373f
C23714 VGND.n2879 0 0.0331f
C23715 VGND.t196 0 0.0792f
C23716 VGND.n2880 0 0.0552f
C23717 VGND.n2881 0 0.0243f
C23718 VGND.n2882 0 0.0166f
C23719 VGND.n2883 0 0.00981f
C23720 VGND.n2884 0 0.00828f
C23721 VGND.n2885 0 0.00509f
C23722 VGND.n2886 0 0.0582f
C23723 VGND.n2887 0 0.02f
C23724 VGND.n2888 0 0.00963f
C23725 VGND.n2889 0 0.0121f
C23726 VGND.n2890 0 0.045f
C23727 VGND.t101 0 0.128f
C23728 VGND.n2891 0 0.155f
C23729 VGND.n2892 0 0.0839f
C23730 VGND.n2893 0 0.00828f
C23731 VGND.n2894 0 0.0172f
C23732 VGND.t173 0 0.0837f
C23733 VGND.n2895 0 0.185f
C23734 VGND.n2896 0 0.0245f
C23735 VGND.n2897 0 0.0294f
C23736 VGND.n2898 0 0.0166f
C23737 VGND.t197 0 0.0792f
C23738 VGND.n2899 0 0.0547f
C23739 VGND.n2900 0 0.00513f
C23740 VGND.n2901 0 0.0166f
C23741 VGND.n2902 0 0.037f
C23742 VGND.n2903 0 0.0166f
C23743 VGND.t57 0 0.0792f
C23744 VGND.n2904 0 0.00463f
C23745 VGND.n2905 0 0.0269f
C23746 VGND.n2906 0 0.0232f
C23747 VGND.n2907 0 0.0251f
C23748 VGND.t326 0 0.0445f
C23749 VGND.n2908 0 0.0166f
C23750 VGND.t303 0 0.0445f
C23751 VGND.n2909 0 0.244f
C23752 VGND.n2910 0 0.00405f
C23753 VGND.n2911 0 0.0104f
C23754 VGND.n2912 0 0.0166f
C23755 VGND.n2913 0 0.0166f
C23756 VGND.n2914 0 0.015f
C23757 VGND.n2915 0 0.00981f
C23758 VGND.n2916 0 0.0291f
C23759 VGND.n2917 0 0.0689f
C23760 VGND.n2918 0 0.0352f
C23761 VGND.n2919 0 0.0331f
C23762 VGND.n2920 0 0.0166f
C23763 VGND.n2921 0 0.0166f
C23764 VGND.n2922 0 0.0166f
C23765 VGND.n2923 0 0.0304f
C23766 VGND.n2924 0 0.02f
C23767 VGND.n2925 0 0.0321f
C23768 VGND.n2926 0 0.0166f
C23769 VGND.n2927 0 0.0149f
C23770 VGND.n2928 0 0.00837f
C23771 VGND.n2929 0 0.0246f
C23772 VGND.n2930 0 0.0281f
C23773 VGND.n2931 0 0.00981f
C23774 VGND.n2932 0 0.0166f
C23775 VGND.n2933 0 0.0243f
C23776 VGND.n2934 0 0.0387f
C23777 VGND.n2935 0 0.0569f
C23778 VGND.n2936 0 0.015f
C23779 VGND.n2937 0 0.00981f
C23780 VGND.n2938 0 0.015f
C23781 VGND.n2939 0 0.00828f
C23782 VGND.n2940 0 0.0037f
C23783 VGND.n2941 0 0.0411f
C23784 VGND.n2942 0 0.00828f
C23785 VGND.n2943 0 0.022f
C23786 VGND.n2944 0 0.00837f
C23787 VGND.n2945 0 0.0292f
C23788 VGND.n2946 0 0.229f
C23789 VGND.n2947 0 0.0935f
C23790 VGND.n2948 0 0.0257f
C23791 VGND.n2949 0 8.57e-19
C23792 VGND.n2950 0 0.00126f
C23793 VGND.n2951 0 0.00135f
C23794 VGND.n2952 0 0.00126f
C23795 VGND.n2953 0 7.2e-19
C23796 VGND.n2954 0 9.9e-19
C23797 VGND.n2955 0 0.00207f
C23798 VGND.n2956 0 0.00315f
C23799 VGND.n2957 0 0.00297f
C23800 VGND.n2958 0 0.00234f
C23801 VGND.n2959 0 0.00824f
C23802 VGND.n2960 0 0.00912f
C23803 VGND.n2961 0 0.025f
C23804 VGND.n2962 0 0.00126f
C23805 VGND.n2963 0 0.00153f
C23806 VGND.n2964 0 0.0127f
C23807 VGND.n2965 0 0.00828f
C23808 VGND.t41 0 0.0792f
C23809 VGND.n2966 0 0.0509f
C23810 VGND.n2967 0 0.0243f
C23811 VGND.n2968 0 0.0153f
C23812 VGND.n2969 0 0.0331f
C23813 VGND.n2970 0 0.0166f
C23814 VGND.n2971 0 0.015f
C23815 VGND.n2972 0 0.0379f
C23816 VGND.n2973 0 0.00485f
C23817 VGND.n2974 0 0.00981f
C23818 VGND.n2975 0 0.0166f
C23819 VGND.n2976 0 0.015f
C23820 VGND.n2977 0 0.00485f
C23821 VGND.n2978 0 0.0291f
C23822 VGND.n2979 0 0.00981f
C23823 VGND.n2980 0 0.0166f
C23824 VGND.n2981 0 0.0515f
C23825 VGND.n2982 0 0.0166f
C23826 VGND.n2983 0 0.015f
C23827 VGND.n2984 0 0.038f
C23828 VGND.n2985 0 0.0287f
C23829 VGND.n2986 0 0.0547f
C23830 VGND.n2987 0 0.0445f
C23831 VGND.n2988 0 0.0166f
C23832 VGND.n2989 0 0.0166f
C23833 VGND.n2990 0 0.015f
C23834 VGND.n2991 0 0.0546f
C23835 VGND.n2992 0 0.045f
C23836 VGND.n2993 0 0.00981f
C23837 VGND.n2994 0 0.0166f
C23838 VGND.n2995 0 0.015f
C23839 VGND.n2996 0 0.0375f
C23840 VGND.n2997 0 0.0287f
C23841 VGND.n2998 0 0.00981f
C23842 VGND.n2999 0 0.0166f
C23843 VGND.n3000 0 0.0358f
C23844 VGND.n3001 0 0.0166f
C23845 VGND.n3002 0 0.0602f
C23846 VGND.n3003 0 0.0149f
C23847 VGND.n3004 0 0.00828f
C23848 VGND.n3005 0 0.00507f
C23849 VGND.n3006 0 0.0467f
C23850 VGND.n3007 0 0.00981f
C23851 VGND.t77 0 0.0792f
C23852 VGND.n3008 0 0.0551f
C23853 VGND.n3009 0 0.0243f
C23854 VGND.n3010 0 0.0166f
C23855 VGND.n3011 0 0.0166f
C23856 VGND.n3012 0 0.0143f
C23857 VGND.n3013 0 0.009f
C23858 VGND.n3014 0 0.026f
C23859 VGND.n3015 0 0.0279f
C23860 VGND.n3016 0 0.00981f
C23861 VGND.t125 0 0.0792f
C23862 VGND.n3017 0 0.0547f
C23863 VGND.n3018 0 0.0243f
C23864 VGND.n3019 0 0.0166f
C23865 VGND.n3020 0 0.0166f
C23866 VGND.n3021 0 0.015f
C23867 VGND.n3022 0 0.0474f
C23868 VGND.n3023 0 0.0182f
C23869 VGND.n3024 0 0.00981f
C23870 VGND.n3025 0 0.0166f
C23871 VGND.n3026 0 0.00446f
C23872 VGND.n3027 0 0.0166f
C23873 VGND.n3028 0 0.0166f
C23874 VGND.n3029 0 0.0268f
C23875 VGND.n3030 0 0.0166f
C23876 VGND.n3031 0 0.00821f
C23877 VGND.n3032 0 0.0166f
C23878 VGND.n3033 0 0.00586f
C23879 VGND.n3034 0 0.0166f
C23880 VGND.n3035 0 0.00504f
C23881 VGND.n3036 0 0.0166f
C23882 VGND.n3037 0 0.0166f
C23883 VGND.n3038 0 0.015f
C23884 VGND.n3039 0 0.00797f
C23885 VGND.n3040 0 0.0488f
C23886 VGND.n3041 0 0.00981f
C23887 VGND.t124 0 0.0792f
C23888 VGND.n3042 0 0.0547f
C23889 VGND.n3043 0 0.0243f
C23890 VGND.n3044 0 0.0166f
C23891 VGND.n3045 0 0.0166f
C23892 VGND.n3046 0 0.0151f
C23893 VGND.n3047 0 0.0384f
C23894 VGND.n3048 0 0.0535f
C23895 VGND.n3049 0 0.00972f
C23896 VGND.n3050 0 0.0142f
C23897 VGND.n3051 0 0.0166f
C23898 VGND.n3052 0 0.0238f
C23899 VGND.n3053 0 0.0166f
C23900 VGND.n3054 0 0.00835f
C23901 VGND.n3055 0 0.0166f
C23902 VGND.n3056 0 0.015f
C23903 VGND.n3057 0 0.00828f
C23904 VGND.n3058 0 0.0127f
C23905 VGND.t99 0 0.0813f
C23906 VGND.n3059 0 0.139f
C23907 VGND.n3060 0 0.0349f
C23908 VGND.n3061 0 0.0118f
C23909 VGND.n3062 0 0.0136f
C23910 VGND.n3063 0 0.00207f
C23911 VGND.n3064 0 0.00315f
C23912 VGND.n3065 0 0.00162f
C23913 VGND.n3066 0 0.00162f
C23914 VGND.n3067 0 0.00189f
C23915 VGND.n3068 0 9.9e-19
C23916 VGND.n3069 0 0.00162f
C23917 VGND.n3070 0 0.00171f
C23918 VGND.n3071 0 9.9e-19
C23919 VGND.n3072 0 0.00189f
C23920 VGND.n3073 0 0.00162f
C23921 VGND.n3074 0 0.00342f
C23922 VGND.n3075 0 0.00387f
C23923 VGND.n3076 0 7.2e-19
C23924 VGND.n3077 0 0.00162f
C23925 VGND.n3078 0 0.00207f
C23926 VGND.n3079 0 0.00207f
C23927 VGND.n3080 0 0.00162f
C23928 VGND.n3081 0 0.00234f
C23929 VGND.n3082 0 0.00234f
C23930 VGND.n3083 0 0.00234f
C23931 VGND.n3084 0 0.00297f
C23932 VGND.n3085 0 0.00144f
C23933 VGND.n3086 0 0.00135f
C23934 VGND.n3087 0 2.7e-19
C23935 VGND.n3088 0 0.00126f
C23936 VGND.n3089 0 0.00207f
C23937 VGND.n3090 0 0.00126f
C23938 VGND.n3091 0 0.00126f
C23939 VGND.n3092 0 0.00701f
C23940 VGND.n3093 0 0.0041f
C23941 VGND.n3094 0 0.018f
C23942 VGND.n3095 0 0.00287f
C23943 VGND.n3096 0 0.00207f
C23944 VGND.n3097 0 0.00274f
C23945 VGND.n3098 0 0.00403f
C23946 VGND.n3099 0 0.00493f
C23947 VGND.n3100 0 0.00126f
C23948 VGND.n3101 0 0.00173f
C23949 VGND.n3103 0 0.317f
C23950 VGND.n3104 0 0.317f
C23951 VGND.n3105 0 0.00207f
C23952 VGND.n3106 0 0.00287f
C23953 VGND.n3107 0 0.00173f
C23954 VGND.n3108 0 0.00269f
C23955 VGND.n3109 0 0.0039f
C23956 VGND.n3110 0 0.00269f
C23957 VGND.n3111 0 0.00173f
C23958 VGND.n3113 0 0.317f
C23959 VGND.n3114 0 0.317f
C23960 VGND.n3115 0 0.00287f
C23961 VGND.n3116 0 0.00207f
C23962 VGND.n3117 0 0.00274f
C23963 VGND.n3118 0 0.00403f
C23964 VGND.n3119 0 0.00493f
C23965 VGND.n3120 0 0.00126f
C23966 VGND.n3121 0 0.00173f
C23967 VGND.n3123 0 0.018f
C23968 VGND.n3124 0 0.00274f
C23969 VGND.n3125 0 0.00173f
C23970 VGND.n3126 0 0.0041f
C23971 VGND.n3127 0 0.00701f
C23972 VGND.n3128 0 0.00207f
C23973 VGND.n3129 0 0.00207f
C23974 VGND.n3130 0 0.00162f
C23975 VGND.n3131 0 0.00234f
C23976 VGND.n3132 0 0.00126f
C23977 VGND.n3133 0 2.7e-19
C23978 VGND.n3134 0 0.00135f
C23979 VGND.n3135 0 0.00144f
C23980 VGND.n3136 0 0.00297f
C23981 VGND.n3137 0 5.1e-19
C23982 VGND.n3138 0 0.00135f
C23983 VGND.n3139 0 0.00186f
C23984 VGND.n3140 0 8.1e-19
C23985 VGND.n3141 0 0.00234f
C23986 VGND.n3142 0 0.00234f
C23987 VGND.n3143 0 0.00234f
C23988 VGND.n3144 0 7.2e-19
C23989 VGND.n3145 0 0.00252f
C23990 VGND.n3146 0 0.00369f
C23991 VGND.n3147 0 0.00189f
C23992 VGND.n3148 0 0.00135f
C23993 VGND.n3149 0 0.00207f
C23994 VGND.n3150 0 0.00126f
C23995 VGND.n3151 0 0.00126f
C23996 VGND.n3152 0 0.00603f
C23997 VGND.t271 0 0.155f
C23998 VGND.t14 0 0.155f
C23999 VGND.n3153 0 0.297f
C24000 VGND.n3154 0 0.0151f
C24001 VGND.n3155 0 0.00545f
C24002 VGND.n3156 0 0.05f
C24003 VGND.n3157 0 0.0439f
C24004 VGND.n3158 0 0.014f
C24005 VGND.n3159 0 0.0449f
C24006 VGND.n3160 0 0.0166f
C24007 VGND.n3161 0 0.059f
C24008 VGND.n3162 0 0.0166f
C24009 VGND.n3163 0 0.059f
C24010 VGND.n3164 0 0.0166f
C24011 VGND.n3165 0 0.059f
C24012 VGND.n3166 0 0.0166f
C24013 VGND.n3167 0 0.0604f
C24014 VGND.n3168 0 0.0166f
C24015 VGND.n3169 0 0.0685f
C24016 VGND.n3170 0 0.0144f
C24017 VGND.n3171 0 0.0104f
C24018 VGND.n3172 0 0.0149f
C24019 VGND.n3173 0 0.0374f
C24020 VGND.n3174 0 0.0332f
C24021 VGND.n3175 0 0.0281f
C24022 VGND.n3176 0 0.00981f
C24023 VGND.n3177 0 0.0166f
C24024 VGND.n3178 0 0.0795f
C24025 VGND.n3179 0 0.0166f
C24026 VGND.n3180 0 0.015f
C24027 VGND.n3181 0 0.0362f
C24028 VGND.n3182 0 0.0371f
C24029 VGND.n3183 0 0.0459f
C24030 VGND.n3184 0 0.012f
C24031 VGND.n3185 0 0.0112f
C24032 VGND.n3186 0 0.0104f
C24033 VGND.n3187 0 0.028f
C24034 VGND.n3188 0 0.0619f
C24035 VGND.n3189 0 0.0471f
C24036 VGND.n3190 0 0.0319f
C24037 VGND.n3191 0 0.0283f
C24038 VGND.n3192 0 0.00981f
C24039 VGND.n3193 0 0.0166f
C24040 VGND.n3194 0 0.0334f
C24041 VGND.n3195 0 0.0166f
C24042 VGND.n3196 0 0.0143f
C24043 VGND.n3197 0 0.0603f
C24044 VGND.n3198 0 0.0254f
C24045 VGND.n3199 0 0.229f
C24046 VGND.n3200 0 0.319f
C24047 VGND.n3201 0 0.0191f
C24048 VGND.n3202 0 7.2e-19
C24049 VGND.n3203 0 0.0118f
C24050 VGND.n3204 0 0.00198f
C24051 VGND.n3205 0 0.00162f
C24052 VGND.n3206 0 0.00189f
C24053 VGND.n3207 0 0.00162f
C24054 VGND.n3208 0 0.00342f
C24055 VGND.n3209 0 0.00387f
C24056 VGND.n3210 0 7.2e-19
C24057 VGND.n3211 0 7.2e-19
C24058 VGND.n3212 0 0.00207f
C24059 VGND.n3213 0 0.00315f
C24060 VGND.n3214 0 0.00162f
C24061 VGND.n3215 0 0.00162f
C24062 VGND.n3216 0 0.00189f
C24063 VGND.n3217 0 9.9e-19
C24064 VGND.n3218 0 0.00162f
C24065 VGND.n3219 0 0.00171f
C24066 VGND.n3220 0 0.00783f
C24067 VGND.n3221 0 0.0331f
C24068 VGND.n3222 0 0.0148f
C24069 VGND.n3223 0 0.0273f
C24070 VGND.n3224 0 0.0275f
C24071 VGND.n3225 0 0.019f
C24072 VGND.n3226 0 0.0494f
C24073 VGND.n3227 0 0.025f
C24074 VGND.n3228 0 0.015f
C24075 VGND.n3229 0 0.0245f
C24076 VGND.n3230 0 0.0114f
C24077 VGND.n3231 0 0.0166f
C24078 VGND.n3232 0 0.0306f
C24079 VGND.n3233 0 0.00478f
C24080 VGND.n3234 0 0.0223f
C24081 VGND.n3235 0 0.00108f
C24082 VGND.n3236 0 0.0166f
C24083 VGND.n3237 0 0.00819f
C24084 VGND.n3238 0 0.0663f
C24085 VGND.n3239 0 0.028f
C24086 VGND.n3240 0 0.009f
C24087 VGND.n3241 0 0.0112f
C24088 VGND.n3242 0 0.045f
C24089 VGND.t218 0 0.128f
C24090 VGND.n3243 0 0.157f
C24091 VGND.n3244 0 0.0772f
C24092 VGND.n3245 0 0.026f
C24093 VGND.n3246 0 0.0191f
C24094 VGND.n3247 0 0.00819f
C24095 VGND.n3248 0 0.0543f
C24096 VGND.n3249 0 0.0499f
C24097 VGND.n3250 0 0.0429f
C24098 VGND.n3251 0 0.0151f
C24099 VGND.n3252 0 0.0166f
C24100 VGND.t47 0 0.0792f
C24101 VGND.n3253 0 0.0547f
C24102 VGND.n3254 0 0.0243f
C24103 VGND.n3255 0 0.0166f
C24104 VGND.n3256 0 0.00972f
C24105 VGND.n3257 0 0.046f
C24106 VGND.n3258 0 0.0371f
C24107 VGND.n3259 0 0.0528f
C24108 VGND.n3260 0 0.015f
C24109 VGND.n3261 0 0.0166f
C24110 VGND.t235 0 0.0792f
C24111 VGND.n3262 0 0.0591f
C24112 VGND.n3263 0 0.0382f
C24113 VGND.n3264 0 0.0166f
C24114 VGND.n3265 0 0.0279f
C24115 VGND.n3266 0 0.00981f
C24116 VGND.n3267 0 0.009f
C24117 VGND.n3268 0 0.0439f
C24118 VGND.n3269 0 0.00376f
C24119 VGND.n3270 0 0.0143f
C24120 VGND.n3271 0 0.0106f
C24121 VGND.n3272 0 0.025f
C24122 VGND.n3273 0 0.042f
C24123 VGND.n3274 0 0.0142f
C24124 VGND.n3275 0 0.046f
C24125 VGND.n3276 0 0.0166f
C24126 VGND.n3277 0 0.0393f
C24127 VGND.n3278 0 0.0166f
C24128 VGND.n3279 0 0.0424f
C24129 VGND.n3280 0 0.0166f
C24130 VGND.n3281 0 0.0458f
C24131 VGND.n3282 0 0.0252f
C24132 VGND.n3283 0 0.0166f
C24133 VGND.n3284 0 0.0166f
C24134 VGND.n3285 0 0.0166f
C24135 VGND.n3286 0 0.00981f
C24136 VGND.n3287 0 0.00837f
C24137 VGND.n3288 0 0.0263f
C24138 VGND.n3289 0 0.0331f
C24139 VGND.n3290 0 0.0149f
C24140 VGND.n3291 0 0.0251f
C24141 VGND.n3292 0 0.0166f
C24142 VGND.n3293 0 0.0289f
C24143 VGND.n3294 0 0.0166f
C24144 VGND.n3295 0 0.00981f
C24145 VGND.n3296 0 0.0268f
C24146 VGND.n3297 0 0.0367f
C24147 VGND.n3298 0 0.015f
C24148 VGND.n3299 0 0.0331f
C24149 VGND.n3300 0 0.0166f
C24150 VGND.t139 0 0.0799f
C24151 VGND.n3301 0 0.0723f
C24152 VGND.n3302 0 0.0241f
C24153 VGND.n3303 0 0.0166f
C24154 VGND.n3304 0 0.00981f
C24155 VGND.n3305 0 0.0192f
C24156 VGND.t225 0 0.0792f
C24157 VGND.n3306 0 0.057f
C24158 VGND.n3307 0 0.0249f
C24159 VGND.n3308 0 0.0825f
C24160 VGND.n3309 0 0.00828f
C24161 VGND.n3310 0 0.015f
C24162 VGND.n3311 0 0.00981f
C24163 VGND.n3312 0 0.00837f
C24164 VGND.n3313 0 0.0375f
C24165 VGND.n3314 0 0.0331f
C24166 VGND.n3315 0 0.0149f
C24167 VGND.n3316 0 0.0273f
C24168 VGND.n3317 0 0.0284f
C24169 VGND.n3318 0 0.0166f
C24170 VGND.n3319 0 0.0145f
C24171 VGND.n3320 0 0.00824f
C24172 VGND.n3321 0 0.00234f
C24173 VGND.n3322 0 0.00297f
C24174 VGND.n3323 0 0.00315f
C24175 VGND.n3324 0 0.00207f
C24176 VGND.n3325 0 9.9e-19
C24177 VGND.n3326 0 0.00261f
C24178 VGND.n3327 0 0.00207f
C24179 VGND.n3328 0 0.00135f
C24180 VGND.n3329 0 7.2e-19
C24181 VGND.n3330 0 0.00126f
C24182 VGND.n3331 0 0.00135f
C24183 VGND.n3332 0 0.00126f
C24184 VGND.n3333 0 0.0254f
C24185 VGND.n3334 0 0.00198f
C24186 VGND.n3335 0 0.00453f
C24187 VGND.n3336 0 0.00153f
C24188 VGND.n3337 0 0.00282f
C24189 VGND.n3338 0 0.00144f
C24190 VGND.n3339 0 0.00651f
C24191 VGND.n3340 0 0.00261f
C24192 VGND.n3341 0 0.00234f
C24193 VGND.n3342 0 0.00234f
C24194 VGND.n3343 0 0.00225f
C24195 VGND.n3344 0 0.00144f
C24196 VGND.n3345 0 0.00148f
C24197 VGND.n3346 0 8.57e-19
C24198 VGND.n3347 0 0.0246f
C24199 VGND.n3348 0 0.229f
C24200 VGND.n3349 0 0.049f
C24201 VGND.n3350 0 0.03f
C24202 VGND.t201 0 0.124f
C24203 VGND.t217 0 0.0837f
C24204 VGND.n3351 0 0.0438f
C24205 VGND.n3352 0 0.0457f
C24206 VGND.n3353 0 0.039f
C24207 VGND.n3354 0 0.0199f
C24208 VGND.n3355 0 0.0457f
C24209 VGND.n3356 0 0.0122f
C24210 VGND.t39 0 0.0812f
C24211 VGND.n3357 0 0.139f
C24212 VGND.t231 0 0.0445f
C24213 VGND.n3358 0 0.14f
C24214 VGND.t278 0 0.0445f
C24215 VGND.t247 0 0.0445f
C24216 VGND.n3359 0 0.243f
C24217 VGND.n3360 0 0.0173f
C24218 VGND.n3361 0 0.0172f
C24219 VGND.n3362 0 0.00981f
C24220 VGND.n3363 0 0.0395f
C24221 VGND.n3364 0 0.0166f
C24222 VGND.n3365 0 0.00707f
C24223 VGND.n3366 0 0.0166f
C24224 VGND.n3367 0 0.015f
C24225 VGND.n3368 0 0.011f
C24226 VGND.n3369 0 0.0291f
C24227 VGND.n3370 0 0.00981f
C24228 VGND.t249 0 0.0792f
C24229 VGND.n3371 0 0.0547f
C24230 VGND.n3372 0 0.0243f
C24231 VGND.n3373 0 0.0166f
C24232 VGND.n3374 0 0.0331f
C24233 VGND.n3375 0 0.0166f
C24234 VGND.n3376 0 0.0379f
C24235 VGND.n3377 0 0.0166f
C24236 VGND.n3378 0 0.0396f
C24237 VGND.n3379 0 0.0166f
C24238 VGND.n3380 0 0.015f
C24239 VGND.n3381 0 0.00828f
C24240 VGND.n3382 0 0.0339f
C24241 VGND.n3383 0 0.0283f
C24242 VGND.n3384 0 0.00981f
C24243 VGND.t341 0 0.0792f
C24244 VGND.n3385 0 0.0547f
C24245 VGND.n3386 0 0.0243f
C24246 VGND.n3387 0 0.0166f
C24247 VGND.n3388 0 0.0166f
C24248 VGND.n3389 0 0.0511f
C24249 VGND.n3390 0 0.0438f
C24250 VGND.n3391 0 0.0149f
C24251 VGND.n3392 0 0.0099f
C24252 VGND.n3393 0 0.00931f
C24253 VGND.n3394 0 0.0166f
C24254 VGND.n3395 0 0.015f
C24255 VGND.n3396 0 0.024f
C24256 VGND.n3397 0 0.0291f
C24257 VGND.n3398 0 0.00981f
C24258 VGND.t293 0 0.0792f
C24259 VGND.n3399 0 0.0689f
C24260 VGND.n3400 0 0.0293f
C24261 VGND.n3401 0 0.0166f
C24262 VGND.n3402 0 0.0166f
C24263 VGND.n3403 0 0.0143f
C24264 VGND.n3404 0 0.00828f
C24265 VGND.n3405 0 0.0229f
C24266 VGND.n3406 0 0.185f
C24267 VGND.n3407 0 0.225f
C24268 VGND.n3408 0 0.0116f
C24269 VGND.n3409 0 0.00382f
C24270 VGND.n3410 0 0.00972f
C24271 VGND.n3411 0 0.0166f
C24272 VGND.n3412 0 0.0166f
C24273 VGND.n3413 0 0.015f
C24274 VGND.n3414 0 0.00437f
C24275 VGND.n3415 0 0.0291f
C24276 VGND.n3416 0 0.00981f
C24277 VGND.t328 0 0.0792f
C24278 VGND.n3417 0 0.0547f
C24279 VGND.n3418 0 0.0243f
C24280 VGND.n3419 0 0.0166f
C24281 VGND.n3420 0 0.0689f
C24282 VGND.n3421 0 0.0166f
C24283 VGND.n3422 0 0.0443f
C24284 VGND.n3423 0 0.0166f
C24285 VGND.n3424 0 0.015f
C24286 VGND.n3425 0 0.00511f
C24287 VGND.n3426 0 0.0391f
C24288 VGND.n3427 0 0.00981f
C24289 VGND.t129 0 0.0792f
C24290 VGND.n3428 0 0.0639f
C24291 VGND.n3429 0 0.0243f
C24292 VGND.n3430 0 0.0166f
C24293 VGND.n3431 0 0.0166f
C24294 VGND.n3432 0 0.0149f
C24295 VGND.n3433 0 0.042f
C24296 VGND.n3434 0 0.0208f
C24297 VGND.n3435 0 0.0099f
C24298 VGND.n3436 0 0.0166f
C24299 VGND.n3437 0 0.014f
C24300 VGND.n3438 0 0.0166f
C24301 VGND.n3439 0 0.0166f
C24302 VGND.n3440 0 0.015f
C24303 VGND.n3441 0 0.00463f
C24304 VGND.n3442 0 0.0291f
C24305 VGND.n3443 0 0.00981f
C24306 VGND.t105 0 0.0792f
C24307 VGND.n3444 0 0.0547f
C24308 VGND.n3445 0 0.0243f
C24309 VGND.n3446 0 0.0166f
C24310 VGND.n3447 0 0.0312f
C24311 VGND.n3448 0 0.0136f
C24312 VGND.n3449 0 0.0063f
C24313 VGND.n3450 0 0.00824f
C24314 VGND.n3451 0 0.00413f
C24315 VGND.n3452 0 0.018f
C24316 VGND.n3453 0 0.00269f
C24317 VGND.n3454 0 0.00207f
C24318 VGND.n3455 0 0.00287f
C24319 VGND.n3456 0 0.00173f
C24320 VGND.n3458 0 0.317f
C24321 VGND.n3459 0 0.317f
C24322 VGND.n3460 0 0.00207f
C24323 VGND.n3461 0 0.00287f
C24324 VGND.n3462 0 0.0039f
C24325 VGND.n3463 0 0.00269f
C24326 VGND.n3464 0 0.00173f
C24327 VGND.n3466 0 0.018f
C24328 VGND.n3467 0 0.00274f
C24329 VGND.n3468 0 0.00173f
C24330 VGND.n3469 0 0.00413f
C24331 VGND.n3470 0 0.00824f
C24332 VGND.n3471 0 0.0123f
C24333 VGND.n3472 0 0.0103f
C24334 VGND.n3473 0 0.0172f
C24335 VGND.n3474 0 0.0674f
C24336 VGND.n3475 0 0.017f
C24337 VGND.n3476 0 0.015f
C24338 VGND.n3477 0 0.0444f
C24339 VGND.n3478 0 0.0166f
C24340 VGND.n3479 0 0.057f
C24341 VGND.n3480 0 0.0167f
C24342 VGND.n3481 0 0.00825f
C24343 VGND.n3482 0 0.0166f
C24344 VGND.n3483 0 0.0536f
C24345 VGND.n3484 0 0.0166f
C24346 VGND.n3485 0 0.00987f
C24347 VGND.n3486 0 0.0387f
C24348 VGND.n3487 0 0.0519f
C24349 VGND.n3488 0 0.0398f
C24350 VGND.n3489 0 0.0151f
C24351 VGND.n3490 0 0.0166f
C24352 VGND.n3491 0 0.0245f
C24353 VGND.n3492 0 0.00972f
C24354 VGND.n3493 0 0.00837f
C24355 VGND.n3494 0 0.0193f
C24356 VGND.t310 0 0.0792f
C24357 VGND.n3495 0 0.0575f
C24358 VGND.n3496 0 0.0243f
C24359 VGND.n3497 0 0.0832f
C24360 VGND.n3498 0 0.015f
C24361 VGND.n3499 0 0.0166f
C24362 VGND.n3500 0 0.00981f
C24363 VGND.n3501 0 0.0477f
C24364 VGND.n3502 0 0.0059f
C24365 VGND.n3503 0 0.015f
C24366 VGND.n3504 0 0.0166f
C24367 VGND.n3505 0 0.0245f
C24368 VGND.n3506 0 0.00586f
C24369 VGND.n3507 0 0.00891f
C24370 VGND.n3508 0 0.00981f
C24371 VGND.n3509 0 0.0144f
C24372 VGND.n3510 0 0.0561f
C24373 VGND.n3511 0 0.0284f
C24374 VGND.n3512 0 0.0934f
C24375 VGND.n3513 0 0.0217f
C24376 VGND.n3514 0 0.0119f
C24377 VGND.t36 0 0.0792f
C24378 VGND.n3515 0 0.0547f
C24379 VGND.n3516 0 0.035f
C24380 VGND.n3517 0 0.0342f
C24381 VGND.n3518 0 0.0511f
C24382 VGND.n3519 0 0.0331f
C24383 VGND.n3520 0 0.00488f
C24384 VGND.n3521 0 0.055f
C24385 VGND.t305 0 0.0409f
C24386 VGND.n3522 0 0.0465f
C24387 VGND.t369 0 0.0445f
C24388 VGND.t339 0 0.0445f
C24389 VGND.n3523 0 0.0222f
C24390 VGND.n3524 0 0.244f
C24391 VGND.n3525 0 0.0163f
C24392 VGND.n3526 0 0.00981f
C24393 VGND.n3527 0 0.015f
C24394 VGND.n3528 0 0.0285f
C24395 VGND.n3529 0 0.0358f
C24396 VGND.n3530 0 0.00981f
C24397 VGND.n3531 0 0.0166f
C24398 VGND.n3532 0 0.0149f
C24399 VGND.n3533 0 0.00837f
C24400 VGND.n3534 0 0.0503f
C24401 VGND.n3535 0 0.037f
C24402 VGND.n3536 0 0.00981f
C24403 VGND.t378 0 0.0792f
C24404 VGND.n3537 0 0.0547f
C24405 VGND.n3538 0 0.0243f
C24406 VGND.n3539 0 0.0166f
C24407 VGND.n3540 0 0.0166f
C24408 VGND.n3541 0 0.015f
C24409 VGND.n3542 0 0.0379f
C24410 VGND.n3543 0 0.00549f
C24411 VGND.n3544 0 0.0356f
C24412 VGND.n3545 0 0.0166f
C24413 VGND.n3546 0 0.0183f
C24414 VGND.n3547 0 0.0166f
C24415 VGND.n3548 0 0.015f
C24416 VGND.n3549 0 0.0261f
C24417 VGND.n3550 0 0.028f
C24418 VGND.n3551 0 0.00981f
C24419 VGND.t66 0 0.0792f
C24420 VGND.n3552 0 0.0547f
C24421 VGND.n3553 0 0.0243f
C24422 VGND.n3554 0 0.0166f
C24423 VGND.n3555 0 0.0166f
C24424 VGND.n3556 0 0.015f
C24425 VGND.n3557 0 0.045f
C24426 VGND.n3558 0 0.00463f
C24427 VGND.n3559 0 0.0166f
C24428 VGND.n3560 0 0.0203f
C24429 VGND.n3561 0 0.0166f
C24430 VGND.n3562 0 0.015f
C24431 VGND.n3563 0 0.0317f
C24432 VGND.n3564 0 0.0415f
C24433 VGND.n3565 0 0.00981f
C24434 VGND.n3566 0 0.0166f
C24435 VGND.n3567 0 0.015f
C24436 VGND.n3568 0 0.0652f
C24437 VGND.n3569 0 0.0157f
C24438 VGND.n3570 0 0.00756f
C24439 VGND.n3571 0 0.009f
C24440 VGND.n3572 0 0.0316f
C24441 VGND.n3573 0 0.094f
C24442 VGND.n3574 0 0.184f
C24443 VGND.n3575 0 0.229f
C24444 VGND.n3576 0 0.0739f
C24445 VGND.n3577 0 0.0192f
C24446 VGND.n3578 0 0.00765f
C24447 VGND.t387 0 0.0799f
C24448 VGND.n3579 0 0.0723f
C24449 VGND.n3580 0 0.0241f
C24450 VGND.n3581 0 0.0104f
C24451 VGND.n3582 0 0.0331f
C24452 VGND.n3583 0 0.0166f
C24453 VGND.n3584 0 0.0537f
C24454 VGND.n3585 0 0.0166f
C24455 VGND.n3586 0 0.0352f
C24456 VGND.n3587 0 0.0166f
C24457 VGND.n3588 0 0.00427f
C24458 VGND.n3589 0 0.015f
C24459 VGND.n3590 0 0.00828f
C24460 VGND.n3591 0 0.00981f
C24461 VGND.n3592 0 0.015f
C24462 VGND.n3593 0 0.00828f
C24463 VGND.n3594 0 0.0563f
C24464 VGND.n3595 0 0.0192f
C24465 VGND.n3596 0 0.00765f
C24466 VGND.n3597 0 0.00891f
C24467 VGND.n3598 0 0.0241f
C24468 VGND.n3599 0 0.0337f
C24469 VGND.n3600 0 0.0553f
C24470 VGND.n3601 0 0.00586f
C24471 VGND.n3602 0 0.00972f
C24472 VGND.n3603 0 0.0432f
C24473 VGND.n3604 0 0.0166f
C24474 VGND.n3605 0 0.0114f
C24475 VGND.n3606 0 0.0166f
C24476 VGND.n3607 0 0.00586f
C24477 VGND.n3608 0 0.0166f
C24478 VGND.n3609 0 0.00586f
C24479 VGND.n3610 0 0.0166f
C24480 VGND.n3611 0 0.00644f
C24481 VGND.n3612 0 0.0166f
C24482 VGND.n3613 0 0.0433f
C24483 VGND.n3614 0 0.0166f
C24484 VGND.n3615 0 0.0132f
C24485 VGND.n3616 0 0.0166f
C24486 VGND.n3617 0 0.015f
C24487 VGND.n3618 0 0.0256f
C24488 VGND.n3619 0 0.0291f
C24489 VGND.n3620 0 0.00981f
C24490 VGND.t65 0 0.0792f
C24491 VGND.n3621 0 0.0547f
C24492 VGND.n3622 0 0.0243f
C24493 VGND.n3623 0 0.0166f
C24494 VGND.n3624 0 0.0148f
C24495 VGND.n3625 0 0.00783f
C24496 VGND.n3626 0 0.00207f
C24497 VGND.n3627 0 0.00315f
C24498 VGND.n3628 0 0.00162f
C24499 VGND.n3629 0 0.00162f
C24500 VGND.n3630 0 0.00189f
C24501 VGND.n3631 0 9.9e-19
C24502 VGND.n3632 0 0.00162f
C24503 VGND.n3633 0 0.00171f
C24504 VGND.n3634 0 0.0573f
C24505 VGND.n3635 0 9.9e-19
C24506 VGND.n3636 0 0.00189f
C24507 VGND.n3637 0 0.00162f
C24508 VGND.n3638 0 0.00342f
C24509 VGND.n3639 0 0.00387f
C24510 VGND.n3640 0 7.2e-19
C24511 VGND.n3641 0 0.00162f
C24512 VGND.n3642 0 0.00207f
C24513 VGND.n3643 0 0.00207f
C24514 VGND.n3644 0 0.00162f
C24515 VGND.n3645 0 0.00234f
C24516 VGND.n3646 0 0.00234f
C24517 VGND.n3647 0 0.00234f
C24518 VGND.n3648 0 0.00297f
C24519 VGND.n3649 0 0.00842f
C24520 VGND.n3650 0 0.00144f
C24521 VGND.n3651 0 0.00135f
C24522 VGND.n3652 0 2.7e-19
C24523 VGND.n3653 0 0.003f
C24524 VGND.n3654 0 0.0179f
C24525 VGND.n3655 0 0.00126f
C24526 VGND.n3656 0 0.00207f
C24527 VGND.n3657 0 0.00126f
C24528 VGND.n3658 0 0.00126f
C24529 VGND.n3659 0 0.00701f
C24530 VGND.n3660 0 0.0041f
C24531 VGND.n3661 0 0.018f
C24532 VGND.n3662 0 0.00287f
C24533 VGND.n3663 0 0.00207f
C24534 VGND.n3664 0 0.00274f
C24535 VGND.n3665 0 0.00403f
C24536 VGND.n3666 0 0.00493f
C24537 VGND.n3667 0 0.00126f
C24538 VGND.n3668 0 0.00173f
C24539 VGND.n3670 0 0.192f
C24540 VGND.n3671 0 0.134f
C24541 VGND.n3672 0 0.308f
C24542 VGND.n3673 0 4.5f
C24543 VGND.n3674 0 3.67f
C24544 VGND.n3675 0 0.134f
C24545 VGND.n3676 0 0.00207f
C24546 VGND.n3677 0 0.00287f
C24547 VGND.n3678 0 0.00173f
C24548 VGND.n3679 0 0.00269f
C24549 VGND.n3680 0 0.0039f
C24550 VGND.n3681 0 0.00269f
C24551 VGND.n3682 0 0.00173f
C24552 VGND.n3684 0 0.317f
C24553 VGND.n3685 0 0.317f
C24554 VGND.n3686 0 0.00287f
C24555 VGND.n3687 0 0.00207f
C24556 VGND.n3688 0 0.00274f
C24557 VGND.n3689 0 0.00403f
C24558 VGND.n3690 0 0.00493f
C24559 VGND.n3691 0 0.00126f
C24560 VGND.n3692 0 0.00173f
C24561 VGND.n3694 0 0.018f
C24562 VGND.n3695 0 0.00274f
C24563 VGND.n3696 0 0.00173f
C24564 VGND.n3697 0 0.0041f
C24565 VGND.n3698 0 0.00701f
C24566 VGND.n3699 0 0.00252f
C24567 VGND.n3700 0 0.00369f
C24568 VGND.n3701 0 0.00189f
C24569 VGND.n3702 0 0.00135f
C24570 VGND.n3703 0 0.00207f
C24571 VGND.n3704 0 0.00126f
C24572 VGND.n3705 0 0.00126f
C24573 VGND.n3706 0 0.00207f
C24574 VGND.n3707 0 0.00126f
C24575 VGND.n3708 0 1.12e-19
C24576 VGND.n3709 0 0.00151f
C24577 VGND.n3710 0 0.00144f
C24578 VGND.n3711 0 0.00297f
C24579 VGND.n3712 0 0.00234f
C24580 VGND.n3713 0 0.00234f
C24581 VGND.n3714 0 0.00234f
C24582 VGND.n3715 0 0.00234f
C24583 VGND.n3716 0 0.00162f
C24584 VGND.n3717 0 0.00207f
C24585 VGND.n3718 0 0.00207f
C24586 VGND.n3719 0 0.00387f
C24587 VGND.n3720 0 0.00342f
C24588 VGND.n3721 0 0.00162f
C24589 VGND.n3722 0 0.00189f
C24590 VGND.n3723 0 9.9e-19
C24591 VGND.n3724 0 0.00459f
C24592 VGND.n3725 0 0.0331f
C24593 VGND.n3726 0 0.0554f
C24594 VGND.n3727 0 0.0331f
C24595 VGND.n3728 0 0.00837f
C24596 VGND.t110 0 0.119f
C24597 VGND.n3729 0 0.053f
C24598 VGND.n3730 0 0.0446f
C24599 VGND.n3731 0 0.0433f
C24600 VGND.n3732 0 0.0374f
C24601 VGND.n3733 0 0.0162f
C24602 VGND.n3734 0 0.00972f
C24603 VGND.n3735 0 0.0166f
C24604 VGND.n3736 0 0.0324f
C24605 VGND.n3737 0 0.0166f
C24606 VGND.n3738 0 0.0331f
C24607 VGND.n3739 0 0.0166f
C24608 VGND.n3740 0 0.0379f
C24609 VGND.n3741 0 0.0144f
C24610 VGND.n3742 0 0.00891f
C24611 VGND.n3743 0 0.00549f
C24612 VGND.n3744 0 0.042f
C24613 VGND.n3745 0 0.00981f
C24614 VGND.n3746 0 0.0298f
C24615 VGND.n3747 0 0.0166f
C24616 VGND.n3748 0 0.015f
C24617 VGND.n3749 0 0.00549f
C24618 VGND.n3750 0 0.0435f
C24619 VGND.n3751 0 0.00981f
C24620 VGND.t366 0 0.0792f
C24621 VGND.n3752 0 0.0658f
C24622 VGND.n3753 0 0.0243f
C24623 VGND.n3754 0 0.0166f
C24624 VGND.n3755 0 0.0166f
C24625 VGND.n3756 0 0.0151f
C24626 VGND.n3757 0 0.0379f
C24627 VGND.n3758 0 0.00488f
C24628 VGND.n3759 0 0.00972f
C24629 VGND.n3760 0 0.043f
C24630 VGND.n3761 0 0.0166f
C24631 VGND.n3762 0 0.00756f
C24632 VGND.n3763 0 0.0166f
C24633 VGND.n3764 0 0.026f
C24634 VGND.n3765 0 0.0166f
C24635 VGND.n3766 0 0.00586f
C24636 VGND.n3767 0 0.0166f
C24637 VGND.n3768 0 0.00586f
C24638 VGND.n3769 0 0.0166f
C24639 VGND.n3770 0 0.00787f
C24640 VGND.n3771 0 0.0166f
C24641 VGND.n3772 0 0.015f
C24642 VGND.n3773 0 0.0497f
C24643 VGND.n3774 0 0.0386f
C24644 VGND.n3775 0 0.00981f
C24645 VGND.t27 0 0.0792f
C24646 VGND.n3776 0 0.0547f
C24647 VGND.n3777 0 0.0243f
C24648 VGND.n3778 0 0.0166f
C24649 VGND.n3779 0 0.0166f
C24650 VGND.n3780 0 0.0144f
C24651 VGND.n3781 0 0.00171f
C24652 VGND.n3782 0 0.00171f
C24653 VGND.n3783 0 0.00162f
C24654 VGND.n3784 0 9.9e-19
C24655 VGND.n3785 0 0.00189f
C24656 VGND.n3786 0 0.00162f
C24657 VGND.n3787 0 0.00162f
C24658 VGND.n3788 0 0.00315f
C24659 VGND.n3789 0 0.00207f
C24660 VGND.n3790 0 7.2e-19
C24661 VGND.n3791 0 7.2e-19
C24662 VGND.n3792 0 0.00162f
C24663 VGND.n3793 0 7.2e-19
C24664 VGND.n3794 0 0.00153f
C24665 VGND.n3795 0 1.46e-19
C24666 VGND.n3796 0 0.00185f
C24667 VGND.n3797 0 9.77e-19
C24668 VGND.n3798 0 0.0301f
C24669 VGND.n3799 0 0.049f
C24670 VGND.n3800 0 0.139f
C24671 VGND.n3801 0 0.0697f
C24672 VGND.n3802 0 0.009f
C24673 VGND.n3803 0 0.0111f
C24674 VGND.n3804 0 0.045f
C24675 VGND.n3805 0 0.0631f
C24676 VGND.n3806 0 0.015f
C24677 VGND.n3807 0 0.035f
C24678 VGND.n3808 0 0.0166f
C24679 VGND.n3809 0 0.0166f
C24680 VGND.n3810 0 0.0166f
C24681 VGND.n3811 0 0.0361f
C24682 VGND.n3812 0 0.0345f
C24683 VGND.n3813 0 0.0271f
C24684 VGND.t134 0 0.0946f
C24685 VGND.n3814 0 0.0183f
C24686 VGND.n3815 0 0.0961f
C24687 VGND.n3816 0 0.0318f
C24688 VGND.n3817 0 0.0378f
C24689 VGND.n3818 0 0.00981f
C24690 VGND.n3819 0 0.00828f
C24691 VGND.n3820 0 0.0448f
C24692 VGND.n3821 0 0.0436f
C24693 VGND.n3822 0 0.0144f
C24694 VGND.n3823 0 0.0525f
C24695 VGND.n3824 0 0.0166f
C24696 VGND.n3825 0 0.0324f
C24697 VGND.n3826 0 0.0166f
C24698 VGND.n3827 0 0.0316f
C24699 VGND.n3828 0 0.0166f
C24700 VGND.n3829 0 0.0166f
C24701 VGND.n3830 0 0.0166f
C24702 VGND.n3831 0 0.0252f
C24703 VGND.n3832 0 0.0391f
C24704 VGND.n3833 0 0.0491f
C24705 VGND.t301 0 0.0946f
C24706 VGND.n3834 0 0.0183f
C24707 VGND.n3835 0 0.0961f
C24708 VGND.n3836 0 0.0252f
C24709 VGND.n3837 0 0.0271f
C24710 VGND.n3838 0 0.00972f
C24711 VGND.n3839 0 0.00837f
C24712 VGND.n3840 0 0.0448f
C24713 VGND.n3841 0 0.0694f
C24714 VGND.n3842 0 0.0144f
C24715 VGND.n3843 0 0.0331f
C24716 VGND.n3844 0 0.0166f
C24717 VGND.n3845 0 0.0166f
C24718 VGND.n3846 0 0.0221f
C24719 VGND.n3847 0 0.0481f
C24720 VGND.n3848 0 0.03f
C24721 VGND.n3849 0 0.0469f
C24722 VGND.n3850 0 0.0372f
C24723 VGND.n3851 0 0.0119f
C24724 VGND.n3852 0 0.0551f
C24725 VGND.n3853 0 0.058f
C24726 VGND.n3854 0 0.0269f
C24727 VGND.n3855 0 0.0166f
C24728 VGND.n3856 0 0.0145f
C24729 VGND.n3857 0 0.00824f
C24730 VGND.n3858 0 0.00234f
C24731 VGND.n3859 0 0.00297f
C24732 VGND.n3860 0 0.00315f
C24733 VGND.n3861 0 0.00207f
C24734 VGND.n3862 0 9.9e-19
C24735 VGND.n3863 0 0.00261f
C24736 VGND.n3864 0 0.00207f
C24737 VGND.n3865 0 0.00135f
C24738 VGND.n3866 0 7.2e-19
C24739 VGND.n3867 0 0.00126f
C24740 VGND.n3868 0 0.00135f
C24741 VGND.n3869 0 0.00126f
C24742 VGND.n3870 0 0.0254f
C24743 VGND.n3871 0 0.00198f
C24744 VGND.n3872 0 0.00453f
C24745 VGND.n3873 0 0.00153f
C24746 VGND.n3874 0 0.00282f
C24747 VGND.n3875 0 0.00144f
C24748 VGND.n3876 0 0.00651f
C24749 VGND.n3877 0 0.00261f
C24750 VGND.n3878 0 0.00234f
C24751 VGND.n3879 0 0.00234f
C24752 VGND.n3880 0 0.00225f
C24753 VGND.n3881 0 0.00144f
C24754 VGND.n3882 0 0.00148f
C24755 VGND.n3883 0 8.57e-19
C24756 VGND.n3884 0 0.0246f
C24757 VGND.n3885 0 0.202f
C24758 VGND.n3886 0 0.094f
C24759 VGND.t133 0 0.128f
C24760 VGND.n3887 0 0.154f
C24761 VGND.n3888 0 0.0441f
C24762 VGND.n3889 0 0.057f
C24763 VGND.n3890 0 0.0375f
C24764 VGND.n3891 0 0.0383f
C24765 VGND.n3892 0 0.0323f
C24766 VGND.n3893 0 0.0331f
C24767 VGND.n3894 0 0.00981f
C24768 VGND.t122 0 0.0792f
C24769 VGND.n3895 0 0.046f
C24770 VGND.t342 0 0.0837f
C24771 VGND.t169 0 0.0837f
C24772 VGND.n3896 0 0.324f
C24773 VGND.t318 0 0.0445f
C24774 VGND.t287 0 0.0445f
C24775 VGND.n3897 0 0.243f
C24776 VGND.n3898 0 0.0173f
C24777 VGND.n3899 0 0.0222f
C24778 VGND.n3900 0 0.00891f
C24779 VGND.n3901 0 0.0253f
C24780 VGND.n3902 0 0.00351f
C24781 VGND.n3903 0 0.00981f
C24782 VGND.n3904 0 0.015f
C24783 VGND.n3905 0 0.0045f
C24784 VGND.n3906 0 0.0435f
C24785 VGND.n3907 0 0.0658f
C24786 VGND.n3908 0 0.0243f
C24787 VGND.n3909 0 0.0166f
C24788 VGND.n3910 0 0.0166f
C24789 VGND.n3911 0 0.0151f
C24790 VGND.n3912 0 0.0373f
C24791 VGND.n3913 0 0.00233f
C24792 VGND.n3914 0 0.00972f
C24793 VGND.n3915 0 0.0166f
C24794 VGND.n3916 0 0.00753f
C24795 VGND.n3917 0 0.0166f
C24796 VGND.n3918 0 0.0441f
C24797 VGND.n3919 0 0.0166f
C24798 VGND.n3920 0 0.0303f
C24799 VGND.n3921 0 0.0166f
C24800 VGND.n3922 0 0.00564f
C24801 VGND.n3923 0 0.0166f
C24802 VGND.n3924 0 0.0107f
C24803 VGND.n3925 0 0.0166f
C24804 VGND.n3926 0 0.015f
C24805 VGND.n3927 0 0.019f
C24806 VGND.n3928 0 0.0275f
C24807 VGND.n3929 0 0.015f
C24808 VGND.n3930 0 0.00756f
C24809 VGND.n3931 0 0.0157f
C24810 VGND.t59 0 0.0818f
C24811 VGND.n3932 0 0.139f
C24812 VGND.n3933 0 0.0316f
C24813 VGND.n3934 0 0.009f
C24814 VGND.n3935 0 0.0112f
C24815 VGND.n3936 0 0.00891f
C24816 VGND.n3937 0 0.00837f
C24817 VGND.n3938 0 0.0385f
C24818 VGND.n3939 0 0.0224f
C24819 VGND.n3940 0 0.00972f
C24820 VGND.n3941 0 0.0166f
C24821 VGND.n3942 0 0.00488f
C24822 VGND.n3943 0 0.0166f
C24823 VGND.n3944 0 0.0245f
C24824 VGND.n3945 0 0.0166f
C24825 VGND.n3946 0 0.015f
C24826 VGND.n3947 0 0.0059f
C24827 VGND.n3948 0 0.0291f
C24828 VGND.n3949 0 0.00981f
C24829 VGND.t58 0 0.0792f
C24830 VGND.n3950 0 0.0547f
C24831 VGND.n3951 0 0.0601f
C24832 VGND.n3952 0 0.0166f
C24833 VGND.n3953 0 0.0166f
C24834 VGND.n3954 0 0.015f
C24835 VGND.n3955 0 0.0375f
C24836 VGND.n3956 0 0.0448f
C24837 VGND.n3957 0 0.00972f
C24838 VGND.n3958 0 0.0321f
C24839 VGND.n3959 0 0.0525f
C24840 VGND.n3960 0 0.0166f
C24841 VGND.t109 0 0.0946f
C24842 VGND.n3961 0 0.0183f
C24843 VGND.n3962 0 0.0961f
C24844 VGND.n3963 0 0.0275f
C24845 VGND.n3964 0 0.0271f
C24846 VGND.n3965 0 0.0166f
C24847 VGND.n3966 0 0.0345f
C24848 VGND.n3967 0 0.0474f
C24849 VGND.n3968 0 0.0166f
C24850 VGND.n3969 0 0.033f
C24851 VGND.n3970 0 0.0166f
C24852 VGND.n3971 0 0.0324f
C24853 VGND.n3972 0 0.0166f
C24854 VGND.n3973 0 0.0166f
C24855 VGND.n3974 0 0.0142f
C24856 VGND.n3975 0 0.012f
C24857 VGND.n3976 0 0.0271f
C24858 VGND.n3977 0 0.00972f
C24859 VGND.n3978 0 0.0446f
C24860 VGND.n3979 0 0.0166f
C24861 VGND.n3980 0 0.0312f
C24862 VGND.n3981 0 0.0136f
C24863 VGND.n3982 0 0.0063f
C24864 VGND.n3983 0 0.00824f
C24865 VGND.n3984 0 0.00413f
C24866 VGND.n3985 0 0.018f
C24867 VGND.n3986 0 0.00269f
C24868 VGND.n3987 0 0.00207f
C24869 VGND.n3988 0 0.00287f
C24870 VGND.n3989 0 0.00173f
C24871 VGND.n3991 0 0.317f
C24872 VGND.n3992 0 0.317f
C24873 VGND.n3993 0 0.00207f
C24874 VGND.n3994 0 0.00287f
C24875 VGND.n3995 0 0.0039f
C24876 VGND.n3996 0 0.00269f
C24877 VGND.n3997 0 0.00173f
C24878 VGND.n3999 0 0.018f
C24879 VGND.n4000 0 0.00274f
C24880 VGND.n4001 0 0.00173f
C24881 VGND.n4002 0 0.00413f
C24882 VGND.n4003 0 0.00824f
C24883 VGND.n4004 0 0.0063f
C24884 VGND.t92 0 0.082f
C24885 VGND.n4005 0 0.0934f
C24886 VGND.n4006 0 0.0261f
C24887 VGND.n4007 0 0.0191f
C24888 VGND.n4008 0 0.0137f
C24889 VGND.n4009 0 0.045f
C24890 VGND.t275 0 0.157f
C24891 VGND.n4010 0 0.199f
C24892 VGND.n4011 0 0.033f
C24893 VGND.n4012 0 0.0291f
C24894 VGND.n4013 0 0.0875f
C24895 VGND.n4014 0 0.015f
C24896 VGND.n4015 0 0.0166f
C24897 VGND.n4016 0 0.0352f
C24898 VGND.n4017 0 0.0172f
C24899 VGND.n4018 0 0.00828f
C24900 VGND.n4019 0 0.0372f
C24901 VGND.n4020 0 0.00389f
C24902 VGND.n4021 0 0.015f
C24903 VGND.n4022 0 0.00981f
C24904 VGND.n4023 0 0.0081f
C24905 VGND.n4024 0 0.0194f
C24906 VGND.n4025 0 0.0247f
C24907 VGND.n4026 0 0.00909f
C24908 VGND.n4027 0 0.0112f
C24909 VGND.n4028 0 0.045f
C24910 VGND.t151 0 0.128f
C24911 VGND.n4029 0 0.154f
C24912 VGND.n4030 0 0.058f
C24913 VGND.n4031 0 0.00828f
C24914 VGND.n4032 0 0.0172f
C24915 VGND.n4033 0 0.015f
C24916 VGND.n4034 0 0.0104f
C24917 VGND.n4035 0 0.00414f
C24918 VGND.n4036 0 0.0384f
C24919 VGND.n4037 0 0.00765f
C24920 VGND.n4038 0 0.0172f
C24921 VGND.n4039 0 0.0166f
C24922 VGND.t274 0 0.0792f
C24923 VGND.n4040 0 0.0394f
C24924 VGND.n4041 0 0.0166f
C24925 VGND.n4042 0 0.0331f
C24926 VGND.n4043 0 0.00981f
C24927 VGND.t324 0 0.0792f
C24928 VGND.n4044 0 0.0287f
C24929 VGND.n4045 0 0.0387f
C24930 VGND.n4046 0 0.00981f
C24931 VGND.t230 0 0.0792f
C24932 VGND.n4047 0 0.0265f
C24933 VGND.n4048 0 0.0329f
C24934 VGND.t262 0 0.0445f
C24935 VGND.t146 0 0.0445f
C24936 VGND.n4049 0 0.243f
C24937 VGND.t383 0 0.0837f
C24938 VGND.n4050 0 0.0173f
C24939 VGND.n4051 0 0.0247f
C24940 VGND.n4052 0 0.186f
C24941 VGND.t187 0 0.126f
C24942 VGND.n4053 0 0.178f
C24943 VGND.n4054 0 0.0453f
C24944 VGND.n4055 0 0.0378f
C24945 VGND.n4056 0 0.015f
C24946 VGND.n4057 0 0.00828f
C24947 VGND.n4058 0 0.025f
C24948 VGND.n4059 0 0.0278f
C24949 VGND.n4060 0 0.0547f
C24950 VGND.n4061 0 0.0442f
C24951 VGND.n4062 0 0.0166f
C24952 VGND.n4063 0 0.0166f
C24953 VGND.n4064 0 0.0152f
C24954 VGND.n4065 0 0.0373f
C24955 VGND.n4066 0 0.00236f
C24956 VGND.n4067 0 0.00963f
C24957 VGND.n4068 0 0.0166f
C24958 VGND.n4069 0 0.015f
C24959 VGND.n4070 0 0.00444f
C24960 VGND.n4071 0 0.0291f
C24961 VGND.n4072 0 0.074f
C24962 VGND.n4073 0 0.0284f
C24963 VGND.n4074 0 0.0166f
C24964 VGND.n4075 0 0.0166f
C24965 VGND.n4076 0 0.0166f
C24966 VGND.n4077 0 0.0373f
C24967 VGND.n4078 0 0.0325f
C24968 VGND.n4079 0 0.0239f
C24969 VGND.n4080 0 0.015f
C24970 VGND.n4081 0 0.00828f
C24971 VGND.n4082 0 0.00981f
C24972 VGND.n4083 0 0.0283f
C24973 VGND.n4084 0 0.0547f
C24974 VGND.n4085 0 0.0243f
C24975 VGND.n4086 0 0.0499f
C24976 VGND.n4087 0 0.0166f
C24977 VGND.n4088 0 0.0143f
C24978 VGND.n4089 0 0.00828f
C24979 VGND.n4090 0 0.03f
C24980 VGND.n4091 0 0.049f
C24981 VGND.n4092 0 0.229f
C24982 VGND.n4093 0 0.094f
C24983 VGND.t84 0 0.0818f
C24984 VGND.n4094 0 0.139f
C24985 VGND.n4095 0 0.0316f
C24986 VGND.n4096 0 0.009f
C24987 VGND.n4097 0 0.0112f
C24988 VGND.n4098 0 0.00891f
C24989 VGND.n4099 0 0.028f
C24990 VGND.n4100 0 0.0384f
C24991 VGND.n4101 0 0.00981f
C24992 VGND.n4102 0 0.0401f
C24993 VGND.n4103 0 0.0166f
C24994 VGND.n4104 0 0.00707f
C24995 VGND.n4105 0 0.0166f
C24996 VGND.n4106 0 0.015f
C24997 VGND.n4107 0 0.011f
C24998 VGND.n4108 0 0.0291f
C24999 VGND.n4109 0 0.00981f
C25000 VGND.t199 0 0.0792f
C25001 VGND.n4110 0 0.0547f
C25002 VGND.n4111 0 0.0243f
C25003 VGND.n4112 0 0.0166f
C25004 VGND.n4113 0 0.0166f
C25005 VGND.n4114 0 0.0151f
C25006 VGND.n4115 0 0.0379f
C25007 VGND.n4116 0 0.0151f
C25008 VGND.n4117 0 0.00972f
C25009 VGND.n4118 0 0.0492f
C25010 VGND.n4119 0 0.0166f
C25011 VGND.n4120 0 0.0112f
C25012 VGND.n4121 0 0.0166f
C25013 VGND.n4122 0 0.00586f
C25014 VGND.n4123 0 0.0166f
C25015 VGND.n4124 0 0.00586f
C25016 VGND.n4125 0 0.0166f
C25017 VGND.n4126 0 0.0285f
C25018 VGND.n4127 0 0.0166f
C25019 VGND.n4128 0 0.00697f
C25020 VGND.n4129 0 0.0166f
C25021 VGND.n4130 0 0.015f
C25022 VGND.n4131 0 0.0386f
C25023 VGND.n4132 0 0.028f
C25024 VGND.n4133 0 0.00981f
C25025 VGND.n4134 0 0.0166f
C25026 VGND.n4135 0 0.015f
C25027 VGND.n4136 0 0.00828f
C25028 VGND.n4137 0 0.0192f
C25029 VGND.t153 0 0.0799f
C25030 VGND.n4138 0 0.0723f
C25031 VGND.n4139 0 0.0241f
C25032 VGND.n4140 0 0.0148f
C25033 VGND.n4141 0 0.00783f
C25034 VGND.n4142 0 0.00207f
C25035 VGND.n4143 0 0.00315f
C25036 VGND.n4144 0 0.00162f
C25037 VGND.n4145 0 0.00162f
C25038 VGND.n4146 0 0.00189f
C25039 VGND.n4147 0 9.9e-19
C25040 VGND.n4148 0 0.00162f
C25041 VGND.n4149 0 0.00171f
C25042 VGND.n4150 0 0.0377f
C25043 VGND.n4151 0 9.9e-19
C25044 VGND.n4152 0 0.00189f
C25045 VGND.n4153 0 0.00162f
C25046 VGND.n4154 0 0.00342f
C25047 VGND.n4155 0 0.00387f
C25048 VGND.n4156 0 7.2e-19
C25049 VGND.n4157 0 0.00162f
C25050 VGND.n4158 0 0.00207f
C25051 VGND.n4159 0 0.00207f
C25052 VGND.n4160 0 0.00162f
C25053 VGND.n4161 0 0.00234f
C25054 VGND.n4162 0 0.00234f
C25055 VGND.n4163 0 0.00234f
C25056 VGND.n4164 0 0.00297f
C25057 VGND.n4165 0 0.00144f
C25058 VGND.n4166 0 0.00151f
C25059 VGND.n4167 0 1.12e-19
C25060 VGND.n4168 0 0.00126f
C25061 VGND.n4169 0 0.00207f
C25062 VGND.n4170 0 0.00126f
C25063 VGND.n4171 0 0.00126f
C25064 VGND.n4172 0 0.00701f
C25065 VGND.n4173 0 0.0041f
C25066 VGND.n4174 0 0.018f
C25067 VGND.n4175 0 0.00287f
C25068 VGND.n4176 0 0.00207f
C25069 VGND.n4177 0 0.00274f
C25070 VGND.n4178 0 0.00403f
C25071 VGND.n4179 0 0.00493f
C25072 VGND.n4180 0 0.00126f
C25073 VGND.n4181 0 0.00173f
C25074 VGND.n4183 0 0.317f
C25075 VGND.n4184 0 0.317f
C25076 VGND.n4185 0 0.00207f
C25077 VGND.n4186 0 0.00287f
C25078 VGND.n4187 0 0.00173f
C25079 VGND.n4188 0 0.00269f
C25080 VGND.n4189 0 0.0039f
C25081 VGND.n4190 0 0.00269f
C25082 VGND.n4191 0 0.00173f
C25083 VGND.n4193 0 0.00162f
C25084 VGND.n4194 0 9.9e-19
C25085 VGND.n4195 0 0.00189f
C25086 VGND.n4196 0 0.00162f
C25087 VGND.n4197 0 0.00162f
C25088 VGND.n4198 0 0.00315f
C25089 VGND.n4199 0 0.00207f
C25090 VGND.n4200 0 7.2e-19
C25091 VGND.n4201 0 7.2e-19
C25092 VGND.n4202 0 0.00162f
C25093 VGND.n4203 0 0.00207f
C25094 VGND.n4204 0 0.00207f
C25095 VGND.n4205 0 0.00162f
C25096 VGND.n4206 0 0.00234f
C25097 VGND.t186 0 0.0837f
C25098 VGND.t313 0 0.0837f
C25099 VGND.n4207 0 0.324f
C25100 VGND.n4208 0 0.0107f
C25101 VGND.t157 0 0.0813f
C25102 VGND.n4209 0 0.139f
C25103 VGND.n4210 0 0.0496f
C25104 VGND.t273 0 0.225f
C25105 VGND.n4211 0 0.336f
C25106 VGND.n4212 0 0.0586f
C25107 VGND.n4213 0 0.0336f
C25108 VGND.n4214 0 0.0526f
C25109 VGND.t206 0 0.082f
C25110 VGND.n4215 0 0.139f
C25111 VGND.t127 0 0.148f
C25112 VGND.n4216 0 0.0882f
C25113 VGND.t258 0 0.121f
C25114 VGND.n4217 0 0.059f
C25115 VGND.n4218 0 0.123f
C25116 VGND.n4219 0 0.0603f
C25117 VGND.n4220 0 0.0271f
C25118 VGND.n4221 0 0.00828f
C25119 VGND.t156 0 0.0812f
C25120 VGND.n4222 0 0.139f
C25121 VGND.t103 0 0.0837f
C25122 VGND.t88 0 0.0445f
C25123 VGND.t73 0 0.0445f
C25124 VGND.n4223 0 0.243f
C25125 VGND.n4224 0 0.032f
C25126 VGND.n4225 0 0.0351f
C25127 VGND.t215 0 0.0837f
C25128 VGND.n4226 0 0.324f
C25129 VGND.n4227 0 0.0243f
C25130 VGND.n4228 0 0.015f
C25131 VGND.n4229 0 0.0265f
C25132 VGND.n4230 0 0.0166f
C25133 VGND.n4231 0 0.00963f
C25134 VGND.n4232 0 0.00476f
C25135 VGND.n4233 0 0.0107f
C25136 VGND.n4234 0 0.0172f
C25137 VGND.n4235 0 0.0349f
C25138 VGND.t242 0 0.0813f
C25139 VGND.n4236 0 0.139f
C25140 VGND.n4237 0 0.0363f
C25141 VGND.n4238 0 0.0245f
C25142 VGND.n4239 0 0.015f
C25143 VGND.n4240 0 0.032f
C25144 VGND.n4241 0 0.00981f
C25145 VGND.n4242 0 0.015f
C25146 VGND.n4243 0 0.00457f
C25147 VGND.n4244 0 0.0697f
C25148 VGND.n4245 0 0.0142f
C25149 VGND.n4246 0 0.0604f
C25150 VGND.n4247 0 0.0166f
C25151 VGND.n4248 0 0.059f
C25152 VGND.n4249 0 0.0166f
C25153 VGND.n4250 0 0.0166f
C25154 VGND.n4251 0 0.0166f
C25155 VGND.n4252 0 0.009f
C25156 VGND.n4253 0 0.00981f
C25157 VGND.n4254 0 0.0327f
C25158 VGND.n4255 0 0.0245f
C25159 VGND.n4256 0 0.0584f
C25160 VGND.n4257 0 0.014f
C25161 VGND.n4258 0 0.00756f
C25162 VGND.n4259 0 0.009f
C25163 VGND.n4260 0 0.0111f
C25164 VGND.n4261 0 0.0447f
C25165 VGND.n4262 0 0.0801f
C25166 VGND.n4263 0 0.015f
C25167 VGND.n4264 0 0.0166f
C25168 VGND.n4265 0 0.0166f
C25169 VGND.n4266 0 0.039f
C25170 VGND.n4267 0 0.0393f
C25171 VGND.n4268 0 0.0449f
C25172 VGND.n4269 0 0.0315f
C25173 VGND.n4270 0 0.015f
C25174 VGND.n4271 0 0.0535f
C25175 VGND.n4272 0 0.0166f
C25176 VGND.n4273 0 0.0166f
C25177 VGND.n4274 0 0.0166f
C25178 VGND.n4275 0 0.0166f
C25179 VGND.n4276 0 0.0176f
C25180 VGND.n4277 0 0.0385f
C25181 VGND.n4278 0 0.0535f
C25182 VGND.t102 0 0.151f
C25183 VGND.n4279 0 0.126f
C25184 VGND.n4280 0 0.0274f
C25185 VGND.n4281 0 0.0385f
C25186 VGND.n4282 0 0.0426f
C25187 VGND.n4283 0 0.0493f
C25188 VGND.n4284 0 0.0475f
C25189 VGND.n4285 0 0.0633f
C25190 VGND.n4286 0 0.00981f
C25191 VGND.n4287 0 0.052f
C25192 VGND.n4288 0 0.0172f
C25193 VGND.n4289 0 0.00828f
C25194 VGND.n4290 0 0.0258f
C25195 VGND.n4291 0 0.0265f
C25196 VGND.n4292 0 0.015f
C25197 VGND.n4293 0 0.0243f
C25198 VGND.n4294 0 0.0328f
C25199 VGND.n4295 0 0.0249f
C25200 VGND.n4296 0 0.009f
C25201 VGND.n4297 0 0.00378f
C25202 VGND.n4298 0 0.00126f
C25203 VGND.n4299 0 0.00207f
C25204 VGND.n4300 0 0.0175f
C25205 VGND.n4301 0 0.0195f
C25206 VGND.n4302 0 0.00126f
C25207 VGND.n4303 0 2.7e-19
C25208 VGND.n4304 0 0.00135f
C25209 VGND.n4305 0 0.0177f
C25210 VGND.n4306 0 0.00414f
C25211 VGND.n4307 0 0.00315f
C25212 VGND.n4308 0 0.0281f
C25213 VGND.t299 0 0.0792f
C25214 VGND.n4309 0 0.034f
C25215 VGND.n4310 0 0.0547f
C25216 VGND.n4311 0 0.00386f
C25217 VGND.n4312 0 0.0324f
C25218 VGND.n4313 0 0.0306f
C25219 VGND.n4314 0 0.0248f
C25220 VGND.n4315 0 0.0155f
C25221 VGND.n4316 0 0.0745f
C25222 VGND.t128 0 0.128f
C25223 VGND.n4317 0 0.156f
C25224 VGND.n4318 0 0.0472f
C25225 VGND.n4319 0 0.0371f
C25226 VGND.t347 0 0.0792f
C25227 VGND.n4320 0 0.0243f
C25228 VGND.n4321 0 0.0547f
C25229 VGND.n4322 0 0.00427f
C25230 VGND.n4323 0 0.0325f
C25231 VGND.t5 0 0.0792f
C25232 VGND.n4324 0 0.0243f
C25233 VGND.n4325 0 0.074f
C25234 VGND.n4326 0 0.00586f
C25235 VGND.t29 0 0.0792f
C25236 VGND.n4327 0 0.0428f
C25237 VGND.n4328 0 0.0547f
C25238 VGND.n4329 0 0.00251f
C25239 VGND.n4330 0 0.00287f
C25240 VGND.n4331 0 0.00207f
C25241 VGND.n4332 0 0.00274f
C25242 VGND.n4333 0 0.00173f
C25243 VGND.n4334 0 0.00415f
C25244 VGND.n4335 0 0.00261f
C25245 VGND.n4336 0 0.00207f
C25246 VGND.n4337 0 0.00135f
C25247 VGND.n4338 0 7.2e-19
C25248 VGND.n4339 0 9.9e-19
C25249 VGND.n4340 0 0.00207f
C25250 VGND.n4341 0 0.00315f
C25251 VGND.n4342 0 0.00297f
C25252 VGND.n4343 0 0.00234f
C25253 VGND.n4344 0 0.00823f
C25254 VGND.n4345 0 0.0111f
C25255 VGND.n4346 0 0.00198f
C25256 VGND.n4347 0 0.003f
C25257 VGND.n4348 0 0.00153f
C25258 VGND.n4349 0 0.00282f
C25259 VGND.n4350 0 0.00144f
C25260 VGND.n4351 0 0.0205f
C25261 VGND.n4352 0 0.00261f
C25262 VGND.n4353 0 0.00234f
C25263 VGND.n4354 0 0.00234f
C25264 VGND.n4355 0 0.00315f
C25265 VGND.n4356 0 0.0286f
C25266 VGND.n4357 0 0.00162f
C25267 VGND.n4358 0 0.00135f
C25268 VGND.n4359 0 9.9e-19
C25269 VGND.n4360 0 0.00943f
C25270 VGND.n4361 0 0.0113f
C25271 VGND.n4362 0 0.00126f
C25272 VGND.n4363 0 0.00135f
C25273 VGND.n4364 0 0.00126f
C25274 VGND.n4365 0 0.00414f
C25275 VGND.n4366 0 0.00351f
C25276 VGND.n4367 0 0.00198f
C25277 VGND.n4368 0 0.00126f
C25278 VGND.n4369 0 0.00153f
C25279 VGND.n4370 0 0.00675f
C25280 VGND.n4371 0 0.0147f
C25281 VGND.n4372 0 0.0356f
C25282 VGND.n4373 0 0.00981f
C25283 VGND.n4374 0 0.0166f
C25284 VGND.n4375 0 0.0376f
C25285 VGND.n4376 0 0.0166f
C25286 VGND.n4377 0 0.0379f
C25287 VGND.n4378 0 0.0166f
C25288 VGND.n4379 0 0.0149f
C25289 VGND.n4380 0 0.0166f
C25290 VGND.n4381 0 0.0427f
C25291 VGND.n4382 0 0.0166f
C25292 VGND.n4383 0 0.00586f
C25293 VGND.n4384 0 0.0166f
C25294 VGND.n4385 0 0.015f
C25295 VGND.n4386 0 0.00828f
C25296 VGND.n4387 0 0.00549f
C25297 VGND.n4388 0 0.0332f
C25298 VGND.n4389 0 0.00981f
C25299 VGND.n4390 0 0.0166f
C25300 VGND.n4391 0 0.0331f
C25301 VGND.n4392 0 0.0166f
C25302 VGND.n4393 0 0.0373f
C25303 VGND.n4394 0 0.0166f
C25304 VGND.n4395 0 0.0166f
C25305 VGND.n4396 0 0.015f
C25306 VGND.n4397 0 0.00828f
C25307 VGND.n4398 0 0.0368f
C25308 VGND.n4399 0 0.0509f
C25309 VGND.n4400 0 0.00981f
C25310 VGND.n4401 0 0.0166f
C25311 VGND.n4402 0 0.0506f
C25312 VGND.n4403 0 0.015f
C25313 VGND.n4404 0 0.00828f
C25314 VGND.n4405 0 0.0166f
C25315 VGND.n4406 0 0.026f
C25316 VGND.n4407 0 0.0112f
C25317 VGND.n4408 0 0.045f
C25318 VGND.t314 0 0.082f
C25319 VGND.n4409 0 0.0934f
C25320 VGND.n4410 0 0.028f
C25321 VGND.n4411 0 0.00819f
C25322 VGND.n4412 0 0.00828f
C25323 VGND.n4413 0 0.00828f
C25324 VGND.t95 0 0.148f
C25325 VGND.n4414 0 0.093f
C25326 VGND.t377 0 0.155f
C25327 VGND.n4415 0 0.0449f
C25328 VGND.n4416 0 0.163f
C25329 VGND.n4417 0 0.0147f
C25330 VGND.n4418 0 0.07f
C25331 VGND.n4419 0 0.0508f
C25332 VGND.n4420 0 0.0482f
C25333 VGND.n4421 0 0.00981f
C25334 VGND.n4422 0 0.0166f
C25335 VGND.n4423 0 0.0166f
C25336 VGND.n4424 0 0.059f
C25337 VGND.n4425 0 0.0166f
C25338 VGND.n4426 0 0.059f
C25339 VGND.n4427 0 0.0166f
C25340 VGND.n4428 0 0.0597f
C25341 VGND.n4429 0 0.0166f
C25342 VGND.n4430 0 0.0878f
C25343 VGND.n4431 0 0.0142f
C25344 VGND.n4432 0 0.00828f
C25345 VGND.n4433 0 0.00909f
C25346 VGND.n4434 0 0.00494f
C25347 VGND.n4435 0 0.00475f
C25348 VGND.n4436 0 0.00981f
C25349 VGND.n4437 0 0.0166f
C25350 VGND.n4438 0 0.0166f
C25351 VGND.n4439 0 0.0166f
C25352 VGND.n4440 0 0.00418f
C25353 VGND.n4441 0 0.0166f
C25354 VGND.n4442 0 0.00586f
C25355 VGND.n4443 0 0.0166f
C25356 VGND.n4444 0 0.015f
C25357 VGND.n4445 0 0.00828f
C25358 VGND.n4446 0 0.0474f
C25359 VGND.n4447 0 0.028f
C25360 VGND.n4448 0 0.00981f
C25361 VGND.n4449 0 0.0166f
C25362 VGND.n4450 0 0.0468f
C25363 VGND.n4451 0 0.0166f
C25364 VGND.n4452 0 0.0379f
C25365 VGND.n4453 0 0.0166f
C25366 VGND.n4454 0 0.00444f
C25367 VGND.n4455 0 0.0166f
C25368 VGND.n4456 0 0.0148f
C25369 VGND.n4457 0 0.00846f
C25370 VGND.n4458 0 8.29e-19
C25371 VGND.n4459 0 0.0289f
C25372 VGND.n4460 0 0.0269f
C25373 VGND.n4461 0 0.0081f
C25374 VGND.n4462 0 0.00783f
C25375 VGND.n4463 0 0.00171f
C25376 VGND.t243 0 0.0792f
C25377 VGND.n4464 0 0.0547f
C25378 VGND.n4465 0 0.0231f
C25379 VGND.n4466 0 9.9e-19
C25380 VGND.n4467 0 0.00189f
C25381 VGND.n4468 0 0.00162f
C25382 VGND.n4469 0 0.00342f
C25383 VGND.n4470 0 0.00387f
C25384 VGND.n4471 0 9.9e-19
C25385 VGND.n4472 0 0.00162f
C25386 VGND.n4473 0 0.0162f
C25387 VGND.n4474 0 0.00198f
C25388 VGND.n4475 0 0.003f
C25389 VGND.n4476 0 7.2e-19
C25390 VGND.n4477 0 9e-19
C25391 VGND.n4478 0 0.00282f
C25392 VGND.n4479 0 0.00135f
C25393 VGND.n4480 0 0.0118f
C25394 VGND.n4481 0 8.1e-19
C25395 VGND.n4482 0 0.00234f
C25396 VGND.n4483 0 0.00234f
C25397 VGND.n4484 0 0.00234f
C25398 VGND.n4485 0 7.2e-19
C25399 VGND.n4486 0 0.00252f
C25400 VGND.n4487 0 0.00369f
C25401 VGND.n4488 0 0.00189f
C25402 VGND.n4489 0 0.00135f
C25403 VGND.n4490 0 0.00207f
C25404 VGND.n4491 0 0.00126f
C25405 VGND.n4492 0 0.007f
C25406 VGND.n4493 0 0.00412f
C25407 VGND.n4494 0 0.00207f
C25408 VGND.n4495 0 0.00274f
C25409 VGND.n4496 0 0.00173f
C25410 VGND.n4497 0 0.00287f
C25411 VGND.n4498 0 0.00207f
C25412 VGND.n4499 0 0.00274f
C25413 VGND.n4500 0 0.00494f
C25414 VGND.n4501 0 0.00126f
C25415 VGND.n4502 0 0.00173f
C25416 VGND.n4503 0 0.00403f
C25417 VGND.n4504 0 0.00287f
C25418 VGND.n4505 0 0.00173f
C25419 VGND.n4506 0 0.00269f
C25420 VGND.n4507 0 0.0039f
C25421 VGND.n4508 0 0.00269f
C25422 VGND.n4509 0 0.00173f
C25423 VGND.n4510 0 0.178f
C25424 VGND.n4512 0 0.018f
C25425 VGND.n4514 0 0.317f
C25426 VGND.n4515 0 0.317f
C25427 VGND.n4516 0 0.00287f
C25428 VGND.n4517 0 0.00207f
C25429 VGND.n4518 0 0.00274f
C25430 VGND.n4519 0 0.00403f
C25431 VGND.n4520 0 0.00493f
C25432 VGND.n4521 0 0.00126f
C25433 VGND.n4522 0 0.00173f
C25434 VGND.n4524 0 0.018f
C25435 VGND.n4525 0 0.00274f
C25436 VGND.n4526 0 0.00173f
C25437 VGND.n4527 0 0.0041f
C25438 VGND.n4528 0 0.00701f
C25439 VGND.n4529 0 0.00207f
C25440 VGND.n4530 0 0.00207f
C25441 VGND.n4531 0 0.00162f
C25442 VGND.n4532 0 0.00234f
C25443 VGND.n4533 0 0.00144f
C25444 VGND.n4534 0 0.00297f
C25445 VGND.n4535 0 0.00234f
C25446 VGND.n4536 0 0.00234f
C25447 VGND.n4537 0 0.00234f
C25448 VGND.n4538 0 7.2e-19
C25449 VGND.n4539 0 0.00252f
C25450 VGND.n4540 0 0.00369f
C25451 VGND.n4541 0 0.00189f
C25452 VGND.n4542 0 0.00135f
C25453 VGND.n4543 0 0.00207f
C25454 VGND.n4544 0 0.00126f
C25455 VGND.n4545 0 0.00126f
C25456 VGND.n4546 0 0.00207f
C25457 VGND.n4547 0 0.00126f
C25458 VGND.n4548 0 1.12e-19
C25459 VGND.n4549 0 0.0382f
C25460 VGND.n4550 0 0.00828f
C25461 VGND.n4551 0 0.0119f
C25462 VGND.n4552 0 0.00981f
C25463 VGND.n4553 0 0.0543f
C25464 VGND.n4554 0 0.0375f
C25465 VGND.n4555 0 0.0324f
C25466 VGND.n4556 0 0.0528f
C25467 VGND.n4557 0 0.00981f
C25468 VGND.n4558 0 0.0166f
C25469 VGND.n4559 0 0.0331f
C25470 VGND.n4560 0 0.0166f
C25471 VGND.n4561 0 0.0379f
C25472 VGND.n4562 0 0.0166f
C25473 VGND.n4563 0 0.00444f
C25474 VGND.n4564 0 0.0166f
C25475 VGND.n4565 0 0.015f
C25476 VGND.n4566 0 0.0274f
C25477 VGND.n4567 0 0.0367f
C25478 VGND.n4568 0 0.186f
C25479 VGND.n4569 0 0.023f
C25480 VGND.n4570 0 0.00981f
C25481 VGND.n4571 0 0.0286f
C25482 VGND.n4572 0 0.0553f
C25483 VGND.n4573 0 0.00547f
C25484 VGND.n4574 0 0.0104f
C25485 VGND.n4575 0 0.0549f
C25486 VGND.n4576 0 0.0166f
C25487 VGND.n4577 0 0.0149f
C25488 VGND.n4578 0 0.0107f
C25489 VGND.n4579 0 0.0345f
C25490 VGND.n4580 0 0.0281f
C25491 VGND.n4581 0 0.00981f
C25492 VGND.n4582 0 0.0166f
C25493 VGND.n4583 0 0.0331f
C25494 VGND.n4584 0 0.0166f
C25495 VGND.n4585 0 0.0143f
C25496 VGND.n4586 0 0.009f
C25497 VGND.n4587 0 0.0336f
C25498 VGND.n4588 0 0.229f
C25499 VGND.n4589 0 0.229f
C25500 VGND.n4590 0 0.0251f
C25501 VGND.n4591 0 9.77e-19
C25502 VGND.n4592 0 0.00185f
C25503 VGND.n4593 0 1.46e-19
C25504 VGND.n4594 0 0.00198f
C25505 VGND.n4595 0 0.00162f
C25506 VGND.n4596 0 0.00189f
C25507 VGND.n4597 0 0.00162f
C25508 VGND.n4598 0 0.00342f
C25509 VGND.n4599 0 0.00387f
C25510 VGND.n4600 0 7.2e-19
C25511 VGND.n4601 0 7.2e-19
C25512 VGND.n4602 0 0.00207f
C25513 VGND.n4603 0 0.00315f
C25514 VGND.n4604 0 0.00162f
C25515 VGND.n4605 0 0.00162f
C25516 VGND.n4606 0 0.00189f
C25517 VGND.n4607 0 9.9e-19
C25518 VGND.n4608 0 0.00162f
C25519 VGND.n4609 0 0.00171f
C25520 VGND.n4610 0 0.00783f
C25521 VGND.n4611 0 0.0387f
C25522 VGND.n4612 0 0.0148f
C25523 VGND.t4 0 0.0792f
C25524 VGND.n4613 0 0.0547f
C25525 VGND.n4614 0 0.0243f
C25526 VGND.n4615 0 0.0166f
C25527 VGND.n4616 0 0.00981f
C25528 VGND.n4617 0 0.0291f
C25529 VGND.n4618 0 0.00437f
C25530 VGND.n4619 0 0.015f
C25531 VGND.n4620 0 0.0254f
C25532 VGND.n4621 0 0.0166f
C25533 VGND.n4622 0 0.00823f
C25534 VGND.n4623 0 0.0166f
C25535 VGND.n4624 0 0.026f
C25536 VGND.n4625 0 0.0166f
C25537 VGND.n4626 0 0.00821f
C25538 VGND.n4627 0 0.0166f
C25539 VGND.n4628 0 0.0285f
C25540 VGND.n4629 0 0.0166f
C25541 VGND.n4630 0 0.00586f
C25542 VGND.n4631 0 0.0166f
C25543 VGND.n4632 0 0.0285f
C25544 VGND.n4633 0 0.0166f
C25545 VGND.n4634 0 0.00821f
C25546 VGND.n4635 0 0.0166f
C25547 VGND.n4636 0 0.026f
C25548 VGND.n4637 0 0.0166f
C25549 VGND.n4638 0 0.00823f
C25550 VGND.n4639 0 0.0166f
C25551 VGND.n4640 0 0.0254f
C25552 VGND.n4641 0 0.0166f
C25553 VGND.n4642 0 0.00475f
C25554 VGND.n4643 0 0.0166f
C25555 VGND.n4644 0 0.00586f
C25556 VGND.n4645 0 0.0166f
C25557 VGND.n4646 0 0.0106f
C25558 VGND.n4647 0 0.00549f
C25559 VGND.n4648 0 0.053f
C25560 VGND.n4649 0 0.0435f
C25561 VGND.n4650 0 0.0142f
C25562 VGND.n4651 0 0.0166f
C25563 VGND.n4652 0 0.0324f
C25564 VGND.n4653 0 0.0166f
C25565 VGND.t375 0 0.157f
C25566 VGND.n4654 0 0.199f
C25567 VGND.n4655 0 0.0257f
C25568 VGND.n4656 0 0.0454f
C25569 VGND.n4657 0 0.0166f
C25570 VGND.n4658 0 0.0163f
C25571 VGND.n4659 0 0.0172f
C25572 VGND.n4660 0 0.009f
C25573 VGND.n4661 0 0.00819f
C25574 VGND.n4662 0 0.0377f
C25575 VGND.n4663 0 0.0772f
C25576 VGND.t190 0 0.125f
C25577 VGND.n4664 0 0.118f
C25578 VGND.n4665 0 0.0213f
C25579 VGND.n4666 0 0.00765f
C25580 VGND.t298 0 0.0792f
C25581 VGND.n4667 0 0.0547f
C25582 VGND.n4668 0 0.0319f
C25583 VGND.n4669 0 0.0874f
C25584 VGND.n4670 0 0.00828f
C25585 VGND.n4671 0 0.015f
C25586 VGND.n4672 0 0.00981f
C25587 VGND.n4673 0 0.00463f
C25588 VGND.n4674 0 0.0268f
C25589 VGND.n4675 0 0.015f
C25590 VGND.n4676 0 0.0299f
C25591 VGND.n4677 0 0.0166f
C25592 VGND.n4678 0 0.0242f
C25593 VGND.n4679 0 0.0328f
C25594 VGND.n4680 0 0.0249f
C25595 VGND.t189 0 0.0837f
C25596 VGND.n4681 0 0.325f
C25597 VGND.n4682 0 0.0312f
C25598 VGND.n4683 0 0.015f
C25599 VGND.n4684 0 0.0199f
C25600 VGND.n4685 0 0.0166f
C25601 VGND.n4686 0 0.0358f
C25602 VGND.n4687 0 0.0166f
C25603 VGND.n4688 0 0.0178f
C25604 VGND.n4689 0 0.0166f
C25605 VGND.n4690 0 0.0494f
C25606 VGND.n4691 0 0.0166f
C25607 VGND.n4692 0 0.0088f
C25608 VGND.n4693 0 0.0166f
C25609 VGND.n4694 0 0.031f
C25610 VGND.n4695 0 0.0166f
C25611 VGND.n4696 0 0.0126f
C25612 VGND.n4697 0 0.0166f
C25613 VGND.n4698 0 0.0317f
C25614 VGND.n4699 0 0.0166f
C25615 VGND.n4700 0 0.00513f
C25616 VGND.n4701 0 0.0166f
C25617 VGND.n4702 0 0.00981f
C25618 VGND.n4703 0 0.03f
C25619 VGND.n4704 0 0.0367f
C25620 VGND.n4705 0 0.015f
C25621 VGND.n4706 0 0.0468f
C25622 VGND.n4707 0 0.0166f
C25623 VGND.t266 0 0.0792f
C25624 VGND.n4708 0 0.0509f
C25625 VGND.n4709 0 0.034f
C25626 VGND.n4710 0 0.0153f
C25627 VGND.n4711 0 0.0127f
C25628 VGND.n4712 0 0.00828f
C25629 VGND.n4713 0 0.00153f
C25630 VGND.n4714 0 0.00423f
C25631 VGND.n4715 0 0.00126f
C25632 VGND.n4716 0 0.00912f
C25633 VGND.n4717 0 0.0101f
C25634 VGND.n4718 0 0.00126f
C25635 VGND.n4719 0 0.00824f
C25636 VGND.n4720 0 0.00234f
C25637 VGND.n4721 0 0.00297f
C25638 VGND.n4722 0 0.00315f
C25639 VGND.n4723 0 0.00207f
C25640 VGND.n4724 0 9.9e-19
C25641 VGND.n4725 0 0.00261f
C25642 VGND.n4726 0 0.00207f
C25643 VGND.n4727 0 0.00135f
C25644 VGND.n4728 0 7.2e-19
C25645 VGND.n4729 0 0.00126f
C25646 VGND.n4730 0 0.00135f
C25647 VGND.n4731 0 0.00126f
C25648 VGND.n4732 0 0.0254f
C25649 VGND.n4733 0 0.00198f
C25650 VGND.n4734 0 0.00453f
C25651 VGND.n4735 0 0.00153f
C25652 VGND.n4736 0 0.00282f
C25653 VGND.n4737 0 0.00144f
C25654 VGND.n4738 0 0.00651f
C25655 VGND.n4739 0 0.00261f
C25656 VGND.n4740 0 0.00234f
C25657 VGND.n4741 0 0.00234f
C25658 VGND.n4742 0 0.00225f
C25659 VGND.n4743 0 0.00144f
C25660 VGND.n4744 0 0.00148f
C25661 VGND.n4745 0 8.57e-19
C25662 VGND.n4746 0 0.0252f
C25663 VGND.n4747 0 0.229f
C25664 VGND.n4748 0 0.229f
C25665 VGND.n4749 0 0.00427f
C25666 VGND.n4750 0 0.0365f
C25667 VGND.t248 0 0.082f
C25668 VGND.n4751 0 0.0934f
C25669 VGND.n4752 0 0.0525f
C25670 VGND.n4753 0 0.038f
C25671 VGND.n4754 0 0.0217f
C25672 VGND.n4755 0 0.051f
C25673 VGND.t381 0 0.0816f
C25674 VGND.n4756 0 0.139f
C25675 VGND.n4757 0 0.0825f
C25676 VGND.n4758 0 0.00981f
C25677 VGND.t30 0 0.0792f
C25678 VGND.t121 0 0.0445f
C25679 VGND.n4759 0 0.0173f
C25680 VGND.t98 0 0.0445f
C25681 VGND.n4760 0 0.244f
C25682 VGND.n4761 0 0.0513f
C25683 VGND.n4762 0 0.057f
C25684 VGND.n4763 0 0.0249f
C25685 VGND.n4764 0 0.015f
C25686 VGND.n4765 0 0.00828f
C25687 VGND.n4766 0 0.00828f
C25688 VGND.n4767 0 0.0192f
C25689 VGND.t250 0 0.0799f
C25690 VGND.n4768 0 0.0723f
C25691 VGND.n4769 0 0.0241f
C25692 VGND.n4770 0 0.0533f
C25693 VGND.n4771 0 0.0166f
C25694 VGND.n4772 0 0.0362f
C25695 VGND.n4773 0 0.0166f
C25696 VGND.n4774 0 0.015f
C25697 VGND.n4775 0 0.00828f
C25698 VGND.n4776 0 0.0471f
C25699 VGND.n4777 0 0.00828f
C25700 VGND.n4778 0 0.0137f
C25701 VGND.n4779 0 0.0221f
C25702 VGND.n4780 0 0.015f
C25703 VGND.n4781 0 0.00828f
C25704 VGND.n4782 0 0.0339f
C25705 VGND.n4783 0 0.0458f
C25706 VGND.n4784 0 0.00981f
C25707 VGND.t64 0 0.0792f
C25708 VGND.n4785 0 0.0551f
C25709 VGND.n4786 0 0.0243f
C25710 VGND.n4787 0 0.0166f
C25711 VGND.n4788 0 0.053f
C25712 VGND.n4789 0 0.0166f
C25713 VGND.n4790 0 0.0423f
C25714 VGND.n4791 0 0.0166f
C25715 VGND.n4792 0 0.0166f
C25716 VGND.n4793 0 0.0149f
C25717 VGND.n4794 0 0.00837f
C25718 VGND.n4795 0 0.0345f
C25719 VGND.n4796 0 0.0281f
C25720 VGND.n4797 0 0.00981f
C25721 VGND.t25 0 0.0792f
C25722 VGND.n4798 0 0.0547f
C25723 VGND.n4799 0 0.034f
C25724 VGND.n4800 0 0.0166f
C25725 VGND.n4801 0 0.0166f
C25726 VGND.n4802 0 0.0143f
C25727 VGND.n4803 0 0.009f
C25728 VGND.n4804 0 0.026f
C25729 VGND.n4805 0 0.044f
C25730 VGND.n4806 0 0.00981f
C25731 VGND.n4807 0 0.0321f
C25732 VGND.n4808 0 0.0432f
C25733 VGND.n4809 0 0.0166f
C25734 VGND.t343 0 0.0946f
C25735 VGND.n4810 0 0.0183f
C25736 VGND.n4811 0 0.0961f
C25737 VGND.n4812 0 0.0341f
C25738 VGND.n4813 0 0.0271f
C25739 VGND.n4814 0 0.0166f
C25740 VGND.n4815 0 0.0345f
C25741 VGND.n4816 0 0.0252f
C25742 VGND.n4817 0 0.0166f
C25743 VGND.n4818 0 0.0316f
C25744 VGND.n4819 0 0.0166f
C25745 VGND.n4820 0 0.0166f
C25746 VGND.n4821 0 0.015f
C25747 VGND.n4822 0 0.00747f
C25748 VGND.n4823 0 0.0213f
C25749 VGND.t280 0 0.125f
C25750 VGND.n4824 0 0.118f
C25751 VGND.n4825 0 0.0391f
C25752 VGND.n4826 0 0.0277f
C25753 VGND.n4827 0 0.00981f
C25754 VGND.n4828 0 0.0166f
C25755 VGND.n4829 0 0.0151f
C25756 VGND.n4830 0 0.0379f
C25757 VGND.n4831 0 0.00437f
C25758 VGND.n4832 0 0.00972f
C25759 VGND.n4833 0 0.0166f
C25760 VGND.n4834 0 0.015f
C25761 VGND.n4835 0 0.0045f
C25762 VGND.n4836 0 0.0291f
C25763 VGND.n4837 0 0.00981f
C25764 VGND.t11 0 0.0792f
C25765 VGND.n4838 0 0.0547f
C25766 VGND.n4839 0 0.0243f
C25767 VGND.n4840 0 0.0166f
C25768 VGND.n4841 0 0.0166f
C25769 VGND.n4842 0 0.015f
C25770 VGND.n4843 0 0.0379f
C25771 VGND.n4844 0 0.0099f
C25772 VGND.n4845 0 0.00981f
C25773 VGND.n4846 0 0.0458f
C25774 VGND.n4847 0 0.0166f
C25775 VGND.n4848 0 0.015f
C25776 VGND.n4849 0 0.00549f
C25777 VGND.n4850 0 0.0435f
C25778 VGND.n4851 0 0.00981f
C25779 VGND.t211 0 0.0792f
C25780 VGND.n4852 0 0.0658f
C25781 VGND.n4853 0 0.0243f
C25782 VGND.n4854 0 0.0166f
C25783 VGND.n4855 0 0.0312f
C25784 VGND.n4856 0 0.0136f
C25785 VGND.n4857 0 0.0063f
C25786 VGND.n4858 0 0.00824f
C25787 VGND.n4859 0 0.00413f
C25788 VGND.n4860 0 0.018f
C25789 VGND.n4861 0 0.00269f
C25790 VGND.n4862 0 0.00207f
C25791 VGND.n4863 0 0.00287f
C25792 VGND.n4864 0 0.00173f
C25793 VGND.n4866 0 0.317f
C25794 VGND.n4867 0 0.317f
C25795 VGND.n4868 0 0.00173f
C25796 VGND.n4869 0 0.00269f
C25797 VGND.n4870 0 0.0039f
C25798 VGND.n4871 0 0.00269f
C25799 VGND.n4872 0 0.00207f
C25800 VGND.n4873 0 0.00287f
C25801 VGND.n4874 0 0.00173f
C25802 VGND.n4876 0 0.018f
C25803 VGND.n4877 0 0.00274f
C25804 VGND.n4878 0 0.00173f
C25805 VGND.n4879 0 0.00413f
C25806 VGND.n4880 0 0.00824f
C25807 VGND.n4881 0 0.0123f
C25808 VGND.t362 0 0.082f
C25809 VGND.n4882 0 0.0921f
C25810 VGND.n4883 0 0.0217f
C25811 VGND.n4884 0 0.0103f
C25812 VGND.n4885 0 0.0119f
C25813 VGND.n4886 0 0.0387f
C25814 VGND.n4887 0 0.00535f
C25815 VGND.n4888 0 0.015f
C25816 VGND.n4889 0 0.0242f
C25817 VGND.n4890 0 0.0166f
C25818 VGND.n4891 0 0.00821f
C25819 VGND.n4892 0 0.0166f
C25820 VGND.n4893 0 0.0285f
C25821 VGND.n4894 0 0.0166f
C25822 VGND.n4895 0 0.00586f
C25823 VGND.n4896 0 0.0166f
C25824 VGND.n4897 0 0.024f
C25825 VGND.n4898 0 0.0166f
C25826 VGND.n4899 0 0.00981f
C25827 VGND.n4900 0 0.00891f
C25828 VGND.n4901 0 0.0194f
C25829 VGND.n4902 0 0.0331f
C25830 VGND.n4903 0 0.0474f
C25831 VGND.n4904 0 0.0144f
C25832 VGND.n4905 0 0.0166f
C25833 VGND.n4906 0 0.0273f
C25834 VGND.n4907 0 0.0275f
C25835 VGND.n4908 0 0.019f
C25836 VGND.n4909 0 0.0316f
C25837 VGND.n4910 0 0.0264f
C25838 VGND.n4911 0 0.015f
C25839 VGND.n4912 0 0.0237f
C25840 VGND.n4913 0 0.0166f
C25841 VGND.n4914 0 0.0242f
C25842 VGND.n4915 0 0.00981f
C25843 VGND.n4916 0 0.023f
C25844 VGND.n4917 0 0.00489f
C25845 VGND.n4918 0 0.0309f
C25846 VGND.n4919 0 0.0251f
C25847 VGND.n4920 0 0.0319f
C25848 VGND.t116 0 0.0792f
C25849 VGND.n4921 0 0.0567f
C25850 VGND.n4922 0 0.0245f
C25851 VGND.n4923 0 0.053f
C25852 VGND.t255 0 0.128f
C25853 VGND.n4924 0 0.154f
C25854 VGND.n4925 0 0.0518f
C25855 VGND.n4926 0 0.0348f
C25856 VGND.t55 0 0.0445f
C25857 VGND.n4927 0 0.14f
C25858 VGND.t81 0 0.0445f
C25859 VGND.t62 0 0.0445f
C25860 VGND.n4928 0 0.243f
C25861 VGND.n4929 0 0.0173f
C25862 VGND.n4930 0 0.019f
C25863 VGND.n4931 0 0.0275f
C25864 VGND.n4932 0 0.015f
C25865 VGND.n4933 0 0.00828f
C25866 VGND.n4934 0 0.0638f
C25867 VGND.n4935 0 0.045f
C25868 VGND.n4936 0 0.00981f
C25869 VGND.n4937 0 0.0166f
C25870 VGND.n4938 0 0.015f
C25871 VGND.n4939 0 0.0375f
C25872 VGND.n4940 0 0.0448f
C25873 VGND.n4941 0 0.00981f
C25874 VGND.n4942 0 0.0446f
C25875 VGND.n4943 0 0.0471f
C25876 VGND.n4944 0 0.0166f
C25877 VGND.t6 0 0.0946f
C25878 VGND.n4945 0 0.0183f
C25879 VGND.n4946 0 0.0961f
C25880 VGND.n4947 0 0.0252f
C25881 VGND.n4948 0 0.0315f
C25882 VGND.n4949 0 0.0166f
C25883 VGND.n4950 0 0.0551f
C25884 VGND.n4951 0 0.0252f
C25885 VGND.n4952 0 0.0166f
C25886 VGND.n4953 0 0.0431f
C25887 VGND.n4954 0 0.0166f
C25888 VGND.n4955 0 0.046f
C25889 VGND.n4956 0 0.0166f
C25890 VGND.n4957 0 0.0166f
C25891 VGND.n4958 0 0.0489f
C25892 VGND.n4959 0 0.0466f
C25893 VGND.n4960 0 0.015f
C25894 VGND.n4961 0 0.0166f
C25895 VGND.n4962 0 0.0149f
C25896 VGND.n4963 0 0.00837f
C25897 VGND.n4964 0 0.0221f
C25898 VGND.n4965 0 0.009f
C25899 VGND.n4966 0 0.0428f
C25900 VGND.n4967 0 0.233f
C25901 VGND.n4968 0 0.229f
C25902 VGND.n4969 0 0.0944f
C25903 VGND.n4970 0 0.049f
C25904 VGND.n4971 0 0.229f
C25905 VGND.n4972 0 0.139f
C25906 VGND.n4973 0 0.094f
C25907 VGND.n4974 0 6.43f
C25908 VGND.n4975 0 7.18f
C25909 VGND.n4976 0 0.0749f
C25910 VGND.n4977 0 0.0707f
C25911 VGND.n4978 0 0.0783f
C25912 VGND.n4979 0 0.0911f
C25913 VGND.n4980 0 0.0849f
C25914 VGND.n4981 0 0.0811f
C25915 VGND.n4982 0 0.0821f
C25916 VGND.n4983 0 0.0778f
C25917 VGND.n4984 0 0.0859f
C25918 VGND.n4985 0 0.0897f
C25919 VGND.n4986 0 0.0441f
C25920 VGND.n4987 0 0.992f
C25921 VGND.n4988 0 0.101f
C25922 VGND.n4989 0 0.178f
C25923 VGND.n4990 0 0.178f
C25924 VGND.n4991 0 0.0835f
C25925 VGND.n4992 0 0.178f
C25926 VGND.n4993 0 0.178f
C25927 VGND.n4994 0 0.0835f
C25928 VGND.n4995 0 0.178f
C25929 VGND.n4996 0 0.178f
C25930 VGND.n4997 0 0.0835f
C25931 VGND.n4998 0 0.178f
C25932 VGND.n4999 0 0.178f
C25933 VGND.n5000 0 0.0835f
C25934 VGND.n5001 0 0.178f
C25935 VGND.n5002 0 0.178f
C25936 VGND.n5003 0 0.0835f
C25937 VGND.n5004 0 0.178f
C25938 VGND.n5005 0 0.178f
C25939 VGND.n5006 0 0.0835f
C25940 VGND.n5007 0 0.178f
C25941 VGND.n5008 0 0.178f
C25942 VGND.n5009 0 0.0835f
C25943 VGND.n5010 0 0.178f
C25944 VGND.n5011 0 0.178f
C25945 VGND.n5012 0 0.0835f
C25946 VGND.n5013 0 0.178f
C25947 VGND.n5014 0 0.178f
C25948 VGND.n5015 0 0.0835f
C25949 VGND.n5016 0 0.178f
C25950 VGND.n5017 0 0.178f
C25951 VGND.n5018 0 0.0835f
C25952 VGND.n5019 0 0.229f
C25953 VGND.n5020 0 0.229f
C25954 VGND.n5021 0 0.0279f
C25955 VGND.n5022 0 8.57e-19
C25956 VGND.n5023 0 0.00126f
C25957 VGND.n5024 0 0.00135f
C25958 VGND.n5025 0 0.00126f
C25959 VGND.n5026 0 7.2e-19
C25960 VGND.n5027 0 9.9e-19
C25961 VGND.n5028 0 0.00207f
C25962 VGND.n5029 0 0.00315f
C25963 VGND.n5030 0 0.00297f
C25964 VGND.n5031 0 0.00234f
C25965 VGND.n5032 0 0.00824f
C25966 VGND.n5033 0 0.00126f
C25967 VGND.n5034 0 0.00153f
C25968 VGND.n5035 0 0.00828f
C25969 VGND.n5036 0 0.0378f
C25970 VGND.n5037 0 0.0108f
C25971 VGND.n5038 0 0.0227f
C25972 VGND.n5039 0 0.0273f
C25973 VGND.n5040 0 0.0271f
C25974 VGND.n5041 0 0.0153f
C25975 VGND.t46 0 0.0946f
C25976 VGND.n5042 0 0.0183f
C25977 VGND.n5043 0 0.0961f
C25978 VGND.n5044 0 0.0252f
C25979 VGND.n5045 0 0.0271f
C25980 VGND.n5046 0 0.0166f
C25981 VGND.n5047 0 0.0345f
C25982 VGND.n5048 0 0.0252f
C25983 VGND.n5049 0 0.0166f
C25984 VGND.n5050 0 0.0453f
C25985 VGND.n5051 0 0.0166f
C25986 VGND.n5052 0 0.0421f
C25987 VGND.n5053 0 0.0166f
C25988 VGND.n5054 0 0.0331f
C25989 VGND.n5055 0 0.0166f
C25990 VGND.n5056 0 0.015f
C25991 VGND.n5057 0 0.0379f
C25992 VGND.n5058 0 0.00437f
C25993 VGND.n5059 0 0.00981f
C25994 VGND.n5060 0 0.0166f
C25995 VGND.n5061 0 0.0104f
C25996 VGND.n5062 0 0.0166f
C25997 VGND.n5063 0 0.0457f
C25998 VGND.n5064 0 0.0166f
C25999 VGND.n5065 0 0.0104f
C26000 VGND.n5066 0 0.0166f
C26001 VGND.n5067 0 0.015f
C26002 VGND.n5068 0 0.00828f
C26003 VGND.n5069 0 0.00437f
C26004 VGND.n5070 0 0.0291f
C26005 VGND.n5071 0 0.00981f
C26006 VGND.n5072 0 0.0166f
C26007 VGND.n5073 0 0.0428f
C26008 VGND.n5074 0 0.0166f
C26009 VGND.n5075 0 0.0508f
C26010 VGND.n5076 0 0.015f
C26011 VGND.n5077 0 0.00981f
C26012 VGND.n5078 0 0.00427f
C26013 VGND.n5079 0 0.0166f
C26014 VGND.n5080 0 0.015f
C26015 VGND.n5081 0 0.0191f
C26016 VGND.n5082 0 0.0273f
C26017 VGND.n5083 0 0.0275f
C26018 VGND.n5084 0 0.0499f
C26019 VGND.n5085 0 0.0166f
C26020 VGND.n5086 0 0.0375f
C26021 VGND.n5087 0 0.0143f
C26022 VGND.n5088 0 0.00828f
C26023 VGND.n5089 0 0.0172f
C26024 VGND.n5090 0 0.0349f
C26025 VGND.n5091 0 0.139f
C26026 VGND.n5092 0 0.0105f
C26027 VGND.n5093 0 0.00837f
C26028 VGND.n5094 0 0.00972f
C26029 VGND.n5095 0 0.0166f
C26030 VGND.n5096 0 0.0166f
C26031 VGND.n5097 0 0.00418f
C26032 VGND.n5098 0 0.0166f
C26033 VGND.n5099 0 0.00586f
C26034 VGND.n5100 0 0.0166f
C26035 VGND.n5101 0 0.00586f
C26036 VGND.n5102 0 0.0166f
C26037 VGND.n5103 0 0.00462f
C26038 VGND.n5104 0 0.0166f
C26039 VGND.n5105 0 0.015f
C26040 VGND.n5106 0 0.0386f
C26041 VGND.n5107 0 0.028f
C26042 VGND.n5108 0 0.00981f
C26043 VGND.t141 0 0.0792f
C26044 VGND.n5109 0 0.074f
C26045 VGND.n5110 0 0.0284f
C26046 VGND.n5111 0 0.0166f
C26047 VGND.n5112 0 0.0166f
C26048 VGND.n5113 0 0.0144f
C26049 VGND.n5114 0 0.0379f
C26050 VGND.n5115 0 0.00549f
C26051 VGND.n5116 0 0.0104f
C26052 VGND.n5117 0 0.0209f
C26053 VGND.n5118 0 0.0166f
C26054 VGND.n5119 0 0.0166f
C26055 VGND.n5120 0 0.00504f
C26056 VGND.n5121 0 0.0166f
C26057 VGND.n5122 0 0.00504f
C26058 VGND.n5123 0 0.0166f
C26059 VGND.n5124 0 0.0166f
C26060 VGND.n5125 0 0.015f
C26061 VGND.n5126 0 0.0205f
C26062 VGND.n5127 0 0.0291f
C26063 VGND.n5128 0 0.00981f
C26064 VGND.t213 0 0.0792f
C26065 VGND.n5129 0 0.0547f
C26066 VGND.n5130 0 0.0243f
C26067 VGND.n5131 0 0.0166f
C26068 VGND.n5132 0 0.0148f
C26069 VGND.n5133 0 0.00783f
C26070 VGND.n5134 0 0.00207f
C26071 VGND.n5135 0 0.00315f
C26072 VGND.n5136 0 0.00162f
C26073 VGND.n5137 0 0.00162f
C26074 VGND.n5138 0 0.00189f
C26075 VGND.n5139 0 9.9e-19
C26076 VGND.n5140 0 0.00162f
C26077 VGND.n5141 0 0.00171f
C26078 VGND.n5142 0 0.0549f
C26079 VGND.n5143 0 9.9e-19
C26080 VGND.n5144 0 0.00189f
C26081 VGND.n5145 0 0.00162f
C26082 VGND.n5146 0 0.00342f
C26083 VGND.n5147 0 0.00387f
C26084 VGND.n5148 0 7.2e-19
C26085 VGND.n5149 0 0.00162f
C26086 VGND.n5150 0 0.00207f
C26087 VGND.n5151 0 0.00207f
C26088 VGND.n5152 0 0.00162f
C26089 VGND.n5153 0 0.00234f
C26090 VGND.n5154 0 0.00234f
C26091 VGND.n5155 0 0.00234f
C26092 VGND.n5156 0 0.00297f
C26093 VGND.n5157 0 0.00887f
C26094 VGND.n5158 0 0.00144f
C26095 VGND.n5159 0 0.00135f
C26096 VGND.n5160 0 2.7e-19
C26097 VGND.n5161 0 0.003f
C26098 VGND.n5162 0 0.0179f
C26099 VGND.n5163 0 0.00126f
C26100 VGND.n5164 0 0.00207f
C26101 VGND.n5165 0 0.00126f
C26102 VGND.n5166 0 0.00126f
C26103 VGND.n5167 0 0.00701f
C26104 VGND.n5168 0 0.0041f
C26105 VGND.n5169 0 0.018f
C26106 VGND.n5170 0 0.00207f
C26107 VGND.n5171 0 0.00287f
C26108 VGND.n5172 0 0.00173f
C26109 VGND.n5173 0 0.00269f
C26110 VGND.n5174 0 0.0039f
C26111 VGND.n5175 0 0.00269f
C26112 VGND.n5176 0 0.00173f
C26113 VGND.n5178 0 0.317f
C26114 VGND.n5179 0 0.317f
C26115 VGND.n5181 0 0.0198f
C26116 VGND.n5183 0 0.018f
C26117 VGND.n5184 0 0.00403f
C26118 VGND.n5185 0 0.00173f
C26119 VGND.n5186 0 0.00274f
C26120 VGND.n5187 0 0.00207f
C26121 VGND.n5188 0 0.00287f
C26122 VGND.n5189 0 0.00173f
C26123 VGND.n5190 0 0.00269f
C26124 VGND.n5191 0 0.0039f
C26125 VGND.n5192 0 0.00269f
C26126 VGND.n5193 0 0.00173f
C26127 VGND.n5194 0 0.00287f
C26128 VGND.n5195 0 0.00207f
C26129 VGND.n5196 0 0.00274f
C26130 VGND.n5197 0 0.00173f
C26131 VGND.n5198 0 0.0041f
C26132 VGND.n5199 0 0.00701f
C26133 VGND.n5200 0 0.0452f
C26134 VGND.n5201 0 0.0278f
C26135 VGND.n5202 0 0.0143f
C26136 VGND.n5203 0 0.0166f
C26137 VGND.t354 0 0.0792f
C26138 VGND.n5204 0 0.0547f
C26139 VGND.n5205 0 0.0243f
C26140 VGND.n5206 0 0.0166f
C26141 VGND.n5207 0 0.00981f
C26142 VGND.n5208 0 0.028f
C26143 VGND.n5209 0 0.0261f
C26144 VGND.n5210 0 0.015f
C26145 VGND.n5211 0 0.00373f
C26146 VGND.n5212 0 0.0166f
C26147 VGND.n5213 0 0.0166f
C26148 VGND.n5214 0 0.00462f
C26149 VGND.n5215 0 0.0331f
C26150 VGND.n5216 0 0.0376f
C26151 VGND.n5217 0 0.015f
C26152 VGND.n5218 0 0.0166f
C26153 VGND.n5219 0 0.0324f
C26154 VGND.n5220 0 0.0166f
C26155 VGND.n5221 0 0.0324f
C26156 VGND.n5222 0 0.0166f
C26157 VGND.n5223 0 0.0324f
C26158 VGND.n5224 0 0.0166f
C26159 VGND.n5225 0 0.0316f
C26160 VGND.n5226 0 0.0166f
C26161 VGND.n5227 0 0.0393f
C26162 VGND.n5228 0 0.0252f
C26163 VGND.n5229 0 0.025f
C26164 VGND.n5230 0 0.0166f
C26165 VGND.n5231 0 0.0176f
C26166 VGND.n5232 0 0.0252f
C26167 VGND.n5233 0 0.035f
C26168 VGND.n5234 0 0.0166f
C26169 VGND.n5235 0 0.035f
C26170 VGND.n5236 0 0.0166f
C26171 VGND.t33 0 0.151f
C26172 VGND.n5237 0 0.126f
C26173 VGND.n5238 0 0.0274f
C26174 VGND.n5239 0 0.0252f
C26175 VGND.n5240 0 0.0279f
C26176 VGND.n5241 0 0.0166f
C26177 VGND.n5242 0 0.0342f
C26178 VGND.n5243 0 0.0323f
C26179 VGND.n5244 0 0.0166f
C26180 VGND.n5245 0 0.00981f
C26181 VGND.n5246 0 0.00459f
C26182 VGND.n5247 0 0.0278f
C26183 VGND.n5248 0 0.015f
C26184 VGND.n5249 0 0.00373f
C26185 VGND.n5250 0 0.0166f
C26186 VGND.n5251 0 0.0261f
C26187 VGND.n5252 0 0.0166f
C26188 VGND.n5253 0 0.0368f
C26189 VGND.n5254 0 0.0166f
C26190 VGND.n5255 0 0.0331f
C26191 VGND.n5256 0 0.0166f
C26192 VGND.t61 0 0.0792f
C26193 VGND.n5257 0 0.0547f
C26194 VGND.n5258 0 0.0243f
C26195 VGND.n5259 0 0.0166f
C26196 VGND.n5260 0 0.0279f
C26197 VGND.n5261 0 0.00981f
C26198 VGND.n5262 0 0.009f
C26199 VGND.n5263 0 0.00378f
C26200 VGND.n5264 0 0.00207f
C26201 VGND.n5265 0 0.00135f
C26202 VGND.n5266 0 2.7e-19
C26203 VGND.n5267 0 0.00219f
C26204 VGND.n5268 0 5.42e-19
C26205 VGND.n5269 0 0.00201f
C26206 VGND.n5270 0 0.00126f
C26207 VGND.n5271 0 0.00207f
C26208 VGND.n5272 0 0.00126f
C26209 VGND.n5273 0 0.00126f
C26210 VGND.n5274 0 0.00207f
C26211 VGND.n5275 0 0.00135f
C26212 VGND.n5276 0 0.00189f
C26213 VGND.n5277 0 0.00369f
C26214 VGND.n5278 0 0.00252f
C26215 VGND.n5279 0 7.2e-19
C26216 VGND.n5280 0 0.00493f
C26217 VGND.n5281 0 0.00126f
C26218 VGND.n5282 0 0.00162f
C26219 VGND.n5283 0 9.9e-19
C26220 VGND.n5284 0 0.00189f
C26221 VGND.n5285 0 0.00162f
C26222 VGND.n5286 0 0.00162f
C26223 VGND.n5287 0 0.00315f
C26224 VGND.n5288 0 0.00207f
C26225 VGND.n5289 0 7.2e-19
C26226 VGND.n5290 0 7.2e-19
C26227 VGND.n5291 0 0.00162f
C26228 VGND.n5292 0 0.00207f
C26229 VGND.n5293 0 0.00207f
C26230 VGND.n5294 0 0.00162f
C26231 VGND.n5295 0 0.00234f
C26232 VGND.n5296 0 0.00234f
C26233 VGND.n5297 0 0.00234f
C26234 VGND.n5298 0 0.00234f
C26235 VGND.n5299 0 0.00699f
C26236 VGND.n5300 0 8.1e-19
C26237 VGND.n5301 0 0.00282f
C26238 VGND.n5302 0 0.00135f
C26239 VGND.n5303 0 9e-19
C26240 VGND.n5304 0 0.00453f
C26241 VGND.n5305 0 7.2e-19
C26242 VGND.n5306 0 0.0254f
C26243 VGND.n5307 0 0.00198f
C26244 VGND.n5308 0 0.00162f
C26245 VGND.n5309 0 9.9e-19
C26246 VGND.n5310 0 0.00387f
C26247 VGND.n5311 0 0.00342f
C26248 VGND.n5312 0 0.00162f
C26249 VGND.n5313 0 0.00189f
C26250 VGND.n5314 0 0.0312f
C26251 VGND.n5315 0 9.9e-19
C26252 VGND.n5316 0 0.00171f
C26253 VGND.n5317 0 0.00783f
C26254 VGND.n5318 0 0.0324f
C26255 VGND.n5319 0 0.0148f
C26256 VGND.n5320 0 0.0316f
C26257 VGND.n5321 0 0.0166f
C26258 VGND.n5322 0 0.0345f
C26259 VGND.n5323 0 0.0252f
C26260 VGND.n5324 0 0.0166f
C26261 VGND.t72 0 0.0946f
C26262 VGND.n5325 0 0.0183f
C26263 VGND.n5326 0 0.0961f
C26264 VGND.n5327 0 0.0252f
C26265 VGND.n5328 0 0.0271f
C26266 VGND.n5329 0 0.0166f
C26267 VGND.n5330 0 0.0321f
C26268 VGND.n5331 0 0.0271f
C26269 VGND.n5332 0 0.0166f
C26270 VGND.n5333 0 0.00981f
C26271 VGND.n5334 0 0.00459f
C26272 VGND.n5335 0 0.0278f
C26273 VGND.n5336 0 0.015f
C26274 VGND.n5337 0 0.00373f
C26275 VGND.n5338 0 0.0166f
C26276 VGND.n5339 0 0.0261f
C26277 VGND.n5340 0 0.0166f
C26278 VGND.n5341 0 0.0368f
C26279 VGND.n5342 0 0.0166f
C26280 VGND.n5343 0 0.0331f
C26281 VGND.n5344 0 0.0166f
C26282 VGND.t268 0 0.0792f
C26283 VGND.n5345 0 0.0547f
C26284 VGND.n5346 0 0.0243f
C26285 VGND.n5347 0 0.0166f
C26286 VGND.n5348 0 0.00981f
C26287 VGND.n5349 0 0.0291f
C26288 VGND.n5350 0 0.00549f
C26289 VGND.n5351 0 0.015f
C26290 VGND.n5352 0 0.00658f
C26291 VGND.n5353 0 0.0166f
C26292 VGND.n5354 0 0.0194f
C26293 VGND.n5355 0 0.0166f
C26294 VGND.n5356 0 0.00619f
C26295 VGND.n5357 0 0.0166f
C26296 VGND.n5358 0 0.00981f
C26297 VGND.n5359 0 0.0225f
C26298 VGND.n5360 0 0.0331f
C26299 VGND.n5361 0 0.0379f
C26300 VGND.n5362 0 0.015f
C26301 VGND.n5363 0 0.0166f
C26302 VGND.n5364 0 0.0273f
C26303 VGND.n5365 0 0.0275f
C26304 VGND.n5366 0 0.019f
C26305 VGND.n5367 0 0.009f
C26306 VGND.n5368 0 0.00456f
C26307 VGND.n5369 0 0.00819f
C26308 VGND.n5370 0 0.0379f
C26309 VGND.n5371 0 0.0144f
C26310 VGND.n5372 0 0.0331f
C26311 VGND.n5373 0 0.0166f
C26312 VGND.n5374 0 0.0324f
C26313 VGND.n5375 0 0.0166f
C26314 VGND.n5376 0 0.0316f
C26315 VGND.n5377 0 0.0166f
C26316 VGND.n5378 0 0.0345f
C26317 VGND.n5379 0 0.0252f
C26318 VGND.n5380 0 0.0166f
C26319 VGND.n5381 0 0.0166f
C26320 VGND.n5382 0 0.0166f
C26321 VGND.n5383 0 0.00981f
C26322 VGND.n5384 0 0.00459f
C26323 VGND.n5385 0 0.0278f
C26324 VGND.n5386 0 0.015f
C26325 VGND.n5387 0 0.00373f
C26326 VGND.n5388 0 0.0166f
C26327 VGND.n5389 0 0.0261f
C26328 VGND.n5390 0 0.0166f
C26329 VGND.n5391 0 0.0368f
C26330 VGND.n5392 0 0.0166f
C26331 VGND.n5393 0 0.0331f
C26332 VGND.n5394 0 0.0166f
C26333 VGND.n5395 0 0.0324f
C26334 VGND.n5396 0 0.0166f
C26335 VGND.n5397 0 0.0316f
C26336 VGND.n5398 0 0.0166f
C26337 VGND.n5399 0 0.0345f
C26338 VGND.n5400 0 0.0252f
C26339 VGND.n5401 0 0.0166f
C26340 VGND.n5402 0 0.0166f
C26341 VGND.n5403 0 0.0166f
C26342 VGND.n5404 0 0.00981f
C26343 VGND.n5405 0 0.0452f
C26344 VGND.n5406 0 0.00439f
C26345 VGND.n5407 0 0.015f
C26346 VGND.n5408 0 0.0287f
C26347 VGND.n5409 0 0.0166f
C26348 VGND.n5410 0 0.00981f
C26349 VGND.n5411 0 0.00444f
C26350 VGND.n5412 0 0.0379f
C26351 VGND.n5413 0 0.015f
C26352 VGND.n5414 0 0.0331f
C26353 VGND.n5415 0 0.0166f
C26354 VGND.n5416 0 0.0166f
C26355 VGND.t322 0 0.0792f
C26356 VGND.n5417 0 0.0243f
C26357 VGND.n5418 0 0.0547f
C26358 VGND.n5419 0 0.0279f
C26359 VGND.n5420 0 0.00981f
C26360 VGND.n5421 0 0.00611f
C26361 VGND.n5422 0 0.0162f
C26362 VGND.n5423 0 0.00198f
C26363 VGND.n5424 0 0.003f
C26364 VGND.n5425 0 0.00153f
C26365 VGND.n5426 0 0.00282f
C26366 VGND.n5427 0 0.00144f
C26367 VGND.n5428 0 0.0118f
C26368 VGND.n5429 0 0.00261f
C26369 VGND.n5430 0 0.00234f
C26370 VGND.n5431 0 0.00234f
C26371 VGND.n5432 0 0.00315f
C26372 VGND.n5433 0 0.0177f
C26373 VGND.n5434 0 0.00162f
C26374 VGND.n5435 0 0.00135f
C26375 VGND.n5436 0 9.9e-19
C26376 VGND.n5437 0 0.00943f
C26377 VGND.n5438 0 0.0102f
C26378 VGND.n5439 0 0.00126f
C26379 VGND.n5440 0 0.00135f
C26380 VGND.n5441 0 0.00126f
C26381 VGND.n5442 0 0.00414f
C26382 VGND.n5443 0 0.00351f
C26383 VGND.n5444 0 0.00198f
C26384 VGND.n5445 0 0.00235f
C26385 VGND.n5446 0 0.00824f
C26386 VGND.n5447 0 0.00413f
C26387 VGND.n5448 0 0.0198f
C26388 VGND.n5449 0 0.00207f
C26389 VGND.n5450 0 0.00287f
C26390 VGND.n5451 0 0.00269f
C26391 VGND.n5452 0 0.00173f
C26392 VGND.n5454 0 0.018f
C26393 VGND.n5455 0 0.00413f
C26394 VGND.n5456 0 0.00824f
C26395 VGND.n5457 0 0.0063f
C26396 VGND.t253 0 0.0792f
C26397 VGND.n5458 0 0.0547f
C26398 VGND.n5459 0 0.0231f
C26399 VGND.n5460 0 0.0136f
C26400 VGND.n5461 0 0.00981f
C26401 VGND.n5462 0 0.028f
C26402 VGND.n5463 0 0.0261f
C26403 VGND.n5464 0 0.015f
C26404 VGND.n5465 0 0.00373f
C26405 VGND.n5466 0 0.0166f
C26406 VGND.n5467 0 0.0166f
C26407 VGND.n5468 0 0.00463f
C26408 VGND.n5469 0 0.0331f
C26409 VGND.n5470 0 0.0379f
C26410 VGND.n5471 0 0.015f
C26411 VGND.n5472 0 0.0166f
C26412 VGND.t295 0 0.0792f
C26413 VGND.n5473 0 0.0547f
C26414 VGND.n5474 0 0.0243f
C26415 VGND.n5475 0 0.0166f
C26416 VGND.n5476 0 0.00981f
C26417 VGND.n5477 0 0.00463f
C26418 VGND.n5478 0 0.0278f
C26419 VGND.n5479 0 0.015f
C26420 VGND.n5480 0 0.00373f
C26421 VGND.n5481 0 0.0166f
C26422 VGND.n5482 0 0.0261f
C26423 VGND.n5483 0 0.0166f
C26424 VGND.n5484 0 0.0368f
C26425 VGND.n5485 0 0.0166f
C26426 VGND.n5486 0 0.0331f
C26427 VGND.n5487 0 0.0166f
C26428 VGND.t330 0 0.0792f
C26429 VGND.n5488 0 0.0547f
C26430 VGND.n5489 0 0.0243f
C26431 VGND.n5490 0 0.0166f
C26432 VGND.n5491 0 0.00981f
C26433 VGND.n5492 0 0.00463f
C26434 VGND.n5493 0 0.0278f
C26435 VGND.n5494 0 0.015f
C26436 VGND.n5495 0 0.00373f
C26437 VGND.n5496 0 0.0166f
C26438 VGND.n5497 0 0.0261f
C26439 VGND.n5498 0 0.0166f
C26440 VGND.n5499 0 0.0368f
C26441 VGND.n5500 0 0.0166f
C26442 VGND.n5501 0 0.0331f
C26443 VGND.n5502 0 0.0166f
C26444 VGND.t227 0 0.0792f
C26445 VGND.n5503 0 0.0547f
C26446 VGND.n5504 0 0.0243f
C26447 VGND.n5505 0 0.0166f
C26448 VGND.n5506 0 0.00981f
C26449 VGND.n5507 0 0.009f
C26450 VGND.n5508 0 0.0331f
C26451 VGND.n5509 0 0.0278f
C26452 VGND.n5510 0 0.0261f
C26453 VGND.n5511 0 0.0278f
C26454 VGND.n5512 0 0.0261f
C26455 VGND.t349 0 0.128f
C26456 VGND.n5513 0 0.154f
C26457 VGND.n5514 0 0.0271f
C26458 VGND.n5515 0 0.0285f
C26459 VGND.n5516 0 0.0362f
C26460 VGND.t276 0 0.0409f
C26461 VGND.n5517 0 0.062f
C26462 VGND.n5518 0 0.0151f
C26463 VGND.n5519 0 0.0166f
C26464 VGND.n5520 0 0.015f
C26465 VGND.n5521 0 0.0191f
C26466 VGND.n5522 0 0.0273f
C26467 VGND.n5523 0 0.0275f
C26468 VGND.n5524 0 0.0331f
C26469 VGND.n5525 0 0.0166f
C26470 VGND.n5526 0 0.0368f
C26471 VGND.n5527 0 0.0166f
C26472 VGND.n5528 0 0.0166f
C26473 VGND.n5529 0 0.00373f
C26474 VGND.n5530 0 0.0166f
C26475 VGND.n5531 0 0.015f
C26476 VGND.n5532 0 0.00463f
C26477 VGND.n5533 0 0.0291f
C26478 VGND.n5534 0 0.00981f
C26479 VGND.t296 0 0.0792f
C26480 VGND.n5535 0 0.0547f
C26481 VGND.n5536 0 0.0243f
C26482 VGND.n5537 0 0.0166f
C26483 VGND.n5538 0 0.0331f
C26484 VGND.n5539 0 0.0166f
C26485 VGND.n5540 0 0.0368f
C26486 VGND.n5541 0 0.0166f
C26487 VGND.n5542 0 0.0166f
C26488 VGND.n5543 0 0.00373f
C26489 VGND.n5544 0 0.0166f
C26490 VGND.n5545 0 0.015f
C26491 VGND.n5546 0 0.00459f
C26492 VGND.n5547 0 0.0452f
C26493 VGND.n5548 0 0.00981f
C26494 VGND.n5549 0 0.0321f
C26495 VGND.n5550 0 0.0271f
C26496 VGND.n5551 0 0.0166f
C26497 VGND.t254 0 0.0946f
C26498 VGND.n5552 0 0.0183f
C26499 VGND.n5553 0 0.0961f
C26500 VGND.n5554 0 0.0252f
C26501 VGND.n5555 0 0.0271f
C26502 VGND.n5556 0 0.0166f
C26503 VGND.n5557 0 0.0345f
C26504 VGND.n5558 0 0.0252f
C26505 VGND.n5559 0 0.0166f
C26506 VGND.n5560 0 0.0316f
C26507 VGND.n5561 0 0.0166f
C26508 VGND.n5562 0 0.0324f
C26509 VGND.n5563 0 0.0166f
C26510 VGND.n5564 0 0.0166f
C26511 VGND.n5565 0 0.0143f
C26512 VGND.n5566 0 0.0367f
C26513 VGND.n5567 0 0.026f
C26514 VGND.n5568 0 0.939f
C26515 VGND.n5569 0 0.524f
C26516 VGND.n5570 0 0.213f
C26517 VGND.n5571 0 0.213f
C26518 VGND.n5572 0 0.524f
C26519 VGND.n5573 0 0.0252f
C26520 VGND.n5574 0 0.009f
C26521 VGND.n5575 0 0.019f
C26522 VGND.n5576 0 0.0273f
C26523 VGND.n5577 0 0.0275f
C26524 VGND.n5578 0 0.0166f
C26525 VGND.n5579 0 0.015f
C26526 VGND.n5580 0 0.0379f
C26527 VGND.n5581 0 0.00463f
C26528 VGND.n5582 0 0.0166f
C26529 VGND.n5583 0 0.00373f
C26530 VGND.n5584 0 0.0166f
C26531 VGND.n5585 0 0.015f
C26532 VGND.n5586 0 0.0261f
C26533 VGND.n5587 0 0.028f
C26534 VGND.n5588 0 0.00981f
C26535 VGND.t10 0 0.0792f
C26536 VGND.n5589 0 0.0547f
C26537 VGND.n5590 0 0.0243f
C26538 VGND.n5591 0 0.0166f
C26539 VGND.n5592 0 0.0166f
C26540 VGND.n5593 0 0.015f
C26541 VGND.n5594 0 0.0379f
C26542 VGND.n5595 0 0.00463f
C26543 VPWR.t374 0 0.0774f
C26544 VPWR.t288 0 0.0417f
C26545 VPWR.t260 0 0.0417f
C26546 VPWR.n0 0 0.383f
C26547 VPWR.n1 0 0.0384f
C26548 VPWR.n2 0 0.0421f
C26549 VPWR.t90 0 0.0774f
C26550 VPWR.n3 0 0.501f
C26551 VPWR.n4 0 0.0809f
C26552 VPWR.n5 0 0.018f
C26553 VPWR.n6 0 0.00429f
C26554 VPWR.n7 0 0.0199f
C26555 VPWR.n8 0 0.114f
C26556 VPWR.n9 0 0.0199f
C26557 VPWR.t10 0 0.0774f
C26558 VPWR.n10 0 0.0276f
C26559 VPWR.t123 0 0.0774f
C26560 VPWR.n11 0 0.0518f
C26561 VPWR.n12 0 0.0457f
C26562 VPWR.n13 0 0.0949f
C26563 VPWR.t111 0 0.0949f
C26564 VPWR.n14 0 0.101f
C26565 VPWR.n15 0 0.0331f
C26566 VPWR.n16 0 0.0369f
C26567 VPWR.n17 0 0.0214f
C26568 VPWR.n18 0 0.0483f
C26569 VPWR.t24 0 0.0876f
C26570 VPWR.n19 0 0.0987f
C26571 VPWR.n20 0 0.0973f
C26572 VPWR.n21 0 0.0973f
C26573 VPWR.n22 0 0.168f
C26574 VPWR.n23 0 0.0772f
C26575 VPWR.n24 0 0.13f
C26576 VPWR.n25 0 0.0271f
C26577 VPWR.n26 0 0.00851f
C26578 VPWR.n27 0 0.0014f
C26579 VPWR.n28 0 0.00151f
C26580 VPWR.n29 0 0.00162f
C26581 VPWR.n30 0 0.00378f
C26582 VPWR.n31 0 0.00497f
C26583 VPWR.n32 0 0.00417f
C26584 VPWR.n33 0 0.00248f
C26585 VPWR.n34 0 0.00335f
C26586 VPWR.n35 0 0.00421f
C26587 VPWR.n36 0 0.00248f
C26588 VPWR.n37 0 5.4e-19
C26589 VPWR.n38 0 0.00119f
C26590 VPWR.n39 0 0.0199f
C26591 VPWR.t147 0 0.0876f
C26592 VPWR.n40 0 0.0651f
C26593 VPWR.n41 0 0.051f
C26594 VPWR.n42 0 0.0199f
C26595 VPWR.n43 0 0.0973f
C26596 VPWR.n44 0 0.0809f
C26597 VPWR.t33 0 0.154f
C26598 VPWR.n45 0 0.41f
C26599 VPWR.t132 0 0.164f
C26600 VPWR.n46 0 0.769f
C26601 VPWR.n47 0 0.0596f
C26602 VPWR.n48 0 0.0445f
C26603 VPWR.n49 0 0.0372f
C26604 VPWR.n50 0 0.0256f
C26605 VPWR.t354 0 0.0671f
C26606 VPWR.n51 0 0.0607f
C26607 VPWR.n52 0 0.0851f
C26608 VPWR.n53 0 0.0376f
C26609 VPWR.n54 0 0.00119f
C26610 VPWR.n55 0 0.00162f
C26611 VPWR.n56 0 0.00215f
C26612 VPWR.n57 0 0.00113f
C26613 VPWR.n58 0 0.0736f
C26614 VPWR.n59 0 0.129f
C26615 VPWR.n60 0 0.13f
C26616 VPWR.n61 0 0.00302f
C26617 VPWR.t72 0 0.116f
C26618 VPWR.n62 0 0.322f
C26619 VPWR.n63 0 0.122f
C26620 VPWR.n64 0 0.0557f
C26621 VPWR.n65 0 0.0751f
C26622 VPWR.n66 0 0.0994f
C26623 VPWR.n67 0 0.0447f
C26624 VPWR.t268 0 0.0774f
C26625 VPWR.t141 0 0.0774f
C26626 VPWR.n68 0 0.0339f
C26627 VPWR.n69 0 0.0625f
C26628 VPWR.t269 0 0.0876f
C26629 VPWR.n70 0 0.113f
C26630 VPWR.n71 0 0.018f
C26631 VPWR.n72 0 0.0199f
C26632 VPWR.n73 0 0.0376f
C26633 VPWR.n74 0 0.0399f
C26634 VPWR.t227 0 0.0726f
C26635 VPWR.n75 0 0.0391f
C26636 VPWR.n76 0 0.267f
C26637 VPWR.n77 0 0.0405f
C26638 VPWR.n78 0 0.0619f
C26639 VPWR.n79 0 0.00164f
C26640 VPWR.n80 0 0.00281f
C26641 VPWR.n81 0 0.0086f
C26642 VPWR.n82 0 0.00529f
C26643 VPWR.n83 0 0.0555f
C26644 VPWR.n84 0 0.0572f
C26645 VPWR.t191 0 0.068f
C26646 VPWR.n85 0 0.0468f
C26647 VPWR.n86 0 0.0701f
C26648 VPWR.n87 0 0.0916f
C26649 VPWR.n88 0 0.0471f
C26650 VPWR.t270 0 0.116f
C26651 VPWR.n89 0 0.322f
C26652 VPWR.n90 0 0.00994f
C26653 VPWR.n91 0 0.0892f
C26654 VPWR.t60 0 0.0876f
C26655 VPWR.n92 0 0.104f
C26656 VPWR.n93 0 0.0397f
C26657 VPWR.n94 0 0.0556f
C26658 VPWR.n95 0 0.0664f
C26659 VPWR.n96 0 0.00259f
C26660 VPWR.n97 0 0.00421f
C26661 VPWR.n98 0 0.00378f
C26662 VPWR.n99 0 0.00162f
C26663 VPWR.n100 0 0.0014f
C26664 VPWR.n101 0 0.0014f
C26665 VPWR.n102 0 0.00208f
C26666 VPWR.n103 0 0.00344f
C26667 VPWR.n104 0 0.00248f
C26668 VPWR.n105 0 0.00329f
C26669 VPWR.n106 0 0.416f
C26670 VPWR.n107 0 0.00248f
C26671 VPWR.n108 0 0.00344f
C26672 VPWR.n109 0 0.00323f
C26673 VPWR.n110 0 0.00468f
C26674 VPWR.n111 0 0.00323f
C26675 VPWR.n112 0 0.00208f
C26676 VPWR.n114 0 0.00329f
C26677 VPWR.n115 0 0.00208f
C26678 VPWR.n116 0 0.00302f
C26679 VPWR.n117 0 0.00248f
C26680 VPWR.n118 0 0.00173f
C26681 VPWR.n119 0 0.0027f
C26682 VPWR.n120 0 0.00248f
C26683 VPWR.n121 0 0.00205f
C26684 VPWR.n122 0 0.00162f
C26685 VPWR.n123 0 0.00335f
C26686 VPWR.n124 0 0.00421f
C26687 VPWR.n125 0 0.00248f
C26688 VPWR.n126 0 7.56e-19
C26689 VPWR.n127 0 8.64e-19
C26690 VPWR.n128 0 0.00108f
C26691 VPWR.n129 0 0.00205f
C26692 VPWR.n130 0 0.00248f
C26693 VPWR.n131 0 0.0027f
C26694 VPWR.n132 0 0.00302f
C26695 VPWR.n133 0 0.00184f
C26696 VPWR.n134 0 9.72e-19
C26697 VPWR.n135 0 0.0014f
C26698 VPWR.n136 0 8.64e-19
C26699 VPWR.n137 0 0.00108f
C26700 VPWR.n138 0 0.00248f
C26701 VPWR.n139 0 0.00389f
C26702 VPWR.n140 0 0.00357f
C26703 VPWR.n141 0 0.00281f
C26704 VPWR.n142 0 0.00265f
C26705 VPWR.n143 0 0.00284f
C26706 VPWR.n144 0 0.00499f
C26707 VPWR.n145 0 0.00281f
C26708 VPWR.n146 0 0.00238f
C26709 VPWR.n147 0 0.00989f
C26710 VPWR.n148 0 0.00496f
C26711 VPWR.n149 0 0.0217f
C26712 VPWR.n151 0 0.00329f
C26713 VPWR.n152 0 0.00208f
C26714 VPWR.n153 0 0.00281f
C26715 VPWR.n154 0 0.00184f
C26716 VPWR.t388 0 0.0726f
C26717 VPWR.n155 0 0.245f
C26718 VPWR.n156 0 0.04f
C26719 VPWR.n157 0 0.0154f
C26720 VPWR.n158 0 0.306f
C26721 VPWR.n159 0 0.0818f
C26722 VPWR.n160 0 0.0715f
C26723 VPWR.t219 0 0.154f
C26724 VPWR.n161 0 0.521f
C26725 VPWR.n162 0 0.13f
C26726 VPWR.t96 0 0.0949f
C26727 VPWR.n163 0 0.0218f
C26728 VPWR.n164 0 0.128f
C26729 VPWR.n165 0 0.0176f
C26730 VPWR.n166 0 0.0483f
C26731 VPWR.n167 0 0.0894f
C26732 VPWR.n168 0 0.053f
C26733 VPWR.n169 0 0.156f
C26734 VPWR.n170 0 0.0856f
C26735 VPWR.n171 0 0.0452f
C26736 VPWR.n172 0 0.187f
C26737 VPWR.n173 0 0.158f
C26738 VPWR.n174 0 0.00119f
C26739 VPWR.n175 0 0.00119f
C26740 VPWR.n176 0 0.00344f
C26741 VPWR.n177 0 0.00248f
C26742 VPWR.n178 0 0.00329f
C26743 VPWR.n179 0 4.86f
C26744 VPWR.n181 0 0.00329f
C26745 VPWR.n182 0 0.00208f
C26746 VPWR.n183 0 0.00259f
C26747 VPWR.t216 0 0.15f
C26748 VPWR.n184 0 0.475f
C26749 VPWR.n185 0 0.165f
C26750 VPWR.t118 0 0.116f
C26751 VPWR.n186 0 0.325f
C26752 VPWR.n187 0 0.0848f
C26753 VPWR.n188 0 0.00352f
C26754 VPWR.n189 0 0.00994f
C26755 VPWR.t306 0 0.0716f
C26756 VPWR.n190 0 0.0306f
C26757 VPWR.n191 0 0.197f
C26758 VPWR.t202 0 0.0407f
C26759 VPWR.n192 0 0.0607f
C26760 VPWR.t161 0 0.0774f
C26761 VPWR.t264 0 0.0774f
C26762 VPWR.n193 0 0.501f
C26763 VPWR.t325 0 0.0417f
C26764 VPWR.t302 0 0.0417f
C26765 VPWR.n194 0 0.383f
C26766 VPWR.n195 0 0.0384f
C26767 VPWR.n196 0 0.0421f
C26768 VPWR.n197 0 0.00994f
C26769 VPWR.n198 0 0.00595f
C26770 VPWR.n199 0 0.05f
C26771 VPWR.n200 0 0.018f
C26772 VPWR.n201 0 0.0199f
C26773 VPWR.n202 0 0.00578f
C26774 VPWR.n203 0 0.189f
C26775 VPWR.n204 0 0.018f
C26776 VPWR.n205 0 0.0118f
C26777 VPWR.n206 0 0.0143f
C26778 VPWR.n207 0 0.125f
C26779 VPWR.n208 0 0.018f
C26780 VPWR.n209 0 0.0199f
C26781 VPWR.n210 0 0.0125f
C26782 VPWR.n211 0 0.115f
C26783 VPWR.t289 0 0.0592f
C26784 VPWR.n212 0 0.0237f
C26785 VPWR.n213 0 0.0906f
C26786 VPWR.n214 0 0.0192f
C26787 VPWR.n215 0 0.115f
C26788 VPWR.n216 0 0.16f
C26789 VPWR.n217 0 0.0246f
C26790 VPWR.n218 0 0.0887f
C26791 VPWR.n219 0 0.0784f
C26792 VPWR.n220 0 0.0135f
C26793 VPWR.n221 0 0.0387f
C26794 VPWR.n222 0 0.0359f
C26795 VPWR.n223 0 0.00184f
C26796 VPWR.t319 0 0.073f
C26797 VPWR.n224 0 0.207f
C26798 VPWR.n225 0 0.0645f
C26799 VPWR.n226 0 0.0387f
C26800 VPWR.n227 0 0.0386f
C26801 VPWR.n228 0 0.0534f
C26802 VPWR.n229 0 0.00497f
C26803 VPWR.n230 0 0.00344f
C26804 VPWR.n231 0 0.00248f
C26805 VPWR.n232 0 0.00329f
C26806 VPWR.n233 0 0.00208f
C26807 VPWR.n234 0 0.00302f
C26808 VPWR.n235 0 0.00248f
C26809 VPWR.n236 0 0.00173f
C26810 VPWR.n237 0 0.014f
C26811 VPWR.n238 0 0.00194f
C26812 VPWR.n239 0 0.0013f
C26813 VPWR.n240 0 0.00108f
C26814 VPWR.n241 0 0.00194f
C26815 VPWR.n242 0 0.00173f
C26816 VPWR.n243 0 0.0014f
C26817 VPWR.n244 0 8.64e-19
C26818 VPWR.n245 0 0.00108f
C26819 VPWR.n246 0 0.00248f
C26820 VPWR.n247 0 0.00378f
C26821 VPWR.n248 0 0.00194f
C26822 VPWR.n249 0 0.00173f
C26823 VPWR.n250 0 0.0027f
C26824 VPWR.n251 0 0.00119f
C26825 VPWR.n252 0 0.00486f
C26826 VPWR.n253 0 0.00389f
C26827 VPWR.n254 0 0.00173f
C26828 VPWR.n255 0 0.0027f
C26829 VPWR.t32 0 0.0876f
C26830 VPWR.n256 0 0.00482f
C26831 VPWR.n257 0 0.0462f
C26832 VPWR.n258 0 0.0261f
C26833 VPWR.n259 0 0.125f
C26834 VPWR.n260 0 0.00119f
C26835 VPWR.n261 0 0.0428f
C26836 VPWR.n262 0 0.028f
C26837 VPWR.t21 0 0.116f
C26838 VPWR.n263 0 0.00467f
C26839 VPWR.t149 0 0.0774f
C26840 VPWR.n264 0 0.114f
C26841 VPWR.n265 0 0.0809f
C26842 VPWR.t261 0 0.0417f
C26843 VPWR.n266 0 0.0208f
C26844 VPWR.t234 0 0.0417f
C26845 VPWR.n267 0 0.383f
C26846 VPWR.t142 0 0.0774f
C26847 VPWR.t365 0 0.0774f
C26848 VPWR.n268 0 0.501f
C26849 VPWR.n269 0 0.0299f
C26850 VPWR.n270 0 0.0394f
C26851 VPWR.n271 0 0.00429f
C26852 VPWR.n272 0 0.0199f
C26853 VPWR.n273 0 0.018f
C26854 VPWR.n274 0 0.0275f
C26855 VPWR.n275 0 0.339f
C26856 VPWR.n276 0 0.432f
C26857 VPWR.n277 0 0.0885f
C26858 VPWR.n278 0 0.0276f
C26859 VPWR.n279 0 0.0118f
C26860 VPWR.n280 0 0.00597f
C26861 VPWR.n281 0 0.0199f
C26862 VPWR.n282 0 0.0199f
C26863 VPWR.n283 0 0.018f
C26864 VPWR.n284 0 0.0059f
C26865 VPWR.n285 0 0.0753f
C26866 VPWR.n286 0 0.0118f
C26867 VPWR.n287 0 0.0671f
C26868 VPWR.n288 0 0.0199f
C26869 VPWR.n289 0 0.0636f
C26870 VPWR.n290 0 0.0199f
C26871 VPWR.n291 0 0.0709f
C26872 VPWR.n292 0 0.018f
C26873 VPWR.n293 0 0.00983f
C26874 VPWR.n294 0 0.00184f
C26875 VPWR.n295 0 0.00881f
C26876 VPWR.n296 0 0.00496f
C26877 VPWR.n297 0 0.381f
C26878 VPWR.n298 0 0.00329f
C26879 VPWR.n299 0 0.0027f
C26880 VPWR.n300 0 0.00497f
C26881 VPWR.n301 0 0.00367f
C26882 VPWR.n302 0 0.00281f
C26883 VPWR.n303 0 0.00162f
C26884 VPWR.n304 0 0.00205f
C26885 VPWR.n305 0 0.00443f
C26886 VPWR.n306 0 0.00302f
C26887 VPWR.n307 0 0.00443f
C26888 VPWR.n308 0 0.00281f
C26889 VPWR.n309 0 8.64e-19
C26890 VPWR.n310 0 0.00238f
C26891 VPWR.t380 0 0.068f
C26892 VPWR.n311 0 0.0701f
C26893 VPWR.n312 0 0.0525f
C26894 VPWR.n313 0 0.0617f
C26895 VPWR.n314 0 0.0856f
C26896 VPWR.n315 0 0.0749f
C26897 VPWR.t75 0 0.0876f
C26898 VPWR.n316 0 0.109f
C26899 VPWR.t391 0 0.068f
C26900 VPWR.n317 0 0.0731f
C26901 VPWR.n318 0 0.0014f
C26902 VPWR.n319 0 0.0014f
C26903 VPWR.n320 0 0.00329f
C26904 VPWR.n321 0 0.00208f
C26905 VPWR.n322 0 0.0605f
C26906 VPWR.n323 0 0.37f
C26907 VPWR.n324 0 0.331f
C26908 VPWR.n325 0 0.00248f
C26909 VPWR.n326 0 0.00344f
C26910 VPWR.n327 0 0.00468f
C26911 VPWR.n328 0 0.00323f
C26912 VPWR.n329 0 0.00208f
C26913 VPWR.n331 0 0.00329f
C26914 VPWR.n332 0 0.00208f
C26915 VPWR.n333 0 0.00481f
C26916 VPWR.n334 0 0.00329f
C26917 VPWR.n335 0 0.00208f
C26918 VPWR.n336 0 0.00302f
C26919 VPWR.n337 0 0.00248f
C26920 VPWR.n338 0 0.00173f
C26921 VPWR.n339 0 0.00306f
C26922 VPWR.n340 0 0.00259f
C26923 VPWR.n341 0 0.0027f
C26924 VPWR.n342 0 0.00248f
C26925 VPWR.n343 0 0.00205f
C26926 VPWR.n344 0 0.00744f
C26927 VPWR.n345 0 0.00266f
C26928 VPWR.n346 0 0.00259f
C26929 VPWR.n347 0 0.00302f
C26930 VPWR.n348 0 0.00162f
C26931 VPWR.n349 0 0.0014f
C26932 VPWR.n350 0 0.0671f
C26933 VPWR.t53 0 0.068f
C26934 VPWR.n351 0 0.0893f
C26935 VPWR.n352 0 0.0391f
C26936 VPWR.n353 0 0.0844f
C26937 VPWR.t257 0 0.068f
C26938 VPWR.n354 0 0.0701f
C26939 VPWR.n355 0 0.0199f
C26940 VPWR.n356 0 0.0118f
C26941 VPWR.n357 0 0.0773f
C26942 VPWR.n358 0 0.0199f
C26943 VPWR.t54 0 0.068f
C26944 VPWR.n359 0 0.0535f
C26945 VPWR.n360 0 0.0199f
C26946 VPWR.t7 0 0.068f
C26947 VPWR.n361 0 0.0855f
C26948 VPWR.n362 0 0.0457f
C26949 VPWR.n363 0 0.0199f
C26950 VPWR.t37 0 0.068f
C26951 VPWR.n364 0 0.0865f
C26952 VPWR.n365 0 0.0199f
C26953 VPWR.n366 0 0.00609f
C26954 VPWR.n367 0 0.0118f
C26955 VPWR.t332 0 0.0876f
C26956 VPWR.n368 0 0.113f
C26957 VPWR.t67 0 0.0718f
C26958 VPWR.n369 0 0.208f
C26959 VPWR.n370 0 0.0963f
C26960 VPWR.t229 0 0.068f
C26961 VPWR.t94 0 0.0711f
C26962 VPWR.n371 0 0.195f
C26963 VPWR.n372 0 0.0877f
C26964 VPWR.n373 0 0.0391f
C26965 VPWR.n374 0 0.0701f
C26966 VPWR.n375 0 0.0118f
C26967 VPWR.n376 0 0.0199f
C26968 VPWR.n377 0 0.018f
C26969 VPWR.n378 0 0.00994f
C26970 VPWR.n379 0 0.049f
C26971 VPWR.n380 0 0.00529f
C26972 VPWR.n381 0 0.0199f
C26973 VPWR.n382 0 0.018f
C26974 VPWR.n383 0 0.00429f
C26975 VPWR.n384 0 0.0569f
C26976 VPWR.n385 0 0.00994f
C26977 VPWR.n386 0 0.0198f
C26978 VPWR.n387 0 0.0107f
C26979 VPWR.n388 0 0.125f
C26980 VPWR.n389 0 0.128f
C26981 VPWR.n390 0 0.106f
C26982 VPWR.n391 0 0.0173f
C26983 VPWR.n392 0 0.0107f
C26984 VPWR.n393 0 0.0118f
C26985 VPWR.n394 0 0.0657f
C26986 VPWR.n395 0 0.0934f
C26987 VPWR.n396 0 0.0443f
C26988 VPWR.n397 0 0.0199f
C26989 VPWR.n398 0 0.018f
C26990 VPWR.n399 0 0.0484f
C26991 VPWR.n400 0 0.0324f
C26992 VPWR.n401 0 0.0605f
C26993 VPWR.n402 0 0.00429f
C26994 VPWR.n403 0 0.0199f
C26995 VPWR.n404 0 0.018f
C26996 VPWR.n405 0 0.0118f
C26997 VPWR.n406 0 0.0199f
C26998 VPWR.n407 0 0.0649f
C26999 VPWR.n408 0 0.0408f
C27000 VPWR.n409 0 0.0939f
C27001 VPWR.n410 0 0.0475f
C27002 VPWR.n411 0 0.0173f
C27003 VPWR.n412 0 0.0107f
C27004 VPWR.n413 0 0.0619f
C27005 VPWR.n414 0 0.0118f
C27006 VPWR.n415 0 0.0199f
C27007 VPWR.n416 0 0.0199f
C27008 VPWR.n417 0 0.051f
C27009 VPWR.n418 0 0.0785f
C27010 VPWR.n419 0 0.049f
C27011 VPWR.n420 0 0.0115f
C27012 VPWR.n421 0 0.0199f
C27013 VPWR.n422 0 0.018f
C27014 VPWR.n423 0 0.00994f
C27015 VPWR.n424 0 0.00706f
C27016 VPWR.n425 0 0.0664f
C27017 VPWR.n426 0 0.0536f
C27018 VPWR.n427 0 0.0391f
C27019 VPWR.n428 0 0.018f
C27020 VPWR.n429 0 0.00994f
C27021 VPWR.n430 0 0.0478f
C27022 VPWR.n431 0 0.0505f
C27023 VPWR.n432 0 0.0117f
C27024 VPWR.n433 0 0.0199f
C27025 VPWR.n434 0 0.0199f
C27026 VPWR.n435 0 0.018f
C27027 VPWR.n436 0 0.0712f
C27028 VPWR.n437 0 0.025f
C27029 VPWR.n438 0 0.0118f
C27030 VPWR.n439 0 0.0671f
C27031 VPWR.n440 0 0.0199f
C27032 VPWR.n441 0 0.0393f
C27033 VPWR.n442 0 0.0199f
C27034 VPWR.n443 0 0.0271f
C27035 VPWR.n444 0 0.0199f
C27036 VPWR.n445 0 0.0575f
C27037 VPWR.n446 0 0.0199f
C27038 VPWR.n447 0 0.0197f
C27039 VPWR.n448 0 0.0199f
C27040 VPWR.n449 0 0.0199f
C27041 VPWR.n450 0 0.018f
C27042 VPWR.n451 0 0.00491f
C27043 VPWR.n452 0 0.0753f
C27044 VPWR.n453 0 0.0118f
C27045 VPWR.n454 0 0.0671f
C27046 VPWR.n455 0 0.0199f
C27047 VPWR.t195 0 0.068f
C27048 VPWR.n456 0 0.045f
C27049 VPWR.n457 0 0.09f
C27050 VPWR.n458 0 0.0391f
C27051 VPWR.n459 0 0.0196f
C27052 VPWR.n460 0 0.00994f
C27053 VPWR.n461 0 0.00482f
C27054 VPWR.n462 0 0.00184f
C27055 VPWR.n463 0 0.014f
C27056 VPWR.n464 0 0.00292f
C27057 VPWR.n465 0 0.00259f
C27058 VPWR.n466 0 0.00259f
C27059 VPWR.n467 0 0.0014f
C27060 VPWR.n468 0 0.00162f
C27061 VPWR.n469 0 0.00335f
C27062 VPWR.n470 0 0.00421f
C27063 VPWR.n471 0 0.00248f
C27064 VPWR.n472 0 7.56e-19
C27065 VPWR.n473 0 8.64e-19
C27066 VPWR.n474 0 0.00108f
C27067 VPWR.n475 0 0.00205f
C27068 VPWR.n476 0 0.00248f
C27069 VPWR.n477 0 0.0027f
C27070 VPWR.n478 0 0.00302f
C27071 VPWR.n479 0 0.00184f
C27072 VPWR.n480 0 9.72e-19
C27073 VPWR.n481 0 0.0014f
C27074 VPWR.n482 0 8.64e-19
C27075 VPWR.n483 0 0.00108f
C27076 VPWR.n484 0 0.00248f
C27077 VPWR.n485 0 0.00389f
C27078 VPWR.n486 0 0.00357f
C27079 VPWR.n487 0 0.00281f
C27080 VPWR.n488 0 0.0575f
C27081 VPWR.n489 0 0.0715f
C27082 VPWR.t348 0 0.0973f
C27083 VPWR.n490 0 0.219f
C27084 VPWR.n491 0 0.113f
C27085 VPWR.n492 0 0.0623f
C27086 VPWR.t367 0 0.0726f
C27087 VPWR.n493 0 0.0391f
C27088 VPWR.n494 0 0.267f
C27089 VPWR.n495 0 0.0391f
C27090 VPWR.t210 0 0.107f
C27091 VPWR.n496 0 0.0612f
C27092 VPWR.n497 0 0.00994f
C27093 VPWR.t265 0 0.068f
C27094 VPWR.n498 0 0.0701f
C27095 VPWR.t188 0 0.069f
C27096 VPWR.n499 0 0.102f
C27097 VPWR.t353 0 0.116f
C27098 VPWR.n500 0 0.322f
C27099 VPWR.t162 0 0.0737f
C27100 VPWR.n501 0 0.3f
C27101 VPWR.n502 0 0.241f
C27102 VPWR.t370 0 0.0774f
C27103 VPWR.n503 0 0.29f
C27104 VPWR.n504 0 0.00417f
C27105 VPWR.n505 0 0.00113f
C27106 VPWR.n506 0 0.00215f
C27107 VPWR.n507 0 0.00184f
C27108 VPWR.n508 0 0.00259f
C27109 VPWR.n509 0 0.00119f
C27110 VPWR.n510 0 0.00421f
C27111 VPWR.n511 0 0.00248f
C27112 VPWR.n512 0 5.4e-19
C27113 VPWR.n513 0 0.00119f
C27114 VPWR.n514 0 0.00302f
C27115 VPWR.n515 0 0.00248f
C27116 VPWR.n516 0 5.4e-19
C27117 VPWR.n517 0 0.00259f
C27118 VPWR.n518 0 8.64e-19
C27119 VPWR.n519 0 0.00227f
C27120 VPWR.n520 0 0.00248f
C27121 VPWR.n521 0 0.00248f
C27122 VPWR.n522 0 0.00194f
C27123 VPWR.n523 0 0.00184f
C27124 VPWR.n524 0 0.00259f
C27125 VPWR.n525 0 0.00119f
C27126 VPWR.n526 0 0.00344f
C27127 VPWR.n527 0 0.00248f
C27128 VPWR.n528 0 0.00329f
C27129 VPWR.n529 0 0.00208f
C27130 VPWR.n530 0 0.00498f
C27131 VPWR.n531 0 0.00891f
C27132 VPWR.n532 0 0.0201f
C27133 VPWR.n533 0 0.0181f
C27134 VPWR.n534 0 0.00994f
C27135 VPWR.n535 0 0.0652f
C27136 VPWR.n536 0 0.00467f
C27137 VPWR.n537 0 0.018f
C27138 VPWR.n538 0 0.0118f
C27139 VPWR.n539 0 0.0998f
C27140 VPWR.n540 0 0.00467f
C27141 VPWR.n541 0 0.00994f
C27142 VPWR.n542 0 0.0267f
C27143 VPWR.n543 0 0.00994f
C27144 VPWR.n544 0 0.0429f
C27145 VPWR.n545 0 0.0958f
C27146 VPWR.n546 0 0.0954f
C27147 VPWR.n547 0 0.018f
C27148 VPWR.n548 0 0.0199f
C27149 VPWR.n549 0 0.0305f
C27150 VPWR.n550 0 0.0118f
C27151 VPWR.n551 0 0.0118f
C27152 VPWR.n552 0 0.0199f
C27153 VPWR.n553 0 0.018f
C27154 VPWR.n554 0 0.0381f
C27155 VPWR.n555 0 0.0967f
C27156 VPWR.n556 0 0.0629f
C27157 VPWR.n557 0 0.0485f
C27158 VPWR.n558 0 0.00994f
C27159 VPWR.n559 0 0.0118f
C27160 VPWR.n560 0 0.0199f
C27161 VPWR.n561 0 0.018f
C27162 VPWR.n562 0 0.0391f
C27163 VPWR.n563 0 0.0696f
C27164 VPWR.n564 0 0.0709f
C27165 VPWR.n565 0 0.0544f
C27166 VPWR.t209 0 0.0724f
C27167 VPWR.n566 0 0.207f
C27168 VPWR.n567 0 0.079f
C27169 VPWR.n568 0 0.0311f
C27170 VPWR.n569 0 0.0429f
C27171 VPWR.n570 0 0.0231f
C27172 VPWR.n571 0 0.0107f
C27173 VPWR.n572 0 0.00918f
C27174 VPWR.n573 0 0.0659f
C27175 VPWR.n574 0 0.0108f
C27176 VPWR.n575 0 0.0172f
C27177 VPWR.n576 0 0.0117f
C27178 VPWR.n577 0 0.041f
C27179 VPWR.n578 0 0.185f
C27180 VPWR.n579 0 0.0386f
C27181 VPWR.n580 0 0.0181f
C27182 VPWR.n581 0 0.0199f
C27183 VPWR.n582 0 0.0199f
C27184 VPWR.n583 0 0.0118f
C27185 VPWR.n584 0 0.0522f
C27186 VPWR.n585 0 0.0535f
C27187 VPWR.n586 0 0.00994f
C27188 VPWR.n587 0 0.00994f
C27189 VPWR.n588 0 0.00994f
C27190 VPWR.n589 0 0.0426f
C27191 VPWR.n590 0 0.00604f
C27192 VPWR.n591 0 0.018f
C27193 VPWR.n592 0 0.0199f
C27194 VPWR.n593 0 0.0199f
C27195 VPWR.t228 0 0.0876f
C27196 VPWR.n594 0 0.0975f
C27197 VPWR.n595 0 0.149f
C27198 VPWR.n596 0 0.13f
C27199 VPWR.n597 0 0.0125f
C27200 VPWR.n598 0 0.0198f
C27201 VPWR.n599 0 0.018f
C27202 VPWR.n600 0 0.0199f
C27203 VPWR.n601 0 0.0118f
C27204 VPWR.n602 0 0.0758f
C27205 VPWR.n603 0 0.00521f
C27206 VPWR.n604 0 0.018f
C27207 VPWR.n605 0 0.0117f
C27208 VPWR.n606 0 0.0514f
C27209 VPWR.n607 0 0.0528f
C27210 VPWR.n608 0 0.0181f
C27211 VPWR.n609 0 0.0199f
C27212 VPWR.n610 0 0.0199f
C27213 VPWR.t256 0 0.068f
C27214 VPWR.n611 0 0.0865f
C27215 VPWR.n612 0 0.0391f
C27216 VPWR.n613 0 0.0751f
C27217 VPWR.n614 0 0.0654f
C27218 VPWR.n615 0 0.0118f
C27219 VPWR.n616 0 0.00258f
C27220 VPWR.n617 0 0.00291f
C27221 VPWR.n618 0 0.00498f
C27222 VPWR.n619 0 0.00281f
C27223 VPWR.n620 0 0.00313f
C27224 VPWR.n621 0 0.00989f
C27225 VPWR.n622 0 0.00496f
C27226 VPWR.n623 0 0.0217f
C27227 VPWR.n624 0 0.00323f
C27228 VPWR.n625 0 0.00248f
C27229 VPWR.n626 0 0.00344f
C27230 VPWR.n627 0 0.00208f
C27231 VPWR.n629 0 0.381f
C27232 VPWR.n630 0 0.381f
C27233 VPWR.n631 0 0.00248f
C27234 VPWR.n632 0 0.00344f
C27235 VPWR.n633 0 0.00468f
C27236 VPWR.n634 0 0.00323f
C27237 VPWR.n635 0 0.00208f
C27238 VPWR.n637 0 0.00323f
C27239 VPWR.n638 0 0.00248f
C27240 VPWR.n639 0 0.00344f
C27241 VPWR.n640 0 0.00208f
C27242 VPWR.n642 0 0.00329f
C27243 VPWR.n643 0 0.00208f
C27244 VPWR.n644 0 0.00281f
C27245 VPWR.n645 0 0.00258f
C27246 VPWR.t340 0 0.068f
C27247 VPWR.n646 0 0.00482f
C27248 VPWR.n647 0 0.013f
C27249 VPWR.n648 0 0.0587f
C27250 VPWR.n649 0 0.00357f
C27251 VPWR.n650 0 0.00389f
C27252 VPWR.n651 0 0.00248f
C27253 VPWR.n652 0 0.00108f
C27254 VPWR.n653 0 0.00302f
C27255 VPWR.n654 0 0.00248f
C27256 VPWR.n655 0 0.00173f
C27257 VPWR.n656 0 8.64e-19
C27258 VPWR.n657 0 0.0014f
C27259 VPWR.n658 0 9.72e-19
C27260 VPWR.n659 0 0.00184f
C27261 VPWR.n660 0 0.00302f
C27262 VPWR.n661 0 0.0027f
C27263 VPWR.n662 0 0.00248f
C27264 VPWR.n663 0 0.00205f
C27265 VPWR.n664 0 0.0027f
C27266 VPWR.n665 0 0.00248f
C27267 VPWR.n666 0 0.00205f
C27268 VPWR.n667 0 0.00162f
C27269 VPWR.n668 0 0.00335f
C27270 VPWR.n669 0 0.00421f
C27271 VPWR.n670 0 0.00248f
C27272 VPWR.n671 0 7.56e-19
C27273 VPWR.n672 0 8.64e-19
C27274 VPWR.n673 0 0.00108f
C27275 VPWR.n674 0 0.00259f
C27276 VPWR.n675 0 0.00162f
C27277 VPWR.n676 0 0.00378f
C27278 VPWR.n677 0 0.0202f
C27279 VPWR.n678 0 0.0427f
C27280 VPWR.n679 0 2.35e-19
C27281 VPWR.n680 0 0.0759f
C27282 VPWR.n681 0 0.0952f
C27283 VPWR.n682 0 0.00983f
C27284 VPWR.n683 0 0.00119f
C27285 VPWR.n684 0 0.00119f
C27286 VPWR.n685 0 0.00344f
C27287 VPWR.n686 0 0.00248f
C27288 VPWR.n687 0 0.00329f
C27289 VPWR.n688 0 0.00214f
C27290 VPWR.n689 0 0.00237f
C27291 VPWR.n690 0 3.59f
C27292 VPWR.n691 0 0.00323f
C27293 VPWR.n692 0 0.00344f
C27294 VPWR.n693 0 0.00208f
C27295 VPWR.n694 0 0.00214f
C27296 VPWR.n695 0 0.00344f
C27297 VPWR.n696 0 0.00468f
C27298 VPWR.n697 0 0.00323f
C27299 VPWR.n698 0 0.00208f
C27300 VPWR.n700 0 0.00259f
C27301 VPWR.n701 0 0.061f
C27302 VPWR.t150 0 0.116f
C27303 VPWR.n702 0 0.0196f
C27304 VPWR.t192 0 0.0775f
C27305 VPWR.n703 0 0.01f
C27306 VPWR.t317 0 0.0417f
C27307 VPWR.t291 0 0.0417f
C27308 VPWR.n704 0 0.384f
C27309 VPWR.n705 0 0.019f
C27310 VPWR.n706 0 0.0246f
C27311 VPWR.n707 0 0.00482f
C27312 VPWR.n708 0 0.303f
C27313 VPWR.n709 0 0.322f
C27314 VPWR.n710 0 0.0953f
C27315 VPWR.n711 0 0.018f
C27316 VPWR.n712 0 0.0541f
C27317 VPWR.n713 0 0.0199f
C27318 VPWR.n714 0 0.13f
C27319 VPWR.n715 0 0.0199f
C27320 VPWR.t220 0 0.069f
C27321 VPWR.n716 0 0.0381f
C27322 VPWR.n717 0 0.102f
C27323 VPWR.n718 0 0.0305f
C27324 VPWR.n719 0 0.0118f
C27325 VPWR.n720 0 0.018f
C27326 VPWR.n721 0 0.0199f
C27327 VPWR.n722 0 0.0118f
C27328 VPWR.n723 0 0.0856f
C27329 VPWR.n724 0 0.0668f
C27330 VPWR.n725 0 0.018f
C27331 VPWR.n726 0 0.00394f
C27332 VPWR.n727 0 0.0199f
C27333 VPWR.n728 0 0.0329f
C27334 VPWR.n729 0 0.0199f
C27335 VPWR.n730 0 0.00482f
C27336 VPWR.n731 0 0.0265f
C27337 VPWR.n732 0 0.162f
C27338 VPWR.n733 0 0.0265f
C27339 VPWR.n734 0 0.0184f
C27340 VPWR.n735 0 0.00552f
C27341 VPWR.n736 0 0.049f
C27342 VPWR.n737 0 0.018f
C27343 VPWR.t221 0 0.068f
C27344 VPWR.n738 0 0.0818f
C27345 VPWR.n739 0 0.049f
C27346 VPWR.n740 0 0.0199f
C27347 VPWR.n741 0 0.0561f
C27348 VPWR.n742 0 0.0563f
C27349 VPWR.n743 0 0.0186f
C27350 VPWR.n744 0 0.00994f
C27351 VPWR.n745 0 0.00184f
C27352 VPWR.n746 0 0.015f
C27353 VPWR.n747 0 0.0156f
C27354 VPWR.n748 0 7.56e-19
C27355 VPWR.n749 0 0.00184f
C27356 VPWR.n750 0 0.0376f
C27357 VPWR.n751 0 0.0385f
C27358 VPWR.n752 0 0.0398f
C27359 VPWR.n753 0 0.0627f
C27360 VPWR.n754 0 0.0027f
C27361 VPWR.n755 0 0.00367f
C27362 VPWR.n756 0 0.00281f
C27363 VPWR.n757 0 0.00859f
C27364 VPWR.t26 0 0.068f
C27365 VPWR.n758 0 0.0701f
C27366 VPWR.n759 0 0.0391f
C27367 VPWR.n760 0 0.0716f
C27368 VPWR.t328 0 0.068f
C27369 VPWR.n761 0 0.0701f
C27370 VPWR.n762 0 0.0391f
C27371 VPWR.n763 0 0.121f
C27372 VPWR.n764 0 0.123f
C27373 VPWR.n765 0 0.0522f
C27374 VPWR.n766 0 0.0535f
C27375 VPWR.n767 0 0.141f
C27376 VPWR.n768 0 0.0246f
C27377 VPWR.t236 0 0.107f
C27378 VPWR.n769 0 0.00305f
C27379 VPWR.n770 0 0.00259f
C27380 VPWR.n771 0 0.0275f
C27381 VPWR.n772 0 0.00275f
C27382 VPWR.n773 0 0.00525f
C27383 VPWR.n774 0 0.00162f
C27384 VPWR.n775 0 0.0014f
C27385 VPWR.n776 0 0.0014f
C27386 VPWR.n777 0 0.00484f
C27387 VPWR.n778 0 0.00214f
C27388 VPWR.n779 0 0.00214f
C27389 VPWR.n780 0 0.00344f
C27390 VPWR.n781 0 0.00468f
C27391 VPWR.n782 0 0.00323f
C27392 VPWR.n783 0 0.00208f
C27393 VPWR.n785 0 0.00302f
C27394 VPWR.n786 0 0.00248f
C27395 VPWR.n787 0 0.00173f
C27396 VPWR.n788 0 0.0027f
C27397 VPWR.n789 0 0.00248f
C27398 VPWR.n790 0 0.00205f
C27399 VPWR.n791 0 0.00162f
C27400 VPWR.n792 0 0.00335f
C27401 VPWR.n793 0 0.00421f
C27402 VPWR.n794 0 0.00248f
C27403 VPWR.n795 0 7.56e-19
C27404 VPWR.n796 0 8.64e-19
C27405 VPWR.n797 0 0.00108f
C27406 VPWR.n798 0 0.00205f
C27407 VPWR.n799 0 0.00248f
C27408 VPWR.n800 0 0.0027f
C27409 VPWR.n801 0 0.00302f
C27410 VPWR.n802 0 0.00184f
C27411 VPWR.n803 0 9.72e-19
C27412 VPWR.n804 0 0.0014f
C27413 VPWR.n805 0 8.64e-19
C27414 VPWR.n806 0 0.00108f
C27415 VPWR.n807 0 0.00248f
C27416 VPWR.n808 0 0.00389f
C27417 VPWR.n809 0 0.00357f
C27418 VPWR.n810 0 0.00281f
C27419 VPWR.n811 0 0.0449f
C27420 VPWR.n812 0 0.0655f
C27421 VPWR.n813 0 0.0617f
C27422 VPWR.t218 0 0.0876f
C27423 VPWR.n814 0 0.0631f
C27424 VPWR.n815 0 0.0181f
C27425 VPWR.t124 0 0.068f
C27426 VPWR.t99 0 0.068f
C27427 VPWR.n816 0 0.0981f
C27428 VPWR.n817 0 0.0391f
C27429 VPWR.n818 0 0.0815f
C27430 VPWR.t164 0 0.0774f
C27431 VPWR.t271 0 0.116f
C27432 VPWR.n819 0 0.432f
C27433 VPWR.n820 0 0.338f
C27434 VPWR.n821 0 0.114f
C27435 VPWR.n822 0 0.0634f
C27436 VPWR.n823 0 0.0391f
C27437 VPWR.n824 0 0.0173f
C27438 VPWR.t178 0 0.107f
C27439 VPWR.n825 0 0.0526f
C27440 VPWR.n826 0 0.00994f
C27441 VPWR.n827 0 0.0118f
C27442 VPWR.n828 0 0.00313f
C27443 VPWR.n829 0 0.00397f
C27444 VPWR.n830 0 0.00151f
C27445 VPWR.n831 0 0.011f
C27446 VPWR.n832 0 0.00162f
C27447 VPWR.n833 0 0.00119f
C27448 VPWR.n834 0 0.00184f
C27449 VPWR.n835 0 0.00259f
C27450 VPWR.n836 0 0.00119f
C27451 VPWR.n837 0 0.00421f
C27452 VPWR.n838 0 0.00248f
C27453 VPWR.n839 0 5.4e-19
C27454 VPWR.n840 0 0.00119f
C27455 VPWR.n841 0 0.00302f
C27456 VPWR.n842 0 0.00248f
C27457 VPWR.n843 0 5.4e-19
C27458 VPWR.n844 0 0.00259f
C27459 VPWR.n845 0 8.64e-19
C27460 VPWR.n846 0 0.00227f
C27461 VPWR.n847 0 0.00248f
C27462 VPWR.n848 0 0.00248f
C27463 VPWR.n849 0 0.00194f
C27464 VPWR.n850 0 0.00184f
C27465 VPWR.n851 0 0.00259f
C27466 VPWR.n852 0 0.00119f
C27467 VPWR.n853 0 0.00484f
C27468 VPWR.n854 0 0.00126f
C27469 VPWR.n855 0 0.00208f
C27470 VPWR.n856 0 1.45e-19
C27471 VPWR.n857 0 0.00891f
C27472 VPWR.n858 0 0.00616f
C27473 VPWR.t297 0 0.068f
C27474 VPWR.n859 0 0.0266f
C27475 VPWR.n860 0 0.0649f
C27476 VPWR.n861 0 0.0399f
C27477 VPWR.n862 0 0.0159f
C27478 VPWR.n863 0 0.0873f
C27479 VPWR.n864 0 0.0199f
C27480 VPWR.n865 0 0.0118f
C27481 VPWR.n866 0 0.0618f
C27482 VPWR.n867 0 0.0869f
C27483 VPWR.n868 0 0.00283f
C27484 VPWR.n869 0 0.00994f
C27485 VPWR.n870 0 0.0107f
C27486 VPWR.n871 0 0.00994f
C27487 VPWR.n872 0 0.0626f
C27488 VPWR.n873 0 0.041f
C27489 VPWR.n874 0 0.185f
C27490 VPWR.t203 0 0.0726f
C27491 VPWR.n875 0 0.267f
C27492 VPWR.n876 0 0.0255f
C27493 VPWR.n877 0 0.0199f
C27494 VPWR.n878 0 0.0199f
C27495 VPWR.n879 0 0.0118f
C27496 VPWR.n880 0 0.0522f
C27497 VPWR.n881 0 0.0487f
C27498 VPWR.n882 0 0.062f
C27499 VPWR.n883 0 0.00994f
C27500 VPWR.n884 0 0.018f
C27501 VPWR.n885 0 0.0118f
C27502 VPWR.n886 0 0.00994f
C27503 VPWR.n887 0 0.00655f
C27504 VPWR.n888 0 0.0395f
C27505 VPWR.n889 0 0.018f
C27506 VPWR.n890 0 0.0601f
C27507 VPWR.n891 0 0.0199f
C27508 VPWR.n892 0 0.0057f
C27509 VPWR.n893 0 0.0199f
C27510 VPWR.n894 0 0.00593f
C27511 VPWR.n895 0 0.0125f
C27512 VPWR.n896 0 0.057f
C27513 VPWR.n897 0 0.0491f
C27514 VPWR.n898 0 0.0107f
C27515 VPWR.n899 0 0.0553f
C27516 VPWR.n900 0 0.0173f
C27517 VPWR.n901 0 0.0199f
C27518 VPWR.n902 0 0.0199f
C27519 VPWR.n903 0 0.0118f
C27520 VPWR.n904 0 0.0711f
C27521 VPWR.n905 0 0.00655f
C27522 VPWR.n906 0 0.018f
C27523 VPWR.n907 0 0.00704f
C27524 VPWR.n908 0 0.0199f
C27525 VPWR.n909 0 0.0057f
C27526 VPWR.n910 0 0.0199f
C27527 VPWR.n911 0 0.0576f
C27528 VPWR.n912 0 0.0199f
C27529 VPWR.n913 0 0.0117f
C27530 VPWR.n914 0 0.00537f
C27531 VPWR.n915 0 0.049f
C27532 VPWR.n916 0 0.0701f
C27533 VPWR.n917 0 0.0391f
C27534 VPWR.n918 0 0.0117f
C27535 VPWR.n919 0 0.0108f
C27536 VPWR.n920 0 0.00918f
C27537 VPWR.n921 0 0.109f
C27538 VPWR.n922 0 0.15f
C27539 VPWR.n923 0 0.018f
C27540 VPWR.n924 0 0.0926f
C27541 VPWR.n925 0 0.0199f
C27542 VPWR.n926 0 0.0199f
C27543 VPWR.n927 0 0.0199f
C27544 VPWR.n928 0 0.0118f
C27545 VPWR.n929 0 0.088f
C27546 VPWR.n930 0 0.0345f
C27547 VPWR.n931 0 0.018f
C27548 VPWR.n932 0 0.011f
C27549 VPWR.n933 0 0.0199f
C27550 VPWR.n934 0 0.0192f
C27551 VPWR.n935 0 0.0199f
C27552 VPWR.n936 0 0.0199f
C27553 VPWR.n937 0 0.0117f
C27554 VPWR.n938 0 0.00399f
C27555 VPWR.n939 0 0.0507f
C27556 VPWR.n940 0 0.0181f
C27557 VPWR.n941 0 0.0199f
C27558 VPWR.n942 0 0.0199f
C27559 VPWR.t235 0 0.068f
C27560 VPWR.n943 0 0.0939f
C27561 VPWR.n944 0 0.0391f
C27562 VPWR.n945 0 0.0535f
C27563 VPWR.n946 0 0.0619f
C27564 VPWR.n947 0 0.0118f
C27565 VPWR.n948 0 0.00258f
C27566 VPWR.n949 0 0.00291f
C27567 VPWR.n950 0 0.00498f
C27568 VPWR.n951 0 0.00281f
C27569 VPWR.n952 0 0.00313f
C27570 VPWR.n953 0 0.00988f
C27571 VPWR.n954 0 0.00496f
C27572 VPWR.n955 0 0.00208f
C27573 VPWR.n956 0 0.00126f
C27574 VPWR.n957 0 0.00237f
C27575 VPWR.n958 0 0.376f
C27576 VPWR.n960 0 0.0108f
C27577 VPWR.n962 0 0.0115f
C27578 VPWR.n963 0 2.79e-20
C27579 VPWR.n964 0 0.00329f
C27580 VPWR.n965 0 0.00208f
C27581 VPWR.n966 0 0.00302f
C27582 VPWR.n967 0 0.00248f
C27583 VPWR.n968 0 0.00173f
C27584 VPWR.n969 0 0.014f
C27585 VPWR.n970 0 0.00194f
C27586 VPWR.n971 0 0.0013f
C27587 VPWR.n972 0 0.00108f
C27588 VPWR.n973 0 0.00194f
C27589 VPWR.n974 0 0.00173f
C27590 VPWR.n975 0 0.0014f
C27591 VPWR.n976 0 8.64e-19
C27592 VPWR.n977 0 0.00108f
C27593 VPWR.n978 0 0.00248f
C27594 VPWR.n979 0 0.00378f
C27595 VPWR.n980 0 0.00194f
C27596 VPWR.n981 0 0.00173f
C27597 VPWR.n982 0 0.0027f
C27598 VPWR.n983 0 0.00119f
C27599 VPWR.n984 0 0.00486f
C27600 VPWR.n985 0 0.00389f
C27601 VPWR.n986 0 0.00173f
C27602 VPWR.n987 0 0.0027f
C27603 VPWR.t36 0 0.068f
C27604 VPWR.n988 0 0.00482f
C27605 VPWR.n989 0 0.0329f
C27606 VPWR.n990 0 0.103f
C27607 VPWR.n991 0 0.0261f
C27608 VPWR.n992 0 0.0214f
C27609 VPWR.n993 0 0.00119f
C27610 VPWR.t66 0 0.068f
C27611 VPWR.n994 0 0.0535f
C27612 VPWR.n995 0 0.0391f
C27613 VPWR.n996 0 0.0701f
C27614 VPWR.t378 0 0.068f
C27615 VPWR.n997 0 0.0695f
C27616 VPWR.n998 0 0.0391f
C27617 VPWR.n999 0 0.0701f
C27618 VPWR.n1000 0 0.0385f
C27619 VPWR.t231 0 0.0417f
C27620 VPWR.t305 0 0.0417f
C27621 VPWR.n1001 0 0.0644f
C27622 VPWR.n1002 0 0.386f
C27623 VPWR.t247 0 0.0417f
C27624 VPWR.t369 0 0.0417f
C27625 VPWR.n1003 0 0.383f
C27626 VPWR.n1004 0 0.0208f
C27627 VPWR.n1005 0 0.0208f
C27628 VPWR.n1006 0 0.0118f
C27629 VPWR.n1007 0 0.0179f
C27630 VPWR.n1008 0 0.01f
C27631 VPWR.n1009 0 0.00537f
C27632 VPWR.n1010 0 0.0675f
C27633 VPWR.n1011 0 0.0118f
C27634 VPWR.n1012 0 0.0199f
C27635 VPWR.n1013 0 0.0199f
C27636 VPWR.n1014 0 0.018f
C27637 VPWR.n1015 0 0.049f
C27638 VPWR.n1016 0 0.00655f
C27639 VPWR.n1017 0 0.0714f
C27640 VPWR.n1018 0 0.0199f
C27641 VPWR.n1019 0 0.023f
C27642 VPWR.n1020 0 0.0199f
C27643 VPWR.n1021 0 0.018f
C27644 VPWR.n1022 0 0.046f
C27645 VPWR.n1023 0 0.0927f
C27646 VPWR.n1024 0 0.0118f
C27647 VPWR.n1025 0 0.0199f
C27648 VPWR.n1026 0 0.0199f
C27649 VPWR.n1027 0 0.018f
C27650 VPWR.n1028 0 0.0469f
C27651 VPWR.n1029 0 0.0342f
C27652 VPWR.n1030 0 0.0672f
C27653 VPWR.n1031 0 0.0199f
C27654 VPWR.n1032 0 0.0189f
C27655 VPWR.n1033 0 0.0199f
C27656 VPWR.n1034 0 0.018f
C27657 VPWR.n1035 0 0.0853f
C27658 VPWR.n1036 0 0.0757f
C27659 VPWR.n1037 0 0.0118f
C27660 VPWR.n1038 0 0.0721f
C27661 VPWR.n1039 0 0.018f
C27662 VPWR.n1040 0 0.00983f
C27663 VPWR.n1041 0 0.00184f
C27664 VPWR.n1042 0 0.00881f
C27665 VPWR.n1043 0 0.00496f
C27666 VPWR.n1044 0 0.00323f
C27667 VPWR.n1045 0 0.00248f
C27668 VPWR.n1046 0 0.00344f
C27669 VPWR.n1047 0 0.00208f
C27670 VPWR.n1049 0 0.00329f
C27671 VPWR.n1050 0 0.00208f
C27672 VPWR.n1051 0 0.0027f
C27673 VPWR.n1052 0 0.00497f
C27674 VPWR.n1053 0 0.00367f
C27675 VPWR.n1054 0 0.00281f
C27676 VPWR.n1055 0 0.00162f
C27677 VPWR.n1056 0 0.00205f
C27678 VPWR.n1057 0 0.00443f
C27679 VPWR.n1058 0 0.00302f
C27680 VPWR.n1059 0 0.00443f
C27681 VPWR.n1060 0 0.00281f
C27682 VPWR.n1061 0 8.64e-19
C27683 VPWR.n1062 0 0.00238f
C27684 VPWR.t363 0 0.0726f
C27685 VPWR.n1063 0 0.0391f
C27686 VPWR.n1064 0 0.267f
C27687 VPWR.n1065 0 0.0391f
C27688 VPWR.n1066 0 0.0917f
C27689 VPWR.n1067 0 0.0639f
C27690 VPWR.t139 0 0.0774f
C27691 VPWR.t18 0 0.0774f
C27692 VPWR.n1068 0 0.502f
C27693 VPWR.n1069 0 0.00259f
C27694 VPWR.n1070 0 0.00275f
C27695 VPWR.n1071 0 0.00525f
C27696 VPWR.n1072 0 0.00162f
C27697 VPWR.n1073 0 0.0014f
C27698 VPWR.n1074 0 0.0014f
C27699 VPWR.n1075 0 0.00344f
C27700 VPWR.n1076 0 0.00248f
C27701 VPWR.n1077 0 0.00329f
C27702 VPWR.n1078 0 0.381f
C27703 VPWR.n1079 0 0.0412f
C27704 VPWR.n1080 0 0.368f
C27705 VPWR.n1081 0 0.347f
C27706 VPWR.n1082 0 0.00248f
C27707 VPWR.n1083 0 0.00344f
C27708 VPWR.n1084 0 0.00208f
C27709 VPWR.n1085 0 0.00323f
C27710 VPWR.n1086 0 0.00468f
C27711 VPWR.n1087 0 0.00323f
C27712 VPWR.n1088 0 0.00208f
C27713 VPWR.n1090 0 0.00329f
C27714 VPWR.n1091 0 0.00208f
C27715 VPWR.n1092 0 0.00302f
C27716 VPWR.n1093 0 0.00248f
C27717 VPWR.n1094 0 0.00173f
C27718 VPWR.n1095 0 0.0027f
C27719 VPWR.n1096 0 0.00248f
C27720 VPWR.n1097 0 0.00205f
C27721 VPWR.n1098 0 0.00162f
C27722 VPWR.n1099 0 0.00335f
C27723 VPWR.n1100 0 0.00421f
C27724 VPWR.n1101 0 0.00248f
C27725 VPWR.n1102 0 7.56e-19
C27726 VPWR.n1103 0 8.64e-19
C27727 VPWR.n1104 0 0.00108f
C27728 VPWR.n1105 0 0.00205f
C27729 VPWR.n1106 0 0.00248f
C27730 VPWR.n1107 0 0.0027f
C27731 VPWR.n1108 0 0.00302f
C27732 VPWR.n1109 0 0.00184f
C27733 VPWR.n1110 0 9.72e-19
C27734 VPWR.n1111 0 0.0014f
C27735 VPWR.n1112 0 8.64e-19
C27736 VPWR.n1113 0 0.00108f
C27737 VPWR.n1114 0 0.00248f
C27738 VPWR.n1115 0 0.00389f
C27739 VPWR.n1116 0 0.00357f
C27740 VPWR.n1117 0 0.00281f
C27741 VPWR.n1118 0 0.00258f
C27742 VPWR.t387 0 0.0722f
C27743 VPWR.n1119 0 0.207f
C27744 VPWR.n1120 0 0.0685f
C27745 VPWR.n1121 0 0.0926f
C27746 VPWR.n1122 0 0.0668f
C27747 VPWR.n1123 0 0.0715f
C27748 VPWR.t14 0 0.111f
C27749 VPWR.n1124 0 0.288f
C27750 VPWR.n1125 0 0.153f
C27751 VPWR.n1126 0 0.044f
C27752 VPWR.n1127 0 0.01f
C27753 VPWR.t40 0 0.116f
C27754 VPWR.n1128 0 0.432f
C27755 VPWR.n1129 0 0.0818f
C27756 VPWR.t359 0 0.0724f
C27757 VPWR.n1130 0 0.0522f
C27758 VPWR.n1131 0 0.00119f
C27759 VPWR.n1132 0 0.00119f
C27760 VPWR.n1133 0 0.00344f
C27761 VPWR.n1134 0 0.00248f
C27762 VPWR.n1135 0 0.00329f
C27763 VPWR.n1137 0 0.00329f
C27764 VPWR.n1138 0 0.00208f
C27765 VPWR.n1139 0 0.00259f
C27766 VPWR.n1140 0 0.00593f
C27767 VPWR.t76 0 0.0774f
C27768 VPWR.n1141 0 0.0534f
C27769 VPWR.t351 0 0.0417f
C27770 VPWR.t327 0 0.0417f
C27771 VPWR.n1142 0 0.384f
C27772 VPWR.n1143 0 0.019f
C27773 VPWR.t50 0 0.068f
C27774 VPWR.t166 0 0.0711f
C27775 VPWR.n1144 0 0.195f
C27776 VPWR.n1145 0 0.0877f
C27777 VPWR.n1146 0 0.0391f
C27778 VPWR.n1147 0 0.0701f
C27779 VPWR.n1148 0 0.0475f
C27780 VPWR.n1149 0 0.0246f
C27781 VPWR.n1150 0 0.0173f
C27782 VPWR.n1151 0 0.0199f
C27783 VPWR.n1152 0 0.0118f
C27784 VPWR.n1153 0 0.00994f
C27785 VPWR.n1154 0 0.0616f
C27786 VPWR.n1155 0 0.00695f
C27787 VPWR.n1156 0 0.018f
C27788 VPWR.n1157 0 0.0526f
C27789 VPWR.n1158 0 0.0199f
C27790 VPWR.n1159 0 0.00816f
C27791 VPWR.n1160 0 0.0199f
C27792 VPWR.n1161 0 0.0117f
C27793 VPWR.n1162 0 0.0276f
C27794 VPWR.t182 0 0.0774f
C27795 VPWR.n1163 0 0.503f
C27796 VPWR.n1164 0 0.0302f
C27797 VPWR.n1165 0 0.018f
C27798 VPWR.n1166 0 0.0578f
C27799 VPWR.n1167 0 0.0199f
C27800 VPWR.n1168 0 0.0314f
C27801 VPWR.n1169 0 0.0199f
C27802 VPWR.n1170 0 0.0148f
C27803 VPWR.n1171 0 0.0199f
C27804 VPWR.n1172 0 0.0117f
C27805 VPWR.n1173 0 0.0342f
C27806 VPWR.n1174 0 0.0613f
C27807 VPWR.n1175 0 0.0181f
C27808 VPWR.t181 0 0.0876f
C27809 VPWR.n1176 0 0.149f
C27810 VPWR.n1177 0 0.0199f
C27811 VPWR.n1178 0 0.0522f
C27812 VPWR.n1179 0 0.0199f
C27813 VPWR.n1180 0 0.0758f
C27814 VPWR.n1181 0 0.0199f
C27815 VPWR.n1182 0 0.0363f
C27816 VPWR.n1183 0 0.0602f
C27817 VPWR.n1184 0 0.0186f
C27818 VPWR.n1185 0 0.00994f
C27819 VPWR.n1186 0 0.00184f
C27820 VPWR.n1187 0 0.015f
C27821 VPWR.n1188 0 0.0357f
C27822 VPWR.n1189 0 7.56e-19
C27823 VPWR.n1190 0 0.0408f
C27824 VPWR.n1191 0 0.00421f
C27825 VPWR.n1192 0 0.00248f
C27826 VPWR.n1193 0 5.4e-19
C27827 VPWR.n1194 0 0.00344f
C27828 VPWR.n1195 0 0.00248f
C27829 VPWR.n1196 0 0.00329f
C27830 VPWR.n1197 0 0.00208f
C27831 VPWR.n1198 0 0.00498f
C27832 VPWR.n1199 0 0.0123f
C27833 VPWR.n1200 0 0.00313f
C27834 VPWR.n1201 0 0.00397f
C27835 VPWR.n1202 0 0.00151f
C27836 VPWR.n1203 0 0.011f
C27837 VPWR.n1204 0 0.00162f
C27838 VPWR.n1205 0 0.00119f
C27839 VPWR.n1206 0 0.00184f
C27840 VPWR.n1207 0 0.00259f
C27841 VPWR.n1208 0 0.00119f
C27842 VPWR.n1209 0 0.00585f
C27843 VPWR.n1210 0 0.0743f
C27844 VPWR.t165 0 0.0774f
C27845 VPWR.n1211 0 0.296f
C27846 VPWR.t135 0 0.0951f
C27847 VPWR.n1212 0 0.333f
C27848 VPWR.t193 0 0.068f
C27849 VPWR.n1213 0 0.0535f
C27850 VPWR.n1214 0 0.0391f
C27851 VPWR.n1215 0 0.0942f
C27852 VPWR.n1216 0 0.049f
C27853 VPWR.t113 0 0.068f
C27854 VPWR.n1217 0 0.0701f
C27855 VPWR.n1218 0 0.0199f
C27856 VPWR.n1219 0 0.306f
C27857 VPWR.n1220 0 0.0725f
C27858 VPWR.n1221 0 0.0118f
C27859 VPWR.t65 0 0.068f
C27860 VPWR.n1222 0 0.0738f
C27861 VPWR.n1223 0 0.0777f
C27862 VPWR.n1224 0 0.0668f
C27863 VPWR.n1225 0 0.0449f
C27864 VPWR.t222 0 0.068f
C27865 VPWR.n1226 0 0.0701f
C27866 VPWR.n1227 0 0.0391f
C27867 VPWR.n1228 0 0.0695f
C27868 VPWR.n1229 0 0.0504f
C27869 VPWR.n1230 0 0.1f
C27870 VPWR.n1231 0 0.0818f
C27871 VPWR.n1232 0 0.0805f
C27872 VPWR.n1233 0 0.0742f
C27873 VPWR.n1234 0 0.00281f
C27874 VPWR.n1235 0 0.00329f
C27875 VPWR.n1236 0 0.00208f
C27876 VPWR.n1237 0 0.00496f
C27877 VPWR.n1238 0 0.00302f
C27878 VPWR.n1239 0 0.00248f
C27879 VPWR.n1240 0 0.00173f
C27880 VPWR.n1241 0 0.0027f
C27881 VPWR.n1242 0 0.00248f
C27882 VPWR.n1243 0 0.00205f
C27883 VPWR.n1244 0 0.00743f
C27884 VPWR.n1245 0 0.00259f
C27885 VPWR.n1246 0 0.00275f
C27886 VPWR.n1247 0 0.00525f
C27887 VPWR.n1248 0 0.00162f
C27888 VPWR.n1249 0 0.0014f
C27889 VPWR.n1250 0 0.0612f
C27890 VPWR.t184 0 0.0863f
C27891 VPWR.n1251 0 0.0993f
C27892 VPWR.n1252 0 0.101f
C27893 VPWR.n1253 0 0.11f
C27894 VPWR.t134 0 0.111f
C27895 VPWR.n1254 0 0.288f
C27896 VPWR.n1255 0 0.0572f
C27897 VPWR.n1256 0 0.119f
C27898 VPWR.n1257 0 0.114f
C27899 VPWR.t285 0 0.068f
C27900 VPWR.n1258 0 0.0701f
C27901 VPWR.n1259 0 0.0512f
C27902 VPWR.n1260 0 0.0656f
C27903 VPWR.n1261 0 0.0619f
C27904 VPWR.n1262 0 0.00258f
C27905 VPWR.n1263 0 0.00498f
C27906 VPWR.n1264 0 0.00291f
C27907 VPWR.n1265 0 0.0504f
C27908 VPWR.n1266 0 0.307f
C27909 VPWR.n1267 0 0.279f
C27910 VPWR.t204 0 0.0876f
C27911 VPWR.n1268 0 0.149f
C27912 VPWR.n1269 0 0.0971f
C27913 VPWR.t109 0 0.116f
C27914 VPWR.n1270 0 0.322f
C27915 VPWR.n1271 0 0.154f
C27916 VPWR.n1272 0 0.0181f
C27917 VPWR.n1273 0 0.128f
C27918 VPWR.n1274 0 0.0535f
C27919 VPWR.n1275 0 0.049f
C27920 VPWR.t310 0 0.068f
C27921 VPWR.n1276 0 0.0942f
C27922 VPWR.n1277 0 0.0391f
C27923 VPWR.n1278 0 0.0535f
C27924 VPWR.t89 0 0.0724f
C27925 VPWR.n1279 0 0.207f
C27926 VPWR.n1280 0 0.0429f
C27927 VPWR.n1281 0 0.0027f
C27928 VPWR.n1282 0 0.00861f
C27929 VPWR.n1283 0 0.00443f
C27930 VPWR.n1284 0 0.00281f
C27931 VPWR.n1285 0 0.00162f
C27932 VPWR.n1286 0 0.00164f
C27933 VPWR.n1287 0 0.0462f
C27934 VPWR.n1288 0 0.0213f
C27935 VPWR.n1289 0 0.00822f
C27936 VPWR.t323 0 0.073f
C27937 VPWR.n1290 0 0.0975f
C27938 VPWR.n1291 0 0.101f
C27939 VPWR.n1292 0 0.131f
C27940 VPWR.n1293 0 0.0552f
C27941 VPWR.n1294 0 0.00212f
C27942 VPWR.n1295 0 0.00302f
C27943 VPWR.n1296 0 0.00248f
C27944 VPWR.n1297 0 0.00173f
C27945 VPWR.n1298 0 0.00329f
C27946 VPWR.n1299 0 0.00208f
C27947 VPWR.n1300 0 0.381f
C27948 VPWR.n1301 0 0.381f
C27949 VPWR.n1302 0 0.00248f
C27950 VPWR.n1303 0 0.00344f
C27951 VPWR.n1304 0 0.00468f
C27952 VPWR.n1305 0 0.00323f
C27953 VPWR.n1306 0 0.00208f
C27954 VPWR.n1308 0 0.00329f
C27955 VPWR.n1309 0 0.00208f
C27956 VPWR.n1310 0 0.00496f
C27957 VPWR.n1311 0 0.00323f
C27958 VPWR.n1312 0 0.00248f
C27959 VPWR.n1313 0 0.00344f
C27960 VPWR.n1314 0 0.00208f
C27961 VPWR.n1316 0 0.00329f
C27962 VPWR.n1317 0 0.00208f
C27963 VPWR.n1318 0 0.0027f
C27964 VPWR.n1319 0 0.00497f
C27965 VPWR.n1320 0 0.00302f
C27966 VPWR.n1321 0 0.00248f
C27967 VPWR.n1322 0 0.00173f
C27968 VPWR.n1323 0 0.00486f
C27969 VPWR.n1324 0 0.00389f
C27970 VPWR.n1325 0 0.00173f
C27971 VPWR.n1326 0 0.0027f
C27972 VPWR.t274 0 0.068f
C27973 VPWR.n1327 0 0.0665f
C27974 VPWR.n1328 0 0.0283f
C27975 VPWR.n1329 0 0.0179f
C27976 VPWR.n1330 0 0.00119f
C27977 VPWR.n1331 0 0.0321f
C27978 VPWR.n1332 0 0.0518f
C27979 VPWR.t230 0 0.068f
C27980 VPWR.n1333 0 0.0701f
C27981 VPWR.n1334 0 0.0199f
C27982 VPWR.n1335 0 0.00655f
C27983 VPWR.n1336 0 0.0118f
C27984 VPWR.t169 0 0.0774f
C27985 VPWR.t383 0 0.0774f
C27986 VPWR.n1337 0 0.501f
C27987 VPWR.t287 0 0.0417f
C27988 VPWR.t262 0 0.0417f
C27989 VPWR.n1338 0 0.383f
C27990 VPWR.n1339 0 0.0208f
C27991 VPWR.n1340 0 0.0267f
C27992 VPWR.n1341 0 0.0107f
C27993 VPWR.n1342 0 0.0447f
C27994 VPWR.n1343 0 0.00621f
C27995 VPWR.n1344 0 0.0892f
C27996 VPWR.n1345 0 0.018f
C27997 VPWR.n1346 0 0.0118f
C27998 VPWR.n1347 0 0.0675f
C27999 VPWR.n1348 0 0.0695f
C28000 VPWR.n1349 0 0.0391f
C28001 VPWR.n1350 0 0.0199f
C28002 VPWR.n1351 0 0.018f
C28003 VPWR.n1352 0 0.0482f
C28004 VPWR.n1353 0 0.00417f
C28005 VPWR.n1354 0 0.0118f
C28006 VPWR.n1355 0 0.0621f
C28007 VPWR.n1356 0 0.0199f
C28008 VPWR.n1357 0 0.018f
C28009 VPWR.n1358 0 0.0201f
C28010 VPWR.n1359 0 0.0748f
C28011 VPWR.n1360 0 0.0118f
C28012 VPWR.n1361 0 0.0771f
C28013 VPWR.n1362 0 0.0199f
C28014 VPWR.n1363 0 0.0391f
C28015 VPWR.n1364 0 0.0199f
C28016 VPWR.t324 0 0.068f
C28017 VPWR.n1365 0 0.0701f
C28018 VPWR.n1366 0 0.0482f
C28019 VPWR.n1367 0 0.0199f
C28020 VPWR.n1368 0 0.0199f
C28021 VPWR.n1369 0 0.018f
C28022 VPWR.n1370 0 0.00994f
C28023 VPWR.n1371 0 0.0686f
C28024 VPWR.n1372 0 0.0704f
C28025 VPWR.n1373 0 0.0118f
C28026 VPWR.n1374 0 0.0886f
C28027 VPWR.n1375 0 0.018f
C28028 VPWR.n1376 0 0.00983f
C28029 VPWR.n1377 0 0.00184f
C28030 VPWR.n1378 0 0.00881f
C28031 VPWR.n1379 0 0.00119f
C28032 VPWR.n1380 0 0.0027f
C28033 VPWR.n1381 0 0.00173f
C28034 VPWR.n1382 0 0.00194f
C28035 VPWR.n1383 0 0.00378f
C28036 VPWR.n1384 0 0.00248f
C28037 VPWR.n1385 0 0.00108f
C28038 VPWR.n1386 0 8.64e-19
C28039 VPWR.n1387 0 0.0014f
C28040 VPWR.n1388 0 4.32e-19
C28041 VPWR.n1389 0 0.00184f
C28042 VPWR.n1390 0 0.00108f
C28043 VPWR.n1391 0 0.0013f
C28044 VPWR.n1392 0 0.00194f
C28045 VPWR.n1393 0 0.00367f
C28046 VPWR.n1394 0 0.00281f
C28047 VPWR.n1395 0 0.00162f
C28048 VPWR.n1396 0 0.00205f
C28049 VPWR.n1397 0 0.00443f
C28050 VPWR.n1398 0 0.00302f
C28051 VPWR.n1399 0 0.00443f
C28052 VPWR.n1400 0 0.00281f
C28053 VPWR.n1401 0 8.64e-19
C28054 VPWR.n1402 0 0.00238f
C28055 VPWR.n1403 0 0.0329f
C28056 VPWR.n1404 0 0.0213f
C28057 VPWR.n1405 0 0.00822f
C28058 VPWR.n1406 0 0.101f
C28059 VPWR.n1407 0 0.0661f
C28060 VPWR.t337 0 0.0954f
C28061 VPWR.n1408 0 0.332f
C28062 VPWR.n1409 0 0.0922f
C28063 VPWR.t31 0 0.0951f
C28064 VPWR.n1410 0 0.333f
C28065 VPWR.t180 0 0.0774f
C28066 VPWR.n1411 0 0.295f
C28067 VPWR.n1412 0 0.0942f
C28068 VPWR.t301 0 0.116f
C28069 VPWR.n1413 0 0.322f
C28070 VPWR.n1414 0 0.118f
C28071 VPWR.t244 0 0.107f
C28072 VPWR.n1415 0 0.00259f
C28073 VPWR.n1416 0 0.00421f
C28074 VPWR.n1417 0 0.00378f
C28075 VPWR.n1418 0 0.00162f
C28076 VPWR.n1419 0 0.0014f
C28077 VPWR.n1420 0 0.0014f
C28078 VPWR.n1421 0 0.00344f
C28079 VPWR.n1422 0 0.00248f
C28080 VPWR.n1423 0 0.00329f
C28081 VPWR.n1424 0 0.378f
C28082 VPWR.n1425 0 0.381f
C28083 VPWR.n1426 0 0.00248f
C28084 VPWR.n1427 0 0.00344f
C28085 VPWR.n1428 0 0.00208f
C28086 VPWR.n1429 0 0.00323f
C28087 VPWR.n1430 0 0.00468f
C28088 VPWR.n1431 0 0.00323f
C28089 VPWR.n1432 0 0.00208f
C28090 VPWR.n1434 0 0.0217f
C28091 VPWR.n1435 0 0.00344f
C28092 VPWR.n1436 0 0.00248f
C28093 VPWR.n1437 0 0.00329f
C28094 VPWR.n1438 0 0.00483f
C28095 VPWR.n1439 0 0.00208f
C28096 VPWR.n1441 0 0.381f
C28097 VPWR.n1442 0 0.381f
C28098 VPWR.n1443 0 0.00248f
C28099 VPWR.n1444 0 0.00344f
C28100 VPWR.n1445 0 0.00208f
C28101 VPWR.n1446 0 0.00323f
C28102 VPWR.n1447 0 0.00468f
C28103 VPWR.n1448 0 0.00323f
C28104 VPWR.n1449 0 0.00208f
C28105 VPWR.n1451 0 0.00329f
C28106 VPWR.n1452 0 0.00208f
C28107 VPWR.n1453 0 0.00302f
C28108 VPWR.n1454 0 0.00248f
C28109 VPWR.n1455 0 0.00173f
C28110 VPWR.n1456 0 0.0027f
C28111 VPWR.n1457 0 0.00248f
C28112 VPWR.n1458 0 0.00205f
C28113 VPWR.n1459 0 0.00162f
C28114 VPWR.n1460 0 0.00335f
C28115 VPWR.n1461 0 0.00421f
C28116 VPWR.n1462 0 0.00248f
C28117 VPWR.n1463 0 7.56e-19
C28118 VPWR.n1464 0 8.64e-19
C28119 VPWR.n1465 0 0.00108f
C28120 VPWR.n1466 0 0.00205f
C28121 VPWR.n1467 0 0.00248f
C28122 VPWR.n1468 0 0.0027f
C28123 VPWR.n1469 0 0.00302f
C28124 VPWR.n1470 0 0.00184f
C28125 VPWR.n1471 0 9.72e-19
C28126 VPWR.n1472 0 0.0014f
C28127 VPWR.n1473 0 8.64e-19
C28128 VPWR.n1474 0 0.00108f
C28129 VPWR.n1475 0 0.00248f
C28130 VPWR.n1476 0 0.00389f
C28131 VPWR.n1477 0 0.00357f
C28132 VPWR.n1478 0 0.00281f
C28133 VPWR.n1479 0 0.00265f
C28134 VPWR.n1480 0 0.00482f
C28135 VPWR.n1481 0 0.013f
C28136 VPWR.n1482 0 0.0404f
C28137 VPWR.n1483 0 0.0202f
C28138 VPWR.n1484 0 0.0262f
C28139 VPWR.n1485 0 0.189f
C28140 VPWR.t338 0 0.0716f
C28141 VPWR.n1486 0 0.196f
C28142 VPWR.n1487 0 0.01f
C28143 VPWR.t223 0 0.068f
C28144 VPWR.n1488 0 0.0476f
C28145 VPWR.n1489 0 0.0701f
C28146 VPWR.n1490 0 0.0841f
C28147 VPWR.n1491 0 0.0799f
C28148 VPWR.t366 0 0.0724f
C28149 VPWR.n1492 0 0.0143f
C28150 VPWR.n1493 0 0.0455f
C28151 VPWR.t27 0 0.0724f
C28152 VPWR.n1494 0 0.0103f
C28153 VPWR.t357 0 0.0774f
C28154 VPWR.t83 0 0.0774f
C28155 VPWR.n1495 0 0.503f
C28156 VPWR.n1496 0 0.0014f
C28157 VPWR.n1497 0 0.00421f
C28158 VPWR.n1498 0 0.00248f
C28159 VPWR.n1499 0 5.4e-19
C28160 VPWR.n1500 0 0.00344f
C28161 VPWR.n1501 0 0.00248f
C28162 VPWR.n1502 0 0.00329f
C28163 VPWR.n1503 0 0.00206f
C28164 VPWR.n1504 0 1.77f
C28165 VPWR.n1505 0 0.933f
C28166 VPWR.n1506 0 0.0629f
C28167 VPWR.n1507 0 1.87f
C28168 VPWR.n1508 0 1.87f
C28169 VPWR.n1509 0 0.0655f
C28170 VPWR.n1510 0 1.87f
C28171 VPWR.n1511 0 1.86f
C28172 VPWR.n1512 0 0.00323f
C28173 VPWR.n1513 0 0.00208f
C28174 VPWR.n1514 0 0.00457f
C28175 VPWR.n1515 0 0.00206f
C28176 VPWR.n1517 0 0.00329f
C28177 VPWR.n1518 0 0.00208f
C28178 VPWR.n1519 0 0.00259f
C28179 VPWR.n1520 0 0.0634f
C28180 VPWR.n1521 0 0.0199f
C28181 VPWR.t384 0 0.0876f
C28182 VPWR.t156 0 0.0716f
C28183 VPWR.n1522 0 0.196f
C28184 VPWR.n1523 0 0.0519f
C28185 VPWR.n1524 0 0.0584f
C28186 VPWR.t385 0 0.0774f
C28187 VPWR.t108 0 0.0417f
C28188 VPWR.t88 0 0.0417f
C28189 VPWR.n1525 0 0.383f
C28190 VPWR.n1526 0 0.0384f
C28191 VPWR.n1527 0 0.0421f
C28192 VPWR.t103 0 0.0774f
C28193 VPWR.n1528 0 0.501f
C28194 VPWR.n1529 0 0.0435f
C28195 VPWR.n1530 0 0.018f
C28196 VPWR.n1531 0 0.05f
C28197 VPWR.n1532 0 0.0199f
C28198 VPWR.n1533 0 0.0118f
C28199 VPWR.n1534 0 0.039f
C28200 VPWR.n1535 0 0.0464f
C28201 VPWR.n1536 0 0.0107f
C28202 VPWR.n1537 0 0.0173f
C28203 VPWR.n1538 0 0.018f
C28204 VPWR.n1539 0 0.0118f
C28205 VPWR.n1540 0 0.134f
C28206 VPWR.n1541 0 0.0952f
C28207 VPWR.n1542 0 0.0552f
C28208 VPWR.n1543 0 0.0995f
C28209 VPWR.n1544 0 0.0118f
C28210 VPWR.n1545 0 0.00994f
C28211 VPWR.n1546 0 0.0108f
C28212 VPWR.n1547 0 0.00621f
C28213 VPWR.n1548 0 0.105f
C28214 VPWR.n1549 0 0.0172f
C28215 VPWR.n1550 0 0.0469f
C28216 VPWR.n1551 0 0.0199f
C28217 VPWR.t127 0 0.107f
C28218 VPWR.n1552 0 0.201f
C28219 VPWR.n1553 0 0.0386f
C28220 VPWR.n1554 0 0.0199f
C28221 VPWR.n1555 0 0.0737f
C28222 VPWR.n1556 0 0.0199f
C28223 VPWR.n1557 0 0.0557f
C28224 VPWR.n1558 0 0.0199f
C28225 VPWR.n1559 0 0.0522f
C28226 VPWR.n1560 0 0.0199f
C28227 VPWR.n1561 0 0.0363f
C28228 VPWR.n1562 0 0.0488f
C28229 VPWR.n1563 0 0.0186f
C28230 VPWR.n1564 0 0.00994f
C28231 VPWR.n1565 0 0.00184f
C28232 VPWR.n1566 0 0.015f
C28233 VPWR.n1567 0 0.0467f
C28234 VPWR.n1568 0 7.56e-19
C28235 VPWR.n1569 0 0.00184f
C28236 VPWR.n1570 0 0.0457f
C28237 VPWR.n1571 0 0.0354f
C28238 VPWR.n1572 0 0.0516f
C28239 VPWR.t79 0 0.068f
C28240 VPWR.n1573 0 0.0701f
C28241 VPWR.n1574 0 0.0607f
C28242 VPWR.n1575 0 0.0571f
C28243 VPWR.n1576 0 0.0619f
C28244 VPWR.n1577 0 0.00497f
C28245 VPWR.n1578 0 0.381f
C28246 VPWR.n1579 0 0.00344f
C28247 VPWR.n1580 0 0.00248f
C28248 VPWR.n1581 0 0.00329f
C28249 VPWR.n1582 0 0.00208f
C28250 VPWR.n1583 0 0.00302f
C28251 VPWR.n1584 0 0.00248f
C28252 VPWR.n1585 0 0.00173f
C28253 VPWR.n1586 0 0.014f
C28254 VPWR.n1587 0 0.00194f
C28255 VPWR.n1588 0 0.0013f
C28256 VPWR.n1589 0 0.00108f
C28257 VPWR.n1590 0 0.00194f
C28258 VPWR.n1591 0 0.00173f
C28259 VPWR.n1592 0 0.0014f
C28260 VPWR.n1593 0 8.64e-19
C28261 VPWR.n1594 0 0.00108f
C28262 VPWR.n1595 0 0.00248f
C28263 VPWR.n1596 0 0.00378f
C28264 VPWR.n1597 0 0.00194f
C28265 VPWR.n1598 0 0.00173f
C28266 VPWR.n1599 0 0.0027f
C28267 VPWR.n1600 0 0.00119f
C28268 VPWR.n1601 0 0.00486f
C28269 VPWR.n1602 0 0.00389f
C28270 VPWR.n1603 0 0.00173f
C28271 VPWR.n1604 0 0.0027f
C28272 VPWR.t138 0 0.068f
C28273 VPWR.n1605 0 0.00482f
C28274 VPWR.n1606 0 0.0466f
C28275 VPWR.n1607 0 0.0879f
C28276 VPWR.n1608 0 0.0261f
C28277 VPWR.n1609 0 0.0179f
C28278 VPWR.n1610 0 0.00119f
C28279 VPWR.n1611 0 0.0199f
C28280 VPWR.n1612 0 0.0107f
C28281 VPWR.n1613 0 0.0199f
C28282 VPWR.n1614 0 0.0699f
C28283 VPWR.n1615 0 0.0199f
C28284 VPWR.t248 0 0.068f
C28285 VPWR.n1616 0 0.0973f
C28286 VPWR.n1617 0 0.0935f
C28287 VPWR.n1618 0 0.0199f
C28288 VPWR.t116 0 0.068f
C28289 VPWR.n1619 0 0.0722f
C28290 VPWR.t250 0 0.068f
C28291 VPWR.n1620 0 0.0701f
C28292 VPWR.n1621 0 0.105f
C28293 VPWR.t55 0 0.0417f
C28294 VPWR.n1622 0 0.296f
C28295 VPWR.t98 0 0.0417f
C28296 VPWR.t81 0 0.0417f
C28297 VPWR.n1623 0 0.383f
C28298 VPWR.n1624 0 0.0208f
C28299 VPWR.n1625 0 0.0144f
C28300 VPWR.n1626 0 0.00994f
C28301 VPWR.n1627 0 0.0118f
C28302 VPWR.n1628 0 0.018f
C28303 VPWR.n1629 0 0.0565f
C28304 VPWR.n1630 0 0.0851f
C28305 VPWR.n1631 0 0.00994f
C28306 VPWR.n1632 0 0.0118f
C28307 VPWR.n1633 0 0.0948f
C28308 VPWR.n1634 0 0.106f
C28309 VPWR.n1635 0 0.0411f
C28310 VPWR.n1636 0 0.018f
C28311 VPWR.n1637 0 0.00994f
C28312 VPWR.n1638 0 0.0118f
C28313 VPWR.n1639 0 0.0691f
C28314 VPWR.n1640 0 0.105f
C28315 VPWR.n1641 0 0.0391f
C28316 VPWR.n1642 0 0.0199f
C28317 VPWR.n1643 0 0.018f
C28318 VPWR.n1644 0 0.0118f
C28319 VPWR.n1645 0 0.0292f
C28320 VPWR.n1646 0 0.0629f
C28321 VPWR.n1647 0 0.0556f
C28322 VPWR.n1648 0 0.0199f
C28323 VPWR.n1649 0 0.0199f
C28324 VPWR.n1650 0 0.0199f
C28325 VPWR.n1651 0 0.0525f
C28326 VPWR.n1652 0 0.0142f
C28327 VPWR.n1653 0 0.0419f
C28328 VPWR.n1654 0 0.0179f
C28329 VPWR.n1655 0 0.01f
C28330 VPWR.n1656 0 0.00372f
C28331 VPWR.n1657 0 0.0753f
C28332 VPWR.n1658 0 0.0118f
C28333 VPWR.n1659 0 0.0622f
C28334 VPWR.n1660 0 0.018f
C28335 VPWR.n1661 0 0.00983f
C28336 VPWR.n1662 0 0.00184f
C28337 VPWR.n1663 0 0.00881f
C28338 VPWR.n1664 0 0.00496f
C28339 VPWR.n1665 0 0.00302f
C28340 VPWR.n1666 0 0.00248f
C28341 VPWR.n1667 0 0.00173f
C28342 VPWR.n1668 0 0.014f
C28343 VPWR.n1669 0 0.00194f
C28344 VPWR.n1670 0 0.0013f
C28345 VPWR.n1671 0 0.00108f
C28346 VPWR.n1672 0 0.00194f
C28347 VPWR.n1673 0 0.00173f
C28348 VPWR.n1674 0 0.0014f
C28349 VPWR.n1675 0 8.64e-19
C28350 VPWR.n1676 0 0.00108f
C28351 VPWR.n1677 0 0.00248f
C28352 VPWR.n1678 0 0.00378f
C28353 VPWR.n1679 0 0.00194f
C28354 VPWR.n1680 0 0.00173f
C28355 VPWR.n1681 0 0.0027f
C28356 VPWR.n1682 0 0.00119f
C28357 VPWR.n1683 0 0.00486f
C28358 VPWR.n1684 0 0.00389f
C28359 VPWR.n1685 0 0.00173f
C28360 VPWR.n1686 0 0.0027f
C28361 VPWR.t25 0 0.068f
C28362 VPWR.n1687 0 0.00482f
C28363 VPWR.n1688 0 0.0329f
C28364 VPWR.n1689 0 0.0702f
C28365 VPWR.n1690 0 0.0261f
C28366 VPWR.n1691 0 0.0564f
C28367 VPWR.n1692 0 0.00119f
C28368 VPWR.n1693 0 0.00409f
C28369 VPWR.n1694 0 0.0667f
C28370 VPWR.n1695 0 0.00711f
C28371 VPWR.n1696 0 0.0533f
C28372 VPWR.n1697 0 0.018f
C28373 VPWR.t187 0 0.0876f
C28374 VPWR.t30 0 0.0726f
C28375 VPWR.n1698 0 0.0405f
C28376 VPWR.n1699 0 0.267f
C28377 VPWR.n1700 0 0.0391f
C28378 VPWR.n1701 0 0.0522f
C28379 VPWR.t146 0 0.0417f
C28380 VPWR.n1702 0 0.0208f
C28381 VPWR.t121 0 0.0417f
C28382 VPWR.n1703 0 0.384f
C28383 VPWR.n1704 0 0.0619f
C28384 VPWR.n1705 0 0.0118f
C28385 VPWR.n1706 0 0.0199f
C28386 VPWR.n1707 0 0.0199f
C28387 VPWR.n1708 0 0.018f
C28388 VPWR.n1709 0 0.15f
C28389 VPWR.n1710 0 0.115f
C28390 VPWR.n1711 0 0.00963f
C28391 VPWR.n1712 0 0.0118f
C28392 VPWR.n1713 0 0.018f
C28393 VPWR.n1714 0 0.0702f
C28394 VPWR.n1715 0 0.0634f
C28395 VPWR.n1716 0 0.0118f
C28396 VPWR.n1717 0 0.0577f
C28397 VPWR.n1718 0 0.0199f
C28398 VPWR.n1719 0 0.0552f
C28399 VPWR.n1720 0 0.0199f
C28400 VPWR.t381 0 0.068f
C28401 VPWR.n1721 0 0.0701f
C28402 VPWR.n1722 0 0.0482f
C28403 VPWR.n1723 0 0.0199f
C28404 VPWR.n1724 0 0.0199f
C28405 VPWR.n1725 0 0.018f
C28406 VPWR.n1726 0 0.00994f
C28407 VPWR.n1727 0 0.0595f
C28408 VPWR.n1728 0 0.0818f
C28409 VPWR.n1729 0 0.0118f
C28410 VPWR.n1730 0 0.0649f
C28411 VPWR.n1731 0 0.0199f
C28412 VPWR.n1732 0 0.0627f
C28413 VPWR.n1733 0 0.0199f
C28414 VPWR.t64 0 0.068f
C28415 VPWR.n1734 0 0.0701f
C28416 VPWR.n1735 0 0.0476f
C28417 VPWR.n1736 0 0.0199f
C28418 VPWR.n1737 0 0.0199f
C28419 VPWR.n1738 0 0.0179f
C28420 VPWR.n1739 0 0.01f
C28421 VPWR.n1740 0 0.0337f
C28422 VPWR.n1741 0 0.071f
C28423 VPWR.n1742 0 0.0118f
C28424 VPWR.n1743 0 0.062f
C28425 VPWR.n1744 0 0.018f
C28426 VPWR.n1745 0 0.00983f
C28427 VPWR.n1746 0 0.00184f
C28428 VPWR.n1747 0 0.00881f
C28429 VPWR.n1748 0 0.00495f
C28430 VPWR.n1749 0 0.00208f
C28431 VPWR.n1750 0 0.00257f
C28432 VPWR.n1751 0 0.00203f
C28433 VPWR.n1752 0 0.0027f
C28434 VPWR.n1753 0 0.00497f
C28435 VPWR.n1754 0 0.00367f
C28436 VPWR.n1755 0 0.00281f
C28437 VPWR.n1756 0 0.00162f
C28438 VPWR.n1757 0 0.00205f
C28439 VPWR.n1758 0 0.00443f
C28440 VPWR.n1759 0 0.00302f
C28441 VPWR.n1760 0 0.00443f
C28442 VPWR.n1761 0 0.00281f
C28443 VPWR.n1762 0 8.64e-19
C28444 VPWR.n1763 0 0.00238f
C28445 VPWR.t185 0 0.0718f
C28446 VPWR.n1764 0 0.208f
C28447 VPWR.t92 0 0.068f
C28448 VPWR.n1765 0 0.0695f
C28449 VPWR.n1766 0 0.0391f
C28450 VPWR.n1767 0 0.0701f
C28451 VPWR.n1768 0 0.0475f
C28452 VPWR.n1769 0 0.0738f
C28453 VPWR.n1770 0 0.0771f
C28454 VPWR.t329 0 0.068f
C28455 VPWR.n1771 0 0.0701f
C28456 VPWR.t115 0 0.068f
C28457 VPWR.n1772 0 0.0701f
C28458 VPWR.n1773 0 0.106f
C28459 VPWR.n1774 0 0.0014f
C28460 VPWR.n1775 0 0.0014f
C28461 VPWR.n1776 0 0.37f
C28462 VPWR.n1777 0 0.014f
C28463 VPWR.n1778 0 0.00461f
C28464 VPWR.n1779 0 0.00323f
C28465 VPWR.n1780 0 0.00208f
C28466 VPWR.n1782 0 0.00302f
C28467 VPWR.n1783 0 0.00248f
C28468 VPWR.n1784 0 0.00173f
C28469 VPWR.n1785 0 0.00162f
C28470 VPWR.n1786 0 0.00302f
C28471 VPWR.n1788 0 0.00259f
C28472 VPWR.n1789 0 0.0027f
C28473 VPWR.n1790 0 0.00248f
C28474 VPWR.n1791 0 0.00205f
C28475 VPWR.n1792 0 0.00162f
C28476 VPWR.n1793 0 0.00335f
C28477 VPWR.n1794 0 0.00421f
C28478 VPWR.n1795 0 0.00248f
C28479 VPWR.n1796 0 7.56e-19
C28480 VPWR.n1797 0 8.64e-19
C28481 VPWR.n1798 0 0.00108f
C28482 VPWR.n1799 0 0.00205f
C28483 VPWR.n1800 0 0.00248f
C28484 VPWR.n1801 0 0.0027f
C28485 VPWR.n1802 0 0.00302f
C28486 VPWR.n1803 0 0.00184f
C28487 VPWR.n1804 0 9.72e-19
C28488 VPWR.n1805 0 0.0014f
C28489 VPWR.n1806 0 8.64e-19
C28490 VPWR.n1807 0 0.00108f
C28491 VPWR.n1808 0 0.00248f
C28492 VPWR.n1809 0 0.00389f
C28493 VPWR.n1810 0 0.00357f
C28494 VPWR.n1811 0 0.00281f
C28495 VPWR.t84 0 0.073f
C28496 VPWR.n1812 0 0.207f
C28497 VPWR.t194 0 0.073f
C28498 VPWR.n1813 0 0.207f
C28499 VPWR.n1814 0 0.0647f
C28500 VPWR.n1815 0 0.0475f
C28501 VPWR.t345 0 0.0724f
C28502 VPWR.n1816 0 0.00463f
C28503 VPWR.t205 0 0.0951f
C28504 VPWR.n1817 0 0.259f
C28505 VPWR.n1818 0 0.0882f
C28506 VPWR.n1819 0 0.00918f
C28507 VPWR.t361 0 0.0954f
C28508 VPWR.n1820 0 0.332f
C28509 VPWR.n1821 0 0.01f
C28510 VPWR.n1822 0 0.0266f
C28511 VPWR.n1823 0 0.00313f
C28512 VPWR.n1824 0 0.00397f
C28513 VPWR.n1825 0 0.00151f
C28514 VPWR.n1826 0 0.011f
C28515 VPWR.n1827 0 0.00162f
C28516 VPWR.n1828 0 0.00119f
C28517 VPWR.n1829 0 0.00184f
C28518 VPWR.n1830 0 0.00259f
C28519 VPWR.n1831 0 0.00119f
C28520 VPWR.n1832 0 0.00421f
C28521 VPWR.n1833 0 0.00248f
C28522 VPWR.n1834 0 5.4e-19
C28523 VPWR.n1835 0 0.00497f
C28524 VPWR.n1836 0 0.00258f
C28525 VPWR.n1837 0 0.00208f
C28526 VPWR.n1838 0 0.00493f
C28527 VPWR.n1839 0 0.00851f
C28528 VPWR.n1840 0 0.00994f
C28529 VPWR.n1841 0 0.0963f
C28530 VPWR.n1842 0 0.0973f
C28531 VPWR.n1843 0 0.0987f
C28532 VPWR.n1844 0 0.108f
C28533 VPWR.t137 0 0.0774f
C28534 VPWR.t163 0 0.0417f
C28535 VPWR.t131 0 0.0417f
C28536 VPWR.n1845 0 0.383f
C28537 VPWR.n1846 0 0.0384f
C28538 VPWR.n1847 0 0.0421f
C28539 VPWR.t241 0 0.0774f
C28540 VPWR.n1848 0 0.501f
C28541 VPWR.n1849 0 0.0897f
C28542 VPWR.n1850 0 0.018f
C28543 VPWR.n1851 0 0.00429f
C28544 VPWR.n1852 0 0.0199f
C28545 VPWR.n1853 0 0.0118f
C28546 VPWR.n1854 0 0.0189f
C28547 VPWR.n1855 0 0.0729f
C28548 VPWR.n1856 0 0.0844f
C28549 VPWR.n1857 0 0.018f
C28550 VPWR.t154 0 0.0876f
C28551 VPWR.t240 0 0.1f
C28552 VPWR.n1858 0 0.113f
C28553 VPWR.n1859 0 0.0978f
C28554 VPWR.n1860 0 0.146f
C28555 VPWR.n1861 0 0.0199f
C28556 VPWR.n1862 0 0.0199f
C28557 VPWR.n1863 0 0.0199f
C28558 VPWR.n1864 0 0.0199f
C28559 VPWR.n1865 0 0.0118f
C28560 VPWR.n1866 0 0.15f
C28561 VPWR.n1867 0 0.0224f
C28562 VPWR.n1868 0 0.0809f
C28563 VPWR.n1869 0 0.018f
C28564 VPWR.n1870 0 0.0316f
C28565 VPWR.n1871 0 0.0199f
C28566 VPWR.n1872 0 0.0159f
C28567 VPWR.n1873 0 0.0199f
C28568 VPWR.n1874 0 0.0341f
C28569 VPWR.n1875 0 0.0199f
C28570 VPWR.n1876 0 0.0117f
C28571 VPWR.n1877 0 0.0051f
C28572 VPWR.n1878 0 0.049f
C28573 VPWR.n1879 0 0.0181f
C28574 VPWR.t272 0 0.068f
C28575 VPWR.n1880 0 0.0701f
C28576 VPWR.n1881 0 0.0391f
C28577 VPWR.n1882 0 0.0199f
C28578 VPWR.n1883 0 0.0494f
C28579 VPWR.n1884 0 0.0706f
C28580 VPWR.n1885 0 0.0186f
C28581 VPWR.n1886 0 0.00994f
C28582 VPWR.n1887 0 0.00184f
C28583 VPWR.n1888 0 0.015f
C28584 VPWR.n1889 0 0.017f
C28585 VPWR.n1890 0 7.56e-19
C28586 VPWR.n1891 0 0.00378f
C28587 VPWR.n1892 0 0.00162f
C28588 VPWR.n1893 0 0.00151f
C28589 VPWR.n1894 0 0.0013f
C28590 VPWR.n1895 0 0.0014f
C28591 VPWR.n1896 0 0.00259f
C28592 VPWR.n1897 0 0.00162f
C28593 VPWR.n1898 0 0.00216f
C28594 VPWR.n1899 0 0.00357f
C28595 VPWR.n1900 0 0.00248f
C28596 VPWR.n1901 0 0.0014f
C28597 VPWR.n1902 0 0.00335f
C28598 VPWR.n1903 0 0.00248f
C28599 VPWR.n1904 0 0.0014f
C28600 VPWR.n1905 0 8.64e-19
C28601 VPWR.n1906 0 0.00173f
C28602 VPWR.n1907 0 0.0014f
C28603 VPWR.n1908 0 0.306f
C28604 VPWR.n1909 0 0.0341f
C28605 VPWR.n1910 0 0.00248f
C28606 VPWR.n1911 0 0.00184f
C28607 VPWR.n1912 0 0.0138f
C28608 VPWR.n1913 0 0.00119f
C28609 VPWR.n1914 0 0.00302f
C28610 VPWR.n1915 0 0.00248f
C28611 VPWR.n1916 0 5.4e-19
C28612 VPWR.n1917 0 0.00259f
C28613 VPWR.n1918 0 8.64e-19
C28614 VPWR.n1919 0 0.00227f
C28615 VPWR.n1920 0 0.00248f
C28616 VPWR.n1921 0 0.00248f
C28617 VPWR.n1922 0 0.00194f
C28618 VPWR.n1923 0 0.00184f
C28619 VPWR.n1924 0 0.00259f
C28620 VPWR.n1925 0 0.00119f
C28621 VPWR.n1926 0 0.00258f
C28622 VPWR.n1927 0 0.00208f
C28623 VPWR.n1928 0 0.00497f
C28624 VPWR.n1929 0 0.00891f
C28625 VPWR.n1930 0 0.00616f
C28626 VPWR.t346 0 0.068f
C28627 VPWR.n1931 0 0.0266f
C28628 VPWR.n1932 0 0.0649f
C28629 VPWR.n1933 0 0.0391f
C28630 VPWR.n1934 0 0.0159f
C28631 VPWR.n1935 0 0.0535f
C28632 VPWR.n1936 0 0.0199f
C28633 VPWR.n1937 0 0.0118f
C28634 VPWR.n1938 0 0.0631f
C28635 VPWR.n1939 0 0.0287f
C28636 VPWR.n1940 0 0.00386f
C28637 VPWR.n1941 0 0.0179f
C28638 VPWR.n1942 0 0.0657f
C28639 VPWR.n1943 0 0.0199f
C28640 VPWR.n1944 0 0.0125f
C28641 VPWR.n1945 0 0.0378f
C28642 VPWR.n1946 0 0.0337f
C28643 VPWR.n1947 0 0.0107f
C28644 VPWR.n1948 0 0.0265f
C28645 VPWR.n1949 0 0.0118f
C28646 VPWR.n1950 0 0.018f
C28647 VPWR.n1951 0 0.0454f
C28648 VPWR.n1952 0 0.0634f
C28649 VPWR.n1953 0 0.00617f
C28650 VPWR.n1954 0 0.018f
C28651 VPWR.n1955 0 0.0626f
C28652 VPWR.n1956 0 0.0199f
C28653 VPWR.n1957 0 0.0049f
C28654 VPWR.n1958 0 0.0199f
C28655 VPWR.n1959 0 0.0688f
C28656 VPWR.n1960 0 0.0199f
C28657 VPWR.n1961 0 0.0657f
C28658 VPWR.n1962 0 0.0199f
C28659 VPWR.n1963 0 0.0117f
C28660 VPWR.n1964 0 0.0143f
C28661 VPWR.n1965 0 0.104f
C28662 VPWR.n1966 0 0.207f
C28663 VPWR.n1967 0 0.0429f
C28664 VPWR.n1968 0 0.0145f
C28665 VPWR.n1969 0 0.00994f
C28666 VPWR.n1970 0 0.00994f
C28667 VPWR.t153 0 0.068f
C28668 VPWR.n1971 0 0.0785f
C28669 VPWR.n1972 0 0.051f
C28670 VPWR.n1973 0 0.0535f
C28671 VPWR.t375 0 0.107f
C28672 VPWR.n1974 0 0.185f
C28673 VPWR.n1975 0 0.0386f
C28674 VPWR.n1976 0 0.0819f
C28675 VPWR.n1977 0 0.0674f
C28676 VPWR.n1978 0 0.0135f
C28677 VPWR.n1979 0 0.0107f
C28678 VPWR.n1980 0 0.115f
C28679 VPWR.n1981 0 0.0528f
C28680 VPWR.n1982 0 0.0118f
C28681 VPWR.n1983 0 0.0199f
C28682 VPWR.n1984 0 0.0199f
C28683 VPWR.n1985 0 0.0452f
C28684 VPWR.n1986 0 0.0199f
C28685 VPWR.n1987 0 0.0172f
C28686 VPWR.n1988 0 0.0794f
C28687 VPWR.n1989 0 0.00655f
C28688 VPWR.n1990 0 0.0126f
C28689 VPWR.n1991 0 0.00704f
C28690 VPWR.n1992 0 0.0199f
C28691 VPWR.n1993 0 0.00933f
C28692 VPWR.n1994 0 0.0199f
C28693 VPWR.n1995 0 0.0589f
C28694 VPWR.n1996 0 0.0199f
C28695 VPWR.n1997 0 0.0426f
C28696 VPWR.n1998 0 0.0199f
C28697 VPWR.n1999 0 0.018f
C28698 VPWR.n2000 0 0.0199f
C28699 VPWR.n2001 0 0.0522f
C28700 VPWR.n2002 0 0.0199f
C28701 VPWR.n2003 0 0.0106f
C28702 VPWR.n2004 0 0.0199f
C28703 VPWR.n2005 0 0.00704f
C28704 VPWR.n2006 0 0.0199f
C28705 VPWR.n2007 0 0.0106f
C28706 VPWR.n2008 0 0.0199f
C28707 VPWR.n2009 0 0.0522f
C28708 VPWR.n2010 0 0.0199f
C28709 VPWR.n2011 0 0.018f
C28710 VPWR.n2012 0 0.0199f
C28711 VPWR.n2013 0 0.0426f
C28712 VPWR.n2014 0 0.0199f
C28713 VPWR.n2015 0 0.0593f
C28714 VPWR.n2016 0 0.0199f
C28715 VPWR.n2017 0 0.018f
C28716 VPWR.n2018 0 0.00839f
C28717 VPWR.n2019 0 0.0634f
C28718 VPWR.n2020 0 0.0118f
C28719 VPWR.n2021 0 0.0199f
C28720 VPWR.n2022 0 0.0199f
C28721 VPWR.n2023 0 0.0173f
C28722 VPWR.n2024 0 0.0107f
C28723 VPWR.n2025 0 0.0375f
C28724 VPWR.n2026 0 0.307f
C28725 VPWR.n2027 0 0.13f
C28726 VPWR.n2028 0 0.0647f
C28727 VPWR.n2029 0 0.00265f
C28728 VPWR.n2030 0 0.00284f
C28729 VPWR.n2031 0 0.00499f
C28730 VPWR.n2032 0 0.00281f
C28731 VPWR.n2033 0 0.00313f
C28732 VPWR.n2034 0 0.00989f
C28733 VPWR.n2035 0 0.00496f
C28734 VPWR.n2036 0 0.00208f
C28735 VPWR.n2037 0 0.00257f
C28736 VPWR.n2038 0 0.00203f
C28737 VPWR.n2039 0 0.0173f
C28738 VPWR.n2040 0 0.00248f
C28739 VPWR.n2041 0 0.00344f
C28740 VPWR.n2042 0 0.00323f
C28741 VPWR.n2043 0 0.00208f
C28742 VPWR.n2045 0 0.00329f
C28743 VPWR.n2046 0 0.00208f
C28744 VPWR.n2047 0 0.00481f
C28745 VPWR.n2048 0 0.00329f
C28746 VPWR.n2049 0 0.00208f
C28747 VPWR.n2050 0 0.00302f
C28748 VPWR.n2051 0 0.00248f
C28749 VPWR.n2052 0 0.00173f
C28750 VPWR.n2053 0 8.64e-19
C28751 VPWR.n2054 0 0.00108f
C28752 VPWR.n2055 0 0.00248f
C28753 VPWR.n2056 0 0.00389f
C28754 VPWR.n2057 0 0.00357f
C28755 VPWR.n2058 0 0.00281f
C28756 VPWR.n2059 0 0.00302f
C28757 VPWR.n2060 0 0.00248f
C28758 VPWR.n2061 0 0.00173f
C28759 VPWR.n2062 0 0.0014f
C28760 VPWR.n2063 0 0.00162f
C28761 VPWR.n2064 0 0.00184f
C28762 VPWR.n2065 0 0.0522f
C28763 VPWR.n2066 0 0.0535f
C28764 VPWR.n2067 0 0.0619f
C28765 VPWR.n2068 0 0.0386f
C28766 VPWR.t333 0 0.068f
C28767 VPWR.n2069 0 0.0701f
C28768 VPWR.n2070 0 0.0391f
C28769 VPWR.n2071 0 0.0535f
C28770 VPWR.n2072 0 0.0619f
C28771 VPWR.t362 0 0.068f
C28772 VPWR.n2073 0 0.0701f
C28773 VPWR.n2074 0 0.0391f
C28774 VPWR.n2075 0 0.0535f
C28775 VPWR.n2076 0 0.00994f
C28776 VPWR.n2077 0 0.062f
C28777 VPWR.n2078 0 0.0275f
C28778 VPWR.t314 0 0.068f
C28779 VPWR.n2079 0 0.00482f
C28780 VPWR.n2080 0 0.0329f
C28781 VPWR.n2081 0 0.0665f
C28782 VPWR.n2082 0 0.00482f
C28783 VPWR.n2083 0 0.0213f
C28784 VPWR.n2084 0 0.0221f
C28785 VPWR.n2085 0 0.0179f
C28786 VPWR.n2086 0 0.00259f
C28787 VPWR.n2087 0 0.00421f
C28788 VPWR.n2088 0 0.00378f
C28789 VPWR.n2089 0 0.00162f
C28790 VPWR.n2090 0 0.0014f
C28791 VPWR.n2091 0 0.0027f
C28792 VPWR.n2092 0 0.00248f
C28793 VPWR.n2093 0 0.00205f
C28794 VPWR.n2094 0 0.0027f
C28795 VPWR.n2095 0 0.00248f
C28796 VPWR.n2096 0 0.00205f
C28797 VPWR.n2097 0 0.00108f
C28798 VPWR.n2098 0 8.64e-19
C28799 VPWR.n2099 0 7.56e-19
C28800 VPWR.n2100 0 0.00248f
C28801 VPWR.n2101 0 0.00421f
C28802 VPWR.n2102 0 0.00335f
C28803 VPWR.n2103 0 0.00162f
C28804 VPWR.n2104 0 0.0014f
C28805 VPWR.n2105 0 0.00745f
C28806 VPWR.n2106 0 0.00259f
C28807 VPWR.n2107 0 0.00259f
C28808 VPWR.n2108 0 0.00292f
C28809 VPWR.n2109 0 0.00184f
C28810 VPWR.n2110 0 0.00994f
C28811 VPWR.n2111 0 0.0115f
C28812 VPWR.n2112 0 0.0611f
C28813 VPWR.n2113 0 0.0457f
C28814 VPWR.n2114 0 0.018f
C28815 VPWR.n2115 0 0.00429f
C28816 VPWR.n2116 0 0.0199f
C28817 VPWR.n2117 0 0.0199f
C28818 VPWR.n2118 0 0.00529f
C28819 VPWR.t347 0 0.068f
C28820 VPWR.n2119 0 0.0535f
C28821 VPWR.n2120 0 0.0391f
C28822 VPWR.n2121 0 0.0701f
C28823 VPWR.n2122 0 0.049f
C28824 VPWR.n2123 0 0.018f
C28825 VPWR.n2124 0 0.0199f
C28826 VPWR.n2125 0 0.0199f
C28827 VPWR.n2126 0 0.0118f
C28828 VPWR.n2127 0 0.0623f
C28829 VPWR.n2128 0 0.0555f
C28830 VPWR.n2129 0 0.00513f
C28831 VPWR.n2130 0 0.018f
C28832 VPWR.n2131 0 0.0533f
C28833 VPWR.n2132 0 0.0199f
C28834 VPWR.t5 0 0.068f
C28835 VPWR.n2133 0 0.0701f
C28836 VPWR.n2134 0 0.0482f
C28837 VPWR.n2135 0 0.0199f
C28838 VPWR.n2136 0 0.0391f
C28839 VPWR.n2137 0 0.0199f
C28840 VPWR.n2138 0 0.0535f
C28841 VPWR.n2139 0 0.0199f
C28842 VPWR.n2140 0 0.0619f
C28843 VPWR.n2141 0 0.0118f
C28844 VPWR.n2142 0 0.00994f
C28845 VPWR.n2143 0 0.0687f
C28846 VPWR.n2144 0 0.018f
C28847 VPWR.n2145 0 0.00631f
C28848 VPWR.n2146 0 0.0199f
C28849 VPWR.n2147 0 0.0464f
C28850 VPWR.n2148 0 0.0199f
C28851 VPWR.n2149 0 0.00533f
C28852 VPWR.n2150 0 0.0199f
C28853 VPWR.n2151 0 0.049f
C28854 VPWR.n2152 0 0.0199f
C28855 VPWR.n2153 0 0.0199f
C28856 VPWR.n2154 0 0.0199f
C28857 VPWR.t29 0 0.068f
C28858 VPWR.n2155 0 0.0701f
C28859 VPWR.n2156 0 0.0391f
C28860 VPWR.n2157 0 0.0535f
C28861 VPWR.n2158 0 0.0619f
C28862 VPWR.n2159 0 0.0118f
C28863 VPWR.n2160 0 0.0107f
C28864 VPWR.n2161 0 0.0475f
C28865 VPWR.n2162 0 0.0173f
C28866 VPWR.n2163 0 0.0199f
C28867 VPWR.n2164 0 0.0199f
C28868 VPWR.n2165 0 0.0118f
C28869 VPWR.n2166 0 0.0634f
C28870 VPWR.n2167 0 0.00521f
C28871 VPWR.n2168 0 0.018f
C28872 VPWR.n2169 0 0.0516f
C28873 VPWR.n2170 0 0.0199f
C28874 VPWR.n2171 0 0.028f
C28875 VPWR.n2172 0 0.0199f
C28876 VPWR.n2173 0 0.0061f
C28877 VPWR.n2174 0 0.0199f
C28878 VPWR.n2175 0 0.0341f
C28879 VPWR.n2176 0 0.0199f
C28880 VPWR.n2177 0 0.00559f
C28881 VPWR.n2178 0 0.0199f
C28882 VPWR.n2179 0 0.00704f
C28883 VPWR.n2180 0 0.0199f
C28884 VPWR.n2181 0 0.00677f
C28885 VPWR.n2182 0 0.0199f
C28886 VPWR.n2183 0 0.0449f
C28887 VPWR.n2184 0 0.0199f
C28888 VPWR.n2185 0 0.00448f
C28889 VPWR.n2186 0 0.0199f
C28890 VPWR.n2187 0 0.0233f
C28891 VPWR.n2188 0 0.0199f
C28892 VPWR.n2189 0 0.0162f
C28893 VPWR.n2190 0 0.0199f
C28894 VPWR.n2191 0 0.00704f
C28895 VPWR.n2192 0 0.0199f
C28896 VPWR.n2193 0 0.00704f
C28897 VPWR.n2194 0 0.0199f
C28898 VPWR.n2195 0 0.00681f
C28899 VPWR.n2196 0 0.0199f
C28900 VPWR.n2197 0 0.0291f
C28901 VPWR.n2198 0 0.0199f
C28902 VPWR.n2199 0 0.00536f
C28903 VPWR.n2200 0 0.0199f
C28904 VPWR.n2201 0 0.00585f
C28905 VPWR.n2202 0 0.0199f
C28906 VPWR.n2203 0 0.04f
C28907 VPWR.n2204 0 0.0199f
C28908 VPWR.n2205 0 0.0118f
C28909 VPWR.n2206 0 0.00521f
C28910 VPWR.n2207 0 0.049f
C28911 VPWR.n2208 0 0.018f
C28912 VPWR.n2209 0 0.0199f
C28913 VPWR.n2210 0 0.0199f
C28914 VPWR.n2211 0 0.0118f
C28915 VPWR.n2212 0 0.00497f
C28916 VPWR.n2213 0 0.381f
C28917 VPWR.n2214 0 0.00208f
C28918 VPWR.n2215 0 0.00323f
C28919 VPWR.n2216 0 0.00468f
C28920 VPWR.n2217 0 0.00323f
C28921 VPWR.n2218 0 0.00248f
C28922 VPWR.n2219 0 0.00344f
C28923 VPWR.n2220 0 0.00208f
C28924 VPWR.n2222 0 0.00329f
C28925 VPWR.n2223 0 0.00208f
C28926 VPWR.n2224 0 0.00302f
C28927 VPWR.n2225 0 0.00248f
C28928 VPWR.n2226 0 0.00173f
C28929 VPWR.n2227 0 0.014f
C28930 VPWR.n2228 0 0.00194f
C28931 VPWR.n2229 0 0.0013f
C28932 VPWR.n2230 0 0.00108f
C28933 VPWR.n2231 0 0.00194f
C28934 VPWR.n2232 0 0.00173f
C28935 VPWR.n2233 0 0.0014f
C28936 VPWR.n2234 0 8.64e-19
C28937 VPWR.n2235 0 0.00108f
C28938 VPWR.n2236 0 0.00248f
C28939 VPWR.n2237 0 0.00378f
C28940 VPWR.n2238 0 0.00194f
C28941 VPWR.n2239 0 0.00173f
C28942 VPWR.n2240 0 0.0027f
C28943 VPWR.n2241 0 0.00119f
C28944 VPWR.n2242 0 0.00486f
C28945 VPWR.n2243 0 0.00389f
C28946 VPWR.n2244 0 0.00173f
C28947 VPWR.n2245 0 0.0027f
C28948 VPWR.t17 0 0.068f
C28949 VPWR.n2246 0 0.00482f
C28950 VPWR.n2247 0 0.0329f
C28951 VPWR.n2248 0 0.0665f
C28952 VPWR.n2249 0 0.0261f
C28953 VPWR.n2250 0 0.0179f
C28954 VPWR.n2251 0 0.00119f
C28955 VPWR.n2252 0 0.062f
C28956 VPWR.n2253 0 0.0482f
C28957 VPWR.n2254 0 0.0413f
C28958 VPWR.t6 0 0.0592f
C28959 VPWR.n2255 0 0.0227f
C28960 VPWR.n2256 0 0.0865f
C28961 VPWR.n2257 0 0.0369f
C28962 VPWR.n2258 0 0.0413f
C28963 VPWR.n2259 0 0.0462f
C28964 VPWR.n2260 0 0.062f
C28965 VPWR.n2261 0 0.0457f
C28966 VPWR.t62 0 0.0336f
C28967 VPWR.n2262 0 0.0983f
C28968 VPWR.n2263 0 0.0651f
C28969 VPWR.n2264 0 0.023f
C28970 VPWR.n2265 0 0.0393f
C28971 VPWR.n2266 0 0.0629f
C28972 VPWR.n2267 0 0.0118f
C28973 VPWR.n2268 0 0.0535f
C28974 VPWR.n2269 0 0.0199f
C28975 VPWR.n2270 0 0.0522f
C28976 VPWR.n2271 0 0.0199f
C28977 VPWR.n2272 0 0.0522f
C28978 VPWR.n2273 0 0.0199f
C28979 VPWR.t255 0 0.0876f
C28980 VPWR.n2274 0 0.149f
C28981 VPWR.n2275 0 0.0199f
C28982 VPWR.n2276 0 0.062f
C28983 VPWR.n2277 0 0.0199f
C28984 VPWR.n2278 0 0.0199f
C28985 VPWR.n2279 0 0.00429f
C28986 VPWR.n2280 0 0.0199f
C28987 VPWR.n2281 0 0.018f
C28988 VPWR.n2282 0 0.00529f
C28989 VPWR.n2283 0 0.0634f
C28990 VPWR.n2284 0 0.0118f
C28991 VPWR.n2285 0 0.0535f
C28992 VPWR.n2286 0 0.0199f
C28993 VPWR.n2287 0 0.0522f
C28994 VPWR.n2288 0 0.0199f
C28995 VPWR.n2289 0 0.0513f
C28996 VPWR.n2290 0 0.0199f
C28997 VPWR.n2291 0 0.0363f
C28998 VPWR.n2292 0 0.0199f
C28999 VPWR.n2293 0 0.0199f
C29000 VPWR.n2294 0 0.0199f
C29001 VPWR.n2295 0 0.018f
C29002 VPWR.n2296 0 0.07f
C29003 VPWR.n2297 0 0.00526f
C29004 VPWR.n2298 0 0.0199f
C29005 VPWR.n2299 0 0.00429f
C29006 VPWR.n2300 0 0.0199f
C29007 VPWR.n2301 0 0.018f
C29008 VPWR.n2302 0 0.0457f
C29009 VPWR.n2303 0 0.062f
C29010 VPWR.n2304 0 0.0118f
C29011 VPWR.n2305 0 0.0487f
C29012 VPWR.n2306 0 0.018f
C29013 VPWR.n2307 0 0.00983f
C29014 VPWR.n2308 0 0.00184f
C29015 VPWR.n2309 0 0.00882f
C29016 VPWR.n2310 0 0.00496f
C29017 VPWR.n2311 0 0.0216f
C29018 VPWR.n2312 0 0.0173f
C29019 VPWR.n2314 0 0.00344f
C29020 VPWR.n2315 0 0.00248f
C29021 VPWR.n2316 0 0.00329f
C29022 VPWR.n2317 0 0.00208f
C29023 VPWR.n2318 0 0.00496f
C29024 VPWR.n2319 0 0.00859f
C29025 VPWR.n2320 0 0.00443f
C29026 VPWR.n2321 0 0.00281f
C29027 VPWR.n2322 0 0.00367f
C29028 VPWR.n2323 0 0.00281f
C29029 VPWR.n2324 0 0.00238f
C29030 VPWR.n2325 0 8.64e-19
C29031 VPWR.n2326 0 0.00302f
C29032 VPWR.n2327 0 0.00443f
C29033 VPWR.n2328 0 0.00205f
C29034 VPWR.n2329 0 0.00162f
C29035 VPWR.n2330 0 0.0027f
C29036 VPWR.n2331 0 0.0013f
C29037 VPWR.n2332 0 0.0013f
C29038 VPWR.n2333 0 0.0027f
C29039 VPWR.n2334 0 0.00162f
C29040 VPWR.n2335 0 0.00164f
C29041 VPWR.n2336 0 0.00212f
C29042 VPWR.n2337 0 0.038f
C29043 VPWR.n2338 0 0.18f
C29044 VPWR.n2339 0 0.18f
C29045 VPWR.n2340 0 0.18f
C29046 VPWR.t299 0 0.068f
C29047 VPWR.n2341 0 0.0701f
C29048 VPWR.n2342 0 0.0391f
C29049 VPWR.n2343 0 0.0535f
C29050 VPWR.n2344 0 0.0634f
C29051 VPWR.n2345 0 0.0634f
C29052 VPWR.n2346 0 0.0619f
C29053 VPWR.n2347 0 0.18f
C29054 VPWR.n2348 0 0.0634f
C29055 VPWR.n2349 0 0.062f
C29056 VPWR.n2350 0 0.0276f
C29057 VPWR.n2351 0 0.00378f
C29058 VPWR.n2352 0 0.00248f
C29059 VPWR.n2353 0 5.4e-19
C29060 VPWR.n2354 0 0.00259f
C29061 VPWR.n2355 0 0.00313f
C29062 VPWR.n2356 0 0.00151f
C29063 VPWR.n2357 0 0.00162f
C29064 VPWR.n2358 0 0.00119f
C29065 VPWR.n2359 0 0.00184f
C29066 VPWR.n2360 0 0.00259f
C29067 VPWR.n2361 0 0.00119f
C29068 VPWR.n2362 0 0.00421f
C29069 VPWR.n2363 0 0.00248f
C29070 VPWR.n2364 0 5.4e-19
C29071 VPWR.n2365 0 8.64e-19
C29072 VPWR.n2366 0 0.00227f
C29073 VPWR.n2367 0 0.00248f
C29074 VPWR.n2368 0 0.00248f
C29075 VPWR.n2369 0 0.00194f
C29076 VPWR.n2370 0 0.00184f
C29077 VPWR.n2371 0 0.00259f
C29078 VPWR.n2372 0 0.00119f
C29079 VPWR.n2373 0 0.00344f
C29080 VPWR.n2374 0 0.00248f
C29081 VPWR.n2375 0 0.00329f
C29082 VPWR.n2376 0 0.00208f
C29083 VPWR.n2377 0 0.381f
C29084 VPWR.n2378 0 0.381f
C29085 VPWR.n2379 0 0.00335f
C29086 VPWR.n2380 0 0.00248f
C29087 VPWR.n2381 0 0.0014f
C29088 VPWR.n2382 0 8.64e-19
C29089 VPWR.n2383 0 0.0014f
C29090 VPWR.n2384 0 0.00248f
C29091 VPWR.n2385 0 0.00357f
C29092 VPWR.n2386 0 0.00216f
C29093 VPWR.n2387 0 0.00162f
C29094 VPWR.n2388 0 0.00259f
C29095 VPWR.n2389 0 0.0522f
C29096 VPWR.n2390 0 0.0535f
C29097 VPWR.n2391 0 0.0619f
C29098 VPWR.n2392 0 0.18f
C29099 VPWR.n2393 0 0.062f
C29100 VPWR.t242 0 0.068f
C29101 VPWR.n2394 0 0.0701f
C29102 VPWR.n2395 0 0.0391f
C29103 VPWR.n2396 0 0.0535f
C29104 VPWR.n2397 0 0.062f
C29105 VPWR.t215 0 0.068f
C29106 VPWR.n2398 0 0.0701f
C29107 VPWR.n2399 0 0.0391f
C29108 VPWR.n2400 0 0.0535f
C29109 VPWR.n2401 0 0.0552f
C29110 VPWR.t73 0 0.0336f
C29111 VPWR.n2402 0 0.0984f
C29112 VPWR.n2403 0 0.0393f
C29113 VPWR.n2404 0 0.0237f
C29114 VPWR.n2405 0 0.0485f
C29115 VPWR.n2406 0 0.0199f
C29116 VPWR.n2407 0 0.0199f
C29117 VPWR.n2408 0 0.0199f
C29118 VPWR.n2409 0 0.0118f
C29119 VPWR.n2410 0 0.062f
C29120 VPWR.n2411 0 0.0457f
C29121 VPWR.n2412 0 0.018f
C29122 VPWR.n2413 0 0.00429f
C29123 VPWR.n2414 0 0.0199f
C29124 VPWR.n2415 0 0.0199f
C29125 VPWR.n2416 0 0.00529f
C29126 VPWR.n2417 0 0.049f
C29127 VPWR.n2418 0 0.018f
C29128 VPWR.n2419 0 0.0199f
C29129 VPWR.n2420 0 0.0199f
C29130 VPWR.n2421 0 0.0118f
C29131 VPWR.n2422 0 0.062f
C29132 VPWR.n2423 0 0.0457f
C29133 VPWR.n2424 0 0.018f
C29134 VPWR.n2425 0 0.00429f
C29135 VPWR.n2426 0 0.0199f
C29136 VPWR.n2427 0 0.0199f
C29137 VPWR.n2428 0 0.00529f
C29138 VPWR.n2429 0 0.0634f
C29139 VPWR.n2430 0 0.018f
C29140 VPWR.t258 0 0.0876f
C29141 VPWR.n2431 0 0.149f
C29142 VPWR.n2432 0 0.0199f
C29143 VPWR.n2433 0 0.0522f
C29144 VPWR.n2434 0 0.0199f
C29145 VPWR.n2435 0 0.0199f
C29146 VPWR.n2436 0 0.0199f
C29147 VPWR.n2437 0 0.0118f
C29148 VPWR.n2438 0 0.0107f
C29149 VPWR.n2439 0 0.038f
C29150 VPWR.n2440 0 0.014f
C29151 VPWR.n2441 0 0.00735f
C29152 VPWR.n2442 0 0.00184f
C29153 VPWR.n2443 0 0.00482f
C29154 VPWR.n2444 0 0.0329f
C29155 VPWR.n2445 0 7.56e-19
C29156 VPWR.n2446 0 0.00194f
C29157 VPWR.n2447 0 0.00184f
C29158 VPWR.t206 0 0.068f
C29159 VPWR.n2448 0 0.0665f
C29160 VPWR.n2449 0 0.00425f
C29161 VPWR.n2450 0 0.00397f
C29162 VPWR.n2451 0 0.0196f
C29163 VPWR.n2452 0 0.0221f
C29164 VPWR.n2453 0 0.0179f
C29165 VPWR.n2454 0 0.00248f
C29166 VPWR.n2455 0 0.0014f
C29167 VPWR.n2456 0 0.00173f
C29168 VPWR.n2457 0 0.00497f
C29169 VPWR.n2458 0 0.00378f
C29170 VPWR.n2459 0 0.00162f
C29171 VPWR.n2460 0 0.00259f
C29172 VPWR.n2461 0 0.0014f
C29173 VPWR.n2462 0 0.0014f
C29174 VPWR.n2463 0 0.0085f
C29175 VPWR.n2464 0 0.00495f
C29176 VPWR.n2465 0 0.00248f
C29177 VPWR.n2466 0 0.00329f
C29178 VPWR.n2467 0 0.00208f
C29179 VPWR.n2469 0 0.00344f
C29180 VPWR.n2470 0 0.00208f
C29181 VPWR.n2471 0 0.00323f
C29182 VPWR.n2472 0 0.00468f
C29183 VPWR.n2473 0 0.00323f
C29184 VPWR.n2474 0 0.00208f
C29185 VPWR.n2475 0 0.0173f
C29186 VPWR.n2477 0 0.0217f
C29187 VPWR.n2478 0 0.00496f
C29188 VPWR.n2479 0 0.00892f
C29189 VPWR.n2480 0 0.00616f
C29190 VPWR.n2481 0 0.00778f
C29191 VPWR.n2482 0 0.0593f
C29192 VPWR.n2483 0 0.0457f
C29193 VPWR.n2484 0 0.018f
C29194 VPWR.n2485 0 0.00429f
C29195 VPWR.n2486 0 0.0199f
C29196 VPWR.n2487 0 0.0199f
C29197 VPWR.n2488 0 0.00525f
C29198 VPWR.t273 0 0.0949f
C29199 VPWR.n2489 0 0.101f
C29200 VPWR.n2490 0 0.0331f
C29201 VPWR.n2491 0 0.0369f
C29202 VPWR.n2492 0 0.0425f
C29203 VPWR.n2493 0 0.0457f
C29204 VPWR.n2494 0 0.0487f
C29205 VPWR.n2495 0 0.071f
C29206 VPWR.n2496 0 0.018f
C29207 VPWR.n2497 0 0.0199f
C29208 VPWR.n2498 0 0.0199f
C29209 VPWR.n2499 0 0.0513f
C29210 VPWR.n2500 0 0.0199f
C29211 VPWR.n2501 0 0.0214f
C29212 VPWR.n2502 0 0.0369f
C29213 VPWR.n2503 0 0.0513f
C29214 VPWR.n2504 0 0.0199f
C29215 VPWR.n2505 0 0.0475f
C29216 VPWR.n2506 0 0.0369f
C29217 VPWR.n2507 0 0.0367f
C29218 VPWR.n2508 0 0.0199f
C29219 VPWR.n2509 0 0.0513f
C29220 VPWR.n2510 0 0.0199f
C29221 VPWR.n2511 0 0.0522f
C29222 VPWR.n2512 0 0.0199f
C29223 VPWR.n2513 0 0.0522f
C29224 VPWR.n2514 0 0.0199f
C29225 VPWR.n2515 0 0.0522f
C29226 VPWR.n2516 0 0.0199f
C29227 VPWR.n2517 0 0.0535f
C29228 VPWR.n2518 0 0.0199f
C29229 VPWR.n2519 0 0.0118f
C29230 VPWR.n2520 0 0.00529f
C29231 VPWR.n2521 0 0.062f
C29232 VPWR.n2522 0 0.018f
C29233 VPWR.n2523 0 0.00429f
C29234 VPWR.n2524 0 0.0199f
C29235 VPWR.n2525 0 0.0457f
C29236 VPWR.n2526 0 0.0199f
C29237 VPWR.t313 0 0.068f
C29238 VPWR.n2527 0 0.0701f
C29239 VPWR.n2528 0 0.0476f
C29240 VPWR.n2529 0 0.0199f
C29241 VPWR.n2530 0 0.0391f
C29242 VPWR.n2531 0 0.0199f
C29243 VPWR.n2532 0 0.0535f
C29244 VPWR.n2533 0 0.0199f
C29245 VPWR.n2534 0 0.0118f
C29246 VPWR.n2535 0 0.0107f
C29247 VPWR.n2536 0 0.0386f
C29248 VPWR.t243 0 0.068f
C29249 VPWR.n2537 0 0.0535f
C29250 VPWR.n2538 0 0.0391f
C29251 VPWR.n2539 0 0.0701f
C29252 VPWR.n2540 0 0.0475f
C29253 VPWR.n2541 0 0.0173f
C29254 VPWR.n2542 0 0.0199f
C29255 VPWR.n2543 0 0.0199f
C29256 VPWR.n2544 0 0.0118f
C29257 VPWR.n2545 0 0.00994f
C29258 VPWR.n2546 0 0.00368f
C29259 VPWR.n2547 0 0.0521f
C29260 VPWR.n2548 0 0.018f
C29261 VPWR.n2549 0 0.00529f
C29262 VPWR.n2550 0 0.0199f
C29263 VPWR.n2551 0 0.049f
C29264 VPWR.n2552 0 0.0199f
C29265 VPWR.n2553 0 0.0199f
C29266 VPWR.n2554 0 0.0199f
C29267 VPWR.n2555 0 0.0118f
C29268 VPWR.n2556 0 0.00994f
C29269 VPWR.n2557 0 0.00655f
C29270 VPWR.n2558 0 0.00704f
C29271 VPWR.n2559 0 0.018f
C29272 VPWR.n2560 0 0.00566f
C29273 VPWR.n2561 0 0.0199f
C29274 VPWR.n2562 0 0.0127f
C29275 VPWR.n2563 0 0.0199f
C29276 VPWR.n2564 0 0.00513f
C29277 VPWR.n2565 0 0.0199f
C29278 VPWR.n2566 0 0.0544f
C29279 VPWR.n2567 0 0.0199f
C29280 VPWR.n2568 0 0.0057f
C29281 VPWR.n2569 0 0.0199f
C29282 VPWR.n2570 0 0.00704f
C29283 VPWR.n2571 0 0.0199f
C29284 VPWR.n2572 0 0.0126f
C29285 VPWR.n2573 0 0.00652f
C29286 VPWR.n2574 0 0.07f
C29287 VPWR.n2575 0 0.0172f
C29288 VPWR.n2576 0 0.0462f
C29289 VPWR.n2577 0 0.0413f
C29290 VPWR.n2578 0 0.0199f
C29291 VPWR.t377 0 0.0592f
C29292 VPWR.n2579 0 0.0227f
C29293 VPWR.n2580 0 0.0865f
C29294 VPWR.n2581 0 0.0369f
C29295 VPWR.n2582 0 0.0413f
C29296 VPWR.n2583 0 0.0199f
C29297 VPWR.n2584 0 0.0482f
C29298 VPWR.n2585 0 0.0363f
C29299 VPWR.n2586 0 0.0199f
C29300 VPWR.n2587 0 0.0513f
C29301 VPWR.n2588 0 0.0199f
C29302 VPWR.n2589 0 0.0199f
C29303 VPWR.n2590 0 0.0199f
C29304 VPWR.n2591 0 0.0118f
C29305 VPWR.n2592 0 0.0107f
C29306 VPWR.n2593 0 0.038f
C29307 VPWR.n2594 0 0.014f
C29308 VPWR.n2595 0 0.00335f
C29309 VPWR.n2596 0 0.00367f
C29310 VPWR.n2597 0 0.00281f
C29311 VPWR.n2598 0 0.00238f
C29312 VPWR.n2599 0 0.0099f
C29313 VPWR.n2600 0 0.00496f
C29314 VPWR.n2601 0 0.0216f
C29315 VPWR.n2602 0 0.00468f
C29316 VPWR.n2603 0 0.00323f
C29317 VPWR.n2604 0 0.00248f
C29318 VPWR.n2605 0 0.00344f
C29319 VPWR.n2606 0 0.00208f
C29320 VPWR.n2608 0 0.381f
C29321 VPWR.n2609 0 0.381f
C29322 VPWR.n2610 0 0.00323f
C29323 VPWR.n2611 0 0.00248f
C29324 VPWR.n2612 0 0.00344f
C29325 VPWR.n2613 0 0.00208f
C29326 VPWR.n2615 0 0.00329f
C29327 VPWR.n2616 0 0.00208f
C29328 VPWR.n2617 0 0.00481f
C29329 VPWR.n2618 0 0.00329f
C29330 VPWR.n2619 0 0.00208f
C29331 VPWR.n2620 0 0.00302f
C29332 VPWR.n2621 0 0.00248f
C29333 VPWR.n2622 0 0.00173f
C29334 VPWR.n2623 0 0.067f
C29335 VPWR.n2624 0 0.0295f
C29336 VPWR.n2625 0 0.00259f
C29337 VPWR.n2626 0 0.0027f
C29338 VPWR.n2627 0 0.00248f
C29339 VPWR.n2628 0 0.00205f
C29340 VPWR.n2629 0 0.00744f
C29341 VPWR.n2630 0 0.00259f
C29342 VPWR.n2631 0 0.00302f
C29343 VPWR.n2632 0 0.00162f
C29344 VPWR.n2633 0 0.0014f
C29345 VPWR.n2634 0 0.025f
C29346 VPWR.n2635 0 0.0549f
C29347 VPWR.t128 0 0.0854f
C29348 VPWR.n2636 0 0.0688f
C29349 VPWR.n2637 0 0.0565f
C29350 VPWR.n2638 0 0.0522f
C29351 VPWR.n2639 0 0.0386f
C29352 VPWR.n2640 0 0.0595f
C29353 VPWR.n2641 0 0.0443f
C29354 VPWR.n2642 0 0.0341f
C29355 VPWR.t266 0 0.068f
C29356 VPWR.n2643 0 0.0672f
C29357 VPWR.n2644 0 0.0633f
C29358 VPWR.n2645 0 0.0856f
C29359 VPWR.t78 0 0.0711f
C29360 VPWR.n2646 0 0.195f
C29361 VPWR.t211 0 0.068f
C29362 VPWR.n2647 0 0.0701f
C29363 VPWR.n2648 0 0.0391f
C29364 VPWR.n2649 0 0.0877f
C29365 VPWR.n2650 0 0.0658f
C29366 VPWR.n2651 0 0.0189f
C29367 VPWR.t168 0 0.0926f
C29368 VPWR.n2652 0 0.335f
C29369 VPWR.n2653 0 0.111f
C29370 VPWR.n2654 0 0.0531f
C29371 VPWR.n2655 0 0.0118f
C29372 VPWR.n2656 0 0.0199f
C29373 VPWR.n2657 0 0.0199f
C29374 VPWR.n2658 0 0.0608f
C29375 VPWR.n2659 0 0.0199f
C29376 VPWR.n2660 0 0.0487f
C29377 VPWR.n2661 0 0.0199f
C29378 VPWR.n2662 0 0.0199f
C29379 VPWR.n2663 0 0.018f
C29380 VPWR.n2664 0 0.0596f
C29381 VPWR.t280 0 0.094f
C29382 VPWR.n2665 0 0.334f
C29383 VPWR.n2666 0 0.019f
C29384 VPWR.n2667 0 0.0347f
C29385 VPWR.n2668 0 0.00907f
C29386 VPWR.n2669 0 0.0107f
C29387 VPWR.n2670 0 0.0479f
C29388 VPWR.n2671 0 0.0039f
C29389 VPWR.n2672 0 0.0184f
C29390 VPWR.n2673 0 0.185f
C29391 VPWR.n2674 0 0.0265f
C29392 VPWR.n2675 0 0.0727f
C29393 VPWR.n2676 0 0.0265f
C29394 VPWR.n2677 0 0.0376f
C29395 VPWR.n2678 0 0.0199f
C29396 VPWR.n2679 0 0.0057f
C29397 VPWR.n2680 0 0.0199f
C29398 VPWR.n2681 0 0.018f
C29399 VPWR.n2682 0 0.00994f
C29400 VPWR.n2683 0 0.0301f
C29401 VPWR.n2684 0 0.0534f
C29402 VPWR.n2685 0 0.0118f
C29403 VPWR.n2686 0 0.0199f
C29404 VPWR.n2687 0 0.0199f
C29405 VPWR.n2688 0 0.0743f
C29406 VPWR.n2689 0 0.0173f
C29407 VPWR.n2690 0 0.0107f
C29408 VPWR.n2691 0 0.0868f
C29409 VPWR.n2692 0 0.0118f
C29410 VPWR.n2693 0 0.0199f
C29411 VPWR.n2694 0 0.0199f
C29412 VPWR.n2695 0 0.018f
C29413 VPWR.n2696 0 0.0669f
C29414 VPWR.n2697 0 0.0321f
C29415 VPWR.n2698 0 0.0118f
C29416 VPWR.n2699 0 0.0199f
C29417 VPWR.n2700 0 0.00559f
C29418 VPWR.n2701 0 0.0199f
C29419 VPWR.n2702 0 0.00704f
C29420 VPWR.n2703 0 0.0199f
C29421 VPWR.n2704 0 0.00677f
C29422 VPWR.n2705 0 0.0199f
C29423 VPWR.n2706 0 0.0199f
C29424 VPWR.n2707 0 0.0199f
C29425 VPWR.n2708 0 0.0192f
C29426 VPWR.n2709 0 0.0199f
C29427 VPWR.n2710 0 0.0593f
C29428 VPWR.n2711 0 0.0199f
C29429 VPWR.n2712 0 0.00852f
C29430 VPWR.n2713 0 0.0199f
C29431 VPWR.n2714 0 0.018f
C29432 VPWR.n2715 0 0.0509f
C29433 VPWR.n2716 0 0.0627f
C29434 VPWR.n2717 0 0.0118f
C29435 VPWR.n2718 0 0.0695f
C29436 VPWR.n2719 0 0.0199f
C29437 VPWR.n2720 0 0.0433f
C29438 VPWR.n2721 0 0.0199f
C29439 VPWR.t189 0 0.068f
C29440 VPWR.n2722 0 0.0701f
C29441 VPWR.n2723 0 0.0474f
C29442 VPWR.n2724 0 0.0199f
C29443 VPWR.n2725 0 0.018f
C29444 VPWR.n2726 0 0.00994f
C29445 VPWR.n2727 0 0.0527f
C29446 VPWR.n2728 0 0.0627f
C29447 VPWR.n2729 0 0.0118f
C29448 VPWR.n2730 0 0.0199f
C29449 VPWR.n2731 0 0.0199f
C29450 VPWR.n2732 0 0.018f
C29451 VPWR.n2733 0 0.044f
C29452 VPWR.n2734 0 0.0578f
C29453 VPWR.n2735 0 0.0269f
C29454 VPWR.n2736 0 0.00994f
C29455 VPWR.n2737 0 0.0024f
C29456 VPWR.n2738 0 0.0031f
C29457 VPWR.n2739 0 0.00259f
C29458 VPWR.n2740 0 0.00259f
C29459 VPWR.n2741 0 0.0014f
C29460 VPWR.n2742 0 0.00162f
C29461 VPWR.n2743 0 0.00335f
C29462 VPWR.n2744 0 0.00421f
C29463 VPWR.n2745 0 0.00248f
C29464 VPWR.n2746 0 7.56e-19
C29465 VPWR.n2747 0 8.64e-19
C29466 VPWR.n2748 0 0.00108f
C29467 VPWR.n2749 0 0.00205f
C29468 VPWR.n2750 0 0.00248f
C29469 VPWR.n2751 0 0.0027f
C29470 VPWR.n2752 0 0.00302f
C29471 VPWR.n2753 0 0.00184f
C29472 VPWR.n2754 0 9.72e-19
C29473 VPWR.n2755 0 0.0014f
C29474 VPWR.n2756 0 8.64e-19
C29475 VPWR.n2757 0 0.00108f
C29476 VPWR.n2758 0 0.00248f
C29477 VPWR.n2759 0 0.00389f
C29478 VPWR.n2760 0 0.00357f
C29479 VPWR.n2761 0 0.00281f
C29480 VPWR.n2762 0 0.0261f
C29481 VPWR.n2763 0 0.00162f
C29482 VPWR.n2764 0 0.00184f
C29483 VPWR.t190 0 0.0973f
C29484 VPWR.t95 0 0.107f
C29485 VPWR.n2765 0 0.185f
C29486 VPWR.n2766 0 0.0386f
C29487 VPWR.n2767 0 0.0819f
C29488 VPWR.n2768 0 0.13f
C29489 VPWR.t4 0 0.068f
C29490 VPWR.n2769 0 0.0701f
C29491 VPWR.n2770 0 0.0607f
C29492 VPWR.n2771 0 0.0571f
C29493 VPWR.t52 0 0.073f
C29494 VPWR.t186 0 0.0724f
C29495 VPWR.n2772 0 0.207f
C29496 VPWR.t16 0 0.073f
C29497 VPWR.n2773 0 0.207f
C29498 VPWR.n2774 0 0.00994f
C29499 VPWR.t157 0 0.0724f
C29500 VPWR.n2775 0 0.207f
C29501 VPWR.n2776 0 0.0787f
C29502 VPWR.t85 0 0.073f
C29503 VPWR.n2777 0 0.207f
C29504 VPWR.n2778 0 0.00265f
C29505 VPWR.n2779 0 0.00119f
C29506 VPWR.n2780 0 0.00302f
C29507 VPWR.n2781 0 0.00248f
C29508 VPWR.n2782 0 5.4e-19
C29509 VPWR.n2783 0 0.00259f
C29510 VPWR.n2784 0 0.00313f
C29511 VPWR.n2785 0 0.00151f
C29512 VPWR.n2786 0 0.00162f
C29513 VPWR.n2787 0 0.00119f
C29514 VPWR.n2788 0 0.00184f
C29515 VPWR.n2789 0 0.00259f
C29516 VPWR.n2790 0 0.00119f
C29517 VPWR.n2791 0 0.00421f
C29518 VPWR.n2792 0 0.00248f
C29519 VPWR.n2793 0 5.4e-19
C29520 VPWR.n2794 0 8.64e-19
C29521 VPWR.n2795 0 0.00227f
C29522 VPWR.n2796 0 0.00248f
C29523 VPWR.n2797 0 0.00248f
C29524 VPWR.n2798 0 0.00194f
C29525 VPWR.n2799 0 0.00184f
C29526 VPWR.n2800 0 0.00259f
C29527 VPWR.n2801 0 0.00119f
C29528 VPWR.n2802 0 0.00344f
C29529 VPWR.n2803 0 0.00248f
C29530 VPWR.n2804 0 0.00329f
C29531 VPWR.n2805 0 0.00208f
C29532 VPWR.n2806 0 0.00498f
C29533 VPWR.n2807 0 0.00891f
C29534 VPWR.n2808 0 0.00616f
C29535 VPWR.n2809 0 0.016f
C29536 VPWR.n2810 0 0.00561f
C29537 VPWR.n2811 0 0.0128f
C29538 VPWR.n2812 0 0.0529f
C29539 VPWR.n2813 0 0.0575f
C29540 VPWR.n2814 0 0.0457f
C29541 VPWR.n2815 0 0.0159f
C29542 VPWR.t102 0 0.0949f
C29543 VPWR.n2816 0 0.101f
C29544 VPWR.n2817 0 0.0331f
C29545 VPWR.n2818 0 0.0369f
C29546 VPWR.n2819 0 0.0425f
C29547 VPWR.n2820 0 0.0199f
C29548 VPWR.n2821 0 0.0513f
C29549 VPWR.n2822 0 0.0199f
C29550 VPWR.n2823 0 0.0214f
C29551 VPWR.n2824 0 0.0369f
C29552 VPWR.n2825 0 0.0513f
C29553 VPWR.n2826 0 0.0199f
C29554 VPWR.n2827 0 0.0475f
C29555 VPWR.n2828 0 0.0369f
C29556 VPWR.n2829 0 0.0534f
C29557 VPWR.n2830 0 0.0199f
C29558 VPWR.n2831 0 0.0547f
C29559 VPWR.n2832 0 0.0199f
C29560 VPWR.n2833 0 0.0522f
C29561 VPWR.n2834 0 0.0199f
C29562 VPWR.n2835 0 0.0819f
C29563 VPWR.n2836 0 0.0199f
C29564 VPWR.n2837 0 0.0118f
C29565 VPWR.n2838 0 0.116f
C29566 VPWR.n2839 0 0.0674f
C29567 VPWR.n2840 0 0.0143f
C29568 VPWR.n2841 0 0.0143f
C29569 VPWR.n2842 0 0.00994f
C29570 VPWR.n2843 0 0.00451f
C29571 VPWR.n2844 0 0.0783f
C29572 VPWR.n2845 0 0.0311f
C29573 VPWR.n2846 0 0.0429f
C29574 VPWR.n2847 0 0.023f
C29575 VPWR.n2848 0 0.00994f
C29576 VPWR.n2849 0 0.078f
C29577 VPWR.n2850 0 0.0512f
C29578 VPWR.n2851 0 0.0246f
C29579 VPWR.n2852 0 0.081f
C29580 VPWR.n2853 0 0.0165f
C29581 VPWR.n2854 0 0.0143f
C29582 VPWR.n2855 0 0.0429f
C29583 VPWR.n2856 0 0.207f
C29584 VPWR.n2857 0 0.0775f
C29585 VPWR.n2858 0 0.0143f
C29586 VPWR.n2859 0 0.0107f
C29587 VPWR.n2860 0 0.0608f
C29588 VPWR.n2861 0 0.0173f
C29589 VPWR.n2862 0 0.0199f
C29590 VPWR.n2863 0 0.0199f
C29591 VPWR.n2864 0 0.0118f
C29592 VPWR.n2865 0 0.0634f
C29593 VPWR.n2866 0 0.00839f
C29594 VPWR.n2867 0 0.018f
C29595 VPWR.n2868 0 0.071f
C29596 VPWR.n2869 0 0.0199f
C29597 VPWR.n2870 0 0.0404f
C29598 VPWR.n2871 0 0.0199f
C29599 VPWR.n2872 0 0.0123f
C29600 VPWR.n2873 0 0.0199f
C29601 VPWR.n2874 0 0.0533f
C29602 VPWR.n2875 0 0.0199f
C29603 VPWR.n2876 0 0.00559f
C29604 VPWR.n2877 0 0.0199f
C29605 VPWR.n2878 0 0.00704f
C29606 VPWR.n2879 0 0.0199f
C29607 VPWR.n2880 0 0.00677f
C29608 VPWR.n2881 0 0.0199f
C29609 VPWR.n2882 0 0.065f
C29610 VPWR.n2883 0 0.0199f
C29611 VPWR.n2884 0 0.00448f
C29612 VPWR.n2885 0 0.0199f
C29613 VPWR.n2886 0 0.0206f
C29614 VPWR.n2887 0 0.0199f
C29615 VPWR.n2888 0 0.0487f
C29616 VPWR.n2889 0 0.0199f
C29617 VPWR.n2890 0 0.0118f
C29618 VPWR.n2891 0 0.0077f
C29619 VPWR.n2892 0 0.00704f
C29620 VPWR.n2893 0 0.018f
C29621 VPWR.n2894 0 0.0126f
C29622 VPWR.n2895 0 0.00655f
C29623 VPWR.n2896 0 0.0794f
C29624 VPWR.n2897 0 0.0172f
C29625 VPWR.n2898 0 0.0452f
C29626 VPWR.n2899 0 0.0199f
C29627 VPWR.n2900 0 0.0199f
C29628 VPWR.n2901 0 0.0199f
C29629 VPWR.n2902 0 0.0118f
C29630 VPWR.n2903 0 0.0207f
C29631 VPWR.n2904 0 0.113f
C29632 VPWR.n2905 0 0.216f
C29633 VPWR.n2906 0 0.018f
C29634 VPWR.n2907 0 0.00335f
C29635 VPWR.n2908 0 0.00367f
C29636 VPWR.n2909 0 0.00281f
C29637 VPWR.n2910 0 0.00313f
C29638 VPWR.n2911 0 0.00989f
C29639 VPWR.n2912 0 0.00496f
C29640 VPWR.n2913 0 0.0217f
C29641 VPWR.n2914 0 0.00248f
C29642 VPWR.n2915 0 0.00344f
C29643 VPWR.n2916 0 0.00468f
C29644 VPWR.n2917 0 0.00323f
C29645 VPWR.n2918 0 0.00208f
C29646 VPWR.n2920 0 0.36f
C29647 VPWR.n2921 0 0.366f
C29648 VPWR.n2922 0 0.0362f
C29649 VPWR.n2923 0 0.00468f
C29650 VPWR.n2924 0 0.00323f
C29651 VPWR.n2925 0 0.00461f
C29652 VPWR.n2926 0 0.00208f
C29653 VPWR.n2928 0 0.0217f
C29654 VPWR.n2929 0 0.00203f
C29655 VPWR.n2930 0 0.00257f
C29656 VPWR.n2931 0 0.00208f
C29657 VPWR.n2932 0 0.00481f
C29658 VPWR.n2933 0 0.00744f
C29659 VPWR.n2934 0 0.00259f
C29660 VPWR.n2935 0 0.00259f
C29661 VPWR.n2936 0 0.0135f
C29662 VPWR.n2937 0 0.00292f
C29663 VPWR.n2938 0 0.00482f
C29664 VPWR.n2939 0 0.00184f
C29665 VPWR.n2940 0 0.00994f
C29666 VPWR.t298 0 0.068f
C29667 VPWR.n2941 0 0.0657f
C29668 VPWR.n2942 0 0.0706f
C29669 VPWR.n2943 0 0.0391f
C29670 VPWR.n2944 0 0.0196f
C29671 VPWR.n2945 0 0.0199f
C29672 VPWR.n2946 0 0.0629f
C29673 VPWR.n2947 0 0.0485f
C29674 VPWR.n2948 0 0.0118f
C29675 VPWR.n2949 0 0.0199f
C29676 VPWR.n2950 0 0.018f
C29677 VPWR.n2951 0 0.0916f
C29678 VPWR.n2952 0 0.0555f
C29679 VPWR.n2953 0 0.0971f
C29680 VPWR.n2954 0 0.0485f
C29681 VPWR.n2955 0 0.0118f
C29682 VPWR.n2956 0 0.0199f
C29683 VPWR.n2957 0 0.018f
C29684 VPWR.n2958 0 0.0916f
C29685 VPWR.n2959 0 0.0555f
C29686 VPWR.n2960 0 0.0971f
C29687 VPWR.t155 0 0.068f
C29688 VPWR.n2961 0 0.0769f
C29689 VPWR.n2962 0 0.0426f
C29690 VPWR.n2963 0 0.107f
C29691 VPWR.n2964 0 0.0485f
C29692 VPWR.n2965 0 0.018f
C29693 VPWR.n2966 0 0.0199f
C29694 VPWR.n2967 0 0.0199f
C29695 VPWR.n2968 0 0.0118f
C29696 VPWR.n2969 0 0.00994f
C29697 VPWR.n2970 0 0.0384f
C29698 VPWR.n2971 0 0.0368f
C29699 VPWR.n2972 0 0.018f
C29700 VPWR.n2973 0 0.00656f
C29701 VPWR.n2974 0 0.0199f
C29702 VPWR.n2975 0 0.0315f
C29703 VPWR.n2976 0 0.0199f
C29704 VPWR.n2977 0 0.01f
C29705 VPWR.n2978 0 0.0199f
C29706 VPWR.n2979 0 0.0544f
C29707 VPWR.n2980 0 0.0199f
C29708 VPWR.n2981 0 0.00521f
C29709 VPWR.n2982 0 0.0199f
C29710 VPWR.t152 0 0.068f
C29711 VPWR.n2983 0 0.0929f
C29712 VPWR.n2984 0 0.0612f
C29713 VPWR.n2985 0 0.0199f
C29714 VPWR.n2986 0 0.0391f
C29715 VPWR.n2987 0 0.0199f
C29716 VPWR.n2988 0 0.0671f
C29717 VPWR.n2989 0 0.0199f
C29718 VPWR.n2990 0 0.0118f
C29719 VPWR.n2991 0 0.0381f
C29720 VPWR.n2992 0 0.0534f
C29721 VPWR.n2993 0 0.0513f
C29722 VPWR.n2994 0 0.105f
C29723 VPWR.t151 0 0.0876f
C29724 VPWR.n2995 0 0.0784f
C29725 VPWR.n2996 0 0.018f
C29726 VPWR.t343 0 0.112f
C29727 VPWR.n2997 0 0.264f
C29728 VPWR.n2998 0 0.0207f
C29729 VPWR.n2999 0 0.0654f
C29730 VPWR.n3000 0 0.236f
C29731 VPWR.n3001 0 0.0681f
C29732 VPWR.n3002 0 0.0133f
C29733 VPWR.n3003 0 0.0126f
C29734 VPWR.n3004 0 0.115f
C29735 VPWR.n3005 0 0.0522f
C29736 VPWR.n3006 0 0.149f
C29737 VPWR.n3007 0 0.0118f
C29738 VPWR.n3008 0 0.0173f
C29739 VPWR.n3009 0 0.0107f
C29740 VPWR.n3010 0 0.0733f
C29741 VPWR.n3011 0 0.00291f
C29742 VPWR.n3012 0 0.0118f
C29743 VPWR.n3013 0 0.0199f
C29744 VPWR.n3014 0 0.018f
C29745 VPWR.n3015 0 0.052f
C29746 VPWR.t136 0 0.0774f
C29747 VPWR.t11 0 0.0774f
C29748 VPWR.n3016 0 0.502f
C29749 VPWR.n3017 0 0.0276f
C29750 VPWR.n3018 0 0.0118f
C29751 VPWR.n3019 0 0.0199f
C29752 VPWR.n3020 0 0.018f
C29753 VPWR.n3021 0 0.0521f
C29754 VPWR.n3022 0 0.0667f
C29755 VPWR.n3023 0 0.0118f
C29756 VPWR.n3024 0 0.0199f
C29757 VPWR.n3025 0 0.0199f
C29758 VPWR.n3026 0 0.0173f
C29759 VPWR.n3027 0 0.0107f
C29760 VPWR.n3028 0 0.0386f
C29761 VPWR.n3029 0 0.307f
C29762 VPWR.n3030 0 0.0725f
C29763 VPWR.n3031 0 0.0495f
C29764 VPWR.n3032 0 0.0012f
C29765 VPWR.n3033 0 0.00164f
C29766 VPWR.n3034 0 0.00162f
C29767 VPWR.n3035 0 0.0027f
C29768 VPWR.n3036 0 0.0013f
C29769 VPWR.n3037 0 0.0013f
C29770 VPWR.n3038 0 0.0086f
C29771 VPWR.n3039 0 0.00494f
C29772 VPWR.n3040 0 0.00208f
C29773 VPWR.n3041 0 0.00257f
C29774 VPWR.n3042 0 0.00203f
C29775 VPWR.n3043 0 0.378f
C29776 VPWR.n3044 0 0.37f
C29777 VPWR.n3045 0 0.014f
C29778 VPWR.n3046 0 0.00461f
C29779 VPWR.n3047 0 0.00323f
C29780 VPWR.n3048 0 0.00208f
C29781 VPWR.n3050 0 0.0217f
C29782 VPWR.n3051 0 0.00468f
C29783 VPWR.n3052 0 0.00323f
C29784 VPWR.n3053 0 0.00461f
C29785 VPWR.n3054 0 0.00208f
C29786 VPWR.n3056 0 0.0362f
C29787 VPWR.n3057 0 0.366f
C29788 VPWR.n3058 0 0.36f
C29789 VPWR.n3059 0 0.00248f
C29790 VPWR.n3060 0 0.00344f
C29791 VPWR.n3061 0 0.00208f
C29792 VPWR.n3062 0 0.00323f
C29793 VPWR.n3063 0 0.00468f
C29794 VPWR.n3064 0 0.00323f
C29795 VPWR.n3065 0 0.00208f
C29796 VPWR.n3067 0 0.0216f
C29797 VPWR.n3069 0 0.00329f
C29798 VPWR.n3070 0 0.00208f
C29799 VPWR.n3071 0 0.00496f
C29800 VPWR.n3072 0 0.00859f
C29801 VPWR.n3073 0 0.00443f
C29802 VPWR.n3074 0 0.00281f
C29803 VPWR.n3075 0 0.00367f
C29804 VPWR.n3076 0 0.00281f
C29805 VPWR.n3077 0 0.00238f
C29806 VPWR.n3078 0 8.64e-19
C29807 VPWR.n3079 0 0.00302f
C29808 VPWR.n3080 0 0.00443f
C29809 VPWR.n3081 0 0.00205f
C29810 VPWR.n3082 0 0.00162f
C29811 VPWR.n3083 0 0.0027f
C29812 VPWR.n3084 0 0.0013f
C29813 VPWR.n3085 0 0.0013f
C29814 VPWR.n3086 0 0.0027f
C29815 VPWR.n3087 0 0.00162f
C29816 VPWR.n3088 0 0.00164f
C29817 VPWR.n3089 0 0.00212f
C29818 VPWR.n3090 0 0.038f
C29819 VPWR.n3091 0 0.307f
C29820 VPWR.n3092 0 0.306f
C29821 VPWR.n3093 0 0.129f
C29822 VPWR.n3094 0 0.306f
C29823 VPWR.n3095 0 0.658f
C29824 VPWR.n3096 0 0.0394f
C29825 VPWR.n3097 0 0.00248f
C29826 VPWR.n3098 0 0.0014f
C29827 VPWR.n3099 0 0.00162f
C29828 VPWR.n3100 0 0.00216f
C29829 VPWR.n3101 0 0.00357f
C29830 VPWR.n3102 0 0.00248f
C29831 VPWR.n3103 0 0.0014f
C29832 VPWR.n3104 0 0.00335f
C29833 VPWR.n3105 0 0.00248f
C29834 VPWR.n3106 0 0.0014f
C29835 VPWR.n3107 0 8.64e-19
C29836 VPWR.n3108 0 0.00173f
C29837 VPWR.n3109 0 0.00497f
C29838 VPWR.n3110 0 0.00378f
C29839 VPWR.n3111 0 0.00162f
C29840 VPWR.n3112 0 0.00151f
C29841 VPWR.n3113 0 0.0013f
C29842 VPWR.n3114 0 0.0014f
C29843 VPWR.n3115 0 0.00851f
C29844 VPWR.n3116 0 0.00493f
C29845 VPWR.n3117 0 0.0217f
C29846 VPWR.n3118 0 0.00248f
C29847 VPWR.n3119 0 0.00344f
C29848 VPWR.n3120 0 0.00208f
C29849 VPWR.n3121 0 0.00323f
C29850 VPWR.n3122 0 0.00468f
C29851 VPWR.n3123 0 0.00323f
C29852 VPWR.n3124 0 0.00208f
C29853 VPWR.n3126 0 0.36f
C29854 VPWR.n3127 0 0.366f
C29855 VPWR.n3128 0 0.0362f
C29856 VPWR.n3130 0 0.127f
C29857 VPWR.n3131 0 0.00457f
C29858 VPWR.n3132 0 0.00468f
C29859 VPWR.n3133 0 0.00323f
C29860 VPWR.n3134 0 0.00208f
C29861 VPWR.n3136 0 0.014f
C29862 VPWR.n3137 0 0.37f
C29863 VPWR.n3138 0 0.378f
C29864 VPWR.n3139 0 0.381f
C29865 VPWR.n3140 0 0.381f
C29866 VPWR.n3141 0 0.00248f
C29867 VPWR.n3142 0 0.00344f
C29868 VPWR.n3143 0 0.00208f
C29869 VPWR.n3144 0 0.00323f
C29870 VPWR.n3145 0 0.00468f
C29871 VPWR.n3146 0 0.00323f
C29872 VPWR.n3147 0 0.00208f
C29873 VPWR.n3149 0 0.00329f
C29874 VPWR.n3150 0 0.00208f
C29875 VPWR.n3151 0 0.00259f
C29876 VPWR.n3152 0 0.0299f
C29877 VPWR.n3153 0 0.0199f
C29878 VPWR.t309 0 0.068f
C29879 VPWR.n3154 0 0.00571f
C29880 VPWR.n3155 0 0.018f
C29881 VPWR.n3156 0 0.0144f
C29882 VPWR.t3 0 0.0951f
C29883 VPWR.t284 0 0.0774f
C29884 VPWR.t304 0 0.0417f
C29885 VPWR.t279 0 0.0417f
C29886 VPWR.n3157 0 0.383f
C29887 VPWR.n3158 0 0.0385f
C29888 VPWR.n3159 0 0.0419f
C29889 VPWR.n3160 0 0.294f
C29890 VPWR.n3161 0 0.333f
C29891 VPWR.n3162 0 0.0701f
C29892 VPWR.n3163 0 0.0602f
C29893 VPWR.n3164 0 0.0416f
C29894 VPWR.n3165 0 0.0107f
C29895 VPWR.n3166 0 0.018f
C29896 VPWR.n3167 0 0.00918f
C29897 VPWR.n3168 0 0.049f
C29898 VPWR.n3169 0 0.0701f
C29899 VPWR.n3170 0 0.0391f
C29900 VPWR.t35 0 0.0711f
C29901 VPWR.n3171 0 0.195f
C29902 VPWR.n3172 0 0.0877f
C29903 VPWR.n3173 0 0.0534f
C29904 VPWR.n3174 0 0.0118f
C29905 VPWR.n3175 0 0.00994f
C29906 VPWR.n3176 0 0.01f
C29907 VPWR.n3177 0 0.0505f
C29908 VPWR.n3178 0 0.028f
C29909 VPWR.n3179 0 0.0179f
C29910 VPWR.n3180 0 0.0184f
C29911 VPWR.n3181 0 0.0199f
C29912 VPWR.n3182 0 0.0403f
C29913 VPWR.n3183 0 0.0199f
C29914 VPWR.n3184 0 0.031f
C29915 VPWR.n3185 0 0.0199f
C29916 VPWR.n3186 0 0.0125f
C29917 VPWR.n3187 0 0.00655f
C29918 VPWR.n3188 0 0.049f
C29919 VPWR.n3189 0 0.0173f
C29920 VPWR.t45 0 0.068f
C29921 VPWR.n3190 0 0.0701f
C29922 VPWR.n3191 0 0.0627f
C29923 VPWR.n3192 0 0.0199f
C29924 VPWR.n3193 0 0.0363f
C29925 VPWR.n3194 0 0.0602f
C29926 VPWR.n3195 0 0.0186f
C29927 VPWR.n3196 0 0.00994f
C29928 VPWR.n3197 0 0.00184f
C29929 VPWR.n3198 0 0.015f
C29930 VPWR.n3199 0 0.0357f
C29931 VPWR.n3200 0 7.56e-19
C29932 VPWR.n3201 0 0.00162f
C29933 VPWR.n3202 0 0.00216f
C29934 VPWR.n3203 0 0.00357f
C29935 VPWR.n3204 0 0.00248f
C29936 VPWR.n3205 0 0.0014f
C29937 VPWR.n3206 0 0.00335f
C29938 VPWR.n3207 0 0.00248f
C29939 VPWR.n3208 0 0.0014f
C29940 VPWR.n3209 0 8.64e-19
C29941 VPWR.n3210 0 0.00173f
C29942 VPWR.n3211 0 0.00497f
C29943 VPWR.n3212 0 0.00378f
C29944 VPWR.n3213 0 0.00162f
C29945 VPWR.n3214 0 0.00151f
C29946 VPWR.n3215 0 0.0013f
C29947 VPWR.n3216 0 0.0014f
C29948 VPWR.n3217 0 0.00851f
C29949 VPWR.n3218 0 0.00493f
C29950 VPWR.n3219 0 0.0217f
C29951 VPWR.n3221 0 0.00208f
C29952 VPWR.n3222 0 0.00498f
C29953 VPWR.n3223 0 0.0123f
C29954 VPWR.n3224 0 0.00313f
C29955 VPWR.n3225 0 0.00397f
C29956 VPWR.n3226 0 0.00151f
C29957 VPWR.n3227 0 0.011f
C29958 VPWR.n3228 0 0.00162f
C29959 VPWR.n3229 0 0.00119f
C29960 VPWR.n3230 0 0.00184f
C29961 VPWR.n3231 0 0.00259f
C29962 VPWR.n3232 0 0.00119f
C29963 VPWR.n3233 0 0.00585f
C29964 VPWR.n3234 0 0.0743f
C29965 VPWR.t283 0 0.0774f
C29966 VPWR.n3235 0 0.0276f
C29967 VPWR.t28 0 0.0774f
C29968 VPWR.n3236 0 0.00555f
C29969 VPWR.n3237 0 0.124f
C29970 VPWR.n3238 0 0.0509f
C29971 VPWR.n3239 0 0.00555f
C29972 VPWR.n3240 0 0.0276f
C29973 VPWR.n3241 0 0.0118f
C29974 VPWR.n3242 0 0.0199f
C29975 VPWR.n3243 0 0.018f
C29976 VPWR.n3244 0 0.052f
C29977 VPWR.n3245 0 0.118f
C29978 VPWR.n3246 0 0.0118f
C29979 VPWR.n3247 0 0.1f
C29980 VPWR.n3248 0 0.0199f
C29981 VPWR.n3249 0 0.0973f
C29982 VPWR.n3250 0 0.0199f
C29983 VPWR.n3251 0 0.0973f
C29984 VPWR.n3252 0 0.0199f
C29985 VPWR.t308 0 0.0876f
C29986 VPWR.t44 0 0.0876f
C29987 VPWR.n3253 0 0.29f
C29988 VPWR.n3254 0 0.0199f
C29989 VPWR.n3255 0 0.118f
C29990 VPWR.n3256 0 0.0199f
C29991 VPWR.n3257 0 0.0199f
C29992 VPWR.n3258 0 0.0179f
C29993 VPWR.n3259 0 0.01f
C29994 VPWR.n3260 0 0.00593f
C29995 VPWR.n3261 0 0.503f
C29996 VPWR.n3262 0 0.00459f
C29997 VPWR.n3263 0 0.0118f
C29998 VPWR.n3264 0 0.0199f
C29999 VPWR.n3265 0 0.018f
C30000 VPWR.n3266 0 0.00994f
C30001 VPWR.n3267 0 0.00704f
C30002 VPWR.n3268 0 0.0831f
C30003 VPWR.n3269 0 0.0118f
C30004 VPWR.n3270 0 0.0535f
C30005 VPWR.n3271 0 0.0199f
C30006 VPWR.t100 0 0.068f
C30007 VPWR.n3272 0 0.0266f
C30008 VPWR.n3273 0 0.0649f
C30009 VPWR.n3274 0 0.0391f
C30010 VPWR.n3275 0 0.0159f
C30011 VPWR.n3276 0 0.00616f
C30012 VPWR.n3277 0 0.00891f
C30013 VPWR.n3278 0 0.00119f
C30014 VPWR.n3279 0 0.00259f
C30015 VPWR.n3280 0 0.00184f
C30016 VPWR.n3281 0 0.00194f
C30017 VPWR.n3282 0 0.00248f
C30018 VPWR.n3283 0 0.00248f
C30019 VPWR.n3284 0 0.00227f
C30020 VPWR.n3285 0 8.64e-19
C30021 VPWR.n3286 0 0.00259f
C30022 VPWR.n3287 0 5.4e-19
C30023 VPWR.n3288 0 0.00248f
C30024 VPWR.n3289 0 0.00302f
C30025 VPWR.n3290 0 0.00266f
C30026 VPWR.n3291 0 0.00119f
C30027 VPWR.n3292 0 0.00184f
C30028 VPWR.n3293 0 0.00248f
C30029 VPWR.n3294 0 0.0408f
C30030 VPWR.n3295 0 0.306f
C30031 VPWR.n3296 0 0.129f
C30032 VPWR.n3297 0 0.0704f
C30033 VPWR.n3298 0 0.0107f
C30034 VPWR.n3299 0 0.00994f
C30035 VPWR.n3300 0 0.00814f
C30036 VPWR.n3301 0 0.0875f
C30037 VPWR.n3302 0 0.207f
C30038 VPWR.t114 0 0.073f
C30039 VPWR.n3303 0 0.132f
C30040 VPWR.n3304 0 0.0429f
C30041 VPWR.n3305 0 0.0143f
C30042 VPWR.n3306 0 0.018f
C30043 VPWR.n3307 0 0.0118f
C30044 VPWR.n3308 0 0.0634f
C30045 VPWR.n3309 0 0.00617f
C30046 VPWR.n3310 0 0.018f
C30047 VPWR.n3311 0 0.0626f
C30048 VPWR.n3312 0 0.0199f
C30049 VPWR.n3313 0 0.0049f
C30050 VPWR.n3314 0 0.0199f
C30051 VPWR.n3315 0 0.0688f
C30052 VPWR.n3316 0 0.0199f
C30053 VPWR.n3317 0 0.0657f
C30054 VPWR.n3318 0 0.0199f
C30055 VPWR.n3319 0 0.0117f
C30056 VPWR.n3320 0 0.00463f
C30057 VPWR.n3321 0 0.104f
C30058 VPWR.n3322 0 0.207f
C30059 VPWR.t199 0 0.073f
C30060 VPWR.n3323 0 0.0455f
C30061 VPWR.n3324 0 0.132f
C30062 VPWR.n3325 0 0.0429f
C30063 VPWR.n3326 0 0.0145f
C30064 VPWR.n3327 0 0.018f
C30065 VPWR.n3328 0 0.0118f
C30066 VPWR.n3329 0 0.0128f
C30067 VPWR.n3330 0 0.062f
C30068 VPWR.n3331 0 0.018f
C30069 VPWR.n3332 0 0.00429f
C30070 VPWR.n3333 0 0.0199f
C30071 VPWR.n3334 0 0.0457f
C30072 VPWR.n3335 0 0.0199f
C30073 VPWR.n3336 0 0.0199f
C30074 VPWR.n3337 0 0.0199f
C30075 VPWR.n3338 0 0.0117f
C30076 VPWR.n3339 0 0.045f
C30077 VPWR.n3340 0 0.142f
C30078 VPWR.n3341 0 0.00284f
C30079 VPWR.n3342 0 0.00499f
C30080 VPWR.n3343 0 0.00281f
C30081 VPWR.n3344 0 0.00313f
C30082 VPWR.n3345 0 0.00989f
C30083 VPWR.n3346 0 0.00496f
C30084 VPWR.n3347 0 0.0217f
C30085 VPWR.n3349 0 0.00208f
C30086 VPWR.n3350 0 0.00483f
C30087 VPWR.n3351 0 0.00743f
C30088 VPWR.n3352 0 0.00259f
C30089 VPWR.n3353 0 0.00259f
C30090 VPWR.n3354 0 0.00292f
C30091 VPWR.n3355 0 0.00184f
C30092 VPWR.n3356 0 0.00184f
C30093 VPWR.n3357 0 0.0136f
C30094 VPWR.n3358 0 0.185f
C30095 VPWR.n3359 0 0.0683f
C30096 VPWR.n3360 0 0.0608f
C30097 VPWR.n3361 0 0.0386f
C30098 VPWR.n3362 0 0.018f
C30099 VPWR.n3363 0 0.0199f
C30100 VPWR.n3364 0 0.0199f
C30101 VPWR.n3365 0 0.0522f
C30102 VPWR.n3366 0 0.0199f
C30103 VPWR.n3367 0 0.0118f
C30104 VPWR.n3368 0 0.0535f
C30105 VPWR.n3369 0 0.0619f
C30106 VPWR.n3370 0 0.00994f
C30107 VPWR.n3371 0 0.00918f
C30108 VPWR.n3372 0 0.0312f
C30109 VPWR.n3373 0 0.0429f
C30110 VPWR.n3374 0 0.033f
C30111 VPWR.n3375 0 0.0125f
C30112 VPWR.n3376 0 0.115f
C30113 VPWR.t259 0 0.073f
C30114 VPWR.n3377 0 0.207f
C30115 VPWR.n3378 0 0.0674f
C30116 VPWR.n3379 0 0.0135f
C30117 VPWR.n3380 0 0.0143f
C30118 VPWR.n3381 0 0.028f
C30119 VPWR.n3382 0 0.0608f
C30120 VPWR.n3383 0 0.018f
C30121 VPWR.n3384 0 0.00429f
C30122 VPWR.n3385 0 0.0199f
C30123 VPWR.n3386 0 0.0447f
C30124 VPWR.n3387 0 0.0118f
C30125 VPWR.n3388 0 0.0276f
C30126 VPWR.n3389 0 0.00994f
C30127 VPWR.n3390 0 0.00994f
C30128 VPWR.t275 0 0.111f
C30129 VPWR.n3391 0 0.288f
C30130 VPWR.n3392 0 0.11f
C30131 VPWR.n3393 0 0.0756f
C30132 VPWR.n3394 0 0.0854f
C30133 VPWR.n3395 0 0.0485f
C30134 VPWR.n3396 0 0.0955f
C30135 VPWR.t198 0 0.068f
C30136 VPWR.t58 0 0.0711f
C30137 VPWR.n3397 0 0.195f
C30138 VPWR.n3398 0 0.0723f
C30139 VPWR.n3399 0 0.0181f
C30140 VPWR.n3400 0 0.0199f
C30141 VPWR.n3401 0 0.0457f
C30142 VPWR.n3402 0 0.00918f
C30143 VPWR.t207 0 0.0724f
C30144 VPWR.n3403 0 0.207f
C30145 VPWR.t59 0 0.073f
C30146 VPWR.n3404 0 0.0975f
C30147 VPWR.n3405 0 0.0429f
C30148 VPWR.n3406 0 0.0135f
C30149 VPWR.n3407 0 0.0107f
C30150 VPWR.n3408 0 0.0338f
C30151 VPWR.n3409 0 0.122f
C30152 VPWR.n3410 0 0.0176f
C30153 VPWR.n3411 0 0.0265f
C30154 VPWR.n3412 0 0.00923f
C30155 VPWR.n3413 0 0.0199f
C30156 VPWR.n3414 0 0.0604f
C30157 VPWR.n3415 0 0.018f
C30158 VPWR.n3416 0 0.00994f
C30159 VPWR.n3417 0 0.0118f
C30160 VPWR.n3418 0 0.0534f
C30161 VPWR.n3419 0 0.0877f
C30162 VPWR.n3420 0 0.0391f
C30163 VPWR.n3421 0 0.0701f
C30164 VPWR.n3422 0 0.048f
C30165 VPWR.n3423 0 0.00983f
C30166 VPWR.n3424 0 0.0118f
C30167 VPWR.n3425 0 0.0199f
C30168 VPWR.n3426 0 0.018f
C30169 VPWR.n3427 0 0.0522f
C30170 VPWR.n3428 0 0.0626f
C30171 VPWR.n3429 0 0.0118f
C30172 VPWR.n3430 0 0.0199f
C30173 VPWR.n3431 0 0.0199f
C30174 VPWR.n3432 0 0.0606f
C30175 VPWR.n3433 0 0.018f
C30176 VPWR.n3434 0 0.0363f
C30177 VPWR.n3435 0 0.0432f
C30178 VPWR.n3436 0 0.0107f
C30179 VPWR.n3437 0 0.0366f
C30180 VPWR.n3438 0 0.424f
C30181 VPWR.n3439 0 0.131f
C30182 VPWR.n3440 0 0.0552f
C30183 VPWR.n3441 0 0.00212f
C30184 VPWR.n3442 0 0.00164f
C30185 VPWR.n3443 0 0.00162f
C30186 VPWR.n3444 0 0.0027f
C30187 VPWR.n3445 0 0.0013f
C30188 VPWR.n3446 0 0.0013f
C30189 VPWR.n3447 0 0.00861f
C30190 VPWR.n3448 0 0.00495f
C30191 VPWR.n3449 0 0.0217f
C30192 VPWR.n3450 0 0.00248f
C30193 VPWR.n3451 0 0.00344f
C30194 VPWR.n3452 0 0.00468f
C30195 VPWR.n3453 0 0.00323f
C30196 VPWR.n3454 0 0.00208f
C30197 VPWR.n3456 0 0.381f
C30198 VPWR.n3457 0 0.381f
C30199 VPWR.n3458 0 0.00323f
C30200 VPWR.n3459 0 0.00248f
C30201 VPWR.n3460 0 0.00344f
C30202 VPWR.n3461 0 0.00208f
C30203 VPWR.n3463 0 0.00329f
C30204 VPWR.n3464 0 0.00208f
C30205 VPWR.n3465 0 0.00495f
C30206 VPWR.n3466 0 0.0217f
C30207 VPWR.n3467 0 0.00496f
C30208 VPWR.n3468 0 0.00486f
C30209 VPWR.n3469 0 0.00389f
C30210 VPWR.n3470 0 0.00173f
C30211 VPWR.n3471 0 0.0027f
C30212 VPWR.t133 0 0.0876f
C30213 VPWR.n3472 0 0.0487f
C30214 VPWR.n3473 0 0.125f
C30215 VPWR.n3474 0 0.00119f
C30216 VPWR.n3475 0 0.0341f
C30217 VPWR.t122 0 0.068f
C30218 VPWR.n3476 0 0.0939f
C30219 VPWR.n3477 0 0.0199f
C30220 VPWR.n3478 0 0.00655f
C30221 VPWR.n3479 0 0.0199f
C30222 VPWR.n3480 0 0.076f
C30223 VPWR.t342 0 0.068f
C30224 VPWR.n3481 0 0.0721f
C30225 VPWR.n3482 0 0.0619f
C30226 VPWR.t339 0 0.0417f
C30227 VPWR.t318 0 0.0417f
C30228 VPWR.n3483 0 0.384f
C30229 VPWR.n3484 0 0.0197f
C30230 VPWR.n3485 0 0.0118f
C30231 VPWR.n3486 0 0.018f
C30232 VPWR.n3487 0 0.0535f
C30233 VPWR.n3488 0 0.0391f
C30234 VPWR.n3489 0 0.0118f
C30235 VPWR.n3490 0 0.0199f
C30236 VPWR.n3491 0 0.0199f
C30237 VPWR.n3492 0 0.0457f
C30238 VPWR.n3493 0 0.00972f
C30239 VPWR.n3494 0 0.0755f
C30240 VPWR.n3495 0 0.018f
C30241 VPWR.n3496 0 0.0118f
C30242 VPWR.n3497 0 0.0634f
C30243 VPWR.n3498 0 0.0535f
C30244 VPWR.n3499 0 0.0391f
C30245 VPWR.n3500 0 0.0199f
C30246 VPWR.n3501 0 0.0181f
C30247 VPWR.n3502 0 0.0499f
C30248 VPWR.n3503 0 0.0157f
C30249 VPWR.n3504 0 0.0117f
C30250 VPWR.n3505 0 0.0394f
C30251 VPWR.n3506 0 0.0199f
C30252 VPWR.n3507 0 0.00704f
C30253 VPWR.n3508 0 0.0199f
C30254 VPWR.n3509 0 0.00704f
C30255 VPWR.n3510 0 0.0199f
C30256 VPWR.n3511 0 0.00559f
C30257 VPWR.n3512 0 0.0199f
C30258 VPWR.n3513 0 0.0199f
C30259 VPWR.n3514 0 0.0331f
C30260 VPWR.n3515 0 0.0199f
C30261 VPWR.n3516 0 0.018f
C30262 VPWR.n3517 0 0.0238f
C30263 VPWR.n3518 0 0.101f
C30264 VPWR.n3519 0 0.0118f
C30265 VPWR.n3520 0 0.0672f
C30266 VPWR.n3521 0 0.0199f
C30267 VPWR.n3522 0 0.0756f
C30268 VPWR.n3523 0 0.0199f
C30269 VPWR.n3524 0 0.0651f
C30270 VPWR.n3525 0 0.018f
C30271 VPWR.n3526 0 0.00983f
C30272 VPWR.n3527 0 0.00184f
C30273 VPWR.n3528 0 0.00881f
C30274 VPWR.n3529 0 0.00119f
C30275 VPWR.n3530 0 0.0027f
C30276 VPWR.n3531 0 0.00173f
C30277 VPWR.n3532 0 0.00194f
C30278 VPWR.n3533 0 0.00378f
C30279 VPWR.n3534 0 0.00248f
C30280 VPWR.n3535 0 0.00108f
C30281 VPWR.n3536 0 8.64e-19
C30282 VPWR.n3537 0 0.0014f
C30283 VPWR.n3538 0 4.32e-19
C30284 VPWR.n3539 0 0.00184f
C30285 VPWR.n3540 0 0.00108f
C30286 VPWR.n3541 0 0.0013f
C30287 VPWR.n3542 0 0.00194f
C30288 VPWR.n3543 0 0.00367f
C30289 VPWR.n3544 0 0.00281f
C30290 VPWR.n3545 0 0.00238f
C30291 VPWR.n3546 0 8.64e-19
C30292 VPWR.n3547 0 0.00302f
C30293 VPWR.n3548 0 0.00443f
C30294 VPWR.n3549 0 0.00205f
C30295 VPWR.n3550 0 0.00162f
C30296 VPWR.n3551 0 0.0027f
C30297 VPWR.n3552 0 0.0013f
C30298 VPWR.n3553 0 0.0013f
C30299 VPWR.n3554 0 0.00497f
C30300 VPWR.n3555 0 0.0143f
C30301 VPWR.n3556 0 0.0145f
C30302 VPWR.n3557 0 0.151f
C30303 VPWR.n3558 0 0.0117f
C30304 VPWR.n3559 0 0.051f
C30305 VPWR.n3560 0 0.0199f
C30306 VPWR.n3561 0 0.00555f
C30307 VPWR.n3562 0 0.0199f
C30308 VPWR.n3563 0 0.018f
C30309 VPWR.n3564 0 0.0542f
C30310 VPWR.n3565 0 0.062f
C30311 VPWR.n3566 0 0.0118f
C30312 VPWR.n3567 0 0.0199f
C30313 VPWR.n3568 0 0.0199f
C30314 VPWR.n3569 0 0.0181f
C30315 VPWR.n3570 0 0.00983f
C30316 VPWR.n3571 0 0.00606f
C30317 VPWR.n3572 0 0.0634f
C30318 VPWR.n3573 0 0.0118f
C30319 VPWR.n3574 0 0.0199f
C30320 VPWR.n3575 0 0.0199f
C30321 VPWR.n3576 0 0.0895f
C30322 VPWR.n3577 0 0.0394f
C30323 VPWR.n3578 0 0.0372f
C30324 VPWR.n3579 0 0.0118f
C30325 VPWR.n3580 0 0.0619f
C30326 VPWR.n3581 0 0.0535f
C30327 VPWR.n3582 0 0.0532f
C30328 VPWR.n3583 0 0.0117f
C30329 VPWR.n3584 0 0.0199f
C30330 VPWR.n3585 0 0.0199f
C30331 VPWR.n3586 0 0.0173f
C30332 VPWR.n3587 0 0.0107f
C30333 VPWR.n3588 0 0.0386f
C30334 VPWR.n3589 0 0.0619f
C30335 VPWR.n3590 0 0.0118f
C30336 VPWR.n3591 0 0.0199f
C30337 VPWR.n3592 0 0.0199f
C30338 VPWR.n3593 0 0.018f
C30339 VPWR.n3594 0 0.0485f
C30340 VPWR.n3595 0 0.0629f
C30341 VPWR.n3596 0 0.0118f
C30342 VPWR.n3597 0 0.0199f
C30343 VPWR.n3598 0 0.0199f
C30344 VPWR.n3599 0 0.0429f
C30345 VPWR.n3600 0 0.0394f
C30346 VPWR.t82 0 0.116f
C30347 VPWR.n3601 0 0.322f
C30348 VPWR.n3602 0 0.167f
C30349 VPWR.n3603 0 0.0373f
C30350 VPWR.n3604 0 0.0107f
C30351 VPWR.n3605 0 0.0556f
C30352 VPWR.n3606 0 0.0619f
C30353 VPWR.n3607 0 0.0117f
C30354 VPWR.n3608 0 0.107f
C30355 VPWR.n3609 0 0.0199f
C30356 VPWR.n3610 0 0.0428f
C30357 VPWR.n3611 0 0.0199f
C30358 VPWR.t183 0 0.068f
C30359 VPWR.n3612 0 0.0701f
C30360 VPWR.n3613 0 0.0919f
C30361 VPWR.n3614 0 0.0199f
C30362 VPWR.n3615 0 0.00735f
C30363 VPWR.n3616 0 0.0199f
C30364 VPWR.n3617 0 0.00704f
C30365 VPWR.n3618 0 0.0199f
C30366 VPWR.n3619 0 0.106f
C30367 VPWR.n3620 0 0.00735f
C30368 VPWR.n3621 0 0.018f
C30369 VPWR.n3622 0 0.0118f
C30370 VPWR.n3623 0 0.0199f
C30371 VPWR.n3624 0 0.0179f
C30372 VPWR.n3625 0 0.105f
C30373 VPWR.n3626 0 0.0606f
C30374 VPWR.n3627 0 0.01f
C30375 VPWR.n3628 0 0.0108f
C30376 VPWR.n3629 0 0.0183f
C30377 VPWR.n3630 0 0.00259f
C30378 VPWR.n3631 0 0.00259f
C30379 VPWR.n3632 0 0.0014f
C30380 VPWR.n3633 0 0.00162f
C30381 VPWR.n3634 0 0.00335f
C30382 VPWR.n3635 0 0.00421f
C30383 VPWR.n3636 0 0.00248f
C30384 VPWR.n3637 0 7.56e-19
C30385 VPWR.n3638 0 8.64e-19
C30386 VPWR.n3639 0 0.00108f
C30387 VPWR.n3640 0 0.00205f
C30388 VPWR.n3641 0 0.00248f
C30389 VPWR.n3642 0 0.0027f
C30390 VPWR.n3643 0 0.00302f
C30391 VPWR.n3644 0 0.00184f
C30392 VPWR.n3645 0 9.72e-19
C30393 VPWR.n3646 0 0.0014f
C30394 VPWR.n3647 0 8.64e-19
C30395 VPWR.n3648 0 0.00108f
C30396 VPWR.n3649 0 0.00248f
C30397 VPWR.n3650 0 0.00389f
C30398 VPWR.n3651 0 0.00357f
C30399 VPWR.n3652 0 0.00281f
C30400 VPWR.n3653 0 0.00989f
C30401 VPWR.n3654 0 0.00313f
C30402 VPWR.n3655 0 0.00918f
C30403 VPWR.n3656 0 0.0328f
C30404 VPWR.n3657 0 0.0958f
C30405 VPWR.n3658 0 0.0125f
C30406 VPWR.n3659 0 0.0199f
C30407 VPWR.n3660 0 0.0199f
C30408 VPWR.t110 0 0.0876f
C30409 VPWR.n3661 0 0.149f
C30410 VPWR.n3662 0 0.0199f
C30411 VPWR.n3663 0 0.0173f
C30412 VPWR.n3664 0 0.0107f
C30413 VPWR.n3665 0 0.00939f
C30414 VPWR.n3666 0 0.012f
C30415 VPWR.n3667 0 0.0118f
C30416 VPWR.n3668 0 0.018f
C30417 VPWR.n3669 0 0.00994f
C30418 VPWR.n3670 0 0.00655f
C30419 VPWR.n3671 0 0.0675f
C30420 VPWR.n3672 0 0.0118f
C30421 VPWR.n3673 0 0.0199f
C30422 VPWR.n3674 0 0.0199f
C30423 VPWR.n3675 0 0.0181f
C30424 VPWR.n3676 0 0.049f
C30425 VPWR.n3677 0 0.00755f
C30426 VPWR.n3678 0 0.0117f
C30427 VPWR.n3679 0 0.0612f
C30428 VPWR.n3680 0 0.0199f
C30429 VPWR.n3681 0 0.0233f
C30430 VPWR.n3682 0 0.0199f
C30431 VPWR.n3683 0 0.00448f
C30432 VPWR.n3684 0 0.0199f
C30433 VPWR.n3685 0 0.0199f
C30434 VPWR.n3686 0 0.00677f
C30435 VPWR.n3687 0 0.0199f
C30436 VPWR.n3688 0 0.0191f
C30437 VPWR.n3689 0 0.0199f
C30438 VPWR.n3690 0 0.0176f
C30439 VPWR.n3691 0 0.0199f
C30440 VPWR.n3692 0 0.018f
C30441 VPWR.n3693 0 0.0337f
C30442 VPWR.n3694 0 0.071f
C30443 VPWR.n3695 0 0.0118f
C30444 VPWR.n3696 0 0.0199f
C30445 VPWR.n3697 0 0.0199f
C30446 VPWR.n3698 0 0.0475f
C30447 VPWR.n3699 0 0.0173f
C30448 VPWR.n3700 0 0.00994f
C30449 VPWR.n3701 0 0.061f
C30450 VPWR.n3702 0 0.0534f
C30451 VPWR.t214 0 0.0711f
C30452 VPWR.n3703 0 0.195f
C30453 VPWR.n3704 0 0.0877f
C30454 VPWR.n3705 0 0.0391f
C30455 VPWR.n3706 0 0.0181f
C30456 VPWR.n3707 0 0.00994f
C30457 VPWR.n3708 0 0.049f
C30458 VPWR.n3709 0 0.00755f
C30459 VPWR.n3710 0 0.0117f
C30460 VPWR.n3711 0 0.0644f
C30461 VPWR.n3712 0 0.0199f
C30462 VPWR.n3713 0 0.011f
C30463 VPWR.n3714 0 0.0199f
C30464 VPWR.n3715 0 0.018f
C30465 VPWR.n3716 0 0.034f
C30466 VPWR.n3717 0 0.0634f
C30467 VPWR.n3718 0 0.0118f
C30468 VPWR.n3719 0 0.0199f
C30469 VPWR.n3720 0 0.0199f
C30470 VPWR.n3721 0 0.0181f
C30471 VPWR.n3722 0 0.00983f
C30472 VPWR.n3723 0 0.00544f
C30473 VPWR.n3724 0 0.0924f
C30474 VPWR.n3725 0 0.0144f
C30475 VPWR.n3726 0 0.0265f
C30476 VPWR.n3727 0 0.0107f
C30477 VPWR.n3728 0 0.00593f
C30478 VPWR.n3729 0 0.0057f
C30479 VPWR.n3730 0 0.0118f
C30480 VPWR.n3731 0 0.0199f
C30481 VPWR.n3732 0 0.018f
C30482 VPWR.n3733 0 0.00994f
C30483 VPWR.n3734 0 0.00704f
C30484 VPWR.n3735 0 0.0831f
C30485 VPWR.n3736 0 0.0118f
C30486 VPWR.n3737 0 0.0535f
C30487 VPWR.n3738 0 0.0199f
C30488 VPWR.t239 0 0.068f
C30489 VPWR.n3739 0 0.0266f
C30490 VPWR.n3740 0 0.0649f
C30491 VPWR.n3741 0 0.0391f
C30492 VPWR.n3742 0 0.0159f
C30493 VPWR.n3743 0 0.00616f
C30494 VPWR.n3744 0 0.00891f
C30495 VPWR.n3745 0 0.00119f
C30496 VPWR.n3746 0 0.00259f
C30497 VPWR.n3747 0 0.00184f
C30498 VPWR.n3748 0 0.00194f
C30499 VPWR.n3749 0 0.00248f
C30500 VPWR.n3750 0 0.00248f
C30501 VPWR.n3751 0 0.00227f
C30502 VPWR.n3752 0 8.64e-19
C30503 VPWR.n3753 0 0.00259f
C30504 VPWR.n3754 0 5.4e-19
C30505 VPWR.n3755 0 0.00248f
C30506 VPWR.n3756 0 0.00302f
C30507 VPWR.n3757 0 0.00266f
C30508 VPWR.n3758 0 0.00119f
C30509 VPWR.n3759 0 0.00184f
C30510 VPWR.n3760 0 0.00248f
C30511 VPWR.n3761 0 0.0014f
C30512 VPWR.n3762 0 0.00162f
C30513 VPWR.n3763 0 0.00216f
C30514 VPWR.n3764 0 0.00357f
C30515 VPWR.n3765 0 0.00248f
C30516 VPWR.n3766 0 0.0014f
C30517 VPWR.n3767 0 0.00335f
C30518 VPWR.n3768 0 0.00248f
C30519 VPWR.n3769 0 0.0014f
C30520 VPWR.n3770 0 8.64e-19
C30521 VPWR.n3771 0 0.00173f
C30522 VPWR.n3772 0 0.00497f
C30523 VPWR.n3773 0 0.00378f
C30524 VPWR.n3774 0 0.00162f
C30525 VPWR.n3775 0 0.00151f
C30526 VPWR.n3776 0 0.0013f
C30527 VPWR.n3777 0 0.0014f
C30528 VPWR.n3778 0 0.00851f
C30529 VPWR.n3779 0 0.00493f
C30530 VPWR.n3780 0 0.0217f
C30531 VPWR.n3781 0 0.00248f
C30532 VPWR.n3782 0 0.00344f
C30533 VPWR.n3783 0 0.00208f
C30534 VPWR.n3784 0 0.00323f
C30535 VPWR.n3785 0 0.00468f
C30536 VPWR.n3786 0 0.00323f
C30537 VPWR.n3787 0 0.00208f
C30538 VPWR.n3789 0 0.381f
C30539 VPWR.n3790 0 0.381f
C30540 VPWR.n3791 0 0.0412f
C30541 VPWR.n3792 0 0.403f
C30542 VPWR.n3793 0 0.347f
C30543 VPWR.n3794 0 0.00248f
C30544 VPWR.n3795 0 0.00344f
C30545 VPWR.n3796 0 0.00208f
C30546 VPWR.n3797 0 0.00323f
C30547 VPWR.n3798 0 0.00468f
C30548 VPWR.n3799 0 0.00323f
C30549 VPWR.n3800 0 0.00208f
C30550 VPWR.n3802 0 0.00329f
C30551 VPWR.n3803 0 0.00208f
C30552 VPWR.n3804 0 0.00259f
C30553 VPWR.t344 0 0.0774f
C30554 VPWR.n3805 0 0.338f
C30555 VPWR.n3806 0 0.209f
C30556 VPWR.t360 0 0.112f
C30557 VPWR.n3807 0 0.253f
C30558 VPWR.t294 0 0.116f
C30559 VPWR.n3808 0 0.325f
C30560 VPWR.n3809 0 0.0848f
C30561 VPWR.n3810 0 0.0522f
C30562 VPWR.n3811 0 0.00994f
C30563 VPWR.t382 0 0.078f
C30564 VPWR.n3812 0 0.0107f
C30565 VPWR.t331 0 0.0774f
C30566 VPWR.t263 0 0.0417f
C30567 VPWR.t379 0 0.0417f
C30568 VPWR.n3813 0 0.383f
C30569 VPWR.n3814 0 0.0384f
C30570 VPWR.n3815 0 0.0421f
C30571 VPWR.t321 0 0.0774f
C30572 VPWR.n3816 0 0.501f
C30573 VPWR.n3817 0 0.102f
C30574 VPWR.n3818 0 0.018f
C30575 VPWR.n3819 0 0.00429f
C30576 VPWR.n3820 0 0.0199f
C30577 VPWR.n3821 0 0.0117f
C30578 VPWR.n3822 0 0.0609f
C30579 VPWR.n3823 0 0.0135f
C30580 VPWR.n3824 0 0.356f
C30581 VPWR.n3825 0 0.018f
C30582 VPWR.n3826 0 0.0199f
C30583 VPWR.n3827 0 0.0199f
C30584 VPWR.n3828 0 0.0126f
C30585 VPWR.n3829 0 0.0958f
C30586 VPWR.n3830 0 0.0328f
C30587 VPWR.n3831 0 0.00907f
C30588 VPWR.n3832 0 0.126f
C30589 VPWR.n3833 0 0.0244f
C30590 VPWR.n3834 0 0.0232f
C30591 VPWR.n3835 0 0.00119f
C30592 VPWR.n3836 0 0.00162f
C30593 VPWR.n3837 0 0.00215f
C30594 VPWR.n3838 0 0.053f
C30595 VPWR.n3839 0 0.00113f
C30596 VPWR.n3840 0 0.00417f
C30597 VPWR.n3841 0 0.00421f
C30598 VPWR.n3842 0 0.00248f
C30599 VPWR.n3843 0 5.4e-19
C30600 VPWR.n3844 0 0.00259f
C30601 VPWR.n3845 0 0.00184f
C30602 VPWR.n3846 0 0.00194f
C30603 VPWR.n3847 0 0.00248f
C30604 VPWR.n3848 0 0.00248f
C30605 VPWR.n3849 0 0.00227f
C30606 VPWR.n3850 0 8.64e-19
C30607 VPWR.n3851 0 0.00259f
C30608 VPWR.n3852 0 5.4e-19
C30609 VPWR.n3853 0 0.00248f
C30610 VPWR.n3854 0 0.00302f
C30611 VPWR.n3855 0 0.00119f
C30612 VPWR.n3856 0 0.00184f
C30613 VPWR.n3857 0 0.13f
C30614 VPWR.n3858 0 0.0364f
C30615 VPWR.n3859 0 0.00248f
C30616 VPWR.n3860 0 0.0014f
C30617 VPWR.n3861 0 0.00162f
C30618 VPWR.n3862 0 0.00216f
C30619 VPWR.n3863 0 0.00357f
C30620 VPWR.n3864 0 0.00248f
C30621 VPWR.n3865 0 0.0014f
C30622 VPWR.n3866 0 0.00335f
C30623 VPWR.n3867 0 0.00248f
C30624 VPWR.n3868 0 0.0014f
C30625 VPWR.n3869 0 8.64e-19
C30626 VPWR.n3870 0 0.00173f
C30627 VPWR.n3871 0 0.00497f
C30628 VPWR.n3872 0 0.00378f
C30629 VPWR.n3873 0 0.00162f
C30630 VPWR.n3874 0 0.00151f
C30631 VPWR.n3875 0 0.0013f
C30632 VPWR.n3876 0 0.0014f
C30633 VPWR.n3877 0 0.00851f
C30634 VPWR.n3878 0 0.00493f
C30635 VPWR.n3879 0 0.0217f
C30636 VPWR.n3881 0 0.00208f
C30637 VPWR.n3882 0 0.00498f
C30638 VPWR.n3883 0 0.00891f
C30639 VPWR.n3884 0 0.00616f
C30640 VPWR.t12 0 0.068f
C30641 VPWR.n3885 0 0.0701f
C30642 VPWR.n3886 0 0.0483f
C30643 VPWR.n3887 0 0.0159f
C30644 VPWR.n3888 0 0.0421f
C30645 VPWR.n3889 0 0.0199f
C30646 VPWR.n3890 0 0.0535f
C30647 VPWR.n3891 0 0.0199f
C30648 VPWR.n3892 0 0.0626f
C30649 VPWR.n3893 0 0.0118f
C30650 VPWR.n3894 0 0.00994f
C30651 VPWR.n3895 0 0.0143f
C30652 VPWR.n3896 0 0.081f
C30653 VPWR.n3897 0 0.207f
C30654 VPWR.t320 0 0.073f
C30655 VPWR.n3898 0 0.207f
C30656 VPWR.n3899 0 0.0429f
C30657 VPWR.n3900 0 0.0143f
C30658 VPWR.n3901 0 0.0144f
C30659 VPWR.n3902 0 0.00994f
C30660 VPWR.n3903 0 0.0932f
C30661 VPWR.t15 0 0.068f
C30662 VPWR.n3904 0 0.0841f
C30663 VPWR.n3905 0 0.0722f
C30664 VPWR.n3906 0 0.0517f
C30665 VPWR.n3907 0 0.018f
C30666 VPWR.n3908 0 0.0118f
C30667 VPWR.n3909 0 0.0107f
C30668 VPWR.n3910 0 0.00918f
C30669 VPWR.n3911 0 0.181f
C30670 VPWR.n3912 0 0.0439f
C30671 VPWR.n3913 0 0.0363f
C30672 VPWR.n3914 0 0.0624f
C30673 VPWR.n3915 0 0.018f
C30674 VPWR.n3916 0 0.0199f
C30675 VPWR.n3917 0 0.0199f
C30676 VPWR.n3918 0 0.0118f
C30677 VPWR.n3919 0 0.0107f
C30678 VPWR.n3920 0 0.0758f
C30679 VPWR.n3921 0 0.0649f
C30680 VPWR.n3922 0 0.062f
C30681 VPWR.t358 0 0.068f
C30682 VPWR.n3923 0 0.0785f
C30683 VPWR.n3924 0 0.0391f
C30684 VPWR.n3925 0 0.0538f
C30685 VPWR.n3926 0 0.00655f
C30686 VPWR.t334 0 0.068f
C30687 VPWR.n3927 0 0.049f
C30688 VPWR.n3928 0 0.0722f
C30689 VPWR.n3929 0 0.0851f
C30690 VPWR.t47 0 0.068f
C30691 VPWR.n3930 0 0.0701f
C30692 VPWR.n3931 0 0.0791f
C30693 VPWR.n3932 0 0.018f
C30694 VPWR.n3933 0 0.023f
C30695 VPWR.n3934 0 0.0311f
C30696 VPWR.n3935 0 0.0118f
C30697 VPWR.n3936 0 0.105f
C30698 VPWR.n3937 0 0.0565f
C30699 VPWR.n3938 0 0.0851f
C30700 VPWR.n3939 0 0.00994f
C30701 VPWR.n3940 0 0.01f
C30702 VPWR.n3941 0 0.0948f
C30703 VPWR.n3942 0 0.0631f
C30704 VPWR.n3943 0 0.0117f
C30705 VPWR.n3944 0 0.0199f
C30706 VPWR.n3945 0 0.0173f
C30707 VPWR.n3946 0 0.0107f
C30708 VPWR.n3947 0 0.00994f
C30709 VPWR.n3948 0 0.00653f
C30710 VPWR.n3949 0 0.0935f
C30711 VPWR.n3950 0 0.0118f
C30712 VPWR.n3951 0 0.0199f
C30713 VPWR.n3952 0 0.0199f
C30714 VPWR.n3953 0 0.018f
C30715 VPWR.n3954 0 0.0608f
C30716 VPWR.n3955 0 0.00529f
C30717 VPWR.n3956 0 0.0199f
C30718 VPWR.n3957 0 0.00814f
C30719 VPWR.n3958 0 0.0199f
C30720 VPWR.n3959 0 0.018f
C30721 VPWR.n3960 0 0.0474f
C30722 VPWR.n3961 0 0.0818f
C30723 VPWR.n3962 0 0.0118f
C30724 VPWR.n3963 0 0.0199f
C30725 VPWR.n3964 0 0.0199f
C30726 VPWR.n3965 0 0.0522f
C30727 VPWR.n3966 0 0.0199f
C30728 VPWR.t51 0 0.0876f
C30729 VPWR.n3967 0 0.149f
C30730 VPWR.n3968 0 0.0199f
C30731 VPWR.n3969 0 0.0173f
C30732 VPWR.n3970 0 0.0682f
C30733 VPWR.n3971 0 0.0568f
C30734 VPWR.n3972 0 0.423f
C30735 VPWR.n3973 0 0.542f
C30736 VPWR.n3974 0 0.078f
C30737 VPWR.n3975 0 0.00291f
C30738 VPWR.n3976 0 0.00498f
C30739 VPWR.n3977 0 0.00281f
C30740 VPWR.n3978 0 0.00313f
C30741 VPWR.n3979 0 0.00989f
C30742 VPWR.n3980 0 0.00496f
C30743 VPWR.n3981 0 0.0217f
C30744 VPWR.n3983 0 0.00208f
C30745 VPWR.n3984 0 0.00483f
C30746 VPWR.n3985 0 0.00743f
C30747 VPWR.n3986 0 0.00259f
C30748 VPWR.n3987 0 0.00259f
C30749 VPWR.n3988 0 0.0183f
C30750 VPWR.t19 0 0.116f
C30751 VPWR.n3989 0 0.322f
C30752 VPWR.n3990 0 0.141f
C30753 VPWR.n3991 0 0.021f
C30754 VPWR.n3992 0 0.0605f
C30755 VPWR.n3993 0 0.0347f
C30756 VPWR.n3994 0 0.0771f
C30757 VPWR.n3995 0 0.0199f
C30758 VPWR.n3996 0 0.0766f
C30759 VPWR.n3997 0 0.0199f
C30760 VPWR.n3998 0 0.0118f
C30761 VPWR.n3999 0 0.0828f
C30762 VPWR.n4000 0 0.0907f
C30763 VPWR.n4001 0 0.018f
C30764 VPWR.n4002 0 0.0226f
C30765 VPWR.n4003 0 0.0199f
C30766 VPWR.n4004 0 0.0531f
C30767 VPWR.n4005 0 0.0199f
C30768 VPWR.n4006 0 0.0039f
C30769 VPWR.n4007 0 0.0265f
C30770 VPWR.n4008 0 0.18f
C30771 VPWR.n4009 0 0.0265f
C30772 VPWR.n4010 0 0.0525f
C30773 VPWR.n4011 0 0.0184f
C30774 VPWR.n4012 0 0.0276f
C30775 VPWR.n4013 0 0.00994f
C30776 VPWR.n4014 0 0.0547f
C30777 VPWR.n4015 0 0.0127f
C30778 VPWR.n4016 0 0.018f
C30779 VPWR.n4017 0 0.0698f
C30780 VPWR.n4018 0 0.0199f
C30781 VPWR.n4019 0 0.0626f
C30782 VPWR.n4020 0 0.0199f
C30783 VPWR.t170 0 0.0876f
C30784 VPWR.n4021 0 0.149f
C30785 VPWR.n4022 0 0.0199f
C30786 VPWR.n4023 0 0.0522f
C30787 VPWR.n4024 0 0.0199f
C30788 VPWR.n4025 0 0.0522f
C30789 VPWR.n4026 0 0.0199f
C30790 VPWR.n4027 0 0.0985f
C30791 VPWR.n4028 0 0.0199f
C30792 VPWR.n4029 0 0.0117f
C30793 VPWR.n4030 0 0.0107f
C30794 VPWR.t386 0 0.068f
C30795 VPWR.t105 0 0.0711f
C30796 VPWR.n4031 0 0.195f
C30797 VPWR.n4032 0 0.0877f
C30798 VPWR.n4033 0 0.0534f
C30799 VPWR.n4034 0 0.0837f
C30800 VPWR.t129 0 0.068f
C30801 VPWR.n4035 0 0.0471f
C30802 VPWR.n4036 0 0.0701f
C30803 VPWR.n4037 0 0.0391f
C30804 VPWR.t364 0 0.068f
C30805 VPWR.n4038 0 0.0701f
C30806 VPWR.n4039 0 0.0391f
C30807 VPWR.n4040 0 0.0656f
C30808 VPWR.n4041 0 0.0261f
C30809 VPWR.t201 0 0.0876f
C30810 VPWR.n4042 0 0.149f
C30811 VPWR.n4043 0 0.0118f
C30812 VPWR.n4044 0 0.0199f
C30813 VPWR.n4045 0 0.0199f
C30814 VPWR.n4046 0 0.0173f
C30815 VPWR.n4047 0 0.0107f
C30816 VPWR.n4048 0 0.0634f
C30817 VPWR.n4049 0 0.0375f
C30818 VPWR.n4050 0 0.0696f
C30819 VPWR.n4051 0 0.0199f
C30820 VPWR.n4052 0 0.00662f
C30821 VPWR.n4053 0 0.0199f
C30822 VPWR.n4054 0 0.0199f
C30823 VPWR.n4055 0 0.00494f
C30824 VPWR.n4056 0 0.0199f
C30825 VPWR.n4057 0 0.018f
C30826 VPWR.n4058 0 0.056f
C30827 VPWR.n4059 0 0.0739f
C30828 VPWR.n4060 0 0.0118f
C30829 VPWR.n4061 0 0.0199f
C30830 VPWR.n4062 0 0.018f
C30831 VPWR.n4063 0 0.01f
C30832 VPWR.n4064 0 0.0948f
C30833 VPWR.n4065 0 0.0631f
C30834 VPWR.n4066 0 0.0117f
C30835 VPWR.n4067 0 0.0199f
C30836 VPWR.n4068 0 0.0179f
C30837 VPWR.n4069 0 0.138f
C30838 VPWR.n4070 0 0.0166f
C30839 VPWR.n4071 0 0.0171f
C30840 VPWR.n4072 0 0.0265f
C30841 VPWR.n4073 0 0.0609f
C30842 VPWR.n4074 0 0.0199f
C30843 VPWR.n4075 0 0.00471f
C30844 VPWR.n4076 0 0.018f
C30845 VPWR.n4077 0 0.00994f
C30846 VPWR.n4078 0 0.0118f
C30847 VPWR.n4079 0 0.0199f
C30848 VPWR.n4080 0 0.0173f
C30849 VPWR.n4081 0 0.0391f
C30850 VPWR.n4082 0 0.0701f
C30851 VPWR.n4083 0 0.0791f
C30852 VPWR.n4084 0 0.248f
C30853 VPWR.n4085 0 0.0725f
C30854 VPWR.n4086 0 0.055f
C30855 VPWR.n4087 0 0.0012f
C30856 VPWR.n4088 0 0.00164f
C30857 VPWR.n4089 0 0.00162f
C30858 VPWR.n4090 0 0.0027f
C30859 VPWR.n4091 0 0.0013f
C30860 VPWR.n4092 0 0.0013f
C30861 VPWR.n4093 0 0.00861f
C30862 VPWR.n4094 0 0.00495f
C30863 VPWR.n4095 0 0.0217f
C30864 VPWR.n4096 0 0.00248f
C30865 VPWR.n4097 0 0.00344f
C30866 VPWR.n4098 0 0.00468f
C30867 VPWR.n4099 0 0.00323f
C30868 VPWR.n4100 0 0.00208f
C30869 VPWR.n4102 0 0.347f
C30870 VPWR.n4103 0 0.368f
C30871 VPWR.n4104 0 0.0412f
C30872 VPWR.n4105 0 0.00468f
C30873 VPWR.n4106 0 0.00323f
C30874 VPWR.n4107 0 0.00214f
C30875 VPWR.n4108 0 0.00344f
C30876 VPWR.n4109 0 0.00208f
C30877 VPWR.n4111 0 0.00484f
C30878 VPWR.n4112 0 1.32e-19
C30879 VPWR.n4113 0 0.00208f
C30880 VPWR.n4114 0 0.00126f
C30881 VPWR.n4115 0 0.00214f
C30882 VPWR.n4116 0 0.00237f
C30883 VPWR.n4117 0 0.00344f
C30884 VPWR.n4118 0 0.00323f
C30885 VPWR.n4119 0 0.00208f
C30886 VPWR.n4120 0 0.00302f
C30887 VPWR.n4121 0 0.00248f
C30888 VPWR.n4122 0 0.00173f
C30889 VPWR.n4123 0 0.0224f
C30890 VPWR.n4124 0 0.00194f
C30891 VPWR.n4125 0 0.0013f
C30892 VPWR.n4126 0 0.00108f
C30893 VPWR.n4127 0 0.00194f
C30894 VPWR.n4128 0 0.00173f
C30895 VPWR.n4129 0 0.0014f
C30896 VPWR.n4130 0 8.64e-19
C30897 VPWR.n4131 0 0.00108f
C30898 VPWR.n4132 0 0.00248f
C30899 VPWR.n4133 0 0.00378f
C30900 VPWR.n4134 0 0.00194f
C30901 VPWR.n4135 0 0.00173f
C30902 VPWR.n4136 0 0.0027f
C30903 VPWR.n4137 0 0.00119f
C30904 VPWR.n4138 0 0.00486f
C30905 VPWR.n4139 0 0.00389f
C30906 VPWR.n4140 0 0.00173f
C30907 VPWR.n4141 0 0.0027f
C30908 VPWR.t34 0 0.0876f
C30909 VPWR.n4142 0 0.0999f
C30910 VPWR.n4143 0 0.0261f
C30911 VPWR.t293 0 0.0726f
C30912 VPWR.n4144 0 0.263f
C30913 VPWR.n4145 0 0.013f
C30914 VPWR.n4146 0 0.0295f
C30915 VPWR.n4147 0 0.00119f
C30916 VPWR.n4148 0 0.00459f
C30917 VPWR.n4149 0 0.092f
C30918 VPWR.n4150 0 0.00804f
C30919 VPWR.n4151 0 0.0351f
C30920 VPWR.n4152 0 0.0605f
C30921 VPWR.t303 0 0.0417f
C30922 VPWR.n4153 0 0.0199f
C30923 VPWR.t278 0 0.0417f
C30924 VPWR.n4154 0 0.384f
C30925 VPWR.n4155 0 0.0619f
C30926 VPWR.n4156 0 0.0118f
C30927 VPWR.n4157 0 0.0558f
C30928 VPWR.n4158 0 0.0199f
C30929 VPWR.n4159 0 0.0791f
C30930 VPWR.n4160 0 0.0199f
C30931 VPWR.t39 0 0.068f
C30932 VPWR.n4161 0 0.0701f
C30933 VPWR.n4162 0 0.0665f
C30934 VPWR.n4163 0 0.0199f
C30935 VPWR.n4164 0 0.044f
C30936 VPWR.n4165 0 0.0199f
C30937 VPWR.n4166 0 0.0199f
C30938 VPWR.n4167 0 0.018f
C30939 VPWR.n4168 0 0.00529f
C30940 VPWR.n4169 0 0.0634f
C30941 VPWR.n4170 0 0.0118f
C30942 VPWR.n4171 0 0.0771f
C30943 VPWR.n4172 0 0.0199f
C30944 VPWR.n4173 0 0.0505f
C30945 VPWR.n4174 0 0.0199f
C30946 VPWR.t249 0 0.068f
C30947 VPWR.n4175 0 0.0701f
C30948 VPWR.n4176 0 0.0677f
C30949 VPWR.n4177 0 0.0199f
C30950 VPWR.n4178 0 0.0563f
C30951 VPWR.n4179 0 0.0199f
C30952 VPWR.n4180 0 0.018f
C30953 VPWR.n4181 0 0.00994f
C30954 VPWR.n4182 0 0.0555f
C30955 VPWR.n4183 0 0.0623f
C30956 VPWR.n4184 0 0.0118f
C30957 VPWR.n4185 0 0.0199f
C30958 VPWR.n4186 0 0.0199f
C30959 VPWR.t341 0 0.068f
C30960 VPWR.n4187 0 0.0695f
C30961 VPWR.n4188 0 0.0433f
C30962 VPWR.n4189 0 0.0701f
C30963 VPWR.n4190 0 0.0474f
C30964 VPWR.n4191 0 0.0179f
C30965 VPWR.n4192 0 0.01f
C30966 VPWR.n4193 0 0.00994f
C30967 VPWR.n4194 0 0.00994f
C30968 VPWR.n4195 0 0.0759f
C30969 VPWR.n4196 0 0.0917f
C30970 VPWR.n4197 0 0.0118f
C30971 VPWR.n4198 0 0.0391f
C30972 VPWR.n4199 0 0.018f
C30973 VPWR.n4200 0 0.00983f
C30974 VPWR.n4201 0 0.00184f
C30975 VPWR.n4202 0 0.0088f
C30976 VPWR.n4203 0 0.00496f
C30977 VPWR.n4204 0 0.00208f
C30978 VPWR.n4205 0 0.00126f
C30979 VPWR.n4206 0 0.00237f
C30980 VPWR.n4207 0 0.0108f
C30981 VPWR.n4208 0 0.94f
C30982 VPWR.n4209 0 0.0655f
C30983 VPWR.n4210 0 1.86f
C30984 VPWR.n4211 0 1.88f
C30985 VPWR.n4212 0 0.0657f
C30986 VPWR.n4213 0 1.87f
C30987 VPWR.n4214 0 0.376f
C30988 VPWR.n4216 0 0.0108f
C30989 VPWR.n4218 0 0.0115f
C30990 VPWR.n4219 0 2.61e-20
C30991 VPWR.n4220 0 0.00323f
C30992 VPWR.n4221 0 0.00344f
C30993 VPWR.n4222 0 0.00208f
C30994 VPWR.n4223 0 0.0108f
C30995 VPWR.n4224 0 0.00237f
C30996 VPWR.n4225 0 0.00126f
C30997 VPWR.n4226 0 0.00208f
C30998 VPWR.n4228 0 0.00743f
C30999 VPWR.n4229 0 0.00259f
C31000 VPWR.n4230 0 0.00259f
C31001 VPWR.n4231 0 0.00184f
C31002 VPWR.n4232 0 0.00292f
C31003 VPWR.n4233 0 6.5e-19
C31004 VPWR.n4234 0 0.00184f
C31005 VPWR.n4235 0 0.0027f
C31006 VPWR.n4236 0 0.0118f
C31007 VPWR.n4237 0 0.0199f
C31008 VPWR.n4238 0 0.0172f
C31009 VPWR.n4239 0 0.0632f
C31010 VPWR.n4240 0 0.0702f
C31011 VPWR.n4241 0 0.187f
C31012 VPWR.n4242 0 0.0386f
C31013 VPWR.t13 0 0.0726f
C31014 VPWR.n4243 0 0.0391f
C31015 VPWR.n4244 0 0.267f
C31016 VPWR.n4245 0 0.0391f
C31017 VPWR.n4246 0 0.0522f
C31018 VPWR.n4247 0 0.018f
C31019 VPWR.n4248 0 0.0199f
C31020 VPWR.n4249 0 0.0199f
C31021 VPWR.n4250 0 0.0917f
C31022 VPWR.n4251 0 0.0118f
C31023 VPWR.n4252 0 0.01f
C31024 VPWR.n4253 0 0.0623f
C31025 VPWR.n4254 0 0.0438f
C31026 VPWR.n4255 0 0.0179f
C31027 VPWR.n4256 0 0.0871f
C31028 VPWR.n4257 0 0.0199f
C31029 VPWR.t42 0 0.068f
C31030 VPWR.n4258 0 0.0701f
C31031 VPWR.n4259 0 0.0476f
C31032 VPWR.n4260 0 0.0199f
C31033 VPWR.n4261 0 0.0391f
C31034 VPWR.n4262 0 0.0199f
C31035 VPWR.n4263 0 0.0854f
C31036 VPWR.n4264 0 0.0199f
C31037 VPWR.n4265 0 0.0118f
C31038 VPWR.n4266 0 0.0853f
C31039 VPWR.n4267 0 0.0597f
C31040 VPWR.n4268 0 0.018f
C31041 VPWR.t225 0 0.068f
C31042 VPWR.n4269 0 0.0701f
C31043 VPWR.n4270 0 0.0479f
C31044 VPWR.n4271 0 0.0199f
C31045 VPWR.n4272 0 0.0391f
C31046 VPWR.n4273 0 0.0199f
C31047 VPWR.n4274 0 0.054f
C31048 VPWR.n4275 0 0.0199f
C31049 VPWR.n4276 0 0.0121f
C31050 VPWR.n4277 0 0.01f
C31051 VPWR.n4278 0 0.0957f
C31052 VPWR.n4279 0 0.0126f
C31053 VPWR.n4280 0 0.00983f
C31054 VPWR.n4281 0 0.0911f
C31055 VPWR.n4282 0 0.018f
C31056 VPWR.n4283 0 0.0199f
C31057 VPWR.n4284 0 0.0199f
C31058 VPWR.t41 0 0.068f
C31059 VPWR.n4285 0 0.0701f
C31060 VPWR.n4286 0 0.0391f
C31061 VPWR.n4287 0 0.125f
C31062 VPWR.n4288 0 0.0966f
C31063 VPWR.n4289 0 0.0118f
C31064 VPWR.n4290 0 0.0107f
C31065 VPWR.n4291 0 0.0406f
C31066 VPWR.n4292 0 0.0173f
C31067 VPWR.n4293 0 0.0126f
C31068 VPWR.n4294 0 0.00655f
C31069 VPWR.n4295 0 0.0634f
C31070 VPWR.n4296 0 0.0172f
C31071 VPWR.n4297 0 0.041f
C31072 VPWR.n4298 0 0.0199f
C31073 VPWR.t43 0 0.107f
C31074 VPWR.n4299 0 0.185f
C31075 VPWR.n4300 0 0.0386f
C31076 VPWR.n4301 0 0.0199f
C31077 VPWR.n4302 0 0.0822f
C31078 VPWR.n4303 0 0.0199f
C31079 VPWR.n4304 0 0.064f
C31080 VPWR.n4305 0 0.0199f
C31081 VPWR.n4306 0 0.0199f
C31082 VPWR.n4307 0 0.0199f
C31083 VPWR.n4308 0 0.0118f
C31084 VPWR.n4309 0 0.0619f
C31085 VPWR.n4310 0 0.0552f
C31086 VPWR.n4311 0 0.018f
C31087 VPWR.n4312 0 0.0434f
C31088 VPWR.n4313 0 0.0199f
C31089 VPWR.n4314 0 0.024f
C31090 VPWR.n4315 0 0.0199f
C31091 VPWR.n4316 0 0.107f
C31092 VPWR.n4317 0 0.0199f
C31093 VPWR.n4318 0 0.0925f
C31094 VPWR.n4319 0 0.0199f
C31095 VPWR.n4320 0 0.0199f
C31096 VPWR.n4321 0 0.0199f
C31097 VPWR.n4322 0 0.0119f
C31098 VPWR.n4323 0 0.00994f
C31099 VPWR.n4324 0 0.0065f
C31100 VPWR.n4325 0 0.086f
C31101 VPWR.n4326 0 0.018f
C31102 VPWR.n4327 0 0.0199f
C31103 VPWR.n4328 0 0.0199f
C31104 VPWR.n4329 0 0.0118f
C31105 VPWR.n4330 0 0.0985f
C31106 VPWR.t217 0 0.068f
C31107 VPWR.n4331 0 0.0965f
C31108 VPWR.n4332 0 0.0411f
C31109 VPWR.n4333 0 0.0722f
C31110 VPWR.n4334 0 0.0935f
C31111 VPWR.n4335 0 0.00994f
C31112 VPWR.n4336 0 0.018f
C31113 VPWR.n4337 0 0.0199f
C31114 VPWR.n4338 0 0.0118f
C31115 VPWR.n4339 0 0.00421f
C31116 VPWR.n4340 0 0.0013f
C31117 VPWR.n4341 0 0.0013f
C31118 VPWR.n4342 0 0.0027f
C31119 VPWR.n4343 0 0.00162f
C31120 VPWR.n4344 0 0.00205f
C31121 VPWR.n4345 0 0.00443f
C31122 VPWR.n4346 0 0.00302f
C31123 VPWR.n4347 0 0.00443f
C31124 VPWR.n4348 0 0.00281f
C31125 VPWR.n4349 0 8.64e-19
C31126 VPWR.n4350 0 0.00238f
C31127 VPWR.n4351 0 0.0321f
C31128 VPWR.n4352 0 0.00259f
C31129 VPWR.n4353 0 0.00173f
C31130 VPWR.n4354 0 4.32e-19
C31131 VPWR.n4355 0 0.00162f
C31132 VPWR.n4356 0 0.0168f
C31133 VPWR.n4357 0 0.0463f
C31134 VPWR.n4358 0 0.306f
C31135 VPWR.n4359 0 0.191f
C31136 VPWR.n4360 0 0.191f
C31137 VPWR.n4361 0 0.307f
C31138 VPWR.n4362 0 0.307f
C31139 VPWR.n4363 0 0.0376f
C31140 VPWR.n4364 0 0.00248f
C31141 VPWR.n4365 0 0.0014f
C31142 VPWR.n4366 0 0.00162f
C31143 VPWR.n4367 0 0.00216f
C31144 VPWR.n4368 0 0.00357f
C31145 VPWR.n4369 0 0.00248f
C31146 VPWR.n4370 0 0.0014f
C31147 VPWR.n4371 0 0.00335f
C31148 VPWR.n4372 0 0.00248f
C31149 VPWR.n4373 0 0.0014f
C31150 VPWR.n4374 0 8.64e-19
C31151 VPWR.n4375 0 0.00173f
C31152 VPWR.n4376 0 0.00497f
C31153 VPWR.n4377 0 0.00378f
C31154 VPWR.n4378 0 0.00162f
C31155 VPWR.n4379 0 0.00151f
C31156 VPWR.n4380 0 0.0013f
C31157 VPWR.n4381 0 0.0014f
C31158 VPWR.n4382 0 0.0085f
C31159 VPWR.n4383 0 0.00494f
C31160 VPWR.n4384 0 0.00208f
C31161 VPWR.n4385 0 0.00126f
C31162 VPWR.n4386 0 0.00237f
C31163 VPWR.n4387 0 0.116f
C31164 VPWR.n4388 0 2.61e-20
C31165 VPWR.n4389 0 0.0115f
C31166 VPWR.n4391 0 0.0108f
C31167 VPWR.n4393 0 0.376f
C31168 VPWR.n4394 0 0.381f
C31169 VPWR.n4396 0 0.00329f
C31170 VPWR.n4397 0 0.00208f
C31171 VPWR.n4398 0 0.00259f
C31172 VPWR.n4399 0 0.061f
C31173 VPWR.t292 0 0.116f
C31174 VPWR.n4400 0 0.00482f
C31175 VPWR.t356 0 0.0775f
C31176 VPWR.n4401 0 0.0197f
C31177 VPWR.t368 0 0.0417f
C31178 VPWR.t336 0 0.0417f
C31179 VPWR.n4402 0 0.384f
C31180 VPWR.n4403 0 0.019f
C31181 VPWR.n4404 0 0.0246f
C31182 VPWR.n4405 0 0.01f
C31183 VPWR.n4406 0 0.303f
C31184 VPWR.n4407 0 0.322f
C31185 VPWR.n4408 0 0.0953f
C31186 VPWR.n4409 0 0.018f
C31187 VPWR.n4410 0 0.0541f
C31188 VPWR.n4411 0 0.0199f
C31189 VPWR.n4412 0 0.13f
C31190 VPWR.n4413 0 0.0199f
C31191 VPWR.t0 0 0.069f
C31192 VPWR.n4414 0 0.0381f
C31193 VPWR.n4415 0 0.102f
C31194 VPWR.n4416 0 0.0305f
C31195 VPWR.n4417 0 0.0118f
C31196 VPWR.n4418 0 0.018f
C31197 VPWR.n4419 0 0.0199f
C31198 VPWR.n4420 0 0.0118f
C31199 VPWR.n4421 0 0.0856f
C31200 VPWR.n4422 0 0.0668f
C31201 VPWR.n4423 0 0.018f
C31202 VPWR.n4424 0 0.00394f
C31203 VPWR.n4425 0 0.0199f
C31204 VPWR.n4426 0 0.0329f
C31205 VPWR.n4427 0 0.0199f
C31206 VPWR.n4428 0 0.00482f
C31207 VPWR.n4429 0 0.0265f
C31208 VPWR.n4430 0 0.162f
C31209 VPWR.n4431 0 0.0265f
C31210 VPWR.n4432 0 0.0184f
C31211 VPWR.n4433 0 0.00552f
C31212 VPWR.n4434 0 0.049f
C31213 VPWR.n4435 0 0.018f
C31214 VPWR.t1 0 0.068f
C31215 VPWR.n4436 0 0.0818f
C31216 VPWR.n4437 0 0.049f
C31217 VPWR.n4438 0 0.0199f
C31218 VPWR.n4439 0 0.0561f
C31219 VPWR.n4440 0 0.0563f
C31220 VPWR.n4441 0 0.0186f
C31221 VPWR.n4442 0 0.00994f
C31222 VPWR.n4443 0 0.00184f
C31223 VPWR.n4444 0 0.015f
C31224 VPWR.n4445 0 0.0156f
C31225 VPWR.n4446 0 7.56e-19
C31226 VPWR.n4447 0 0.0376f
C31227 VPWR.n4448 0 0.00421f
C31228 VPWR.n4449 0 0.00248f
C31229 VPWR.n4450 0 5.4e-19
C31230 VPWR.n4451 0 0.00344f
C31231 VPWR.n4452 0 0.00248f
C31232 VPWR.n4453 0 0.00329f
C31233 VPWR.n4454 0 0.00208f
C31234 VPWR.n4455 0 0.00498f
C31235 VPWR.n4456 0 0.0118f
C31236 VPWR.n4457 0 0.00313f
C31237 VPWR.n4458 0 0.00397f
C31238 VPWR.n4459 0 0.00151f
C31239 VPWR.n4460 0 0.011f
C31240 VPWR.n4461 0 0.00162f
C31241 VPWR.n4462 0 0.00119f
C31242 VPWR.n4463 0 0.00184f
C31243 VPWR.n4464 0 0.00259f
C31244 VPWR.n4465 0 0.00119f
C31245 VPWR.t63 0 0.068f
C31246 VPWR.n4466 0 0.0266f
C31247 VPWR.n4467 0 0.0649f
C31248 VPWR.n4468 0 0.0399f
C31249 VPWR.n4469 0 0.00688f
C31250 VPWR.n4470 0 0.00521f
C31251 VPWR.n4471 0 0.0167f
C31252 VPWR.n4472 0 0.0504f
C31253 VPWR.t307 0 0.0737f
C31254 VPWR.n4473 0 0.299f
C31255 VPWR.n4474 0 0.307f
C31256 VPWR.n4475 0 0.0354f
C31257 VPWR.n4476 0 0.0386f
C31258 VPWR.n4477 0 0.0646f
C31259 VPWR.n4478 0 0.0535f
C31260 VPWR.n4479 0 0.0627f
C31261 VPWR.n4480 0 0.0027f
C31262 VPWR.n4481 0 0.00367f
C31263 VPWR.n4482 0 0.00281f
C31264 VPWR.n4483 0 0.381f
C31265 VPWR.n4484 0 0.00344f
C31266 VPWR.n4485 0 0.00248f
C31267 VPWR.n4486 0 0.00329f
C31268 VPWR.n4487 0 0.00208f
C31269 VPWR.n4488 0 0.00302f
C31270 VPWR.n4489 0 0.00248f
C31271 VPWR.n4490 0 0.00173f
C31272 VPWR.n4491 0 0.013f
C31273 VPWR.n4492 0 0.00194f
C31274 VPWR.n4493 0 0.0013f
C31275 VPWR.n4494 0 0.00108f
C31276 VPWR.n4495 0 0.00194f
C31277 VPWR.n4496 0 0.00173f
C31278 VPWR.n4497 0 0.0014f
C31279 VPWR.n4498 0 8.64e-19
C31280 VPWR.n4499 0 0.00108f
C31281 VPWR.n4500 0 0.00248f
C31282 VPWR.n4501 0 0.00378f
C31283 VPWR.n4502 0 0.00194f
C31284 VPWR.n4503 0 0.00173f
C31285 VPWR.n4504 0 0.0027f
C31286 VPWR.n4505 0 0.00119f
C31287 VPWR.n4506 0 0.00486f
C31288 VPWR.n4507 0 0.00389f
C31289 VPWR.n4508 0 0.00173f
C31290 VPWR.n4509 0 0.0027f
C31291 VPWR.t173 0 0.0711f
C31292 VPWR.n4510 0 0.195f
C31293 VPWR.n4511 0 0.00482f
C31294 VPWR.n4512 0 0.0261f
C31295 VPWR.n4513 0 0.0277f
C31296 VPWR.n4514 0 0.0636f
C31297 VPWR.n4515 0 0.00119f
C31298 VPWR.n4516 0 0.0382f
C31299 VPWR.n4517 0 0.0416f
C31300 VPWR.n4518 0 0.0287f
C31301 VPWR.n4519 0 0.0184f
C31302 VPWR.n4520 0 0.0596f
C31303 VPWR.t179 0 0.0417f
C31304 VPWR.n4521 0 0.239f
C31305 VPWR.t350 0 0.0417f
C31306 VPWR.t326 0 0.0417f
C31307 VPWR.n4522 0 0.383f
C31308 VPWR.n4523 0 0.0199f
C31309 VPWR.n4524 0 0.023f
C31310 VPWR.n4525 0 0.0312f
C31311 VPWR.n4526 0 0.0501f
C31312 VPWR.n4527 0 0.0754f
C31313 VPWR.n4528 0 0.0118f
C31314 VPWR.n4529 0 0.0617f
C31315 VPWR.n4530 0 0.0199f
C31316 VPWR.n4531 0 0.0571f
C31317 VPWR.n4532 0 0.0199f
C31318 VPWR.t57 0 0.068f
C31319 VPWR.n4533 0 0.0772f
C31320 VPWR.n4534 0 0.049f
C31321 VPWR.n4535 0 0.0199f
C31322 VPWR.n4536 0 0.034f
C31323 VPWR.n4537 0 0.0199f
C31324 VPWR.n4538 0 0.011f
C31325 VPWR.n4539 0 0.0199f
C31326 VPWR.n4540 0 0.043f
C31327 VPWR.n4541 0 0.0199f
C31328 VPWR.n4542 0 0.0179f
C31329 VPWR.n4543 0 0.01f
C31330 VPWR.n4544 0 0.0142f
C31331 VPWR.n4545 0 0.0811f
C31332 VPWR.n4546 0 0.0118f
C31333 VPWR.n4547 0 0.0199f
C31334 VPWR.n4548 0 0.0199f
C31335 VPWR.t197 0 0.068f
C31336 VPWR.n4549 0 0.0535f
C31337 VPWR.n4550 0 0.0391f
C31338 VPWR.n4551 0 0.0701f
C31339 VPWR.n4552 0 0.0487f
C31340 VPWR.n4553 0 0.018f
C31341 VPWR.n4554 0 0.0118f
C31342 VPWR.n4555 0 0.00451f
C31343 VPWR.n4556 0 0.0199f
C31344 VPWR.n4557 0 0.0199f
C31345 VPWR.n4558 0 0.018f
C31346 VPWR.n4559 0 0.00994f
C31347 VPWR.n4560 0 0.0299f
C31348 VPWR.n4561 0 0.0482f
C31349 VPWR.n4562 0 0.00994f
C31350 VPWR.n4563 0 0.00983f
C31351 VPWR.n4564 0 0.00184f
C31352 VPWR.n4565 0 0.00881f
C31353 VPWR.n4566 0 0.00496f
C31354 VPWR.n4567 0 0.381f
C31355 VPWR.n4568 0 0.00248f
C31356 VPWR.n4569 0 0.00344f
C31357 VPWR.n4570 0 0.00208f
C31358 VPWR.n4571 0 0.00323f
C31359 VPWR.n4572 0 0.00468f
C31360 VPWR.n4573 0 0.00323f
C31361 VPWR.n4574 0 0.00208f
C31362 VPWR.n4576 0 0.0216f
C31363 VPWR.n4578 0 0.00329f
C31364 VPWR.n4579 0 0.00208f
C31365 VPWR.n4580 0 0.00496f
C31366 VPWR.n4581 0 0.00859f
C31367 VPWR.n4582 0 0.0199f
C31368 VPWR.t286 0 0.116f
C31369 VPWR.n4583 0 0.322f
C31370 VPWR.t196 0 0.0737f
C31371 VPWR.n4584 0 0.299f
C31372 VPWR.n4585 0 0.01f
C31373 VPWR.n4586 0 0.00907f
C31374 VPWR.t167 0 0.116f
C31375 VPWR.n4587 0 0.0561f
C31376 VPWR.n4588 0 0.322f
C31377 VPWR.t232 0 0.068f
C31378 VPWR.n4589 0 0.0734f
C31379 VPWR.n4590 0 0.062f
C31380 VPWR.n4591 0 0.0322f
C31381 VPWR.t208 0 0.068f
C31382 VPWR.n4592 0 0.0329f
C31383 VPWR.n4593 0 0.0665f
C31384 VPWR.t77 0 0.0711f
C31385 VPWR.n4594 0 0.195f
C31386 VPWR.n4595 0 0.039f
C31387 VPWR.n4596 0 0.0213f
C31388 VPWR.n4597 0 0.0221f
C31389 VPWR.n4598 0 0.0179f
C31390 VPWR.n4599 0 0.00259f
C31391 VPWR.n4600 0 0.00421f
C31392 VPWR.n4601 0 0.00378f
C31393 VPWR.n4602 0 0.00162f
C31394 VPWR.n4603 0 0.0014f
C31395 VPWR.n4604 0 0.0014f
C31396 VPWR.n4605 0 0.00329f
C31397 VPWR.n4606 0 0.00208f
C31398 VPWR.n4607 0 0.381f
C31399 VPWR.n4608 0 0.381f
C31400 VPWR.n4609 0 0.00248f
C31401 VPWR.n4610 0 0.00344f
C31402 VPWR.n4611 0 0.00468f
C31403 VPWR.n4612 0 0.00323f
C31404 VPWR.n4613 0 0.00208f
C31405 VPWR.n4615 0 0.381f
C31406 VPWR.n4616 0 0.00323f
C31407 VPWR.n4617 0 0.00248f
C31408 VPWR.n4618 0 0.00344f
C31409 VPWR.n4619 0 0.00208f
C31410 VPWR.n4621 0 0.00329f
C31411 VPWR.n4622 0 0.00208f
C31412 VPWR.n4623 0 0.00302f
C31413 VPWR.n4624 0 0.00248f
C31414 VPWR.n4625 0 0.00173f
C31415 VPWR.n4626 0 0.0027f
C31416 VPWR.n4627 0 0.00248f
C31417 VPWR.n4628 0 0.00205f
C31418 VPWR.n4629 0 0.00162f
C31419 VPWR.n4630 0 0.00335f
C31420 VPWR.n4631 0 0.00421f
C31421 VPWR.n4632 0 0.00248f
C31422 VPWR.n4633 0 7.56e-19
C31423 VPWR.n4634 0 8.64e-19
C31424 VPWR.n4635 0 0.00108f
C31425 VPWR.n4636 0 0.00205f
C31426 VPWR.n4637 0 0.00248f
C31427 VPWR.n4638 0 0.0027f
C31428 VPWR.n4639 0 0.00302f
C31429 VPWR.n4640 0 0.00184f
C31430 VPWR.n4641 0 9.72e-19
C31431 VPWR.n4642 0 0.0014f
C31432 VPWR.n4643 0 8.64e-19
C31433 VPWR.n4644 0 0.00108f
C31434 VPWR.n4645 0 0.00248f
C31435 VPWR.n4646 0 0.00389f
C31436 VPWR.n4647 0 0.00357f
C31437 VPWR.n4648 0 0.00281f
C31438 VPWR.n4649 0 0.00162f
C31439 VPWR.n4650 0 0.00184f
C31440 VPWR.n4651 0 0.0535f
C31441 VPWR.t125 0 0.069f
C31442 VPWR.n4652 0 0.0429f
C31443 VPWR.n4653 0 0.0819f
C31444 VPWR.n4654 0 0.0964f
C31445 VPWR.t174 0 0.116f
C31446 VPWR.n4655 0 0.322f
C31447 VPWR.n4656 0 0.0799f
C31448 VPWR.n4657 0 0.0939f
C31449 VPWR.n4658 0 0.0459f
C31450 VPWR.t355 0 0.0973f
C31451 VPWR.n4659 0 0.219f
C31452 VPWR.n4660 0 0.0654f
C31453 VPWR.n4661 0 0.0198f
C31454 VPWR.n4662 0 0.018f
C31455 VPWR.n4663 0 0.0199f
C31456 VPWR.n4664 0 0.0118f
C31457 VPWR.n4665 0 0.0807f
C31458 VPWR.n4666 0 0.0661f
C31459 VPWR.n4667 0 0.018f
C31460 VPWR.n4668 0 0.0341f
C31461 VPWR.n4669 0 0.0199f
C31462 VPWR.n4670 0 0.00559f
C31463 VPWR.n4671 0 0.0199f
C31464 VPWR.n4672 0 0.00704f
C31465 VPWR.n4673 0 0.0199f
C31466 VPWR.n4674 0 0.00704f
C31467 VPWR.n4675 0 0.0199f
C31468 VPWR.n4676 0 0.0444f
C31469 VPWR.n4677 0 0.0199f
C31470 VPWR.n4678 0 0.0499f
C31471 VPWR.n4679 0 0.0199f
C31472 VPWR.n4680 0 0.0119f
C31473 VPWR.n4681 0 0.0233f
C31474 VPWR.n4682 0 0.0162f
C31475 VPWR.n4683 0 0.0179f
C31476 VPWR.n4684 0 0.00593f
C31477 VPWR.n4685 0 0.0126f
C31478 VPWR.n4686 0 0.0372f
C31479 VPWR.n4687 0 0.0394f
C31480 VPWR.n4688 0 0.0199f
C31481 VPWR.n4689 0 0.0118f
C31482 VPWR.n4690 0 0.00994f
C31483 VPWR.n4691 0 0.0305f
C31484 VPWR.n4692 0 0.104f
C31485 VPWR.n4693 0 0.0881f
C31486 VPWR.n4694 0 0.00983f
C31487 VPWR.n4695 0 0.0181f
C31488 VPWR.n4696 0 0.0118f
C31489 VPWR.n4697 0 0.112f
C31490 VPWR.n4698 0 0.0154f
C31491 VPWR.n4699 0 0.00335f
C31492 VPWR.n4700 0 0.00367f
C31493 VPWR.n4701 0 0.00281f
C31494 VPWR.n4702 0 0.00313f
C31495 VPWR.n4703 0 0.00989f
C31496 VPWR.n4704 0 0.00496f
C31497 VPWR.n4705 0 0.0217f
C31498 VPWR.n4706 0 0.00481f
C31499 VPWR.n4707 0 0.00744f
C31500 VPWR.n4708 0 0.00259f
C31501 VPWR.n4709 0 0.00259f
C31502 VPWR.n4710 0 0.00292f
C31503 VPWR.n4711 0 0.00184f
C31504 VPWR.n4712 0 0.00994f
C31505 VPWR.n4713 0 0.0275f
C31506 VPWR.n4714 0 0.0525f
C31507 VPWR.n4715 0 0.0115f
C31508 VPWR.n4716 0 0.00994f
C31509 VPWR.n4717 0 0.01f
C31510 VPWR.n4718 0 0.0892f
C31511 VPWR.n4719 0 0.00949f
C31512 VPWR.n4720 0 0.0179f
C31513 VPWR.n4721 0 0.0112f
C31514 VPWR.n4722 0 0.0199f
C31515 VPWR.n4723 0 0.0567f
C31516 VPWR.n4724 0 0.0199f
C31517 VPWR.n4725 0 0.0125f
C31518 VPWR.n4726 0 0.00769f
C31519 VPWR.t93 0 0.068f
C31520 VPWR.n4727 0 0.0654f
C31521 VPWR.n4728 0 0.0391f
C31522 VPWR.n4729 0 0.0701f
C31523 VPWR.n4730 0 0.049f
C31524 VPWR.n4731 0 0.0173f
C31525 VPWR.n4732 0 0.0199f
C31526 VPWR.n4733 0 0.0199f
C31527 VPWR.n4734 0 0.0118f
C31528 VPWR.n4735 0 0.0769f
C31529 VPWR.n4736 0 0.0518f
C31530 VPWR.n4737 0 0.018f
C31531 VPWR.n4738 0 0.0317f
C31532 VPWR.n4739 0 0.0199f
C31533 VPWR.n4740 0 0.0199f
C31534 VPWR.n4741 0 0.00529f
C31535 VPWR.t126 0 0.068f
C31536 VPWR.n4742 0 0.0617f
C31537 VPWR.n4743 0 0.0571f
C31538 VPWR.n4744 0 0.0772f
C31539 VPWR.n4745 0 0.049f
C31540 VPWR.n4746 0 0.018f
C31541 VPWR.n4747 0 0.0199f
C31542 VPWR.n4748 0 0.0199f
C31543 VPWR.n4749 0 0.0118f
C31544 VPWR.n4750 0 0.0754f
C31545 VPWR.n4751 0 0.0507f
C31546 VPWR.n4752 0 0.018f
C31547 VPWR.n4753 0 0.0309f
C31548 VPWR.n4754 0 0.0199f
C31549 VPWR.n4755 0 0.0568f
C31550 VPWR.n4756 0 0.0199f
C31551 VPWR.t300 0 0.068f
C31552 VPWR.n4757 0 0.0701f
C31553 VPWR.n4758 0 0.0481f
C31554 VPWR.n4759 0 0.0199f
C31555 VPWR.n4760 0 0.0391f
C31556 VPWR.n4761 0 0.0199f
C31557 VPWR.n4762 0 0.0547f
C31558 VPWR.n4763 0 0.0199f
C31559 VPWR.n4764 0 0.0885f
C31560 VPWR.n4765 0 0.0118f
C31561 VPWR.n4766 0 0.0107f
C31562 VPWR.n4767 0 0.0939f
C31563 VPWR.n4768 0 0.00907f
C31564 VPWR.n4769 0 0.0126f
C31565 VPWR.n4770 0 0.0181f
C31566 VPWR.n4771 0 0.0391f
C31567 VPWR.n4772 0 0.044f
C31568 VPWR.n4773 0 0.191f
C31569 VPWR.n4774 0 0.0243f
C31570 VPWR.n4775 0 0.0265f
C31571 VPWR.n4776 0 0.0919f
C31572 VPWR.n4777 0 0.0199f
C31573 VPWR.n4778 0 0.0535f
C31574 VPWR.n4779 0 0.0199f
C31575 VPWR.n4780 0 0.0118f
C31576 VPWR.n4781 0 0.0634f
C31577 VPWR.n4782 0 0.00529f
C31578 VPWR.n4783 0 0.018f
C31579 VPWR.n4784 0 0.0528f
C31580 VPWR.n4785 0 0.0199f
C31581 VPWR.n4786 0 0.00291f
C31582 VPWR.n4787 0 0.0118f
C31583 VPWR.n4788 0 0.0266f
C31584 VPWR.n4789 0 0.018f
C31585 VPWR.n4790 0 0.0429f
C31586 VPWR.n4791 0 0.0954f
C31587 VPWR.n4792 0 0.0309f
C31588 VPWR.n4793 0 0.0118f
C31589 VPWR.n4794 0 0.00994f
C31590 VPWR.n4795 0 0.025f
C31591 VPWR.n4796 0 0.0549f
C31592 VPWR.t101 0 0.0854f
C31593 VPWR.n4797 0 0.0688f
C31594 VPWR.n4798 0 0.0672f
C31595 VPWR.n4799 0 0.0479f
C31596 VPWR.n4800 0 0.018f
C31597 VPWR.n4801 0 0.045f
C31598 VPWR.n4802 0 0.0199f
C31599 VPWR.n4803 0 0.0199f
C31600 VPWR.n4804 0 0.0199f
C31601 VPWR.n4805 0 0.0117f
C31602 VPWR.n4806 0 0.00497f
C31603 VPWR.n4807 0 0.0013f
C31604 VPWR.n4808 0 0.0013f
C31605 VPWR.n4809 0 0.0027f
C31606 VPWR.n4810 0 0.00162f
C31607 VPWR.n4811 0 0.00205f
C31608 VPWR.n4812 0 0.00443f
C31609 VPWR.n4813 0 0.00302f
C31610 VPWR.n4814 0 0.00443f
C31611 VPWR.n4815 0 0.00281f
C31612 VPWR.n4816 0 8.64e-19
C31613 VPWR.n4817 0 0.00238f
C31614 VPWR.t315 0 0.068f
C31615 VPWR.n4818 0 0.0604f
C31616 VPWR.n4819 0 0.0224f
C31617 VPWR.n4820 0 0.00259f
C31618 VPWR.n4821 0 0.00173f
C31619 VPWR.n4822 0 4.32e-19
C31620 VPWR.n4823 0 0.00162f
C31621 VPWR.n4824 0 0.0168f
C31622 VPWR.n4825 0 0.0463f
C31623 VPWR.n4826 0 0.248f
C31624 VPWR.n4827 0 0.131f
C31625 VPWR.n4828 0 0.248f
C31626 VPWR.n4829 0 0.248f
C31627 VPWR.t2 0 0.116f
C31628 VPWR.n4830 0 0.266f
C31629 VPWR.n4831 0 0.204f
C31630 VPWR.n4832 0 0.0497f
C31631 VPWR.n4833 0 0.0107f
C31632 VPWR.n4834 0 0.0276f
C31633 VPWR.n4835 0 0.0117f
C31634 VPWR.n4836 0 0.018f
C31635 VPWR.n4837 0 0.00994f
C31636 VPWR.n4838 0 0.0544f
C31637 VPWR.n4839 0 0.0623f
C31638 VPWR.n4840 0 0.0118f
C31639 VPWR.n4841 0 0.0535f
C31640 VPWR.n4842 0 0.0199f
C31641 VPWR.n4843 0 0.0391f
C31642 VPWR.n4844 0 0.0199f
C31643 VPWR.t252 0 0.068f
C31644 VPWR.n4845 0 0.0701f
C31645 VPWR.n4846 0 0.0693f
C31646 VPWR.n4847 0 0.0199f
C31647 VPWR.n4848 0 0.018f
C31648 VPWR.n4849 0 0.00707f
C31649 VPWR.n4850 0 0.108f
C31650 VPWR.n4851 0 0.0118f
C31651 VPWR.n4852 0 0.0535f
C31652 VPWR.n4853 0 0.0199f
C31653 VPWR.n4854 0 0.0421f
C31654 VPWR.n4855 0 0.0199f
C31655 VPWR.t49 0 0.068f
C31656 VPWR.n4856 0 0.0701f
C31657 VPWR.n4857 0 0.049f
C31658 VPWR.n4858 0 0.0199f
C31659 VPWR.n4859 0 0.018f
C31660 VPWR.n4860 0 0.00994f
C31661 VPWR.n4861 0 0.0292f
C31662 VPWR.n4862 0 0.0627f
C31663 VPWR.n4863 0 0.0118f
C31664 VPWR.n4864 0 0.0199f
C31665 VPWR.n4865 0 0.0199f
C31666 VPWR.t251 0 0.068f
C31667 VPWR.n4866 0 0.0535f
C31668 VPWR.n4867 0 0.0391f
C31669 VPWR.n4868 0 0.0701f
C31670 VPWR.n4869 0 0.0474f
C31671 VPWR.n4870 0 0.018f
C31672 VPWR.n4871 0 0.00983f
C31673 VPWR.n4872 0 0.01f
C31674 VPWR.n4873 0 0.0373f
C31675 VPWR.n4874 0 0.0618f
C31676 VPWR.n4875 0 0.0118f
C31677 VPWR.n4876 0 0.0873f
C31678 VPWR.n4877 0 0.0199f
C31679 VPWR.n4878 0 0.0159f
C31680 VPWR.n4879 0 0.00616f
C31681 VPWR.n4880 0 0.00891f
C31682 VPWR.n4881 0 0.00119f
C31683 VPWR.n4882 0 0.00259f
C31684 VPWR.n4883 0 0.00184f
C31685 VPWR.n4884 0 0.00194f
C31686 VPWR.n4885 0 0.00248f
C31687 VPWR.n4886 0 0.00248f
C31688 VPWR.n4887 0 0.00227f
C31689 VPWR.n4888 0 8.64e-19
C31690 VPWR.n4889 0 0.00259f
C31691 VPWR.n4890 0 5.4e-19
C31692 VPWR.n4891 0 0.00248f
C31693 VPWR.n4892 0 0.00302f
C31694 VPWR.n4893 0 0.00119f
C31695 VPWR.n4894 0 0.00184f
C31696 VPWR.n4895 0 0.00248f
C31697 VPWR.n4896 0 0.0014f
C31698 VPWR.n4897 0 0.00162f
C31699 VPWR.n4898 0 0.00216f
C31700 VPWR.n4899 0 0.00357f
C31701 VPWR.n4900 0 0.00248f
C31702 VPWR.n4901 0 0.0014f
C31703 VPWR.n4902 0 0.00335f
C31704 VPWR.n4903 0 0.00248f
C31705 VPWR.n4904 0 0.0014f
C31706 VPWR.n4905 0 8.64e-19
C31707 VPWR.n4906 0 0.00173f
C31708 VPWR.n4907 0 0.00497f
C31709 VPWR.n4908 0 0.00378f
C31710 VPWR.n4909 0 0.00162f
C31711 VPWR.n4910 0 0.00151f
C31712 VPWR.n4911 0 0.0013f
C31713 VPWR.n4912 0 0.0014f
C31714 VPWR.n4913 0 0.00851f
C31715 VPWR.n4914 0 0.00493f
C31716 VPWR.n4915 0 0.0217f
C31717 VPWR.n4916 0 0.00248f
C31718 VPWR.n4917 0 0.00344f
C31719 VPWR.n4918 0 0.00208f
C31720 VPWR.n4919 0 0.00323f
C31721 VPWR.n4920 0 0.00468f
C31722 VPWR.n4921 0 0.00323f
C31723 VPWR.n4922 0 0.00208f
C31724 VPWR.n4924 0 0.381f
C31725 VPWR.n4925 0 0.381f
C31726 VPWR.n4926 0 0.381f
C31727 VPWR.n4927 0 0.381f
C31728 VPWR.n4928 0 0.00248f
C31729 VPWR.n4929 0 0.00344f
C31730 VPWR.n4930 0 0.00208f
C31731 VPWR.n4931 0 0.00323f
C31732 VPWR.n4932 0 0.00468f
C31733 VPWR.n4933 0 0.00323f
C31734 VPWR.n4934 0 0.00208f
C31735 VPWR.n4936 0 0.00329f
C31736 VPWR.n4937 0 0.00208f
C31737 VPWR.n4938 0 0.00259f
C31738 VPWR.t9 0 0.107f
C31739 VPWR.n4939 0 0.101f
C31740 VPWR.n4940 0 0.00994f
C31741 VPWR.t22 0 0.0711f
C31742 VPWR.n4941 0 0.195f
C31743 VPWR.n4942 0 0.0877f
C31744 VPWR.n4943 0 0.0534f
C31745 VPWR.n4944 0 0.0199f
C31746 VPWR.t373 0 0.0973f
C31747 VPWR.t120 0 0.0718f
C31748 VPWR.n4945 0 0.208f
C31749 VPWR.n4946 0 0.018f
C31750 VPWR.t277 0 0.0417f
C31751 VPWR.t246 0 0.0417f
C31752 VPWR.n4947 0 0.383f
C31753 VPWR.n4948 0 0.019f
C31754 VPWR.n4949 0 0.0191f
C31755 VPWR.n4950 0 0.0246f
C31756 VPWR.n4951 0 0.0198f
C31757 VPWR.n4952 0 0.0657f
C31758 VPWR.n4953 0 0.219f
C31759 VPWR.n4954 0 0.0779f
C31760 VPWR.n4955 0 0.057f
C31761 VPWR.n4956 0 0.114f
C31762 VPWR.n4957 0 0.0118f
C31763 VPWR.n4958 0 0.0107f
C31764 VPWR.n4959 0 0.00579f
C31765 VPWR.t143 0 0.068f
C31766 VPWR.n4960 0 0.0391f
C31767 VPWR.n4961 0 0.0701f
C31768 VPWR.n4962 0 0.0958f
C31769 VPWR.n4963 0 0.00918f
C31770 VPWR.n4964 0 0.018f
C31771 VPWR.n4965 0 0.0199f
C31772 VPWR.n4966 0 0.0118f
C31773 VPWR.n4967 0 0.0534f
C31774 VPWR.n4968 0 0.0882f
C31775 VPWR.n4969 0 0.0523f
C31776 VPWR.n4970 0 0.018f
C31777 VPWR.n4971 0 0.00513f
C31778 VPWR.n4972 0 0.0199f
C31779 VPWR.n4973 0 0.0118f
C31780 VPWR.n4974 0 0.0544f
C31781 VPWR.n4975 0 0.0903f
C31782 VPWR.n4976 0 0.0107f
C31783 VPWR.n4977 0 0.0173f
C31784 VPWR.n4978 0 0.0118f
C31785 VPWR.n4979 0 0.041f
C31786 VPWR.n4980 0 0.185f
C31787 VPWR.n4981 0 0.0386f
C31788 VPWR.n4982 0 0.018f
C31789 VPWR.n4983 0 0.0391f
C31790 VPWR.n4984 0 0.0199f
C31791 VPWR.t144 0 0.0726f
C31792 VPWR.n4985 0 0.267f
C31793 VPWR.n4986 0 0.0261f
C31794 VPWR.n4987 0 0.0357f
C31795 VPWR.n4988 0 0.0186f
C31796 VPWR.n4989 0 0.00994f
C31797 VPWR.n4990 0 0.00184f
C31798 VPWR.n4991 0 0.00482f
C31799 VPWR.n4992 0 0.0934f
C31800 VPWR.n4993 0 7.56e-19
C31801 VPWR.n4994 0 0.00194f
C31802 VPWR.n4995 0 8.64e-19
C31803 VPWR.n4996 0 0.00215f
C31804 VPWR.n4997 0 0.131f
C31805 VPWR.n4998 0 0.079f
C31806 VPWR.n4999 0 0.00113f
C31807 VPWR.n5000 0 0.00417f
C31808 VPWR.n5001 0 0.00421f
C31809 VPWR.n5002 0 0.00248f
C31810 VPWR.n5003 0 5.4e-19
C31811 VPWR.n5004 0 0.00259f
C31812 VPWR.n5005 0 0.00184f
C31813 VPWR.n5006 0 0.00194f
C31814 VPWR.n5007 0 0.00248f
C31815 VPWR.n5008 0 0.00248f
C31816 VPWR.n5009 0 0.00227f
C31817 VPWR.n5010 0 8.64e-19
C31818 VPWR.n5011 0 0.00259f
C31819 VPWR.n5012 0 5.4e-19
C31820 VPWR.n5013 0 0.00248f
C31821 VPWR.n5014 0 0.00302f
C31822 VPWR.n5015 0 0.00119f
C31823 VPWR.n5016 0 0.00184f
C31824 VPWR.n5017 0 0.00248f
C31825 VPWR.n5018 0 0.0014f
C31826 VPWR.n5019 0 0.00162f
C31827 VPWR.n5020 0 0.00216f
C31828 VPWR.n5021 0 0.00357f
C31829 VPWR.n5022 0 0.00248f
C31830 VPWR.n5023 0 0.0014f
C31831 VPWR.n5024 0 0.00335f
C31832 VPWR.n5025 0 0.00248f
C31833 VPWR.n5026 0 0.0014f
C31834 VPWR.n5027 0 8.64e-19
C31835 VPWR.n5028 0 0.00173f
C31836 VPWR.n5029 0 0.00497f
C31837 VPWR.n5030 0 0.00378f
C31838 VPWR.n5031 0 0.00162f
C31839 VPWR.n5032 0 0.00151f
C31840 VPWR.n5033 0 0.0013f
C31841 VPWR.n5034 0 0.0014f
C31842 VPWR.n5035 0 0.00851f
C31843 VPWR.n5036 0 0.00493f
C31844 VPWR.n5037 0 0.0217f
C31845 VPWR.n5039 0 0.00208f
C31846 VPWR.n5040 0 0.00498f
C31847 VPWR.n5041 0 0.00891f
C31848 VPWR.n5042 0 0.00616f
C31849 VPWR.n5043 0 0.00789f
C31850 VPWR.n5044 0 0.00544f
C31851 VPWR.t145 0 0.107f
C31852 VPWR.n5045 0 0.0386f
C31853 VPWR.n5046 0 0.185f
C31854 VPWR.n5047 0 0.0946f
C31855 VPWR.n5048 0 0.0671f
C31856 VPWR.n5049 0 0.0172f
C31857 VPWR.n5050 0 0.0199f
C31858 VPWR.n5051 0 0.0199f
C31859 VPWR.t48 0 0.0726f
C31860 VPWR.n5052 0 0.267f
C31861 VPWR.n5053 0 0.0391f
C31862 VPWR.n5054 0 0.0199f
C31863 VPWR.n5055 0 0.0391f
C31864 VPWR.n5056 0 0.0199f
C31865 VPWR.n5057 0 0.0118f
C31866 VPWR.n5058 0 0.118f
C31867 VPWR.n5059 0 0.01f
C31868 VPWR.n5060 0 0.103f
C31869 VPWR.n5061 0 0.0579f
C31870 VPWR.n5062 0 0.018f
C31871 VPWR.t87 0 0.068f
C31872 VPWR.n5063 0 0.085f
C31873 VPWR.n5064 0 0.0475f
C31874 VPWR.n5065 0 0.0199f
C31875 VPWR.n5066 0 0.0554f
C31876 VPWR.n5067 0 0.0199f
C31877 VPWR.n5068 0 0.0535f
C31878 VPWR.n5069 0 0.0199f
C31879 VPWR.n5070 0 0.0118f
C31880 VPWR.n5071 0 0.0679f
C31881 VPWR.n5072 0 0.0809f
C31882 VPWR.n5073 0 0.018f
C31883 VPWR.n5074 0 0.00856f
C31884 VPWR.n5075 0 0.0199f
C31885 VPWR.n5076 0 0.031f
C31886 VPWR.n5077 0 0.0199f
C31887 VPWR.n5078 0 0.0078f
C31888 VPWR.n5079 0 0.0199f
C31889 VPWR.n5080 0 0.0712f
C31890 VPWR.n5081 0 0.0199f
C31891 VPWR.n5082 0 0.0599f
C31892 VPWR.n5083 0 0.0199f
C31893 VPWR.n5084 0 0.0118f
C31894 VPWR.n5085 0 0.0321f
C31895 VPWR.t71 0 0.0876f
C31896 VPWR.n5086 0 0.0522f
C31897 VPWR.n5087 0 0.166f
C31898 VPWR.n5088 0 0.0731f
C31899 VPWR.n5089 0 0.018f
C31900 VPWR.n5090 0 0.0199f
C31901 VPWR.n5091 0 0.0199f
C31902 VPWR.n5092 0 0.0522f
C31903 VPWR.n5093 0 0.0199f
C31904 VPWR.n5094 0 0.0546f
C31905 VPWR.n5095 0 0.0199f
C31906 VPWR.n5096 0 0.0118f
C31907 VPWR.t23 0 0.068f
C31908 VPWR.n5097 0 0.0721f
C31909 VPWR.n5098 0 0.0179f
C31910 VPWR.n5099 0 0.0487f
C31911 VPWR.t171 0 0.114f
C31912 VPWR.n5100 0 0.472f
C31913 VPWR.n5101 0 0.111f
C31914 VPWR.t148 0 0.116f
C31915 VPWR.n5102 0 0.359f
C31916 VPWR.n5103 0 0.0935f
C31917 VPWR.n5104 0 0.018f
C31918 VPWR.t371 0 0.068f
C31919 VPWR.n5105 0 0.0722f
C31920 VPWR.n5106 0 0.0411f
C31921 VPWR.n5107 0 0.106f
C31922 VPWR.t74 0 0.068f
C31923 VPWR.n5108 0 0.0565f
C31924 VPWR.n5109 0 0.0335f
C31925 VPWR.t112 0 0.073f
C31926 VPWR.n5110 0 0.198f
C31927 VPWR.t8 0 0.0724f
C31928 VPWR.n5111 0 0.207f
C31929 VPWR.n5112 0 0.0429f
C31930 VPWR.n5113 0 0.0145f
C31931 VPWR.n5114 0 0.0133f
C31932 VPWR.n5115 0 0.0107f
C31933 VPWR.n5116 0 0.0656f
C31934 VPWR.n5117 0 0.105f
C31935 VPWR.n5118 0 0.0118f
C31936 VPWR.n5119 0 0.018f
C31937 VPWR.n5120 0 0.00994f
C31938 VPWR.n5121 0 0.0851f
C31939 VPWR.n5122 0 0.0701f
C31940 VPWR.n5123 0 0.0948f
C31941 VPWR.n5124 0 0.0118f
C31942 VPWR.n5125 0 0.0199f
C31943 VPWR.n5126 0 0.018f
C31944 VPWR.n5127 0 0.00994f
C31945 VPWR.n5128 0 0.0118f
C31946 VPWR.n5129 0 0.106f
C31947 VPWR.n5130 0 0.0565f
C31948 VPWR.n5131 0 0.09f
C31949 VPWR.n5132 0 0.00994f
C31950 VPWR.n5133 0 0.0435f
C31951 VPWR.n5134 0 0.0503f
C31952 VPWR.n5135 0 0.00907f
C31953 VPWR.n5136 0 0.142f
C31954 VPWR.n5137 0 0.0619f
C31955 VPWR.n5138 0 0.0118f
C31956 VPWR.n5139 0 0.018f
C31957 VPWR.n5140 0 0.0118f
C31958 VPWR.n5141 0 0.0173f
C31959 VPWR.n5142 0 0.0107f
C31960 VPWR.n5143 0 0.0387f
C31961 VPWR.n5144 0 0.179f
C31962 VPWR.n5145 0 0.131f
C31963 VPWR.n5146 0 0.0586f
C31964 VPWR.n5147 0 0.00291f
C31965 VPWR.n5148 0 0.00498f
C31966 VPWR.n5149 0 0.00281f
C31967 VPWR.n5150 0 0.00313f
C31968 VPWR.n5151 0 0.00989f
C31969 VPWR.n5152 0 0.00496f
C31970 VPWR.n5153 0 0.0217f
C31971 VPWR.n5154 0 0.00481f
C31972 VPWR.n5155 0 0.00744f
C31973 VPWR.n5156 0 0.00259f
C31974 VPWR.n5157 0 0.00259f
C31975 VPWR.n5158 0 0.00292f
C31976 VPWR.n5159 0 0.00184f
C31977 VPWR.n5160 0 0.00994f
C31978 VPWR.n5161 0 0.0261f
C31979 VPWR.n5162 0 0.0527f
C31980 VPWR.n5163 0 0.0196f
C31981 VPWR.n5164 0 0.0118f
C31982 VPWR.n5165 0 0.0634f
C31983 VPWR.n5166 0 0.0893f
C31984 VPWR.n5167 0 0.018f
C31985 VPWR.n5168 0 0.0213f
C31986 VPWR.n5169 0 0.0199f
C31987 VPWR.n5170 0 0.0118f
C31988 VPWR.n5171 0 0.0117f
C31989 VPWR.n5172 0 0.018f
C31990 VPWR.n5173 0 0.0979f
C31991 VPWR.n5174 0 0.0701f
C31992 VPWR.n5175 0 0.0391f
C31993 VPWR.n5176 0 0.0631f
C31994 VPWR.n5177 0 0.0108f
C31995 VPWR.n5178 0 0.00918f
C31996 VPWR.n5179 0 0.00994f
C31997 VPWR.n5180 0 0.149f
C31998 VPWR.n5181 0 0.0577f
C31999 VPWR.n5182 0 0.0522f
C32000 VPWR.n5183 0 0.0819f
C32001 VPWR.n5184 0 0.018f
C32002 VPWR.n5185 0 0.0199f
C32003 VPWR.n5186 0 0.0199f
C32004 VPWR.n5187 0 0.0118f
C32005 VPWR.n5188 0 0.0794f
C32006 VPWR.n5189 0 0.00655f
C32007 VPWR.n5190 0 0.018f
C32008 VPWR.n5191 0 0.00704f
C32009 VPWR.n5192 0 0.0199f
C32010 VPWR.n5193 0 0.00704f
C32011 VPWR.n5194 0 0.0199f
C32012 VPWR.n5195 0 0.0587f
C32013 VPWR.n5196 0 0.0199f
C32014 VPWR.n5197 0 0.0338f
C32015 VPWR.n5198 0 0.0199f
C32016 VPWR.n5199 0 0.00448f
C32017 VPWR.n5200 0 0.0199f
C32018 VPWR.n5201 0 0.112f
C32019 VPWR.n5202 0 0.0199f
C32020 VPWR.n5203 0 0.0117f
C32021 VPWR.n5204 0 0.00628f
C32022 VPWR.t177 0 0.068f
C32023 VPWR.n5205 0 0.0751f
C32024 VPWR.n5206 0 0.0427f
C32025 VPWR.n5207 0 0.0701f
C32026 VPWR.n5208 0 0.049f
C32027 VPWR.n5209 0 0.0181f
C32028 VPWR.n5210 0 0.0199f
C32029 VPWR.n5211 0 0.0199f
C32030 VPWR.n5212 0 0.0118f
C32031 VPWR.n5213 0 0.0107f
C32032 VPWR.t91 0 0.0876f
C32033 VPWR.t372 0 0.0726f
C32034 VPWR.n5214 0 0.267f
C32035 VPWR.n5215 0 0.0391f
C32036 VPWR.n5216 0 0.149f
C32037 VPWR.n5217 0 0.0615f
C32038 VPWR.n5218 0 0.0626f
C32039 VPWR.n5219 0 0.041f
C32040 VPWR.t70 0 0.0726f
C32041 VPWR.t172 0 0.107f
C32042 VPWR.n5220 0 0.185f
C32043 VPWR.n5221 0 0.0255f
C32044 VPWR.n5222 0 0.267f
C32045 VPWR.n5223 0 0.0391f
C32046 VPWR.n5224 0 0.00621f
C32047 VPWR.n5225 0 0.018f
C32048 VPWR.n5226 0 0.0199f
C32049 VPWR.n5227 0 0.0118f
C32050 VPWR.n5228 0 0.0199f
C32051 VPWR.n5229 0 0.0199f
C32052 VPWR.n5230 0 0.0911f
C32053 VPWR.n5231 0 0.018f
C32054 VPWR.n5232 0 0.00994f
C32055 VPWR.n5233 0 0.0118f
C32056 VPWR.n5234 0 0.0645f
C32057 VPWR.n5235 0 0.0867f
C32058 VPWR.n5236 0 0.0522f
C32059 VPWR.n5237 0 0.0522f
C32060 VPWR.n5238 0 0.0118f
C32061 VPWR.n5239 0 0.0199f
C32062 VPWR.n5240 0 0.0199f
C32063 VPWR.n5241 0 0.0173f
C32064 VPWR.n5242 0 0.00983f
C32065 VPWR.n5243 0 0.0634f
C32066 VPWR.n5244 0 0.00655f
C32067 VPWR.n5245 0 0.0126f
C32068 VPWR.n5246 0 0.0181f
C32069 VPWR.n5247 0 0.00704f
C32070 VPWR.n5248 0 0.00666f
C32071 VPWR.n5249 0 0.0117f
C32072 VPWR.n5250 0 0.0199f
C32073 VPWR.n5251 0 0.0173f
C32074 VPWR.n5252 0 0.0199f
C32075 VPWR.n5253 0 0.033f
C32076 VPWR.n5254 0 0.0199f
C32077 VPWR.n5255 0 0.0179f
C32078 VPWR.n5256 0 0.0788f
C32079 VPWR.n5257 0 0.0258f
C32080 VPWR.n5258 0 0.00994f
C32081 VPWR.n5259 0 0.0917f
C32082 VPWR.n5260 0 0.0118f
C32083 VPWR.n5261 0 0.0391f
C32084 VPWR.n5262 0 0.0199f
C32085 VPWR.n5263 0 0.0199f
C32086 VPWR.n5264 0 0.0199f
C32087 VPWR.n5265 0 0.0173f
C32088 VPWR.n5266 0 0.00994f
C32089 VPWR.n5267 0 0.0516f
C32090 VPWR.n5268 0 0.0461f
C32091 VPWR.n5269 0 0.129f
C32092 VPWR.n5270 0 0.424f
C32093 VPWR.n5271 0 0.0394f
C32094 VPWR.n5272 0 0.00212f
C32095 VPWR.n5273 0 0.00164f
C32096 VPWR.n5274 0 0.00162f
C32097 VPWR.n5275 0 0.0027f
C32098 VPWR.n5276 0 0.0013f
C32099 VPWR.n5277 0 0.0013f
C32100 VPWR.n5278 0 0.00859f
C32101 VPWR.n5279 0 0.00496f
C32102 VPWR.n5280 0 0.00208f
C32103 VPWR.n5282 0 0.0216f
C32104 VPWR.n5283 0 0.00248f
C32105 VPWR.n5284 0 0.00344f
C32106 VPWR.n5285 0 0.00208f
C32107 VPWR.n5286 0 0.00323f
C32108 VPWR.n5287 0 0.00468f
C32109 VPWR.n5288 0 0.00323f
C32110 VPWR.n5289 0 0.00208f
C32111 VPWR.n5291 0 0.381f
C32112 VPWR.n5292 0 0.381f
C32113 VPWR.n5293 0 0.00344f
C32114 VPWR.n5294 0 0.00248f
C32115 VPWR.n5295 0 0.00329f
C32116 VPWR.n5296 0 0.00208f
C32117 VPWR.n5297 0 0.00302f
C32118 VPWR.n5298 0 0.00248f
C32119 VPWR.n5299 0 0.00173f
C32120 VPWR.n5300 0 0.014f
C32121 VPWR.n5301 0 0.00194f
C32122 VPWR.n5302 0 0.0013f
C32123 VPWR.n5303 0 0.00108f
C32124 VPWR.n5304 0 0.00194f
C32125 VPWR.n5305 0 0.00173f
C32126 VPWR.n5306 0 0.0014f
C32127 VPWR.n5307 0 8.64e-19
C32128 VPWR.n5308 0 0.00108f
C32129 VPWR.n5309 0 0.00248f
C32130 VPWR.n5310 0 0.00378f
C32131 VPWR.n5311 0 0.00194f
C32132 VPWR.n5312 0 0.00173f
C32133 VPWR.n5313 0 0.0027f
C32134 VPWR.n5314 0 0.00119f
C32135 VPWR.n5315 0 0.00486f
C32136 VPWR.n5316 0 0.00389f
C32137 VPWR.n5317 0 0.00173f
C32138 VPWR.n5318 0 0.0027f
C32139 VPWR.t311 0 0.068f
C32140 VPWR.n5319 0 0.00482f
C32141 VPWR.n5320 0 0.0329f
C32142 VPWR.n5321 0 0.0702f
C32143 VPWR.n5322 0 0.0261f
C32144 VPWR.n5323 0 0.0564f
C32145 VPWR.n5324 0 0.00119f
C32146 VPWR.n5325 0 0.062f
C32147 VPWR.t312 0 0.0876f
C32148 VPWR.n5326 0 0.0641f
C32149 VPWR.n5327 0 0.162f
C32150 VPWR.n5328 0 0.0535f
C32151 VPWR.n5329 0 0.00386f
C32152 VPWR.n5330 0 0.0657f
C32153 VPWR.t376 0 0.0716f
C32154 VPWR.n5331 0 0.196f
C32155 VPWR.n5332 0 0.0771f
C32156 VPWR.n5333 0 0.0118f
C32157 VPWR.t106 0 0.0876f
C32158 VPWR.n5334 0 0.0559f
C32159 VPWR.t316 0 0.0417f
C32160 VPWR.t290 0 0.0417f
C32161 VPWR.n5335 0 0.107f
C32162 VPWR.n5336 0 0.0619f
C32163 VPWR.n5337 0 0.384f
C32164 VPWR.n5338 0 0.0199f
C32165 VPWR.n5339 0 0.0118f
C32166 VPWR.n5340 0 0.0199f
C32167 VPWR.n5341 0 0.0179f
C32168 VPWR.n5342 0 0.01f
C32169 VPWR.n5343 0 0.0522f
C32170 VPWR.n5344 0 0.134f
C32171 VPWR.n5345 0 0.0519f
C32172 VPWR.n5346 0 0.039f
C32173 VPWR.n5347 0 0.018f
C32174 VPWR.n5348 0 0.0164f
C32175 VPWR.n5349 0 0.0265f
C32176 VPWR.n5350 0 0.0179f
C32177 VPWR.n5351 0 0.01f
C32178 VPWR.n5352 0 0.0287f
C32179 VPWR.n5353 0 0.0631f
C32180 VPWR.n5354 0 0.0118f
C32181 VPWR.n5355 0 0.0535f
C32182 VPWR.n5356 0 0.0199f
C32183 VPWR.n5357 0 0.0522f
C32184 VPWR.n5358 0 0.0199f
C32185 VPWR.n5359 0 0.0199f
C32186 VPWR.n5360 0 0.0199f
C32187 VPWR.n5361 0 0.0173f
C32188 VPWR.n5362 0 0.0107f
C32189 VPWR.n5363 0 0.0516f
C32190 VPWR.n5364 0 0.00551f
C32191 VPWR.n5365 0 0.0199f
C32192 VPWR.n5366 0 0.00429f
C32193 VPWR.n5367 0 0.0199f
C32194 VPWR.n5368 0 0.018f
C32195 VPWR.n5369 0 0.0708f
C32196 VPWR.n5370 0 0.0701f
C32197 VPWR.n5371 0 0.0118f
C32198 VPWR.n5372 0 0.062f
C32199 VPWR.n5373 0 0.018f
C32200 VPWR.n5374 0 0.00983f
C32201 VPWR.n5375 0 0.00184f
C32202 VPWR.n5376 0 0.00881f
C32203 VPWR.n5377 0 0.00496f
C32204 VPWR.n5378 0 0.00329f
C32205 VPWR.n5379 0 0.00208f
C32206 VPWR.n5380 0 0.0027f
C32207 VPWR.n5381 0 0.00497f
C32208 VPWR.n5382 0 4.32e-19
C32209 VPWR.t200 0 0.0726f
C32210 VPWR.n5383 0 0.0391f
C32211 VPWR.n5384 0 0.267f
C32212 VPWR.n5385 0 0.0405f
C32213 VPWR.t68 0 0.116f
C32214 VPWR.n5386 0 0.00593f
C32215 VPWR.t175 0 0.0726f
C32216 VPWR.n5387 0 0.0312f
C32217 VPWR.n5388 0 0.0718f
C32218 VPWR.n5389 0 0.00367f
C32219 VPWR.n5390 0 0.00281f
C32220 VPWR.n5391 0 0.00162f
C32221 VPWR.n5392 0 0.00205f
C32222 VPWR.n5393 0 0.00443f
C32223 VPWR.n5394 0 0.00302f
C32224 VPWR.n5395 0 0.00443f
C32225 VPWR.n5396 0 0.00281f
C32226 VPWR.n5397 0 8.64e-19
C32227 VPWR.n5398 0 0.00238f
C32228 VPWR.n5399 0 0.0292f
C32229 VPWR.n5400 0 0.00259f
C32230 VPWR.n5401 0 0.00173f
C32231 VPWR.n5402 0 0.0312f
C32232 VPWR.n5403 0 0.129f
C32233 VPWR.n5404 0 0.307f
C32234 VPWR.n5405 0 0.0107f
C32235 VPWR.t46 0 0.116f
C32236 VPWR.n5406 0 0.322f
C32237 VPWR.n5407 0 0.0793f
C32238 VPWR.n5408 0 0.0231f
C32239 VPWR.n5409 0 0.00398f
C32240 VPWR.n5410 0 0.00259f
C32241 VPWR.n5411 0 0.00298f
C32242 VPWR.n5412 0 0.00421f
C32243 VPWR.n5413 0 0.00378f
C32244 VPWR.n5414 0 0.00162f
C32245 VPWR.n5415 0 0.0014f
C32246 VPWR.n5416 0 0.0027f
C32247 VPWR.n5417 0 0.00248f
C32248 VPWR.n5418 0 0.00205f
C32249 VPWR.n5419 0 0.00352f
C32250 VPWR.n5420 0 0.00162f
C32251 VPWR.n5421 0 0.0013f
C32252 VPWR.n5422 0 0.00357f
C32253 VPWR.n5423 0 0.00389f
C32254 VPWR.n5424 0 0.00248f
C32255 VPWR.n5425 0 0.00108f
C32256 VPWR.n5426 0 8.64e-19
C32257 VPWR.n5427 0 0.00302f
C32258 VPWR.n5428 0 0.00248f
C32259 VPWR.n5429 0 0.00173f
C32260 VPWR.n5430 0 7.56e-19
C32261 VPWR.n5431 0 0.00184f
C32262 VPWR.n5432 0 0.00302f
C32263 VPWR.n5433 0 0.0027f
C32264 VPWR.n5434 0 0.00248f
C32265 VPWR.n5435 0 0.00205f
C32266 VPWR.n5436 0 0.00108f
C32267 VPWR.n5437 0 8.64e-19
C32268 VPWR.n5438 0 7.56e-19
C32269 VPWR.n5439 0 0.00248f
C32270 VPWR.n5440 0 0.00421f
C32271 VPWR.n5441 0 0.00335f
C32272 VPWR.n5442 0 0.00162f
C32273 VPWR.n5443 0 0.0014f
C32274 VPWR.n5444 0 0.00208f
C32275 VPWR.n5445 0 0.00344f
C32276 VPWR.n5446 0 0.00248f
C32277 VPWR.n5447 0 0.00329f
C32278 VPWR.n5448 0 0.00208f
C32279 VPWR.n5449 0 0.00483f
C32280 VPWR.n5450 0 0.00743f
C32281 VPWR.n5451 0 0.00259f
C32282 VPWR.n5452 0 0.00259f
C32283 VPWR.n5453 0 0.0149f
C32284 VPWR.n5454 0 0.00292f
C32285 VPWR.n5455 0 0.0308f
C32286 VPWR.n5456 0 0.00184f
C32287 VPWR.n5457 0 0.00176f
C32288 VPWR.n5458 0 0.00994f
C32289 VPWR.t86 0 0.0726f
C32290 VPWR.n5459 0 0.245f
C32291 VPWR.n5460 0 0.0186f
C32292 VPWR.n5461 0 0.0196f
C32293 VPWR.n5462 0 0.0118f
C32294 VPWR.n5463 0 0.0148f
C32295 VPWR.n5464 0 0.0341f
C32296 VPWR.n5465 0 0.018f
C32297 VPWR.n5466 0 0.00559f
C32298 VPWR.n5467 0 0.0199f
C32299 VPWR.n5468 0 0.00704f
C32300 VPWR.n5469 0 0.0199f
C32301 VPWR.n5470 0 0.0454f
C32302 VPWR.n5471 0 0.0199f
C32303 VPWR.n5472 0 0.0592f
C32304 VPWR.n5473 0 0.0199f
C32305 VPWR.n5474 0 0.0265f
C32306 VPWR.n5475 0 0.0199f
C32307 VPWR.n5476 0 0.0687f
C32308 VPWR.n5477 0 0.0199f
C32309 VPWR.n5478 0 0.0117f
C32310 VPWR.n5479 0 0.0162f
C32311 VPWR.n5480 0 0.00704f
C32312 VPWR.n5481 0 0.0181f
C32313 VPWR.t80 0 0.0726f
C32314 VPWR.n5482 0 0.245f
C32315 VPWR.n5483 0 0.00528f
C32316 VPWR.n5484 0 0.0199f
C32317 VPWR.n5485 0 0.00528f
C32318 VPWR.n5486 0 0.0199f
C32319 VPWR.n5487 0 0.0118f
C32320 VPWR.n5488 0 0.00994f
C32321 VPWR.n5489 0 0.0119f
C32322 VPWR.n5490 0 0.0356f
C32323 VPWR.n5491 0 0.018f
C32324 VPWR.n5492 0 0.04f
C32325 VPWR.n5493 0 0.0199f
C32326 VPWR.n5494 0 0.00525f
C32327 VPWR.n5495 0 0.0118f
C32328 VPWR.n5496 0 0.0382f
C32329 VPWR.n5497 0 0.0548f
C32330 VPWR.n5498 0 0.0394f
C32331 VPWR.n5499 0 0.0657f
C32332 VPWR.n5500 0 0.0199f
C32333 VPWR.n5501 0 0.0649f
C32334 VPWR.n5502 0 0.0199f
C32335 VPWR.n5503 0 0.0118f
C32336 VPWR.n5504 0 0.0855f
C32337 VPWR.n5505 0 0.0386f
C32338 VPWR.t389 0 0.068f
C32339 VPWR.n5506 0 0.0751f
C32340 VPWR.n5507 0 0.0427f
C32341 VPWR.n5508 0 0.0701f
C32342 VPWR.n5509 0 0.0475f
C32343 VPWR.n5510 0 0.0173f
C32344 VPWR.n5511 0 0.0199f
C32345 VPWR.n5512 0 0.0199f
C32346 VPWR.n5513 0 0.0749f
C32347 VPWR.n5514 0 0.0118f
C32348 VPWR.n5515 0 0.0165f
C32349 VPWR.n5516 0 0.018f
C32350 VPWR.n5517 0 0.0555f
C32351 VPWR.n5518 0 0.0199f
C32352 VPWR.n5519 0 0.0254f
C32353 VPWR.n5520 0 0.0199f
C32354 VPWR.n5521 0 0.00704f
C32355 VPWR.n5522 0 0.0199f
C32356 VPWR.n5523 0 0.0118f
C32357 VPWR.n5524 0 0.00528f
C32358 VPWR.n5525 0 0.245f
C32359 VPWR.n5526 0 0.00528f
C32360 VPWR.n5527 0 0.018f
C32361 VPWR.n5528 0 0.0118f
C32362 VPWR.n5529 0 0.0265f
C32363 VPWR.n5530 0 0.094f
C32364 VPWR.n5531 0 0.322f
C32365 VPWR.n5532 0 0.0429f
C32366 VPWR.n5533 0 0.018f
C32367 VPWR.n5534 0 0.0199f
C32368 VPWR.n5535 0 0.0199f
C32369 VPWR.n5536 0 0.0118f
C32370 VPWR.n5537 0 0.0634f
C32371 VPWR.n5538 0 0.00521f
C32372 VPWR.n5539 0 0.018f
C32373 VPWR.n5540 0 0.0859f
C32374 VPWR.n5541 0 0.0199f
C32375 VPWR.n5542 0 0.028f
C32376 VPWR.n5543 0 0.0199f
C32377 VPWR.n5544 0 0.0118f
C32378 VPWR.n5545 0 0.00656f
C32379 VPWR.n5546 0 0.0286f
C32380 VPWR.n5547 0 0.018f
C32381 VPWR.n5548 0 0.00883f
C32382 VPWR.n5549 0 0.0199f
C32383 VPWR.t117 0 0.0726f
C32384 VPWR.n5550 0 0.245f
C32385 VPWR.n5551 0 0.00528f
C32386 VPWR.n5552 0 0.0199f
C32387 VPWR.n5553 0 0.0118f
C32388 VPWR.n5554 0 0.00689f
C32389 VPWR.n5555 0 0.00352f
C32390 VPWR.n5556 0 0.00162f
C32391 VPWR.n5557 0 0.0027f
C32392 VPWR.n5558 0 0.0013f
C32393 VPWR.n5559 0 0.0013f
C32394 VPWR.n5560 0 0.00861f
C32395 VPWR.n5561 0 0.00495f
C32396 VPWR.n5562 0 0.416f
C32397 VPWR.n5564 0 0.00344f
C32398 VPWR.n5565 0 0.00248f
C32399 VPWR.n5566 0 0.00329f
C32400 VPWR.n5567 0 0.00208f
C32401 VPWR.n5568 0 0.00443f
C32402 VPWR.n5569 0 0.00302f
C32403 VPWR.n5570 0 0.00248f
C32404 VPWR.n5571 0 0.00173f
C32405 VPWR.n5572 0 0.00367f
C32406 VPWR.n5573 0 0.00194f
C32407 VPWR.n5574 0 0.0017f
C32408 VPWR.n5575 0 6.82e-19
C32409 VPWR.n5576 0 0.00194f
C32410 VPWR.n5577 0 0.00173f
C32411 VPWR.n5578 0 0.0014f
C32412 VPWR.n5579 0 8.64e-19
C32413 VPWR.n5580 0 0.00108f
C32414 VPWR.n5581 0 0.00248f
C32415 VPWR.n5582 0 0.00378f
C32416 VPWR.n5583 0 0.00194f
C32417 VPWR.n5584 0 0.00173f
C32418 VPWR.n5585 0 0.0027f
C32419 VPWR.n5586 0 0.00119f
C32420 VPWR.n5587 0 0.00486f
C32421 VPWR.n5588 0 0.00389f
C32422 VPWR.n5589 0 0.00173f
C32423 VPWR.n5590 0 0.0027f
C32424 VPWR.n5591 0 0.00119f
C32425 VPWR.t176 0 0.0737f
C32426 VPWR.n5592 0 0.299f
C32427 VPWR.n5593 0 0.0457f
C32428 VPWR.n5594 0 0.062f
C32429 VPWR.n5595 0 0.0619f
C32430 VPWR.t276 0 0.0417f
C32431 VPWR.t245 0 0.0417f
C32432 VPWR.n5596 0 0.384f
C32433 VPWR.n5597 0 0.0197f
C32434 VPWR.n5598 0 0.0118f
C32435 VPWR.n5599 0 0.018f
C32436 VPWR.n5600 0 0.0535f
C32437 VPWR.n5601 0 0.0528f
C32438 VPWR.n5602 0 0.0118f
C32439 VPWR.n5603 0 0.0819f
C32440 VPWR.n5604 0 0.0199f
C32441 VPWR.t349 0 0.0876f
C32442 VPWR.n5605 0 0.149f
C32443 VPWR.n5606 0 0.0199f
C32444 VPWR.n5607 0 0.0691f
C32445 VPWR.n5608 0 0.0199f
C32446 VPWR.n5609 0 0.0553f
C32447 VPWR.n5610 0 0.0199f
C32448 VPWR.n5611 0 0.00775f
C32449 VPWR.n5612 0 0.0199f
C32450 VPWR.n5613 0 0.018f
C32451 VPWR.n5614 0 0.00529f
C32452 VPWR.n5615 0 0.0753f
C32453 VPWR.n5616 0 0.0118f
C32454 VPWR.n5617 0 0.0671f
C32455 VPWR.n5618 0 0.0199f
C32456 VPWR.n5619 0 0.0391f
C32457 VPWR.n5620 0 0.0199f
C32458 VPWR.t296 0 0.068f
C32459 VPWR.n5621 0 0.0929f
C32460 VPWR.n5622 0 0.0597f
C32461 VPWR.n5623 0 0.0199f
C32462 VPWR.n5624 0 0.0199f
C32463 VPWR.n5625 0 0.00429f
C32464 VPWR.n5626 0 0.0199f
C32465 VPWR.n5627 0 0.018f
C32466 VPWR.n5628 0 0.0605f
C32467 VPWR.n5629 0 0.0324f
C32468 VPWR.n5630 0 0.071f
C32469 VPWR.n5631 0 0.0118f
C32470 VPWR.n5632 0 0.0199f
C32471 VPWR.n5633 0 0.0199f
C32472 VPWR.t254 0 0.116f
C32473 VPWR.n5634 0 0.322f
C32474 VPWR.n5635 0 0.0668f
C32475 VPWR.n5636 0 0.0926f
C32476 VPWR.n5637 0 0.0447f
C32477 VPWR.n5638 0 0.018f
C32478 VPWR.n5639 0 0.0128f
C32479 VPWR.n5640 0 0.0161f
C32480 VPWR.n5641 0 0.00881f
C32481 VPWR.n5642 0 0.00496f
C32482 VPWR.n5643 0 0.0217f
C32483 VPWR.n5644 0 0.00495f
C32484 VPWR.n5645 0 0.00208f
C32485 VPWR.n5646 0 0.00329f
C32486 VPWR.n5647 0 0.00248f
C32487 VPWR.n5648 0 0.00344f
C32488 VPWR.n5649 0 0.00208f
C32489 VPWR.n5650 0 0.00323f
C32490 VPWR.n5651 0 0.00468f
C32491 VPWR.n5652 0 0.00323f
C32492 VPWR.n5653 0 0.00208f
C32493 VPWR.n5655 0 0.381f
C32494 VPWR.n5656 0 0.381f
C32495 VPWR.n5657 0 0.00248f
C32496 VPWR.n5658 0 0.00344f
C32497 VPWR.n5659 0 0.00323f
C32498 VPWR.n5660 0 0.00208f
C32499 VPWR.n5662 0 0.00329f
C32500 VPWR.n5663 0 0.00208f
C32501 VPWR.n5664 0 0.00119f
C32502 VPWR.n5665 0 0.0119f
C32503 VPWR.n5666 0 0.00194f
C32504 VPWR.n5667 0 0.0013f
C32505 VPWR.n5668 0 6.5e-19
C32506 VPWR.n5669 0 0.00108f
C32507 VPWR.n5670 0 0.00352f
C32508 VPWR.n5671 0 0.00194f
C32509 VPWR.n5672 0 0.00173f
C32510 VPWR.n5673 0 0.00302f
C32511 VPWR.n5674 0 0.00248f
C32512 VPWR.n5675 0 0.00173f
C32513 VPWR.n5676 0 0.0027f
C32514 VPWR.n5677 0 0.00173f
C32515 VPWR.n5678 0 0.00194f
C32516 VPWR.n5679 0 0.00378f
C32517 VPWR.n5680 0 0.00248f
C32518 VPWR.n5681 0 0.00108f
C32519 VPWR.n5682 0 8.64e-19
C32520 VPWR.n5683 0 6.48e-19
C32521 VPWR.n5684 0 0.00454f
C32522 VPWR.n5685 0 0.00389f
C32523 VPWR.n5686 0 0.00173f
C32524 VPWR.n5687 0 0.0027f
C32525 VPWR.n5688 0 0.00398f
C32526 VPWR.n5689 0 0.00119f
C32527 VPWR.n5690 0 0.0108f
C32528 VPWR.n5691 0 0.067f
C32529 VPWR.n5692 0 0.114f
C32530 VPWR.n5693 0 0.0809f
C32531 VPWR.t224 0 0.0417f
C32532 VPWR.n5694 0 0.0208f
C32533 VPWR.t335 0 0.0417f
C32534 VPWR.n5695 0 0.383f
C32535 VPWR.t390 0 0.0774f
C32536 VPWR.t282 0 0.0774f
C32537 VPWR.n5696 0 0.501f
C32538 VPWR.n5697 0 0.0299f
C32539 VPWR.n5698 0 0.0394f
C32540 VPWR.n5699 0 0.00429f
C32541 VPWR.n5700 0 0.0199f
C32542 VPWR.n5701 0 0.018f
C32543 VPWR.n5702 0 0.00524f
C32544 VPWR.n5703 0 0.119f
C32545 VPWR.n5704 0 0.0118f
C32546 VPWR.n5705 0 0.1f
C32547 VPWR.n5706 0 0.0199f
C32548 VPWR.n5707 0 0.0199f
C32549 VPWR.n5708 0 0.0199f
C32550 VPWR.n5709 0 0.0199f
C32551 VPWR.n5710 0 0.0389f
C32552 VPWR.t160 0 0.1f
C32553 VPWR.n5711 0 0.125f
C32554 VPWR.t20 0 0.0876f
C32555 VPWR.n5712 0 0.0973f
C32556 VPWR.n5713 0 0.0973f
C32557 VPWR.n5714 0 0.167f
C32558 VPWR.n5715 0 0.0876f
C32559 VPWR.n5716 0 0.0585f
C32560 VPWR.n5717 0 0.0173f
C32561 VPWR.n5718 0 0.0107f
C32562 VPWR.n5719 0 0.00352f
C32563 VPWR.n5720 0 0.0306f
C32564 VPWR.n5721 0 0.00659f
C32565 VPWR.n5722 0 0.0118f
C32566 VPWR.n5723 0 0.0903f
C32567 VPWR.n5724 0 0.0199f
C32568 VPWR.n5725 0 0.0179f
C32569 VPWR.n5726 0 0.01f
C32570 VPWR.n5727 0 0.0112f
C32571 VPWR.n5728 0 0.0231f
C32572 VPWR.n5729 0 0.0118f
C32573 VPWR.n5730 0 0.00704f
C32574 VPWR.n5731 0 0.0199f
C32575 VPWR.n5732 0 0.00528f
C32576 VPWR.n5733 0 0.0199f
C32577 VPWR.t159 0 0.105f
C32578 VPWR.n5734 0 0.376f
C32579 VPWR.n5735 0 0.00528f
C32580 VPWR.n5736 0 0.0199f
C32581 VPWR.n5737 0 0.0152f
C32582 VPWR.n5738 0 0.018f
C32583 VPWR.n5739 0 0.0201f
C32584 VPWR.n5740 0 0.00983f
C32585 VPWR.n5741 0 0.00184f
C32586 VPWR.n5742 0 0.00882f
C32587 VPWR.n5743 0 0.00496f
C32588 VPWR.n5744 0 0.0217f
C32589 VPWR.n5745 0 0.00468f
C32590 VPWR.n5746 0 0.00323f
C32591 VPWR.n5747 0 0.00248f
C32592 VPWR.n5748 0 0.00344f
C32593 VPWR.n5749 0 0.00208f
C32594 VPWR.n5751 0 0.0605f
C32595 VPWR.n5752 0 2.85f
C32596 VPWR.n5753 0 0.37f
C32597 VPWR.n5754 0 0.331f
C32598 VPWR.n5755 0 0.00248f
C32599 VPWR.n5756 0 0.00344f
C32600 VPWR.n5757 0 0.00208f
C32601 VPWR.n5758 0 0.00323f
C32602 VPWR.n5759 0 0.00468f
C32603 VPWR.n5760 0 0.00323f
C32604 VPWR.n5761 0 0.00208f
C32605 VPWR.n5763 0 0.0216f
C32606 VPWR.n5765 0 0.00329f
C32607 VPWR.n5766 0 0.00208f
C32608 VPWR.n5767 0 0.00496f
C32609 VPWR.n5768 0 0.00859f
C32610 VPWR.n5769 0 0.00443f
C32611 VPWR.n5770 0 0.00281f
C32612 VPWR.n5771 0 0.00367f
C32613 VPWR.n5772 0 0.00281f
C32614 VPWR.n5773 0 0.00238f
C32615 VPWR.n5774 0 8.64e-19
C32616 VPWR.n5775 0 0.00302f
C32617 VPWR.n5776 0 0.00443f
C32618 VPWR.n5777 0 0.00205f
C32619 VPWR.n5778 0 0.00162f
C32620 VPWR.n5779 0 0.0027f
C32621 VPWR.n5780 0 0.0013f
C32622 VPWR.n5781 0 0.0013f
C32623 VPWR.n5782 0 0.0027f
C32624 VPWR.n5783 0 0.00162f
C32625 VPWR.n5784 0 0.00164f
C32626 VPWR.n5785 0 0.0012f
C32627 VPWR.n5786 0 0.0604f
C32628 VPWR.n5787 0 0.0725f
C32629 VPWR.n5788 0 0.307f
C32630 VPWR.n5789 0 0.13f
C32631 VPWR.n5790 0 0.131f
C32632 VPWR.n5791 0 0.307f
C32633 VPWR.n5792 0 0.05f
C32634 VPWR.n5793 0 0.00248f
C32635 VPWR.n5794 0 0.0014f
C32636 VPWR.n5795 0 0.00162f
C32637 VPWR.n5796 0 0.00216f
C32638 VPWR.n5797 0 0.00357f
C32639 VPWR.n5798 0 0.00248f
C32640 VPWR.n5799 0 0.0014f
C32641 VPWR.n5800 0 0.00335f
C32642 VPWR.n5801 0 0.00248f
C32643 VPWR.n5802 0 0.0014f
C32644 VPWR.n5803 0 8.64e-19
C32645 VPWR.n5804 0 0.00173f
C32646 VPWR.n5805 0 0.00497f
C32647 VPWR.n5806 0 0.00378f
C32648 VPWR.n5807 0 0.00162f
C32649 VPWR.n5808 0 0.00151f
C32650 VPWR.n5809 0 0.0013f
C32651 VPWR.n5810 0 0.0014f
C32652 VPWR.n5811 0 0.00851f
C32653 VPWR.n5812 0 0.00493f
C32654 VPWR.n5813 0 0.0217f
C32655 VPWR.n5814 0 0.00248f
C32656 VPWR.n5815 0 0.00344f
C32657 VPWR.n5816 0 0.00208f
C32658 VPWR.n5817 0 0.00323f
C32659 VPWR.n5818 0 0.00468f
C32660 VPWR.n5819 0 0.00323f
C32661 VPWR.n5820 0 0.00208f
C32662 VPWR.n5822 0 0.331f
C32663 VPWR.n5823 0 3.04f
C32664 VPWR.n5824 0 0.0605f
C32665 VPWR.n5825 0 0.416f
C32666 VPWR.n5827 0 0.00498f
C32667 VPWR.n5828 0 0.00208f
C32668 VPWR.n5829 0 0.00329f
C32669 VPWR.n5830 0 0.00248f
C32670 VPWR.n5831 0 0.00344f
C32671 VPWR.n5832 0 0.00208f
C32672 VPWR.n5833 0 0.00323f
C32673 VPWR.n5834 0 0.00468f
C32674 VPWR.n5835 0 0.00323f
C32675 VPWR.n5836 0 0.00208f
C32676 VPWR.n5837 0 0.00344f
C32677 VPWR.n5838 0 0.00248f
C32678 VPWR.n5839 0 0.00329f
C32679 VPWR.n5840 0 0.00208f
C32680 VPWR.n5841 0 0.00493f
C32681 VPWR.n5842 0 0.0217f
C32682 VPWR.n5844 0 0.381f
C32683 VPWR.n5845 0 0.381f
C32684 VPWR.n5846 0 0.00248f
C32685 VPWR.n5847 0 0.00344f
C32686 VPWR.n5848 0 0.00208f
C32687 VPWR.n5849 0 0.00323f
C32688 VPWR.n5850 0 0.00468f
C32689 VPWR.n5851 0 0.00323f
C32690 VPWR.n5852 0 0.00208f
C32691 VPWR.n5854 0 0.00329f
C32692 VPWR.n5855 0 0.00208f
C32693 VPWR.n5856 0 0.00259f
C32694 VPWR.n5857 0 0.074f
C32695 VPWR.n5858 0 0.0537f
C32696 VPWR.t69 0 0.0718f
C32697 VPWR.n5859 0 0.208f
C32698 VPWR.n5860 0 0.113f
C32699 VPWR.n5861 0 0.0312f
C32700 VPWR.t237 0 0.116f
C32701 VPWR.n5862 0 0.00994f
C32702 VPWR.t212 0 0.0407f
C32703 VPWR.t38 0 0.068f
C32704 VPWR.n5863 0 0.0475f
C32705 VPWR.n5864 0 0.0701f
C32706 VPWR.n5865 0 0.222f
C32707 VPWR.t233 0 0.0417f
C32708 VPWR.t352 0 0.0417f
C32709 VPWR.n5866 0 0.384f
C32710 VPWR.n5867 0 0.019f
C32711 VPWR.n5868 0 0.0319f
C32712 VPWR.n5869 0 0.0199f
C32713 VPWR.n5870 0 0.0118f
C32714 VPWR.n5871 0 0.044f
C32715 VPWR.n5872 0 0.213f
C32716 VPWR.n5873 0 0.322f
C32717 VPWR.n5874 0 0.121f
C32718 VPWR.n5875 0 0.0207f
C32719 VPWR.n5876 0 0.00994f
C32720 VPWR.n5877 0 0.0646f
C32721 VPWR.n5878 0 0.0515f
C32722 VPWR.n5879 0 0.018f
C32723 VPWR.n5880 0 0.0118f
C32724 VPWR.n5881 0 0.00994f
C32725 VPWR.n5882 0 0.0107f
C32726 VPWR.n5883 0 0.0812f
C32727 VPWR.n5884 0 0.107f
C32728 VPWR.n5885 0 0.0591f
C32729 VPWR.n5886 0 0.0173f
C32730 VPWR.t238 0 0.1f
C32731 VPWR.n5887 0 0.13f
C32732 VPWR.n5888 0 0.0876f
C32733 VPWR.n5889 0 0.0487f
C32734 VPWR.n5890 0 0.0199f
C32735 VPWR.n5891 0 0.0199f
C32736 VPWR.n5892 0 0.0199f
C32737 VPWR.n5893 0 0.0199f
C32738 VPWR.t56 0 0.107f
C32739 VPWR.n5894 0 0.208f
C32740 VPWR.n5895 0 0.0719f
C32741 VPWR.n5896 0 0.0973f
C32742 VPWR.n5897 0 0.0987f
C32743 VPWR.n5898 0 0.176f
C32744 VPWR.n5899 0 0.0118f
C32745 VPWR.n5900 0 0.0121f
C32746 VPWR.n5901 0 0.00966f
C32747 VPWR.n5902 0 0.00119f
C32748 VPWR.n5903 0 0.00162f
C32749 VPWR.n5904 0 0.00119f
C32750 VPWR.n5905 0 0.00162f
C32751 VPWR.n5906 0 0.00151f
C32752 VPWR.n5907 0 0.00313f
C32753 VPWR.n5908 0 0.00421f
C32754 VPWR.n5909 0 0.00248f
C32755 VPWR.n5910 0 5.4e-19
C32756 VPWR.n5911 0 0.00259f
C32757 VPWR.n5912 0 0.00184f
C32758 VPWR.n5913 0 0.00194f
C32759 VPWR.n5914 0 0.00248f
C32760 VPWR.n5915 0 0.00248f
C32761 VPWR.n5916 0 0.00227f
C32762 VPWR.n5917 0 8.64e-19
C32763 VPWR.n5918 0 0.00259f
C32764 VPWR.n5919 0 5.4e-19
C32765 VPWR.n5920 0 0.00248f
C32766 VPWR.n5921 0 0.00302f
C32767 VPWR.n5922 0 0.00119f
C32768 VPWR.n5923 0 0.00184f
C32769 VPWR.n5924 0 0.129f
C32770 VPWR.n5925 0 0.133f
C32771 VPWR.n5926 0 0.00601f
C32772 VPWR.n5927 0 0.00561f
C32773 VPWR.n5928 0 0.0276f
C32774 VPWR.n5929 0 0.0256f
C32775 VPWR.t226 0 0.0949f
C32776 VPWR.n5930 0 0.101f
C32777 VPWR.n5931 0 0.0371f
C32778 VPWR.n5932 0 0.00681f
C32779 VPWR.n5933 0 0.0616f
C32780 VPWR.n5934 0 0.00248f
C32781 VPWR.n5935 0 0.0014f
C32782 VPWR.n5936 0 0.00162f
C32783 VPWR.n5937 0 0.00216f
C32784 VPWR.n5938 0 0.00357f
C32785 VPWR.n5939 0 0.00248f
C32786 VPWR.n5940 0 0.0014f
C32787 VPWR.n5941 0 0.00335f
C32788 VPWR.n5942 0 0.00248f
C32789 VPWR.n5943 0 0.0014f
C32790 VPWR.n5944 0 8.64e-19
C32791 VPWR.n5945 0 0.00173f
C32792 VPWR.n5946 0 0.00497f
C32793 VPWR.n5947 0 0.00378f
C32794 VPWR.n5948 0 0.00162f
C32795 VPWR.n5949 0 0.00151f
C32796 VPWR.n5950 0 0.0013f
C32797 VPWR.n5951 0 0.0014f
C32798 VPWR.n5952 0 0.00851f
C32799 VPWR.n5953 0 0.00493f
C32800 VPWR.n5954 0 0.0217f
C32801 VPWR.n5956 0 0.00208f
C32802 VPWR.n5957 0 0.00498f
C32803 VPWR.n5958 0 0.00891f
C32804 VPWR.n5959 0 0.00616f
C32805 VPWR.n5960 0 0.02f
C32806 VPWR.n5961 0 0.0214f
C32807 VPWR.n5962 0 0.0333f
C32808 VPWR.n5963 0 0.0576f
C32809 VPWR.n5964 0 0.0357f
C32810 VPWR.n5965 0 0.0159f
C32811 VPWR.n5966 0 0.0475f
C32812 VPWR.n5967 0 0.018f
C32813 VPWR.n5968 0 0.21f
C32814 VPWR.n5969 0 0.0148f
C32815 VPWR.n5970 0 0.0265f
C32816 VPWR.t104 0 0.0721f
C32817 VPWR.n5971 0 0.196f
C32818 VPWR.n5972 0 0.0523f
C32819 VPWR.n5973 0 0.0164f
C32820 VPWR.n5974 0 0.0275f
C32821 VPWR.n5975 0 0.0531f
C32822 VPWR.n5976 0 0.0259f
C32823 VPWR.n5977 0 0.0518f
C32824 VPWR.n5978 0 0.0118f
C32825 VPWR.n5979 0 0.0437f
C32826 VPWR.n5980 0 0.0668f
C32827 VPWR.n5981 0 0.0926f
C32828 VPWR.n5982 0 0.054f
C32829 VPWR.n5983 0 0.018f
C32830 VPWR.n5984 0 0.0199f
C32831 VPWR.n5985 0 0.0199f
C32832 VPWR.n5986 0 0.0118f
C32833 VPWR.n5987 0 0.01f
C32834 VPWR.n5988 0 0.0281f
C32835 VPWR.n5989 0 0.00909f
C32836 VPWR.n5990 0 0.0179f
C32837 VPWR.n5991 0 0.0667f
C32838 VPWR.n5992 0 0.0199f
C32839 VPWR.t267 0 0.068f
C32840 VPWR.n5993 0 0.0701f
C32841 VPWR.n5994 0 0.0476f
C32842 VPWR.n5995 0 0.0199f
C32843 VPWR.n5996 0 0.0627f
C32844 VPWR.n5997 0 0.0199f
C32845 VPWR.n5998 0 0.0649f
C32846 VPWR.n5999 0 0.0199f
C32847 VPWR.n6000 0 0.0118f
C32848 VPWR.n6001 0 0.0107f
C32849 VPWR.n6002 0 0.0436f
C32850 VPWR.t213 0 0.068f
C32851 VPWR.n6003 0 0.0535f
C32852 VPWR.n6004 0 0.0391f
C32853 VPWR.n6005 0 0.0701f
C32854 VPWR.n6006 0 0.049f
C32855 VPWR.n6007 0 0.0173f
C32856 VPWR.n6008 0 0.0199f
C32857 VPWR.n6009 0 0.0199f
C32858 VPWR.n6010 0 0.00656f
C32859 VPWR.n6011 0 0.0822f
C32860 VPWR.n6012 0 0.0118f
C32861 VPWR.n6013 0 0.018f
C32862 VPWR.n6014 0 0.0516f
C32863 VPWR.n6015 0 0.0199f
C32864 VPWR.n6016 0 0.0491f
C32865 VPWR.n6017 0 0.0199f
C32866 VPWR.n6018 0 0.0118f
C32867 VPWR.n6019 0 0.0107f
C32868 VPWR.n6020 0 0.0341f
C32869 VPWR.n6021 0 0.00559f
C32870 VPWR.n6022 0 0.0173f
C32871 VPWR.n6023 0 0.00704f
C32872 VPWR.n6024 0 0.0199f
C32873 VPWR.n6025 0 0.00528f
C32874 VPWR.n6026 0 0.0199f
C32875 VPWR.t158 0 0.105f
C32876 VPWR.n6027 0 0.376f
C32877 VPWR.n6028 0 0.0289f
C32878 VPWR.n6029 0 0.0199f
C32879 VPWR.n6030 0 0.0184f
C32880 VPWR.n6031 0 0.0199f
C32881 VPWR.n6032 0 0.0118f
C32882 VPWR.n6033 0 0.0206f
C32883 VPWR.n6034 0 0.0189f
C32884 VPWR.n6035 0 0.018f
C32885 VPWR.n6036 0 0.00704f
C32886 VPWR.n6037 0 0.0199f
C32887 VPWR.n6038 0 0.00704f
C32888 VPWR.n6039 0 0.0199f
C32889 VPWR.n6040 0 0.0456f
C32890 VPWR.n6041 0 0.0199f
C32891 VPWR.n6042 0 0.0433f
C32892 VPWR.n6043 0 0.0199f
C32893 VPWR.n6044 0 0.0273f
C32894 VPWR.n6045 0 0.0199f
C32895 VPWR.n6046 0 0.0513f
C32896 VPWR.n6047 0 0.0199f
C32897 VPWR.n6048 0 0.0117f
C32898 VPWR.n6049 0 0.01f
C32899 VPWR.n6050 0 0.0057f
C32900 VPWR.n6051 0 0.00528f
C32901 VPWR.n6052 0 0.018f
C32902 VPWR.t140 0 0.0726f
C32903 VPWR.n6053 0 0.245f
C32904 VPWR.n6054 0 0.00352f
C32905 VPWR.n6055 0 0.0199f
C32906 VPWR.n6056 0 0.0118f
C32907 VPWR.n6057 0 0.00482f
C32908 VPWR.n6058 0 0.00352f
C32909 VPWR.n6059 0 0.00335f
C32910 VPWR.n6060 0 0.00367f
C32911 VPWR.n6061 0 0.00281f
C32912 VPWR.n6062 0 0.00313f
C32913 VPWR.n6063 0 0.00989f
C32914 VPWR.n6064 0 0.00496f
C32915 VPWR.n6065 0 0.0217f
C32916 VPWR.n6066 0 0.00248f
C32917 VPWR.n6067 0 0.00344f
C32918 VPWR.n6068 0 0.00323f
C32919 VPWR.n6069 0 0.00468f
C32920 VPWR.n6070 0 0.00323f
C32921 VPWR.n6071 0 0.00208f
C32922 VPWR.n6073 0 0.381f
C32923 VPWR.n6074 0 0.381f
C32924 VPWR.n6076 0 0.00208f
C32925 VPWR.n6077 0 0.00483f
C32926 VPWR.n6078 0 0.00743f
C32927 VPWR.n6079 0 0.00259f
C32928 VPWR.n6080 0 0.00259f
C32929 VPWR.n6081 0 0.00292f
C32930 VPWR.n6082 0 0.00184f
C32931 VPWR.n6083 0 0.00994f
C32932 VPWR.t281 0 0.107f
C32933 VPWR.n6084 0 0.0254f
C32934 VPWR.n6085 0 0.206f
C32935 VPWR.n6086 0 0.0719f
C32936 VPWR.n6087 0 0.0196f
C32937 VPWR.n6088 0 0.0973f
C32938 VPWR.n6089 0 0.0199f
C32939 VPWR.n6090 0 0.0987f
C32940 VPWR.n6091 0 0.0199f
C32941 VPWR.n6092 0 0.18f
C32942 VPWR.n6093 0 0.0118f
C32943 VPWR.n6094 0 0.0143f
C32944 VPWR.n6095 0 0.0546f
C32945 VPWR.t97 0 0.068f
C32946 VPWR.n6096 0 0.0782f
C32947 VPWR.n6097 0 0.0411f
C32948 VPWR.n6098 0 0.0723f
C32949 VPWR.n6099 0 0.0981f
C32950 VPWR.n6100 0 0.018f
C32951 VPWR.n6101 0 0.0199f
C32952 VPWR.n6102 0 0.0199f
C32953 VPWR.n6103 0 0.0118f
C32954 VPWR.n6104 0 0.154f
C32955 VPWR.n6105 0 0.0245f
C32956 VPWR.n6106 0 0.0265f
C32957 VPWR.n6107 0 0.0682f
C32958 VPWR.n6108 0 0.0199f
C32959 VPWR.n6109 0 0.0535f
C32960 VPWR.n6110 0 0.0199f
C32961 VPWR.n6111 0 0.0118f
C32962 VPWR.n6112 0 0.0634f
C32963 VPWR.n6113 0 0.00655f
C32964 VPWR.n6114 0 0.018f
C32965 VPWR.n6115 0 0.0621f
C32966 VPWR.n6116 0 0.0199f
C32967 VPWR.n6117 0 0.0118f
C32968 VPWR.n6118 0 0.0201f
C32969 VPWR.t322 0 0.068f
C32970 VPWR.n6119 0 0.0535f
C32971 VPWR.n6120 0 0.0513f
C32972 VPWR.n6121 0 0.0929f
C32973 VPWR.n6122 0 0.049f
C32974 VPWR.n6123 0 0.018f
C32975 VPWR.n6124 0 0.0199f
C32976 VPWR.n6125 0 0.0199f
C32977 VPWR.n6126 0 0.0619f
C32978 VPWR.n6127 0 0.0118f
C32979 VPWR.n6128 0 0.0107f
C32980 VPWR.t253 0 0.068f
C32981 VPWR.n6129 0 0.0668f
C32982 VPWR.n6130 0 0.0473f
C32983 VPWR.n6131 0 0.0701f
C32984 VPWR.n6132 0 0.0713f
C32985 VPWR.n6133 0 0.0173f
C32986 VPWR.n6134 0 0.0199f
C32987 VPWR.n6135 0 0.0199f
C32988 VPWR.n6136 0 0.0465f
C32989 VPWR.n6137 0 0.103f
C32990 VPWR.n6138 0 0.0118f
C32991 VPWR.n6139 0 0.018f
C32992 VPWR.n6140 0 0.0199f
C32993 VPWR.n6141 0 0.0199f
C32994 VPWR.n6142 0 0.0631f
C32995 VPWR.t295 0 0.068f
C32996 VPWR.n6143 0 0.0927f
C32997 VPWR.n6144 0 0.0701f
C32998 VPWR.n6145 0 0.0948f
C32999 VPWR.n6146 0 0.00994f
C33000 VPWR.n6147 0 0.018f
C33001 VPWR.n6148 0 0.0199f
C33002 VPWR.n6149 0 0.0117f
C33003 VPWR.n6150 0 0.0629f
C33004 VPWR.t119 0 0.068f
C33005 VPWR.n6151 0 0.0916f
C33006 VPWR.n6152 0 0.0701f
C33007 VPWR.n6153 0 0.0485f
C33008 VPWR.n6154 0 0.018f
C33009 VPWR.n6155 0 0.0199f
C33010 VPWR.n6156 0 0.0118f
C33011 VPWR.n6157 0 0.0971f
C33012 VPWR.n6158 0 0.073f
C33013 VPWR.n6159 0 0.018f
C33014 VPWR.n6160 0 0.0199f
C33015 VPWR.n6161 0 0.0199f
C33016 VPWR.t330 0 0.068f
C33017 VPWR.n6162 0 0.0761f
C33018 VPWR.n6163 0 0.0402f
C33019 VPWR.n6164 0 0.0659f
C33020 VPWR.n6165 0 0.0634f
C33021 VPWR.n6166 0 0.0118f
C33022 VPWR.n6167 0 0.0107f
C33023 VPWR.n6168 0 0.062f
C33024 VPWR.n6169 0 0.0636f
C33025 VPWR.n6170 0 0.0173f
C33026 VPWR.t107 0 0.0876f
C33027 VPWR.n6171 0 0.183f
C33028 VPWR.n6172 0 0.0199f
C33029 VPWR.n6173 0 0.0522f
C33030 VPWR.n6174 0 0.0199f
C33031 VPWR.n6175 0 0.0199f
C33032 VPWR.n6176 0 0.0199f
C33033 VPWR.n6177 0 0.0118f
C33034 VPWR.n6178 0 0.00497f
C33035 VPWR.n6179 0 0.00162f
C33036 VPWR.n6180 0 0.0027f
C33037 VPWR.n6181 0 0.0013f
C33038 VPWR.n6182 0 0.0013f
C33039 VPWR.n6183 0 0.0027f
C33040 VPWR.n6184 0 0.00162f
C33041 VPWR.n6185 0 0.00205f
C33042 VPWR.n6186 0 0.00443f
C33043 VPWR.n6187 0 0.00302f
C33044 VPWR.n6188 0 0.00281f
C33045 VPWR.n6189 0 8.64e-19
C33046 VPWR.n6190 0 0.00238f
C33047 VPWR.n6191 0 0.00212f
C33048 VPWR.n6192 0 0.0672f
C33049 VPWR.n6193 0 0.321f
C33050 VPWR.n6194 0 0.307f
C33051 VPWR.n6195 0 0.0716f
C33052 VPWR.n6196 0 0.0725f
C33053 VPWR.t130 0 0.0718f
C33054 VPWR.n6197 0 0.208f
C33055 VPWR.n6198 0 0.0491f
C33056 VPWR.n6199 0 0.00994f
C33057 VPWR.n6200 0 0.0208f
C33058 VPWR.n6201 0 0.0117f
C33059 VPWR.n6202 0 0.13f
C33060 VPWR.n6203 0 0.194f
C33061 VPWR.n6204 0 0.0854f
C33062 VPWR.n6205 0 0.00441f
C33063 VPWR.n6206 0 0.0118f
C33064 VPWR.n6207 0 0.0199f
C33065 VPWR.n6208 0 0.0199f
C33066 VPWR.n6209 0 0.00455f
C33067 VPWR.n6210 0 0.0199f
C33068 VPWR.n6211 0 0.018f
C33069 VPWR.n6212 0 0.00593f
C33070 VPWR.n6213 0 0.502f
C33071 VPWR.n6214 0 0.0267f
C33072 VPWR.n6215 0 0.0125f
C33073 VPWR.n6216 0 0.00784f
C33074 VPWR.n6217 0 0.0199f
C33075 VPWR.n6218 0 0.018f
C33076 VPWR.n6219 0 0.0263f
C33077 VPWR.n6220 0 0.0651f
C33078 VPWR.n6221 0 0.0118f
C33079 VPWR.n6222 0 0.0199f
C33080 VPWR.n6223 0 0.0199f
C33081 VPWR.n6224 0 0.0429f
C33082 VPWR.n6225 0 0.0394f
C33083 VPWR.n6226 0 0.0373f
C33084 VPWR.n6227 0 0.00994f
C33085 VPWR.n6228 0 0.0107f
C33086 VPWR.n6229 0 0.0387f
C33087 VPWR.n6230 0 0.0619f
C33088 VPWR.n6231 0 0.0118f
C33089 VPWR.n6232 0 0.0535f
C33090 VPWR.n6233 0 0.0199f
C33091 VPWR.n6234 0 0.051f
C33092 VPWR.n6235 0 0.0199f
C33093 VPWR.t61 0 0.068f
C33094 VPWR.n6236 0 0.0785f
C33095 VPWR.n6237 0 0.0476f
C33096 VPWR.n6238 0 0.0199f
C33097 VPWR.n6239 0 0.0199f
C33098 VPWR.n6240 0 0.018f
C33099 VPWR.n6241 0 0.00994f
C33100 VPWR.n6242 0 0.0225f
C33101 VPWR.n6243 0 0.15f
C33102 VPWR.n6244 0 0.0118f
C33103 VPWR.n6245 0 0.0987f
C33104 VPWR.n6246 0 0.0199f
C33105 VPWR.n6247 0 0.0973f
C33106 VPWR.n6248 0 0.0199f
C33107 VPWR.n6249 0 0.0199f
C33108 VPWR.n6250 0 0.0518f
C33109 VPWR.n6251 0 0.0531f
C33110 VPWR.n6252 0 0.00994f
C33111 VPWR.n6253 0 0.096f
C33112 VPWR.n6254 0 0.105f
C33113 VPWR.n6255 0 0.0545f
C33114 VPWR.n6256 0 0.182f
C33115 VPWR.n6257 0 0.018f
C33116 VPWR.n6258 0 0.00778f
C33117 VPWR.n6259 0 0.00616f
C33118 VPWR.n6260 0 0.00891f
C33119 VPWR.n6261 0 0.00119f
C33120 VPWR.n6262 0 0.00259f
C33121 VPWR.n6263 0 0.00184f
C33122 VPWR.n6264 0 0.00194f
C33123 VPWR.n6265 0 0.00248f
C33124 VPWR.n6266 0 0.00248f
C33125 VPWR.n6267 0 0.00227f
C33126 VPWR.n6268 0 8.64e-19
C33127 VPWR.n6269 0 0.00259f
C33128 VPWR.n6270 0 5.4e-19
C33129 VPWR.n6271 0 0.00248f
C33130 VPWR.n6272 0 0.00302f
C33131 VPWR.n6273 0 0.00119f
C33132 VPWR.n6274 0 0.00184f
C33133 VPWR.n6275 0 0.00248f
C33134 VPWR.n6276 0 0.0014f
C33135 VPWR.n6277 0 0.00173f
C33136 VPWR.n6278 0 8.64e-19
C33137 VPWR.n6279 0 0.0014f
C33138 VPWR.n6280 0 0.00248f
C33139 VPWR.n6281 0 0.00357f
C33140 VPWR.n6282 0 0.00216f
C33141 VPWR.n6283 0 0.00162f
C33142 VPWR.n6284 0 0.00259f
C33143 VPWR.n6285 0 0.0014f
C33144 VPWR.n6286 0 0.0013f
C33145 VPWR.n6287 0 0.00172f
C33146 VPWR.n6288 0 0.00702f
C33147 VPWR.n6289 0 0.0107f
C33148 VPWR.n6290 0 0.125f
C33149 VPWR.n6291 0 0.11f
C33150 VPWR.n6292 0 0.0118f
C33151 VPWR.n6293 0 0.0199f
C33152 VPWR.n6294 0 0.0199f
C33153 VPWR.n6295 0 0.0199f
C33154 VPWR.n6296 0 0.0199f
C33155 VPWR.n6297 0 0.0191f
C33156 VPWR.n6298 0 0.0692f
C33157 VPWR.n6299 0 0.0423f
C33158 VPWR.n6300 0 0.0513f
C33159 VPWR.n6301 0 0.0199f
C33160 VPWR.n6302 0 0.0199f
C33161 VPWR.n6303 0 0.018f
C33162 VPWR.n6304 0 0.103f
C33163 VPWR.n6305 0 0.503f
C33164 VPWR.n6306 0 0.00467f
C33165 sample 0 0.104f
C33166 _286_/Y 0 0.221f
C33167 output30/a_27_7# 0 0.32f
C33168 valid 0 0.113f
C33169 _298_/X 0 0.191f
C33170 output41/a_27_7# 0 0.32f
C33171 VGND 0 0.325p
C33172 ctln[0] 0 0.227f
C33173 VPWR 0 0.671p
C33174 _269_/Y 0 0.199f
C33175 output6/a_27_7# 0 0.32f
C33176 _201_/a_27_7# 0 0.32f
C33177 _347_/D 0 0.174f
C33178 _347_/a_651_373# 0 0.00469f
C33179 _347_/a_448_7# 0 0.0139f
C33180 _347_/a_1108_7# 0 0.139f
C33181 _347_/a_1283_n19# 0 0.299f
C33182 _347_/a_543_7# 0 0.158f
C33183 _347_/a_761_249# 0 0.121f
C33184 _347_/a_193_7# 0 0.274f
C33185 _347_/a_27_7# 0 0.496f
C33186 _278_/a_68_257# 0 0.154f
C33187 _295_/a_512_7# 0 0.0326f
C33188 _295_/a_79_n19# 0 0.158f
C33189 clkc 0 0.221f
C33190 _297_/Y 0 0.183f
C33191 output5/a_27_7# 0 0.208f
C33192 trimb[4] 0 0.17f
C33193 output40/a_27_7# 0 0.32f
C33194 _336_/D 0 0.172f
C33195 _284_/A 0 0.659f
C33196 _202_/a_250_257# 0 0.0278f
C33197 _202_/a_93_n19# 0 0.151f
C33198 _279_/A 0 0.424f
C33199 _150_/a_27_7# 0 0.499f
C33200 _296_/a_213_83# 0 0.0371f
C33201 _296_/a_109_7# 0 0.0115f
C33202 _147_/Y 0 0.652f
C33203 _203_/a_209_257# 0 0.00621f
C33204 _203_/a_80_n19# 0 0.211f
C33205 _328_/D 0 0.185f
C33206 _220_/a_250_257# 0 0.0278f
C33207 _220_/a_93_n19# 0 0.151f
C33208 _297_/a_27_257# 0 0.0647f
C33209 _190_/A 0 0.718f
C33210 _333_/Q 0 0.726f
C33211 _332_/Q 0 0.73f
C33212 _204_/a_277_7# 0 0.00976f
C33213 _204_/a_27_7# 0 0.0193f
C33214 _204_/a_27_257# 0 0.0672f
C33215 _153_/B 0 0.335f
C33216 _327_/D 0 0.182f
C33217 _328_/Q 0 0.509f
C33218 _221_/a_250_257# 0 0.0278f
C33219 _221_/a_93_n19# 0 0.151f
C33220 _298_/A 0 0.779f
C33221 _298_/a_27_7# 0 0.177f
C33222 _204_/Y 0 0.245f
C33223 _335_/Q 0 0.254f
C33224 _205_/a_297_7# 0 0.0348f
C33225 _205_/a_79_n19# 0 0.158f
C33226 _154_/A 0 0.176f
C33227 _153_/A 0 0.353f
C33228 _153_/a_215_257# 0 0.414f
C33229 _153_/a_109_53# 0 0.148f
C33230 _217_/X 0 0.57f
C33231 _212_/X 0 0.617f
C33232 _327_/Q 0 0.535f
C33233 _222_/a_250_257# 0 0.0278f
C33234 _222_/a_93_n19# 0 0.151f
C33235 _299_/a_215_7# 0 0.0357f
C33236 _299_/a_78_159# 0 0.154f
C33237 _346_/D 0 0.139f
C33238 _170_/a_489_373# 0 0.0254f
C33239 _170_/a_226_7# 0 0.162f
C33240 _170_/a_76_159# 0 0.141f
C33241 _207_/C 0 0.31f
C33242 _206_/A 0 0.64f
C33243 _254_/B 0 0.597f
C33244 _154_/a_27_7# 0 0.208f
C33245 _325_/D 0 0.165f
C33246 _223_/a_250_257# 0 0.0278f
C33247 _223_/a_93_n19# 0 0.151f
C33248 _172_/B 0 0.157f
C33249 _171_/a_215_7# 0 0.0357f
C33250 _171_/a_78_159# 0 0.154f
C33251 _319_/D 0 0.18f
C33252 _207_/a_27_7# 0 0.177f
C33253 _324_/D 0 0.172f
C33254 _217_/A 0 0.492f
C33255 _304_/X 0 0.728f
C33256 _224_/a_250_257# 0 0.0278f
C33257 _224_/a_93_n19# 0 0.151f
C33258 _241_/a_113_257# 0 0.034f
C33259 _310_/Q 0 0.292f
C33260 _310_/D 0 0.174f
C33261 _310_/a_651_373# 0 0.00469f
C33262 _310_/a_448_7# 0 0.0139f
C33263 _310_/a_1108_7# 0 0.139f
C33264 _310_/a_1283_n19# 0 0.299f
C33265 _310_/a_543_7# 0 0.158f
C33266 _310_/a_761_249# 0 0.121f
C33267 _310_/a_193_7# 0 0.274f
C33268 _310_/a_27_7# 0 0.496f
C33269 _207_/X 0 0.133f
C33270 _208_/a_215_7# 0 0.0357f
C33271 _208_/a_78_159# 0 0.154f
C33272 _225_/B 0 0.351f
C33273 _336_/Q 0 0.414f
C33274 _225_/a_59_35# 0 0.177f
C33275 _156_/a_39_257# 0 0.229f
C33276 _311_/Q 0 0.267f
C33277 _311_/D 0 0.187f
C33278 _311_/a_651_373# 0 0.00469f
C33279 _311_/a_448_7# 0 0.0139f
C33280 _311_/a_1108_7# 0 0.139f
C33281 _311_/a_1283_n19# 0 0.299f
C33282 _311_/a_543_7# 0 0.158f
C33283 _311_/a_761_249# 0 0.121f
C33284 _311_/a_193_7# 0 0.274f
C33285 _311_/a_27_7# 0 0.496f
C33286 _172_/Y 0 0.123f
C33287 _345_/D 0 0.137f
C33288 _345_/Q 0 0.502f
C33289 _173_/a_489_373# 0 0.0254f
C33290 _173_/a_226_7# 0 0.162f
C33291 _173_/a_76_159# 0 0.141f
C33292 _318_/D 0 0.163f
C33293 _242_/B 0 0.141f
C33294 _190_/a_27_7# 0 0.32f
C33295 _209_/a_109_257# 0 0.00274f
C33296 _209_/a_27_257# 0 0.19f
C33297 _157_/a_27_7# 0 0.32f
C33298 _226_/X 0 0.161f
C33299 _150_/C 0 0.887f
C33300 _225_/X 0 0.131f
C33301 _147_/A 0 0.618f
C33302 _226_/a_297_7# 0 0.0348f
C33303 _226_/a_79_n19# 0 0.158f
C33304 _344_/D 0 0.13f
C33305 _344_/Q 0 0.459f
C33306 _174_/a_109_257# 0 0.00274f
C33307 _174_/a_27_257# 0 0.19f
C33308 _312_/Q 0 0.304f
C33309 _312_/D 0 0.179f
C33310 _312_/a_651_373# 0 0.00469f
C33311 _312_/a_448_7# 0 0.0139f
C33312 _312_/a_1108_7# 0 0.139f
C33313 _312_/a_1283_n19# 0 0.299f
C33314 _312_/a_543_7# 0 0.158f
C33315 _312_/a_761_249# 0 0.121f
C33316 _312_/a_193_7# 0 0.274f
C33317 _312_/a_27_7# 0 0.496f
C33318 _326_/Q 0 0.638f
C33319 _243_/a_113_257# 0 0.034f
C33320 _192_/B 0 0.443f
C33321 _323_/Q 0 0.361f
C33322 _191_/B 0 0.426f
C33323 _260_/a_27_257# 0 0.0647f
C33324 _313_/a_651_373# 0 0.00469f
C33325 _313_/a_448_7# 0 0.0139f
C33326 _313_/a_1108_7# 0 0.139f
C33327 _313_/a_1283_n19# 0 0.299f
C33328 _313_/a_543_7# 0 0.158f
C33329 _313_/a_761_249# 0 0.121f
C33330 _313_/a_193_7# 0 0.274f
C33331 _313_/a_27_7# 0 0.496f
C33332 _317_/D 0 0.19f
C33333 _244_/B 0 0.168f
C33334 _175_/Y 0 0.274f
C33335 _194_/A 0 0.338f
C33336 _305_/X 0 0.122f
C33337 _192_/a_68_257# 0 0.154f
C33338 _261_/A 0 0.141f
C33339 _267_/A 0 0.614f
C33340 _330_/a_651_373# 0 0.00469f
C33341 _330_/a_448_7# 0 0.0139f
C33342 _330_/a_1108_7# 0 0.139f
C33343 _330_/a_1283_n19# 0 0.299f
C33344 _330_/a_543_7# 0 0.158f
C33345 _330_/a_761_249# 0 0.121f
C33346 _330_/a_193_7# 0 0.274f
C33347 _330_/a_27_7# 0 0.496f
C33348 _228_/A 0 0.387f
C33349 _160_/A 0 0.244f
C33350 _162_/A 0 0.504f
C33351 _298_/C 0 0.62f
C33352 _343_/Q 0 0.37f
C33353 _176_/a_27_7# 0 0.208f
C33354 _314_/Q 0 0.247f
C33355 _314_/D 0 0.195f
C33356 _297_/B 0 1.59f
C33357 _314_/a_651_373# 0 0.00469f
C33358 _314_/a_448_7# 0 0.0139f
C33359 _314_/a_1108_7# 0 0.139f
C33360 _314_/a_1283_n19# 0 0.299f
C33361 _314_/a_543_7# 0 0.158f
C33362 _314_/a_761_249# 0 0.121f
C33363 _314_/a_193_7# 0 0.274f
C33364 _314_/a_27_7# 0 0.496f
C33365 _246_/B 0 0.135f
C33366 _245_/a_113_257# 0 0.034f
C33367 _262_/a_113_257# 0 0.034f
C33368 _331_/a_651_373# 0 0.00469f
C33369 _331_/a_448_7# 0 0.0139f
C33370 _331_/a_1108_7# 0 0.139f
C33371 _331_/a_1283_n19# 0 0.299f
C33372 _331_/a_543_7# 0 0.158f
C33373 _331_/a_761_249# 0 0.121f
C33374 _331_/a_193_7# 0 0.274f
C33375 _331_/a_27_7# 0 0.496f
C33376 _248_/A 0 0.813f
C33377 _229_/a_489_373# 0 0.0254f
C33378 _229_/a_226_7# 0 0.162f
C33379 _229_/a_76_159# 0 0.141f
C33380 _177_/A 0 0.441f
C33381 _177_/a_27_7# 0 0.32f
C33382 _315_/D 0 0.242f
C33383 _315_/a_651_373# 0 0.00469f
C33384 _315_/a_448_7# 0 0.0139f
C33385 _315_/a_1108_7# 0 0.139f
C33386 _315_/a_1283_n19# 0 0.299f
C33387 _315_/a_543_7# 0 0.158f
C33388 _315_/a_761_249# 0 0.121f
C33389 _315_/a_193_7# 0 0.274f
C33390 _315_/a_27_7# 0 0.496f
C33391 _263_/B 0 0.127f
C33392 _194_/a_27_7# 0 0.208f
C33393 _332_/D 0 0.18f
C33394 _340_/CLK 0 1.76f
C33395 _332_/a_651_373# 0 0.00469f
C33396 _332_/a_448_7# 0 0.0139f
C33397 _332_/a_1108_7# 0 0.135f
C33398 _332_/a_1283_n19# 0 0.564f
C33399 _332_/a_543_7# 0 0.158f
C33400 _332_/a_761_249# 0 0.121f
C33401 _332_/a_193_7# 0 0.273f
C33402 _332_/a_27_7# 0 0.496f
C33403 _281_/A 0 0.441f
C33404 _280_/a_68_257# 0 0.154f
C33405 _178_/a_27_7# 0 0.499f
C33406 _248_/B 0 0.151f
C33407 _232_/A 0 0.554f
C33408 _247_/a_113_257# 0 0.034f
C33409 _316_/D 0 0.0256f
C33410 _331_/CLK 0 2.04f
C33411 _316_/a_651_373# 0 0.00469f
C33412 _316_/a_448_7# 0 0.0139f
C33413 _316_/a_1108_7# 0 0.139f
C33414 _316_/a_1283_n19# 0 0.299f
C33415 _316_/a_543_7# 0 0.158f
C33416 _316_/a_761_249# 0 0.121f
C33417 _316_/a_193_7# 0 0.274f
C33418 _316_/a_27_7# 0 0.496f
C33419 _265_/B 0 0.148f
C33420 _264_/a_113_257# 0 0.034f
C33421 _333_/D 0 0.175f
C33422 _333_/a_651_373# 0 0.00469f
C33423 _333_/a_448_7# 0 0.0139f
C33424 _333_/a_1108_7# 0 0.135f
C33425 _333_/a_1283_n19# 0 0.564f
C33426 _333_/a_543_7# 0 0.158f
C33427 _333_/a_761_249# 0 0.121f
C33428 _333_/a_193_7# 0 0.273f
C33429 _333_/a_27_7# 0 0.496f
C33430 _340_/D 0 0.221f
C33431 _193_/Y 0 0.517f
C33432 _306_/S 0 1.15f
C33433 _340_/Q 0 0.405f
C33434 _194_/X 0 0.593f
C33435 _195_/a_109_257# 0 0.00274f
C33436 _195_/a_27_257# 0 0.19f
C33437 _179_/a_27_7# 0 0.32f
C33438 _317_/a_651_373# 0 0.00469f
C33439 _317_/a_448_7# 0 0.0139f
C33440 _317_/a_1108_7# 0 0.139f
C33441 _317_/a_1283_n19# 0 0.299f
C33442 _317_/a_543_7# 0 0.158f
C33443 _317_/a_761_249# 0 0.121f
C33444 _317_/a_193_7# 0 0.274f
C33445 _317_/a_27_7# 0 0.496f
C33446 _334_/Q 0 0.415f
C33447 _334_/D 0 0.198f
C33448 _343_/CLK 0 2.18f
C33449 _334_/a_651_373# 0 0.00469f
C33450 _334_/a_448_7# 0 0.0139f
C33451 _334_/a_1108_7# 0 0.139f
C33452 _334_/a_1283_n19# 0 0.299f
C33453 _334_/a_543_7# 0 0.158f
C33454 _334_/a_761_249# 0 0.121f
C33455 _334_/a_193_7# 0 0.274f
C33456 _334_/a_27_7# 0 0.496f
C33457 _282_/a_39_257# 0 0.229f
C33458 _318_/a_651_373# 0 0.00469f
C33459 _318_/a_448_7# 0 0.0139f
C33460 _318_/a_1108_7# 0 0.139f
C33461 _318_/a_1283_n19# 0 0.299f
C33462 _318_/a_543_7# 0 0.158f
C33463 _318_/a_761_249# 0 0.121f
C33464 _318_/a_193_7# 0 0.274f
C33465 _318_/a_27_7# 0 0.496f
C33466 _309_/Q 0 0.268f
C33467 _266_/a_113_257# 0 0.034f
C33468 _260_/A 0 0.442f
C33469 _197_/a_27_7# 0 0.32f
C33470 _335_/D 0 0.237f
C33471 _335_/a_651_373# 0 0.00469f
C33472 _335_/a_448_7# 0 0.0139f
C33473 _335_/a_1108_7# 0 0.139f
C33474 _335_/a_1283_n19# 0 0.299f
C33475 _335_/a_543_7# 0 0.158f
C33476 _335_/a_761_249# 0 0.121f
C33477 _335_/a_193_7# 0 0.274f
C33478 _335_/a_27_7# 0 0.496f
C33479 _283_/A 0 0.468f
C33480 clkbuf_1_0_0_clk/a_75_172# 0 0.21f
C33481 _319_/a_651_373# 0 0.00469f
C33482 _319_/a_448_7# 0 0.0139f
C33483 _319_/a_1108_7# 0 0.139f
C33484 _319_/a_1283_n19# 0 0.299f
C33485 _319_/a_543_7# 0 0.158f
C33486 _319_/a_761_249# 0 0.121f
C33487 _319_/a_193_7# 0 0.274f
C33488 _319_/a_27_7# 0 0.496f
C33489 _336_/a_651_373# 0 0.00469f
C33490 _336_/a_448_7# 0 0.0139f
C33491 _336_/a_1108_7# 0 0.139f
C33492 _336_/a_1283_n19# 0 0.299f
C33493 _336_/a_543_7# 0 0.158f
C33494 _336_/a_761_249# 0 0.121f
C33495 _336_/a_193_7# 0 0.274f
C33496 _336_/a_27_7# 0 0.496f
C33497 _309_/D 0 0.183f
C33498 _267_/B 0 0.136f
C33499 _198_/a_250_257# 0 0.0278f
C33500 _198_/a_93_n19# 0 0.151f
C33501 _284_/a_39_257# 0 0.229f
C33502 _199_/a_250_257# 0 0.0278f
C33503 _199_/a_93_n19# 0 0.151f
C33504 _337_/Q 0 0.491f
C33505 _337_/D 0 0.169f
C33506 _337_/a_651_373# 0 0.00469f
C33507 _337_/a_448_7# 0 0.0139f
C33508 _337_/a_1108_7# 0 0.139f
C33509 _337_/a_1283_n19# 0 0.299f
C33510 _337_/a_543_7# 0 0.158f
C33511 _337_/a_761_249# 0 0.121f
C33512 _337_/a_193_7# 0 0.274f
C33513 _337_/a_27_7# 0 0.496f
C33514 _268_/a_39_257# 0 0.229f
C33515 clkbuf_1_1_0_clk/a_75_172# 0 0.21f
C33516 _285_/Y 0 0.179f
C33517 _269_/A 0 0.596f
C33518 _338_/Q 0 0.468f
C33519 _346_/SET_B 0 5.25f
C33520 _338_/D 0 0.19f
C33521 _338_/a_651_373# 0 0.00469f
C33522 _338_/a_448_7# 0 0.0139f
C33523 _338_/a_1108_7# 0 0.139f
C33524 _338_/a_1283_n19# 0 0.299f
C33525 _338_/a_543_7# 0 0.158f
C33526 _338_/a_761_249# 0 0.121f
C33527 _338_/a_193_7# 0 0.274f
C33528 _338_/a_27_7# 0 0.496f
C33529 _339_/Q 0 0.479f
C33530 _339_/D 0 0.194f
C33531 _339_/a_651_373# 0 0.00469f
C33532 _339_/a_448_7# 0 0.0139f
C33533 _339_/a_1108_7# 0 0.139f
C33534 _339_/a_1283_n19# 0 0.299f
C33535 _339_/a_543_7# 0 0.158f
C33536 _339_/a_761_249# 0 0.121f
C33537 _339_/a_193_7# 0 0.274f
C33538 _339_/a_27_7# 0 0.496f
C33539 _209_/X 0 0.121f
C33540 _210_/a_27_7# 0 0.0465f
C33541 _287_/a_39_257# 0 0.229f
C33542 _149_/A 0 0.314f
C33543 _197_/X 0 0.651f
C33544 _211_/a_109_257# 0 0.00274f
C33545 _211_/a_27_257# 0 0.19f
C33546 rstn 0 1.64f
C33547 input4/a_27_7# 0 0.208f
C33548 _288_/Y 0 0.152f
C33549 _144_/A 0 0.152f
C33550 _143_/a_27_7# 0 0.177f
C33551 _212_/a_27_7# 0 0.208f
C33552 _289_/a_39_257# 0 0.229f
C33553 _227_/A 0 0.753f
C33554 en 0 0.225f
C33555 input3/a_27_7# 0 0.32f
C33556 _160_/a_27_7# 0 0.32f
C33557 _144_/a_27_7# 0 0.208f
C33558 comp 0 0.778f
C33559 input2/a_27_7# 0 0.208f
C33560 _161_/Y 0 0.39f
C33561 _242_/A 0 0.691f
C33562 _230_/a_27_7# 0 0.32f
C33563 _304_/S 0 0.561f
C33564 _331_/D 0 0.186f
C33565 _214_/a_109_257# 0 0.00274f
C33566 _214_/a_27_257# 0 0.19f
C33567 input1/X 0 0.179f
C33568 cal 0 3.95f
C33569 input1/a_75_172# 0 0.21f
C33570 _300_/Y 0 0.126f
C33571 _160_/X 0 0.561f
C33572 _347_/Q 0 0.542f
C33573 _299_/X 0 0.405f
C33574 _300_/a_735_7# 0 0.00532f
C33575 _300_/a_383_7# 0 0.00406f
C33576 _300_/a_301_257# 0 0.0376f
C33577 _300_/a_27_257# 0 0.0292f
C33578 _162_/a_27_7# 0 0.32f
C33579 _162_/X 0 0.621f
C33580 _231_/a_512_7# 0 0.0326f
C33581 _231_/a_79_n19# 0 0.158f
C33582 _215_/A 0 0.361f
C33583 _146_/C 0 0.282f
C33584 _146_/a_29_271# 0 0.271f
C33585 _301_/a_240_7# 0 0.0138f
C33586 _301_/a_149_7# 0 0.00821f
C33587 _301_/a_51_257# 0 0.207f
C33588 _158_/Y 0 0.235f
C33589 _163_/a_215_7# 0 0.0357f
C33590 _163_/a_78_159# 0 0.154f
C33591 _232_/X 0 0.948f
C33592 _232_/a_27_7# 0 0.32f
C33593 _180_/a_29_13# 0 0.18f
C33594 clkbuf_2_1_0_clk/A 0 0.332f
C33595 clkbuf_2_0_0_clk/a_75_172# 0 0.21f
C33596 ctlp[5] 0 0.385f
C33597 output19/a_27_7# 0 0.32f
C33598 _216_/a_27_7# 0 0.32f
C33599 _164_/Y 0 0.219f
C33600 _164_/A 0 0.317f
C33601 _303_/A 0 0.262f
C33602 _301_/X 0 0.135f
C33603 _302_/a_227_7# 0 0.0309f
C33604 _302_/a_77_159# 0 0.147f
C33605 _331_/Q 0 0.613f
C33606 _322_/Q 0 0.484f
C33607 _233_/a_113_257# 0 0.034f
C33608 _250_/X 0 0.143f
C33609 _216_/A 0 0.614f
C33610 _250_/a_215_7# 0 0.0357f
C33611 _250_/a_78_159# 0 0.154f
C33612 _181_/a_27_7# 0 0.32f
C33613 result[7] 0 0.919f
C33614 output29/a_27_7# 0 0.32f
C33615 ctlp[4] 0 0.386f
C33616 output18/a_27_7# 0 0.32f
C33617 _298_/B 0 0.325f
C33618 _341_/Q 0 0.665f
C33619 _217_/a_27_7# 0 0.32f
C33620 _165_/a_215_7# 0 0.0357f
C33621 _165_/a_78_159# 0 0.154f
C33622 clkbuf_2_1_0_clk/a_75_172# 0 0.21f
C33623 _322_/D 0 0.19f
C33624 _234_/B 0 0.13f
C33625 _182_/X 0 0.163f
C33626 _181_/X 0 0.871f
C33627 _196_/A 0 0.747f
C33628 _286_/B 0 1.18f
C33629 _182_/a_215_7# 0 0.0101f
C33630 _182_/a_79_n19# 0 0.225f
C33631 _251_/X 0 0.119f
C33632 _251_/a_215_7# 0 0.0101f
C33633 _251_/a_79_n19# 0 0.225f
C33634 _320_/a_651_373# 0 0.00469f
C33635 _320_/a_448_7# 0 0.0139f
C33636 _320_/a_1108_7# 0 0.139f
C33637 _320_/a_1283_n19# 0 0.299f
C33638 _320_/a_543_7# 0 0.158f
C33639 _320_/a_761_249# 0 0.121f
C33640 _320_/a_193_7# 0 0.274f
C33641 _320_/a_27_7# 0 0.496f
C33642 result[6] 0 0.244f
C33643 output28/a_27_7# 0 0.32f
C33644 ctlp[3] 0 0.353f
C33645 output17/a_27_7# 0 0.32f
C33646 trimb[3] 0 0.615f
C33647 output39/a_27_7# 0 0.32f
C33648 _149_/a_27_7# 0 0.32f
C33649 _330_/D 0 0.204f
C33650 _218_/a_250_257# 0 0.0278f
C33651 _218_/a_93_n19# 0 0.151f
C33652 _166_/Y 0 0.233f
C33653 _346_/Q 0 0.485f
C33654 _216_/X 0 0.608f
C33655 _304_/a_257_159# 0 0.216f
C33656 _304_/a_79_n19# 0 0.227f
C33657 _330_/Q 0 0.798f
C33658 _321_/Q 0 0.503f
C33659 _235_/a_113_257# 0 0.034f
C33660 _324_/Q 0 1.06f
C33661 _157_/A 0 0.653f
C33662 _183_/a_471_7# 0 0.0538f
C33663 _183_/a_27_7# 0 0.0485f
C33664 _183_/a_553_257# 0 0.00146f
C33665 _297_/A 0 0.347f
C33666 _252_/a_27_7# 0 0.0311f
C33667 _321_/a_651_373# 0 0.00469f
C33668 _321_/a_448_7# 0 0.0139f
C33669 _321_/a_1108_7# 0 0.139f
C33670 _321_/a_1283_n19# 0 0.299f
C33671 _321_/a_543_7# 0 0.158f
C33672 _321_/a_761_249# 0 0.121f
C33673 _321_/a_193_7# 0 0.274f
C33674 _321_/a_27_7# 0 0.496f
C33675 clkbuf_2_3_0_clk/A 0 0.302f
C33676 clkbuf_2_2_0_clk/a_75_172# 0 0.21f
C33677 clkbuf_0_clk/X 0 0.385f
C33678 clk 0 3.57f
C33679 clkbuf_0_clk/a_110_7# 0 1.73f
C33680 result[5] 0 0.105f
C33681 output27/a_27_7# 0 0.32f
C33682 trimb[2] 0 0.156f
C33683 output38/a_27_7# 0 0.32f
C33684 ctlp[2] 0 0.337f
C33685 output16/a_27_7# 0 0.32f
C33686 _329_/D 0 0.182f
C33687 _219_/a_250_257# 0 0.0278f
C33688 _219_/a_93_n19# 0 0.151f
C33689 _305_/a_505_n19# 0 0.247f
C33690 _305_/a_76_159# 0 0.139f
C33691 _167_/a_109_257# 0 0.00274f
C33692 _167_/a_27_257# 0 0.19f
C33693 _321_/D 0 0.195f
C33694 _236_/B 0 0.155f
C33695 _188_/S 0 0.602f
C33696 _184_/a_505_n19# 0 0.247f
C33697 _184_/a_76_159# 0 0.139f
C33698 _322_/a_651_373# 0 0.00469f
C33699 _322_/a_448_7# 0 0.0139f
C33700 _322_/a_1108_7# 0 0.139f
C33701 _322_/a_1283_n19# 0 0.299f
C33702 _322_/a_543_7# 0 0.158f
C33703 _322_/a_761_249# 0 0.121f
C33704 _322_/a_193_7# 0 0.274f
C33705 _322_/a_27_7# 0 0.496f
C33706 _325_/Q 0 0.467f
C33707 _270_/a_39_257# 0 0.229f
C33708 clkbuf_2_3_0_clk/a_75_172# 0 0.21f
C33709 trimb[1] 0 0.136f
C33710 output37/a_27_7# 0 0.32f
C33711 result[4] 0 0.11f
C33712 output26/a_27_7# 0 0.32f
C33713 ctlp[1] 0 0.36f
C33714 output15/a_27_7# 0 0.32f
C33715 _306_/a_505_n19# 0 0.247f
C33716 _306_/a_76_159# 0 0.139f
C33717 _165_/X 0 0.375f
C33718 _167_/X 0 0.311f
C33719 _168_/a_397_257# 0 0.0287f
C33720 _168_/a_109_7# 0 0.148f
C33721 _238_/B 0 0.15f
C33722 _329_/Q 0 0.459f
C33723 _320_/Q 0 0.521f
C33724 _237_/a_113_257# 0 0.034f
C33725 _254_/A 0 0.604f
C33726 _323_/D 0 0.197f
C33727 _323_/a_651_373# 0 0.00469f
C33728 _323_/a_448_7# 0 0.0139f
C33729 _323_/a_1108_7# 0 0.139f
C33730 _323_/a_1283_n19# 0 0.299f
C33731 _323_/a_543_7# 0 0.158f
C33732 _323_/a_761_249# 0 0.121f
C33733 _323_/a_193_7# 0 0.274f
C33734 _323_/a_27_7# 0 0.496f
C33735 _343_/D 0 0.166f
C33736 _185_/A 0 0.252f
C33737 _340_/a_651_373# 0 0.00469f
C33738 _340_/a_448_7# 0 0.0139f
C33739 _340_/a_1108_7# 0 0.139f
C33740 _340_/a_1283_n19# 0 0.299f
C33741 _340_/a_543_7# 0 0.158f
C33742 _340_/a_761_249# 0 0.121f
C33743 _340_/a_193_7# 0 0.274f
C33744 _340_/a_27_7# 0 0.496f
C33745 _271_/Y 0 0.188f
C33746 _271_/A 0 0.432f
C33747 result[3] 0 0.11f
C33748 _318_/Q 0 0.465f
C33749 output25/a_27_7# 0 0.32f
C33750 trimb[0] 0 0.146f
C33751 output36/a_27_7# 0 0.32f
C33752 ctlp[0] 0 0.394f
C33753 output14/a_27_7# 0 0.32f
C33754 _169_/Y 0 0.13f
C33755 _169_/B 0 0.124f
C33756 _145_/A 0 0.296f
C33757 _296_/Y 0 0.161f
C33758 _307_/a_505_n19# 0 0.247f
C33759 _307_/a_76_159# 0 0.139f
C33760 _320_/D 0 0.178f
C33761 _308_/X 0 0.145f
C33762 _172_/A 0 0.696f
C33763 _186_/a_297_7# 0 0.0348f
C33764 _186_/a_79_n19# 0 0.158f
C33765 _255_/X 0 0.117f
C33766 _342_/Q 0 0.725f
C33767 _255_/B 0 0.567f
C33768 _255_/a_30_13# 0 0.267f
C33769 _324_/a_651_373# 0 0.00469f
C33770 _324_/a_448_7# 0 0.0139f
C33771 _324_/a_1108_7# 0 0.137f
C33772 _324_/a_1283_n19# 0 0.389f
C33773 _324_/a_543_7# 0 0.158f
C33774 _324_/a_761_249# 0 0.121f
C33775 _324_/a_193_7# 0 0.273f
C33776 _324_/a_27_7# 0 0.496f
C33777 _341_/D 0 0.184f
C33778 _341_/a_651_373# 0 0.00469f
C33779 _341_/a_448_7# 0 0.0139f
C33780 _341_/a_1108_7# 0 0.135f
C33781 _341_/a_1283_n19# 0 0.564f
C33782 _341_/a_543_7# 0 0.158f
C33783 _341_/a_761_249# 0 0.121f
C33784 _341_/a_193_7# 0 0.273f
C33785 _341_/a_27_7# 0 0.496f
C33786 _272_/a_39_257# 0 0.229f
C33787 repeater43/X 0 5.28f
C33788 input4/X 0 0.576f
C33789 repeater43/a_27_7# 0 0.839f
C33790 trim[4] 0 0.17f
C33791 output35/a_27_7# 0 0.32f
C33792 ctln[7] 0 0.0154f
C33793 _283_/Y 0 1.46f
C33794 output13/a_27_7# 0 0.32f
C33795 result[2] 0 0.149f
C33796 _317_/Q 0 0.447f
C33797 output24/a_27_7# 0 0.32f
C33798 _308_/S 0 0.476f
C33799 _308_/a_505_n19# 0 0.247f
C33800 _308_/a_76_159# 0 0.139f
C33801 _240_/B 0 0.106f
C33802 _319_/Q 0 0.515f
C33803 _239_/a_113_257# 0 0.034f
C33804 _260_/B 0 0.304f
C33805 _256_/a_209_257# 0 0.00621f
C33806 _256_/a_80_n19# 0 0.211f
C33807 _187_/a_27_7# 0 0.208f
C33808 _325_/a_651_373# 0 0.00469f
C33809 _325_/a_448_7# 0 0.0139f
C33810 _325_/a_1108_7# 0 0.139f
C33811 _325_/a_1283_n19# 0 0.299f
C33812 _325_/a_543_7# 0 0.158f
C33813 _325_/a_761_249# 0 0.121f
C33814 _325_/a_193_7# 0 0.274f
C33815 _325_/a_27_7# 0 0.496f
C33816 _342_/D 0 0.194f
C33817 _342_/a_651_373# 0 0.00469f
C33818 _342_/a_448_7# 0 0.0139f
C33819 _342_/a_1108_7# 0 0.135f
C33820 _342_/a_1283_n19# 0 0.564f
C33821 _342_/a_543_7# 0 0.158f
C33822 _342_/a_761_249# 0 0.121f
C33823 _342_/a_193_7# 0 0.273f
C33824 _342_/a_27_7# 0 0.496f
C33825 _273_/Y 0 0.196f
C33826 _273_/A 0 0.521f
C33827 repeater42/a_27_7# 0 0.839f
C33828 _290_/Y 0 0.164f
C33829 ctln[6] 0 0.222f
C33830 _281_/Y 0 0.178f
C33831 output12/a_27_7# 0 0.32f
C33832 trim[3] 0 0.47f
C33833 _292_/A 0 0.447f
C33834 output34/a_27_7# 0 0.32f
C33835 result[1] 0 0.169f
C33836 _316_/Q 0 0.528f
C33837 output23/a_27_7# 0 0.32f
C33838 _309_/a_651_373# 0 0.00469f
C33839 _309_/a_448_7# 0 0.0139f
C33840 _309_/a_1108_7# 0 0.139f
C33841 _309_/a_1283_n19# 0 0.299f
C33842 _309_/a_543_7# 0 0.158f
C33843 _309_/a_761_249# 0 0.121f
C33844 _309_/a_193_7# 0 0.274f
C33845 _309_/a_27_7# 0 0.496f
C33846 _307_/X 0 0.156f
C33847 _188_/a_505_n19# 0 0.247f
C33848 _188_/a_76_159# 0 0.139f
C33849 _254_/Y 0 0.106f
C33850 _257_/a_448_7# 0 0.0324f
C33851 _257_/a_222_53# 0 0.159f
C33852 _257_/a_79_159# 0 0.148f
C33853 _326_/D 0 0.184f
C33854 _326_/a_651_373# 0 0.00469f
C33855 _326_/a_448_7# 0 0.0139f
C33856 _326_/a_1108_7# 0 0.139f
C33857 _326_/a_1283_n19# 0 0.299f
C33858 _326_/a_543_7# 0 0.158f
C33859 _326_/a_761_249# 0 0.121f
C33860 _326_/a_193_7# 0 0.274f
C33861 _326_/a_27_7# 0 0.496f
C33862 _343_/a_651_373# 0 0.00469f
C33863 _343_/a_448_7# 0 0.0139f
C33864 _343_/a_1108_7# 0 0.139f
C33865 _343_/a_1283_n19# 0 0.299f
C33866 _343_/a_543_7# 0 0.158f
C33867 _343_/a_761_249# 0 0.121f
C33868 _343_/a_193_7# 0 0.274f
C33869 _343_/a_27_7# 0 0.496f
C33870 _275_/A 0 0.415f
C33871 _274_/a_39_257# 0 0.229f
C33872 _291_/a_39_257# 0 0.229f
C33873 ctln[5] 0 0.204f
C33874 _279_/Y 0 0.235f
C33875 output11/a_27_7# 0 0.32f
C33876 ctln[3] 0 0.228f
C33877 _275_/Y 0 0.205f
C33878 output9/a_27_7# 0 0.32f
C33879 trim[2] 0 0.129f
C33880 _290_/A 0 0.445f
C33881 output33/a_27_7# 0 0.32f
C33882 result[0] 0 0.116f
C33883 _315_/Q 0 0.507f
C33884 output22/a_27_7# 0 0.32f
C33885 _306_/X 0 0.151f
C33886 _313_/Q 0 0.313f
C33887 _313_/D 0 0.184f
C33888 _258_/a_505_n19# 0 0.247f
C33889 _258_/a_76_159# 0 0.139f
C33890 _189_/a_27_7# 0 0.32f
C33891 _327_/a_651_373# 0 0.00469f
C33892 _327_/a_448_7# 0 0.0139f
C33893 _327_/a_1108_7# 0 0.139f
C33894 _327_/a_1283_n19# 0 0.299f
C33895 _327_/a_543_7# 0 0.158f
C33896 _327_/a_761_249# 0 0.121f
C33897 _327_/a_193_7# 0 0.274f
C33898 _327_/a_27_7# 0 0.496f
C33899 _344_/a_381_7# 0 0.0203f
C33900 _344_/a_1602_7# 0 0.126f
C33901 _344_/a_1032_373# 0 0.305f
C33902 _344_/a_1182_221# 0 0.128f
C33903 _344_/a_476_7# 0 0.286f
C33904 _344_/a_652_n19# 0 0.119f
C33905 _344_/a_193_7# 0 0.322f
C33906 _344_/a_27_7# 0 0.437f
C33907 _292_/Y 0 0.175f
C33908 trim[1] 0 0.126f
C33909 _288_/A 0 0.393f
C33910 output32/a_27_7# 0 0.32f
C33911 ctln[4] 0 0.178f
C33912 _277_/Y 0 0.203f
C33913 output10/a_27_7# 0 0.32f
C33914 ctln[2] 0 0.226f
C33915 output8/a_27_7# 0 0.32f
C33916 ctlp[7] 0 0.338f
C33917 output21/a_27_7# 0 0.32f
C33918 _258_/S 0 0.752f
C33919 _259_/a_113_257# 0 0.034f
C33920 _328_/a_651_373# 0 0.00469f
C33921 _328_/a_448_7# 0 0.0139f
C33922 _328_/a_1108_7# 0 0.139f
C33923 _328_/a_1283_n19# 0 0.299f
C33924 _328_/a_543_7# 0 0.158f
C33925 _328_/a_761_249# 0 0.121f
C33926 _328_/a_193_7# 0 0.274f
C33927 _328_/a_27_7# 0 0.496f
C33928 _345_/a_381_7# 0 0.0203f
C33929 _345_/a_1602_7# 0 0.126f
C33930 _345_/a_1032_373# 0 0.305f
C33931 _345_/a_1182_221# 0 0.128f
C33932 _345_/a_476_7# 0 0.286f
C33933 _345_/a_652_n19# 0 0.119f
C33934 _345_/a_193_7# 0 0.322f
C33935 _345_/a_27_7# 0 0.437f
C33936 _276_/a_68_257# 0 0.154f
C33937 _293_/a_39_257# 0 0.229f
C33938 trim[0] 0 0.151f
C33939 _285_/A 0 0.65f
C33940 output31/a_27_7# 0 0.32f
C33941 ctln[1] 0 0.199f
C33942 output7/a_27_7# 0 0.32f
C33943 ctlp[6] 0 0.379f
C33944 output20/a_27_7# 0 0.32f
C33945 _329_/a_651_373# 0 0.00469f
C33946 _329_/a_448_7# 0 0.0139f
C33947 _329_/a_1108_7# 0 0.139f
C33948 _329_/a_1283_n19# 0 0.299f
C33949 _329_/a_543_7# 0 0.158f
C33950 _329_/a_761_249# 0 0.121f
C33951 _329_/a_193_7# 0 0.274f
C33952 _329_/a_27_7# 0 0.496f
C33953 _200_/a_250_257# 0 0.0278f
C33954 _200_/a_93_n19# 0 0.151f
C33955 _277_/A 0 0.421f
C33956 _346_/a_381_7# 0 0.0203f
C33957 _346_/a_1602_7# 0 0.126f
C33958 _346_/a_1032_373# 0 0.305f
C33959 _346_/a_1182_221# 0 0.128f
C33960 _346_/a_476_7# 0 0.286f
C33961 _346_/a_652_n19# 0 0.119f
C33962 _346_/a_193_7# 0 0.322f
C33963 _346_/a_27_7# 0 0.437f
C33964 _294_/Y 0 0.151f
C33965 _294_/A 0 0.547f
.ends

