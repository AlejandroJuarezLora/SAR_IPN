magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 1970 542
<< pwell >>
rect 273 117 457 161
rect 1673 141 1857 163
rect 1390 117 1857 141
rect 1 -19 1857 117
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 109 91
rect 163 7 193 91
rect 351 7 381 135
rect 446 7 476 79
rect 556 7 586 79
rect 652 7 682 91
rect 766 7 796 91
rect 838 7 868 91
rect 1026 7 1056 91
rect 1098 7 1128 91
rect 1194 7 1224 91
rect 1266 7 1296 91
rect 1342 7 1372 91
rect 1466 7 1496 115
rect 1654 7 1684 91
rect 1749 7 1779 137
<< scpmoshvt >>
rect 79 323 109 451
rect 163 323 193 451
rect 351 289 381 457
rect 448 373 478 457
rect 532 373 562 457
rect 652 373 682 457
rect 758 373 788 457
rect 842 373 872 457
rect 926 373 956 457
rect 1002 373 1032 457
rect 1110 373 1140 457
rect 1182 373 1212 457
rect 1370 373 1400 457
rect 1466 289 1496 457
rect 1654 329 1684 457
rect 1749 257 1779 457
<< ndiff >>
rect 27 79 79 91
rect 27 45 35 79
rect 69 45 79 79
rect 27 7 79 45
rect 109 53 163 91
rect 109 19 119 53
rect 153 19 163 53
rect 109 7 163 19
rect 193 79 245 91
rect 193 45 203 79
rect 237 45 245 79
rect 193 7 245 45
rect 299 53 351 135
rect 299 19 307 53
rect 341 19 351 53
rect 299 7 351 19
rect 381 79 431 135
rect 1416 91 1466 115
rect 601 79 652 91
rect 381 71 446 79
rect 381 37 391 71
rect 425 37 446 71
rect 381 7 446 37
rect 476 53 556 79
rect 476 19 501 53
rect 535 19 556 53
rect 476 7 556 19
rect 586 7 652 79
rect 682 49 766 91
rect 682 15 722 49
rect 756 15 766 49
rect 682 7 766 15
rect 796 7 838 91
rect 868 69 920 91
rect 868 35 878 69
rect 912 35 920 69
rect 868 7 920 35
rect 974 53 1026 91
rect 974 19 982 53
rect 1016 19 1026 53
rect 974 7 1026 19
rect 1056 7 1098 91
rect 1128 55 1194 91
rect 1128 21 1144 55
rect 1178 21 1194 55
rect 1128 7 1194 21
rect 1224 7 1266 91
rect 1296 7 1342 91
rect 1372 73 1466 91
rect 1372 39 1402 73
rect 1436 39 1466 73
rect 1372 7 1466 39
rect 1496 80 1548 115
rect 1699 91 1749 137
rect 1496 46 1506 80
rect 1540 46 1548 80
rect 1496 7 1548 46
rect 1602 79 1654 91
rect 1602 45 1610 79
rect 1644 45 1654 79
rect 1602 7 1654 45
rect 1684 53 1749 91
rect 1684 19 1705 53
rect 1739 19 1749 53
rect 1684 7 1749 19
rect 1779 103 1831 137
rect 1779 69 1789 103
rect 1823 69 1831 103
rect 1779 7 1831 69
<< pdiff >>
rect 27 437 79 451
rect 27 403 35 437
rect 69 403 79 437
rect 27 369 79 403
rect 27 335 35 369
rect 69 335 79 369
rect 27 323 79 335
rect 109 421 163 451
rect 109 387 119 421
rect 153 387 163 421
rect 109 323 163 387
rect 193 437 245 451
rect 193 403 203 437
rect 237 403 245 437
rect 193 369 245 403
rect 193 335 203 369
rect 237 335 245 369
rect 193 323 245 335
rect 299 421 351 457
rect 299 387 307 421
rect 341 387 351 421
rect 299 289 351 387
rect 381 437 448 457
rect 381 403 391 437
rect 425 403 448 437
rect 381 373 448 403
rect 478 444 532 457
rect 478 410 488 444
rect 522 410 532 444
rect 478 373 532 410
rect 562 373 652 457
rect 682 445 758 457
rect 682 411 702 445
rect 736 411 758 445
rect 682 373 758 411
rect 788 419 842 457
rect 788 385 798 419
rect 832 385 842 419
rect 788 373 842 385
rect 872 445 926 457
rect 872 411 882 445
rect 916 411 926 445
rect 872 373 926 411
rect 956 373 1002 457
rect 1032 443 1110 457
rect 1032 409 1042 443
rect 1076 409 1110 443
rect 1032 373 1110 409
rect 1140 373 1182 457
rect 1212 445 1264 457
rect 1212 411 1222 445
rect 1256 411 1264 445
rect 1212 373 1264 411
rect 1318 419 1370 457
rect 1318 385 1326 419
rect 1360 385 1370 419
rect 1318 373 1370 385
rect 1400 419 1466 457
rect 1400 385 1422 419
rect 1456 385 1466 419
rect 1400 373 1466 385
rect 381 369 433 373
rect 381 335 391 369
rect 425 335 433 369
rect 381 289 433 335
rect 1415 289 1466 373
rect 1496 419 1548 457
rect 1496 385 1506 419
rect 1540 385 1548 419
rect 1496 351 1548 385
rect 1496 317 1506 351
rect 1540 317 1548 351
rect 1602 445 1654 457
rect 1602 411 1610 445
rect 1644 411 1654 445
rect 1602 377 1654 411
rect 1602 343 1610 377
rect 1644 343 1654 377
rect 1602 329 1654 343
rect 1684 445 1749 457
rect 1684 411 1705 445
rect 1739 411 1749 445
rect 1684 377 1749 411
rect 1684 343 1705 377
rect 1739 343 1749 377
rect 1684 329 1749 343
rect 1496 289 1548 317
rect 1699 257 1749 329
rect 1779 409 1831 457
rect 1779 375 1789 409
rect 1823 375 1831 409
rect 1779 341 1831 375
rect 1779 307 1789 341
rect 1823 307 1831 341
rect 1779 257 1831 307
<< ndiffc >>
rect 35 45 69 79
rect 119 19 153 53
rect 203 45 237 79
rect 307 19 341 53
rect 391 37 425 71
rect 501 19 535 53
rect 722 15 756 49
rect 878 35 912 69
rect 982 19 1016 53
rect 1144 21 1178 55
rect 1402 39 1436 73
rect 1506 46 1540 80
rect 1610 45 1644 79
rect 1705 19 1739 53
rect 1789 69 1823 103
<< pdiffc >>
rect 35 403 69 437
rect 35 335 69 369
rect 119 387 153 421
rect 203 403 237 437
rect 203 335 237 369
rect 307 387 341 421
rect 391 403 425 437
rect 488 410 522 444
rect 702 411 736 445
rect 798 385 832 419
rect 882 411 916 445
rect 1042 409 1076 443
rect 1222 411 1256 445
rect 1326 385 1360 419
rect 1422 385 1456 419
rect 391 335 425 369
rect 1506 385 1540 419
rect 1506 317 1540 351
rect 1610 411 1644 445
rect 1610 343 1644 377
rect 1705 411 1739 445
rect 1705 343 1739 377
rect 1789 375 1823 409
rect 1789 307 1823 341
<< poly >>
rect 79 451 109 477
rect 163 451 193 477
rect 351 457 381 483
rect 448 457 478 483
rect 532 457 562 483
rect 652 457 682 483
rect 758 457 788 483
rect 842 457 872 483
rect 926 457 956 483
rect 1002 457 1032 483
rect 1110 457 1140 483
rect 1182 457 1212 483
rect 1370 457 1400 483
rect 1466 457 1496 483
rect 1654 457 1684 483
rect 1749 457 1779 483
rect 79 308 109 323
rect 46 278 109 308
rect 46 240 76 278
rect 22 224 76 240
rect 163 234 193 323
rect 22 190 32 224
rect 66 190 76 224
rect 22 174 76 190
rect 118 224 193 234
rect 351 227 381 289
rect 448 239 478 373
rect 532 335 562 373
rect 652 341 682 373
rect 520 325 586 335
rect 520 291 536 325
rect 570 291 586 325
rect 520 281 586 291
rect 652 325 716 341
rect 652 291 672 325
rect 706 291 716 325
rect 652 275 716 291
rect 118 190 134 224
rect 168 190 193 224
rect 118 180 193 190
rect 46 136 76 174
rect 46 106 109 136
rect 79 91 109 106
rect 163 91 193 180
rect 344 211 398 227
rect 344 177 354 211
rect 388 177 398 211
rect 448 209 586 239
rect 344 161 398 177
rect 556 179 586 209
rect 351 135 381 161
rect 446 151 514 167
rect 446 117 470 151
rect 504 117 514 151
rect 446 101 514 117
rect 556 163 610 179
rect 556 129 566 163
rect 600 129 610 163
rect 556 113 610 129
rect 446 79 476 101
rect 556 79 586 113
rect 652 91 682 275
rect 758 189 788 373
rect 842 273 872 373
rect 926 273 956 373
rect 1002 335 1032 373
rect 1002 325 1068 335
rect 1002 291 1018 325
rect 1052 291 1068 325
rect 1002 281 1068 291
rect 830 257 956 273
rect 830 223 840 257
rect 874 223 956 257
rect 1110 251 1140 373
rect 1098 239 1140 251
rect 830 207 956 223
rect 1034 229 1140 239
rect 728 173 788 189
rect 728 139 738 173
rect 772 153 788 173
rect 772 139 796 153
rect 728 123 796 139
rect 766 91 796 123
rect 838 143 868 207
rect 1034 195 1050 229
rect 1084 221 1140 229
rect 1182 325 1212 373
rect 1182 309 1246 325
rect 1182 275 1202 309
rect 1236 275 1246 309
rect 1370 297 1400 373
rect 1182 251 1246 275
rect 1366 267 1400 297
rect 1182 221 1296 251
rect 1084 195 1128 221
rect 1034 185 1128 195
rect 838 107 1056 143
rect 838 91 868 107
rect 1026 91 1056 107
rect 1098 91 1128 185
rect 1170 163 1224 179
rect 1170 129 1180 163
rect 1214 129 1224 163
rect 1170 113 1224 129
rect 1194 91 1224 113
rect 1266 91 1296 221
rect 1366 189 1396 267
rect 1466 245 1496 289
rect 1654 245 1684 329
rect 1342 173 1396 189
rect 1438 229 1684 245
rect 1438 195 1448 229
rect 1482 195 1684 229
rect 1749 225 1779 257
rect 1438 179 1684 195
rect 1342 139 1352 173
rect 1386 139 1396 173
rect 1342 123 1396 139
rect 1342 91 1372 123
rect 1466 115 1496 179
rect 1654 91 1684 179
rect 1726 209 1780 225
rect 1726 175 1736 209
rect 1770 175 1780 209
rect 1726 159 1780 175
rect 1749 137 1779 159
rect 79 -19 109 7
rect 163 -19 193 7
rect 351 -19 381 7
rect 446 -19 476 7
rect 556 -19 586 7
rect 652 -19 682 7
rect 766 -19 796 7
rect 838 -19 868 7
rect 1026 -19 1056 7
rect 1098 -19 1128 7
rect 1194 -19 1224 7
rect 1266 -19 1296 7
rect 1342 -19 1372 7
rect 1466 -19 1496 7
rect 1654 -19 1684 7
rect 1749 -19 1779 7
<< polycont >>
rect 32 190 66 224
rect 536 291 570 325
rect 672 291 706 325
rect 134 190 168 224
rect 354 177 388 211
rect 470 117 504 151
rect 566 129 600 163
rect 1018 291 1052 325
rect 840 223 874 257
rect 738 139 772 173
rect 1050 195 1084 229
rect 1202 275 1236 309
rect 1180 129 1214 163
rect 1448 195 1482 229
rect 1352 139 1386 173
rect 1736 175 1770 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1133 521
rect 1167 487 1225 521
rect 1259 487 1317 521
rect 1351 487 1409 521
rect 1443 487 1501 521
rect 1535 487 1593 521
rect 1627 487 1685 521
rect 1719 487 1777 521
rect 1811 487 1869 521
rect 1903 487 1932 521
rect 35 437 69 453
rect 35 369 69 403
rect 103 421 169 487
rect 103 387 119 421
rect 153 387 169 421
rect 203 437 248 453
rect 237 403 248 437
rect 203 369 248 403
rect 291 421 357 487
rect 291 387 307 421
rect 341 387 357 421
rect 391 437 425 453
rect 686 445 762 487
rect 472 410 488 444
rect 522 410 638 444
rect 686 411 702 445
rect 736 411 762 445
rect 866 445 932 487
rect 798 419 832 435
rect 69 351 168 353
rect 69 335 122 351
rect 35 319 122 335
rect 156 317 168 351
rect 18 224 88 285
rect 18 190 32 224
rect 66 190 88 224
rect 18 155 88 190
rect 122 224 168 317
rect 122 190 134 224
rect 122 121 168 190
rect 35 87 168 121
rect 237 335 248 369
rect 391 369 425 403
rect 203 147 248 335
rect 203 113 214 147
rect 35 79 69 87
rect 203 79 248 113
rect 286 335 391 353
rect 286 319 425 335
rect 286 125 320 319
rect 470 317 494 351
rect 528 325 570 351
rect 528 317 536 325
rect 470 291 536 317
rect 354 211 436 285
rect 388 177 436 211
rect 354 161 436 177
rect 470 275 570 291
rect 470 151 514 275
rect 604 241 638 410
rect 866 411 882 445
rect 916 411 932 445
rect 1188 445 1272 487
rect 1026 409 1042 443
rect 1076 409 1152 443
rect 1188 411 1222 445
rect 1256 411 1272 445
rect 1312 419 1360 435
rect 1026 393 1152 409
rect 798 377 832 385
rect 1118 377 1152 393
rect 1312 385 1326 419
rect 1312 377 1360 385
rect 672 327 946 377
rect 672 325 722 327
rect 706 291 722 325
rect 672 275 722 291
rect 824 257 874 273
rect 824 241 840 257
rect 604 223 840 241
rect 604 207 874 223
rect 604 199 688 207
rect 286 87 425 125
rect 504 117 514 151
rect 470 101 514 117
rect 550 129 566 163
rect 600 147 620 163
rect 550 113 586 129
rect 550 89 620 113
rect 35 29 69 45
rect 103 19 119 53
rect 153 19 169 53
rect 237 45 248 79
rect 391 71 425 87
rect 203 29 248 45
rect 103 -23 169 19
rect 291 19 307 53
rect 341 19 357 53
rect 654 53 688 199
rect 908 173 946 327
rect 722 139 738 173
rect 772 147 804 173
rect 722 113 770 139
rect 722 107 804 113
rect 862 105 946 173
rect 980 351 1084 353
rect 980 325 1050 351
rect 980 291 1018 325
rect 1052 291 1084 317
rect 1118 343 1360 377
rect 1406 419 1472 487
rect 1696 445 1753 487
rect 1406 385 1422 419
rect 1456 385 1472 419
rect 1406 349 1472 385
rect 1506 419 1540 435
rect 1506 351 1540 385
rect 980 139 1014 291
rect 1048 229 1084 255
rect 1048 181 1050 229
rect 1118 241 1152 343
rect 1594 411 1610 445
rect 1644 411 1660 445
rect 1594 377 1660 411
rect 1594 343 1610 377
rect 1644 343 1660 377
rect 1506 313 1540 317
rect 1506 309 1570 313
rect 1186 275 1202 309
rect 1236 275 1570 309
rect 1118 229 1498 241
rect 1118 207 1448 229
rect 1048 173 1084 181
rect 1164 139 1180 163
rect 980 129 1180 139
rect 1214 129 1230 163
rect 980 105 1230 129
rect 862 69 912 105
rect 391 21 425 37
rect 291 -23 357 19
rect 485 19 501 53
rect 535 19 688 53
rect 485 13 688 19
rect 722 49 804 65
rect 756 15 804 49
rect 862 35 878 69
rect 862 19 912 35
rect 952 53 1016 69
rect 1264 55 1298 207
rect 1432 195 1448 207
rect 1482 195 1498 229
rect 1336 139 1352 173
rect 1386 161 1402 173
rect 1386 147 1468 161
rect 1386 139 1422 147
rect 1336 113 1422 139
rect 1456 113 1468 147
rect 1336 107 1468 113
rect 1532 96 1570 275
rect 1506 80 1570 96
rect 952 19 982 53
rect 1128 21 1144 55
rect 1178 21 1298 55
rect 1338 39 1402 73
rect 1436 39 1470 73
rect 722 -23 804 15
rect 952 -23 1016 19
rect 1338 -23 1470 39
rect 1540 46 1570 80
rect 1506 30 1570 46
rect 1610 225 1660 343
rect 1696 411 1705 445
rect 1739 411 1753 445
rect 1696 377 1753 411
rect 1696 343 1705 377
rect 1739 343 1753 377
rect 1696 327 1753 343
rect 1789 409 1840 425
rect 1823 375 1840 409
rect 1789 341 1840 375
rect 1823 307 1840 341
rect 1789 291 1840 307
rect 1610 209 1770 225
rect 1610 175 1736 209
rect 1610 159 1770 175
rect 1610 79 1660 159
rect 1804 119 1840 291
rect 1644 45 1660 79
rect 1789 103 1840 119
rect 1823 69 1840 103
rect 1610 29 1660 45
rect 1696 53 1753 69
rect 1696 19 1705 53
rect 1739 19 1753 53
rect 1696 -23 1753 19
rect 1789 13 1840 69
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1133 -23
rect 1167 -57 1225 -23
rect 1259 -57 1317 -23
rect 1351 -57 1409 -23
rect 1443 -57 1501 -23
rect 1535 -57 1593 -23
rect 1627 -57 1685 -23
rect 1719 -57 1777 -23
rect 1811 -57 1869 -23
rect 1903 -57 1932 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 857 487 891 521
rect 949 487 983 521
rect 1041 487 1075 521
rect 1133 487 1167 521
rect 1225 487 1259 521
rect 1317 487 1351 521
rect 1409 487 1443 521
rect 1501 487 1535 521
rect 1593 487 1627 521
rect 1685 487 1719 521
rect 1777 487 1811 521
rect 1869 487 1903 521
rect 122 317 156 351
rect 214 113 248 147
rect 494 317 528 351
rect 586 129 600 147
rect 600 129 620 147
rect 586 113 620 129
rect 770 139 772 147
rect 772 139 804 147
rect 770 113 804 139
rect 1050 325 1084 351
rect 1050 317 1052 325
rect 1052 317 1084 325
rect 1050 195 1084 215
rect 1050 181 1084 195
rect 1422 113 1456 147
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
rect 857 -57 891 -23
rect 949 -57 983 -23
rect 1041 -57 1075 -23
rect 1133 -57 1167 -23
rect 1225 -57 1259 -23
rect 1317 -57 1351 -23
rect 1409 -57 1443 -23
rect 1501 -57 1535 -23
rect 1593 -57 1627 -23
rect 1685 -57 1719 -23
rect 1777 -57 1811 -23
rect 1869 -57 1903 -23
<< metal1 >>
rect 0 521 1932 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1133 521
rect 1167 487 1225 521
rect 1259 487 1317 521
rect 1351 487 1409 521
rect 1443 487 1501 521
rect 1535 487 1593 521
rect 1627 487 1685 521
rect 1719 487 1777 521
rect 1811 487 1869 521
rect 1903 487 1932 521
rect 0 456 1932 487
rect 110 351 168 357
rect 110 317 122 351
rect 156 348 168 351
rect 482 351 540 357
rect 482 348 494 351
rect 156 320 494 348
rect 156 317 168 320
rect 110 311 168 317
rect 482 317 494 320
rect 528 348 540 351
rect 1038 351 1096 357
rect 1038 348 1050 351
rect 528 320 1050 348
rect 528 317 540 320
rect 482 311 540 317
rect 1038 317 1050 320
rect 1084 317 1096 351
rect 1038 311 1096 317
rect 1038 215 1096 221
rect 1038 212 1050 215
rect 589 184 1050 212
rect 589 153 632 184
rect 1038 181 1050 184
rect 1084 181 1096 215
rect 1038 175 1096 181
rect 202 147 260 153
rect 202 113 214 147
rect 248 144 260 147
rect 574 147 632 153
rect 574 144 586 147
rect 248 116 586 144
rect 248 113 260 116
rect 202 107 260 113
rect 574 113 586 116
rect 620 113 632 147
rect 574 107 632 113
rect 758 147 816 153
rect 758 113 770 147
rect 804 144 816 147
rect 1410 147 1468 153
rect 1410 144 1422 147
rect 804 116 1422 144
rect 804 113 816 116
rect 758 107 816 113
rect 1410 113 1422 116
rect 1456 113 1468 147
rect 1410 107 1468 113
rect 0 -23 1932 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1133 -23
rect 1167 -57 1225 -23
rect 1259 -57 1317 -23
rect 1351 -57 1409 -23
rect 1443 -57 1501 -23
rect 1535 -57 1593 -23
rect 1627 -57 1685 -23
rect 1719 -57 1777 -23
rect 1811 -57 1869 -23
rect 1903 -57 1932 -23
rect 0 -88 1932 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 dfstp_1
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel nwell s 46 504 46 504 3 FreeSans 400 0 0 0 VPB
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel pwell s 46 -40 46 -40 3 FreeSans 400 0 0 0 VNB
flabel locali s 402 249 436 283 0 FreeSans 200 0 0 0 D
port 9 nsew
flabel locali s 402 181 436 215 0 FreeSans 200 0 0 0 D
port 9 nsew
flabel locali s 29 487 63 521 3 FreeSans 400 0 0 0 VPWR
port 2 nsew
flabel locali s 1794 385 1828 419 0 FreeSans 400 0 0 0 Q
port 7 nsew
flabel locali s 1794 317 1828 351 0 FreeSans 400 0 0 0 Q
port 7 nsew
flabel locali s 1794 45 1828 79 0 FreeSans 400 0 0 0 Q
port 7 nsew
flabel locali s 770 113 804 147 0 FreeSans 400 0 0 0 SET_B
port 8 nsew
flabel locali s 30 249 64 283 0 FreeSans 400 0 0 0 CLK
port 10 nsew
flabel locali s 30 181 64 215 0 FreeSans 400 0 0 0 CLK
port 10 nsew
flabel locali s 29 -57 63 -23 3 FreeSans 400 0 0 0 VGND
port 3 nsew
<< properties >>
string FIXED_BBOX 0 -40 1932 504
<< end >>
