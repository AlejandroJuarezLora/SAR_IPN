* SPICE3 file created from sarlogic.ext - technology: sky130B

.subckt sar_logic VGND VPWR cal clk clkc comp ctln[0] ctln[1] ctln[2] ctln[3] ctln[4]
+ ctln[5] ctln[6] ctln[7] ctlp[0] ctlp[1] ctlp[2] ctlp[3] ctlp[4] ctlp[5] ctlp[6]
+ ctlp[7] en result[0] result[1] result[2] result[3] result[4] result[5] result[6]
+ result[7] rstn sample trim[0] trim[1] trim[2] trim[3] trim[4] trimb[0] trimb[1]
+ trimb[2] trimb[3] trimb[4] valid
X0 clknet_0_clk a_8022_7119# VPWR.t1605 VPWR.t1604 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1 VGND.t343 clknet_0_clk a_2857_7637# VGND.t342 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_745_10933# a_579_10933# VPWR.t1336 VPWR.t1335 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3 VGND.t1586 VPWR.t3333 VGND.t1585 VGND.t1584 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4 a_7710_9839# a_6633_9845# a_7548_10217# VPWR.t2809 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 trimb[4].t3 a_15023_8751# VPWR.t2716 VPWR.t2715 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6 VPWR.t2033 a_4677_7882# net15 VPWR.t2032 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X7 a_14172_1513# a_13257_1141# a_13825_1109# VGND.t2773 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X8 VGND.t2375 _066_ a_11045_5807# VGND.t2374 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X9 a_12612_8725# a_12436_9129# a_12756_9117# VGND.t462 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 a_11856_2589# _026_ VGND.t2438 VGND.t2437 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X11 a_10329_1921# a_10111_1679# VGND.t2743 VGND.t2742 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X12 VPWR.t1029 clknet_2_2__leaf_clk a_9595_1679# VPWR.t1028 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X13 _096_ _095_ a_4725_5487# VPWR.t1742 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X14 _011_ _086_ a_1137_11721# VPWR.t1030 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X15 VGND.t601 _104_ a_11321_3855# VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X16 VPWR.t2419 net2 a_14807_8359# VPWR.t2418 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_5340_6031# a_4425_6031# a_4993_6273# VGND.t3088 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X18 VGND.t2864 a_3339_2767# net45 VGND.t2863 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 a_9195_10357# net47 VPWR.t1710 VPWR.t1709 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X20 VGND.t2136 mask\[3\] a_2368_9955# VGND.t2135 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VGND.t2080 clknet_2_1__leaf_clk.t32 a_2787_9845# VGND.t2079 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X22 VGND.t3197 _082_ _007_ VGND.t3196 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 a_12061_7669# a_11895_7669# VGND.t1914 VGND.t1913 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VPWR.t942 net16 net8 VPWR.t941 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X25 mask\[5\] a_7999_11231# VGND.t3184 VGND.t3183 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X26 net23 a_1651_7093# VPWR.t2776 VPWR.t2775 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X27 VPWR.t1859 a_9802_4007# a_9478_4105# VPWR.t1858 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.28 ps=2.56 w=1 l=0.15
X28 VPWR.t2 VGND.t3254 VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X29 _063_.t3 a_8307_6575# VPWR.t2340 VPWR.t2339 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X30 a_3224_2601# a_2143_2229# a_2877_2197# VPWR.t2384 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X31 a_7197_7119# a_6007_7119# a_7088_7119# VGND.t300 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X32 _012_ a_855_4105# VPWR.t2035 VPWR.t2034 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X33 a_5535_8181# _077_ VGND.t3189 VGND.t3188 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X34 VGND.t1583 VPWR.t3334 VGND.t1582 VGND.t1581 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X35 a_3751_4765# _048_.t12 a_3388_4631# VGND.t2321 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X36 a_9099_3689# a_8583_3317# a_9004_3677# VGND.t2643 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X37 a_8083_8181# _072_ VPWR.t2801 VPWR.t2800 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X38 a_14071_3689# a_13625_3317# a_13975_3689# VGND.t2277 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X39 VGND.t1580 VPWR.t3335 VGND.t1579 VGND.t1578 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X40 VPWR.t2298 a_3868_10217# a_4043_10143# VPWR.t2297 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X41 VGND.t2015 _125_ a_15159_9269# VGND.t2014 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X42 VGND.t1577 VPWR.t3336 VGND.t1576 VGND.t1575 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X43 a_14485_7663# _132_ _133_ VPWR.t2592 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X44 VGND.t1574 VPWR.t3337 VGND.t1573 VGND.t1400 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X45 VPWR.t763 a_11059_7356# a_10990_7485# VPWR.t762 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.129 ps=1.18 w=0.84 l=0.15
X46 VGND.t1693 net47 a_10621_7119# VGND.t1692 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.064 ps=0.725 w=0.42 l=0.15
X47 a_2787_10927# _101_ a_2869_11247# VGND.t797 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X48 VPWR.t2350 _048_.t13 a_4091_5309# VPWR.t2349 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X49 VGND.t2386 net2 a_14788_7369# VGND.t2385 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X50 VPWR.t3070 net34.t2 net39 VPWR.t3069 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X51 a_4091_5309# a_4308_4917# a_4266_4943# VGND.t580 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X52 a_1000_12381# _011_ VPWR.t936 VPWR.t935 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X53 a_10676_1679# a_9761_1679# a_10329_1921# VGND.t2497 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X54 a_7902_10205# net44 VGND.t2808 VGND.t2807 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X55 VPWR.t5 VGND.t3255 VPWR.t4 VPWR.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X56 a_10903_7261# clknet_2_3__leaf_clk VGND.t1897 VGND.t1896 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X57 a_6619_7119# a_6173_7119# a_6523_7119# VGND.t808 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X58 a_9007_2601# a_8657_2229# a_8912_2589# VPWR.t1499 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X59 sample.t3 a_455_5747# VPWR.t2563 VPWR.t2562 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X60 _085_ net28 VGND.t3077 VGND.t3076 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X61 a_6181_10383# mask\[4\] VGND.t2639 VGND.t2638 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X62 _058_ a_10188_4105# VPWR.t2910 VPWR.t2909 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X63 ctlp[4].t1 a_10752_12533# VPWR.t2304 VPWR.t2303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X64 net17 a_11803_10383# VGND.t2630 VGND.t2629 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X65 a_7010_3311# trim_mask\[4\] a_6927_3311# VPWR.t1907 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X66 a_9889_6873# cal_itt\[0\] VGND.t2510 VGND.t2509 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X67 a_14335_4020# _108_ VPWR.t1537 VPWR.t1536 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X68 VGND.t2828 a_2283_4020# _013_ VGND.t2827 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X69 VGND.t1572 VPWR.t3338 VGND.t1571 VGND.t1030 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X70 a_9103_2601# a_8657_2229# a_9007_2601# VGND.t747 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X71 trim_val\[0\] a_14347_4917# VGND.t545 VGND.t544 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X72 a_1279_9129# a_763_8757# a_1184_9117# VGND.t85 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X73 a_7891_3617# _050_ VPWR.t2623 VPWR.t2622 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X74 a_2815_9447# mask\[2\] a_2961_9545# VPWR.t3190 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X75 net22 a_1651_6005# VPWR.t2892 VPWR.t2891 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X76 _092_ a_10005_6031# VGND.t71 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X77 VPWR.t2621 _050_ a_6763_5193# VPWR.t2620 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X78 VPWR.t1332 a_4863_4917# _095_ VPWR.t1331 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X79 VPWR.t8 VGND.t3256 VPWR.t7 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X80 VPWR.t11 VGND.t3257 VPWR.t10 VPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X81 a_14564_6397# a_14379_6397# VPWR.t2788 VPWR.t2787 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0767 ps=0.785 w=0.42 l=0.15
X82 a_7942_2223# a_7223_2465# a_7379_2197# VGND.t2369 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X83 a_11233_4405# a_11067_4405# VPWR.t2598 VPWR.t2597 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X84 a_10137_4943# net30.t4 _118_ VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X85 VGND.t2516 a_7723_10143# a_7657_10217# VGND.t2515 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X86 trim[1].t7 a_15083_4659# VGND.t2253 VGND.t2252 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X87 ctlp[6].t7 a_6927_12559# VGND.t2245 VGND.t2244 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X88 VGND.t2450 a_448_9269# result[3].t3 VGND.t2449 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X89 VPWR.t14 VGND.t3258 VPWR.t13 VPWR.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X90 net52 a_5691_7637# VPWR.t2639 VPWR.t2638 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X91 a_7715_3285# a_7891_3617# a_7843_3677# VGND.t2461 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X92 a_1638_6397# a_561_6031# a_1476_6031# VPWR.t2625 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X93 VPWR.t1519 a_14172_4943# a_14347_4917# VPWR.t1518 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X94 a_2014_12381# net43.t8 VGND.t626 VGND.t625 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X95 VPWR.t2431 net52 a_2225_7663# VPWR.t2430 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X96 VPWR.t1438 a_2857_5461# clknet_2_0__leaf_clk VPWR.t1437 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X97 VGND.t1570 VPWR.t3339 VGND.t1569 VGND.t854 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X98 VGND.t1624 a_10747_8970# _035_ VGND.t1623 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X99 net7 net15 VGND.t1869 VGND.t1868 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X100 a_3977_7119# a_2787_7119# a_3868_7119# VGND.t2832 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X101 VPWR.t2155 a_8298_5487# clknet_2_3__leaf_clk VPWR.t2154 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X102 VGND.t684 a_2857_5461# clknet_2_0__leaf_clk VGND.t683 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X103 VGND.t715 net9 a_12631_591# VGND.t714 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X104 a_13881_2741# trim_val\[1\] VGND.t176 VGND.t175 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X105 VPWR.t2896 a_13059_4631# _111_ VPWR.t2895 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X106 clknet_2_1__leaf_clk.t31 a_2857_7637# VGND.t375 VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X107 a_13142_8725# a_12992_8751# VPWR.t1291 VPWR.t1290 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X108 VPWR.t2609 _053_ a_11098_6691# VPWR.t2608 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X109 result[6].t7 a_455_12533# VGND.t2446 VGND.t2445 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X110 VGND.t1568 VPWR.t3340 VGND.t1567 VGND.t1566 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X111 a_1493_5487# net22 _079_ VPWR.t3169 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X112 VPWR.t2103 clknet_2_1__leaf_clk.t33 a_3431_10933# VPWR.t2102 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X113 VPWR.t2969 a_13519_4007# _113_ VPWR.t2968 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X114 a_4609_9295# a_4443_9295# VPWR.t1935 VPWR.t1934 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X115 a_8270_8029# net43.t9 VGND.t628 VGND.t627 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X116 VPWR.t1603 a_8022_7119# clknet_0_clk VPWR.t1602 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X117 _096_ _092_ VGND.t2824 VGND.t2823 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X118 a_14249_8725# _125_ VGND.t2013 VGND.t2012 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X119 a_14181_6031# _134_ VGND.t1839 VGND.t1838 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X120 VPWR.t1080 clknet_0_clk a_8298_2767# VPWR.t1079 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X121 a_9207_3311# net46 VPWR.t995 VPWR.t994 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X122 VGND.t2495 net45 a_4995_7119# VGND.t2494 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X123 a_4886_4399# net54 VPWR.t1404 VPWR.t1403 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X124 VGND.t2608 a_1835_12319# a_1769_12393# VGND.t2607 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X125 a_3781_8207# a_3615_8207# VGND.t1669 VGND.t1668 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X126 VPWR.t2534 a_14981_4020# net31 VPWR.t2533 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X127 VPWR.t1921 clknet_2_3__leaf_clk a_14379_6397# VPWR.t1920 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.109 ps=1.36 w=0.42 l=0.15
X128 VGND.t1691 net47 a_8717_10383# VGND.t1690 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X129 VPWR.t17 VGND.t3259 VPWR.t16 VPWR.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X130 ctln[6].t7 a_6927_591# VGND.t1788 VGND.t1787 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X131 _022_ a_2787_10927# VPWR.t1788 VPWR.t1787 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X132 a_1007_10217# a_561_9845# a_911_10217# VGND.t3111 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X133 a_4239_8573# a_3615_8207# a_4131_8207# VPWR.t1686 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X134 a_9458_9661# a_8381_9295# a_9296_9295# VPWR.t3309 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X135 VPWR.t2051 a_15023_10927# trimb[0].t3 VPWR.t2050 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X136 a_4775_6031# a_4425_6031# a_4680_6031# VPWR.t3161 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X137 VPWR.t3183 net11 a_8767_591# VPWR.t3182 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X138 _126_ a_14236_8457# VGND.t2556 VGND.t2555 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X139 VGND.t2354 _065_.t4 _101_ VGND.t2353 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X140 a_14335_2442# _108_ VPWR.t1535 VPWR.t1534 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X141 a_13512_4943# _029_ VPWR.t748 VPWR.t747 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X142 _103_ _092_ VGND.t2822 VGND.t2821 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X143 a_3557_5193# _092_ a_3461_5193# VPWR.t2868 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X144 VPWR.t20 VGND.t3260 VPWR.t19 VPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X145 a_7223_2465# clknet_2_2__leaf_clk VGND.t290 VGND.t289 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X146 _098_ a_6210_4989# VGND.t3094 VGND.t3093 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X147 _104_ net30.t5 VPWR.t765 VPWR.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X148 VPWR.t2569 a_1476_10217# a_1651_10143# VPWR.t2568 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X149 a_13100_8751# a_12153_8757# a_12992_8751# VPWR.t1239 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X150 trim_mask\[0\] a_12323_4703# VPWR.t3256 VPWR.t3255 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X151 VGND.t288 clknet_2_2__leaf_clk a_9595_1679# VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X152 VPWR.t1027 clknet_2_2__leaf_clk a_13459_3317# VPWR.t1026 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X153 VPWR.t23 VGND.t3261 VPWR.t22 VPWR.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X154 trim_val\[2\] a_14347_1439# VGND.t3195 VGND.t3194 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X155 a_9503_4399# _107_ _108_ VPWR.t1682 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X156 VGND.t257 net46 a_13869_4943# VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X157 VGND.t1565 VPWR.t3341 VGND.t1564 VGND.t1563 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X158 VPWR.t26 VGND.t3262 VPWR.t25 VPWR.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X159 VGND.t1562 VPWR.t3342 VGND.t1561 VGND.t1560 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X160 VGND.t1559 VPWR.t3343 VGND.t1558 VGND.t1557 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X161 VGND.t341 clknet_0_clk a_8298_5487# VGND.t340 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X162 VPWR.t29 VGND.t3263 VPWR.t28 VPWR.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X163 VGND.t2670 a_15023_8751# trimb[4].t7 VGND.t2669 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X164 a_6909_10933# a_6743_10933# VPWR.t2573 VPWR.t2572 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X165 a_12169_2197# a_11951_2601# VPWR.t928 VPWR.t927 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X166 trim_mask\[2\] a_12691_2527# VPWR.t955 VPWR.t954 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X167 a_1095_11305# a_745_10933# a_1000_11293# VPWR.t1720 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X168 a_2601_3285# a_2383_3689# VPWR.t1810 VPWR.t1809 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X169 VPWR.t2072 a_5363_12559# ctlp[7].t3 VPWR.t2071 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X170 a_8105_10383# a_7939_10383# VPWR.t946 VPWR.t945 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X171 clknet_2_1__leaf_clk.t15 a_2857_7637# VPWR.t1112 VPWR.t1111 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X172 a_14335_4020# _108_ VGND.t781 VGND.t780 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X173 a_12522_8751# a_11987_8757# a_12436_9129# VPWR.t2937 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X174 a_9459_7895# _067_ VPWR.t924 VPWR.t923 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.34 w=0.42 l=0.15
X175 a_14199_7369# _129_ VPWR.t1564 VPWR.t1563 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X176 a_4959_1679# a_4609_1679# a_4864_1679# VPWR.t2914 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X177 VGND.t59 trim_val\[3\] a_11292_1251# VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X178 a_4883_6397# a_4259_6031# a_4775_6031# VPWR.t1048 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X179 VPWR.t32 VGND.t3264 VPWR.t31 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X180 VGND.t2460 a_4687_11231# a_4621_11305# VGND.t2459 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X181 clknet_0_clk a_8022_7119# VPWR.t1601 VPWR.t1600 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X182 net5 a_15023_6031# VPWR.t1392 VPWR.t1391 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X183 VPWR.t35 VGND.t3265 VPWR.t34 VPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X184 VGND.t2655 a_448_10357# result[4].t3 VGND.t2654 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X185 a_8298_2767# clknet_0_clk VPWR.t1078 VPWR.t1077 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X186 VGND.t1556 VPWR.t3344 VGND.t1555 VGND.t1554 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X187 a_4864_9295# _019_ VGND.t2877 VGND.t2876 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X188 VPWR.t38 VGND.t3266 VPWR.t37 VPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X189 a_5177_1921# a_4959_1679# VPWR.t2797 VPWR.t2796 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X190 a_9503_4399# _106_ VPWR.t757 VPWR.t756 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X191 a_12257_4777# a_11067_4405# a_12148_4777# VGND.t2560 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X192 VPWR.t2651 a_1835_12319# a_1822_12015# VPWR.t2650 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X193 _034_ a_4167_6575# VPWR.t3264 VPWR.t3263 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X194 VGND.t816 a_10055_2767# net46 VGND.t815 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X195 a_6633_9845# a_6467_9845# VPWR.t2489 VPWR.t2488 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X196 VGND.t1553 VPWR.t3345 VGND.t1552 VGND.t1367 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X197 a_7442_7119# net44 VGND.t2806 VGND.t2805 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X198 VPWR.t41 VGND.t3267 VPWR.t40 VPWR.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X199 VPWR.t44 VGND.t3268 VPWR.t43 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X200 VGND.t1551 VPWR.t3346 VGND.t1550 VGND.t1549 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X201 VPWR.t47 VGND.t3269 VPWR.t46 VPWR.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X202 VPWR.t2547 cal_itt\[0\] a_9957_7663# VPWR.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X203 VPWR.t50 VGND.t3270 VPWR.t49 VPWR.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X204 VPWR.t53 VGND.t3271 VPWR.t52 VPWR.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X205 VPWR.t2703 a_8949_9537# a_8839_9661# VPWR.t2702 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X206 VPWR.t3250 a_14249_8725# _129_ VPWR.t3249 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X207 a_11575_8790# _123_.t3 a_11116_8983# VPWR.t1654 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X208 _051_.t5 a_3933_2767# VPWR.t1251 VPWR.t1250 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X209 VPWR.t2365 a_13697_4373# _109_ VPWR.t2364 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X210 VGND.t2547 a_5691_2741# _050_ VGND.t2546 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X211 a_9839_3615# a_9664_3689# a_10018_3677# VGND.t2744 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X212 a_12516_2601# a_11435_2229# a_12169_2197# VPWR.t1754 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X213 _094_ mask\[0\] VGND.t2994 VGND.t2993 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X214 _059_ net55 VGND.t2965 VGND.t2964 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X215 VPWR.t56 VGND.t3272 VPWR.t55 VPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X216 a_2948_3689# a_1867_3317# a_2601_3285# VPWR.t1947 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X217 VPWR.t59 VGND.t3273 VPWR.t58 VPWR.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X218 a_5691_7637# net51 VGND.t392 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X219 a_14335_2442# _108_ VGND.t779 VGND.t778 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X220 VPWR.t2967 _045_ a_6191_12559# VPWR.t2966 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X221 VGND.t2432 a_8298_2767# clknet_2_2__leaf_clk VGND.t2431 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X222 VGND.t2499 a_14981_4020# net31 VGND.t2498 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X223 VPWR.t1919 clknet_2_3__leaf_clk a_11987_8757# VPWR.t1918 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X224 a_1129_9813# a_911_10217# VPWR.t2815 VPWR.t2814 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X225 net26 a_7723_10143# VGND.t2514 VGND.t2513 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X226 a_13607_1513# a_13257_1141# a_13512_1501# VPWR.t2819 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X227 VPWR.t62 VGND.t3274 VPWR.t61 VPWR.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X228 clknet_2_1__leaf_clk.t14 a_2857_7637# VPWR.t1110 VPWR.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X229 a_11679_4777# a_11233_4405# a_11583_4777# VGND.t1854 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X230 a_11479_9117# _122_ a_11116_8983# VGND.t2072 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X231 cal_count\[3\] a_12231_6005# VPWR.t904 VPWR.t903 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X232 VGND.t3222 a_12599_3615# a_12533_3689# VGND.t3221 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X233 a_11244_9661# a_10405_9295# a_11268_9295# VGND.t1820 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X234 VPWR.t65 VGND.t3275 VPWR.t64 VPWR.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X235 _044_ a_8072_11721# VPWR.t2203 VPWR.t2202 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X236 a_845_7663# _080_ _005_ VPWR.t2965 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X237 a_3388_4631# _048_.t14 a_3530_4438# VPWR.t2351 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X238 a_8298_5487# clknet_0_clk VGND.t339 VGND.t338 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X239 trimb[4].t6 a_15023_8751# VGND.t2668 VGND.t2667 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X240 a_8307_4719# _103_ VGND.t1696 VGND.t1695 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X241 a_2689_8751# net24 _081_ VPWR.t3236 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X242 VPWR.t68 VGND.t3276 VPWR.t67 VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X243 a_13975_3689# a_13625_3317# a_13880_3677# VPWR.t2306 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X244 a_11859_3689# a_11509_3317# a_11764_3677# VPWR.t2283 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X245 VPWR.t2186 a_15023_12015# trimb[2].t3 VPWR.t2185 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X246 a_5915_11721# mask\[5\] VPWR.t2502 VPWR.t2501 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X247 VPWR.t3285 a_7088_7119# a_7263_7093# VPWR.t3284 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X248 a_3057_4719# a_2865_4460# _014_ VGND.t2981 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X249 VPWR.t3328 a_15023_9839# trimb[1].t3 VPWR.t3327 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X250 net44 a_4995_7119# VGND.t23 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X251 VPWR.t1640 cal_itt\[1\] _063_.t1 VPWR.t1639 sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X252 _090_ _089_ VGND.t1734 VGND.t1733 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X253 _024_ a_10975_4105# VPWR.t1148 VPWR.t1147 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X254 _108_ _107_ VGND.t1665 VGND.t1664 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X255 VGND.t1548 VPWR.t3347 VGND.t1547 VGND.t1546 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X256 a_8301_8207# cal_itt\[2\] VGND.t2987 VGND.t2986 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X257 VPWR.t3200 a_7939_3855# net30.t1 VPWR.t3199 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X258 VGND.t203 net16 a_14471_12559# VGND.t202 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X259 VPWR.t1965 a_1660_11305# a_1835_11231# VPWR.t1964 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X260 VPWR.t71 VGND.t3277 VPWR.t70 VPWR.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X261 VPWR.t3090 a_1276_565# ctln[0].t1 VPWR.t3089 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X262 a_4175_4943# _048_.t15 a_4091_4943# VGND.t2322 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.0567 ps=0.69 w=0.42 l=0.15
X263 VPWR.t74 VGND.t3278 VPWR.t73 VPWR.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X264 VPWR.t1235 a_15023_5487# trim[4].t3 VPWR.t1234 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X265 valid.t7 a_455_3571# VGND.t2169 VGND.t2168 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X266 a_8381_9295# a_8215_9295# VGND.t1936 VGND.t1935 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X267 a_13142_7271# _123_.t4 a_13356_7369# VPWR.t1655 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X268 VPWR.t2725 _135_ a_13783_6183# VPWR.t2724 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X269 a_11149_3017# trim_mask\[3\] a_11067_3017# VPWR.t2101 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X270 a_1313_11989# a_1095_12393# VGND.t2624 VGND.t2623 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X271 VGND.t1545 VPWR.t3348 VGND.t1544 VGND.t1394 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X272 VPWR.t2898 a_9889_6873# a_9919_6614# VPWR.t2897 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X273 a_3748_6281# _120_ VGND.t2904 VGND.t2903 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X274 a_12056_6031# a_11141_6031# a_11709_6273# VGND.t2737 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X275 _048_.t5 a_3667_3829# VPWR.t3299 VPWR.t3298 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X276 ctlp[6].t6 a_6927_12559# VGND.t2243 VGND.t2242 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X277 a_1476_10217# a_395_9845# a_1129_9813# VPWR.t2115 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X278 trim[3].t3 a_15023_1135# VPWR.t2738 VPWR.t2737 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X279 a_4864_1679# _015_ VGND.t395 VGND.t394 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X280 a_13715_1135# a_13091_1141# a_13607_1513# VPWR.t1277 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X281 a_4801_9839# net53 VPWR.t1851 VPWR.t1850 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X282 a_3530_4438# _096_ VPWR.t1044 VPWR.t1043 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X283 VGND.t1895 clknet_2_3__leaf_clk a_11895_7669# VGND.t1894 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X284 VGND.t2804 net44 a_7153_12381# VGND.t2803 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X285 a_1467_7923# net45 VPWR.t2530 VPWR.t2529 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X286 a_14000_4719# trim_mask\[0\] a_13697_4373# VGND.t1876 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X287 VPWR.t1436 a_2857_5461# clknet_2_0__leaf_clk VPWR.t1435 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X288 VGND.t1543 VPWR.t3349 VGND.t1542 VGND.t1352 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X289 a_10207_1679# a_9761_1679# a_10111_1679# VGND.t2496 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X290 VGND.t682 a_2857_5461# clknet_2_0__leaf_clk VGND.t681 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X291 a_7569_7637# a_7351_8041# VPWR.t1253 VPWR.t1252 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X292 VGND.t459 a_2313_6183# _039_ VGND.t458 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X293 a_15111_9295# _126_ VGND.t75 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X294 cal_itt\[2\] a_8091_7967# VPWR.t1855 VPWR.t1854 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X295 a_3273_4943# en_co_clk VPWR.t2661 VPWR.t2660 sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.42 as=0.345 ps=2.69 w=1 l=0.15
X296 a_14318_8457# cal_count\[1\] a_14236_8457# VPWR.t2201 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X297 a_14184_1679# trim_mask\[2\] a_13881_1653# VGND.t2842 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X298 a_6737_4719# calibrate VGND.t743 VGND.t742 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X299 VGND.t377 net12 a_6927_591# VGND.t376 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X300 a_11967_3311# a_11343_3317# a_11859_3689# VPWR.t2263 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X301 a_9747_2527# a_9572_2601# a_9926_2589# VGND.t2907 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X302 a_10405_9295# a_10239_9295# VGND.t3018 VGND.t3017 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X303 VGND.t1541 VPWR.t3350 VGND.t1540 VGND.t1539 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X304 a_2857_7637# clknet_0_clk VGND.t337 VGND.t336 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X305 a_3399_10217# a_2953_9845# a_3303_10217# VGND.t1943 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X306 a_1045_9545# _074_ VPWR.t890 VPWR.t889 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X307 _074_ a_5423_9011# VGND.t3036 VGND.t3035 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X308 VPWR.t2714 a_15023_8751# trimb[4].t2 VPWR.t2713 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X309 a_1660_12393# a_745_12021# a_1313_11989# VGND.t3144 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X310 VGND.t1538 VPWR.t3351 VGND.t1537 VGND.t1536 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X311 VPWR.t77 VGND.t3279 VPWR.t76 VPWR.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X312 VGND.t1926 a_6885_8372# net51 VGND.t1925 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X313 VPWR.t2930 a_4471_4007# _015_ VPWR.t2929 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X314 VPWR.t1210 a_1461_10357# _023_ VPWR.t1209 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X315 _021_ a_5915_10927# VPWR.t783 VPWR.t782 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X316 _001_ _069_ VGND.t3024 VGND.t3023 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X317 a_12410_6031# net46 VGND.t255 VGND.t254 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X318 VGND.t3253 a_5087_3855# net54 VGND.t3252 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X319 VGND.t2324 _048_.t16 _049_ VGND.t2323 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X320 a_4043_10143# a_3868_10217# a_4222_10205# VGND.t2270 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X321 a_6428_7119# _003_ VPWR.t2084 VPWR.t2083 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X322 _098_ calibrate VGND.t741 VGND.t740 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X323 VGND.t2260 net36 a_15023_10927# VGND.t2259 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X324 VGND.t2622 net33 a_15023_2223# VGND.t80 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X325 a_5578_12131# net28 a_5496_12131# VPWR.t3142 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X326 a_8178_11293# net44 VGND.t2802 VGND.t2801 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X327 VGND.t1535 VPWR.t3352 VGND.t1534 VGND.t848 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X328 trimb[1].t2 a_15023_9839# VPWR.t3326 VPWR.t3325 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X329 a_14422_7093# _131_ VGND.t3022 VGND.t3021 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.136 ps=1.1 w=0.42 l=0.15
X330 result[0].t1 a_448_6549# VPWR.t2772 VPWR.t2771 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X331 a_4471_4007# _100_ a_4617_4105# VPWR.t3064 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X332 ctlp[7].t2 a_5363_12559# VPWR.t2070 VPWR.t2069 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X333 a_4425_6031# a_4259_6031# VPWR.t1047 VPWR.t1046 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X334 a_7456_12393# a_6375_12021# a_7109_11989# VPWR.t3063 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X335 VPWR.t79 VGND.t3280 VPWR.t78 VPWR.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X336 _041_ a_3840_8867# VPWR.t2259 VPWR.t2258 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X337 a_10569_1109# trim_val\[3\] VGND.t57 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X338 a_7916_8041# a_6835_7669# a_7569_7637# VPWR.t792 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X339 a_4165_10901# a_3947_11305# VGND.t1705 VGND.t1704 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X340 a_2953_9845# a_2787_9845# VPWR.t1009 VPWR.t1008 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X341 a_10864_9269# net47 VPWR.t1708 VPWR.t1707 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X342 _136_ a_13783_6183# VPWR.t2720 VPWR.t2719 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.36 ps=2.72 w=1 l=0.15
X343 VGND.t335 clknet_0_clk a_2857_5461# VGND.t334 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X344 a_4043_7093# net43.t10 VPWR.t1380 VPWR.t1379 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X345 VGND.t1533 VPWR.t3353 VGND.t1532 VGND.t1531 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X346 a_4091_5309# a_3891_4943# VPWR.t1943 VPWR.t1942 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0588 ps=0.7 w=0.42 l=0.15
X347 VPWR.t1780 clknet_2_0__leaf_clk a_6007_7119# VPWR.t1779 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X348 a_11168_9661# a_10688_9295# VPWR.t894 VPWR.t893 sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X349 VPWR.t1808 a_6927_591# ctln[6].t3 VPWR.t1807 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X350 VPWR.t82 VGND.t3281 VPWR.t81 VPWR.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X351 a_3116_12533# net15 VGND.t1867 VGND.t1866 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X352 VGND.t1530 VPWR.t3354 VGND.t1529 VGND.t1528 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X353 VPWR.t2706 a_14807_8359# _125_ VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X354 VPWR.t85 VGND.t3282 VPWR.t84 VPWR.t83 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X355 VGND.t1527 VPWR.t3355 VGND.t1526 VGND.t1525 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X356 VPWR.t2561 a_455_5747# sample.t2 VPWR.t2560 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X357 net9 net17 VPWR.t2825 VPWR.t2824 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X358 VGND.t1524 VPWR.t3356 VGND.t1523 VGND.t1522 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X359 ctln[5].t3 a_8767_591# VGND.t2360 VGND.t2359 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X360 VPWR.t3175 a_7379_2197# a_7310_2223# VPWR.t3174 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.129 ps=1.18 w=0.84 l=0.15
X361 a_4658_3427# state\[0\] a_4576_3427# VPWR.t1459 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X362 a_7010_3311# _104_ a_7010_3631# VGND.t599 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.0683 ps=0.86 w=0.65 l=0.15
X363 VGND.t1715 a_4871_8181# a_4805_8207# VGND.t1714 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X364 a_911_4777# a_561_4405# a_816_4765# VPWR.t1951 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X365 a_10781_3311# trim_mask\[1\] VPWR.t872 VPWR.t871 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X366 VGND.t373 a_2857_7637# clknet_2_1__leaf_clk.t30 VGND.t372 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X367 a_7262_5461# _051_.t12 VPWR.t2758 VPWR.t2757 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.176 ps=1.39 w=0.42 l=0.15
X368 trimb[4].t1 a_15023_8751# VPWR.t2712 VPWR.t2711 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X369 a_4393_8207# a_4349_8449# a_4227_8207# VGND.t2974 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X370 VGND.t1521 VPWR.t3357 VGND.t1520 VGND.t1519 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X371 VGND.t2251 a_15083_4659# trim[1].t6 VGND.t2250 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X372 trim_val\[3\] a_10851_1653# VPWR.t1152 VPWR.t1151 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X373 a_10781_5487# _092_ a_10699_5487# VPWR.t2867 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X374 a_7088_7119# a_6007_7119# a_6741_7361# VPWR.t1037 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X375 a_1019_6397# a_395_6031# a_911_6031# VPWR.t1301 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X376 a_7715_3285# _051_.t13 VPWR.t2760 VPWR.t2759 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X377 ctlp[5].t1 a_8820_12533# VPWR.t3244 VPWR.t3243 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X378 result[4].t2 a_448_10357# VGND.t2653 VGND.t2652 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X379 VPWR.t88 VGND.t3283 VPWR.t87 VPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X380 a_10689_2543# _104_ VGND.t598 VGND.t597 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X381 VPWR.t2924 a_5547_5603# _075_ VPWR.t2923 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X382 _092_ a_10005_6031# VGND.t69 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X383 _057_ a_11292_1251# VPWR.t2587 VPWR.t2586 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X384 clknet_2_0__leaf_clk a_2857_5461# VGND.t680 VGND.t679 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X385 VGND.t3052 _078_ a_2775_9071# VGND.t3051 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X386 VGND.t371 a_2857_7637# clknet_2_1__leaf_clk.t29 VGND.t370 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X387 VPWR.t91 VGND.t3284 VPWR.t90 VPWR.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X388 a_10018_3677# net46 VGND.t253 VGND.t252 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X389 a_4617_3855# _060_ VGND.t2206 VGND.t2205 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X390 net18 a_9871_10383# VPWR.t1297 VPWR.t1296 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X391 VPWR.t2685 mask\[4\] a_4801_9839# VPWR.t2684 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X392 a_10005_6031# _091_ VGND.t565 VGND.t564 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X393 VGND.t847 a_8022_7119# clknet_0_clk VGND.t846 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X394 VGND.t1518 VPWR.t3358 VGND.t1517 VGND.t1516 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X395 VPWR.t1446 _028_ a_7942_2223# VPWR.t1445 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X396 VPWR.t761 a_4995_7119# net44 VPWR.t760 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X397 VGND.t688 a_14471_591# ctln[2].t3 VGND.t687 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X398 VPWR.t1146 _055_ a_15299_3311# VPWR.t1145 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X399 VPWR.t2904 _113_ a_13183_3311# VPWR.t2903 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X400 a_13349_6031# net2 VGND.t2384 VGND.t2383 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X401 clknet_2_2__leaf_clk a_8298_2767# VPWR.t2465 VPWR.t2464 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X402 VGND.t3203 a_7019_4407# net55 VGND.t3202 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X403 a_5536_4399# _048_.t17 a_5363_4719# VGND.t2325 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X404 VGND.t1515 VPWR.t3359 VGND.t1514 VGND.t1513 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X405 VGND.t1689 net47 a_13256_9117# VGND.t1688 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
X406 VPWR.t1786 a_2948_3689# a_3123_3615# VPWR.t1785 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X407 VPWR.t2207 a_7201_9813# a_7091_9839# VPWR.t2206 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X408 VPWR.t1778 clknet_2_0__leaf_clk a_2787_7119# VPWR.t1777 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X409 ctln[7].t7 a_5363_591# VGND.t1849 VGND.t1848 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X410 VGND.t476 net32 net37.t3 VGND.t475 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X411 a_8495_6895# cal_itt\[2\] a_8745_6895# VGND.t2985 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X412 VGND.t1512 VPWR.t3360 VGND.t1511 VGND.t1510 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X413 a_3840_8867# net24 VGND.t3160 VGND.t3159 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X414 a_9374_10383# net47 VGND.t1687 VGND.t1686 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X415 a_11030_1679# net46 VGND.t251 VGND.t250 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X416 VPWR.t94 VGND.t3285 VPWR.t93 VPWR.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X417 a_11488_4765# _024_ VPWR.t2107 VPWR.t2106 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X418 net6 net14 VPWR.t1959 VPWR.t1958 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X419 _104_ _103_ VPWR.t1714 VPWR.t1713 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X420 a_11023_5108# _108_ VPWR.t1533 VPWR.t1532 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X421 a_2869_10927# mask\[7\] VPWR.t3029 VPWR.t3028 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X422 _017_ a_2971_8457# VGND.t1767 VGND.t1766 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X423 VPWR.t97 VGND.t3286 VPWR.t96 VPWR.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X424 a_7104_3855# _052_ VGND.t384 VGND.t383 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X425 a_6987_12393# a_6541_12021# a_6891_12393# VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X426 VGND.t1509 VPWR.t3361 VGND.t1508 VGND.t1507 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X427 _054_ a_7190_3855# VPWR.t1949 VPWR.t1948 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X428 VGND.t2812 a_1651_10143# a_1585_10217# VGND.t2811 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X429 a_11599_6397# a_10975_6031# a_11491_6031# VPWR.t2211 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X430 a_11801_4373# a_11583_4777# VPWR.t2928 VPWR.t2927 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X431 VPWR.t1178 a_5699_9269# a_5686_9661# VPWR.t1177 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X432 a_3053_8207# mask\[1\] VGND.t1780 VGND.t1779 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X433 VPWR.t3270 a_14564_6397# _061_ VPWR.t3269 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X434 _043_ a_8992_9955# VPWR.t2718 VPWR.t2717 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X435 a_10688_9295# a_10405_9295# a_10593_9295# VPWR.t1844 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X436 VPWR.t2233 _044_ a_8767_11471# VPWR.t2232 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X437 VGND.t2007 a_11116_8983# _124_ VGND.t2006 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X438 a_4239_8573# net44 VPWR.t2855 VPWR.t2854 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X439 a_3868_7119# a_2787_7119# a_3521_7361# VPWR.t2876 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X440 VGND.t2493 net45 a_6941_2589# VGND.t2492 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.064 ps=0.725 w=0.42 l=0.15
X441 a_3388_4631# _090_ a_3530_4765# VGND.t400 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X442 a_7245_10205# a_7201_9813# a_7079_10217# VGND.t2180 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X443 VGND.t1506 VPWR.t3362 VGND.t1505 VGND.t1504 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X444 a_7631_12319# a_7456_12393# a_7810_12381# VGND.t2285 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X445 VPWR.t2795 net8 a_14471_591# VPWR.t2794 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X446 _066_ _065_.t5 VGND.t2356 VGND.t2355 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X447 VPWR.t1541 a_4043_7093# a_4030_7485# VPWR.t1540 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X448 trim[1].t5 a_15083_4659# VGND.t2249 VGND.t2248 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X449 VPWR.t1187 a_6056_8359# _077_ VPWR.t1186 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X450 a_6198_8534# _076_ VPWR.t1226 VPWR.t1225 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X451 a_9369_3855# _108_ VGND.t777 VGND.t776 sky130_fd_pr__nfet_01v8 ad=0.275 pd=1.5 as=0.0878 ps=0.92 w=0.65 l=0.15
X452 a_8820_6005# cal_itt\[1\] a_9043_6031# VGND.t1620 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X453 VPWR.t100 VGND.t3287 VPWR.t99 VPWR.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X454 _105_ _048_.t18 VPWR.t2353 VPWR.t2352 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X455 clknet_2_3__leaf_clk a_8298_5487# VGND.t2130 VGND.t2129 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X456 ctlp[0].t7 a_1099_12533# VGND.t723 VGND.t722 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X457 VGND.t1503 VPWR.t3363 VGND.t1502 VGND.t1501 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X458 a_11845_4765# a_11801_4373# a_11679_4777# VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X459 trimb[2].t7 a_15023_12015# VGND.t2159 VGND.t2158 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X460 a_5177_9537# a_4959_9295# VGND.t87 VGND.t86 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X461 a_13825_5185# a_13607_4943# VPWR.t2285 VPWR.t2284 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X462 VPWR.t1324 a_4308_4917# a_4091_5309# VPWR.t1323 sky130_fd_pr__pfet_01v8_hvt ad=0.331 pd=1.71 as=0.0672 ps=0.74 w=0.42 l=0.15
X463 _064_ _062_.t8 VGND.t2228 VGND.t2227 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X464 a_4030_9839# a_2953_9845# a_3868_10217# VPWR.t1971 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X465 VPWR.t2386 _065_.t6 a_9761_8457# VPWR.t2385 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X466 a_6198_8207# _076_ VGND.t485 VGND.t484 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X467 VPWR.t1108 a_2857_7637# clknet_2_1__leaf_clk.t13 VPWR.t1107 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X468 VGND.t1500 VPWR.t3364 VGND.t1499 VGND.t1498 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X469 VPWR.t2153 a_8298_5487# clknet_2_3__leaf_clk VPWR.t2152 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X470 VPWR.t1170 a_12520_7637# a_12430_7663# VPWR.t1169 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X471 a_3852_12381# _010_ VGND.t2826 VGND.t2825 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X472 VPWR.t1485 a_5535_8181# _078_ VPWR.t1484 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X473 VPWR.t103 VGND.t3288 VPWR.t102 VPWR.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X474 a_1585_4777# a_395_4405# a_1476_4777# VGND.t2200 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X475 a_10195_1354# _117_ VGND.t1622 VGND.t1621 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X476 VPWR.t106 VGND.t3289 VPWR.t105 VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X477 VGND.t511 a_3933_2767# _051_.t11 VGND.t510 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X478 a_14715_3615# a_14540_3689# a_14894_3677# VGND.t2837 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X479 a_12599_3615# a_12424_3689# a_12778_3677# VGND.t2231 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X480 a_14604_2339# trim_mask\[2\] VGND.t2841 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X481 a_3399_2527# net45 VPWR.t2528 VPWR.t2527 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X482 _103_ net42 a_7393_5193# VPWR.t773 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X483 net5 a_15023_6031# VGND.t639 VGND.t638 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X484 VGND.t2192 net20.t2 a_6927_12559# VGND.t2191 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X485 cal_count\[1\] a_13562_8751# VPWR.t1503 VPWR.t1502 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X486 VGND.t1764 clknet_2_0__leaf_clk a_6007_7119# VGND.t1763 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X487 a_9503_4399# _106_ VPWR.t755 VPWR.t754 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X488 VPWR.t1599 a_8022_7119# clknet_0_clk VPWR.t1598 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X489 a_12148_4777# a_11067_4405# a_11801_4373# VPWR.t2596 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X490 a_12249_7663# _037_ VGND.t97 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X491 VPWR.t1076 clknet_0_clk a_8298_2767# VPWR.t1075 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X492 a_1357_12381# a_1313_11989# a_1191_12393# VGND.t2693 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X493 a_8563_10749# net47 VPWR.t1706 VPWR.t1705 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X494 a_455_12533# net28 VGND.t3075 VGND.t3074 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X495 a_11488_4765# _024_ VGND.t2082 VGND.t2081 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X496 a_3947_12393# a_3597_12021# a_3852_12381# VPWR.t3021 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X497 a_5997_11247# mask\[5\] VGND.t2467 VGND.t2466 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X498 VGND.t3124 _114_ a_13393_1707# VGND.t3123 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X499 VGND.t410 _055_ a_15299_3311# VGND.t409 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X500 VGND.t2860 _113_ a_13183_3311# VGND.t2859 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X501 VPWR.t1345 _104_ a_10781_3311# VPWR.t1344 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X502 VPWR.t949 trim_val\[0\] a_15054_5193# VPWR.t948 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X503 a_4871_8181# net44 VPWR.t2853 VPWR.t2852 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X504 _034_ a_4167_6575# VGND.t3187 VGND.t3186 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X505 VGND.t1497 VPWR.t3365 VGND.t1496 VGND.t1495 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X506 VGND.t2820 _092_ a_4498_4373# VGND.t2819 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.123 ps=1.03 w=0.65 l=0.15
X507 VPWR.t2318 _048_.t19 a_5536_4399# VPWR.t2317 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.195 ps=1.39 w=1 l=0.15
X508 VPWR.t109 VGND.t3290 VPWR.t108 VPWR.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X509 a_9719_1473# _110_.t2 VPWR.t2164 VPWR.t2163 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X510 VPWR.t837 a_1129_4373# a_1019_4399# VPWR.t836 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X511 VPWR.t112 VGND.t3291 VPWR.t111 VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X512 VGND.t3050 _078_ a_1763_9295# VGND.t3049 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X513 ctln[7].t3 a_5363_591# VPWR.t1873 VPWR.t1872 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X514 VPWR.t2105 clknet_2_1__leaf_clk.t34 a_579_12021# VPWR.t2104 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X515 VPWR.t115 VGND.t3292 VPWR.t114 VPWR.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X516 _063_.t0 cal_itt\[1\] VPWR.t1638 VPWR.t1637 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.37 ps=1.74 w=1 l=0.15
X517 a_5524_9295# a_4609_9295# a_5177_9537# VGND.t261 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X518 a_1229_8457# _074_ VPWR.t888 VPWR.t887 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X519 _099_ _098_ a_6197_4399# VPWR.t1033 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X520 VPWR.t118 VGND.t3293 VPWR.t117 VPWR.t116 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X521 VGND.t1494 VPWR.t3366 VGND.t1493 VGND.t931 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X522 mask\[4\] a_9195_10357# VGND.t2764 VGND.t2763 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X523 VGND.t1652 a_9471_9269# a_9405_9295# VGND.t1651 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X524 VPWR.t121 VGND.t3294 VPWR.t120 VPWR.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X525 VPWR.t2271 a_6927_12559# ctlp[6].t3 VPWR.t2270 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X526 a_9595_5193# _063_.t10 _064_ VPWR.t2171 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X527 VPWR.t2708 a_13881_2741# _112_ VPWR.t2707 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X528 VPWR.t1794 a_7916_8041# a_8091_7967# VPWR.t1793 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X529 a_6515_6794# _073_ VPWR.t2549 VPWR.t2548 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X530 a_11601_2229# a_11435_2229# VPWR.t1753 VPWR.t1752 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X531 VPWR.t124 VGND.t3295 VPWR.t123 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X532 VPWR.t1489 a_14471_12559# ctlp[2].t1 VPWR.t1488 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X533 cal_itt\[0\] a_9471_9269# VPWR.t1672 VPWR.t1671 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.301 ps=2.66 w=1 l=0.15
X534 a_11023_5108# _108_ VGND.t775 VGND.t774 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X535 VGND.t333 clknet_0_clk a_8298_5487# VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X536 VGND.t3218 a_3667_3829# _048_.t11 VGND.t3217 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X537 trimb[3].t7 a_15023_12559# VGND.t2348 VGND.t2158 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X538 VPWR.t3189 mask\[2\] a_2689_8751# VPWR.t3188 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X539 VGND.t785 a_4043_7093# a_3977_7119# VGND.t784 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X540 VPWR.t2253 _062_.t9 a_10245_5193# VPWR.t2252 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X541 trim_mask\[3\] a_9747_2527# VGND.t404 VGND.t403 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X542 a_4512_12393# a_3431_12021# a_4165_11989# VPWR.t1174 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X543 result[6].t3 a_455_12533# VPWR.t2479 VPWR.t2478 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X544 VGND.t1492 VPWR.t3367 VGND.t1491 VGND.t1490 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X545 a_8745_4943# _053_ a_8307_4943# VGND.t2569 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X546 VGND.t1762 clknet_2_0__leaf_clk a_2787_7119# VGND.t1761 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X547 a_5177_1921# a_4959_1679# VGND.t2755 VGND.t2754 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X548 VPWR.t1354 a_3521_9813# a_3411_9839# VPWR.t1353 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X549 a_8820_12533# net19 VGND.t3136 VGND.t3135 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X550 a_4043_12393# a_3597_12021# a_3947_12393# VGND.t2968 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X551 a_4209_11293# a_4165_10901# a_4043_11305# VGND.t1611 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X552 VGND.t1489 VPWR.t3368 VGND.t1488 VGND.t1487 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X553 VGND.t3048 _078_ a_1211_7983# VGND.t3047 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X554 VGND.t2910 cal_itt\[3\] a_8307_6575# VGND.t2909 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X555 VPWR.t127 VGND.t3296 VPWR.t126 VPWR.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X556 VPWR.t3114 _078_ a_6007_9839# VPWR.t3113 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X557 VPWR.t2766 net13 a_5363_591# VPWR.t2765 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X558 VPWR.t2774 a_1651_7093# a_1638_7485# VPWR.t2773 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X559 a_929_8757# a_763_8757# VGND.t84 VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X560 clknet_0_clk a_8022_7119# VPWR.t1597 VPWR.t1596 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X561 a_8749_3317# a_8583_3317# VPWR.t2689 VPWR.t2688 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X562 a_10752_12533# net18 VGND.t93 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X563 net47 a_9463_8725# VPWR.t1547 VPWR.t1546 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X564 trim[4].t2 a_15023_5487# VPWR.t1233 VPWR.t1232 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X565 a_561_6031# a_395_6031# VPWR.t1300 VPWR.t1299 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X566 VGND.t2167 a_455_3571# valid.t6 VGND.t2166 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X567 VPWR.t130 VGND.t3297 VPWR.t129 VPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X568 VPWR.t132 VGND.t3298 VPWR.t131 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X569 a_4815_3031# state\[2\] VPWR.t1989 VPWR.t1988 sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X570 a_9084_4515# _106_ VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X571 a_7256_8029# _002_ VPWR.t1727 VPWR.t1726 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X572 VPWR.t2736 a_15023_1135# trim[3].t2 VPWR.t2735 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X573 VPWR.t135 VGND.t3299 VPWR.t134 VPWR.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X574 VPWR.t1562 _129_ a_14485_7663# VPWR.t1561 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.105 ps=1.21 w=1 l=0.15
X575 VPWR.t138 VGND.t3300 VPWR.t137 VPWR.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X576 net39 net34.t3 VPWR.t3072 VPWR.t3071 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X577 VPWR.t2388 _065_.t7 a_5363_7369# VPWR.t2387 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X578 a_3947_12393# a_3431_12021# a_3852_12381# VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X579 a_8022_7119# clk.t0 VPWR.t3157 VPWR.t3156 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X580 a_14686_3017# trim_mask\[1\] a_14604_3017# VPWR.t870 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X581 VGND.t1486 VPWR.t3369 VGND.t1485 VGND.t1484 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X582 a_2143_7663# _101_ a_2225_7663# VPWR.t1554 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X583 VPWR.t1987 state\[2\] a_7019_4407# VPWR.t1986 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X584 a_11374_1251# trim_mask\[3\] a_11292_1251# VPWR.t2100 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X585 a_1125_7663# net23 _080_ VPWR.t1653 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X586 VGND.t42 net48 a_14184_1679# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X587 VGND.t1960 state\[2\] a_5691_2741# VGND.t1959 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X588 VPWR.t1166 a_14063_7093# _134_ VPWR.t1165 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X589 a_2659_2601# a_2143_2229# a_2564_2589# VGND.t2352 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X590 VPWR.t141 VGND.t3301 VPWR.t140 VPWR.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X591 VPWR.t1871 a_5363_591# ctln[7].t2 VPWR.t1870 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X592 net55 a_7019_4407# VPWR.t3281 VPWR.t3280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X593 VPWR.t1704 net47 a_11244_9661# VPWR.t1703 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X594 a_2971_8457# _101_ a_3053_8457# VPWR.t1553 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X595 VGND.t1483 VPWR.t3370 VGND.t1482 VGND.t1481 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X596 a_5524_1679# a_4609_1679# a_5177_1921# VGND.t2869 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X597 a_1493_5487# _078_ VPWR.t3112 VPWR.t3111 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X598 VGND.t446 _084_ _009_ VGND.t445 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X599 VGND.t3034 a_5423_9011# _074_ VGND.t3033 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X600 clknet_2_2__leaf_clk a_8298_2767# VPWR.t2463 VPWR.t2462 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X601 VPWR.t144 VGND.t3302 VPWR.t143 VPWR.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X602 VPWR.t147 VGND.t3303 VPWR.t146 VPWR.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X603 VGND.t1480 VPWR.t3371 VGND.t1479 VGND.t908 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X604 VPWR.t150 VGND.t3304 VPWR.t149 VPWR.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X605 _102_ net52 VGND.t2398 VGND.t2397 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X606 a_4674_10927# a_3597_10933# a_4512_11305# VPWR.t2054 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X607 VGND.t1478 VPWR.t3372 VGND.t1477 VGND.t1476 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X608 _131_ cal_count\[2\] VPWR.t2216 VPWR.t2215 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X609 ctln[1].t1 a_3063_591# VPWR.t779 VPWR.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X610 VGND.t1475 VPWR.t3373 VGND.t1474 VGND.t1473 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X611 VPWR.t2647 cal_count\[3\] a_13111_6031# VPWR.t2646 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X612 net33 a_15023_1679# VPWR.t2074 VPWR.t2073 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X613 a_7460_5807# _048_.t20 VGND.t2287 VGND.t2286 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X614 _099_ _087_ VGND.t116 VGND.t115 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X615 VPWR.t3196 a_4165_11989# a_4055_12015# VPWR.t3195 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X616 a_10851_1653# a_10676_1679# a_11030_1679# VGND.t2768 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X617 VPWR.t1840 a_10569_1109# _116_ VPWR.t1839 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X618 a_5536_4399# _059_ a_5445_4399# VPWR.t1730 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.153 ps=1.3 w=1 l=0.15
X619 a_6999_12015# net44 VPWR.t2851 VPWR.t2850 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X620 a_11141_6031# a_10975_6031# VPWR.t2210 VPWR.t2209 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X621 VGND.t2430 a_8298_2767# clknet_2_2__leaf_clk VGND.t2429 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X622 VGND.t249 net46 a_9269_2589# VGND.t248 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X623 _046_ a_2828_12131# VGND.t2222 VGND.t2221 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X624 VPWR.t2811 a_1476_6031# a_1651_6005# VPWR.t2810 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X625 VGND.t2902 a_4498_4373# _093_ VGND.t2901 sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X626 VPWR.t153 VGND.t3305 VPWR.t152 VPWR.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X627 VGND.t2031 a_12631_12559# ctlp[3].t3 VGND.t2030 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X628 net26 a_7723_10143# VPWR.t2553 VPWR.t2552 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X629 a_4680_6031# _034_ VGND.t2436 VGND.t2435 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X630 VPWR.t1496 calibrate a_6927_3311# VPWR.t1495 sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.185 ps=1.37 w=1 l=0.15
X631 VGND.t1472 VPWR.t3374 VGND.t1471 VGND.t1470 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X632 a_9074_9955# net26 a_8992_9955# VPWR.t900 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X633 a_937_4105# calibrate VPWR.t1494 VPWR.t1493 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X634 _050_ a_5691_2741# VPWR.t2585 VPWR.t2584 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X635 a_1764_10383# mask\[7\] a_1461_10357# VGND.t2973 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X636 _122_ a_11016_6691# VGND.t124 VGND.t123 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X637 valid.t5 a_455_3571# VGND.t2165 VGND.t2164 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X638 VGND.t1469 VPWR.t3375 VGND.t1468 VGND.t1415 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X639 a_7477_10901# a_7259_11305# VPWR.t2314 VPWR.t2313 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X640 VGND.t2735 a_1651_7093# a_1585_7119# VGND.t2734 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X641 a_13783_6183# _135_ a_14181_6031# VGND.t2678 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X642 VGND.t3071 a_12612_8725# a_12546_9129# VGND.t3070 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X643 trim[3].t1 a_15023_1135# VPWR.t2734 VPWR.t2733 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X644 _000_ _068_ VPWR.t2251 VPWR.t2250 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X645 clknet_2_3__leaf_clk a_8298_5487# VGND.t2128 VGND.t2127 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X646 a_13279_8207# cal_count\[1\] VGND.t2175 VGND.t2174 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X647 a_7001_7669# a_6835_7669# VPWR.t791 VPWR.t790 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X648 a_1173_7119# a_1129_7361# a_1007_7119# VGND.t531 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X649 _056_ a_14604_2339# VGND.t1771 VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X650 VPWR.t156 VGND.t3306 VPWR.t155 VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X651 _107_ a_5536_4399# VGND.t537 VGND.t536 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X652 trimb[2].t6 a_15023_12015# VGND.t2157 VGND.t2156 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X653 a_12612_8725# net47 VPWR.t1702 VPWR.t1701 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X654 a_6927_3311# _104_ a_7010_3311# VPWR.t1343 sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.14 ps=1.28 w=1 l=0.15
X655 VGND.t678 a_2857_5461# clknet_2_0__leaf_clk VGND.t677 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X656 a_1644_12533# net29 VPWR.t2902 VPWR.t2901 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X657 VPWR.t1106 a_2857_7637# clknet_2_1__leaf_clk.t12 VPWR.t1105 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X658 VGND.t46 a_13142_8359# _036_ VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X659 VGND.t1467 VPWR.t3376 VGND.t1466 VGND.t1465 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X660 VGND.t1464 VPWR.t3377 VGND.t1463 VGND.t1462 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X661 a_14236_8457# cal_count\[1\] VGND.t2173 VGND.t2172 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X662 VGND.t1828 net53 a_6261_11247# VGND.t1827 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X663 a_8455_10383# a_8105_10383# a_8360_10383# VPWR.t2880 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X664 a_2857_7637# clknet_0_clk VGND.t331 VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X665 a_10688_9295# a_10239_9295# a_10593_9295# VGND.t3016 sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X666 VPWR.t1857 a_13142_8725# a_13100_8751# VPWR.t1856 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X667 a_14347_1439# a_14172_1513# a_14526_1501# VGND.t3078 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X668 VPWR.t2461 a_8298_2767# clknet_2_2__leaf_clk VPWR.t2460 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X669 _092_ a_10005_6031# VGND.t67 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X670 a_5931_4105# _087_ VPWR.t856 VPWR.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X671 VGND.t2098 a_4091_5309# _065_.t3 VGND.t2097 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X672 a_7250_7485# a_6173_7119# a_7088_7119# VPWR.t1566 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X673 a_11067_3017# _064_ a_11149_2767# VGND.t1608 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X674 a_3521_9813# a_3303_10217# VGND.t2914 VGND.t2913 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X675 a_11116_8983# _123_.t5 a_11258_9117# VGND.t1635 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X676 VGND.t2049 a_9460_6807# _068_ VGND.t2048 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X677 a_7256_8029# _002_ VGND.t1707 VGND.t1706 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X678 a_11016_6691# _065_.t8 VGND.t3230 VGND.t3229 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X679 a_9099_3689# a_8749_3317# a_9004_3677# VPWR.t2918 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X680 ctln[0].t0 a_1276_565# VPWR.t3088 VPWR.t3087 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X681 a_9662_3855# trim_val\[4\] a_9003_3829# VGND.t108 sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.104 ps=0.97 w=0.65 l=0.15
X682 net18 a_9871_10383# VGND.t555 VGND.t554 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X683 VGND.t73 _126_ a_14552_9071# VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X684 VPWR.t159 VGND.t3307 VPWR.t158 VPWR.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X685 a_6741_7361# a_6523_7119# VPWR.t2370 VPWR.t2369 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X686 a_10977_2543# _064_ a_10543_2455# VGND.t1607 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X687 VGND.t1461 VPWR.t3378 VGND.t1460 VGND.t1270 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X688 a_1201_3855# calibrate a_855_4105# VGND.t739 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X689 VGND.t2846 a_1651_6005# a_1585_6031# VGND.t2845 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X690 mask\[6\] a_4687_11231# VGND.t2458 VGND.t2457 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X691 _038_ a_10699_5487# VPWR.t1461 VPWR.t1460 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X692 _067_ trim_mask\[0\] a_10138_5807# VGND.t1875 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X693 a_1549_6794# _039_ VPWR.t3218 VPWR.t3217 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X694 a_3302_3677# net45 VGND.t2491 VGND.t2490 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X695 VPWR.t1818 _042_.t2 a_11803_10383# VPWR.t1817 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X696 mask\[0\] a_4043_7093# VGND.t783 VGND.t782 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X697 a_1173_6031# a_1129_6273# a_1007_6031# VGND.t3130 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X698 a_4905_3855# _096_ a_4471_4007# VGND.t307 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X699 VPWR.t162 VGND.t3308 VPWR.t161 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X700 VPWR.t2697 a_5699_1653# a_5686_2045# VPWR.t2696 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X701 VGND.t2023 a_15023_10927# trimb[0].t7 VGND.t2022 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X702 _123_.t2 _063_.t11 VPWR.t2173 VPWR.t2172 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X703 VGND.t286 clknet_2_2__leaf_clk a_8583_3317# VGND.t285 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X704 a_10781_3631# trim_mask\[2\] VGND.t2840 VGND.t2839 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X705 VPWR.t2269 a_6927_12559# ctlp[6].t2 VPWR.t2268 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X706 VPWR.t1074 clknet_0_clk a_2857_7637# VPWR.t1073 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X707 a_1019_7485# net43.t11 VPWR.t1382 VPWR.t1381 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X708 calibrate a_1651_4703# VPWR.t2979 VPWR.t2978 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X709 a_8301_8207# _072_ a_8083_8181# VGND.t2758 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X710 VGND.t2614 a_15259_7637# net2 VGND.t2613 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X711 VGND.t2992 mask\[0\] a_2313_6183# VGND.t2991 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X712 VPWR.t165 VGND.t3309 VPWR.t164 VPWR.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X713 a_9020_10383# a_7939_10383# a_8673_10625# VPWR.t944 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X714 clknet_0_clk a_8022_7119# VPWR.t1595 VPWR.t1594 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X715 _060_ a_4576_3427# VGND.t464 VGND.t463 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X716 VPWR.t3068 a_10383_7093# cal_itt\[1\] VPWR.t3067 sky130_fd_pr__pfet_01v8_hvt ad=0.301 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X717 a_2921_2589# a_2877_2197# a_2755_2601# VGND.t187 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X718 VGND.t2126 a_8298_5487# clknet_2_3__leaf_clk VGND.t2125 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X719 _042_.t1 a_2368_9955# VGND.t2518 VGND.t2517 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X720 VGND.t1459 VPWR.t3379 VGND.t1458 VGND.t1457 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X721 a_7190_3855# _049_ a_7104_3855# VGND.t457 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X722 ctlp[2].t0 a_14471_12559# VPWR.t1487 VPWR.t1486 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X723 a_6999_12015# a_6375_12021# a_6891_12393# VPWR.t3062 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X724 a_1276_565# net6 VPWR.t1744 VPWR.t1743 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X725 trimb[3].t6 a_15023_12559# VGND.t2347 VGND.t2156 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X726 VPWR.t168 VGND.t3310 VPWR.t167 VPWR.t166 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X727 VPWR.t1700 net47 a_11204_7485# VPWR.t1699 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.109 ps=1.36 w=0.42 l=0.15
X728 VPWR.t171 VGND.t3311 VPWR.t170 VPWR.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X729 a_9207_3311# a_8583_3317# a_9099_3689# VPWR.t2687 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X730 a_8495_6895# a_8307_6575# _063_.t5 VGND.t2313 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X731 VGND.t2208 _044_ a_8767_11471# VGND.t2207 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X732 result[6].t2 a_455_12533# VPWR.t2477 VPWR.t2476 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X733 VPWR.t3004 a_10752_565# ctln[4].t1 VPWR.t3003 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X734 VGND.t2996 net4.t2 a_10055_2767# VGND.t2995 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X735 a_13050_7637# a_12900_7663# VPWR.t3228 VPWR.t3227 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X736 a_12424_3689# a_11509_3317# a_12077_3285# VGND.t2256 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X737 VPWR.t1824 a_11545_9049# a_11575_8790# VPWR.t1823 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X738 VGND.t1456 VPWR.t3380 VGND.t1455 VGND.t1454 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X739 VPWR.t174 VGND.t3312 VPWR.t173 VPWR.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X740 a_15159_9269# _125_ VPWR.t2043 VPWR.t2042 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X741 a_6007_9839# mask\[4\] VPWR.t2683 VPWR.t2682 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X742 a_9115_2223# net46 VPWR.t993 VPWR.t992 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X743 a_3057_4719# _092_ VGND.t2818 VGND.t2817 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X744 VPWR.t177 VGND.t3313 VPWR.t176 VPWR.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X745 a_9677_8457# _070_ _001_ VPWR.t2001 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X746 VPWR.t180 VGND.t3314 VPWR.t179 VPWR.t178 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X747 VPWR.t2983 a_9020_10383# a_9195_10357# VPWR.t2982 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X748 VPWR.t1875 a_10655_2932# _033_ VPWR.t1874 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X749 VPWR.t2312 a_6741_7361# a_6631_7485# VPWR.t2311 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X750 a_1476_6031# a_395_6031# a_1129_6273# VPWR.t1298 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X751 net8 net16 VGND.t201 VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X752 a_3521_7361# a_3303_7119# VPWR.t1509 VPWR.t1508 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X753 a_2309_2229# a_2143_2229# VGND.t2351 VGND.t2350 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X754 VPWR.t1917 clknet_2_3__leaf_clk a_8215_9295# VPWR.t1916 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X755 a_12436_9129# a_12153_8757# a_12341_8751# VPWR.t1238 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X756 VGND.t509 a_3933_2767# _051_.t10 VGND.t508 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X757 VGND.t2692 a_15023_1135# trim[3].t7 VGND.t2691 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X758 mask\[2\] a_4043_10143# VPWR.t2792 VPWR.t2791 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X759 clknet_2_1__leaf_clk.t11 a_2857_7637# VPWR.t1104 VPWR.t1103 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X760 VGND.t1453 VPWR.t3381 VGND.t1452 VGND.t1451 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X761 a_9471_9269# a_9296_9295# a_9650_9295# VGND.t769 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X762 a_5423_9011# _065_.t9 VPWR.t3311 VPWR.t3310 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X763 a_1579_5807# mask\[0\] _079_ VGND.t2990 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X764 a_13557_7369# _122_ a_13142_7271# VPWR.t2095 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X765 VGND.t247 net46 a_14237_3677# VGND.t246 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X766 VPWR.t3303 a_12599_3615# a_12586_3311# VPWR.t3302 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X767 a_13519_4007# _112_ VPWR.t1746 VPWR.t1745 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X768 a_12310_4399# a_11233_4405# a_12148_4777# VPWR.t1879 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X769 a_816_7119# _005_ VGND.t2929 VGND.t2928 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X770 a_8298_2767# clknet_0_clk VPWR.t1072 VPWR.t1071 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X771 VGND.t390 net51 _101_ VGND.t389 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X772 a_2948_3689# a_2033_3317# a_2601_3285# VGND.t754 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X773 a_13519_4007# _110_.t3 a_13693_3883# VGND.t2137 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X774 a_10621_7119# a_10586_7371# a_10383_7093# VGND.t570 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X775 a_11297_7119# net47 VGND.t1685 VGND.t1684 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.135 ps=1.15 w=0.42 l=0.15
X776 clkc.t0 a_15299_6575# VPWR.t1660 VPWR.t1659 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X777 a_9317_3285# a_9099_3689# VGND.t2610 VGND.t2609 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X778 a_7379_2197# a_7223_2465# a_7524_2223# VPWR.t2402 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.116 ps=0.97 w=0.42 l=0.15
X779 VPWR.t2619 _050_ _062_.t7 VPWR.t2618 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X780 a_14099_1929# trim_val\[2\] a_13881_1653# VPWR.t2678 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X781 _045_ a_5496_12131# VPWR.t1609 VPWR.t1608 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X782 a_1677_9545# net25 _082_ VPWR.t3132 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X783 a_9296_9295# a_8215_9295# a_8949_9537# VPWR.t1963 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X784 VGND.t2597 a_5691_7637# net52 VGND.t2596 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X785 VPWR.t1543 a_13111_6031# _135_ VPWR.t1542 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X786 VPWR.t183 VGND.t3315 VPWR.t182 VPWR.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X787 VPWR.t1070 clknet_0_clk a_2857_5461# VPWR.t1069 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X788 VPWR.t186 VGND.t3316 VPWR.t185 VPWR.t184 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X789 VGND.t1450 VPWR.t3382 VGND.t1449 VGND.t1448 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X790 VPWR.t2302 a_10752_12533# ctlp[4].t0 VPWR.t2301 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X791 _106_ a_8307_4943# VGND.t497 VGND.t496 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102 ps=0.965 w=0.65 l=0.15
X792 a_1173_10205# a_1129_9813# a_1007_10217# VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X793 a_12231_6005# net46 VPWR.t991 VPWR.t990 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X794 VGND.t2955 a_8820_6005# _071_ VGND.t2954 sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X795 a_9595_5193# _062_.t10 VPWR.t2235 VPWR.t2234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X796 _093_ a_4498_4373# VPWR.t2947 VPWR.t2946 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X797 a_911_10217# a_561_9845# a_816_10205# VPWR.t3181 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X798 a_13142_7271# _133_ a_13279_7119# VGND.t3101 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X799 a_6737_3855# _052_ VGND.t382 VGND.t381 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X800 VPWR.t2912 a_5340_6031# a_5515_6005# VPWR.t2911 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X801 VGND.t630 net43.t12 a_4209_12381# VGND.t629 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X802 ctlp[3].t2 a_12631_12559# VGND.t2029 VGND.t2028 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X803 a_6515_6794# _073_ VGND.t2512 VGND.t2511 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X804 ctln[2].t2 a_14471_591# VGND.t686 VGND.t685 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X805 a_3513_12809# _085_ _010_ VPWR.t2038 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X806 VPWR.t809 a_10005_6031# _092_ VPWR.t808 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X807 _062_.t3 a_7262_5461# VPWR.t1613 VPWR.t1612 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X808 a_8298_5487# clknet_0_clk VGND.t329 VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X809 a_816_6031# _004_ VGND.t1613 VGND.t1612 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X810 VGND.t1447 VPWR.t3383 VGND.t1446 VGND.t1445 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X811 a_9225_2197# a_9007_2601# VPWR.t2404 VPWR.t2403 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X812 VGND.t1805 clknet_2_1__leaf_clk.t35 a_579_10933# VGND.t1804 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X813 _028_ a_7010_3311# VPWR.t2485 VPWR.t2484 sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.243 ps=1.49 w=1 l=0.15
X814 VPWR.t189 VGND.t3317 VPWR.t188 VPWR.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X815 a_7942_2223# a_7184_2339# a_7379_2197# VPWR.t2742 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0724 ps=0.765 w=0.42 l=0.15
X816 a_3597_10933# a_3431_10933# VPWR.t1666 VPWR.t1665 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X817 VGND.t3020 _131_ a_15289_7119# VGND.t3019 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X818 VPWR.t2986 _130_ a_14199_7369# VPWR.t2985 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X819 VPWR.t2332 a_7715_3285# _052_ VPWR.t2331 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X820 a_1099_12533# net14 VGND.t1932 VGND.t1931 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X821 a_4055_12015# a_3431_12021# a_3947_12393# VPWR.t1173 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X822 a_2961_9545# net52 VPWR.t2429 VPWR.t2428 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X823 VPWR.t2996 cal_count\[0\] a_14377_9545# VPWR.t2995 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X824 VPWR.t192 VGND.t3318 VPWR.t191 VPWR.t190 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X825 VPWR.t1593 a_8022_7119# clknet_0_clk VPWR.t1592 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X826 _133_ a_14335_7895# VPWR.t2998 VPWR.t2997 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.36 ps=2.72 w=1 l=0.15
X827 VPWR.t1231 a_15023_5487# trim[4].t1 VPWR.t1230 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X828 a_11753_6031# a_11709_6273# a_11587_6031# VGND.t1818 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X829 VPWR.t1718 a_12631_591# ctln[3].t1 VPWR.t1717 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X830 a_11057_4105# trim_mask\[0\] VPWR.t1902 VPWR.t1901 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X831 net29 a_1835_12319# VPWR.t2649 VPWR.t2648 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X832 a_8455_10383# a_7939_10383# a_8360_10383# VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X833 VPWR.t1826 clknet_2_1__leaf_clk.t36 a_395_9845# VPWR.t1825 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X834 a_12625_2601# a_11435_2229# a_12516_2601# VGND.t1738 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X835 VGND.t1850 a_10655_2932# _033_ VGND.t597 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X836 a_2033_3317# a_1867_3317# VPWR.t1946 VPWR.t1945 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X837 VGND.t2554 _132_ a_14377_7983# VGND.t2553 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X838 VGND.t107 trim_val\[4\] a_10188_4105# VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X839 VPWR.t2151 a_8298_5487# clknet_2_3__leaf_clk VPWR.t2150 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X840 a_13356_8457# _128_ VPWR.t3000 VPWR.t2999 sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X841 a_7617_2589# net45 VGND.t2489 VGND.t2488 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.135 ps=1.15 w=0.42 l=0.15
X842 net42 a_7571_4943# VPWR.t2916 VPWR.t2915 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X843 a_4222_10205# net43.t13 VGND.t632 VGND.t631 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X844 a_4858_8573# a_3781_8207# a_4696_8207# VPWR.t1792 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X845 VPWR.t2392 a_8767_591# ctln[5].t1 VPWR.t2391 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X846 a_4687_11231# a_4512_11305# a_4866_11293# VGND.t693 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X847 VGND.t1444 VPWR.t3384 VGND.t1443 VGND.t1442 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X848 net35 a_14655_4399# VPWR.t1314 VPWR.t1313 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X849 VPWR.t195 VGND.t3319 VPWR.t194 VPWR.t193 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X850 VGND.t2779 net17 net9 VGND.t2778 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X851 a_12454_8041# a_12061_7669# a_12344_8041# VGND.t1951 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X852 VGND.t773 _108_ a_14000_4719# VGND.t772 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X853 a_4709_2773# state\[1\] VPWR.t3126 VPWR.t3125 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X854 a_2019_9055# net43.t14 VPWR.t2746 VPWR.t2745 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X855 VPWR.t1800 mask\[1\] a_1125_7663# VPWR.t1799 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X856 a_9572_2601# a_8491_2229# a_9225_2197# VPWR.t2361 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X857 a_8761_7983# _071_ VGND.t2976 VGND.t2975 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X858 VPWR.t819 net31 net36 VPWR.t818 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X859 _006_ _074_ VGND.t151 VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X860 VGND.t1441 VPWR.t3385 VGND.t1440 VGND.t1439 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X861 a_3303_7119# a_2953_7119# a_3208_7119# VPWR.t2003 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X862 a_11396_6031# _038_ VGND.t1639 VGND.t1638 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X863 VPWR.t3159 a_12169_2197# a_12059_2223# VPWR.t3158 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X864 clknet_0_clk a_8022_7119# VGND.t845 VGND.t844 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X865 VGND.t3014 a_5515_6005# a_5449_6031# VGND.t3013 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X866 VPWR.t787 a_10195_1354# _032_ VPWR.t786 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X867 VGND.t2749 a_4043_10143# a_3977_10217# VGND.t2748 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X868 a_8949_9537# a_8731_9295# VPWR.t1820 VPWR.t1819 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X869 a_7379_2197# a_7184_2339# a_7689_2589# VGND.t2695 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.14 ps=1.1 w=0.36 l=0.15
X870 clknet_2_0__leaf_clk a_2857_5461# VPWR.t1434 VPWR.t1433 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X871 a_5037_6031# a_4993_6273# a_4871_6031# VGND.t3206 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X872 VGND.t1893 clknet_2_3__leaf_clk a_11987_8757# VGND.t1892 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X873 VGND.t731 a_5535_8181# _078_ VGND.t730 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X874 VGND.t2545 a_5691_2741# _050_ VGND.t2544 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X875 VGND.t1760 clknet_2_0__leaf_clk a_395_4405# VGND.t1759 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X876 net16 a_13919_8751# VPWR.t3146 VPWR.t3145 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X877 VPWR.t1738 a_6519_4631# _100_ VPWR.t1737 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X878 a_455_5747# net30.t6 VGND.t28 VGND.t27 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X879 VGND.t2800 net44 a_4393_8207# VGND.t2799 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X880 a_11045_5807# cal_count\[3\] a_10699_5487# VGND.t2604 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X881 VPWR.t1953 a_6885_8372# net51 VPWR.t1952 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X882 VGND.t2900 a_4498_4373# _093_ VGND.t2899 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X883 a_3852_11293# _022_ VPWR.t896 VPWR.t895 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X884 VPWR.t198 VGND.t3320 VPWR.t197 VPWR.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X885 VGND.t1438 VPWR.t3386 VGND.t1437 VGND.t1220 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X886 VGND.t1969 net50 a_10872_1455# VGND.t1968 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X887 _050_ a_5691_2741# VPWR.t2583 VPWR.t2582 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X888 VGND.t705 state\[0\] a_3667_3829# VGND.t704 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X889 clknet_2_2__leaf_clk a_8298_2767# VGND.t2428 VGND.t2427 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X890 VGND.t1436 VPWR.t3387 VGND.t1435 VGND.t1262 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X891 a_911_7119# a_395_7119# a_816_7119# VGND.t1796 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X892 a_11321_3855# trim_mask\[0\] a_10975_4105# VGND.t1874 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X893 VGND.t149 _074_ _005_ VGND.t148 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X894 VPWR.t902 a_12231_6005# a_12218_6397# VPWR.t901 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X895 VPWR.t845 a_3116_12533# ctlp[1].t1 VPWR.t844 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X896 a_3053_8457# mask\[2\] VPWR.t3187 VPWR.t3186 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X897 VPWR.t2021 a_2601_3285# a_2491_3311# VPWR.t2020 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X898 a_8078_7663# a_7001_7669# a_7916_8041# VPWR.t1452 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X899 VPWR.t201 VGND.t3321 VPWR.t200 VPWR.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X900 VGND.t1434 VPWR.t3388 VGND.t1433 VGND.t1432 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X901 a_8473_5193# net55 a_8389_5193# VPWR.t3017 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X902 VPWR.t2882 a_14540_3689# a_14715_3615# VPWR.t2881 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X903 trim[4].t0 a_15023_5487# VPWR.t1229 VPWR.t1228 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X904 VGND.t2163 a_455_3571# valid.t4 VGND.t2162 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X905 a_3411_7485# a_2787_7119# a_3303_7119# VPWR.t2875 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X906 VGND.t1431 VPWR.t3389 VGND.t1430 VGND.t1429 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X907 VGND.t1711 _059_ net41 VGND.t1710 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X908 VPWR.t204 VGND.t3322 VPWR.t203 VPWR.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X909 a_1203_10927# a_579_10933# a_1095_11305# VPWR.t1334 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X910 a_13059_4631# _110_.t4 VPWR.t2166 VPWR.t2165 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X911 VGND.t1428 VPWR.t3390 VGND.t1427 VGND.t1321 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X912 VPWR.t841 a_1129_9813# a_1019_9839# VPWR.t840 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X913 VGND.t1634 net23 a_2092_8457# VGND.t1633 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X914 state\[1\] a_3399_2527# VGND.t517 VGND.t516 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X915 VGND.t456 _049_ _076_ VGND.t455 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X916 VGND.t2699 net43.t15 a_1173_10205# VGND.t2698 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X917 VGND.t2701 net43.t16 a_1541_9117# VGND.t2700 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X918 a_3847_4438# _090_ a_3388_4631# VPWR.t1136 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X919 VGND.t1426 VPWR.t3391 VGND.t1425 VGND.t1424 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X920 a_2019_9055# a_1844_9129# a_2198_9117# VGND.t2263 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X921 VGND.t122 a_4815_3031# _053_ VGND.t121 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X922 clknet_2_0__leaf_clk a_2857_5461# VGND.t676 VGND.t675 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X923 VPWR.t2500 mask\[5\] a_8154_11721# VPWR.t2499 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X924 a_5998_11471# _078_ VGND.t3046 VGND.t3045 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X925 VGND.t1423 VPWR.t3392 VGND.t1422 VGND.t1421 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X926 a_5931_4105# _089_ _090_ VPWR.t1750 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X927 VGND.t1420 VPWR.t3393 VGND.t1419 VGND.t1418 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X928 a_937_3855# net1 VGND.t1986 VGND.t1985 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X929 _048_.t4 a_3667_3829# VPWR.t3297 VPWR.t3296 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X930 VPWR.t207 VGND.t3323 VPWR.t206 VPWR.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X931 VGND.t1417 VPWR.t3394 VGND.t1416 VGND.t1415 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X932 a_911_6031# a_395_6031# a_816_6031# VGND.t559 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X933 _098_ _050_ VGND.t2581 VGND.t2580 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X934 clknet_2_2__leaf_clk a_8298_2767# VPWR.t2459 VPWR.t2458 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X935 VGND.t1414 VPWR.t3395 VGND.t1413 VGND.t1412 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X936 a_10747_8970# _124_ VPWR.t1444 VPWR.t1443 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X937 net42 a_7571_4943# VGND.t2871 VGND.t2870 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X938 _091_ a_9443_6059# VGND.t768 VGND.t767 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X939 VPWR.t2380 a_15023_12559# trimb[3].t3 VPWR.t2379 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X940 VPWR.t209 VGND.t3324 VPWR.t208 VPWR.t196 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X941 a_3057_3689# a_1867_3317# a_2948_3689# VGND.t1920 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X942 a_9802_4007# _108_ VGND.t771 VGND.t770 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.109 ps=0.985 w=0.65 l=0.15
X943 VGND.t1411 VPWR.t3396 VGND.t1410 VGND.t1409 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X944 VPWR.t886 _074_ a_3513_12809# VPWR.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X945 a_4901_2773# a_4709_2773# a_4815_3031# VGND.t3061 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X946 VPWR.t2052 a_6519_3829# _089_ VPWR.t1737 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X947 VPWR.t212 VGND.t3325 VPWR.t211 VPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X948 a_6906_2355# a_7184_2339# a_7140_2223# VPWR.t2741 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X949 VGND.t596 _104_ a_11413_2767# VGND.t595 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X950 VPWR.t1623 _064_ a_10055_5487# VPWR.t1622 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X951 clknet_2_1__leaf_clk.t28 a_2857_7637# VGND.t369 VGND.t368 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X952 VPWR.t1863 _134_ a_13933_6281# VPWR.t1862 sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.105 ps=1.21 w=1 l=0.15
X953 VGND.t2426 a_8298_2767# clknet_2_2__leaf_clk VGND.t2425 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X954 VPWR.t215 VGND.t3326 VPWR.t214 VPWR.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X955 a_455_3571# net41 VPWR.t2336 VPWR.t2335 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X956 VGND.t2373 _066_ _067_ VGND.t2372 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X957 VPWR.t218 VGND.t3327 VPWR.t217 VPWR.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X958 VGND.t1798 _042_.t3 a_11803_10383# VGND.t1797 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X959 VGND.t1408 VPWR.t3397 VGND.t1407 VGND.t1406 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X960 a_12341_8751# _036_ VGND.t2684 VGND.t2683 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X961 a_1549_6794# _039_ VGND.t3142 VGND.t3141 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X962 VGND.t1807 clknet_2_1__leaf_clk.t37 a_6743_10933# VGND.t1806 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X963 a_7810_12381# net44 VGND.t2798 VGND.t2797 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X964 net13 net21 VGND.t2269 VGND.t2268 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X965 VGND.t1405 VPWR.t3398 VGND.t1404 VGND.t1403 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X966 a_13825_1109# a_13607_1513# VPWR.t1142 VPWR.t1141 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X967 VGND.t1402 VPWR.t3399 VGND.t1401 VGND.t1400 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X968 a_6261_11247# mask\[6\] a_5915_10927# VGND.t607 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X969 VPWR.t2205 a_4655_10071# _019_ VPWR.t2204 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X970 VPWR.t3283 a_7569_7637# a_7459_7663# VPWR.t3282 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X971 VGND.t2568 _053_ a_7190_3855# VGND.t2567 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X972 ctln[4].t0 a_10752_565# VPWR.t3002 VPWR.t3001 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X973 VGND.t515 a_3399_2527# a_3333_2601# VGND.t514 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X974 a_2479_3689# a_2033_3317# a_2383_3689# VGND.t753 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X975 net54 a_5087_3855# VPWR.t3332 VPWR.t3331 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X976 VPWR.t1865 _043_ a_9871_10383# VPWR.t1864 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X977 clknet_2_3__leaf_clk a_8298_5487# VGND.t2124 VGND.t2123 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X978 a_11491_6031# a_10975_6031# a_11396_6031# VGND.t2184 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X979 VGND.t612 a_7631_12319# a_7565_12393# VGND.t611 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X980 result[2].t7 a_455_8181# VGND.t2320 VGND.t1629 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X981 VGND.t1786 a_6927_591# ctln[6].t6 VGND.t1785 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X982 a_2659_2601# a_2309_2229# a_2564_2589# VPWR.t741 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X983 VPWR.t221 VGND.t3328 VPWR.t220 VPWR.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X984 _025_ a_10699_3311# VGND.t1903 VGND.t1902 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X985 VPWR.t224 VGND.t3329 VPWR.t223 VPWR.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X986 VPWR.t1102 a_2857_7637# clknet_2_1__leaf_clk.t10 VPWR.t1101 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X987 VGND.t1399 VPWR.t3400 VGND.t1398 VGND.t1397 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X988 a_3365_4943# _092_ VGND.t2816 VGND.t2815 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X989 VGND.t2045 a_5363_12559# ctlp[7].t7 VGND.t2044 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X990 VPWR.t1995 a_7824_11305# a_7999_11231# VPWR.t1994 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X991 a_10861_7119# a_10383_7093# VGND.t3010 VGND.t3009 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.125 ps=1.01 w=0.42 l=0.15
X992 VPWR.t3216 a_15023_2223# trim[2].t3 VPWR.t3215 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X993 VGND.t2731 a_448_6549# result[0].t3 VGND.t2730 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X994 a_9926_2589# net46 VGND.t245 VGND.t244 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X995 a_1000_11293# _023_ VGND.t2161 VGND.t2160 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X996 clknet_2_1__leaf_clk.t27 a_2857_7637# VGND.t367 VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X997 VPWR.t2427 net52 a_3053_8457# VPWR.t2426 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X998 a_4131_8207# a_3781_8207# a_4036_8207# VPWR.t1791 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X999 a_3208_10205# _018_ VPWR.t1607 VPWR.t1606 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1000 _083_ net26 a_6007_9839# VPWR.t899 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1001 a_11059_7356# a_10903_7261# a_11204_7485# VPWR.t1517 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.116 ps=0.97 w=0.42 l=0.15
X1002 VGND.t3090 _079_ _004_ VGND.t3089 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1003 VGND.t1396 VPWR.t3401 VGND.t1395 VGND.t1394 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1004 VGND.t495 a_15023_5487# trim[4].t7 VGND.t494 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1005 a_14172_1513# a_13091_1141# a_13825_1109# VPWR.t1276 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1006 VGND.t1683 net47 a_13164_8029# VGND.t1682 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
X1007 a_14335_7895# _132_ a_14733_7983# VGND.t2552 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X1008 a_4801_9839# _101_ a_4655_10071# VPWR.t1552 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X1009 en_co_clk a_5515_6005# VGND.t3012 VGND.t3011 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1010 VGND.t588 a_4863_4917# _095_ VGND.t587 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1011 a_10752_565# net10 VPWR.t1156 VPWR.t1155 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1012 VPWR.t227 VGND.t3330 VPWR.t226 VPWR.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1013 _119_ a_9003_3829# VGND.t427 VGND.t426 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1014 VPWR.t230 VGND.t3331 VPWR.t229 VPWR.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1015 trim[3].t6 a_15023_1135# VGND.t2690 VGND.t2689 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1016 VGND.t1681 net47 a_8993_9295# VGND.t1680 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1017 VPWR.t1322 a_6793_8970# net53 VPWR.t1321 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1018 net52 a_5691_7637# VPWR.t2637 VPWR.t2636 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1019 a_9460_6807# _067_ a_9602_6941# VGND.t186 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1020 clknet_2_2__leaf_clk a_8298_2767# VGND.t2424 VGND.t2423 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1021 a_3425_11721# _078_ VPWR.t3110 VPWR.t3109 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X1022 a_1129_6273# a_911_6031# VPWR.t1617 VPWR.t1616 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1023 a_7657_10217# a_6467_9845# a_7548_10217# VGND.t2456 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1024 VGND.t3113 net11 a_8767_591# VGND.t3112 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1025 clknet_0_clk a_8022_7119# VGND.t843 VGND.t842 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1026 a_2767_2223# a_2143_2229# a_2659_2601# VPWR.t2383 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1027 result[7].t3 a_1644_12533# VGND.t529 VGND.t528 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1028 a_14335_7895# _129_ VPWR.t1560 VPWR.t1559 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.365 ps=1.73 w=1 l=0.15
X1029 VPWR.t233 VGND.t3332 VPWR.t232 VPWR.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1030 VGND.t2595 a_5691_7637# net52 VGND.t2594 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1031 cal_itt\[3\] a_7263_7093# VPWR.t1969 VPWR.t1968 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1032 VPWR.t1025 clknet_2_2__leaf_clk a_11343_3317# VPWR.t1024 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1033 VPWR.t3016 net55 _059_ VPWR.t3015 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1034 net36 net31 VPWR.t817 VPWR.t816 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1035 a_4609_1679# a_4443_1679# VPWR.t1977 VPWR.t1976 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1036 VPWR.t1023 clknet_2_2__leaf_clk a_13091_4943# VPWR.t1022 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1037 clkc.t1 a_15299_6575# VGND.t1641 VGND.t1640 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1038 VGND.t1393 VPWR.t3402 VGND.t1392 VGND.t1391 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1039 a_11057_3855# trim_mask\[1\] VGND.t132 VGND.t131 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1040 a_14347_4917# a_14172_4943# a_14526_4943# VGND.t764 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1041 a_5054_4399# _090_ a_4970_4399# VPWR.t1135 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X1042 VPWR.t2162 mask\[3\] a_1677_9545# VPWR.t2161 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X1043 VPWR.t3208 net19 net11 VPWR.t3207 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1044 clknet_0_clk a_8022_7119# VPWR.t1591 VPWR.t1590 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1045 a_7088_7119# a_6173_7119# a_6741_7361# VGND.t807 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1046 a_11622_7485# a_10864_7387# a_11059_7356# VPWR.t951 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0724 ps=0.765 w=0.42 l=0.15
X1047 a_2857_5461# clknet_0_clk VPWR.t1068 VPWR.t1067 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1048 a_1467_7923# net45 VGND.t2487 VGND.t2486 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X1049 _093_ a_4498_4373# VPWR.t2945 VPWR.t2944 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1050 VGND.t1809 clknet_2_1__leaf_clk.t38 a_7939_10383# VGND.t1808 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1051 VPWR.t1265 a_1467_7923# net43.t3 VPWR.t1264 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1052 VPWR.t1150 a_10851_1653# a_10838_2045# VPWR.t1149 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1053 a_816_4765# _012_ VPWR.t2433 VPWR.t2432 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1054 net23 a_1651_7093# VGND.t2733 VGND.t2732 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1055 VGND.t1390 VPWR.t3403 VGND.t1389 VGND.t1388 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1056 VPWR.t1358 a_7631_12319# a_7618_12015# VPWR.t1357 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1057 VGND.t806 _129_ a_14377_7983# VGND.t805 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1058 a_1769_12393# a_579_12021# a_1660_12393# VGND.t569 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1059 VPWR.t913 trim_val\[1\] a_14686_3017# VPWR.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1060 _086_ net29 VGND.t2858 VGND.t2857 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1061 VPWR.t236 VGND.t3333 VPWR.t235 VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1062 a_13441_6281# cal_count\[3\] VPWR.t2645 VPWR.t2644 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X1063 a_3521_7361# a_3303_7119# VGND.t756 VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1064 trim[1].t3 a_15083_4659# VPWR.t2279 VPWR.t2278 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1065 ctlp[1].t0 a_3116_12533# VPWR.t843 VPWR.t842 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1066 net37.t1 net32 VPWR.t1216 VPWR.t1215 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1067 VPWR.t1306 _091_ a_10005_6031# VPWR.t1305 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1068 VPWR.t797 trim_val\[3\] a_11374_1251# VPWR.t796 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1069 a_9004_3677# _033_ VPWR.t1877 VPWR.t1876 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1070 cal_count\[2\] a_13470_7663# VPWR.t930 VPWR.t929 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1071 VPWR.t3242 a_8820_12533# ctlp[5].t0 VPWR.t3241 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1072 VPWR.t239 VGND.t3334 VPWR.t238 VPWR.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1073 VPWR.t1776 clknet_2_0__leaf_clk a_1867_3317# VPWR.t1775 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1074 net11 net19 VGND.t3134 VGND.t3133 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1075 VGND.t2179 a_4655_10071# _019_ VGND.t2178 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1076 a_7310_2223# a_7184_2339# a_6906_2355# VGND.t2694 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1077 VGND.t507 a_3933_2767# _051_.t9 VGND.t506 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1078 a_2910_12131# net29 a_2828_12131# VPWR.t2900 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1079 a_1137_11721# _074_ VPWR.t884 VPWR.t883 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1080 VGND.t1387 VPWR.t3404 VGND.t1386 VGND.t1385 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1081 VGND.t1384 VPWR.t3405 VGND.t1383 VGND.t1382 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1082 _055_ a_14604_3017# VGND.t118 VGND.t117 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1083 a_1313_10901# a_1095_11305# VPWR.t2878 VPWR.t2877 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1084 a_7723_10143# net44 VPWR.t2849 VPWR.t2848 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1085 VGND.t1381 VPWR.t3406 VGND.t1380 VGND.t1379 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1086 a_4609_9295# a_4443_9295# VGND.t1910 VGND.t1909 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1087 a_10543_2455# trim_mask\[4\] a_10689_2223# VPWR.t1906 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1088 VGND.t1930 net14 net6 VGND.t1929 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1089 VGND.t1378 VPWR.t3407 VGND.t1377 VGND.t1376 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1090 state\[0\] a_3123_3615# VPWR.t2964 VPWR.t2963 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1091 VGND.t1375 VPWR.t3408 VGND.t1374 VGND.t1373 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1092 a_5363_4719# _059_ VGND.t1709 VGND.t1708 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.0878 ps=0.92 w=0.65 l=0.15
X1093 VPWR.t2372 net37.t4 a_15023_9839# VPWR.t2371 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1094 a_1638_7485# a_561_7119# a_1476_7119# VPWR.t1003 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1095 a_12436_9129# a_11987_8757# a_12341_8751# VGND.t2892 sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X1096 VGND.t2071 _122_ a_13279_7119# VGND.t2070 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X1097 VPWR.t242 VGND.t3335 VPWR.t241 VPWR.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1098 VPWR.t1516 a_10903_7261# a_10864_7387# VPWR.t1515 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1099 VPWR.t245 VGND.t3336 VPWR.t244 VPWR.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1100 net22 a_1651_6005# VGND.t2844 VGND.t2843 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1101 a_13193_6031# net2 a_13111_6031# VGND.t2382 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X1102 VPWR.t1164 a_9003_3829# _119_ VPWR.t1163 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1103 a_10699_3311# _064_ a_10781_3631# VGND.t1606 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1104 a_5089_10159# _101_ a_4655_10071# VGND.t796 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1105 VGND.t1372 VPWR.t3409 VGND.t1371 VGND.t1370 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1106 a_3868_7119# a_2953_7119# a_3521_7361# VGND.t1975 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1107 a_2476_6281# net22 VPWR.t3168 VPWR.t3167 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.34 w=0.42 l=0.15
X1108 VPWR.t2546 cal_itt\[0\] a_8949_6281# VPWR.t2545 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1109 a_9317_3285# a_9099_3689# VPWR.t2653 VPWR.t2652 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1110 a_6316_5193# _048_.t21 a_6566_5193# VPWR.t2319 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1111 clknet_2_0__leaf_clk a_2857_5461# VGND.t674 VGND.t673 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1112 net25 a_1651_10143# VPWR.t2859 VPWR.t2858 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1113 VGND.t1369 VPWR.t3410 VGND.t1368 VGND.t1367 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1114 _063_.t7 cal_itt\[0\] VPWR.t2544 VPWR.t2543 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X1115 clknet_2_3__leaf_clk a_8298_5487# VPWR.t2149 VPWR.t2148 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1116 VPWR.t2681 mask\[4\] a_9074_9955# VPWR.t2680 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1117 a_8025_8041# a_6835_7669# a_7916_8041# VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1118 VGND.t1366 VPWR.t3411 VGND.t1365 VGND.t1364 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1119 VPWR.t3151 clk.t1 a_8022_7119# VPWR.t3150 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1120 net35 a_14655_4399# VGND.t571 VGND.t544 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1121 VPWR.t1432 a_2857_5461# clknet_2_0__leaf_clk VPWR.t1431 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1122 net43.t2 a_1467_7923# VPWR.t1263 VPWR.t1262 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1123 VPWR.t2526 net45 a_4995_7119# VPWR.t2525 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1124 net16 a_13919_8751# VGND.t3080 VGND.t3079 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1125 a_9734_2223# a_8657_2229# a_9572_2601# VPWR.t1498 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1126 a_5915_10927# _101_ a_5997_10927# VPWR.t1551 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1127 a_1835_12319# net43.t17 VPWR.t2748 VPWR.t2747 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1128 trimb[1].t7 a_15023_9839# VGND.t3249 VGND.t3248 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1129 VGND.t2703 net43.t18 a_1173_7119# VGND.t2702 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1130 a_4805_8207# a_3615_8207# a_4696_8207# VGND.t1667 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1131 ctlp[7].t6 a_5363_12559# VGND.t2043 VGND.t2042 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1132 VGND.t841 a_8022_7119# clknet_0_clk VGND.t840 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1133 VPWR.t248 VGND.t3337 VPWR.t247 VPWR.t246 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1134 VPWR.t1430 a_2857_5461# clknet_2_0__leaf_clk VPWR.t1429 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1135 VPWR.t251 VGND.t3338 VPWR.t250 VPWR.t249 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1136 VPWR.t746 net40 a_15023_8751# VPWR.t745 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1137 VPWR.t807 a_10005_6031# _092_ VPWR.t806 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1138 VPWR.t254 VGND.t3339 VPWR.t253 VPWR.t252 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1139 VGND.t2051 _116_ a_9805_1473# VGND.t2050 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1140 VGND.t3216 a_3667_3829# _048_.t10 VGND.t3215 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1141 VPWR.t257 VGND.t3340 VPWR.t256 VPWR.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1142 a_8657_2229# a_8491_2229# VPWR.t2360 VPWR.t2359 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1143 a_7548_10217# a_6633_9845# a_7201_9813# VGND.t2766 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1144 cal_count\[0\] a_11814_9295# VPWR.t1283 VPWR.t1282 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X1145 VPWR.t1729 _059_ a_5537_4105# VPWR.t1728 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1146 a_12121_3677# a_12077_3285# a_11955_3689# VGND.t1801 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1147 VPWR.t1589 a_8022_7119# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1148 VPWR.t2981 a_8673_10625# a_8563_10749# VPWR.t2980 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1149 ctln[6].t2 a_6927_591# VPWR.t1806 VPWR.t1805 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1150 a_9664_3689# a_8583_3317# a_9317_3285# VPWR.t2686 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1151 VGND.t2444 a_455_12533# result[6].t6 VGND.t2443 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1152 VGND.t2422 a_8298_2767# clknet_2_2__leaf_clk VGND.t2421 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1153 net27 a_7631_12319# VGND.t610 VGND.t609 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1154 VGND.t1663 _107_ _108_ VGND.t1662 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1155 a_5067_9661# a_4443_9295# a_4959_9295# VPWR.t1933 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1156 a_13016_9117# a_12436_9129# VGND.t461 VGND.t460 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1157 VPWR.t260 VGND.t3341 VPWR.t259 VPWR.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1158 _130_ a_14788_7369# VPWR.t2308 VPWR.t2307 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1159 a_4609_1679# a_4443_1679# VGND.t1949 VGND.t1948 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1160 a_14894_3677# net46 VGND.t243 VGND.t242 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1161 a_12778_3677# net46 VGND.t241 VGND.t240 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1162 VPWR.t1674 a_995_3530# net1 VPWR.t1673 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1163 a_12047_2601# a_11601_2229# a_11951_2601# VGND.t408 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1164 a_6927_3311# _049_ VPWR.t1196 VPWR.t1195 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.225 ps=1.45 w=1 l=0.15
X1165 _026_ a_11067_3017# VPWR.t1923 VPWR.t1922 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1166 VPWR.t3295 a_3667_3829# _048_.t3 VPWR.t3294 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1167 _101_ net51 a_5363_7369# VPWR.t1128 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1168 VGND.t2972 mask\[7\] a_2828_12131# VGND.t2971 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1169 VGND.t2621 net33 net38 VGND.t2620 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1170 VPWR.t2287 net36 a_15023_10927# VPWR.t2286 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1171 VGND.t1363 VPWR.t3412 VGND.t1362 VGND.t1361 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1172 _090_ _087_ VGND.t114 VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1173 a_7999_11231# net44 VPWR.t2847 VPWR.t2846 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1174 VGND.t1360 VPWR.t3413 VGND.t1359 VGND.t1358 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1175 a_14686_2339# trim_mask\[2\] a_14604_2339# VPWR.t2888 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1176 VGND.t2485 net45 a_1173_6031# VGND.t2484 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1177 VGND.t1357 VPWR.t3414 VGND.t1356 VGND.t1355 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1178 VGND.t801 a_4687_12319# a_4621_12393# VGND.t800 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1179 VPWR.t1021 clknet_2_2__leaf_clk a_13091_1141# VPWR.t1020 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1180 VPWR.t2147 a_8298_5487# clknet_2_3__leaf_clk VPWR.t2146 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1181 VPWR.t2551 a_7723_10143# a_7710_9839# VPWR.t2550 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1182 a_14807_8359# cal_count\[1\] VPWR.t2200 VPWR.t2199 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X1183 VPWR.t2401 a_7223_2465# a_7184_2339# VPWR.t2400 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1184 a_10747_8970# _124_ VGND.t690 VGND.t689 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1185 VGND.t3172 a_448_11445# result[5].t3 VGND.t3171 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X1186 a_2645_3677# a_2601_3285# a_2479_3689# VGND.t1991 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1187 a_745_12021# a_579_12021# VPWR.t1310 VPWR.t1309 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1188 _011_ _074_ VGND.t147 VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1189 VGND.t1354 VPWR.t3415 VGND.t1353 VGND.t1352 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1190 a_1651_4703# net45 VPWR.t2524 VPWR.t2523 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1191 VGND.t1351 VPWR.t3416 VGND.t1350 VGND.t1349 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1192 a_1203_10927# net43.t19 VPWR.t2750 VPWR.t2749 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1193 a_7259_11305# a_6743_10933# a_7164_11293# VGND.t2535 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1194 a_8551_10383# a_8105_10383# a_8455_10383# VGND.t2836 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1195 _128_ a_14347_9480# VGND.t561 VGND.t560 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1196 a_14063_7093# _129_ a_14282_7119# VGND.t804 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.091 ps=0.93 w=0.65 l=0.15
X1197 VGND.t2483 net45 a_2921_2589# VGND.t2482 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1198 a_10219_2045# net46 VPWR.t989 VPWR.t988 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1199 VGND.t1901 a_13881_1653# _114_ VGND.t1900 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1200 a_3399_2527# a_3224_2601# a_3578_2589# VGND.t2925 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1201 _029_ a_12723_4943# VPWR.t1406 VPWR.t1405 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1202 _120_ a_3273_4943# VPWR.t2117 VPWR.t2116 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.195 ps=1.39 w=1 l=0.15
X1203 a_5829_9839# _074_ VPWR.t882 VPWR.t881 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1204 VPWR.t263 VGND.t3342 VPWR.t262 VPWR.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1205 clknet_0_clk a_8022_7119# VGND.t839 VGND.t838 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1206 VPWR.t831 net18 net10 VPWR.t830 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1207 a_12148_4777# a_11233_4405# a_11801_4373# VGND.t1853 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1208 VPWR.t2457 a_8298_2767# clknet_2_2__leaf_clk VPWR.t2456 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1209 VGND.t1348 VPWR.t3417 VGND.t1347 VGND.t1346 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1210 VPWR.t3027 mask\[7\] a_2910_12131# VPWR.t3026 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1211 a_2288_3677# _013_ VGND.t2434 VGND.t2433 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1212 a_7310_2223# a_7223_2465# a_6906_2355# VPWR.t2399 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.0588 ps=0.7 w=0.42 l=0.15
X1213 VPWR.t266 VGND.t3343 VPWR.t265 VPWR.t264 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1214 VGND.t763 a_10903_7261# a_10864_7387# VGND.t762 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1215 ctln[3].t0 a_12631_591# VPWR.t1716 VPWR.t1715 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X1216 VPWR.t269 VGND.t3344 VPWR.t268 VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1217 VGND.t365 a_2857_7637# clknet_2_1__leaf_clk.t26 VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1218 _132_ _130_ VPWR.t2984 VPWR.t2656 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1219 VGND.t433 a_12520_7637# a_12454_8041# VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1220 clknet_2_2__leaf_clk a_8298_2767# VGND.t2420 VGND.t2419 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1221 a_5691_2741# state\[2\] VPWR.t1985 VPWR.t1984 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1222 VPWR.t272 VGND.t3345 VPWR.t271 VPWR.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1223 VGND.t2579 _050_ a_5547_5603# VGND.t2578 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X1224 a_4621_12393# a_3431_12021# a_4512_12393# VGND.t435 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1225 VPWR.t2068 a_5363_12559# ctlp[7].t1 VPWR.t2067 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1226 a_12520_7637# net47 VPWR.t1698 VPWR.t1697 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X1227 a_911_6031# a_561_6031# a_816_6031# VPWR.t2624 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1228 VGND.t1345 VPWR.t3418 VGND.t1344 VGND.t1343 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1229 a_3530_4765# _096_ VGND.t306 VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1230 VGND.t3044 _078_ a_1579_11471# VGND.t3043 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X1231 a_14347_9480# cal_count\[0\] VGND.t2947 VGND.t2946 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1232 VPWR.t275 VGND.t3346 VPWR.t274 VPWR.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1233 a_7618_12015# a_6541_12021# a_7456_12393# VPWR.t794 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1234 VPWR.t278 VGND.t3347 VPWR.t277 VPWR.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1235 VGND.t1654 a_995_3530# net1 VGND.t1653 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1236 _065_.t1 a_4091_5309# VPWR.t2123 VPWR.t2122 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.331 ps=1.71 w=1 l=0.15
X1237 net40 net35 VGND.t577 VGND.t576 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1238 a_12916_8751# a_12436_9129# VPWR.t1202 VPWR.t1201 sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X1239 VPWR.t1289 a_12992_8751# a_13562_8751# VPWR.t1288 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1240 cal_count\[3\] a_12231_6005# VGND.t166 VGND.t165 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1241 VGND.t1841 _043_ a_9871_10383# VGND.t1840 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1242 VPWR.t3230 a_13050_7637# a_13008_7663# VPWR.t3229 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1243 a_10851_1653# net46 VPWR.t987 VPWR.t986 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1244 clknet_2_3__leaf_clk a_8298_5487# VPWR.t2145 VPWR.t2144 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1245 VGND.t1847 a_5363_591# ctln[7].t6 VGND.t1846 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1246 VGND.t2122 a_8298_5487# clknet_2_3__leaf_clk VGND.t2121 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1247 VPWR.t940 net16 a_14471_12559# VPWR.t939 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1248 a_11369_7119# a_10990_7485# a_11297_7119# VGND.t1915 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1249 a_9166_4515# _106_ a_9084_4515# VPWR.t753 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1250 VGND.t2319 a_455_8181# result[2].t6 VGND.t2318 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1251 a_13142_8359# _123_.t6 a_13356_8457# VPWR.t1656 sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.117 ps=1.24 w=1 l=0.15
X1252 mask\[5\] a_7999_11231# VPWR.t3260 VPWR.t3259 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1253 VGND.t1342 VPWR.t3419 VGND.t1341 VGND.t1140 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1254 a_7001_7669# a_6835_7669# VGND.t52 VGND.t51 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1255 VGND.t1679 net47 a_11508_9295# VGND.t1678 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
X1256 clknet_2_1__leaf_clk.t9 a_2857_7637# VPWR.t1100 VPWR.t1099 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1257 VGND.t1340 VPWR.t3420 VGND.t1339 VGND.t1338 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1258 trim[2].t2 a_15023_2223# VPWR.t3214 VPWR.t3213 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1259 VGND.t1865 net15 net7 VGND.t1864 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1260 VGND.t1337 VPWR.t3421 VGND.t1336 VGND.t1335 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1261 VGND.t579 a_6793_8970# net53 VGND.t578 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1262 VPWR.t1881 a_7109_11989# a_6999_12015# VPWR.t1880 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1263 net52 a_5691_7637# VPWR.t2635 VPWR.t2634 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1264 a_9405_9295# a_8215_9295# a_9296_9295# VGND.t1934 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1265 _094_ _049_ a_3529_6281# VPWR.t1194 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1266 a_3933_2767# state\[1\] VGND.t3060 VGND.t3059 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1267 VGND.t2396 net52 _102_ VGND.t2395 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1268 VPWR.t2493 a_4687_11231# a_4674_10927# VPWR.t2492 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1269 VGND.t40 a_3063_591# ctln[1].t3 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1270 VGND.t1334 VPWR.t3422 VGND.t1333 VGND.t1134 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1271 VPWR.t2762 _051_.t14 a_7800_4631# VPWR.t2761 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1272 trim[4].t6 a_15023_5487# VGND.t493 VGND.t492 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1273 VGND.t1724 _095_ _096_ VGND.t1723 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1274 VPWR.t1828 clknet_2_1__leaf_clk.t39 a_3431_12021# VPWR.t1827 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1275 a_14334_1135# a_13257_1141# a_14172_1513# VPWR.t2818 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1276 a_14184_2767# trim_mask\[1\] a_13881_2741# VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X1277 VPWR.t2932 _054_ a_7939_3855# VPWR.t2931 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1278 VGND.t284 clknet_2_2__leaf_clk a_8491_2229# VGND.t283 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1279 a_11491_6031# a_11141_6031# a_11396_6031# VPWR.t2778 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1280 a_9125_4943# _048_.t22 _105_ VGND.t2288 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1281 a_8673_10625# a_8455_10383# VGND.t36 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1282 VGND.t2688 a_15023_1135# trim[3].t5 VGND.t2687 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1283 a_5445_4399# net54 VPWR.t1402 VPWR.t1401 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X1284 VPWR.t2009 a_7527_4631# _088_ VPWR.t2008 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X1285 a_14552_9071# cal_count\[0\] a_14249_8725# VGND.t2945 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X1286 a_3511_11471# mask\[6\] _085_ VGND.t606 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1287 VGND.t1332 VPWR.t3423 VGND.t1331 VGND.t1330 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1288 VGND.t2418 a_8298_2767# clknet_2_2__leaf_clk VGND.t2417 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1289 VGND.t1718 a_6519_4631# _100_ VGND.t1717 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1290 a_15083_4659# net32 VGND.t474 VGND.t473 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X1291 _029_ a_12723_4943# VGND.t652 VGND.t651 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1292 a_9957_7663# _067_ VPWR.t922 VPWR.t921 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X1293 a_8935_6895# cal_itt\[1\] a_8745_6895# VGND.t1619 sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0878 ps=0.92 w=0.65 l=0.15
X1294 VPWR.t281 VGND.t3348 VPWR.t280 VPWR.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1295 VPWR.t284 VGND.t3349 VPWR.t283 VPWR.t282 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1296 VPWR.t3025 mask\[7\] a_1493_11721# VPWR.t3024 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X1297 a_8827_9295# a_8381_9295# a_8731_9295# VGND.t3228 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1298 VGND.t34 net42 _103_ VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1299 VPWR.t2184 a_15023_12015# trimb[2].t2 VPWR.t2183 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1300 a_10016_1679# _032_ VGND.t3148 VGND.t3147 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1301 a_9115_2223# a_8491_2229# a_9007_2601# VPWR.t2358 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1302 VPWR.t287 VGND.t3350 VPWR.t286 VPWR.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1303 trimb[1].t6 a_15023_9839# VGND.t3247 VGND.t3246 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1304 net47 a_9463_8725# VGND.t790 VGND.t789 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1305 VGND.t1987 net38 a_15023_12015# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1306 VPWR.t3254 a_12323_4703# trim_mask\[0\] VPWR.t3253 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1307 result[1].t1 a_448_7637# VPWR.t3240 VPWR.t3239 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1308 VPWR.t290 VGND.t3351 VPWR.t289 VPWR.t288 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1309 VGND.t2241 a_6927_12559# ctlp[6].t5 VGND.t2240 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1310 VGND.t1329 VPWR.t3424 VGND.t1328 VGND.t1327 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1311 a_6056_8359# _065_.t10 a_6198_8534# VPWR.t3312 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1312 VGND.t1326 VPWR.t3425 VGND.t1325 VGND.t1324 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1313 VGND.t440 a_5699_9269# a_5633_9295# VGND.t439 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1314 VGND.t211 trim_val\[0\] a_14972_5193# VGND.t210 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1315 a_3399_7119# a_2953_7119# a_3303_7119# VGND.t1974 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1316 VPWR.t1588 a_8022_7119# clknet_0_clk VPWR.t1587 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1317 a_2767_2223# net45 VPWR.t2522 VPWR.t2521 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1318 a_4165_11989# a_3947_12393# VGND.t466 VGND.t465 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1319 a_10689_2223# _064_ a_10543_2455# VPWR.t1621 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X1320 VGND.t1323 VPWR.t3426 VGND.t1322 VGND.t1321 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1321 VPWR.t3314 _065_.t11 a_3830_6281# VPWR.t3313 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1322 VGND.t2753 net8 a_14471_591# VGND.t2752 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1323 VPWR.t293 VGND.t3352 VPWR.t292 VPWR.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1324 trim_val\[4\] a_9839_3615# VPWR.t3037 VPWR.t3036 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1325 a_7153_12381# a_7109_11989# a_6987_12393# VGND.t1855 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1326 result[2].t5 a_455_8181# VGND.t2317 VGND.t2316 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X1327 VPWR.t296 VGND.t3353 VPWR.t295 VPWR.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1328 VGND.t431 _056_ a_15023_1679# VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1329 a_7689_2589# a_7310_2223# a_7617_2589# VGND.t3154 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1330 VGND.t2442 a_455_12533# result[6].t5 VGND.t2441 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1331 a_12344_8041# a_12061_7669# a_12249_7663# VPWR.t1979 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.125 ps=1.17 w=0.42 l=0.15
X1332 VGND.t1320 VPWR.t3427 VGND.t1319 VGND.t1318 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1333 a_3116_12533# net15 VPWR.t1893 VPWR.t1892 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1334 VPWR.t2520 net45 a_7524_2223# VPWR.t2519 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.109 ps=1.36 w=0.42 l=0.15
X1335 VPWR.t2277 a_15083_4659# trim[1].t2 VPWR.t2276 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1336 a_1095_12393# a_745_12021# a_1000_12381# VPWR.t3220 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1337 a_7824_11305# a_6743_10933# a_7477_10901# VPWR.t2571 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1338 a_8105_10383# a_7939_10383# VGND.t206 VGND.t205 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1339 VGND.t1317 VPWR.t3428 VGND.t1316 VGND.t1315 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1340 _123_.t1 _053_ a_10877_7983# VGND.t2566 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1341 a_14526_1501# net46 VGND.t239 VGND.t238 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1342 VGND.t2143 _063_.t12 _064_ VGND.t2142 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1343 a_4866_11293# net43.t20 VGND.t2705 VGND.t2704 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1344 a_14467_8751# _125_ a_14249_8725# VPWR.t2041 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1345 a_2288_3677# _013_ VPWR.t2467 VPWR.t2466 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1346 a_13915_4399# trim_val\[0\] a_13697_4373# VPWR.t947 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1347 a_9443_6059# _053_ VPWR.t2607 VPWR.t2606 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1348 a_2828_12131# net29 VGND.t2856 VGND.t2855 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1349 net2 a_15259_7637# VPWR.t2657 VPWR.t2656 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1350 ctlp[0].t3 a_1099_12533# VPWR.t1477 VPWR.t1476 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1351 a_4512_12393# a_3597_12021# a_4165_11989# VGND.t2967 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1352 a_1585_10217# a_395_9845# a_1476_10217# VGND.t2090 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1353 VPWR.t1904 a_13825_1109# a_13715_1135# VPWR.t1903 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1354 VPWR.t299 VGND.t3354 VPWR.t298 VPWR.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1355 a_9225_2197# a_9007_2601# VGND.t2371 VGND.t2370 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1356 trimb[0].t2 a_15023_10927# VPWR.t2049 VPWR.t2048 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1357 VPWR.t302 VGND.t3355 VPWR.t301 VPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1358 trim_val\[1\] a_14715_3615# VGND.t1628 VGND.t1627 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1359 trim_mask\[1\] a_12599_3615# VGND.t3220 VGND.t3219 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1360 a_1279_9129# a_929_8757# a_1184_9117# VPWR.t2768 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1361 VPWR.t3202 a_1129_6273# a_1019_6397# VPWR.t3201 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1362 trim[3].t4 a_15023_1135# VGND.t2686 VGND.t2685 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1363 a_10137_4943# _062_.t11 VGND.t2210 VGND.t2209 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.107 ps=0.98 w=0.65 l=0.15
X1364 a_5455_4943# _075_ VPWR.t1386 VPWR.t1385 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1365 VPWR.t1830 clknet_2_1__leaf_clk.t40 a_763_8757# VPWR.t1829 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1366 VGND.t2850 a_13059_4631# _111_ VGND.t2849 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1367 VPWR.t305 VGND.t3356 VPWR.t304 VPWR.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1368 VGND.t1314 VPWR.t3429 VGND.t1313 VGND.t1312 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1369 VGND.t2660 a_14807_8359# _125_ VGND.t2659 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1370 a_1019_7485# a_395_7119# a_911_7119# VPWR.t1816 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1371 VPWR.t2321 _048_.t23 _062_.t1 VPWR.t2320 sky130_fd_pr__pfet_01v8_hvt ad=0.176 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X1372 _079_ net22 VGND.t3100 VGND.t3099 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1373 result[5].t2 a_448_11445# VGND.t3170 VGND.t3169 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1374 VPWR.t1162 a_9003_3829# _119_ VPWR.t1161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1375 VGND.t1311 VPWR.t3430 VGND.t1310 VGND.t1309 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1376 a_8563_10749# a_7939_10383# a_8455_10383# VPWR.t943 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1377 a_6316_5193# a_6210_4989# _098_ VPWR.t3164 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1378 _050_ a_5691_2741# VGND.t2543 VGND.t2542 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1379 VGND.t3 net39 a_15023_12559# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1380 a_4498_4373# net54 VGND.t650 VGND.t649 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.123 ps=1.03 w=0.65 l=0.15
X1381 VGND.t1308 VPWR.t3431 VGND.t1307 VGND.t1306 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1382 VGND.t388 net51 a_5691_7637# VGND.t387 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1383 VGND.t672 a_2857_5461# clknet_2_0__leaf_clk VGND.t671 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1384 mask\[2\] a_4043_10143# VGND.t2747 VGND.t2746 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1385 a_1585_7119# a_395_7119# a_1476_7119# VGND.t1795 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1386 VPWR.t2237 _062_.t12 a_5455_4943# VPWR.t2236 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1387 VPWR.t2143 a_8298_5487# clknet_2_3__leaf_clk VPWR.t2142 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1388 VPWR.t308 VGND.t3357 VPWR.t307 VPWR.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1389 _051_.t4 a_3933_2767# VPWR.t1249 VPWR.t1248 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1390 a_11233_4405# a_11067_4405# VGND.t2559 VGND.t2558 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1391 VPWR.t3074 net34.t4 a_15023_1135# VPWR.t3073 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1392 a_8022_7119# clk.t2 VPWR.t3153 VPWR.t3152 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1393 a_13059_4631# _109_ a_13233_4737# VGND.t3069 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1394 a_2857_5461# clknet_0_clk VPWR.t1066 VPWR.t1065 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1395 VGND.t1305 VPWR.t3432 VGND.t1304 VGND.t1303 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1396 VPWR.t1261 a_1467_7923# net43.t1 VPWR.t1260 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1397 VGND.t2651 a_5699_1653# a_5633_1679# VGND.t2650 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1398 VGND.t2145 _063_.t13 a_9529_6059# VGND.t2144 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1399 VGND.t363 a_2857_7637# clknet_2_1__leaf_clk.t25 VGND.t362 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1400 a_9826_3311# a_8749_3317# a_9664_3689# VPWR.t2917 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1401 a_2368_9955# net25 VGND.t3067 VGND.t3066 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1402 _042_.t0 a_2368_9955# VPWR.t2555 VPWR.t2554 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1403 trim_mask\[0\] a_12323_4703# VGND.t3180 VGND.t3179 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X1404 _104_ net30.t7 a_8307_4719# VGND.t29 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1405 a_1387_8751# a_763_8757# a_1279_9129# VPWR.t823 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1406 VPWR.t805 a_10005_6031# _092_ VPWR.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1407 VGND.t21 a_4995_7119# net44 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X1408 a_5067_2045# a_4443_1679# a_4959_1679# VPWR.t1975 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1409 trim[1].t1 a_15083_4659# VPWR.t2275 VPWR.t2274 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1410 VGND.t1661 _107_ _108_ VGND.t1660 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1411 VGND.t168 a_7723_6807# _073_ VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1412 clknet_2_2__leaf_clk a_8298_2767# VPWR.t2455 VPWR.t2454 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1413 VGND.t1302 VPWR.t3433 VGND.t1301 VGND.t1300 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1414 a_1095_12393# a_579_12021# a_1000_12381# VGND.t568 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1415 VPWR.t311 VGND.t3358 VPWR.t310 VPWR.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1416 a_11258_9117# cal_count\[0\] VGND.t2944 VGND.t2943 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X1417 a_4677_7882# _040_ VGND.t2675 VGND.t2674 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1418 a_10975_4105# _064_ a_11057_4105# VPWR.t1620 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1419 a_14347_9480# _127_ a_14733_9545# VPWR.t3149 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1420 ctln[7].t1 a_5363_591# VPWR.t1869 VPWR.t1868 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1421 a_14649_3689# a_13459_3317# a_14540_3689# VGND.t180 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1422 a_2865_4460# _095_ VGND.t1722 VGND.t1721 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1423 VPWR.t1631 a_1660_12393# a_1835_12319# VPWR.t1630 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1424 VPWR.t1774 clknet_2_0__leaf_clk a_3615_8207# VPWR.t1773 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1425 VGND.t81 net31 a_15023_2767# VGND.t80 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1426 VPWR.t314 VGND.t3359 VPWR.t313 VPWR.t312 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1427 a_10593_9295# _035_ VGND.t766 VGND.t765 sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X1428 VPWR.t2218 net20.t3 net12 VPWR.t2217 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1429 VGND.t1299 VPWR.t3434 VGND.t1298 VGND.t1297 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1430 a_9650_9295# net47 VGND.t1677 VGND.t1676 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1431 a_1585_6031# a_395_6031# a_1476_6031# VGND.t558 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1432 a_4973_2773# state\[2\] a_4901_2773# VGND.t1958 sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X1433 valid.t3 a_455_3571# VPWR.t2196 VPWR.t2195 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1434 net25 a_1651_10143# VGND.t2810 VGND.t2809 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1435 VGND.t1296 VPWR.t3435 VGND.t1295 VGND.t1294 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1436 VGND.t3191 a_14564_6397# _061_ VGND.t574 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.0878 ps=0.92 w=0.65 l=0.15
X1437 VGND.t1293 VPWR.t3436 VGND.t1292 VGND.t1291 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1438 net41 _060_ VGND.t2204 VGND.t2203 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1439 VPWR.t317 VGND.t3360 VPWR.t316 VPWR.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1440 VGND.t327 clknet_0_clk a_2857_7637# VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1441 a_7447_8041# a_7001_7669# a_7351_8041# VGND.t697 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1442 a_10820_7485# a_10383_7093# VPWR.t3066 VPWR.t3065 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1443 _115_ a_13307_1707# VPWR.t932 VPWR.t931 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1444 VGND.t282 clknet_2_2__leaf_clk a_13459_3317# VGND.t281 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1445 VGND.t17 _106_ _108_ VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1446 VPWR.t320 VGND.t3361 VPWR.t319 VPWR.t318 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1447 a_5067_9661# net44 VPWR.t2845 VPWR.t2844 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1448 a_9003_3829# _118_ a_9478_4105# VPWR.t2407 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.3 ps=2.6 w=1 l=0.15
X1449 clknet_2_3__leaf_clk a_8298_5487# VPWR.t2141 VPWR.t2140 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1450 clknet_2_0__leaf_clk a_2857_5461# VGND.t670 VGND.t669 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1451 VGND.t448 a_6056_8359# _077_ VGND.t447 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X1452 clknet_2_1__leaf_clk.t8 a_2857_7637# VPWR.t1098 VPWR.t1097 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1453 a_3411_9839# net43.t21 VPWR.t2752 VPWR.t2751 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1454 net24 a_2019_9055# VGND.t1979 VGND.t1978 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1455 net45 a_3339_2767# VGND.t2862 VGND.t2861 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1456 clknet_2_3__leaf_clk a_8298_5487# VGND.t2120 VGND.t2119 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1457 a_4696_8207# a_3615_8207# a_4349_8449# VPWR.t1685 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1458 net10 net18 VPWR.t829 VPWR.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1459 a_1476_4777# a_561_4405# a_1129_4373# VGND.t1924 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1460 VGND.t1290 VPWR.t3437 VGND.t1289 VGND.t1288 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1461 VGND.t1650 a_9471_9269# cal_itt\[0\] VGND.t1649 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1462 VPWR.t323 VGND.t3362 VPWR.t322 VPWR.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1463 _084_ net27 a_5915_11721# VPWR.t1885 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1464 VGND.t2226 _068_ _000_ VGND.t2225 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1465 VGND.t1287 VPWR.t3438 VGND.t1286 VGND.t1285 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1466 a_816_10205# _007_ VPWR.t2894 VPWR.t2893 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1467 VPWR.t1760 _058_ a_14655_4399# VPWR.t1759 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1468 VGND.t2337 a_13697_4373# _109_ VGND.t2336 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1469 VGND.t3232 _065_.t12 _001_ VGND.t3231 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1470 VGND.t729 a_5535_8181# _078_ VGND.t728 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1471 a_14083_3311# a_13459_3317# a_13975_3689# VPWR.t917 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1472 a_1476_10217# a_561_9845# a_1129_9813# VGND.t3110 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1473 net32 a_15299_3311# VPWR.t2310 VPWR.t2309 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1474 VPWR.t1696 net47 a_12900_7663# VPWR.t1695 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X1475 VPWR.t1257 a_3399_2527# a_3386_2223# VPWR.t1256 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1476 VPWR.t1501 a_5524_9295# a_5699_9269# VPWR.t1500 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1477 VGND.t837 a_8022_7119# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1478 a_7677_4759# trim_mask\[0\] VGND.t1873 VGND.t1872 sky130_fd_pr__nfet_01v8 ad=0.0536 pd=0.675 as=0.122 ps=1.08 w=0.42 l=0.15
X1479 VPWR.t1394 a_3388_4631# _097_ VPWR.t1393 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1480 VGND.t126 a_10864_9269# a_10798_9295# VGND.t125 sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.0671 ps=0.75 w=0.42 l=0.15
X1481 a_2869_11247# mask\[6\] VGND.t605 VGND.t604 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1482 VGND.t721 a_1099_12533# ctlp[0].t6 VGND.t720 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1483 a_14788_7369# cal_count\[2\] VGND.t2190 VGND.t2189 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1484 _007_ _074_ VGND.t145 VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1485 VGND.t2239 a_6927_12559# ctlp[6].t4 VGND.t2238 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1486 a_2225_7983# mask\[0\] VGND.t2989 VGND.t2988 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1487 a_4425_6031# a_4259_6031# VGND.t311 VGND.t310 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1488 a_745_10933# a_579_10933# VGND.t592 VGND.t591 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1489 VPWR.t3262 a_3868_7119# a_4043_7093# VPWR.t3261 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1490 a_9823_6941# _062_.t13 a_9460_6807# VGND.t2211 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X1491 VPWR.t2933 a_2815_9447# _018_ VPWR.t1833 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X1492 VPWR.t1586 a_8022_7119# clknet_0_clk VPWR.t1585 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1493 clknet_2_1__leaf_clk.t24 a_2857_7637# VGND.t361 VGND.t360 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1494 _069_ cal_itt\[1\] VGND.t1618 VGND.t1617 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1495 a_10872_1455# trim_mask\[3\] a_10569_1109# VGND.t2078 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X1496 net7 net15 VPWR.t1891 VPWR.t1890 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1497 a_14565_9295# _127_ _128_ VGND.t3083 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.25 ps=1.42 w=0.65 l=0.15
X1498 a_5423_9011# _065_.t13 VGND.t3234 VGND.t3233 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X1499 VPWR.t1842 a_11709_6273# a_11599_6397# VPWR.t1841 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1500 VPWR.t326 VGND.t3363 VPWR.t325 VPWR.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1501 a_7613_8029# a_7569_7637# a_7447_8041# VGND.t3204 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1502 a_14807_8359# net2 a_14981_8235# VGND.t2381 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1503 VPWR.t329 VGND.t3364 VPWR.t328 VPWR.t327 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1504 a_13715_5309# net46 VPWR.t985 VPWR.t984 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1505 a_14422_7093# _131_ VPWR.t3085 VPWR.t3084 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1506 a_7723_6807# cal_itt\[3\] a_7897_6913# VGND.t2908 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1507 a_13307_1707# _110_.t5 VPWR.t2168 VPWR.t2167 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1508 a_13825_1109# a_13607_1513# VGND.t406 VGND.t405 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1509 VGND.t1826 net53 a_6445_10383# VGND.t1825 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1510 _016_ a_2143_7663# VGND.t2875 VGND.t2874 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1511 VGND.t2577 _050_ a_7891_3617# VGND.t2576 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1512 VGND.t1284 VPWR.t3439 VGND.t1283 VGND.t1282 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1513 a_6763_5193# calibrate a_6566_5193# VPWR.t1492 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1514 VPWR.t332 VGND.t3365 VPWR.t331 VPWR.t330 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1515 VGND.t1281 VPWR.t3440 VGND.t1280 VGND.t1279 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1516 VPWR.t335 VGND.t3366 VPWR.t334 VPWR.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1517 VPWR.t1019 clknet_2_2__leaf_clk a_11067_4405# VPWR.t1018 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1518 a_3817_4697# _096_ VPWR.t1042 VPWR.t1041 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1519 a_4864_9295# _019_ VPWR.t2922 VPWR.t2921 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1520 result[3].t2 a_448_9269# VGND.t2448 VGND.t2447 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1521 VGND.t3140 a_15023_2223# trim[2].t7 VGND.t1998 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1522 a_4209_12381# a_4165_11989# a_4043_12393# VGND.t3125 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1523 a_14193_3285# a_13975_3689# VGND.t259 VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1524 VPWR.t2139 a_8298_5487# clknet_2_3__leaf_clk VPWR.t2138 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1525 a_8820_12533# net19 VPWR.t3206 VPWR.t3205 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1526 a_3667_3829# state\[0\] VPWR.t1458 VPWR.t1457 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1527 a_14347_4917# net46 VPWR.t983 VPWR.t982 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1528 a_6796_12381# _009_ VPWR.t2243 VPWR.t2242 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1529 VPWR.t338 VGND.t3367 VPWR.t337 VPWR.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1530 a_10699_5487# _136_ a_10781_5487# VPWR.t788 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1531 a_8673_10625# a_8455_10383# VPWR.t775 VPWR.t774 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1532 a_561_7119# a_395_7119# VPWR.t1815 VPWR.t1814 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1533 trimb[0].t1 a_15023_10927# VPWR.t2047 VPWR.t2046 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1534 a_10752_12533# net18 VPWR.t827 VPWR.t826 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1535 a_2961_9545# _101_ a_2815_9447# VPWR.t1550 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X1536 VPWR.t341 VGND.t3368 VPWR.t340 VPWR.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1537 a_8745_6895# cal_itt\[1\] a_8935_6895# VGND.t1616 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1538 VPWR.t3212 a_15023_2223# trim[2].t1 VPWR.t3211 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1539 a_1830_7119# net43.t22 VGND.t2707 VGND.t2706 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1540 a_5699_9269# a_5524_9295# a_5878_9295# VGND.t748 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1541 VGND.t1837 _134_ a_13825_6031# VGND.t1836 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1542 a_12691_2527# net46 VPWR.t981 VPWR.t980 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1543 VPWR.t2786 a_9664_3689# a_9839_3615# VPWR.t2785 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1544 VGND.t1278 VPWR.t3441 VGND.t1277 VGND.t1276 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1545 VGND.t1275 VPWR.t3442 VGND.t1274 VGND.t1273 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1546 a_4349_8449# a_4131_8207# VPWR.t3277 VPWR.t3276 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1547 clknet_0_clk a_8022_7119# VGND.t836 VGND.t835 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1548 VPWR.t343 VGND.t3369 VPWR.t342 VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1549 VGND.t1758 clknet_2_0__leaf_clk a_3615_8207# VGND.t1757 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1550 VPWR.t1694 net47 a_10383_7093# VPWR.t1693 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1551 trim_val\[2\] a_14347_1439# VPWR.t3274 VPWR.t3273 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1552 net32 a_15299_3311# VGND.t2281 VGND.t2280 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1553 a_9773_3689# a_8583_3317# a_9664_3689# VGND.t2642 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1554 VGND.t491 a_15023_5487# trim[4].t5 VGND.t490 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1555 _083_ mask\[4\] a_6090_10159# VGND.t2637 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X1556 a_11352_9661# a_10405_9295# a_11244_9661# VPWR.t1843 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X1557 VGND.t2658 net49 a_14184_2767# VGND.t2657 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1558 a_13825_6031# a_13783_6183# _136_ VGND.t2673 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.195 ps=1.9 w=0.65 l=0.15
X1559 a_7355_11305# a_6909_10933# a_7259_11305# VGND.t2628 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1560 _053_ a_4815_3031# VPWR.t862 VPWR.t861 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X1561 VGND.t3118 mask\[2\] a_3840_8867# VGND.t3117 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1562 _101_ _065_.t14 VGND.t3236 VGND.t3235 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1563 VGND.t1272 VPWR.t3443 VGND.t1271 VGND.t1270 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1564 VGND.t553 a_6703_2197# trim_mask\[4\] VGND.t552 sky130_fd_pr__nfet_01v8 ad=0.209 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1565 a_8022_7119# clk.t3 VGND.t3085 VGND.t3084 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1566 clknet_2_2__leaf_clk a_8298_2767# VGND.t2416 VGND.t2415 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1567 a_14604_3017# trim_mask\[1\] VGND.t129 VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1568 VGND.t429 a_14063_7093# _134_ VGND.t428 sky130_fd_pr__nfet_01v8 ad=0.258 pd=1.45 as=0.169 ps=1.82 w=0.65 l=0.15
X1569 a_1830_10205# net43.t23 VGND.t2709 VGND.t2708 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1570 a_1276_565# net6 VGND.t1726 VGND.t1725 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1571 VGND.t1811 clknet_2_1__leaf_clk.t41 a_3431_10933# VGND.t1810 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1572 a_6983_10217# a_6633_9845# a_6888_10205# VPWR.t2808 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1573 VPWR.t1001 a_14335_4020# net49 VPWR.t1000 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1574 a_10774_9661# a_10239_9295# a_10688_9295# VPWR.t3082 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X1575 VGND.t1269 VPWR.t3444 VGND.t1268 VGND.t1237 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1576 VPWR.t1005 a_1476_7119# a_1651_7093# VPWR.t1004 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1577 a_6785_7119# a_6741_7361# a_6619_7119# VGND.t2282 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1578 a_1953_9129# a_763_8757# a_1844_9129# VGND.t82 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1579 _020_ a_6099_10633# VPWR.t1991 VPWR.t1990 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1580 a_3565_10205# a_3521_9813# a_3399_10217# VGND.t608 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1581 a_13821_7119# cal_count\[2\] VGND.t2188 VGND.t2187 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1582 a_1830_6031# net45 VGND.t2481 VGND.t2480 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1583 VGND.t2603 cal_count\[3\] a_13193_6031# VGND.t2602 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0683 ps=0.86 w=0.65 l=0.15
X1584 a_10838_2045# a_9761_1679# a_10676_1679# VPWR.t2532 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1585 VGND.t1267 VPWR.t3445 VGND.t1266 VGND.t1265 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1586 a_14281_4943# a_13091_4943# a_14172_4943# VGND.t584 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1587 VGND.t2565 _053_ _066_ VGND.t2564 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1588 a_2313_6183# mask\[0\] a_2476_6281# VPWR.t3053 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1589 a_1651_10143# net43.t24 VPWR.t2754 VPWR.t2753 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1590 VGND.t1264 VPWR.t3446 VGND.t1263 VGND.t1262 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1591 VPWR.t2643 cal_count\[3\] _105_ VPWR.t2642 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1592 _074_ a_5423_9011# VPWR.t3098 VPWR.t3097 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1593 VGND.t2315 a_455_8181# result[2].t4 VGND.t2314 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1594 VPWR.t346 VGND.t3370 VPWR.t345 VPWR.t344 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1595 a_2198_9117# net43.t25 VGND.t2711 VGND.t2710 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1596 VPWR.t2231 _060_ a_5455_4943# VPWR.t2230 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1597 a_7367_10927# net44 VPWR.t2843 VPWR.t2842 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1598 a_2450_9955# net25 a_2368_9955# VPWR.t3131 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1599 a_2689_8751# _078_ VPWR.t3108 VPWR.t3107 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X1600 a_9621_8029# _067_ VGND.t185 VGND.t184 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X1601 net12 net20.t4 VPWR.t2220 VPWR.t2219 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1602 trim[2].t0 a_15023_2223# VPWR.t3210 VPWR.t3209 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1603 VGND.t2213 _062_.t14 _064_ VGND.t2212 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1604 VPWR.t349 VGND.t3371 VPWR.t348 VPWR.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1605 VPWR.t880 _074_ a_845_7663# VPWR.t879 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1606 VGND.t1261 VPWR.t3447 VGND.t1260 VGND.t1259 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1607 _119_ a_9003_3829# VGND.t425 VGND.t424 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1608 a_6428_7119# _003_ VGND.t2057 VGND.t2056 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1609 a_5449_6031# a_4259_6031# a_5340_6031# VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1610 a_5691_7637# net51 VPWR.t1127 VPWR.t1126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1611 VPWR.t351 VGND.t3372 VPWR.t350 VPWR.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1612 VPWR.t354 VGND.t3373 VPWR.t353 VPWR.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1613 _051_.t8 a_3933_2767# VGND.t505 VGND.t504 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1614 VGND.t2633 trim_val\[2\] a_14604_2339# VGND.t173 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1615 VPWR.t2952 a_9572_2601# a_9747_2527# VPWR.t2951 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1616 a_5699_1653# a_5524_1679# a_5878_1679# VGND.t636 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1617 VGND.t3178 a_12323_4703# a_12257_4777# VGND.t3177 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1618 VPWR.t752 _106_ a_9503_4399# VPWR.t751 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1619 a_10781_5807# _092_ VGND.t2814 VGND.t2813 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1620 trim[4].t4 a_15023_5487# VGND.t489 VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X1621 a_1497_8725# a_1279_9129# VGND.t1742 VGND.t1741 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1622 VPWR.t1832 clknet_2_1__leaf_clk.t42 a_6467_9845# VPWR.t1831 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1623 a_4043_7093# a_3868_7119# a_4222_7119# VGND.t3185 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1624 VPWR.t3124 state\[1\] a_3933_2767# VPWR.t3123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1625 a_561_4405# a_395_4405# VPWR.t2226 VPWR.t2225 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1626 a_13703_4943# a_13257_4943# a_13607_4943# VGND.t1730 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1627 VPWR.t2803 _093_ a_937_4105# VPWR.t2802 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1628 _075_ a_5547_5603# a_5726_5807# VGND.t2878 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1629 clknet_2_0__leaf_clk a_2857_5461# VGND.t668 VGND.t667 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1630 VGND.t1258 VPWR.t3448 VGND.t1257 VGND.t1256 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1631 VPWR.t1287 a_14347_4917# a_14334_5309# VPWR.t1286 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1632 VGND.t280 clknet_2_2__leaf_clk a_13091_1141# VGND.t279 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1633 VPWR.t1662 a_4696_8207# a_4871_8181# VPWR.t1661 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1634 VPWR.t357 VGND.t3374 VPWR.t356 VPWR.t355 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1635 VGND.t302 a_9459_7895# _070_ VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1636 VGND.t237 net46 a_12121_3677# VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1637 a_6909_10933# a_6743_10933# VGND.t2534 VGND.t2533 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1638 VPWR.t2078 _116_ a_9719_1473# VPWR.t2077 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1639 a_3224_2601# a_2309_2229# a_2877_2197# VGND.t1 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1640 VPWR.t1741 _095_ a_2865_4460# VPWR.t1740 sky130_fd_pr__pfet_01v8_hvt ad=0.178 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X1641 VGND.t2267 net21 net13 VGND.t2266 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1642 VPWR.t2617 _050_ a_5547_5603# VPWR.t2616 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.109 ps=1.36 w=0.42 l=0.15
X1643 VGND.t1255 VPWR.t3449 VGND.t1254 VGND.t1253 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1644 VGND.t2394 net52 a_3133_11247# VGND.t2393 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1645 a_11951_2601# a_11435_2229# a_11856_2589# VGND.t1737 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1646 VPWR.t1997 a_14335_2442# net48 VPWR.t1996 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1647 a_6631_7485# net44 VPWR.t2841 VPWR.t2840 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1648 VPWR.t953 a_12691_2527# a_12678_2223# VPWR.t952 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1649 VPWR.t2037 a_11116_8983# _124_ VPWR.t2036 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X1650 a_448_6549# net22 VPWR.t3166 VPWR.t3165 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1651 VGND.t1252 VPWR.t3450 VGND.t1251 VGND.t1056 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1652 VPWR.t360 VGND.t3375 VPWR.t359 VPWR.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1653 net38 net33 VGND.t2619 VGND.t2618 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1654 VGND.t2894 a_14983_9269# _127_ VGND.t2893 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X1655 VPWR.t1320 net35 a_15023_5487# VPWR.t1319 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1656 net28 a_4687_12319# VGND.t799 VGND.t798 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1657 VPWR.t1915 clknet_2_3__leaf_clk a_10239_9295# VPWR.t1914 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1658 a_561_7119# a_395_7119# VGND.t1794 VGND.t1793 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1659 VPWR.t363 VGND.t3376 VPWR.t362 VPWR.t361 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1660 VGND.t1250 VPWR.t3451 VGND.t1249 VGND.t1173 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1661 a_4883_6397# net44 VPWR.t2839 VPWR.t2838 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1662 a_11244_9661# a_10239_9295# a_11168_9661# VPWR.t3081 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X1663 a_8912_2589# _027_ VPWR.t2744 VPWR.t2743 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1664 VGND.t719 a_1099_12533# ctlp[0].t5 VGND.t718 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1665 VPWR.t2677 trim_val\[2\] a_14686_2339# VPWR.t2676 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1666 VPWR.t366 VGND.t3377 VPWR.t365 VPWR.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1667 VPWR.t3155 clk.t4 a_8022_7119# VPWR.t3154 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1668 VGND.t1694 _103_ a_8307_4719# VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1669 VGND.t2155 a_15023_12015# trimb[2].t5 VGND.t2154 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1670 VPWR.t369 VGND.t3378 VPWR.t368 VPWR.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1671 VGND.t1248 VPWR.t3452 VGND.t1247 VGND.t1246 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1672 net43.t0 a_1467_7923# VPWR.t1259 VPWR.t1258 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1673 _007_ _082_ a_1045_9545# VPWR.t3275 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1674 VGND.t2593 a_5691_7637# net52 VGND.t2592 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1675 a_4036_8207# _017_ VPWR.t2691 VPWR.t2690 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1676 _048_.t9 a_3667_3829# VGND.t3214 VGND.t3213 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1677 a_3110_3311# a_2033_3317# a_2948_3689# VPWR.t1507 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1678 net30.t0 a_7939_3855# VPWR.t3198 VPWR.t3197 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.33 w=1 l=0.15
X1679 VGND.t263 a_14335_4020# net49 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1680 VPWR.t2273 a_15083_4659# trim[1].t0 VPWR.t2272 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1681 a_9460_6807# _062_.t15 a_9602_6614# VPWR.t2238 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X1682 VPWR.t2453 a_8298_2767# clknet_2_2__leaf_clk VPWR.t2452 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1683 clknet_2_0__leaf_clk a_2857_5461# VPWR.t1428 VPWR.t1427 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1684 VPWR.t2417 net2 a_14318_8457# VPWR.t2416 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1685 a_1835_11231# a_1660_11305# a_2014_11293# VGND.t1937 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1686 VGND.t1891 clknet_2_3__leaf_clk a_8215_9295# VGND.t1890 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1687 a_1387_8751# net43.t26 VPWR.t2756 VPWR.t2755 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1688 VPWR.t1208 _061_ a_15023_6031# VPWR.t1207 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1689 VGND.t1245 VPWR.t3453 VGND.t1244 VGND.t1243 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1690 a_13415_2442# _115_ VPWR.t934 VPWR.t933 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1691 a_5997_10927# mask\[5\] a_5915_10927# VPWR.t2498 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1692 VPWR.t1545 a_9463_8725# net47 VPWR.t1544 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1693 a_7263_7093# net44 VPWR.t2837 VPWR.t2836 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1694 clknet_0_clk a_8022_7119# VGND.t834 VGND.t833 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1695 a_5067_2045# net45 VPWR.t2518 VPWR.t2517 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1696 VGND.t3008 a_10383_7093# cal_itt\[1\] VGND.t3007 sky130_fd_pr__nfet_01v8 ad=0.209 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1697 VPWR.t372 VGND.t3379 VPWR.t371 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1698 VGND.t2290 _048_.t24 a_9084_4515# VGND.t2289 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1699 VPWR.t2334 _121_ a_4167_6575# VPWR.t2333 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1700 a_561_6031# a_395_6031# VGND.t557 VGND.t556 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1701 a_6485_8181# _076_ VPWR.t1224 VPWR.t1223 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1702 VPWR.t2194 a_455_3571# valid.t2 VPWR.t2193 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1703 a_6181_10633# mask\[4\] a_6099_10633# VPWR.t2679 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1704 a_1476_7119# a_395_7119# a_1129_7361# VPWR.t1813 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1705 VGND.t2292 _048_.t25 a_6737_4719# VGND.t2291 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X1706 VGND.t527 a_1644_12533# result[7].t2 VGND.t526 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X1707 a_3425_11721# net28 _085_ VPWR.t3141 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1708 VGND.t648 net54 a_4576_3427# VGND.t647 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1709 _012_ a_855_4105# VGND.t2005 VGND.t2004 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1710 VGND.t15 _106_ _108_ VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1711 a_2971_8457# _101_ a_3053_8207# VGND.t795 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1712 _040_ a_2092_8457# VPWR.t910 VPWR.t909 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1713 a_6485_8181# _076_ VGND.t483 VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X1714 a_1651_7093# a_1476_7119# a_1830_7119# VGND.t266 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1715 a_10787_1135# trim_val\[3\] a_10569_1109# VPWR.t795 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1716 net4.t0 a_395_591# VPWR.t3305 VPWR.t3304 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1717 VGND.t1242 VPWR.t3454 VGND.t1241 VGND.t1240 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1718 VGND.t1239 VPWR.t3455 VGND.t1238 VGND.t1237 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1719 a_9602_6614# cal_itt\[0\] VPWR.t2542 VPWR.t2541 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X1720 a_4680_6031# _034_ VPWR.t2469 VPWR.t2468 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1721 a_13557_8457# _122_ a_13142_8359# VPWR.t2094 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X1722 VGND.t1967 a_14335_2442# net48 VGND.t1966 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1723 VGND.t2713 net43.t27 a_3565_10205# VGND.t2712 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1724 VGND.t2340 _083_ _008_ VGND.t2339 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1725 VPWR.t1388 a_5524_1679# a_5699_1653# VPWR.t1387 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1726 a_11149_3017# trim_mask\[2\] VPWR.t2887 VPWR.t2886 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X1727 a_14526_4943# net46 VGND.t235 VGND.t234 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1728 VGND.t1822 _094_ a_5081_4943# VGND.t1821 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X1729 VGND.t666 a_2857_5461# clknet_2_0__leaf_clk VGND.t665 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1730 VPWR.t375 VGND.t3380 VPWR.t374 VPWR.t373 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1731 a_11394_9509# a_11244_9661# VGND.t713 VGND.t712 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X1732 VPWR.t1096 a_2857_7637# clknet_2_1__leaf_clk.t7 VPWR.t1095 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1733 VGND.t2021 a_15023_10927# trimb[0].t6 VGND.t2020 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1734 VPWR.t2483 a_448_9269# result[3].t1 VPWR.t2482 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1735 VGND.t1973 _070_ _001_ VGND.t1972 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1736 VPWR.t378 VGND.t3381 VPWR.t377 VPWR.t376 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1737 VGND.t2118 a_8298_5487# clknet_2_3__leaf_clk VGND.t2117 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1738 VGND.t2346 a_15023_12559# trimb[3].t5 VGND.t2154 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1739 VPWR.t2415 net2 _131_ VPWR.t2414 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1740 VGND.t1236 VPWR.t3456 VGND.t1235 VGND.t1234 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1741 clknet_2_0__leaf_clk a_2857_5461# VPWR.t1426 VPWR.t1425 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1742 a_6523_7119# a_6007_7119# a_6428_7119# VGND.t299 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1743 a_4674_12015# a_3597_12021# a_4512_12393# VPWR.t3020 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1744 VPWR.t3122 state\[1\] a_5087_3855# VPWR.t3121 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1745 VGND.t1744 _058_ a_14655_4399# VGND.t1743 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1746 VPWR.t2475 a_455_12533# result[6].t1 VPWR.t2474 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1747 a_8839_9661# a_8215_9295# a_8731_9295# VPWR.t1962 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1748 VGND.t359 a_2857_7637# clknet_2_1__leaf_clk.t23 VGND.t358 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1749 a_4617_4105# _096_ a_4471_4007# VPWR.t1040 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.253 ps=2.52 w=1 l=0.15
X1750 a_11691_4399# net46 VPWR.t979 VPWR.t978 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1751 VGND.t296 _098_ _099_ VGND.t295 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1752 _058_ a_10188_4105# VGND.t2866 VGND.t2865 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1753 VPWR.t2323 _048_.t26 a_9166_4515# VPWR.t2322 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1754 net46 a_10055_2767# VPWR.t1574 VPWR.t1573 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1755 VPWR.t1834 clknet_2_1__leaf_clk.t43 a_2787_9845# VPWR.t1833 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1756 a_12924_8029# a_12344_8041# VGND.t2365 VGND.t2364 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1757 VGND.t1233 VPWR.t3457 VGND.t1232 VGND.t1231 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1758 a_11141_6031# a_10975_6031# VGND.t2183 VGND.t2182 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1759 VPWR.t1772 clknet_2_0__leaf_clk a_2143_2229# VPWR.t1771 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1760 VPWR.t2581 a_5691_2741# _050_ VPWR.t2580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1761 VPWR.t1400 net54 a_4658_3427# VPWR.t1399 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1762 VGND.t1230 VPWR.t3458 VGND.t1229 VGND.t1228 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1763 VGND.t1227 VPWR.t3459 VGND.t1226 VGND.t1225 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1764 VPWR.t381 VGND.t3382 VPWR.t380 VPWR.t379 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1765 a_14083_3311# net46 VPWR.t977 VPWR.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1766 a_11967_3311# net46 VPWR.t975 VPWR.t974 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X1767 a_1007_4777# a_561_4405# a_911_4777# VGND.t1923 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1768 a_6541_12021# a_6375_12021# VPWR.t3061 VPWR.t3060 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1769 VGND.t1224 VPWR.t3460 VGND.t1223 VGND.t1152 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1770 a_13142_8359# _128_ a_13279_8207# VGND.t2949 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1771 a_4864_1679# _015_ VPWR.t1132 VPWR.t1131 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1772 a_4871_8181# a_4696_8207# a_5050_8207# VGND.t1642 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1773 clknet_0_clk a_8022_7119# VPWR.t1584 VPWR.t1583 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1774 VPWR.t384 VGND.t3383 VPWR.t383 VPWR.t382 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1775 a_1651_6005# a_1476_6031# a_1830_6031# VGND.t2767 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1776 VPWR.t387 VGND.t3384 VPWR.t386 VPWR.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1777 a_7259_11305# a_6909_10933# a_7164_11293# VPWR.t2673 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1778 mask\[3\] a_5699_9269# VGND.t438 VGND.t437 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1779 VGND.t1222 VPWR.t3461 VGND.t1221 VGND.t1220 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1780 net21 a_4167_11471# VPWR.t1981 VPWR.t1980 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1781 a_3922_8867# net24 a_3840_8867# VPWR.t3235 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1782 a_10689_2223# _104_ VPWR.t1342 VPWR.t1341 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X1783 a_10219_2045# a_9595_1679# a_10111_1679# VPWR.t2567 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X1784 a_13415_2442# _115_ VGND.t195 VGND.t194 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1785 VPWR.t3144 a_14172_1513# a_14347_1439# VPWR.t3143 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1786 a_6983_10217# a_6467_9845# a_6888_10205# VGND.t2455 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1787 VPWR.t1692 net47 a_12992_8751# VPWR.t1691 sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X1788 VPWR.t1770 clknet_2_0__leaf_clk a_4259_6031# VPWR.t1769 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1789 VPWR.t1736 a_9317_3285# a_9207_3311# VPWR.t1735 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1790 a_7460_5807# _050_ a_7210_5807# VGND.t2575 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1791 a_5340_6031# a_4259_6031# a_4993_6273# VPWR.t1045 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1792 a_11413_2767# trim_mask\[2\] a_11067_3017# VGND.t2838 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1793 valid.t1 a_455_3571# VPWR.t2192 VPWR.t2191 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1794 VPWR.t390 VGND.t3385 VPWR.t389 VPWR.t388 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1795 VGND.t2025 a_6519_3829# _089_ VGND.t2024 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1796 a_3148_4399# _099_ _014_ VPWR.t1497 sky130_fd_pr__pfet_01v8_hvt ad=0.127 pd=1.25 as=0.153 ps=1.3 w=1 l=0.15
X1797 a_1191_12393# a_745_12021# a_1095_12393# VGND.t3143 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1798 VGND.t1219 VPWR.t3462 VGND.t1218 VGND.t1217 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1799 VGND.t1813 clknet_2_1__leaf_clk.t44 a_579_12021# VGND.t1812 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1800 VGND.t1216 VPWR.t3463 VGND.t1215 VGND.t1214 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1801 VGND.t416 a_10851_1653# a_10785_1679# VGND.t415 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1802 VGND.t2924 a_13519_4007# _113_ VGND.t2923 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1803 VPWR.t2257 a_12424_3689# a_12599_3615# VPWR.t2256 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1804 trim[2].t6 a_15023_2223# VGND.t3139 VGND.t1996 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1805 VGND.t325 clknet_0_clk a_8298_2767# VGND.t324 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1806 VPWR.t393 VGND.t3386 VPWR.t392 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1807 a_10373_1679# a_10329_1921# a_10207_1679# VGND.t1906 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1808 a_12323_4703# net46 VPWR.t973 VPWR.t972 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1809 a_1660_11305# a_579_10933# a_1313_10901# VPWR.t1333 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1810 VGND.t2265 net21 a_5363_12559# VGND.t2264 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1811 _102_ net52 VPWR.t2425 VPWR.t2424 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1812 VGND.t1213 VPWR.t3464 VGND.t1212 VGND.t1211 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1813 a_5625_4943# _062_.t16 a_5537_4943# VGND.t2214 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1814 clknet_2_3__leaf_clk a_8298_5487# VPWR.t2137 VPWR.t2136 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1815 clknet_2_1__leaf_clk.t6 a_2857_7637# VPWR.t1094 VPWR.t1093 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1816 VPWR.t396 VGND.t3387 VPWR.t395 VPWR.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1817 VPWR.t3047 cal_itt\[2\] _063_.t9 VPWR.t3046 sky130_fd_pr__pfet_01v8_hvt ad=0.37 pd=1.74 as=0.135 ps=1.27 w=1 l=0.15
X1818 _075_ _051_.t15 VPWR.t2764 VPWR.t2763 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.146 ps=1.34 w=1 l=0.15
X1819 _049_ _048_.t27 VPWR.t2325 VPWR.t2324 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1820 VGND.t65 a_10005_6031# _092_ VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1821 a_4655_10071# mask\[4\] a_4801_10159# VGND.t2636 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X1822 VPWR.t1967 a_7263_7093# a_7250_7485# VPWR.t1966 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1823 a_11601_2229# a_11435_2229# VGND.t1736 VGND.t1735 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1824 VGND.t2202 _060_ a_5731_4943# VGND.t2201 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1825 VGND.t1210 VPWR.t3465 VGND.t1209 VGND.t1208 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1826 VGND.t1207 VPWR.t3466 VGND.t1206 VGND.t1205 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1827 a_3461_5193# _095_ a_3273_4943# VPWR.t1739 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.213 ps=1.42 w=1 l=0.15
X1828 a_13512_1501# _031_ VPWR.t2926 VPWR.t2925 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1829 VPWR.t399 VGND.t3388 VPWR.t398 VPWR.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1830 a_14282_7119# _130_ VGND.t2938 VGND.t2937 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.258 ps=1.45 w=0.65 l=0.15
X1831 VPWR.t402 VGND.t3389 VPWR.t401 VPWR.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1832 a_4687_12319# a_4512_12393# a_4866_12381# VGND.t2966 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1833 a_12516_2601# a_11601_2229# a_12169_2197# VGND.t407 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1834 VPWR.t405 VGND.t3390 VPWR.t404 VPWR.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1835 VPWR.t408 VGND.t3391 VPWR.t407 VPWR.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1836 VGND.t233 net46 a_11845_4765# VGND.t232 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1837 a_7758_4759# net55 a_7677_4759# VGND.t2963 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0536 ps=0.675 w=0.42 l=0.15
X1838 net55 a_7019_4407# VGND.t3201 VGND.t3200 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1839 a_9463_8725# net4.t3 VPWR.t3055 VPWR.t3054 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X1840 VGND.t832 a_8022_7119# clknet_0_clk VGND.t831 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1841 VGND.t3042 _078_ a_1579_5807# VGND.t3041 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X1842 a_6445_10383# mask\[5\] a_6099_10633# VGND.t2465 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1843 VPWR.t2701 a_448_10357# result[4].t1 VPWR.t2700 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1844 VGND.t110 _102_ a_1764_10383# VGND.t109 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1845 a_9004_3677# _033_ VGND.t1852 VGND.t1851 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1846 a_11764_3677# _025_ VPWR.t1929 VPWR.t1928 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1847 a_1822_10927# a_745_10933# a_1660_11305# VPWR.t1719 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1848 VPWR.t411 VGND.t3392 VPWR.t410 VPWR.t409 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1849 a_13880_3677# _030_ VPWR.t1625 VPWR.t1624 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1850 a_6197_12015# _074_ VPWR.t878 VPWR.t877 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1851 a_8749_3317# a_8583_3317# VGND.t2641 VGND.t2640 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1852 a_12824_7663# a_12344_8041# VPWR.t2398 VPWR.t2397 sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X1853 VPWR.t1340 _104_ a_11057_4105# VPWR.t1339 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1854 VGND.t1204 VPWR.t3467 VGND.t1203 VGND.t1202 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1855 a_1461_10357# _074_ VGND.t143 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X1856 VPWR.t3226 a_12900_7663# a_13470_7663# VPWR.t3225 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X1857 VPWR.t1582 a_8022_7119# clknet_0_clk VPWR.t1581 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1858 VPWR.t2029 a_15023_2767# trim[0].t3 VPWR.t2028 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1859 VPWR.t2908 a_3339_2767# net45 VPWR.t2907 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1860 a_14193_3285# a_13975_3689# VPWR.t997 VPWR.t996 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1861 VGND.t1201 VPWR.t3468 VGND.t1200 VGND.t1199 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1862 a_5686_9661# a_4609_9295# a_5524_9295# VPWR.t999 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1863 state\[2\] a_5699_1653# VGND.t2649 VGND.t2648 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1864 VPWR.t2007 a_2019_9055# a_2006_8751# VPWR.t2006 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1865 a_13869_1501# a_13825_1109# a_13703_1513# VGND.t1877 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1866 a_1137_5487# _074_ VPWR.t876 VPWR.t875 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1867 a_8745_6895# cal_itt\[2\] a_8495_6895# VGND.t2984 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1868 VGND.t2037 a_3817_4697# a_3751_4765# VGND.t2036 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1869 VGND.t1198 VPWR.t3469 VGND.t1197 VGND.t1009 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1870 VPWR.t1182 a_1313_10901# a_1203_10927# VPWR.t1181 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1871 VPWR.t1849 net53 a_5997_10927# VPWR.t1848 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1872 VGND.t1196 VPWR.t3470 VGND.t1195 VGND.t1194 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1873 a_8298_2767# clknet_0_clk VGND.t323 VGND.t322 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1874 net3.t0 a_395_2767# VPWR.t2031 VPWR.t2030 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1875 VPWR.t414 VGND.t3393 VPWR.t413 VPWR.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1876 VGND.t292 _086_ _011_ VGND.t291 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1877 VPWR.t3096 a_5423_9011# _074_ VPWR.t3095 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1878 _061_ a_14564_6397# VPWR.t3268 VPWR.t3267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.229 ps=1.75 w=1 l=0.15
X1879 VGND.t1193 VPWR.t3471 VGND.t1192 VGND.t1191 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1880 VGND.t199 net16 net8 VGND.t198 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1881 VGND.t2933 a_1651_4703# a_1585_4777# VGND.t2932 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1882 VPWR.t417 VGND.t3394 VPWR.t416 VPWR.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1883 VGND.t1190 VPWR.t3472 VGND.t1189 VGND.t1188 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1884 _051_.t7 a_3933_2767# VGND.t503 VGND.t502 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1885 a_14467_8751# _126_ VPWR.t813 VPWR.t812 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1886 a_10752_565# net10 VGND.t419 VGND.t418 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1887 a_3578_2589# net45 VGND.t2479 VGND.t2478 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X1888 a_14540_3689# a_13459_3317# a_14193_3285# VPWR.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X1889 VPWR.t750 _106_ a_9503_4399# VPWR.t749 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1890 mask\[6\] a_4687_11231# VPWR.t2491 VPWR.t2490 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1891 a_1173_4765# a_1129_4373# a_1007_4777# VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X1892 a_4030_7485# a_2953_7119# a_3868_7119# VPWR.t2002 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1893 VGND.t7 net40 a_15023_8751# VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1894 _006_ _081_ a_1229_8457# VPWR.t1227 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1895 VPWR.t420 VGND.t3395 VPWR.t419 VPWR.t418 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1896 VPWR.t2170 _110_.t6 a_13519_4007# VPWR.t2169 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1897 a_11583_4777# a_11067_4405# a_11488_4765# VGND.t2557 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1898 VPWR.t3252 a_12323_4703# a_12310_4399# VPWR.t3251 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1899 a_7565_12393# a_6375_12021# a_7456_12393# VGND.t3004 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1900 a_9182_10749# a_8105_10383# a_9020_10383# VPWR.t2879 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1901 VGND.t664 a_2857_5461# clknet_2_0__leaf_clk VGND.t663 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1902 VGND.t1187 VPWR.t3473 VGND.t1186 VGND.t1185 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1903 _110_.t0 a_9084_4515# VPWR.t1505 VPWR.t1504 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1904 VPWR.t423 VGND.t3396 VPWR.t422 VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1905 VGND.t1184 VPWR.t3474 VGND.t1183 VGND.t1182 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1906 _078_ a_5535_8181# VPWR.t1483 VPWR.t1482 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1907 _008_ _074_ VGND.t141 VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1908 VGND.t1181 VPWR.t3475 VGND.t1180 VGND.t1179 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1909 a_816_6031# _004_ VPWR.t1629 VPWR.t1628 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1910 VGND.t1178 VPWR.t3476 VGND.t1177 VGND.t1176 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1911 _038_ a_10699_5487# VGND.t707 VGND.t706 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1912 a_448_9269# net25 VPWR.t3130 VPWR.t3129 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X1913 trim_mask\[3\] a_9747_2527# VPWR.t1140 VPWR.t1139 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X1914 a_14099_3017# trim_val\[1\] a_13881_2741# VPWR.t911 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1915 VPWR.t1463 a_11023_5108# net50 VPWR.t1462 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1916 mask\[7\] a_1835_11231# VGND.t2086 VGND.t2085 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1917 VPWR.t2473 a_455_12533# result[6].t0 VPWR.t2472 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1918 _024_ a_10975_4105# VGND.t412 VGND.t411 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X1919 ctlp[4].t3 a_10752_12533# VGND.t2275 VGND.t2274 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X1920 VGND.t2715 net43.t28 a_1357_11293# VGND.t2714 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1921 VPWR.t1271 a_12056_6031# a_12231_6005# VPWR.t1270 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1922 VPWR.t2885 trim_mask\[2\] a_14099_1929# VPWR.t2884 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1923 VPWR.t1114 net12 a_6927_591# VPWR.t1113 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1924 a_7164_11293# _021_ VGND.t2053 VGND.t2052 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1925 a_1125_7663# _078_ VPWR.t3106 VPWR.t3105 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X1926 VGND.t3129 a_7939_3855# net30.t3 VGND.t3128 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1927 _064_ _063_.t14 a_9595_5193# VPWR.t2174 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1928 VGND.t3116 mask\[2\] a_3249_9295# VGND.t3115 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1929 a_13279_7119# _123_.t7 a_13142_7271# VGND.t1636 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X1930 VPWR.t1017 clknet_2_2__leaf_clk a_11435_2229# VPWR.t1016 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1931 calibrate a_1651_4703# VGND.t2931 VGND.t2930 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X1932 VGND.t2294 _048_.t28 _098_ VGND.t2293 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1933 a_11149_2767# trim_mask\[3\] VGND.t2077 VGND.t2076 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1934 VGND.t1175 VPWR.t3477 VGND.t1174 VGND.t1173 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1935 _048_.t8 a_3667_3829# VGND.t3212 VGND.t3211 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1936 VPWR.t2780 a_8083_8181# _002_ VPWR.t2779 sky130_fd_pr__pfet_01v8_hvt ad=0.327 pd=1.65 as=0.28 ps=2.56 w=1 l=0.15
X1937 a_10111_1679# a_9595_1679# a_10016_1679# VGND.t2530 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1938 VPWR.t1836 clknet_2_1__leaf_clk.t45 a_6375_12021# VPWR.t1835 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1939 VPWR.t1611 a_7262_5461# _062_.t2 VPWR.t1610 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1940 a_5515_6005# a_5340_6031# a_5694_6031# VGND.t2867 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X1941 VGND.t1172 VPWR.t3478 VGND.t1171 VGND.t1170 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1942 VGND.t2617 en_co_clk a_14649_6031# VGND.t2616 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1943 a_8154_11721# net27 a_8072_11721# VPWR.t1884 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1944 VGND.t1169 VPWR.t3479 VGND.t1168 VGND.t1167 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1945 a_1660_11305# a_745_10933# a_1313_10901# VGND.t1702 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1946 a_2283_4020# _097_ VPWR.t2060 VPWR.t2059 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1947 ctln[6].t5 a_6927_591# VGND.t1784 VGND.t1783 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1948 VPWR.t1424 a_2857_5461# clknet_2_0__leaf_clk VPWR.t1423 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1949 a_3133_11247# mask\[7\] a_2787_10927# VGND.t2970 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1950 a_11396_6031# _038_ VPWR.t1658 VPWR.t1657 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X1951 VGND.t2327 a_10543_2455# _027_ VGND.t2326 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1952 a_3597_12021# a_3431_12021# VPWR.t1172 VPWR.t1171 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1953 a_8636_9295# _000_ VGND.t1600 VGND.t1599 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1954 VPWR.t1768 clknet_2_0__leaf_clk a_395_6031# VPWR.t1767 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1955 VGND.t48 a_10195_1354# _032_ VGND.t47 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1956 VGND.t1166 VPWR.t3480 VGND.t1165 VGND.t1164 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1957 VGND.t468 _061_ a_15023_6031# VGND.t467 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1958 VPWR.t1189 a_3521_7361# a_3411_7485# VPWR.t1188 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X1959 net3.t1 a_395_2767# VGND.t2001 VGND.t2000 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1960 _009_ _084_ a_6197_12015# VPWR.t1185 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1961 VGND.t3164 a_448_7637# result[1].t3 VGND.t3163 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X1962 VPWR.t3128 a_4709_2773# a_4815_3031# VPWR.t3127 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1963 a_7631_12319# net44 VPWR.t2835 VPWR.t2834 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1964 VGND.t1163 VPWR.t3481 VGND.t1162 VGND.t1161 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1965 VGND.t2344 net37.t5 a_15023_9839# VGND.t2343 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X1966 VGND.t2884 a_4471_4007# _015_ VGND.t2883 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1967 a_1000_12381# _011_ VGND.t197 VGND.t196 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X1968 a_6515_8534# net2 a_6056_8359# VPWR.t2413 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X1969 clknet_2_1__leaf_clk.t5 a_2857_7637# VPWR.t1092 VPWR.t1091 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1970 VGND.t1160 VPWR.t3482 VGND.t1159 VGND.t1158 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1971 VGND.t1157 VPWR.t3483 VGND.t1156 VGND.t1155 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1972 VPWR.t2589 _057_ a_14931_591# VPWR.t2588 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1973 VPWR.t2378 a_15023_12559# trimb[3].t2 VPWR.t2377 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1974 VGND.t2309 _121_ a_4167_6575# VGND.t2308 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1975 VGND.t2777 net17 a_12631_12559# VGND.t2776 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1976 VGND.t539 a_6485_8181# a_6419_8207# VGND.t538 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1977 VGND.t1815 clknet_2_1__leaf_clk.t46 a_763_8757# VGND.t1814 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1978 ctln[5].t0 a_8767_591# VPWR.t2390 VPWR.t2389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X1979 _046_ a_2828_12131# VPWR.t2247 VPWR.t2246 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1980 VPWR.t426 VGND.t3397 VPWR.t425 VPWR.t424 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1981 VGND.t164 a_12231_6005# a_12165_6031# VGND.t163 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X1982 VPWR.t1804 a_6927_591# ctln[6].t1 VPWR.t1803 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1983 a_7262_5461# _051_.t16 VGND.t2719 VGND.t2718 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.12 ps=1.04 w=0.42 l=0.15
X1984 a_7109_11989# a_6891_12393# VGND.t2682 VGND.t2681 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X1985 VGND.t3006 _100_ a_4905_3855# VGND.t3005 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X1986 net4.t1 a_395_591# VGND.t3224 VGND.t3223 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1987 a_4677_7882# _040_ VPWR.t2722 VPWR.t2721 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1988 VGND.t2717 net43.t29 a_7613_8029# VGND.t2716 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1989 _072_ _067_ a_8761_7983# VGND.t183 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1990 a_11622_7485# a_10903_7261# a_11059_7356# VGND.t761 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1991 VGND.t2392 net52 a_3317_8207# VGND.t2391 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X1992 VGND.t549 a_12992_8751# a_13562_8751# VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X1993 a_1129_7361# a_911_7119# VPWR.t2357 VPWR.t2356 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X1994 a_14377_9545# a_14347_9480# _128_ VPWR.t1302 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X1995 VPWR.t429 VGND.t3398 VPWR.t428 VPWR.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1996 VPWR.t1448 a_4512_11305# a_4687_11231# VPWR.t1447 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1997 a_9020_10383# a_8105_10383# a_8673_10625# VGND.t2835 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1998 VPWR.t2956 cal_itt\[3\] a_7723_6807# VPWR.t2955 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1999 _122_ a_11016_6691# VPWR.t864 VPWR.t863 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X2000 a_816_4765# _012_ VGND.t2400 VGND.t2399 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2001 result[4].t0 a_448_10357# VPWR.t2699 VPWR.t2698 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2002 VPWR.t2627 a_6515_6794# _003_ VPWR.t2626 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2003 VPWR.t1318 net35 net40 VPWR.t1317 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2004 VPWR.t1913 clknet_2_3__leaf_clk a_10975_6031# VPWR.t1912 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2005 VGND.t278 clknet_2_2__leaf_clk a_13091_4943# VGND.t277 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2006 VGND.t709 a_11023_5108# net50 VGND.t708 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2007 a_8360_10383# _020_ VGND.t1964 VGND.t1963 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2008 clknet_2_1__leaf_clk.t22 a_2857_7637# VGND.t357 VGND.t356 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2009 _056_ a_14604_2339# VPWR.t1790 VPWR.t1789 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X2010 a_7456_12393# a_6541_12021# a_7109_11989# VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2011 _093_ a_4498_4373# VGND.t2898 VGND.t2897 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2012 VPWR.t2579 a_5691_2741# _050_ VPWR.t2578 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2013 VPWR.t1064 clknet_0_clk a_8298_5487# VPWR.t1063 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2014 VPWR.t432 VGND.t3399 VPWR.t431 VPWR.t430 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2015 VPWR.t1467 a_11244_9661# a_11814_9295# VPWR.t1466 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2016 VGND.t1154 VPWR.t3484 VGND.t1153 VGND.t1152 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2017 _120_ a_3273_4943# VGND.t2092 VGND.t2091 sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.127 ps=1.04 w=0.65 l=0.15
X2018 VPWR.t435 VGND.t3400 VPWR.t434 VPWR.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2019 a_3852_12381# _010_ VPWR.t2870 VPWR.t2869 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2020 VPWR.t1442 a_14471_591# ctln[2].t1 VPWR.t1441 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2021 VGND.t2041 a_5363_12559# ctlp[7].t5 VGND.t2040 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2022 VPWR.t2451 a_8298_2767# clknet_2_2__leaf_clk VPWR.t2450 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2023 a_14870_7369# cal_count\[2\] a_14788_7369# VPWR.t2214 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2024 cal_itt\[3\] a_7263_7093# VGND.t1941 VGND.t1940 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2025 VGND.t1151 VPWR.t3485 VGND.t1150 VGND.t1149 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2026 a_13607_4943# a_13257_4943# a_13512_4943# VPWR.t1748 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2027 a_10699_5487# _136_ a_10781_5807# VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2028 VPWR.t839 a_13142_7271# _037_ VPWR.t838 sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X2029 VGND.t1148 VPWR.t3486 VGND.t1147 VGND.t1146 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2030 VGND.t217 a_12691_2527# a_12625_2601# VGND.t216 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2031 a_8389_5193# _105_ a_8473_5193# VPWR.t1725 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2032 _062_.t5 a_7262_5461# a_7210_5807# VGND.t1598 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2033 net21 a_4167_11471# VGND.t1953 VGND.t1952 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2034 VPWR.t1838 clknet_2_1__leaf_clk.t47 a_6835_7669# VPWR.t1837 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2035 VPWR.t2076 a_9460_6807# _068_ VPWR.t2075 sky130_fd_pr__pfet_01v8_hvt ad=0.158 pd=1.39 as=0.26 ps=2.52 w=1 l=0.15
X2036 a_11436_9295# a_10239_9295# a_11244_9661# VGND.t3015 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2037 clknet_0_clk a_8022_7119# VGND.t830 VGND.t829 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2038 a_12056_6031# a_10975_6031# a_11709_6273# VPWR.t2208 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2039 _117_ a_9719_1473# VGND.t442 VGND.t441 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X2040 VPWR.t3014 net55 a_5166_5193# VPWR.t3013 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X2041 a_1651_6005# net45 VPWR.t2516 VPWR.t2515 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2042 a_12213_2589# a_12169_2197# a_12047_2601# VGND.t3086 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2043 a_11951_2601# a_11601_2229# a_11856_2589# VPWR.t1144 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2044 a_2283_4020# _097_ VGND.t2033 VGND.t2032 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2045 a_5502_6397# a_4425_6031# a_5340_6031# VPWR.t3160 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2046 VPWR.t2190 a_455_3571# valid.t0 VPWR.t2189 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2047 _090_ _089_ a_5931_4105# VPWR.t1749 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2048 a_1203_12015# a_579_12021# a_1095_12393# VPWR.t1308 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2049 VPWR.t438 VGND.t3401 VPWR.t437 VPWR.t436 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2050 a_6906_2355# a_7223_2465# a_7181_2589# VGND.t2368 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2051 VPWR.t2659 en_co_clk a_14564_6397# VPWR.t2658 sky130_fd_pr__pfet_01v8_hvt ad=0.229 pd=1.75 as=0.0609 ps=0.71 w=0.42 l=0.15
X2052 a_13184_9117# a_11987_8757# a_12992_8751# VGND.t2891 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2053 a_455_8181# net24 VPWR.t3234 VPWR.t3233 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2054 VGND.t2980 a_9839_3615# a_9773_3689# VGND.t2979 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2055 VPWR.t441 VGND.t3402 VPWR.t440 VPWR.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2056 VGND.t563 _091_ a_10005_6031# VGND.t562 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2057 VGND.t3138 a_15023_2223# trim[2].t5 VGND.t1994 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2058 clknet_2_2__leaf_clk a_8298_2767# VGND.t2414 VGND.t2413 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2059 _065_.t2 a_4091_5309# VGND.t2096 VGND.t2095 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2060 net20.t1 a_6191_12559# VGND.t95 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2061 VPWR.t444 VGND.t3403 VPWR.t443 VPWR.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2062 a_4993_6273# a_4775_6031# VPWR.t2782 VPWR.t2781 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2063 a_4349_8449# a_4131_8207# VGND.t3199 VGND.t3198 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2064 VGND.t2069 _122_ a_13279_8207# VGND.t2068 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.114 ps=1 w=0.65 l=0.15
X2065 VPWR.t1475 a_1099_12533# ctlp[0].t2 VPWR.t1474 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2066 VPWR.t1090 a_2857_7637# clknet_2_1__leaf_clk.t4 VPWR.t1089 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2067 a_10781_3311# trim_mask\[2\] a_10699_3311# VPWR.t2883 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2068 VGND.t2116 a_8298_5487# clknet_2_3__leaf_clk VGND.t2115 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2069 a_13715_5309# a_13091_4943# a_13607_4943# VPWR.t1328 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2070 a_9761_1679# a_9595_1679# VPWR.t2566 VPWR.t2565 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2071 VPWR.t447 VGND.t3404 VPWR.t446 VPWR.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2072 VPWR.t3031 a_4349_8449# a_4239_8573# VPWR.t3030 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2073 VGND.t2796 net44 a_6785_7119# VGND.t2795 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2074 _044_ a_8072_11721# VGND.t2177 VGND.t2176 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2075 a_9471_9269# net47 VPWR.t1690 VPWR.t1689 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2076 a_10864_9269# a_10688_9295# a_11008_9295# VGND.t154 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2077 VPWR.t1330 _041_ a_13919_8751# VPWR.t1329 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2078 VPWR.t2540 cal_itt\[0\] a_9459_7895# VPWR.t2539 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X2079 VPWR.t1168 _056_ a_15023_1679# VPWR.t1167 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2080 _060_ a_4576_3427# VPWR.t1204 VPWR.t1203 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X2081 a_8731_9295# a_8215_9295# a_8636_9295# VGND.t1933 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2082 _084_ mask\[5\] a_5998_11471# VGND.t2464 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X2083 a_2006_8751# a_929_8757# a_1844_9129# VPWR.t2767 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2084 _054_ a_7190_3855# VGND.t1922 VGND.t1921 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X2085 VPWR.t2338 a_8307_6575# _063_.t2 VPWR.t2337 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2086 a_8298_5487# clknet_0_clk VPWR.t1062 VPWR.t1061 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2087 VGND.t2230 _001_ a_11622_7485# VGND.t2229 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2088 a_5686_2045# a_4609_1679# a_5524_1679# VPWR.t2913 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2089 VPWR.t2222 net20.t5 a_6927_12559# VPWR.t2221 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2090 VPWR.t2160 mask\[3\] a_2961_9545# VPWR.t2159 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X2091 a_7916_8041# a_7001_7669# a_7569_7637# VGND.t696 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2092 a_9693_8029# cal_itt\[0\] a_9621_8029# VGND.t2508 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X2093 a_5633_9295# a_4443_9295# a_5524_9295# VGND.t1908 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2094 VGND.t3028 a_1276_565# ctln[0].t3 VGND.t3027 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2095 VPWR.t450 VGND.t3405 VPWR.t449 VPWR.t448 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2096 a_455_12533# net28 VPWR.t3140 VPWR.t3139 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2097 net2 a_15259_7637# VGND.t2612 VGND.t2611 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2098 VPWR.t2213 cal_count\[2\] a_13557_7369# VPWR.t2212 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2099 a_2313_6183# net22 VGND.t3098 VGND.t3097 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X2100 a_9043_6031# cal_itt\[0\] a_8949_6031# VGND.t2507 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2101 VPWR.t453 VGND.t3406 VPWR.t452 VPWR.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2102 a_2033_3317# a_1867_3317# VGND.t1919 VGND.t1918 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2103 clknet_0_clk a_8022_7119# VPWR.t1580 VPWR.t1579 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2104 trim[0].t2 a_15023_2767# VPWR.t2027 VPWR.t2026 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2105 VGND.t2301 clk.t5 a_8022_7119# VGND.t2300 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2106 VPWR.t3330 a_5087_3855# net54 VPWR.t3329 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2107 a_4165_10901# a_3947_11305# VPWR.t1724 VPWR.t1723 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2108 a_4801_10159# net53 VGND.t1824 VGND.t1823 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X2109 a_4696_8207# a_3781_8207# a_4349_8449# VGND.t1773 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2110 a_1677_9545# _078_ VPWR.t3104 VPWR.t3103 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2111 VPWR.t456 VGND.t3407 VPWR.t455 VPWR.t454 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2112 _063_.t4 a_8307_6575# a_8495_6895# VGND.t2312 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2113 VPWR.t3012 net55 a_7527_4631# VPWR.t3011 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X2114 _074_ a_5423_9011# VPWR.t3094 VPWR.t3093 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2115 a_12756_9117# net47 VGND.t1675 VGND.t1674 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X2116 VPWR.t3287 a_4993_6273# a_4883_6397# VPWR.t3286 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2117 VPWR.t866 a_10864_9269# a_10774_9661# VPWR.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X2118 VPWR.t459 VGND.t3408 VPWR.t458 VPWR.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2119 a_10270_4105# trim_mask\[4\] a_10188_4105# VPWR.t1905 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2120 mask\[4\] a_9195_10357# VPWR.t2807 VPWR.t2806 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2121 a_10781_5487# cal_count\[3\] VPWR.t2641 VPWR.t2640 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2122 VPWR.t1422 a_2857_5461# clknet_2_0__leaf_clk VPWR.t1421 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2123 trim[2].t4 a_15023_2223# VGND.t3137 VGND.t1992 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2124 VGND.t321 clknet_0_clk a_8298_2767# VGND.t320 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2125 VGND.t745 _099_ a_3057_4719# VGND.t744 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X2126 a_5915_10927# _101_ a_5997_11247# VGND.t794 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2127 VGND.t63 a_10005_6031# _092_ VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2128 a_13008_7663# a_12061_7669# a_12900_7663# VPWR.t1978 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X2129 VGND.t2506 cal_itt\[0\] a_8935_6895# VGND.t2505 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X2130 VPWR.t462 VGND.t3409 VPWR.t461 VPWR.t460 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2131 VGND.t1590 net34.t5 net39 VGND.t1589 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2132 VGND.t470 a_1461_10357# _023_ VGND.t469 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2133 a_8820_6005# _062_.t17 a_8949_6281# VPWR.t2239 sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X2134 VPWR.t2633 a_5691_7637# net52 VPWR.t2632 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2135 VGND.t828 a_8022_7119# clknet_0_clk VGND.t827 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2136 VGND.t1145 VPWR.t3487 VGND.t1144 VGND.t1143 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2137 a_4655_10071# mask\[3\] a_4801_9839# VPWR.t2158 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2138 VGND.t1142 VPWR.t3488 VGND.t1141 VGND.t1140 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2139 VGND.t1139 VPWR.t3489 VGND.t1138 VGND.t1137 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2140 a_11258_8790# cal_count\[0\] VPWR.t2994 VPWR.t2993 sky130_fd_pr__pfet_01v8_hvt ad=0.0767 pd=0.785 as=0.158 ps=1.39 w=0.42 l=0.15
X2141 VPWR.t2977 a_1651_4703# a_1638_4399# VPWR.t2976 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2142 a_7010_3631# trim_mask\[4\] VGND.t1883 VGND.t1882 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.172 ps=1.83 w=0.65 l=0.15
X2143 _130_ a_14788_7369# VGND.t2279 VGND.t2278 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2144 a_14702_3311# a_13625_3317# a_14540_3689# VPWR.t2305 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2145 a_12586_3311# a_11509_3317# a_12424_3689# VPWR.t2282 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2146 VGND.t1136 VPWR.t3490 VGND.t1135 VGND.t1134 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2147 a_3977_10217# a_2787_9845# a_3868_10217# VGND.t270 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2148 _101_ net51 VGND.t386 VGND.t385 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2149 _078_ a_5535_8181# VPWR.t1481 VPWR.t1480 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2150 a_855_4105# _074_ a_937_4105# VPWR.t874 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2151 a_6633_9845# a_6467_9845# VGND.t2454 VGND.t2453 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2152 VGND.t1133 VPWR.t3491 VGND.t1132 VGND.t1131 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2153 a_7527_4631# trim_mask\[0\] VPWR.t1900 VPWR.t1899 sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.142 ps=1.34 w=0.42 l=0.15
X2154 VGND.t2662 a_13881_2741# _112_ VGND.t2661 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2155 a_4970_4399# _049_ a_4886_4399# VPWR.t1193 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2156 a_14983_9269# _126_ VPWR.t811 VPWR.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X2157 net52 a_5691_7637# VGND.t2591 VGND.t2590 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2158 a_5633_1679# a_4443_1679# a_5524_1679# VGND.t1947 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2159 a_13625_3317# a_13459_3317# VPWR.t915 VPWR.t914 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2160 a_11509_3317# a_11343_3317# VPWR.t2262 VPWR.t2261 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2161 a_13257_4943# a_13091_4943# VPWR.t1327 VPWR.t1326 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2162 VGND.t1130 VPWR.t3492 VGND.t1129 VGND.t1128 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2163 VGND.t2390 net52 a_2489_7983# VGND.t2389 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2164 a_10138_5807# _064_ VGND.t1605 VGND.t1604 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X2165 a_4043_11305# a_3597_10933# a_3947_11305# VGND.t2027 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2166 a_4687_11231# net43.t30 VPWR.t1360 VPWR.t1359 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2167 VGND.t1127 VPWR.t3493 VGND.t1126 VGND.t1125 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2168 VPWR.t1060 clknet_0_clk a_2857_5461# VPWR.t1059 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2169 a_11098_6691# _065_.t15 a_11016_6691# VPWR.t3315 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2170 VGND.t231 net46 a_11753_6031# VGND.t230 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2171 VPWR.t1670 a_9471_9269# a_9458_9661# VPWR.t1669 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2172 a_8360_10383# _020_ VPWR.t1993 VPWR.t1992 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2173 net9 net17 VGND.t2775 VGND.t2774 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2174 a_4617_4105# _060_ VPWR.t2229 VPWR.t2228 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X2175 a_7091_9839# net44 VPWR.t2833 VPWR.t2832 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2176 a_14099_1929# net48 VPWR.t781 VPWR.t780 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2177 VGND.t1983 _088_ a_6737_3855# VGND.t1982 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X2178 VPWR.t1134 _090_ a_3557_5193# VPWR.t1133 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.135 ps=1.27 w=1 l=0.15
X2179 VGND.t3092 a_6210_4989# _098_ VGND.t3091 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2180 VPWR.t465 VGND.t3410 VPWR.t464 VPWR.t463 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2181 VPWR.t767 net30.t8 _104_ VPWR.t766 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2182 VPWR.t468 VGND.t3411 VPWR.t467 VPWR.t466 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2183 a_9761_1679# a_9595_1679# VGND.t2529 VGND.t2528 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2184 VPWR.t471 VGND.t3412 VPWR.t470 VPWR.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2185 a_6523_7119# a_6173_7119# a_6428_7119# VPWR.t1565 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2186 VPWR.t2040 net7 a_3063_591# VPWR.t2039 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2187 clknet_2_1__leaf_clk.t21 a_2857_7637# VGND.t355 VGND.t354 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2188 a_3947_11305# a_3431_10933# a_3852_11293# VGND.t1646 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2189 trim_val\[3\] a_10851_1653# VGND.t414 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2190 VPWR.t1214 net32 net37.t0 VPWR.t1213 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2191 a_911_7119# a_561_7119# a_816_7119# VPWR.t1002 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2192 a_8949_9537# a_8731_9295# VGND.t1800 VGND.t1799 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2193 a_10593_9295# _035_ VPWR.t1521 VPWR.t1520 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X2194 a_10676_1679# a_9595_1679# a_10329_1921# VPWR.t2564 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2195 VPWR.t473 VGND.t3413 VPWR.t472 VPWR.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2196 ctlp[5].t3 a_8820_12533# VGND.t3168 VGND.t3167 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2197 a_5221_9295# a_5177_9537# a_5055_9295# VGND.t393 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2198 VPWR.t476 VGND.t3414 VPWR.t475 VPWR.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2199 a_5455_4943# net3.t2 VPWR.t1676 VPWR.t1675 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X2200 VPWR.t479 VGND.t3415 VPWR.t478 VPWR.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2201 VPWR.t1722 a_7548_10217# a_7723_10143# VPWR.t1721 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2202 a_15289_7119# _130_ _132_ VGND.t2936 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2203 _108_ _107_ a_9503_4399# VPWR.t1681 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2204 VGND.t2794 net44 a_5037_6031# VGND.t2793 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2205 VPWR.t1122 _052_ a_7021_4105# VPWR.t1121 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2206 VGND.t2998 net4.t4 a_3339_2767# VGND.t2997 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2207 a_1313_11989# a_1095_12393# VPWR.t2669 VPWR.t2668 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2208 a_7181_2589# a_6703_2197# VGND.t551 VGND.t550 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.125 ps=1.01 w=0.42 l=0.15
X2209 a_4055_10927# net43.t31 VPWR.t1362 VPWR.t1361 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2210 a_5878_9295# net44 VGND.t2792 VGND.t2791 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2211 _072_ _071_ VPWR.t3033 VPWR.t3032 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2212 a_13869_4943# a_13825_5185# a_13703_4943# VGND.t444 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2213 a_14063_7093# a_14422_7093# a_14199_7369# VPWR.t2726 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2214 clknet_2_0__leaf_clk a_2857_5461# VPWR.t1420 VPWR.t1419 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2215 sample.t7 a_455_5747# VGND.t2526 VGND.t2525 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2216 VPWR.t2058 a_12631_12559# ctlp[3].t1 VPWR.t2057 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2217 a_10798_9295# a_10405_9295# a_10688_9295# VGND.t1819 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X2218 _121_ a_3748_6281# VPWR.t2793 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X2219 a_14377_7983# a_14335_7895# _133_ VGND.t2948 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.195 ps=1.9 w=0.65 l=0.15
X2220 a_10188_4105# trim_mask\[4\] VGND.t1881 VGND.t1880 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2221 clknet_2_2__leaf_clk a_8298_2767# VGND.t2412 VGND.t2411 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2222 VPWR.t3023 mask\[7\] a_1679_10633# VPWR.t3022 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2223 a_12900_7663# a_12061_7669# a_12924_8029# VGND.t1950 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2224 a_9369_4105# _108_ VPWR.t1531 VPWR.t1530 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2225 VPWR.t2406 _066_ a_10781_5487# VPWR.t1532 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2226 VGND.t2551 _057_ a_14931_591# VGND.t2550 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2227 VPWR.t1088 a_2857_7637# clknet_2_1__leaf_clk.t3 VPWR.t1087 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2228 VPWR.t482 VGND.t3416 VPWR.t481 VPWR.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2229 VGND.t1124 VPWR.t3494 VGND.t1123 VGND.t905 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2230 VPWR.t1473 a_1099_12533# ctlp[0].t1 VPWR.t1472 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2231 a_6631_7485# a_6007_7119# a_6523_7119# VPWR.t1036 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2232 VPWR.t2538 cal_itt\[0\] _063_.t6 VPWR.t2537 sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=2.8 as=0.135 ps=1.27 w=1 l=0.15
X2233 trim_mask\[2\] a_12691_2527# VGND.t215 VGND.t214 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2234 a_10787_1135# net50 VPWR.t1999 VPWR.t1998 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2235 VPWR.t1867 a_5363_591# ctln[7].t0 VPWR.t1866 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2236 a_9296_9295# a_8381_9295# a_8949_9537# VGND.t3227 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2237 VPWR.t3185 mask\[2\] a_3922_8867# VPWR.t3184 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2238 VPWR.t1247 a_3933_2767# _051_.t3 VPWR.t1246 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2239 a_3597_10933# a_3431_10933# VGND.t1645 VGND.t1644 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2240 a_12691_2527# a_12516_2601# a_12870_2589# VGND.t2780 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2241 VGND.t454 _049_ _094_ VGND.t453 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2242 net46 a_10055_2767# VPWR.t1572 VPWR.t1571 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2243 VPWR.t2064 a_3817_4697# a_3847_4438# VPWR.t2063 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2244 VGND.t2962 net55 _059_ VGND.t2961 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2245 VGND.t1122 VPWR.t3495 VGND.t1121 VGND.t1120 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2246 VPWR.t1390 a_7477_10901# a_7367_10927# VPWR.t1389 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2247 a_6885_8372# _076_ VGND.t481 VGND.t480 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2248 VPWR.t485 VGND.t3417 VPWR.t484 VPWR.t483 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2249 VPWR.t488 VGND.t3418 VPWR.t487 VPWR.t486 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2250 VPWR.t491 VGND.t3419 VPWR.t490 VPWR.t489 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2251 _050_ a_5691_2741# VGND.t2541 VGND.t2540 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2252 a_12153_8757# a_11987_8757# VPWR.t2936 VPWR.t2935 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2253 a_4498_4373# _090_ VGND.t399 VGND.t398 sky130_fd_pr__nfet_01v8 ad=0.123 pd=1.03 as=0.0878 ps=0.92 w=0.65 l=0.15
X2254 VGND.t1119 VPWR.t3496 VGND.t1118 VGND.t1117 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2255 _093_ a_4498_4373# VGND.t2896 VGND.t2895 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.179 ps=1.85 w=0.65 l=0.15
X2256 VPWR.t494 VGND.t3420 VPWR.t493 VPWR.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2257 a_3868_10217# a_2953_9845# a_3521_9813# VGND.t1942 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2258 VGND.t229 net46 a_10373_1679# VGND.t228 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2259 a_10043_7983# cal_itt\[0\] _069_ VGND.t2504 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X2260 VGND.t2585 a_6515_6794# _003_ VGND.t2584 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2261 a_12218_6397# a_11141_6031# a_12056_6031# VPWR.t2777 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2262 state\[1\] a_3399_2527# VPWR.t1255 VPWR.t1254 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2263 VPWR.t497 VGND.t3421 VPWR.t496 VPWR.t495 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2264 a_5221_1679# a_5177_1921# a_5055_1679# VGND.t2771 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2265 clknet_2_3__leaf_clk a_8298_5487# VPWR.t2135 VPWR.t2134 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2266 _047_ a_14972_5193# VPWR.t3307 VPWR.t3306 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X2267 a_11583_4777# a_11233_4405# a_11488_4765# VPWR.t1878 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2268 a_8389_5193# net42 a_8307_4943# VPWR.t772 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2269 a_1019_4399# net45 VPWR.t2514 VPWR.t2513 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2270 VGND.t1116 VPWR.t3497 VGND.t1115 VGND.t1114 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2271 a_11268_9295# a_10688_9295# VGND.t153 VGND.t152 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2272 a_5878_1679# net45 VGND.t2477 VGND.t2476 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2273 VGND.t2410 a_8298_2767# clknet_2_2__leaf_clk VGND.t2409 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2274 VGND.t112 _087_ _090_ VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X2275 a_4222_7119# net43.t32 VGND.t614 VGND.t613 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2276 a_12533_3689# a_11343_3317# a_12424_3689# VGND.t2237 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2277 VGND.t276 clknet_2_2__leaf_clk a_11343_3317# VGND.t275 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2278 VPWR.t2015 net38 a_15023_12015# VPWR.t2014 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2279 VPWR.t500 VGND.t3422 VPWR.t499 VPWR.t498 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2280 _005_ _080_ VGND.t2920 VGND.t2919 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2281 VGND.t826 a_8022_7119# clknet_0_clk VGND.t825 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2282 a_11067_3017# _064_ a_11149_3017# VPWR.t1619 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2283 VGND.t1113 VPWR.t3498 VGND.t1112 VGND.t1111 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2284 VGND.t3238 _065_.t16 a_3748_6281# VGND.t3237 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2285 a_13257_1141# a_13091_1141# VPWR.t1275 VPWR.t1274 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2286 VPWR.t3293 a_3667_3829# _048_.t2 VPWR.t3292 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2287 a_4866_12381# net43.t33 VGND.t616 VGND.t615 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2288 VPWR.t1032 _098_ a_7571_4943# VPWR.t1031 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2289 a_1129_7361# a_911_7119# VGND.t2329 VGND.t2328 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2290 a_7223_2465# clknet_2_2__leaf_clk VPWR.t1015 VPWR.t1014 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2291 VGND.t3245 a_15023_9839# trimb[1].t5 VGND.t3244 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2292 a_4227_8207# a_3781_8207# a_4131_8207# VGND.t1772 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2293 VPWR.t502 VGND.t3423 VPWR.t501 VPWR.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2294 VPWR.t1273 a_1129_7361# a_1019_7485# VPWR.t1272 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2295 a_11709_6273# a_11491_6031# VPWR.t2671 VPWR.t2670 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2296 VGND.t586 _041_ a_13919_8751# VGND.t585 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2297 VGND.t738 calibrate _098_ VGND.t737 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2298 a_8992_9955# net26 VGND.t162 VGND.t161 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2299 a_10975_4105# _064_ a_11057_3855# VGND.t1603 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2300 a_1203_12015# net43.t34 VPWR.t1364 VPWR.t1363 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2301 a_9681_2601# a_8491_2229# a_9572_2601# VGND.t2333 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2302 VPWR.t2495 a_7891_3617# a_7715_3285# VPWR.t2494 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X2303 a_9919_6614# _067_ a_9460_6807# VPWR.t920 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.193 ps=1.34 w=0.42 l=0.15
X2304 a_11955_3689# a_11509_3317# a_11859_3689# VGND.t2255 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2305 VGND.t2918 a_3123_3615# a_3057_3689# VGND.t2917 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2306 a_11691_4399# a_11067_4405# a_11583_4777# VPWR.t2595 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2307 VPWR.t2615 _050_ a_3891_4943# VPWR.t2614 sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.109 ps=1.36 w=0.42 l=0.15
X2308 VGND.t1756 clknet_2_0__leaf_clk a_1867_3317# VGND.t1755 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2309 VGND.t735 a_14471_12559# ctlp[2].t3 VGND.t734 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X2310 cal_itt\[0\] a_9471_9269# VGND.t1648 VGND.t1647 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.209 ps=2.02 w=0.65 l=0.15
X2311 a_13050_7637# a_12900_7663# VGND.t3152 VGND.t3151 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X2312 net8 net16 VPWR.t938 VPWR.t937 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2313 VGND.t2059 clknet_2_1__leaf_clk.t48 a_6467_9845# VGND.t2058 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2314 VGND.t1110 VPWR.t3499 VGND.t1109 VGND.t1108 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2315 a_9129_10383# a_7939_10383# a_9020_10383# VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2316 a_455_3571# net41 VGND.t2311 VGND.t2310 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X2317 a_911_10217# a_395_9845# a_816_10205# VGND.t2089 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2318 cal_itt\[2\] a_8091_7967# VGND.t1832 VGND.t1831 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2319 VGND.t1107 VPWR.t3500 VGND.t1106 VGND.t1105 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2320 VPWR.t2667 net33 a_15023_2223# VPWR.t2666 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2321 _030_ a_13183_3311# VPWR.t2693 VPWR.t2692 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2322 _025_ a_10699_3311# VPWR.t1927 VPWR.t1926 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2323 VPWR.t1058 clknet_0_clk a_8298_5487# VPWR.t1057 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2324 a_7824_11305# a_6909_10933# a_7477_10901# VGND.t2627 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2325 VPWR.t505 VGND.t3424 VPWR.t504 VPWR.t503 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2326 VPWR.t2281 a_9225_2197# a_9115_2223# VPWR.t2280 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2327 VPWR.t1983 state\[2\] a_5691_2741# VPWR.t1982 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2328 a_4043_10143# net43.t35 VPWR.t1366 VPWR.t1365 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2329 a_1476_7119# a_561_7119# a_1129_7361# VGND.t265 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2330 VPWR.t2770 a_448_6549# result[0].t0 VPWR.t2769 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2331 a_12059_2223# a_11435_2229# a_11951_2601# VPWR.t1751 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2332 VGND.t2725 net13 a_5363_591# VGND.t2724 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2333 a_8485_4943# net55 VGND.t2960 VGND.t2959 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.107 ps=0.98 w=0.65 l=0.15
X2334 a_1129_6273# a_911_6031# VGND.t1602 VGND.t1601 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2335 VPWR.t2665 net33 net38 VPWR.t2664 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2336 a_4091_5309# net3.t3 VPWR.t1678 VPWR.t1677 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X2337 a_1000_11293# _023_ VPWR.t2188 VPWR.t2187 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2338 a_8949_6281# cal_itt\[2\] VPWR.t3045 VPWR.t3044 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X2339 a_7140_2223# a_6703_2197# VPWR.t1295 VPWR.t1294 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2340 VGND.t2475 net45 a_1173_4765# VGND.t2474 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2341 VGND.t319 clknet_0_clk a_2857_5461# VGND.t318 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2342 mask\[1\] a_4871_8181# VPWR.t1734 VPWR.t1733 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2343 VPWR.t2954 cal_itt\[3\] a_8307_6575# VPWR.t2953 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2344 a_13607_4943# a_13091_4943# a_13512_4943# VGND.t583 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2345 VGND.t1104 VPWR.t3501 VGND.t1103 VGND.t1102 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2346 _022_ a_2787_10927# VGND.t1770 VGND.t1769 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2347 VPWR.t2025 a_15023_2767# trim[0].t1 VPWR.t2024 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2348 a_12077_3285# a_11859_3689# VGND.t2055 VGND.t2054 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2349 a_6173_7119# a_6007_7119# VPWR.t1035 VPWR.t1034 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2350 a_8022_7119# clk.t6 VGND.t2303 VGND.t2302 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2351 a_6099_10633# _101_ a_6181_10633# VPWR.t1549 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2352 a_14983_9269# a_15159_9269# a_15111_9295# VGND.t1765 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X2353 VPWR.t508 VGND.t3425 VPWR.t507 VPWR.t506 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2354 VPWR.t3092 a_5423_9011# _074_ VPWR.t3091 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2355 VPWR.t511 VGND.t3426 VPWR.t510 VPWR.t509 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2356 VPWR.t2449 a_8298_2767# clknet_2_2__leaf_clk VPWR.t2448 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2357 VGND.t1101 VPWR.t3502 VGND.t1100 VGND.t1099 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2358 VGND.t1098 VPWR.t3503 VGND.t1097 VGND.t1096 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2359 result[0].t2 a_448_6549# VGND.t2729 VGND.t2728 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2360 VPWR.t2176 _063_.t15 a_8473_5193# VPWR.t2175 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X2361 VGND.t61 a_10005_6031# _092_ VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2362 VGND.t1095 VPWR.t3504 VGND.t1094 VGND.t1093 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2363 VGND.t1092 VPWR.t3505 VGND.t1091 VGND.t1090 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2364 net43.t7 a_1467_7923# VGND.t525 VGND.t524 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2365 a_8298_2767# clknet_0_clk VGND.t317 VGND.t316 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2366 VPWR.t2631 a_5691_7637# net52 VPWR.t2630 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2367 a_6737_4719# _052_ a_6519_4631# VGND.t380 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2368 a_6763_5193# _050_ VPWR.t2613 VPWR.t2612 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2369 ctlp[3].t0 a_12631_12559# VPWR.t2056 VPWR.t2055 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2370 VPWR.t514 VGND.t3427 VPWR.t513 VPWR.t512 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2371 a_8912_2589# _027_ VGND.t2697 VGND.t2696 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2372 a_1476_6031# a_561_6031# a_1129_6273# VGND.t2583 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2373 _135_ net2 a_13441_6281# VPWR.t2412 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X2374 ctln[2].t0 a_14471_591# VPWR.t1440 VPWR.t1439 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2375 ctln[1].t2 a_3063_591# VGND.t38 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2376 VGND.t294 _098_ a_7571_4943# VGND.t293 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2377 a_5537_4943# net3.t4 a_5455_4943# VGND.t1655 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X2378 VPWR.t1558 a_4687_12319# a_4674_12015# VPWR.t1557 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2379 a_448_10357# net26 VPWR.t898 VPWR.t897 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2380 VPWR.t517 VGND.t3428 VPWR.t516 VPWR.t515 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2381 a_3208_7119# _016_ VPWR.t2363 VPWR.t2362 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2382 a_8657_2229# a_8491_2229# VGND.t2332 VGND.t2331 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2383 a_2601_3285# a_2383_3689# VGND.t1790 VGND.t1789 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2384 a_3521_9813# a_3303_10217# VPWR.t2960 VPWR.t2959 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2385 VGND.t1089 VPWR.t3506 VGND.t1088 VGND.t1087 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2386 VGND.t2601 cal_count\[3\] a_9125_4943# VGND.t2600 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2387 VPWR.t2086 clknet_2_1__leaf_clk.t49 a_4443_9295# VPWR.t2085 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2388 VPWR.t519 VGND.t3429 VPWR.t518 VPWR.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2389 ctlp[7].t0 a_5363_12559# VPWR.t2066 VPWR.t2065 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2390 a_9839_3615# net46 VPWR.t971 VPWR.t970 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2391 a_1099_12533# net14 VPWR.t1957 VPWR.t1956 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2392 VPWR.t521 VGND.t3430 VPWR.t520 VPWR.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2393 _059_ net55 VPWR.t3010 VPWR.t3009 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2394 VGND.t2114 a_8298_5487# clknet_2_3__leaf_clk VGND.t2113 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2395 VPWR.t524 VGND.t3431 VPWR.t523 VPWR.t522 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2396 _030_ a_13183_3311# VGND.t2647 VGND.t2646 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2397 _118_ net30.t9 VPWR.t769 VPWR.t768 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X2398 VGND.t1086 VPWR.t3507 VGND.t1085 VGND.t1084 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2399 VPWR.t527 VGND.t3432 VPWR.t526 VPWR.t525 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2400 VGND.t1083 VPWR.t3508 VGND.t1082 VGND.t1081 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2401 VGND.t788 a_9463_8725# net47 VGND.t787 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X2402 net11 net19 VPWR.t3204 VPWR.t3203 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2403 a_2953_7119# a_2787_7119# VPWR.t2874 VPWR.t2873 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2404 a_4709_2773# state\[1\] VGND.t3058 VGND.t3057 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X2405 VPWR.t530 VGND.t3433 VPWR.t529 VPWR.t528 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2406 VGND.t1080 VPWR.t3509 VGND.t1079 VGND.t1048 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2407 a_5050_8207# net44 VGND.t2790 VGND.t2789 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2408 VPWR.t533 VGND.t3434 VPWR.t532 VPWR.t531 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2409 a_3817_4697# _096_ VGND.t304 VGND.t303 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X2410 trim[0].t0 a_15023_2767# VPWR.t2023 VPWR.t2022 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2411 a_9369_4105# trim_val\[4\] a_9003_3829# VPWR.t848 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X2412 _057_ a_11292_1251# VGND.t2549 VGND.t2548 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2413 VPWR.t2823 net17 net9 VPWR.t2822 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2414 VGND.t2367 a_7223_2465# a_7184_2339# VGND.t2366 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2415 VPWR.t536 VGND.t3435 VPWR.t535 VPWR.t534 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2416 VGND.t3174 a_14249_8725# _129_ VGND.t3173 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2417 VPWR.t1955 net14 net6 VPWR.t1954 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2418 VPWR.t1712 _103_ _104_ VPWR.t1711 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2419 a_5524_9295# a_4443_9295# a_5177_9537# VPWR.t1932 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2420 VPWR.t1281 a_6485_8181# a_6515_8534# VPWR.t1280 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2421 a_745_12021# a_579_12021# VGND.t567 VGND.t566 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2422 a_448_10357# net26 VGND.t160 VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2423 VGND.t692 _028_ a_7942_2223# VGND.t691 sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2424 clknet_2_0__leaf_clk a_2857_5461# VGND.t662 VGND.t661 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X2425 a_3868_10217# a_2787_9845# a_3521_9813# VPWR.t1007 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2426 _014_ a_2865_4460# VPWR.t3039 VPWR.t3038 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.178 ps=1.4 w=1 l=0.15
X2427 clknet_2_3__leaf_clk a_8298_5487# VPWR.t2133 VPWR.t2132 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2428 _108_ _107_ a_9503_4399# VPWR.t1680 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2429 VPWR.t2790 a_4043_10143# a_4030_9839# VPWR.t2789 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2430 VGND.t1078 VPWR.t3510 VGND.t1077 VGND.t1076 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2431 VGND.t1075 VPWR.t3511 VGND.t1074 VGND.t1073 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2432 _087_ a_5455_4943# VPWR.t1973 VPWR.t1972 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X2433 VGND.t1072 VPWR.t3512 VGND.t1071 VGND.t1070 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2434 VPWR.t538 VGND.t3436 VPWR.t537 VPWR.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2435 VPWR.t1418 a_2857_5461# clknet_2_0__leaf_clk VPWR.t1417 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2436 VPWR.t2423 net52 _102_ VPWR.t2422 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2437 VGND.t353 a_2857_7637# clknet_2_1__leaf_clk.t20 VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2438 a_7459_7663# a_6835_7669# a_7351_8041# VPWR.t789 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2439 VPWR.t541 VGND.t3437 VPWR.t540 VPWR.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2440 VPWR.t2512 net45 a_6703_2197# VPWR.t2511 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2441 VPWR.t544 VGND.t3438 VPWR.t543 VPWR.t542 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2442 a_7367_10927# a_6743_10933# a_7259_11305# VPWR.t2570 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2443 net6 net14 VGND.t1928 VGND.t1927 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2444 VGND.t824 a_8022_7119# clknet_0_clk VGND.t823 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2445 ctln[0].t2 a_1276_565# VGND.t3026 VGND.t3025 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2446 VGND.t1069 VPWR.t3513 VGND.t1068 VGND.t1039 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2447 _081_ net24 VGND.t3158 VGND.t3157 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X2448 VGND.t1067 VPWR.t3514 VGND.t1066 VGND.t1065 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2449 a_11292_1251# trim_mask\[3\] VGND.t2075 VGND.t2074 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2450 a_14281_1513# a_13091_1141# a_14172_1513# VGND.t535 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2451 a_7021_4105# _049_ VPWR.t1192 VPWR.t1191 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X2452 a_7521_11293# a_7477_10901# a_7355_11305# VGND.t637 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2453 VPWR.t2992 cal_count\[0\] a_14467_8751# VPWR.t2991 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2454 VPWR.t1898 trim_mask\[0\] a_13915_4399# VPWR.t1897 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2455 trimb[2].t1 a_15023_12015# VPWR.t2182 VPWR.t2181 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2456 a_5535_8181# _077_ VPWR.t3266 VPWR.t3265 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2457 VPWR.t547 VGND.t3439 VPWR.t546 VPWR.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2458 VPWR.t3057 net4.t5 a_10055_2767# VPWR.t3056 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2459 a_2787_10927# _101_ a_2869_10927# VPWR.t1548 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2460 VGND.t1064 VPWR.t3515 VGND.t1063 VGND.t1062 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2461 VPWR.t1491 calibrate a_6822_4399# VPWR.t1119 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X2462 VGND.t2524 a_455_5747# sample.t6 VGND.t2523 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2463 VPWR.t2111 a_1835_11231# a_1822_10927# VPWR.t2110 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2464 VPWR.t2971 a_3224_2601# a_3399_2527# VPWR.t2970 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2465 a_6173_7119# a_6007_7119# VGND.t298 VGND.t297 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2466 a_11394_9509# a_11244_9661# VPWR.t1465 VPWR.t1464 sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.123 ps=1.17 w=0.84 l=0.15
X2467 a_11204_7485# a_10990_7485# VPWR.t1941 VPWR.t1940 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0703 ps=0.755 w=0.42 l=0.15
X2468 VGND.t2721 _051_.t17 a_7800_4631# VGND.t2720 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X2469 a_6566_5193# _048_.t29 a_6316_5193# VPWR.t2326 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2470 a_11709_6273# a_11491_6031# VGND.t2626 VGND.t2625 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2471 VPWR.t550 VGND.t3440 VPWR.t549 VPWR.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2472 VPWR.t553 VGND.t3441 VPWR.t552 VPWR.t551 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2473 VGND.t1061 VPWR.t3516 VGND.t1060 VGND.t1059 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2474 net46 a_10055_2767# VGND.t814 VGND.t813 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2475 VPWR.t2411 net2 a_14870_7369# VPWR.t2410 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2476 a_3303_10217# a_2787_9845# a_3208_10205# VGND.t269 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2477 VGND.t1981 a_7527_4631# _088_ VGND.t1980 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X2478 VGND.t646 net54 a_5363_4719# VGND.t645 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2479 a_13703_1513# a_13257_1141# a_13607_1513# VGND.t2772 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2480 VPWR.t1245 a_3933_2767# _051_.t2 VPWR.t1244 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2481 _050_ a_5691_2741# VGND.t2539 VGND.t2538 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2482 ctlp[2].t2 a_14471_12559# VGND.t733 VGND.t732 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2483 net27 a_7631_12319# VPWR.t1356 VPWR.t1355 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2484 a_4871_6031# a_4425_6031# a_4775_6031# VGND.t3087 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2485 a_13825_5185# a_13607_4943# VGND.t2258 VGND.t2257 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2486 VGND.t227 net46 a_12213_2589# VGND.t226 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2487 a_9664_3689# a_8749_3317# a_9317_3285# VGND.t2873 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2488 VPWR.t3102 _078_ a_5915_11721# VPWR.t3101 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X2489 a_10785_1679# a_9595_1679# a_10676_1679# VGND.t2527 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2490 VGND.t2953 a_10752_565# ctln[4].t3 VGND.t2952 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2491 VPWR.t2131 a_8298_5487# clknet_2_3__leaf_clk VPWR.t2130 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2492 a_6888_10205# _008_ VGND.t170 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2493 VGND.t1058 VPWR.t3517 VGND.t1057 VGND.t1056 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2494 VGND.t2473 net45 a_2645_3677# VGND.t2472 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2495 VPWR.t1570 a_10055_2767# net46 VPWR.t1569 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2496 VGND.t3176 a_12323_4703# trim_mask\[0\] VGND.t3175 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2497 a_12992_8751# a_11987_8757# a_12916_8751# VPWR.t2934 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X2498 VGND.t2574 _050_ a_3891_4943# VGND.t2573 sky130_fd_pr__nfet_01v8 ad=0.0924 pd=0.86 as=0.109 ps=1.36 w=0.42 l=0.15
X2499 result[2].t3 a_455_8181# VPWR.t2348 VPWR.t2347 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2500 _092_ a_10005_6031# VPWR.t803 VPWR.t802 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2501 clknet_2_1__leaf_clk.t19 a_2857_7637# VGND.t351 VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2502 a_2564_2589# _014_ VPWR.t3320 VPWR.t3319 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2503 a_5177_9537# a_4959_9295# VPWR.t825 VPWR.t824 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2504 a_13256_9117# a_13142_8725# a_13184_9117# VGND.t1833 sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X2505 VGND.t594 _104_ a_11045_3631# VGND.t593 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X2506 VPWR.t556 VGND.t3442 VPWR.t555 VPWR.t554 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2507 VPWR.t2045 a_15023_10927# trimb[0].t0 VPWR.t2044 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2508 _021_ a_5915_10927# VGND.t44 VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2509 VGND.t2060 clknet_2_1__leaf_clk.t50 a_3431_12021# VGND.t2008 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2510 VPWR.t559 VGND.t3443 VPWR.t558 VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2511 VGND.t1055 VPWR.t3518 VGND.t1054 VGND.t1024 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2512 VPWR.t562 VGND.t3444 VPWR.t561 VPWR.t560 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2513 a_6891_12393# a_6541_12021# a_6796_12381# VPWR.t793 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2514 VPWR.t2857 a_1651_10143# a_1638_9839# VPWR.t2856 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2515 VGND.t1971 _070_ a_8301_8207# VGND.t1970 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.101 ps=0.96 w=0.65 l=0.15
X2516 a_1844_9129# a_929_8757# a_1497_8725# VGND.t2727 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2517 a_9463_8725# net4.t6 VGND.t3000 VGND.t2999 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X2518 _041_ a_3840_8867# VGND.t2233 VGND.t2232 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2519 VGND.t1732 _089_ _090_ VGND.t1731 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2520 net13 net21 VPWR.t2296 VPWR.t2295 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2521 a_2953_7119# a_2787_7119# VGND.t2831 VGND.t2830 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2522 _048_.t7 a_3667_3829# VGND.t3210 VGND.t3209 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2523 a_15054_5193# trim_mask\[0\] a_14972_5193# VPWR.t1896 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2524 a_4091_4943# net3.t5 VGND.t1657 VGND.t1656 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0924 ps=0.86 w=0.42 l=0.15
X2525 sample.t5 a_455_5747# VGND.t2522 VGND.t2521 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2526 a_6090_10159# _078_ VGND.t3040 VGND.t3039 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X2527 VPWR.t1120 _052_ a_6822_4105# VPWR.t1119 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X2528 VPWR.t565 VGND.t3445 VPWR.t564 VPWR.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2529 a_14172_4943# a_13257_4943# a_13825_5185# VGND.t1729 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2530 a_13783_6183# _134_ VPWR.t1861 VPWR.t1860 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.365 ps=1.73 w=1 l=0.15
X2531 VPWR.t2805 a_9195_10357# a_9182_10749# VPWR.t2804 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2532 a_13697_4373# trim_val\[0\] VGND.t209 VGND.t208 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X2533 a_2014_11293# net43.t36 VGND.t618 VGND.t617 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2534 VGND.t1053 VPWR.t3519 VGND.t1052 VGND.t1051 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2535 _008_ _083_ a_5829_9839# VPWR.t2368 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2536 clknet_2_2__leaf_clk a_8298_2767# VGND.t2408 VGND.t2407 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2537 a_13880_3677# _030_ VGND.t1610 VGND.t1609 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2538 a_11764_3677# _025_ VGND.t1905 VGND.t1904 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2539 VGND.t1050 VPWR.t3520 VGND.t1049 VGND.t1048 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2540 a_13142_8725# a_12992_8751# VGND.t547 VGND.t546 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.6 as=0.114 ps=1.01 w=0.54 l=0.15
X2541 a_8731_9295# a_8381_9295# a_8636_9295# VPWR.t3308 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2542 a_5731_4943# _075_ a_5625_4943# VGND.t635 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X2543 VGND.t3150 a_12900_7663# a_13470_7663# VGND.t3149 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2544 a_10586_7371# a_10864_7387# a_10820_7485# VPWR.t950 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2545 a_13881_1653# trim_val\[2\] VGND.t2632 VGND.t2631 sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X2546 a_9459_7895# cal_itt\[1\] a_9693_8029# VGND.t1615 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2547 VPWR.t567 VGND.t3446 VPWR.t566 VPWR.t327 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2548 _082_ net25 VGND.t3065 VGND.t3064 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X2549 a_9889_6873# cal_itt\[0\] VPWR.t2536 VPWR.t2535 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2550 _126_ a_14236_8457# VPWR.t2594 VPWR.t2593 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X2551 VGND.t2273 a_10752_12533# ctlp[4].t2 VGND.t2272 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2552 VPWR.t570 VGND.t3447 VPWR.t569 VPWR.t568 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2553 a_5363_7369# _065_.t17 VPWR.t3317 VPWR.t3316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2554 VGND.t2296 _048_.t30 a_7460_5807# VGND.t2295 sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.04 as=0.0878 ps=0.92 w=0.65 l=0.15
X2555 VGND.t1889 clknet_2_3__leaf_clk a_10239_9295# VGND.t1888 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2556 VGND.t2084 a_1835_11231# a_1769_11305# VGND.t2083 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2557 VGND.t1999 a_15023_2767# trim[0].t7 VGND.t1998 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2558 VPWR.t573 VGND.t3448 VPWR.t572 VPWR.t571 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2559 a_7079_10217# a_6633_9845# a_6983_10217# VGND.t2765 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2560 VGND.t1047 VPWR.t3521 VGND.t1046 VGND.t1045 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2561 VGND.t3032 a_5423_9011# _074_ VGND.t3031 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2562 a_15259_7637# comp.t0 VPWR.t2119 VPWR.t2118 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.162 ps=1.33 w=1 l=0.15
X2563 a_2383_3689# a_1867_3317# a_2288_3677# VGND.t1917 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2564 VPWR.t576 VGND.t3449 VPWR.t575 VPWR.t574 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2565 a_10111_1679# a_9761_1679# a_10016_1679# VPWR.t2531 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2566 VPWR.t3279 a_7019_4407# net55 VPWR.t3278 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2567 a_10245_5193# net40 _118_ VPWR.t744 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X2568 VGND.t1044 VPWR.t3522 VGND.t1043 VGND.t1042 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2569 VPWR.t847 trim_val\[4\] a_10270_4105# VPWR.t846 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2570 net54 a_5087_3855# VGND.t3251 VGND.t3250 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X2571 VGND.t1041 VPWR.t3523 VGND.t1040 VGND.t1039 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2572 _010_ _085_ VGND.t2009 VGND.t2008 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2573 a_448_7637# net23 VPWR.t1652 VPWR.t1651 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X2574 _049_ _048_.t31 VGND.t2298 VGND.t2297 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2575 net39 net34.t6 VGND.t1592 VGND.t1591 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2576 VPWR.t2245 _046_ a_4167_11471# VPWR.t2244 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2577 VGND.t3105 a_7379_2197# a_7310_2223# VGND.t3104 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2578 VGND.t2788 net44 a_7521_11293# VGND.t2787 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2579 VGND.t1720 _095_ a_3365_4943# VGND.t1719 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X2580 VPWR.t579 VGND.t3450 VPWR.t578 VPWR.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2581 a_14981_8235# cal_count\[1\] VGND.t2171 VGND.t2170 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2582 a_5694_6031# net44 VGND.t2786 VGND.t2785 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2583 VPWR.t582 VGND.t3451 VPWR.t581 VPWR.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2584 VPWR.t584 VGND.t3452 VPWR.t583 VPWR.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2585 _080_ net23 VGND.t1632 VGND.t1631 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X2586 a_8298_5487# clknet_0_clk VPWR.t1056 VPWR.t1055 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2587 VGND.t1038 VPWR.t3524 VGND.t1037 VGND.t1036 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2588 VPWR.t1889 net15 net7 VPWR.t1888 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2589 a_2961_9295# net52 VGND.t2388 VGND.t2387 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.101 ps=0.96 w=0.65 l=0.15
X2590 VGND.t2942 cal_count\[0\] a_14565_9295# VGND.t2941 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2591 VGND.t1035 VPWR.t3525 VGND.t1034 VGND.t1033 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2592 result[7].t1 a_1644_12533# VPWR.t1269 VPWR.t1268 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2593 a_6891_12393# a_6375_12021# a_6796_12381# VGND.t3003 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2594 VGND.t1032 VPWR.t3526 VGND.t1031 VGND.t1030 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2595 VPWR.t3194 _114_ a_13307_1707# VPWR.t3193 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2596 VPWR.t2316 a_7456_12393# a_7631_12319# VPWR.t2315 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2597 a_2857_5461# clknet_0_clk VGND.t315 VGND.t314 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2598 VPWR.t892 a_10688_9295# a_10864_9269# VPWR.t891 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2599 a_13092_8029# a_11895_7669# a_12900_7663# VGND.t1912 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2600 VGND.t1700 a_12631_591# ctln[3].t3 VGND.t1699 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X2601 VGND.t402 a_9747_2527# a_9681_2601# VGND.t401 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2602 VPWR.t587 VGND.t3453 VPWR.t586 VPWR.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2603 VPWR.t2577 a_5691_2741# _050_ VPWR.t2576 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2604 a_11425_5487# _065_.t18 _066_ VPWR.t3318 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2605 VGND.t1830 a_8091_7967# a_8025_8041# VGND.t1829 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2606 a_12059_2223# net46 VPWR.t969 VPWR.t968 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2607 a_1497_8725# a_1279_9129# VPWR.t1758 VPWR.t1757 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2608 VGND.t2305 clk.t7 a_8022_7119# VGND.t2304 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2609 a_9602_6941# cal_itt\[0\] VGND.t2503 VGND.t2502 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.113 ps=1.04 w=0.42 l=0.15
X2610 VGND.t2358 a_8767_591# ctln[5].t2 VGND.t2357 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0878 ps=0.92 w=0.65 l=0.15
X2611 net24 a_2019_9055# VPWR.t2005 VPWR.t2004 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2612 VGND.t1817 a_10569_1109# _116_ VGND.t1816 sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2613 a_9269_2589# a_9225_2197# a_9103_2601# VGND.t2254 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2614 a_2491_3311# net45 VPWR.t2510 VPWR.t2509 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2615 a_1835_12319# a_1660_12393# a_2014_12381# VGND.t1614 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2616 VGND.t2061 clknet_2_1__leaf_clk.t51 a_6835_7669# VGND.t1925 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2617 VPWR.t1456 state\[0\] a_3667_3829# VPWR.t1455 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2618 a_11545_9049# cal_count\[0\] VGND.t2940 VGND.t2939 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.145 ps=1.11 w=0.42 l=0.15
X2619 VPWR.t2249 _068_ _000_ VPWR.t2248 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2620 a_12546_9129# a_12153_8757# a_12436_9129# VGND.t499 sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X2621 VPWR.t590 VGND.t3454 VPWR.t589 VPWR.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2622 clknet_2_2__leaf_clk a_8298_2767# VPWR.t2447 VPWR.t2446 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2623 VGND.t1029 VPWR.t3527 VGND.t1028 VGND.t1027 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2624 a_1007_7119# a_561_7119# a_911_7119# VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2625 VGND.t79 net31 net36 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2626 VPWR.t1200 a_12436_9129# a_12612_8725# VPWR.t1199 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2627 a_1493_11721# net29 _086_ VPWR.t2899 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2628 a_7200_3631# calibrate a_7010_3311# VGND.t736 sky130_fd_pr__nfet_01v8 ad=0.146 pd=1.1 as=0.143 ps=1.09 w=0.65 l=0.15
X2629 trimb[2].t0 a_15023_12015# VPWR.t2180 VPWR.t2179 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2630 VGND.t523 a_1467_7923# net43.t6 VGND.t522 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2631 VGND.t2380 net2 a_14236_8457# VGND.t2379 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2632 VPWR.t1513 _111_ a_12723_4943# VPWR.t1512 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X2633 VPWR.t2827 a_12516_2601# a_12691_2527# VPWR.t2826 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2634 a_10655_2932# _119_ VPWR.t2017 VPWR.t2016 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2635 a_2869_10927# mask\[6\] a_2787_10927# VPWR.t1352 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2636 VPWR.t593 VGND.t3455 VPWR.t592 VPWR.t591 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2637 VPWR.t596 VGND.t3456 VPWR.t595 VPWR.t594 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2638 VPWR.t1469 net9 a_12631_591# VPWR.t1468 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2639 VGND.t1026 VPWR.t3528 VGND.t1025 VGND.t1024 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2640 a_1769_11305# a_579_10933# a_1660_11305# VGND.t590 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2641 a_1638_4399# a_561_4405# a_1476_4777# VPWR.t1950 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2642 VGND.t2563 _053_ a_11016_6691# VGND.t2562 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2643 a_4498_4373# _092_ a_5054_4399# VPWR.t2866 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.19 ps=1.38 w=1 l=0.15
X2644 VGND.t2677 _135_ a_13825_6031# VGND.t2676 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2645 VGND.t2153 a_15023_12015# trimb[2].t4 VGND.t2152 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2646 a_1844_9129# a_763_8757# a_1497_8725# VPWR.t822 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2647 VPWR.t860 a_4815_3031# _053_ VPWR.t859 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2648 a_455_5747# net30.t10 VPWR.t771 VPWR.t770 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2649 VGND.t105 a_3116_12533# ctlp[1].t3 VGND.t104 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2650 VPWR.t599 VGND.t3457 VPWR.t598 VPWR.t597 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2651 VPWR.t602 VGND.t3458 VPWR.t601 VPWR.t600 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2652 VGND.t2784 net44 a_5221_9295# VGND.t2783 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2653 a_12344_8041# a_11895_7669# a_12249_7663# VGND.t1911 sky130_fd_pr__nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X2654 net44 a_4995_7119# VPWR.t759 VPWR.t758 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X2655 VPWR.t605 VGND.t3459 VPWR.t604 VPWR.t603 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2656 cal_count\[1\] a_13562_8751# VGND.t750 VGND.t749 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2657 a_5524_1679# a_4443_1679# a_5177_1921# VPWR.t1974 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2658 VGND.t174 trim_val\[1\] a_14604_3017# VGND.t173 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2659 a_937_4105# net1 a_855_4105# VPWR.t2013 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2660 a_12323_4703# a_12148_4777# a_12502_4765# VGND.t2338 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2661 VGND.t641 a_3388_4631# _097_ VGND.t640 sky130_fd_pr__nfet_01v8 ad=0.113 pd=1.04 as=0.169 ps=1.82 w=0.65 l=0.15
X2662 trim_val\[0\] a_14347_4917# VPWR.t1285 VPWR.t1284 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2663 a_3123_3615# net45 VPWR.t2508 VPWR.t2507 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2664 clknet_2_3__leaf_clk a_8298_5487# VGND.t2112 VGND.t2111 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2665 _040_ a_2092_8457# VGND.t172 VGND.t171 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2666 a_1019_9839# net43.t37 VPWR.t1368 VPWR.t1367 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2667 VPWR.t3043 cal_itt\[2\] a_8386_8457# VPWR.t3042 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.153 ps=1.3 w=1 l=0.15
X2668 a_12664_8029# net47 VGND.t1673 VGND.t1672 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X2669 net37.t2 net32 VGND.t472 VGND.t471 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2670 VPWR.t608 VGND.t3460 VPWR.t607 VPWR.t606 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2671 VGND.t2762 a_9195_10357# a_9129_10383# VGND.t2761 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2672 VPWR.t2605 _053_ _123_.t0 VPWR.t2604 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2673 a_1007_6031# a_561_6031# a_911_6031# VGND.t2582 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2674 a_6703_2197# a_6906_2355# VPWR.t2012 VPWR.t2011 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X2675 VPWR.t611 VGND.t3461 VPWR.t610 VPWR.t609 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2676 a_6210_4989# _051_.t18 VGND.t2723 VGND.t2722 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X2677 VGND.t660 a_2857_5461# clknet_2_0__leaf_clk VGND.t659 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2678 VPWR.t1054 clknet_0_clk a_2857_7637# VPWR.t1053 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2679 clknet_2_1__leaf_clk.t18 a_2857_7637# VGND.t349 VGND.t348 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2680 a_11856_2589# _026_ VPWR.t2471 VPWR.t2470 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2681 VGND.t1023 VPWR.t3529 VGND.t1022 VGND.t1021 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2682 a_9802_4007# _108_ VPWR.t1529 VPWR.t1528 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.162 ps=1.33 w=1 l=0.15
X2683 VPWR.t1338 _104_ a_11149_3017# VPWR.t1337 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2684 a_12077_3285# a_11859_3689# VPWR.t2082 VPWR.t2081 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X2685 a_5166_5193# _094_ a_4863_4917# VPWR.t1845 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X2686 _131_ net2 a_13821_7119# VGND.t2378 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2687 trim_mask\[1\] a_12599_3615# VPWR.t3301 VPWR.t3300 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2688 VGND.t1020 VPWR.t3530 VGND.t1019 VGND.t1018 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2689 trim_val\[1\] a_14715_3615# VPWR.t1648 VPWR.t1647 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2690 a_13349_6031# cal_count\[3\] VGND.t2599 VGND.t2598 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2691 VPWR.t614 VGND.t3462 VPWR.t613 VPWR.t612 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2692 a_6419_8207# _065_.t19 a_6056_8359# VGND.t3239 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0997 ps=0.895 w=0.42 l=0.15
X2693 VPWR.t2445 a_8298_2767# clknet_2_2__leaf_clk VPWR.t2444 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2694 VGND.t1017 VPWR.t3531 VGND.t1016 VGND.t1015 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2695 VGND.t658 a_2857_5461# clknet_2_0__leaf_clk VGND.t657 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2696 VPWR.t1198 a_2313_6183# _039_ VPWR.t1197 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.34 ps=2.68 w=1 l=0.15
X2697 a_12165_6031# a_10975_6031# a_12056_6031# VGND.t2181 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2698 VPWR.t616 VGND.t3463 VPWR.t615 VPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2699 VGND.t2463 mask\[5\] a_8072_11721# VGND.t2462 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2700 VGND.t1939 a_7263_7093# a_7197_7119# VGND.t1938 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2701 VGND.t1014 VPWR.t3532 VGND.t1013 VGND.t1012 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2702 a_1313_10901# a_1095_11305# VGND.t2834 VGND.t2833 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2703 VGND.t1011 VPWR.t3533 VGND.t1010 VGND.t1009 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2704 a_9195_3689# a_8749_3317# a_9099_3689# VGND.t2872 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2705 a_10877_7983# _063_.t16 VGND.t2147 VGND.t2146 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2706 a_11059_7356# a_10864_7387# a_11369_7119# VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.14 ps=1.1 w=0.36 l=0.15
X2707 a_14972_5193# trim_mask\[0\] VGND.t1871 VGND.t1870 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2708 _064_ _063_.t17 VGND.t2149 VGND.t2148 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2709 clknet_2_0__leaf_clk a_2857_5461# VPWR.t1416 VPWR.t1415 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2710 VGND.t158 net26 _083_ VGND.t157 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2711 net43.t5 a_1467_7923# VGND.t521 VGND.t520 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X2712 VGND.t423 a_9003_3829# _119_ VGND.t422 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2713 ctlp[6].t1 a_6927_12559# VPWR.t2267 VPWR.t2266 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2714 VPWR.t1125 net51 a_5691_7637# VPWR.t1124 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2715 a_7190_3855# _053_ a_7021_4105# VPWR.t2603 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X2716 a_561_9845# a_395_9845# VGND.t2088 VGND.t2087 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2717 a_9761_8457# _069_ a_9677_8457# VPWR.t3086 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2718 clknet_0_clk a_8022_7119# VGND.t822 VGND.t821 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2719 a_2775_9071# mask\[2\] _081_ VGND.t3114 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X2720 a_13512_1501# _031_ VGND.t2880 VGND.t2879 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2721 a_7459_7663# net43.t38 VPWR.t1370 VPWR.t1369 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2722 a_8381_9295# a_8215_9295# VPWR.t1961 VPWR.t1960 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2723 a_11587_6031# a_11141_6031# a_11491_6031# VGND.t2736 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2724 VGND.t2345 a_15023_12559# trimb[3].t4 VGND.t2152 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2725 a_13257_1141# a_13091_1141# VGND.t534 VGND.t533 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2726 VGND.t1008 VPWR.t3534 VGND.t1007 VGND.t1006 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2727 VPWR.t2099 trim_mask\[3\] a_10689_2223# VPWR.t2098 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X2728 a_12424_3689# a_11343_3317# a_12077_3285# VPWR.t2260 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2729 VPWR.t619 VGND.t3464 VPWR.t618 VPWR.t617 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2730 a_10016_1679# _032_ VPWR.t3224 VPWR.t3223 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2731 _098_ a_6210_4989# a_6316_5193# VPWR.t3163 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2732 a_10586_7371# a_10903_7261# a_10861_7119# VGND.t760 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2733 a_3947_11305# a_3597_10933# a_3852_11293# VPWR.t2053 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2734 VGND.t759 _111_ a_12723_4943# VGND.t758 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2735 a_1375_9129# a_929_8757# a_1279_9129# VGND.t2726 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2736 VGND.t2471 net45 a_5221_1679# VGND.t2470 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2737 a_10655_2932# _119_ VGND.t1989 VGND.t1988 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2738 VGND.t2110 a_8298_5487# clknet_2_3__leaf_clk VGND.t2109 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2739 a_448_9269# net25 VGND.t3063 VGND.t3062 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2740 a_13393_1707# _110_.t7 a_13307_1707# VGND.t2138 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X2741 VPWR.t906 a_7723_6807# _073_ VPWR.t905 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X2742 a_1830_4765# net45 VGND.t2469 VGND.t2468 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2743 a_14172_4943# a_13091_4943# a_13825_5185# VPWR.t1325 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2744 a_2143_7663# _101_ a_2225_7983# VGND.t793 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2745 VGND.t1782 a_6927_591# ctln[6].t4 VGND.t1781 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2746 a_7091_9839# a_6467_9845# a_6983_10217# VPWR.t2487 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2747 ctln[4].t2 a_10752_565# VGND.t2951 VGND.t2950 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2748 VPWR.t622 VGND.t3465 VPWR.t621 VPWR.t620 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2749 VGND.t274 clknet_2_2__leaf_clk a_11067_4405# VGND.t273 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2750 VPWR.t2088 clknet_2_1__leaf_clk.t52 a_579_10933# VPWR.t2087 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2751 a_8993_9295# a_8949_9537# a_8827_9295# VGND.t2656 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2752 a_10405_9295# a_10239_9295# VPWR.t3080 VPWR.t3079 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2753 _062_.t0 _048_.t32 VPWR.t2328 VPWR.t2327 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2754 VPWR.t3248 a_448_11445# result[5].t1 VPWR.t3247 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2755 a_9529_6059# _053_ a_9443_6059# VGND.t2561 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X2756 _119_ a_9003_3829# VPWR.t1160 VPWR.t1159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2757 clknet_2_2__leaf_clk a_8298_2767# VPWR.t2443 VPWR.t2442 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2758 _043_ a_8992_9955# VGND.t2672 VGND.t2671 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2759 a_10195_1354# _117_ VPWR.t1642 VPWR.t1641 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2760 clknet_2_1__leaf_clk.t2 a_2857_7637# VPWR.t1086 VPWR.t1085 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2761 VGND.t1005 VPWR.t3535 VGND.t1004 VGND.t1003 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2762 clknet_2_3__leaf_clk a_8298_5487# VPWR.t2129 VPWR.t2128 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2763 VPWR.t1925 a_13881_1653# _114_ VPWR.t1924 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2764 a_12992_8751# a_12153_8757# a_13016_9117# VGND.t498 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2765 a_3565_7119# a_3521_7361# a_3399_7119# VGND.t449 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2766 _026_ a_11067_3017# VGND.t1899 VGND.t1898 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X2767 VGND.t3208 a_3667_3829# _048_.t6 VGND.t3207 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2768 VPWR.t2962 a_3123_3615# a_3110_3311# VPWR.t2961 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2769 VPWR.t2943 a_4498_4373# _093_ VPWR.t2942 sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X2770 VPWR.t2346 a_455_8181# result[2].t2 VPWR.t2345 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2771 net20.t0 a_6191_12559# VPWR.t833 VPWR.t832 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2772 a_8091_7967# net43.t39 VPWR.t1372 VPWR.t1371 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2773 VGND.t1002 VPWR.t3536 VGND.t1001 VGND.t1000 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2774 VGND.t999 VPWR.t3537 VGND.t998 VGND.t997 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2775 VGND.t347 a_2857_7637# clknet_2_1__leaf_clk.t17 VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2776 VGND.t1626 a_14715_3615# a_14649_3689# VGND.t1625 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2777 a_11057_4105# trim_mask\[1\] a_10975_4105# VPWR.t869 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2778 a_13233_4737# _110_.t8 VGND.t2140 VGND.t2139 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2779 _045_ a_5496_12131# VGND.t1596 VGND.t1595 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X2780 a_6885_8372# _076_ VPWR.t1222 VPWR.t1221 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2781 VGND.t996 VPWR.t3538 VGND.t995 VGND.t994 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2782 a_4512_11305# a_3431_10933# a_4165_10901# VPWR.t1664 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2783 a_3317_8207# mask\[2\] a_2971_8457# VGND.t358 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2784 a_14237_3677# a_14193_3285# a_14071_3689# VGND.t2271 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2785 VPWR.t1931 a_10329_1921# a_10219_2045# VPWR.t1930 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2786 a_4863_4917# net54 VPWR.t1398 VPWR.t1397 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X2787 VGND.t820 a_8022_7119# clknet_0_clk VGND.t819 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2788 VGND.t993 VPWR.t3539 VGND.t992 VGND.t991 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2789 VPWR.t3258 a_7999_11231# a_7986_10927# VPWR.t3257 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2790 _092_ a_10005_6031# VPWR.t801 VPWR.t800 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2791 a_3208_7119# _016_ VGND.t2335 VGND.t2334 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2792 VGND.t711 a_11244_9661# a_11814_9295# VGND.t710 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2793 VGND.t3038 _078_ a_3511_11471# VGND.t3037 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X2794 a_10005_6031# _091_ VPWR.t1304 VPWR.t1303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2795 VPWR.t1013 clknet_2_2__leaf_clk a_8583_3317# VPWR.t1012 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2796 VGND.t2520 a_455_5747# sample.t4 VGND.t2519 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2797 a_1493_11721# _078_ VPWR.t3100 VPWR.t3099 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.147 ps=1.29 w=1 l=0.15
X2798 VGND.t990 VPWR.t3540 VGND.t989 VGND.t988 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2799 VPWR.t2421 net52 a_2869_10927# VPWR.t2420 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2800 VPWR.t1578 a_8022_7119# clknet_0_clk VPWR.t1577 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2801 a_14733_9545# cal_count\[0\] VPWR.t2990 VPWR.t2989 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2802 VPWR.t624 VGND.t3466 VPWR.t623 VPWR.t382 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2803 _108_ _106_ VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2804 clknet_2_3__leaf_clk a_8298_5487# VGND.t2108 VGND.t2107 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X2805 net36 net31 VGND.t77 VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2806 VGND.t2406 a_8298_2767# clknet_2_2__leaf_clk VGND.t2405 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2807 net38 net33 VPWR.t2663 VPWR.t2662 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2808 ctlp[0].t4 a_1099_12533# VGND.t717 VGND.t716 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2809 VGND.t2782 net44 a_7245_10205# VGND.t2781 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2810 a_2174_8457# mask\[1\] a_2092_8457# VPWR.t1798 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2811 a_8307_4943# _105_ a_8485_4943# VGND.t29 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0683 ps=0.86 w=0.65 l=0.15
X2812 a_10990_7485# a_10903_7261# a_10586_7371# VPWR.t1514 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.0588 ps=0.7 w=0.42 l=0.15
X2813 VPWR.t627 VGND.t3467 VPWR.t626 VPWR.t625 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2814 VPWR.t1243 a_3933_2767# _051_.t1 VPWR.t1242 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2815 a_561_9845# a_395_9845# VPWR.t2114 VPWR.t2113 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2816 a_6197_6281# _075_ VPWR.t1384 VPWR.t1383 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2817 _055_ a_14604_3017# VPWR.t858 VPWR.t857 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X2818 VPWR.t630 VGND.t3468 VPWR.t629 VPWR.t628 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2819 a_11801_4373# a_11583_4777# VGND.t2882 VGND.t2881 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2820 a_1763_9295# mask\[3\] _082_ VGND.t2134 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X2821 _000_ _068_ VGND.t2224 VGND.t2223 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2822 a_2225_7663# mask\[0\] a_2143_7663# VPWR.t3052 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2823 a_12061_7669# a_11895_7669# VPWR.t1939 VPWR.t1938 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2824 a_5081_4943# net55 VGND.t2958 VGND.t2957 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2825 a_4621_11305# a_3431_10933# a_4512_11305# VGND.t1643 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2826 VPWR.t633 VGND.t3469 VPWR.t632 VPWR.t631 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2827 VPWR.t1732 a_4871_8181# a_4858_8573# VPWR.t1731 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2828 _028_ a_7010_3311# VGND.t2452 VGND.t2451 sky130_fd_pr__nfet_01v8 ad=0.214 pd=1.96 as=0.167 ps=1.16 w=0.65 l=0.15
X2829 _017_ a_2971_8457# VPWR.t1784 VPWR.t1783 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2830 VPWR.t2097 trim_mask\[3\] a_10787_1135# VPWR.t2096 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X2831 _061_ a_14564_6397# VGND.t3190 VGND.t576 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.102 ps=0.99 w=0.65 l=0.15
X2832 a_3303_10217# a_2953_9845# a_3208_10205# VPWR.t1970 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2833 VPWR.t636 VGND.t3470 VPWR.t635 VPWR.t634 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2834 a_9957_7663# cal_itt\[1\] _069_ VPWR.t1636 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2835 a_5691_2741# state\[2\] VGND.t1957 VGND.t1956 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2836 a_5997_10927# mask\[6\] VPWR.t1351 VPWR.t1350 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X2837 a_3411_7485# net43.t40 VPWR.t1374 VPWR.t1373 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X2838 VGND.t2307 a_7715_3285# _052_ VGND.t2306 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X2839 a_3386_2223# a_2309_2229# a_3224_2601# VPWR.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2840 VGND.t987 VPWR.t3541 VGND.t986 VGND.t985 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2841 a_5699_9269# net44 VPWR.t2831 VPWR.t2830 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2842 a_3053_8457# mask\[1\] a_2971_8457# VPWR.t1797 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2843 trim[0].t6 a_15023_2767# VGND.t1997 VGND.t1996 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2844 a_10055_5487# trim_mask\[0\] VPWR.t1895 VPWR.t1894 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.147 ps=1.29 w=1 l=0.15
X2845 VPWR.t2290 a_1844_9129# a_2019_9055# VPWR.t2289 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2846 _016_ a_2143_7663# VPWR.t2920 VPWR.t2919 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2847 a_816_7119# _005_ VPWR.t2975 VPWR.t2974 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2848 VGND.t984 VPWR.t3542 VGND.t983 VGND.t982 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2849 VGND.t981 VPWR.t3543 VGND.t980 VGND.t979 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2850 a_4959_9295# a_4443_9295# a_4864_9295# VGND.t1907 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2851 VGND.t978 VPWR.t3544 VGND.t977 VGND.t976 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2852 VPWR.t1568 a_10055_2767# net46 VPWR.t1567 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2853 VGND.t487 _081_ _006_ VGND.t486 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2854 a_8091_7967# a_7916_8041# a_8270_8029# VGND.t1774 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2855 VPWR.t639 VGND.t3471 VPWR.t638 VPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2856 VPWR.t777 a_3063_591# ctln[1].t0 VPWR.t776 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2857 ctlp[1].t2 a_3116_12533# VGND.t103 VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X2858 result[2].t1 a_455_8181# VPWR.t2344 VPWR.t2343 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2859 net29 a_1835_12319# VGND.t2606 VGND.t2605 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X2860 a_13111_6031# net2 VPWR.t2409 VPWR.t2408 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X2861 VGND.t3166 a_8820_12533# ctlp[5].t2 VGND.t3165 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0878 ps=0.92 w=0.65 l=0.15
X2862 VGND.t620 net43.t41 a_1357_12381# VGND.t619 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2863 VPWR.t1627 a_4165_10901# a_4055_10927# VPWR.t1626 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2864 VGND.t975 VPWR.t3545 VGND.t974 VGND.t973 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2865 a_2309_2229# a_2143_2229# VPWR.t2382 VPWR.t2381 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2866 a_6737_3855# _048_.t33 a_6519_3829# VGND.t2299 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2867 VGND.t2220 _046_ a_4167_11471# VGND.t2219 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2868 a_12153_8757# a_11987_8757# VGND.t2890 VGND.t2889 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2869 _078_ a_5535_8181# VGND.t727 VGND.t726 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2870 a_8949_6281# cal_itt\[1\] VPWR.t1635 VPWR.t1634 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2871 a_561_4405# a_395_4405# VGND.t2199 VGND.t2198 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2872 VGND.t2003 a_4677_7882# net15 VGND.t2002 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2873 a_13279_8207# _123_.t8 a_13142_8359# VGND.t1637 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.0878 ps=0.92 w=0.65 l=0.15
X2874 VPWR.t3134 a_11394_9509# a_11352_9661# VPWR.t3133 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2875 VPWR.t1349 mask\[6\] a_3425_11721# VPWR.t1348 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X2876 a_1211_7983# mask\[1\] _080_ VGND.t1778 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X2877 a_7897_6913# _072_ VGND.t2757 VGND.t2756 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X2878 VPWR.t3136 _109_ a_13059_4631# VPWR.t3135 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2879 a_7210_5807# _050_ a_7460_5807# VGND.t2572 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2880 VPWR.t2255 _001_ a_11622_7485# VPWR.t2254 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2881 a_3411_9839# a_2787_9845# a_3303_10217# VPWR.t1006 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2882 VGND.t972 VPWR.t3546 VGND.t971 VGND.t970 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2883 VGND.t1754 clknet_2_0__leaf_clk a_4259_6031# VGND.t1753 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2884 a_1184_9117# _006_ VPWR.t3222 VPWR.t3221 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X2885 VGND.t2922 _045_ a_6191_12559# VGND.t2921 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X2886 VPWR.t1853 a_8091_7967# a_8078_7663# VPWR.t1852 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2887 VGND.t969 VPWR.t3547 VGND.t968 VGND.t967 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2888 _107_ a_5536_4399# VPWR.t1279 VPWR.t1278 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.327 ps=1.65 w=1 l=0.15
X2889 trimb[0].t5 a_15023_10927# VGND.t2019 VGND.t2018 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2890 VPWR.t3291 a_3667_3829# _048_.t1 VPWR.t3290 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2891 VGND.t966 VPWR.t3548 VGND.t965 VGND.t964 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2892 VGND.t1803 a_11545_9049# a_11479_9117# VGND.t1802 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2893 VGND.t2886 _054_ a_7939_3855# VGND.t2885 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X2894 ctlp[6].t0 a_6927_12559# VPWR.t2265 VPWR.t2264 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2895 VPWR.t2367 a_12148_4777# a_12323_4703# VPWR.t2366 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2896 a_3852_11293# _022_ VGND.t156 VGND.t155 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2897 VPWR.t1766 clknet_2_0__leaf_clk a_395_7119# VPWR.t1765 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2898 ctln[7].t5 a_5363_591# VGND.t1845 VGND.t1844 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X2899 a_1660_12393# a_579_12021# a_1313_11989# VPWR.t1307 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X2900 VGND.t2063 clknet_2_1__leaf_clk.t53 a_395_9845# VGND.t2062 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2901 VPWR.t2441 a_8298_2767# clknet_2_2__leaf_clk VPWR.t2440 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2902 VGND.t703 state\[0\] a_4973_2773# VGND.t702 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.1 as=0.0536 ps=0.675 w=0.42 l=0.15
X2903 VPWR.t2330 _048_.t34 _049_ VPWR.t2329 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2904 clknet_2_0__leaf_clk a_2857_5461# VPWR.t1414 VPWR.t1413 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2905 VPWR.t1293 a_6703_2197# trim_mask\[4\] VPWR.t1292 sky130_fd_pr__pfet_01v8_hvt ad=0.301 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X2906 a_6566_5193# calibrate a_6763_5193# VPWR.t1490 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2907 VGND.t963 VPWR.t3549 VGND.t962 VGND.t961 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2908 VPWR.t2090 clknet_2_1__leaf_clk.t54 a_6743_10933# VPWR.t2089 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2909 a_1357_11293# a_1313_10901# a_1191_11305# VGND.t443 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2910 a_12870_2589# net46 VGND.t225 VGND.t224 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X2911 VPWR.t3051 mask\[0\] a_1493_5487# VPWR.t3050 sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.29 as=0.14 ps=1.28 w=1 l=0.15
X2912 VPWR.t926 a_2877_2197# a_2767_2223# VPWR.t925 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2913 VPWR.t1118 _052_ a_6927_3311# VPWR.t1117 sky130_fd_pr__pfet_01v8_hvt ad=0.243 pd=1.49 as=0.165 ps=1.33 w=1 l=0.15
X2914 a_10383_7093# a_10586_7371# VPWR.t1312 VPWR.t1311 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.113 ps=1.38 w=0.42 l=0.15
X2915 VPWR.t854 _087_ a_5931_4105# VPWR.t853 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2916 VGND.t1955 state\[2\] a_7019_4407# VGND.t1954 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X2917 VPWR.t2821 net17 a_12631_12559# VPWR.t2820 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X2918 ctln[6].t0 a_6927_591# VPWR.t1802 VPWR.t1801 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2919 VPWR.t642 VGND.t3472 VPWR.t641 VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2920 VPWR.t2157 mask\[3\] a_2450_9955# VPWR.t2156 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2921 a_10990_7485# a_10864_7387# a_10586_7371# VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2922 a_4959_1679# a_4443_1679# a_4864_1679# VGND.t1946 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2923 VGND.t960 VPWR.t3550 VGND.t959 VGND.t958 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2924 a_9361_3677# a_9317_3285# a_9195_3689# VGND.t1716 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2925 a_7201_9813# a_6983_10217# VGND.t2362 VGND.t2361 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X2926 a_12249_7663# _037_ VPWR.t835 VPWR.t834 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X2927 a_3303_7119# a_2787_7119# a_3208_7119# VGND.t2829 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2928 a_1019_4399# a_395_4405# a_911_4777# VPWR.t2224 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X2929 cal_count\[0\] a_11814_9295# VGND.t541 VGND.t540 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2930 a_6793_8970# _076_ VPWR.t1220 VPWR.t1219 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2931 a_1651_4703# a_1476_4777# a_1830_4765# VGND.t477 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2932 VGND.t957 VPWR.t3551 VGND.t956 VGND.t955 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2933 a_11008_9295# net47 VGND.t1671 VGND.t1670 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X2934 a_7263_7093# a_7088_7119# a_7442_7119# VGND.t3205 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2935 a_2815_9447# mask\[3\] a_2961_9295# VGND.t2133 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X2936 a_1822_12015# a_745_12021# a_1660_12393# VPWR.t3219 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2937 VPWR.t645 VGND.t3473 VPWR.t644 VPWR.t643 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2938 VPWR.t648 VGND.t3474 VPWR.t647 VPWR.t646 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2939 VPWR.t651 VGND.t3475 VPWR.t650 VPWR.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2940 result[5].t0 a_448_11445# VPWR.t3246 VPWR.t3245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2941 a_4036_8207# _017_ VGND.t2645 VGND.t2644 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2942 VPWR.t654 VGND.t3476 VPWR.t653 VPWR.t652 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2943 VPWR.t2865 _092_ a_3148_4399# VPWR.t2864 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.127 ps=1.25 w=1 l=0.15
X2944 VGND.t2106 a_8298_5487# clknet_2_3__leaf_clk VGND.t2105 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2945 a_4512_11305# a_3597_10933# a_4165_10901# VGND.t2026 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2946 VGND.t954 VPWR.t3552 VGND.t953 VGND.t952 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2947 VGND.t951 VPWR.t3553 VGND.t950 VGND.t949 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2948 VPWR.t743 net39 a_15023_12559# VPWR.t742 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2949 a_4725_5487# _092_ VPWR.t2863 VPWR.t2862 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2950 a_6099_10633# _101_ a_6181_10383# VGND.t792 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X2951 VGND.t1594 net34.t7 a_15023_1135# VGND.t1593 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X2952 a_2857_5461# clknet_0_clk VGND.t313 VGND.t312 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2953 a_2857_7637# clknet_0_clk VPWR.t1052 VPWR.t1051 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2954 a_10543_2455# trim_mask\[3\] a_10689_2543# VGND.t2073 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X2955 VGND.t345 a_2857_7637# clknet_2_1__leaf_clk.t16 VGND.t344 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2956 a_1541_9117# a_1497_8725# a_1375_9129# VGND.t1990 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X2957 VGND.t603 mask\[6\] a_5496_12131# VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2958 VPWR.t2740 a_1313_11989# a_1203_12015# VPWR.t2739 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X2959 VGND.t25 a_11059_7356# a_10990_7485# VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2960 VGND.t3193 a_14347_1439# a_14281_1513# VGND.t3192 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2961 a_4471_4007# net55 a_4617_3855# VGND.t2956 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.114 ps=1 w=0.65 l=0.15
X2962 VGND.t5 net40 a_10137_4943# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.0878 ps=0.92 w=0.65 l=0.15
X2963 VPWR.t785 a_13142_8359# _036_ VPWR.t784 sky130_fd_pr__pfet_01v8_hvt ad=0.373 pd=1.75 as=0.28 ps=2.56 w=1 l=0.15
X2964 VPWR.t657 VGND.t3477 VPWR.t656 VPWR.t655 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2965 a_11116_8983# _122_ a_11258_8790# VPWR.t2093 sky130_fd_pr__pfet_01v8_hvt ad=0.193 pd=1.34 as=0.0767 ps=0.785 w=0.42 l=0.15
X2966 clknet_2_2__leaf_clk a_8298_2767# VPWR.t2439 VPWR.t2438 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2967 VPWR.t2890 a_1651_6005# a_1638_6397# VPWR.t2889 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2968 a_2489_7983# mask\[1\] a_2143_7663# VGND.t1777 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2969 VPWR.t1039 a_9459_7895# _070_ VPWR.t1038 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.26 ps=2.52 w=1 l=0.15
X2970 VGND.t421 a_9003_3829# _119_ VGND.t420 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2971 VGND.t3182 a_7999_11231# a_7933_11305# VGND.t3181 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X2972 a_7723_10143# a_7548_10217# a_7902_10205# VGND.t1703 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X2973 VGND.t2635 mask\[4\] a_8992_9955# VGND.t2634 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2974 VGND.t2739 a_8083_8181# _002_ VGND.t2738 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2975 a_1651_7093# net43.t42 VPWR.t1376 VPWR.t1375 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2976 VGND.t1843 a_5363_591# ctln[7].t4 VGND.t1842 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2977 a_995_3530# cal.t0 VPWR.t1756 VPWR.t1755 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2978 VGND.t397 _090_ a_3365_4943# VGND.t396 sky130_fd_pr__nfet_01v8 ad=0.127 pd=1.04 as=0.0878 ps=0.92 w=0.65 l=0.15
X2979 VGND.t948 VPWR.t3554 VGND.t947 VGND.t946 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2980 net19 a_8767_11471# VPWR.t2973 VPWR.t2972 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X2981 a_1184_9117# _006_ VGND.t3146 VGND.t3145 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X2982 a_9747_2527# net46 VPWR.t967 VPWR.t966 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2983 VGND.t91 net18 net10 VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X2984 VGND.t519 a_1467_7923# net43.t4 VGND.t518 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2985 VPWR.t659 VGND.t3478 VPWR.t658 VPWR.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2986 VPWR.t1764 clknet_2_0__leaf_clk a_395_4405# VPWR.t1763 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X2987 net28 a_4687_12319# VPWR.t1556 VPWR.t1555 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X2988 a_13933_6281# _135_ _136_ VPWR.t2723 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X2989 a_4266_4943# a_3891_4943# a_4175_4943# VGND.t1916 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.064 ps=0.725 w=0.42 l=0.15
X2990 a_5726_5807# _051_.t19 VGND.t3120 VGND.t3119 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.1 ps=0.985 w=0.65 l=0.15
X2991 VGND.t1752 clknet_2_0__leaf_clk a_2143_2229# VGND.t1751 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2992 VPWR.t2591 _132_ a_14335_7895# VPWR.t2590 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X2993 _051_.t6 a_3933_2767# VGND.t501 VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X2994 VGND.t945 VPWR.t3555 VGND.t944 VGND.t943 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2995 net46 a_10055_2767# VGND.t812 VGND.t811 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2996 VGND.t942 VPWR.t3556 VGND.t941 VGND.t940 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2997 a_6541_12021# a_6375_12021# VGND.t3002 VGND.t3001 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2998 ctln[3].t2 a_12631_591# VGND.t1698 VGND.t1697 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2999 VPWR.t1347 mask\[6\] a_5578_12131# VPWR.t1346 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3000 a_13915_4399# _108_ VPWR.t1527 VPWR.t1526 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3001 VGND.t939 VPWR.t3557 VGND.t938 VGND.t937 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3002 VPWR.t2629 a_5691_7637# net52 VPWR.t2628 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3003 VPWR.t662 VGND.t3479 VPWR.t661 VPWR.t660 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3004 a_12678_2223# a_11601_2229# a_12516_2601# VPWR.t1143 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3005 a_1095_11305# a_579_10933# a_1000_11293# VGND.t589 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3006 a_13693_3883# _112_ VGND.t1728 VGND.t1727 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X3007 VPWR.t1812 a_1549_6794# net14 VPWR.t1811 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3008 VGND.t936 VPWR.t3558 VGND.t935 VGND.t934 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X3009 clknet_2_3__leaf_clk a_8298_5487# VGND.t2104 VGND.t2103 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3010 a_3933_2767# state\[1\] VPWR.t3120 VPWR.t3119 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3011 VGND.t933 VPWR.t3559 VGND.t932 VGND.t931 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3012 a_455_8181# net24 VGND.t3156 VGND.t3155 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0703 ps=0.755 w=0.42 l=0.15
X3013 VGND.t1750 clknet_2_0__leaf_clk a_395_7119# VGND.t1749 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3014 clknet_2_2__leaf_clk a_8298_2767# VGND.t2404 VGND.t2403 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3015 _062_.t6 _050_ VPWR.t2611 VPWR.t2610 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3016 VGND.t930 VPWR.t3560 VGND.t929 VGND.t928 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3017 a_14334_5309# a_13257_4943# a_14172_4943# VPWR.t1747 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3018 a_7109_11989# a_6891_12393# VPWR.t2728 VPWR.t2727 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3019 VPWR.t1084 a_2857_7637# clknet_2_1__leaf_clk.t1 VPWR.t1083 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3020 VPWR.t868 trim_mask\[1\] a_14099_3017# VPWR.t867 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3021 VGND.t927 VPWR.t3561 VGND.t926 VGND.t925 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3022 VPWR.t1668 a_9471_9269# cal_itt\[0\] VPWR.t1667 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3023 VGND.t2011 net7 a_3063_591# VGND.t2010 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X3024 VPWR.t664 VGND.t3480 VPWR.t663 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3025 net52 a_5691_7637# VGND.t2589 VGND.t2588 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3026 a_12231_6005# a_12056_6031# a_12410_6031# VGND.t530 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3027 VGND.t2666 a_15023_8751# trimb[4].t5 VGND.t2665 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3028 VPWR.t2198 cal_count\[1\] a_13557_8457# VPWR.t2197 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3029 VPWR.t667 VGND.t3481 VPWR.t666 VPWR.t665 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3030 VPWR.t2241 _062_.t18 a_9595_5193# VPWR.t2240 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3031 VGND.t924 VPWR.t3562 VGND.t923 VGND.t922 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3032 VPWR.t2941 a_4498_4373# _093_ VPWR.t2940 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3033 VPWR.t670 VGND.t3482 VPWR.t669 VPWR.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3034 VPWR.t2437 a_8298_2767# clknet_2_2__leaf_clk VPWR.t2436 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3035 VPWR.t1130 a_5177_9537# a_5067_9661# VPWR.t1129 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3036 VPWR.t1082 a_2857_7637# clknet_2_1__leaf_clk.t0 VPWR.t1081 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3037 VPWR.t2127 a_8298_5487# clknet_2_3__leaf_clk VPWR.t2126 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3038 a_5515_6005# net44 VPWR.t2829 VPWR.t2828 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3039 a_855_4105# _074_ a_937_3855# VGND.t139 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3040 VGND.t921 VPWR.t3563 VGND.t920 VGND.t896 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3041 a_14733_7983# _129_ VGND.t803 VGND.t802 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.86 as=0.0878 ps=0.92 w=0.65 l=0.15
X3042 a_7351_8041# a_6835_7669# a_7256_8029# VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3043 VPWR.t2958 rstn.t0 a_395_591# VPWR.t2957 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3044 VPWR.t673 VGND.t3483 VPWR.t672 VPWR.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3045 a_13975_3689# a_13459_3317# a_13880_3677# VGND.t179 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3046 a_11859_3689# a_11343_3317# a_11764_3677# VGND.t2236 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3047 a_995_3530# cal.t1 VGND.t1740 VGND.t1739 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3048 VGND.t919 VPWR.t3564 VGND.t918 VGND.t917 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3049 a_13279_7119# cal_count\[2\] VGND.t2186 VGND.t2185 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3050 _092_ a_10005_6031# VPWR.t799 VPWR.t798 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3051 a_9003_3829# _118_ a_9369_3855# VGND.t2376 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.275 ps=1.5 w=0.65 l=0.15
X3052 a_1644_12533# net29 VGND.t2854 VGND.t2853 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3053 VGND.t3132 net19 net11 VGND.t3131 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3054 trimb[0].t4 a_15023_10927# VGND.t2017 VGND.t2016 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X3055 VPWR.t676 VGND.t3484 VPWR.t675 VPWR.t674 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3056 VPWR.t1911 clknet_2_3__leaf_clk a_11895_7669# VPWR.t1910 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3057 a_2877_2197# a_2659_2601# VGND.t695 VGND.t694 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3058 a_1638_9839# a_561_9845# a_1476_10217# VPWR.t3180 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3059 a_4131_8207# a_3615_8207# a_4036_8207# VGND.t1666 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3060 clknet_0_clk a_8022_7119# VGND.t818 VGND.t817 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3061 VGND.t1748 clknet_2_0__leaf_clk a_395_6031# VGND.t1747 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3062 a_4055_10927# a_3431_10933# a_3947_11305# VPWR.t1663 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3063 VPWR.t679 VGND.t3485 VPWR.t678 VPWR.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3064 VGND.t100 a_13142_7271# _037_ VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3065 VPWR.t682 VGND.t3486 VPWR.t681 VPWR.t680 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3066 VGND.t916 VPWR.t3565 VGND.t915 VGND.t914 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X3067 a_14377_9545# _127_ VPWR.t3148 VPWR.t3147 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3068 a_4576_3427# state\[0\] VGND.t701 VGND.t700 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3069 _108_ _106_ VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3070 _047_ a_14972_5193# VGND.t3226 VGND.t3225 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3071 mask\[7\] a_1835_11231# VPWR.t2109 VPWR.t2108 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3072 a_1129_4373# a_911_4777# VGND.t2906 VGND.t2905 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3073 a_1579_11471# mask\[7\] _086_ VGND.t2969 sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X3074 VPWR.t1847 net53 a_6181_10633# VPWR.t1846 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3075 VGND.t32 net42 a_8307_4943# VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3076 mask\[0\] a_4043_7093# VPWR.t1539 VPWR.t1538 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3077 a_9007_2601# a_8491_2229# a_8912_2589# VGND.t2330 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3078 a_816_10205# _007_ VGND.t2848 VGND.t2847 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3079 VGND.t2102 a_8298_5487# clknet_2_3__leaf_clk VGND.t2101 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3080 a_14379_6397# clknet_2_3__leaf_clk VGND.t1887 VGND.t1886 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3081 VPWR.t1138 a_9747_2527# a_9734_2223# VPWR.t1137 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3082 a_15083_4659# net32 VPWR.t1212 VPWR.t1211 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X3083 cal_count\[2\] a_13470_7663# VGND.t191 VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3084 a_5699_1653# net45 VPWR.t2506 VPWR.t2505 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3085 a_4308_4917# net54 VPWR.t1396 VPWR.t1395 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.141 ps=1.33 w=0.42 l=0.15
X3086 VGND.t913 VPWR.t3566 VGND.t912 VGND.t911 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3087 VPWR.t684 VGND.t3487 VPWR.t683 VPWR.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3088 result[3].t0 a_448_9269# VPWR.t2481 VPWR.t2480 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3089 a_12900_7663# a_11895_7669# a_12824_7663# VPWR.t1937 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X3090 _110_.t1 a_9084_4515# VGND.t752 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3091 VGND.t910 VPWR.t3567 VGND.t909 VGND.t908 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3092 VGND.t907 VPWR.t3568 VGND.t906 VGND.t905 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3093 VPWR.t1184 a_13825_5185# a_13715_5309# VPWR.t1183 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3094 VPWR.t3173 net5 a_15299_6575# VPWR.t3172 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3095 a_7524_2223# a_7310_2223# VPWR.t3232 VPWR.t3231 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0703 ps=0.755 w=0.42 l=0.15
X3096 VGND.t904 VPWR.t3569 VGND.t903 VGND.t902 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3097 VGND.t2132 mask\[3\] a_5089_10159# VGND.t2131 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3098 a_13164_8029# a_13050_7637# a_13092_8029# VGND.t3153 sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X3099 VGND.t2216 _062_.t19 a_8820_6005# VGND.t2215 sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X3100 VGND.t1879 trim_mask\[4\] a_10977_2543# VGND.t1878 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0747 ps=0.88 w=0.65 l=0.15
X3101 VPWR.t687 VGND.t3488 VPWR.t686 VPWR.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3102 state\[0\] a_3123_3615# VGND.t2916 VGND.t2915 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3103 VPWR.t3019 a_4512_12393# a_4687_12319# VPWR.t3018 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3104 a_7843_3677# _051_.t20 VGND.t3122 VGND.t3121 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X3105 a_13512_4943# _029_ VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3106 a_6888_10205# _008_ VPWR.t908 VPWR.t907 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X3107 VPWR.t2602 _053_ a_11425_5487# VPWR.t2601 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3108 a_6056_8359# net2 a_6198_8207# VGND.t2377 sky130_fd_pr__nfet_01v8 ad=0.0997 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3109 a_10329_1921# a_10111_1679# VPWR.t2784 VPWR.t2783 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3110 a_8473_5193# _053_ VPWR.t2600 VPWR.t2599 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3111 a_13257_4943# a_13091_4943# VGND.t582 VGND.t581 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3112 VPWR.t3324 a_15023_9839# trimb[1].t1 VPWR.t3323 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3113 a_13715_1135# net46 VPWR.t965 VPWR.t964 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3114 VGND.t1995 a_15023_2767# trim[0].t5 VGND.t1994 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3115 _067_ _066_ a_10055_5487# VPWR.t2405 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3116 a_7477_10901# a_7259_11305# VGND.t2284 VGND.t2283 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3117 VGND.t1885 clknet_2_3__leaf_clk a_10975_6031# VGND.t1884 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3118 a_7201_9813# a_6983_10217# VPWR.t2394 VPWR.t2393 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3119 a_1019_6397# net45 VPWR.t2504 VPWR.t2503 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3120 _050_ a_5691_2741# VPWR.t2575 VPWR.t2574 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3121 VPWR.t2342 a_455_8181# result[2].t0 VPWR.t2341 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3122 _078_ a_5535_8181# VGND.t725 VGND.t724 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3123 VPWR.t690 VGND.t3489 VPWR.t689 VPWR.t688 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3124 net34.t0 a_14931_591# VPWR.t3179 VPWR.t3178 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3125 a_3667_3829# state\[0\] VGND.t699 VGND.t698 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3126 a_6210_4989# _051_.t21 VPWR.t3192 VPWR.t3191 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3127 trimb[3].t1 a_15023_12559# VPWR.t2376 VPWR.t2375 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3128 a_14347_1439# net46 VPWR.t963 VPWR.t962 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3129 VPWR.t2062 a_13415_2442# _031_ VPWR.t2061 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3130 a_7210_5807# a_7262_5461# _062_.t4 VGND.t1597 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3131 a_5496_12131# net28 VGND.t3073 VGND.t3072 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3132 VPWR.t692 VGND.t3490 VPWR.t691 VPWR.t448 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3133 sample.t1 a_455_5747# VPWR.t2559 VPWR.t2558 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3134 VPWR.t695 VGND.t3491 VPWR.t694 VPWR.t693 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3135 VPWR.t698 VGND.t3492 VPWR.t697 VPWR.t696 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3136 VPWR.t1218 a_1476_4777# a_1651_4703# VPWR.t1217 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3137 VPWR.t3078 a_5515_6005# a_5502_6397# VPWR.t3077 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3138 a_14715_3615# net46 VPWR.t961 VPWR.t960 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3139 a_12599_3615# net46 VPWR.t959 VPWR.t958 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3140 a_6822_4399# _048_.t35 a_6519_4631# VPWR.t2010 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X3141 VPWR.t700 VGND.t3493 VPWR.t699 VPWR.t228 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3142 VGND.t901 VPWR.t3570 VGND.t900 VGND.t899 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3143 VPWR.t3008 net55 a_4617_4105# VPWR.t3007 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X3144 a_3249_9295# _101_ a_2815_9447# VGND.t791 sky130_fd_pr__nfet_01v8 ad=0.0747 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3145 a_8839_9661# net47 VPWR.t1688 VPWR.t1687 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3146 VPWR.t1454 state\[0\] a_4815_3031# VPWR.t1453 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0744 ps=0.815 w=0.42 l=0.15
X3147 a_5363_7369# net51 _101_ VPWR.t1123 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3148 a_7527_4631# a_7800_4631# a_7758_4759# VGND.t757 sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3149 VPWR.t702 VGND.t3494 VPWR.t701 VPWR.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3150 a_7548_10217# a_6467_9845# a_7201_9813# VPWR.t2486 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3151 VPWR.t2710 a_15023_8751# trimb[4].t0 VPWR.t2709 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3152 a_448_6549# net22 VGND.t3096 VGND.t3095 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3153 _004_ _079_ a_1137_5487# VPWR.t3162 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3154 a_2092_8457# mask\[1\] VGND.t1776 VGND.t1775 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3155 a_12520_7637# a_12344_8041# a_12664_8029# VGND.t2363 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3156 _076_ _075_ VGND.t634 VGND.t633 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3157 VGND.t272 clknet_2_2__leaf_clk a_11435_2229# VGND.t271 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3158 VPWR.t815 net31 a_15023_2767# VPWR.t814 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3159 _053_ a_4815_3031# VGND.t120 VGND.t119 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.127 ps=1.1 w=0.65 l=0.15
X3160 a_10699_3311# _064_ a_10781_3311# VPWR.t1618 sky130_fd_pr__pfet_01v8_hvt ad=0.253 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3161 VPWR.t1412 a_2857_5461# clknet_2_0__leaf_clk VPWR.t1411 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3162 a_2383_3689# a_2033_3317# a_2288_3677# VPWR.t1506 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3163 a_6793_8970# _076_ VGND.t479 VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3164 VGND.t898 VPWR.t3571 VGND.t897 VGND.t896 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3165 VPWR.t1525 a_9296_9295# a_9471_9269# VPWR.t1524 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3166 a_9459_7895# cal_itt\[1\] VPWR.t1633 VPWR.t1632 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3167 a_7320_3631# _049_ a_7200_3631# VGND.t452 sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.146 ps=1.1 w=0.65 l=0.15
X3168 VGND.t2151 _063_.t18 a_8745_4943# VGND.t2150 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.965 as=0.107 ps=0.98 w=0.65 l=0.15
X3169 VGND.t2065 clknet_2_1__leaf_clk.t55 a_6375_12021# VGND.t2064 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3170 VPWR.t3006 a_8820_6005# _071_ VPWR.t3005 sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X3171 ctlp[7].t4 a_5363_12559# VGND.t2039 VGND.t2038 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3172 trim[0].t4 a_15023_2767# VGND.t1993 VGND.t1992 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0703 ps=0.755 w=0.42 l=0.15
X3173 a_8072_11721# net27 VGND.t1861 VGND.t1860 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3174 VGND.t2680 a_14422_7093# a_14063_7093# VGND.t2679 sky130_fd_pr__nfet_01v8 ad=0.136 pd=1.1 as=0.0878 ps=0.92 w=0.65 l=0.15
X3175 _063_.t8 cal_itt\[2\] VPWR.t3041 VPWR.t3040 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3176 _121_ a_3748_6281# VGND.t2751 VGND.t2750 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3177 VGND.t223 net46 a_13869_1501# VGND.t222 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3178 a_3333_2601# a_2143_2229# a_3224_2601# VGND.t2349 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3179 a_5537_4105# _060_ net41 VPWR.t2227 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3180 _074_ a_5423_9011# VGND.t3030 VGND.t3029 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.122 ps=1.42 w=0.42 l=0.15
X3181 VPWR.t705 VGND.t3495 VPWR.t704 VPWR.t703 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3182 VPWR.t1782 a_15159_9269# a_14983_9269# VPWR.t1781 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X3183 VPWR.t708 VGND.t3496 VPWR.t707 VPWR.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3184 VGND.t2571 _050_ _098_ VGND.t2570 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3185 VPWR.t711 VGND.t3497 VPWR.t710 VPWR.t709 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3186 a_3597_12021# a_3431_12021# VGND.t434 VGND.t135 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3187 VGND.t3082 _127_ a_14347_9480# VGND.t3081 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3188 net45 a_3339_2767# VPWR.t2906 VPWR.t2905 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.33 w=1 l=0.15
X3189 VGND.t575 net35 net40 VGND.t574 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3190 VPWR.t714 VGND.t3498 VPWR.t713 VPWR.t712 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X3191 VGND.t2194 net20.t6 net12 VGND.t2193 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3192 VGND.t895 VPWR.t3572 VGND.t894 VGND.t893 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3193 VPWR.t2813 a_10676_1679# a_10851_1653# VPWR.t2812 sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3194 VPWR.t3083 _131_ _132_ VPWR.t2654 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3195 VPWR.t2294 net21 net13 VPWR.t2293 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3196 VGND.t622 net43.t43 a_4209_11293# VGND.t621 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3197 VGND.t573 net35 a_15023_5487# VGND.t572 sky130_fd_pr__nfet_01v8 ad=0.0703 pd=0.755 as=0.111 ps=1.37 w=0.42 l=0.15
X3198 VGND.t2035 a_13415_2442# _031_ VGND.t2034 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3199 a_14981_4020# _047_ VPWR.t1887 VPWR.t1886 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3200 a_7527_4631# a_7800_4631# VPWR.t1511 VPWR.t1510 sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3201 a_4165_11989# a_3947_12393# VPWR.t1206 VPWR.t1205 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3202 a_8636_9295# _000_ VPWR.t1615 VPWR.t1614 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X3203 a_2755_2601# a_2309_2229# a_2659_2601# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3204 a_2491_3311# a_1867_3317# a_2383_3689# VPWR.t1944 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3205 a_6822_4105# _088_ a_6519_3829# VPWR.t2010 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X3206 net17 a_11803_10383# VPWR.t2675 VPWR.t2674 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3207 VGND.t1977 a_2019_9055# a_1953_9129# VGND.t1976 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3208 a_12341_8751# _036_ VPWR.t2730 VPWR.t2729 sky130_fd_pr__pfet_01v8_hvt ad=0.125 pd=1.17 as=0.218 ps=2.2 w=0.84 l=0.15
X3209 a_7999_11231# a_7824_11305# a_8178_11293# VGND.t1965 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3210 VPWR.t2939 a_14983_9269# _127_ VPWR.t2938 sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X3211 VPWR.t2396 a_12344_8041# a_12520_7637# VPWR.t2395 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3212 a_1129_4373# a_911_4777# VPWR.t2950 VPWR.t2949 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3213 VPWR.t717 VGND.t3499 VPWR.t716 VPWR.t715 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3214 _115_ a_13307_1707# VGND.t193 VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X3215 VPWR.t2121 a_4091_5309# _065_.t0 VPWR.t2120 sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3216 a_6741_7361# a_6523_7119# VGND.t2342 VGND.t2341 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3217 VGND.t3056 state\[1\] a_3933_2767# VGND.t3055 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3218 VGND.t2247 a_15083_4659# trim[1].t4 VGND.t2246 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3219 VGND.t2760 _093_ a_1201_3855# VGND.t2759 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.114 ps=1 w=0.65 l=0.15
X3220 a_6181_10633# mask\[5\] VPWR.t2497 VPWR.t2496 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X3221 a_13607_1513# a_13091_1141# a_13512_1501# VGND.t532 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3222 net10 net18 VGND.t89 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3223 net33 a_15023_1679# VGND.t2047 VGND.t2046 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3224 a_12169_2197# a_11951_2601# VGND.t189 VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3225 a_8935_6895# cal_itt\[0\] VGND.t2501 VGND.t2500 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3226 VGND.t2852 a_9889_6873# a_9823_6941# VGND.t2851 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3227 VPWR.t3272 a_14347_1439# a_14334_1135# VPWR.t3271 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3228 VGND.t1859 net27 _084_ VGND.t1858 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3229 clknet_2_0__leaf_clk a_2857_5461# VPWR.t1410 VPWR.t1409 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X3230 a_3208_10205# _018_ VGND.t1588 VGND.t1587 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3231 VGND.t892 VPWR.t3573 VGND.t891 VGND.t890 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3232 clknet_2_3__leaf_clk a_8298_5487# VPWR.t2125 VPWR.t2124 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3233 clknet_2_0__leaf_clk a_2857_5461# VGND.t656 VGND.t655 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3234 a_1129_9813# a_911_10217# VGND.t2770 VGND.t2769 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3235 a_4775_6031# a_4259_6031# a_4680_6031# VGND.t308 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3236 a_5081_4943# net54 a_4863_4917# VGND.t644 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3237 net19 a_8767_11471# VGND.t2927 VGND.t2926 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3238 a_5055_9295# a_4609_9295# a_4959_9295# VGND.t260 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3239 a_14540_3689# a_13625_3317# a_14193_3285# VGND.t2276 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3240 VGND.t889 VPWR.t3574 VGND.t888 VGND.t887 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3241 a_6519_4631# _052_ VPWR.t1116 VPWR.t1115 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X3242 a_13356_7369# _133_ VPWR.t3171 VPWR.t3170 sky130_fd_pr__pfet_01v8_hvt ad=0.117 pd=1.24 as=0.373 ps=1.75 w=1 l=0.15
X3243 VPWR.t1646 a_14715_3615# a_14702_3311# VPWR.t1645 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3244 _087_ a_5455_4943# VGND.t1945 VGND.t1944 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X3245 _004_ _074_ VGND.t138 VGND.t137 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3246 clknet_0_clk a_8022_7119# VPWR.t1576 VPWR.t1575 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3247 VPWR.t720 VGND.t3500 VPWR.t719 VPWR.t718 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3248 a_11599_6397# net46 VPWR.t957 VPWR.t956 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3249 VPWR.t722 VGND.t3501 VPWR.t721 VPWR.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3250 a_7164_11293# _021_ VPWR.t2080 VPWR.t2079 sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X3251 a_2564_2589# _014_ VGND.t3241 VGND.t3240 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3252 VGND.t136 _074_ _010_ VGND.t135 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3253 VGND.t624 net43.t44 a_3565_7119# VGND.t623 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3254 a_2953_9845# a_2787_9845# VGND.t268 VGND.t267 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3255 _135_ a_13111_6031# a_13349_6031# VGND.t786 sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.0878 ps=0.92 w=0.65 l=0.15
X3256 VPWR.t1644 a_10747_8970# _035_ VPWR.t1643 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3257 VPWR.t1479 a_5535_8181# _078_ VPWR.t1478 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3258 VGND.t810 a_10055_2767# net46 VGND.t809 sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3259 VGND.t886 VPWR.t3575 VGND.t885 VGND.t884 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3260 a_1476_4777# a_395_4405# a_1129_4373# VPWR.t2223 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X3261 VGND.t2888 a_2815_9447# _018_ VGND.t2887 sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3262 VPWR.t3138 a_12612_8725# a_12522_8751# VPWR.t3137 sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X3263 a_7351_8041# a_7001_7669# a_7256_8029# VPWR.t1451 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3264 VGND.t883 VPWR.t3576 VGND.t882 VGND.t881 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3265 a_9572_2601# a_8657_2229# a_9225_2197# VGND.t746 sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3266 VPWR.t1267 a_1644_12533# result[7].t0 VPWR.t1266 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3267 VPWR.t2019 a_1497_8725# a_1387_8751# VPWR.t2018 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3268 a_3529_6281# mask\[0\] VPWR.t3049 VPWR.t3048 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3269 a_4687_12319# net43.t45 VPWR.t1378 VPWR.t1377 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3270 net30.t2 a_7939_3855# VGND.t3127 VGND.t3126 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0683 ps=0.745 w=0.42 l=0.15
X3271 a_448_7637# net23 VGND.t1630 VGND.t1629 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3272 net52 a_5691_7637# VGND.t2587 VGND.t2586 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3273 a_4308_4917# net54 VGND.t643 VGND.t642 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3274 VPWR.t1762 clknet_2_0__leaf_clk a_4443_1679# VPWR.t1761 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3275 VGND.t1792 a_1549_6794# net14 VGND.t1791 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3276 VPWR.t2817 a_5177_1921# a_5067_2045# VPWR.t2816 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3277 VGND.t2402 a_8298_2767# clknet_2_2__leaf_clk VGND.t2401 sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3278 VPWR.t2355 a_10543_2455# _027_ VPWR.t2354 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X3279 _098_ _048_.t36 VGND.t2262 VGND.t2261 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3280 clknet_2_0__leaf_clk a_2857_5461# VGND.t654 VGND.t653 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3281 VPWR.t2092 clknet_2_1__leaf_clk.t56 a_7939_10383# VPWR.t2091 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3282 VPWR.t724 VGND.t3502 VPWR.t723 VPWR.t222 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3283 a_2857_7637# clknet_0_clk VPWR.t1050 VPWR.t1049 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3284 a_14099_3017# net49 VPWR.t2705 VPWR.t2704 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3285 VGND.t880 VPWR.t3577 VGND.t879 VGND.t878 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3286 _009_ _074_ VGND.t134 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3287 VPWR.t3238 a_448_7637# result[1].t0 VPWR.t3237 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3288 a_1651_10143# a_1476_10217# a_1830_10205# VGND.t2531 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3289 trimb[4].t4 a_15023_8751# VGND.t2664 VGND.t2663 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3290 VPWR.t1650 net23 a_2174_8457# VPWR.t1649 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X3291 VPWR.t3177 en.t0 a_395_2767# VPWR.t3176 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3292 trimb[3].t0 a_15023_12559# VPWR.t2374 VPWR.t2373 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3293 a_14649_6031# a_14379_6397# a_14564_6397# VGND.t2745 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3294 _076_ _049_ a_6197_6281# VPWR.t1190 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3295 clknet_2_2__leaf_clk a_8298_2767# VPWR.t2435 VPWR.t2434 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3296 VGND.t877 VPWR.t3578 VGND.t876 VGND.t875 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3297 a_9195_10357# a_9020_10383# a_9374_10383# VGND.t2935 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3298 VGND.t182 _067_ a_10043_7983# VGND.t181 sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0959 ps=0.945 w=0.65 l=0.15
X3299 a_14981_4020# _047_ VGND.t1863 VGND.t1862 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3300 a_9503_4399# _107_ _108_ VPWR.t1679 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3301 a_12430_7663# a_11895_7669# a_12344_8041# VPWR.t1936 sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X3302 a_929_8757# a_763_8757# VPWR.t821 VPWR.t820 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3303 VGND.t874 VPWR.t3579 VGND.t873 VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3304 VGND.t2912 rstn.t1 a_395_591# VGND.t2911 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3305 VPWR.t726 VGND.t3503 VPWR.t725 VPWR.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3306 VGND.t3243 a_15023_9839# trimb[1].t4 VGND.t3242 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3307 a_6519_3829# _048_.t37 VPWR.t2288 VPWR.t1115 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.327 ps=1.65 w=1 l=0.15
X3308 a_15259_7637# comp.t1 VGND.t2094 VGND.t2093 sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0683 ps=0.745 w=0.42 l=0.15
X3309 VGND.t871 VPWR.t3580 VGND.t870 VGND.t869 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3310 result[1].t2 a_448_7637# VGND.t3162 VGND.t3161 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.172 ps=1.83 w=0.65 l=0.15
X3311 VPWR.t919 _067_ _072_ VPWR.t918 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3312 a_5055_1679# a_4609_1679# a_4959_1679# VGND.t2868 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3313 VPWR.t3059 net4.t7 a_3339_2767# VPWR.t3058 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X3314 mask\[1\] a_4871_8181# VGND.t1713 VGND.t1712 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3315 a_8949_6031# cal_itt\[2\] VGND.t2983 VGND.t2982 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X3316 a_4055_12015# net43.t46 VPWR.t3116 VPWR.t3115 sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X3317 _091_ a_9443_6059# VPWR.t1523 VPWR.t1522 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X3318 VGND.t2067 clknet_2_1__leaf_clk.t57 a_4443_9295# VGND.t2066 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3319 a_1019_9839# a_395_9845# a_911_10217# VPWR.t2112 sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X3320 VPWR.t2178 _063_.t19 a_9443_6059# VPWR.t2177 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3321 VPWR.t2655 a_15259_7637# net2 VPWR.t2654 sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3322 trim_val\[4\] a_9839_3615# VGND.t2978 VGND.t2977 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.209 ps=2.02 w=0.65 l=0.15
X3323 mask\[3\] a_5699_9269# VPWR.t1176 VPWR.t1175 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3324 VGND.t543 a_14347_4917# a_14281_4943# VGND.t542 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X3325 VGND.t868 VPWR.t3581 VGND.t867 VGND.t866 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3326 a_4959_9295# a_4609_9295# a_4864_9295# VPWR.t998 sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3327 a_11045_3631# trim_mask\[1\] a_10699_3311# VGND.t127 sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3328 a_3365_4943# en_co_clk a_3273_4943# VGND.t2615 sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.201 ps=1.92 w=0.65 l=0.15
X3329 VPWR.t729 VGND.t3504 VPWR.t728 VPWR.t727 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3330 VGND.t3054 state\[1\] a_5087_3855# VGND.t3053 sky130_fd_pr__nfet_01v8 ad=0.0683 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X3331 result[6].t4 a_455_12533# VGND.t2440 VGND.t2439 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3332 _106_ a_8307_4943# VPWR.t1237 VPWR.t1236 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.157 ps=1.32 w=1 l=0.15
X3333 a_7569_7637# a_7351_8041# VGND.t513 VGND.t512 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3334 VGND.t865 VPWR.t3582 VGND.t864 VGND.t863 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3335 a_448_11445# net27 VPWR.t1883 VPWR.t1882 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.149 ps=1.33 w=0.64 l=0.15
X3336 VPWR.t1822 a_12077_3285# a_11967_3311# VPWR.t1821 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3337 a_11508_9295# a_11394_9509# a_11436_9295# VGND.t3068 sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X3338 VPWR.t2300 a_14193_3285# a_14083_3311# VPWR.t2299 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3339 a_12502_4765# net46 VGND.t221 VGND.t220 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X3340 _119_ a_9003_3829# VPWR.t1158 VPWR.t1157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3341 clknet_2_3__leaf_clk a_8298_5487# VGND.t2100 VGND.t2099 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3342 a_8386_8457# _070_ a_8083_8181# VPWR.t2000 sky130_fd_pr__pfet_01v8_hvt ad=0.153 pd=1.3 as=0.195 ps=1.39 w=1 l=0.15
X3343 a_11545_9049# cal_count\[0\] VPWR.t2988 VPWR.t2987 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3344 a_10903_7261# clknet_2_3__leaf_clk VPWR.t1909 VPWR.t1908 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3345 _051_.t0 a_3933_2767# VPWR.t1241 VPWR.t1240 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3346 a_7986_10927# a_6909_10933# a_7824_11305# VPWR.t2672 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3347 VGND.t2537 a_5691_2741# _050_ VGND.t2536 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3348 VPWR.t1154 a_11801_4373# a_11691_4399# VPWR.t1153 sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X3349 VPWR.t731 VGND.t3505 VPWR.t730 VPWR.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3350 a_3830_6281# _120_ a_3748_6281# VPWR.t2948 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X3351 VGND.t451 _049_ a_4498_4373# VGND.t450 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3352 VGND.t862 VPWR.t3583 VGND.t861 VGND.t860 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3353 a_7723_6807# _072_ VPWR.t2799 VPWR.t2798 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X3354 a_6941_2589# a_6906_2355# a_6703_2197# VGND.t1984 sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.109 ps=1.36 w=0.42 l=0.15
X3355 a_911_4777# a_395_4405# a_816_4765# VGND.t2197 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3356 VPWR.t2292 net21 a_5363_12559# VPWR.t2291 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3357 a_6796_12381# _009_ VGND.t2218 VGND.t2217 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X3358 a_7933_11305# a_6743_10933# a_7824_11305# VGND.t2532 sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3359 _020_ a_6099_10633# VGND.t1962 VGND.t1961 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.96 w=0.65 l=0.15
X3360 VGND.t3103 net5 a_15299_6575# VGND.t3102 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3361 VPWR.t734 VGND.t3506 VPWR.t733 VPWR.t732 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3362 VGND.t379 _052_ a_7320_3631# VGND.t378 sky130_fd_pr__nfet_01v8 ad=0.167 pd=1.16 as=0.0975 ps=0.95 w=0.65 l=0.15
X3363 VGND.t859 VPWR.t3584 VGND.t858 VGND.t857 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3364 a_1191_11305# a_745_10933# a_1095_11305# VGND.t1701 sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3365 a_1835_11231# net43.t47 VPWR.t3118 VPWR.t3117 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3366 _117_ a_9719_1473# VPWR.t1180 VPWR.t1179 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X3367 a_7393_5193# _092_ VPWR.t2861 VPWR.t2860 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3368 VGND.t856 VPWR.t3585 VGND.t855 VGND.t854 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3369 trimb[1].t0 a_15023_9839# VPWR.t3322 VPWR.t3321 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3370 VPWR.t3035 a_9839_3615# a_9826_3311# VPWR.t3034 sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3371 net12 net20.t7 VGND.t2196 VGND.t2195 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3372 a_3123_3615# a_2948_3689# a_3302_3677# VGND.t1768 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X3373 a_8307_4719# net30.t11 _104_ VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X3374 VPWR.t737 VGND.t3507 VPWR.t736 VPWR.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X3375 VPWR.t2872 a_2283_4020# _013_ VPWR.t2871 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3376 a_9805_1473# _110_.t9 a_9719_1473# VGND.t2141 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X3377 a_448_11445# net27 VGND.t1857 VGND.t1856 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3378 VPWR.t1011 clknet_2_2__leaf_clk a_8491_2229# VPWR.t1010 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X3379 a_1679_10633# _102_ VPWR.t850 VPWR.t849 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3380 net34.t1 a_14931_591# VGND.t3109 VGND.t3108 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3381 net40 net35 VPWR.t1316 VPWR.t1315 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3382 a_4993_6273# a_4775_6031# VGND.t2741 VGND.t2740 sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X3383 a_2225_7663# mask\[1\] VPWR.t1796 VPWR.t1795 sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.253 ps=2.52 w=1 l=0.15
X3384 VGND.t853 VPWR.t3586 VGND.t852 VGND.t851 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3385 ctlp[0].t0 a_1099_12533# VPWR.t1471 VPWR.t1470 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3386 a_8717_10383# a_8673_10625# a_8551_10383# VGND.t2934 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3387 en_co_clk a_5515_6005# VPWR.t3076 VPWR.t3075 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3388 VGND.t3107 en.t1 a_395_2767# VGND.t3106 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X3389 a_1679_10633# _074_ a_1461_10357# VPWR.t873 sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3390 VPWR.t739 VGND.t3508 VPWR.t738 VPWR.t503 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3391 VPWR.t2732 a_15023_1135# trim[3].t0 VPWR.t2731 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3392 a_2877_2197# a_2659_2601# VPWR.t1450 VPWR.t1449 sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
X3393 a_13625_3317# a_13459_3317# VGND.t178 VGND.t177 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3394 a_11509_3317# a_11343_3317# VGND.t2235 VGND.t2234 sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3395 _108_ _107_ VGND.t1659 VGND.t1658 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3396 VGND.t219 net46 a_9361_3677# VGND.t218 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3397 a_6197_4399# _087_ VPWR.t852 VPWR.t851 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3398 a_3781_8207# a_3615_8207# VPWR.t1684 VPWR.t1683 sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3399 VGND.t1746 clknet_2_0__leaf_clk a_4443_1679# VGND.t1745 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X3400 clknet_2_0__leaf_clk a_2857_5461# VPWR.t1408 VPWR.t1407 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3401 VPWR.t2557 a_455_5747# sample.t0 VPWR.t2556 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3402 state\[2\] a_5699_1653# VPWR.t2695 VPWR.t2694 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.301 ps=2.66 w=1 l=0.15
X3403 _048_.t0 a_3667_3829# VPWR.t3289 VPWR.t3288 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3404 VGND.t1835 a_9802_4007# a_9662_3855# VGND.t1834 sky130_fd_pr__nfet_01v8 ad=0.109 pd=0.985 as=0.26 ps=1.45 w=0.65 l=0.15
X3405 VGND.t850 VPWR.t3587 VGND.t849 VGND.t848 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
R0 VPWR.t142 VPWR 1719.47
R1 VPWR.t119 VPWR 1719.47
R2 VPWR VPWR.t454 1719.47
R3 VPWR.t668 VPWR 1716.51
R4 VPWR VPWR.t142 1547.82
R5 VPWR VPWR.t119 1547.82
R6 VPWR VPWR.t668 1547.82
R7 VPWR.t454 VPWR 1547.82
R8 VPWR.n4536 VPWR.n4485 1409.47
R9 VPWR.n7279 VPWR.t469 1225.23
R10 VPWR.t577 VPWR 1180.84
R11 VPWR VPWR.t577 1003.27
R12 VPWR.t469 VPWR 1003.27
R13 VPWR VPWR.t213 975.178
R14 VPWR.t213 VPWR 877.827
R15 VPWR VPWR.t480 820.76
R16 VPWR VPWR.t2303 742.836
R17 VPWR.t406 VPWR 723.41
R18 VPWR.t2379 VPWR.t718 713.24
R19 VPWR.t2476 VPWR.t175 713.24
R20 VPWR.t842 VPWR.t12 689.564
R21 VPWR.n7281 VPWR.t430 680.686
R22 VPWR.t89 VPWR 669.701
R23 VPWR VPWR.t554 666.343
R24 VPWR VPWR.t190 666.343
R25 VPWR VPWR.t545 664.664
R26 VPWR.t433 VPWR 636.293
R27 VPWR VPWR.t512 636.293
R28 VPWR VPWR.t27 636.293
R29 VPWR.t98 VPWR.t148 617.668
R30 VPWR.t306 VPWR.t660 617.668
R31 VPWR.t528 VPWR.t542 617.668
R32 VPWR.t210 VPWR.t712 617.668
R33 VPWR.t57 VPWR.t445 617.668
R34 VPWR.t703 VPWR.t486 617.668
R35 VPWR.t107 VPWR.t674 617.668
R36 VPWR.t495 VPWR.t318 617.668
R37 VPWR VPWR.n6955 597.819
R38 VPWR.n1783 VPWR.t1611 580.938
R39 VPWR.n5282 VPWR.t2611 580.938
R40 VPWR.n4671 VPWR.t2924 579.029
R41 VPWR.n1785 VPWR.t1613 578.254
R42 VPWR VPWR.t489 568.994
R43 VPWR.t727 VPWR 568.994
R44 VPWR.t625 VPWR 568.994
R45 VPWR VPWR.t75 568.994
R46 VPWR VPWR.t225 568.994
R47 VPWR VPWR.t571 568.994
R48 VPWR VPWR.t261 568.994
R49 VPWR.t568 VPWR 568.994
R50 VPWR.n6627 VPWR.t3148 549.573
R51 VPWR.n541 VPWR.t2600 546.317
R52 VPWR.n5123 VPWR.t3200 543.624
R53 VPWR.n621 VPWR.t2591 541.831
R54 VPWR.n8425 VPWR.t1547 541.275
R55 VPWR.n5863 VPWR.t397 540.46
R56 VPWR.n615 VPWR.t2657 540.376
R57 VPWR.n1890 VPWR.t3330 540.376
R58 VPWR.n1372 VPWR.t2409 538.203
R59 VPWR.n1320 VPWR.t2725 538.203
R60 VPWR.n1309 VPWR.t111 521.032
R61 VPWR.n3886 VPWR.t182 519.641
R62 VPWR.n6288 VPWR.t286 519.641
R63 VPWR.n486 VPWR.t710 519.641
R64 VPWR.n452 VPWR.t395 519.641
R65 VPWR.n4074 VPWR.t481 519.418
R66 VPWR.n5490 VPWR.t369 519.418
R67 VPWR.n4771 VPWR.t22 519.418
R68 VPWR VPWR.t436 515.284
R69 VPWR VPWR.t45 515.284
R70 VPWR.n3635 VPWR.t644 515.067
R71 VPWR.n3027 VPWR.t183 515.048
R72 VPWR.n7757 VPWR.t308 515.048
R73 VPWR.n6264 VPWR.t287 515.048
R74 VPWR.n6644 VPWR.t109 515.048
R75 VPWR.n4029 VPWR.t555 514.981
R76 VPWR.n3638 VPWR.t26 514.981
R77 VPWR.n9179 VPWR.t1206 514.263
R78 VPWR.n1163 VPWR.t1509 514.011
R79 VPWR.n2214 VPWR.t997 514.011
R80 VPWR.n6228 VPWR.t59 513.976
R81 VPWR.n4407 VPWR.t118 513.976
R82 VPWR.n5969 VPWR.t488 513.923
R83 VPWR.n7637 VPWR.t426 513.457
R84 VPWR.n6255 VPWR.t704 513.004
R85 VPWR.n6952 VPWR.t120 512.231
R86 VPWR.n7473 VPWR.t121 512.231
R87 VPWR.n7570 VPWR.t143 512.231
R88 VPWR.n6941 VPWR.t144 512.231
R89 VPWR.n6956 VPWR.t669 512.231
R90 VPWR.n7030 VPWR.t670 512.231
R91 VPWR.n3870 VPWR.t666 512.231
R92 VPWR.n3049 VPWR.t667 512.231
R93 VPWR.n3287 VPWR.t170 512.231
R94 VPWR.n3144 VPWR.t171 512.231
R95 VPWR.n3208 VPWR.t99 512.231
R96 VPWR.n3152 VPWR.t100 512.231
R97 VPWR.n3151 VPWR.t149 512.231
R98 VPWR.n3153 VPWR.t150 512.231
R99 VPWR.n3912 VPWR.t428 512.231
R100 VPWR.n4001 VPWR.t429 512.231
R101 VPWR.n4054 VPWR.t627 512.231
R102 VPWR.n2996 VPWR.t556 512.231
R103 VPWR.n4032 VPWR.t626 512.231
R104 VPWR.n4086 VPWR.t482 512.231
R105 VPWR.n4075 VPWR.t407 512.231
R106 VPWR.n4127 VPWR.t408 512.231
R107 VPWR.n6013 VPWR.t305 512.231
R108 VPWR.n6018 VPWR.t32 512.231
R109 VPWR.n6029 VPWR.t304 512.231
R110 VPWR.n7821 VPWR.t31 512.231
R111 VPWR.n6019 VPWR.t633 512.231
R112 VPWR.n6009 VPWR.t714 512.231
R113 VPWR.n7810 VPWR.t632 512.231
R114 VPWR.n7792 VPWR.t713 512.231
R115 VPWR.n6113 VPWR.t212 512.231
R116 VPWR.n6116 VPWR.t544 512.231
R117 VPWR.n7783 VPWR.t211 512.231
R118 VPWR.n6121 VPWR.t543 512.231
R119 VPWR.n6118 VPWR.t530 512.231
R120 VPWR.n6119 VPWR.t529 512.231
R121 VPWR.n7751 VPWR.t662 512.231
R122 VPWR.n6129 VPWR.t307 512.231
R123 VPWR.n7679 VPWR.t661 512.231
R124 VPWR.n7655 VPWR.t425 512.231
R125 VPWR.n6226 VPWR.t447 512.231
R126 VPWR.n6870 VPWR.t58 512.231
R127 VPWR.n6258 VPWR.t487 512.231
R128 VPWR.n5967 VPWR.t705 512.231
R129 VPWR.n7903 VPWR.t5 512.231
R130 VPWR.n7902 VPWR.t4 512.231
R131 VPWR.n8979 VPWR.t363 512.231
R132 VPWR.n8065 VPWR.t362 512.231
R133 VPWR.n8016 VPWR.t167 512.231
R134 VPWR.n5964 VPWR.t168 512.231
R135 VPWR.n8986 VPWR.t681 512.231
R136 VPWR.n9015 VPWR.t682 512.231
R137 VPWR.n9019 VPWR.t345 512.231
R138 VPWR.n8975 VPWR.t346 512.231
R139 VPWR.n6192 VPWR.t446 512.231
R140 VPWR.n6641 VPWR.t676 512.231
R141 VPWR.n6792 VPWR.t108 512.231
R142 VPWR.n6759 VPWR.t374 512.231
R143 VPWR.n6648 VPWR.t375 512.231
R144 VPWR.n6651 VPWR.t441 512.231
R145 VPWR.n6649 VPWR.t440 512.231
R146 VPWR.n5946 VPWR.t10 512.231
R147 VPWR.n5949 VPWR.t11 512.231
R148 VPWR.n6635 VPWR.t675 512.231
R149 VPWR.n6810 VPWR.t602 512.231
R150 VPWR.n6617 VPWR.t601 512.231
R151 VPWR.n8485 VPWR.t399 512.231
R152 VPWR.n8461 VPWR.t398 512.231
R153 VPWR.n6353 VPWR.t392 512.231
R154 VPWR.n8373 VPWR.t393 512.231
R155 VPWR.n6379 VPWR.t134 512.231
R156 VPWR.n6356 VPWR.t135 512.231
R157 VPWR.n1370 VPWR.t112 512.231
R158 VPWR.n1514 VPWR.t377 512.231
R159 VPWR.n1376 VPWR.t378 512.231
R160 VPWR.n1378 VPWR.t444 512.231
R161 VPWR.n1377 VPWR.t443 512.231
R162 VPWR.n5467 VPWR.t368 512.231
R163 VPWR.n472 VPWR.t711 512.231
R164 VPWR.n5614 VPWR.t322 512.231
R165 VPWR.n455 VPWR.t323 512.231
R166 VPWR.n401 VPWR.t396 512.231
R167 VPWR.n4786 VPWR.t23 512.231
R168 VPWR.n4787 VPWR.t386 512.231
R169 VPWR.n4793 VPWR.t387 512.231
R170 VPWR.n558 VPWR.t236 512.231
R171 VPWR.n1639 VPWR.t235 512.231
R172 VPWR.n1670 VPWR.t496 512.231
R173 VPWR.n1686 VPWR.t319 512.231
R174 VPWR.n557 VPWR.t497 512.231
R175 VPWR.n1710 VPWR.t320 512.231
R176 VPWR.n1794 VPWR.t245 512.231
R177 VPWR.n1787 VPWR.t244 512.231
R178 VPWR.n2182 VPWR.t93 512.231
R179 VPWR.n2121 VPWR.t94 512.231
R180 VPWR.n2727 VPWR.t117 512.231
R181 VPWR.n2020 VPWR.t357 512.231
R182 VPWR.n2700 VPWR.t356 512.231
R183 VPWR.n2305 VPWR.t292 512.231
R184 VPWR.n2306 VPWR.t293 512.231
R185 VPWR.n4532 VPWR.t102 512.231
R186 VPWR.n4490 VPWR.t103 512.231
R187 VPWR.n4242 VPWR.t340 512.231
R188 VPWR.n2886 VPWR.t341 512.231
R189 VPWR.n2888 VPWR.t683 512.231
R190 VPWR.n2889 VPWR.t684 512.231
R191 VPWR.n2889 VPWR.t215 512.231
R192 VPWR.n2888 VPWR.t214 512.231
R193 VPWR.n2834 VPWR.t152 512.231
R194 VPWR.n2793 VPWR.t153 512.231
R195 VPWR.n2788 VPWR.t645 512.231
R196 VPWR.n3632 VPWR.t25 512.231
R197 VPWR.n3595 VPWR.t549 512.231
R198 VPWR.n3522 VPWR.t550 512.231
R199 VPWR.n3506 VPWR.t126 512.231
R200 VPWR.n3509 VPWR.t127 512.231
R201 VPWR.n2800 VPWR.t247 512.231
R202 VPWR.n2828 VPWR.t248 512.231
R203 VPWR.n7081 VPWR.t455 512.231
R204 VPWR.n7049 VPWR.t456 512.231
R205 VPWR VPWR.t631 511.926
R206 VPWR VPWR.t574 511.926
R207 VPWR VPWR.t163 511.926
R208 VPWR VPWR.t69 511.926
R209 VPWR.n3286 VPWR.t1142 511.072
R210 VPWR.n101 VPWR.t2669 511.072
R211 VPWR.n6095 VPWR.t2728 511.072
R212 VPWR.n8015 VPWR.t2314 511.072
R213 VPWR.n250 VPWR.t2878 511.072
R214 VPWR.n9000 VPWR.t1724 511.072
R215 VPWR.n7932 VPWR.t775 511.072
R216 VPWR.n8864 VPWR.t2815 511.072
R217 VPWR.n8159 VPWR.t2960 511.072
R218 VPWR.n8327 VPWR.t1820 511.072
R219 VPWR.n5942 VPWR.t2394 511.072
R220 VPWR.n8192 VPWR.t825 511.072
R221 VPWR.n8783 VPWR.t1758 511.072
R222 VPWR.n8666 VPWR.t3277 511.072
R223 VPWR.n5817 VPWR.t2357 511.072
R224 VPWR.n1014 VPWR.t2370 511.072
R225 VPWR.n992 VPWR.t1253 511.072
R226 VPWR.n811 VPWR.t763 511.072
R227 VPWR.n437 VPWR.t1617 511.072
R228 VPWR.n5592 VPWR.t2782 511.072
R229 VPWR.n1472 VPWR.t2671 511.072
R230 VPWR.n1581 VPWR.t2285 511.072
R231 VPWR.n4913 VPWR.t2950 511.072
R232 VPWR.n2165 VPWR.t2928 511.072
R233 VPWR.n2354 VPWR.t2082 511.072
R234 VPWR.n2097 VPWR.t2653 511.072
R235 VPWR.n2003 VPWR.t1810 511.072
R236 VPWR.n2853 VPWR.t1450 511.072
R237 VPWR.n3583 VPWR.t2404 511.072
R238 VPWR.n3505 VPWR.t928 511.072
R239 VPWR.n3679 VPWR.t2784 511.072
R240 VPWR.n3630 VPWR.t3175 511.072
R241 VPWR.n4253 VPWR.t2797 511.072
R242 VPWR.n8053 VPWR.t2497 497.185
R243 VPWR.n8057 VPWR.t1351 497.185
R244 VPWR.n8173 VPWR.t2160 497.185
R245 VPWR.n8133 VPWR.t2685 497.185
R246 VPWR.n1716 VPWR.t2641 497.185
R247 VPWR.n1921 VPWR.t3008 497.185
R248 VPWR.n2122 VPWR.t1902 497.185
R249 VPWR.n2326 VPWR.t872 497.185
R250 VPWR.n2312 VPWR.t2887 497.185
R251 VPWR.n3517 VPWR.t2099 497.185
R252 VPWR.t640 VPWR 494.238
R253 VPWR VPWR.t557 494.238
R254 VPWR.n9038 VPWR.t3029 494.12
R255 VPWR.n8637 VPWR.t3187 494.12
R256 VPWR.n384 VPWR.t1796 494.12
R257 VPWR.n4943 VPWR.t1494 494.12
R258 VPWR.n6111 VPWR 491.784
R259 VPWR VPWR.n8012 491.784
R260 VPWR.n722 VPWR.t1086 490.902
R261 VPWR.n1727 VPWR.t2143 490.902
R262 VPWR.n4642 VPWR.t1434 487.971
R263 VPWR.n935 VPWR.t1603 486.873
R264 VPWR.n2662 VPWR.t2441 486.873
R265 VPWR.t1476 VPWR 485.358
R266 VPWR.n593 VPWR.t2998 477.421
R267 VPWR.n1513 VPWR.t1543 474.63
R268 VPWR.n1360 VPWR.t2720 474.123
R269 VPWR.t1268 VPWR 467.601
R270 VPWR.t631 VPWR.t30 463.252
R271 VPWR.t339 VPWR.t620 463.252
R272 VPWR VPWR.t3243 461.683
R273 VPWR.n7989 VPWR.t535 459.474
R274 VPWR.n3062 VPWR.t96 459.192
R275 VPWR.n3065 VPWR.t490 459.192
R276 VPWR.n3033 VPWR.t298 459.192
R277 VPWR.n3910 VPWR.t728 459.192
R278 VPWR.n4008 VPWR.t686 459.192
R279 VPWR.n4115 VPWR.t586 459.192
R280 VPWR.n4114 VPWR.t587 459.192
R281 VPWR.n4093 VPWR.t733 459.192
R282 VPWR.n9201 VPWR.t241 459.192
R283 VPWR.n9133 VPWR.t452 459.192
R284 VPWR.n7762 VPWR.t311 459.192
R285 VPWR.n7759 VPWR.t310 459.192
R286 VPWR.n7636 VPWR.t76 459.192
R287 VPWR.n6290 VPWR.t161 459.192
R288 VPWR.n6236 VPWR.t331 459.192
R289 VPWR.n6235 VPWR.t332 459.192
R290 VPWR.n8966 VPWR.t64 459.192
R291 VPWR.n6156 VPWR.t572 459.192
R292 VPWR.n6159 VPWR.t226 459.192
R293 VPWR.n337 VPWR.t561 459.192
R294 VPWR.n6751 VPWR.t262 459.192
R295 VPWR.n6666 VPWR.t114 459.192
R296 VPWR.n8622 VPWR.t656 459.192
R297 VPWR.n5865 VPWR.t140 459.192
R298 VPWR.n5867 VPWR.t635 459.192
R299 VPWR.n6361 VPWR.t49 459.192
R300 VPWR.n822 VPWR.t595 459.192
R301 VPWR.n813 VPWR.t158 459.192
R302 VPWR.n495 VPWR.t458 459.192
R303 VPWR.n465 VPWR.t464 459.192
R304 VPWR.n404 VPWR.t607 459.192
R305 VPWR.n4639 VPWR.t592 459.192
R306 VPWR.n4636 VPWR.t593 459.192
R307 VPWR.n1539 VPWR.t716 459.192
R308 VPWR.n5003 VPWR.t40 459.192
R309 VPWR.n1902 VPWR.t613 459.192
R310 VPWR.n2296 VPWR.t200 459.192
R311 VPWR.n1995 VPWR.t313 459.192
R312 VPWR VPWR.t433 458.724
R313 VPWR.t430 VPWR 458.724
R314 VPWR.t512 VPWR 458.724
R315 VPWR.t27 VPWR 458.724
R316 VPWR.t1274 VPWR.t2925 448.146
R317 VPWR.t2079 VPWR.t2572 448.146
R318 VPWR.t895 VPWR.t1665 448.146
R319 VPWR.t1752 VPWR.t2470 448.146
R320 VPWR.t2743 VPWR.t2359 448.146
R321 VPWR.t2400 VPWR.t1445 448.146
R322 VPWR.t1131 VPWR.t1976 448.146
R323 VPWR.t3319 VPWR.t2381 448.146
R324 VPWR.t234 VPWR.t747 438.075
R325 VPWR.n2991 VPWR.t105 432.673
R326 VPWR.n3147 VPWR.t590 432.673
R327 VPWR.n3056 VPWR.t254 432.673
R328 VPWR.n3028 VPWR.t129 432.673
R329 VPWR.n4101 VPWR.t701 432.673
R330 VPWR.n4096 VPWR.t275 432.673
R331 VPWR.n3246 VPWR.t342 432.673
R332 VPWR.n3242 VPWR.t156 432.673
R333 VPWR.n77 VPWR.t699 432.673
R334 VPWR.n74 VPWR.t230 432.673
R335 VPWR.n65 VPWR.t422 432.673
R336 VPWR.n7643 VPWR.t501 432.673
R337 VPWR.n7640 VPWR.t17 432.673
R338 VPWR.n7651 VPWR.t1 432.673
R339 VPWR.n6015 VPWR.t334 432.673
R340 VPWR.n6274 VPWR.t348 432.673
R341 VPWR.n6165 VPWR.t552 432.673
R342 VPWR.n6172 VPWR.t301 432.673
R343 VPWR.n6168 VPWR.t521 432.673
R344 VPWR.n220 VPWR.t478 432.673
R345 VPWR.n217 VPWR.t722 432.673
R346 VPWR.n8295 VPWR.t523 432.673
R347 VPWR.n8878 VPWR.t197 432.673
R348 VPWR.n8875 VPWR.t209 432.673
R349 VPWR.n6653 VPWR.t132 432.673
R350 VPWR.n8146 VPWR.t7 432.673
R351 VPWR.n6592 VPWR.t73 432.673
R352 VPWR.n6589 VPWR.t79 432.673
R353 VPWR.n8744 VPWR.t723 432.673
R354 VPWR.n8740 VPWR.t224 432.673
R355 VPWR.n5874 VPWR.t232 432.673
R356 VPWR.n8616 VPWR.t62 432.673
R357 VPWR.n6496 VPWR.t615 432.673
R358 VPWR.n6492 VPWR.t88 432.673
R359 VPWR.n6485 VPWR.t269 432.673
R360 VPWR.n5789 VPWR.t504 432.673
R361 VPWR.n5786 VPWR.t739 432.673
R362 VPWR.n727 VPWR.t186 432.673
R363 VPWR.n801 VPWR.t251 432.673
R364 VPWR.n606 VPWR.t383 432.673
R365 VPWR.n603 VPWR.t624 432.673
R366 VPWR.n596 VPWR.t317 432.673
R367 VPWR.n1443 VPWR.t638 432.673
R368 VPWR.n416 VPWR.t137 432.673
R369 VPWR.n413 VPWR.t538 432.673
R370 VPWR.n1280 VPWR.t730 432.673
R371 VPWR.n1277 VPWR.t417 432.673
R372 VPWR.n1288 VPWR.t271 432.673
R373 VPWR.n4643 VPWR.t516 432.673
R374 VPWR.n4798 VPWR.t658 432.673
R375 VPWR.n4794 VPWR.t326 432.673
R376 VPWR.n1550 VPWR.t518 432.673
R377 VPWR.n1546 VPWR.t204 432.673
R378 VPWR.n530 VPWR.t173 432.673
R379 VPWR.n1905 VPWR.t698 432.673
R380 VPWR.n4926 VPWR.t663 432.673
R381 VPWR.n4922 VPWR.t124 432.673
R382 VPWR.n1835 VPWR.t84 432.673
R383 VPWR.n1841 VPWR.t484 432.673
R384 VPWR.n2117 VPWR.t581 432.673
R385 VPWR.n2437 VPWR.t540 432.673
R386 VPWR.n2434 VPWR.t726 432.673
R387 VPWR.n2219 VPWR.t328 432.673
R388 VPWR.n2215 VPWR.t567 432.673
R389 VPWR.n2013 VPWR.t629 432.673
R390 VPWR.n2028 VPWR.t52 432.673
R391 VPWR.n2024 VPWR.t280 432.673
R392 VPWR.n2010 VPWR.t527 432.673
R393 VPWR.n4500 VPWR.t449 432.673
R394 VPWR.n4497 VPWR.t692 432.673
R395 VPWR.n2894 VPWR.t217 432.673
R396 VPWR.n2890 VPWR.t473 432.673
R397 VPWR.n3375 VPWR.t81 432.673
R398 VPWR.n3372 VPWR.t351 432.673
R399 VPWR.n3383 VPWR.t353 432.673
R400 VPWR.n3510 VPWR.t468 432.673
R401 VPWR.n6371 VPWR.t2730 426.039
R402 VPWR.n943 VPWR.n942 425.026
R403 VPWR.n1846 VPWR.n1845 424.32
R404 VPWR VPWR.t2662 422.969
R405 VPWR.t1643 VPWR 419.611
R406 VPWR.t1292 VPWR 419.611
R407 VPWR.t2057 VPWR.n6943 417.291
R408 VPWR.n6650 VPWR.t1521 416.543
R409 VPWR.n834 VPWR.t835 416.543
R410 VPWR.t309 VPWR 414.577
R411 VPWR.t30 VPWR 414.577
R412 VPWR.t330 VPWR 414.577
R413 VPWR.t21 VPWR 414.577
R414 VPWR.t163 VPWR 414.577
R415 VPWR.t620 VPWR 414.577
R416 VPWR VPWR.t885 411.372
R417 VPWR.t2735 VPWR.t154 404.505
R418 VPWR.t2185 VPWR.t15 404.505
R419 VPWR.t2044 VPWR.t300 404.505
R420 VPWR.t2713 VPWR.t86 404.505
R421 VPWR.t1230 VPWR.t202 404.505
R422 VPWR.t3211 VPWR.t80 404.505
R423 VPWR.n4424 VPWR.t3126 395.644
R424 VPWR.t252 VPWR.t3203 392.757
R425 VPWR.t3221 VPWR 391.079
R426 VPWR VPWR.t2270 390.654
R427 VPWR VPWR.t2071 390.654
R428 VPWR.t1179 VPWR.t786 389.399
R429 VPWR.t2187 VPWR 389.399
R430 VPWR.t315 VPWR.t2656 389.399
R431 VPWR.t1659 VPWR.t415 389.399
R432 VPWR.t2468 VPWR 389.399
R433 VPWR.t2309 VPWR.t327 389.399
R434 VPWR.t2582 VPWR.t628 389.399
R435 VPWR.n3880 VPWR.t297 386.043
R436 VPWR.n6227 VPWR.t160 386.043
R437 VPWR.n500 VPWR.t2607 382.793
R438 VPWR.n3737 VPWR.t2168 382.793
R439 VPWR.n3043 VPWR.t2164 378.908
R440 VPWR.n6516 VPWR.t2419 378.908
R441 VPWR.n5442 VPWR.t2956 378.908
R442 VPWR.n2554 VPWR.t3136 378.908
R443 VPWR.n2530 VPWR.t2170 378.908
R444 VPWR.n8985 VPWR.t1448 376.663
R445 VPWR.n1488 VPWR.t1271 376.663
R446 VPWR.n8920 VPWR.t2569 376.26
R447 VPWR.n3514 VPWR.t2813 376.202
R448 VPWR.n5119 VPWR.t2762 376.103
R449 VPWR.n975 VPWR.t1794 375.445
R450 VPWR.n8871 VPWR.t2894 375.277
R451 VPWR.n8171 VPWR.t1607 375.277
R452 VPWR.n8135 VPWR.t2922 375.277
R453 VPWR.n5781 VPWR.t2975 375.277
R454 VPWR.n1010 VPWR.t1727 375.277
R455 VPWR.n1457 VPWR.t1658 375.277
R456 VPWR.n4936 VPWR.t2433 375.277
R457 VPWR.n2288 VPWR.t1625 375.277
R458 VPWR.n3554 VPWR.t3224 375.277
R459 VPWR.n8242 VPWR.t1501 375.252
R460 VPWR.n5832 VPWR.t1005 375.252
R461 VPWR.n1000 VPWR.t3285 375.252
R462 VPWR.n1577 VPWR.t1519 375.252
R463 VPWR.n2240 VPWR.t2882 375.252
R464 VPWR.n2367 VPWR.t2257 375.252
R465 VPWR.n3546 VPWR.t2952 375.252
R466 VPWR.n816 VPWR.t2255 373.76
R467 VPWR.n426 VPWR.t1629 373.236
R468 VPWR.n2336 VPWR.t1929 373.072
R469 VPWR.n5251 VPWR.t3192 372.974
R470 VPWR.n8125 VPWR.t2298 372.079
R471 VPWR.n805 VPWR.t1312 372.079
R472 VPWR.n8674 VPWR.t1662 372.079
R473 VPWR.n3268 VPWR.t3144 371.954
R474 VPWR.n34 VPWR.t3019 371.954
R475 VPWR.n6010 VPWR.t2316 371.954
R476 VPWR.n263 VPWR.t1965 371.954
R477 VPWR.n7915 VPWR.t1995 371.954
R478 VPWR.n7948 VPWR.t2983 371.954
R479 VPWR.n8298 VPWR.t1722 371.954
R480 VPWR.n8686 VPWR.t2290 371.954
R481 VPWR.n1142 VPWR.t3262 371.954
R482 VPWR.n448 VPWR.t2811 371.954
R483 VPWR.n5578 VPWR.t2912 371.954
R484 VPWR.n1964 VPWR.t1218 371.954
R485 VPWR.n2181 VPWR.t2367 371.954
R486 VPWR.n2683 VPWR.t2786 371.954
R487 VPWR.n2006 VPWR.t1786 371.954
R488 VPWR.n2837 VPWR.t2971 371.954
R489 VPWR.n3729 VPWR.t2827 371.954
R490 VPWR.n3647 VPWR.t2012 371.954
R491 VPWR.n4277 VPWR.t1388 371.954
R492 VPWR.n68 VPWR.t936 371.825
R493 VPWR.n1998 VPWR.t2467 371.57
R494 VPWR.n3226 VPWR.t2926 370.925
R495 VPWR.n47 VPWR.t2870 370.925
R496 VPWR.n6082 VPWR.t2243 370.925
R497 VPWR.n8034 VPWR.t2080 370.925
R498 VPWR.n235 VPWR.t2188 370.925
R499 VPWR.n9018 VPWR.t896 370.925
R500 VPWR.n7916 VPWR.t1993 370.925
R501 VPWR.n5925 VPWR.t1615 370.925
R502 VPWR.n8269 VPWR.t908 370.925
R503 VPWR.n8767 VPWR.t3222 370.925
R504 VPWR.n8649 VPWR.t2691 370.925
R505 VPWR.n1184 VPWR.t2363 370.925
R506 VPWR.n1033 VPWR.t2084 370.925
R507 VPWR.n5598 VPWR.t2469 370.925
R508 VPWR.n1647 VPWR.t748 370.925
R509 VPWR.n2148 VPWR.t2107 370.925
R510 VPWR.n2074 VPWR.t1877 370.925
R511 VPWR.n4241 VPWR.t3320 370.925
R512 VPWR.n3598 VPWR.t2744 370.925
R513 VPWR.n3620 VPWR.t1446 370.925
R514 VPWR.n3700 VPWR.t2471 370.925
R515 VPWR.n2805 VPWR.t1132 370.925
R516 VPWR.n4685 VPWR.t1676 370.341
R517 VPWR.n9136 VPWR.t1631 368.192
R518 VPWR.n6669 VPWR.t1525 368.192
R519 VPWR.n6453 VPWR.t1857 367.724
R520 VPWR.t914 VPWR 367.579
R521 VPWR.n6721 VPWR.t3134 364.812
R522 VPWR.t1488 VPWR 364.019
R523 VPWR VPWR.t832 364.019
R524 VPWR.n497 VPWR.t2954 363.233
R525 VPWR VPWR.t585 360.866
R526 VPWR.t2982 VPWR.t2806 360.866
R527 VPWR.t2108 VPWR.t1964 360.866
R528 VPWR.t2891 VPWR.t2810 360.866
R529 VPWR.t1518 VPWR.t1284 360.866
R530 VPWR.t2978 VPWR.t1217 360.866
R531 VPWR VPWR.t403 360.866
R532 VPWR VPWR.t609 360.866
R533 VPWR.t2694 VPWR.t1387 360.866
R534 VPWR.t1254 VPWR.t2970 360.866
R535 VPWR.n626 VPWR.t3085 360.43
R536 VPWR.t1654 VPWR.t2093 359.188
R537 VPWR.t2413 VPWR.t3312 359.188
R538 VPWR VPWR.t727 357.51
R539 VPWR.t660 VPWR 357.51
R540 VPWR VPWR.t528 357.51
R541 VPWR VPWR.t210 357.51
R542 VPWR.t445 VPWR 357.51
R543 VPWR VPWR.t703 357.51
R544 VPWR.t674 VPWR 357.51
R545 VPWR.t261 VPWR 357.51
R546 VPWR VPWR.t693 357.51
R547 VPWR VPWR.t42 357.51
R548 VPWR VPWR.t495 357.51
R549 VPWR.t358 VPWR 357.51
R550 VPWR VPWR.t98 355.83
R551 VPWR VPWR.t685 355.83
R552 VPWR.n1208 VPWR.t3230 355.822
R553 VPWR.t1383 VPWR.t3075 342.404
R554 VPWR.t2171 VPWR.t768 342.404
R555 VPWR.n3879 VPWR 339.046
R556 VPWR VPWR.n1373 339.046
R557 VPWR.n5016 VPWR 339.046
R558 VPWR.n8498 VPWR.n5860 337.3
R559 VPWR.n6393 VPWR.n6392 337.3
R560 VPWR.n1410 VPWR.n1409 337.3
R561 VPWR.n1939 VPWR.n1938 337.3
R562 VPWR VPWR.t72 334.012
R563 VPWR VPWR.t382 334.012
R564 VPWR VPWR.t539 334.012
R565 VPWR.t964 VPWR.t1141 330.654
R566 VPWR.t1705 VPWR.t774 330.654
R567 VPWR.t2313 VPWR.t2842 330.654
R568 VPWR.t1699 VPWR.t762 330.654
R569 VPWR.t1616 VPWR.t2503 330.654
R570 VPWR.t984 VPWR.t2284 330.654
R571 VPWR.t978 VPWR.t2927 330.654
R572 VPWR.t968 VPWR.t927 330.654
R573 VPWR.t2403 VPWR.t992 330.654
R574 VPWR.t1449 VPWR.t2521 330.654
R575 VPWR.n1846 VPWR.n1844 330.091
R576 VPWR.t2319 VPWR.t1490 327.298
R577 VPWR VPWR.t640 322.587
R578 VPWR.t557 VPWR 322.587
R579 VPWR.t12 VPWR 322.587
R580 VPWR.t175 VPWR 322.587
R581 VPWR.n934 VPWR.n933 321.457
R582 VPWR.t193 VPWR.t1960 318.906
R583 VPWR.t2488 VPWR.t9 318.906
R584 VPWR.n1179 VPWR.n1178 318.623
R585 VPWR.n1174 VPWR.n1173 318.623
R586 VPWR.n4710 VPWR.n4709 318.623
R587 VPWR.n4707 VPWR.n4706 318.623
R588 VPWR.n4704 VPWR.n4703 318.623
R589 VPWR.n528 VPWR.n527 318.623
R590 VPWR.n947 VPWR.n763 318.361
R591 VPWR.n2084 VPWR.n2083 318.361
R592 VPWR.n1782 VPWR.n1780 318.01
R593 VPWR.n1191 VPWR.n1190 317.599
R594 VPWR.n523 VPWR.n522 317.599
R595 VPWR.n941 VPWR.n940 317.348
R596 VPWR.n2638 VPWR.n2637 317.348
R597 VPWR.n1166 VPWR.n1165 317.115
R598 VPWR.n1162 VPWR.n1161 317.115
R599 VPWR.n1156 VPWR.n1155 317.115
R600 VPWR.n4726 VPWR.n4725 317.115
R601 VPWR.n5304 VPWR.n5303 317.115
R602 VPWR.n758 VPWR.n757 316.87
R603 VPWR.n2078 VPWR.n2077 316.87
R604 VPWR.n2067 VPWR.n2066 316.87
R605 VPWR.n7280 VPWR 316.668
R606 VPWR.n4701 VPWR.n4699 316.342
R607 VPWR.n9255 VPWR.n9254 316.132
R608 VPWR.n354 VPWR.n353 316.132
R609 VPWR.n1726 VPWR.n1725 316.132
R610 VPWR.t1302 VPWR.t3147 315.548
R611 VPWR.t1464 VPWR.t1466 315.548
R612 VPWR.t3133 VPWR.t1703 315.548
R613 VPWR.t2339 VPWR.t2953 315.548
R614 VPWR.t3191 VPWR.t3163 315.548
R615 VPWR.t1924 VPWR.t2678 315.548
R616 VPWR.n533 VPWR.n529 314.873
R617 VPWR.n4713 VPWR.n4712 314.776
R618 VPWR.n5952 VPWR.n5951 314.118
R619 VPWR.n1185 VPWR.n1183 313.921
R620 VPWR.n760 VPWR.n759 313.921
R621 VPWR.n951 VPWR.n948 313.921
R622 VPWR.n535 VPWR.n534 313.921
R623 VPWR.n2098 VPWR.n2096 313.921
R624 VPWR.n2089 VPWR.n2088 313.921
R625 VPWR.n51 VPWR.n50 313.849
R626 VPWR.n972 VPWR.n971 312.685
R627 VPWR.n967 VPWR.n755 312.685
R628 VPWR.n4730 VPWR.n4729 312.685
R629 VPWR.n540 VPWR.n539 312.685
R630 VPWR.n538 VPWR.n537 312.685
R631 VPWR.n2073 VPWR.n2072 312.685
R632 VPWR.n6348 VPWR.n6347 312.283
R633 VPWR.t3028 VPWR.t1548 312.192
R634 VPWR.t1553 VPWR.t3186 312.192
R635 VPWR.t394 VPWR.t2891 312.192
R636 VPWR.t2640 VPWR.t788 312.192
R637 VPWR VPWR.t3191 312.192
R638 VPWR.n3280 VPWR.n3279 311.957
R639 VPWR.n6058 VPWR.n6057 311.957
R640 VPWR.n7906 VPWR.n7905 311.957
R641 VPWR.n8203 VPWR.n8202 311.957
R642 VPWR.n351 VPWR.n350 311.957
R643 VPWR.n1006 VPWR.n1005 311.957
R644 VPWR.n983 VPWR.n982 311.957
R645 VPWR.n3534 VPWR.n3533 311.957
R646 VPWR.n3516 VPWR.n3515 311.957
R647 VPWR.n70 VPWR.n69 311.894
R648 VPWR.n51 VPWR.n49 311.894
R649 VPWR.n230 VPWR.n215 311.894
R650 VPWR.n7908 VPWR.n7907 311.894
R651 VPWR.n8873 VPWR.n8872 311.894
R652 VPWR.n8179 VPWR.n8177 311.894
R653 VPWR.n8142 VPWR.n8126 311.894
R654 VPWR.n8762 VPWR.n8737 311.894
R655 VPWR.n8621 VPWR.n8620 311.894
R656 VPWR.n5783 VPWR.n5782 311.894
R657 VPWR.n721 VPWR.n720 311.894
R658 VPWR.n409 VPWR.n408 311.894
R659 VPWR.n5605 VPWR.n463 311.894
R660 VPWR.n1382 VPWR.n1381 311.894
R661 VPWR.n2124 VPWR.n2123 311.894
R662 VPWR.n2310 VPWR.n2309 311.894
R663 VPWR.n2064 VPWR.n2062 311.894
R664 VPWR.n3575 VPWR.n3574 311.894
R665 VPWR.n7540 VPWR.n7539 311.575
R666 VPWR.n7059 VPWR.n7058 311.575
R667 VPWR.n7285 VPWR.n7284 311.575
R668 VPWR.n8604 VPWR.n8602 311.575
R669 VPWR.n5779 VPWR.n5778 311.575
R670 VPWR.n1558 VPWR.n1545 311.575
R671 VPWR.n2448 VPWR.n2431 311.575
R672 VPWR.n2230 VPWR.n2229 311.575
R673 VPWR.n2034 VPWR.n2033 311.575
R674 VPWR.n4508 VPWR.n4493 311.575
R675 VPWR.n7149 VPWR.n7148 311.575
R676 VPWR.n7154 VPWR.n7153 311.575
R677 VPWR.n593 VPWR.n592 311.118
R678 VPWR.n6602 VPWR.n6600 310.606
R679 VPWR.n102 VPWR.n100 310.551
R680 VPWR.n8912 VPWR.n8909 310.551
R681 VPWR.n5812 VPWR.n5809 310.551
R682 VPWR.n884 VPWR.n882 310.551
R683 VPWR.n4831 VPWR.n4830 310.551
R684 VPWR VPWR.t2586 310.512
R685 VPWR VPWR.t2202 310.512
R686 VPWR.t1789 VPWR 310.512
R687 VPWR.n6602 VPWR.n6601 309.955
R688 VPWR.n8898 VPWR.n8897 309.925
R689 VPWR.n6657 VPWR.n6656 309.729
R690 VPWR.n1024 VPWR.n1023 309.509
R691 VPWR.n2293 VPWR.n2292 309.241
R692 VPWR.n95 VPWR.n94 309.18
R693 VPWR.n244 VPWR.n243 309.18
R694 VPWR.n8320 VPWR.n8319 309.18
R695 VPWR.n1170 VPWR.n1169 309.18
R696 VPWR.n6647 VPWR.n6646 308.986
R697 VPWR.n1214 VPWR.n1213 308.986
R698 VPWR.t685 VPWR.t364 308.834
R699 VPWR.t554 VPWR.t625 308.834
R700 VPWR.t585 VPWR.t732 308.834
R701 VPWR VPWR.t2246 308.834
R702 VPWR.t545 VPWR.t367 308.834
R703 VPWR.n8125 VPWR.n8124 308.83
R704 VPWR.n8674 VPWR.n8673 308.83
R705 VPWR.n805 VPWR.n804 308.83
R706 VPWR.n445 VPWR.n444 308.69
R707 VPWR.n3219 VPWR.n3218 308.598
R708 VPWR.n6070 VPWR.n6066 308.598
R709 VPWR.n5963 VPWR.n5962 308.598
R710 VPWR.n8977 VPWR.n8976 308.598
R711 VPWR.n5948 VPWR.n5947 308.598
R712 VPWR.n843 VPWR.n842 308.598
R713 VPWR.n841 VPWR.n817 308.598
R714 VPWR.n1089 VPWR.n1088 308.598
R715 VPWR.n1018 VPWR.n1017 308.598
R716 VPWR.n1656 VPWR.n1655 308.598
R717 VPWR.n4915 VPWR.n4914 308.598
R718 VPWR.n4545 VPWR.n4544 308.598
R719 VPWR.n4234 VPWR.n4232 308.598
R720 VPWR.n3607 VPWR.n3606 308.598
R721 VPWR.n3613 VPWR.n3524 308.598
R722 VPWR.n3508 VPWR.n3507 308.598
R723 VPWR.n2814 VPWR.n2813 308.598
R724 VPWR.n4417 VPWR.n4415 308.363
R725 VPWR.n1543 VPWR.n1542 308.248
R726 VPWR.n6360 VPWR.n6359 308.149
R727 VPWR.n5450 VPWR.n5449 307.805
R728 VPWR.n110 VPWR.n109 307.604
R729 VPWR.n9186 VPWR.n37 307.604
R730 VPWR.n8990 VPWR.n8989 307.604
R731 VPWR.n7943 VPWR.n7942 307.604
R732 VPWR.n8911 VPWR.n8910 307.604
R733 VPWR.n8337 VPWR.n8336 307.604
R734 VPWR.n8290 VPWR.n5936 307.604
R735 VPWR.n5776 VPWR.n5775 307.604
R736 VPWR.n1150 VPWR.n1149 307.604
R737 VPWR.n5582 VPWR.n5581 307.604
R738 VPWR.n1483 VPWR.n1482 307.604
R739 VPWR.n4963 VPWR.n4962 307.604
R740 VPWR.n2176 VPWR.n2175 307.604
R741 VPWR.n2244 VPWR.n2243 307.604
R742 VPWR.n2663 VPWR.n2661 307.604
R743 VPWR.n2304 VPWR.n2303 307.604
R744 VPWR.n4465 VPWR.n4464 307.604
R745 VPWR.n2843 VPWR.n2842 307.604
R746 VPWR.n3725 VPWR.n3724 307.604
R747 VPWR.n3654 VPWR.n3653 307.604
R748 VPWR.n4263 VPWR.n4262 307.604
R749 VPWR.n2031 VPWR.n2027 307.558
R750 VPWR.n5422 VPWR.n5421 307.433
R751 VPWR.n3992 VPWR.n3991 307.308
R752 VPWR.n3893 VPWR.n3892 307.308
R753 VPWR.n3240 VPWR.n3236 307.308
R754 VPWR.n7648 VPWR.n7647 307.308
R755 VPWR.n6163 VPWR.n6162 307.308
R756 VPWR.n8755 VPWR.n8752 307.308
R757 VPWR.n6510 VPWR.n6506 307.308
R758 VPWR.n4807 VPWR.n4806 307.308
R759 VPWR.n3380 VPWR.n3379 307.308
R760 VPWR.t3001 VPWR.t1839 307.156
R761 VPWR.n1315 VPWR.n1314 306.659
R762 VPWR.n469 VPWR.n468 306.526
R763 VPWR.n3299 VPWR.n3298 305.882
R764 VPWR.n9174 VPWR.n9173 305.882
R765 VPWR.n6061 VPWR.n6059 305.882
R766 VPWR.n8022 VPWR.n8021 305.882
R767 VPWR.n9006 VPWR.n9005 305.882
R768 VPWR.n7927 VPWR.n7926 305.882
R769 VPWR.n8120 VPWR.n8118 305.882
R770 VPWR.n5945 VPWR.n5944 305.882
R771 VPWR.n8113 VPWR.n8112 305.882
R772 VPWR.n8778 VPWR.n8777 305.882
R773 VPWR.n8661 VPWR.n8660 305.882
R774 VPWR.n5811 VPWR.n5810 305.882
R775 VPWR.n997 VPWR.n996 305.882
R776 VPWR.n808 VPWR.n807 305.882
R777 VPWR.n437 VPWR.n436 305.882
R778 VPWR.n1467 VPWR.n1466 305.882
R779 VPWR.n1603 VPWR.n1602 305.882
R780 VPWR.n4947 VPWR.n4946 305.882
R781 VPWR.n2160 VPWR.n2159 305.882
R782 VPWR.n2259 VPWR.n2258 305.882
R783 VPWR.n2348 VPWR.n2347 305.882
R784 VPWR.n2091 VPWR.n2090 305.882
R785 VPWR.n4478 VPWR.n1999 305.882
R786 VPWR.n2859 VPWR.n2858 305.882
R787 VPWR.n3580 VPWR.n3579 305.882
R788 VPWR.n3713 VPWR.n3712 305.882
R789 VPWR.n2791 VPWR.n2790 305.882
R790 VPWR.n3520 VPWR.n3519 305.882
R791 VPWR.n3627 VPWR.n3625 305.882
R792 VPWR.t2648 VPWR.t451 305.478
R793 VPWR.t1671 VPWR.t113 305.478
R794 VPWR.n6711 VPWR.n6710 303.942
R795 VPWR.n821 VPWR.n819 303.942
R796 VPWR.n4732 VPWR.n4731 303.942
R797 VPWR.n4694 VPWR.n4692 303.942
R798 VPWR.n4679 VPWR.n4678 303.942
R799 VPWR.n5150 VPWR.n5149 303.942
R800 VPWR.n2708 VPWR.n2707 303.942
R801 VPWR.n6360 VPWR.n6358 302.661
R802 VPWR.n6705 VPWR.n6704 302.438
R803 VPWR.n821 VPWR.n820 302.438
R804 VPWR.n1306 VPWR.n1305 300.767
R805 VPWR.n4738 VPWR.n4737 300.474
R806 VPWR.t784 VPWR.t2999 300.442
R807 VPWR.n5932 VPWR.n5931 299.541
R808 VPWR.n6378 VPWR.n6377 299.205
R809 VPWR.n1304 VPWR.n1273 297.748
R810 VPWR VPWR.t2719 297.086
R811 VPWR.n290 VPWR.n289 296.56
R812 VPWR.t1862 VPWR.t1860 295.406
R813 VPWR.t2646 VPWR.t2644 295.406
R814 VPWR.n595 VPWR.n594 292.5
R815 VPWR.n629 VPWR.n628 292.5
R816 VPWR VPWR.t2864 288.693
R817 VPWR VPWR.t2987 287.014
R818 VPWR.t1661 VPWR.n8677 287.014
R819 VPWR.t875 VPWR 287.014
R820 VPWR.n2301 VPWR.t2256 287.014
R821 VPWR.t742 VPWR.t2373 284.113
R822 VPWR.t2264 VPWR.t2221 284.113
R823 VPWR.t2069 VPWR.t2291 284.113
R824 VPWR.t1956 VPWR.t1474 284.113
R825 VPWR.t3139 VPWR.t2474 284.113
R826 VPWR.t2466 VPWR.t312 283.658
R827 VPWR.t1282 VPWR.t373 281.979
R828 VPWR VPWR.t1522 281.979
R829 VPWR.t939 VPWR.t1486 281.154
R830 VPWR.t2820 VPWR.t2055 281.154
R831 VPWR.t2301 VPWR.t826 281.154
R832 VPWR.t3241 VPWR.t3205 281.154
R833 VPWR.t1892 VPWR.t844 281.154
R834 VPWR.t2901 VPWR.t1266 281.154
R835 VPWR VPWR.t128 280.3
R836 VPWR VPWR.t273 280.3
R837 VPWR VPWR.t347 280.3
R838 VPWR VPWR.t196 280.3
R839 VPWR VPWR.t222 280.3
R840 VPWR VPWR.t503 280.3
R841 VPWR VPWR.t136 280.3
R842 VPWR VPWR.t324 280.3
R843 VPWR VPWR.t122 280.3
R844 VPWR VPWR.t448 280.3
R845 VPWR VPWR.t216 280.3
R846 VPWR VPWR.t228 278.623
R847 VPWR VPWR.t477 278.623
R848 VPWR.t2230 VPWR.t1972 278.623
R849 VPWR.t1606 VPWR.t2159 276.943
R850 VPWR.t1737 VPWR.t1115 270.231
R851 VPWR.t2250 VPWR 266.873
R852 VPWR.t3067 VPWR 265.195
R853 VPWR.t2929 VPWR 265.195
R854 VPWR.t1874 VPWR 265.195
R855 VPWR.t2424 VPWR 263.517
R856 VPWR.t2626 VPWR 263.517
R857 VPWR.t1673 VPWR 263.517
R858 VPWR.t3087 VPWR 261.837
R859 VPWR VPWR.t424 261.837
R860 VPWR.t457 VPWR 261.837
R861 VPWR.t492 VPWR 261.837
R862 VPWR.t832 VPWR.t2966 260.437
R863 VPWR.t148 VPWR 260.159
R864 VPWR.t364 VPWR 260.159
R865 VPWR VPWR.t306 260.159
R866 VPWR.t542 VPWR 260.159
R867 VPWR.t712 VPWR 260.159
R868 VPWR VPWR.t57 260.159
R869 VPWR.t486 VPWR 260.159
R870 VPWR.t361 VPWR 260.159
R871 VPWR VPWR.t107 260.159
R872 VPWR VPWR.t706 260.159
R873 VPWR.t693 VPWR 260.159
R874 VPWR.t294 VPWR 260.159
R875 VPWR.t367 VPWR 260.159
R876 VPWR.t45 VPWR 260.159
R877 VPWR.t42 VPWR 260.159
R878 VPWR.t318 VPWR 260.159
R879 VPWR VPWR.t336 260.159
R880 VPWR VPWR.t358 260.159
R881 VPWR.t609 VPWR 260.159
R882 VPWR.t69 VPWR 260.159
R883 VPWR VPWR.t2297 258.481
R884 VPWR.t2004 VPWR.t909 258.481
R885 VPWR.t2775 VPWR 258.481
R886 VPWR.t2366 VPWR 258.481
R887 VPWR.t2490 VPWR 256.803
R888 VPWR VPWR.t600 256.803
R889 VPWR.t2858 VPWR 256.803
R890 VPWR.t2729 VPWR 256.803
R891 VPWR.t2356 VPWR.t3105 256.803
R892 VPWR VPWR.t903 256.803
R893 VPWR.t355 VPWR 256.803
R894 VPWR VPWR.t1530 255.125
R895 VPWR.t871 VPWR 255.125
R896 VPWR.t2375 VPWR.t2379 254.518
R897 VPWR.t2377 VPWR.t2375 254.518
R898 VPWR.t2373 VPWR.t2377 254.518
R899 VPWR.t2270 VPWR.t2266 254.518
R900 VPWR.t2266 VPWR.t2268 254.518
R901 VPWR.t2268 VPWR.t2264 254.518
R902 VPWR.t2071 VPWR.t2065 254.518
R903 VPWR.t2065 VPWR.t2067 254.518
R904 VPWR.t2067 VPWR.t2069 254.518
R905 VPWR.t1474 VPWR.t1470 254.518
R906 VPWR.t1470 VPWR.t1472 254.518
R907 VPWR.t1472 VPWR.t1476 254.518
R908 VPWR.t2474 VPWR.t2478 254.518
R909 VPWR.t2478 VPWR.t2472 254.518
R910 VPWR.t2472 VPWR.t2476 254.518
R911 VPWR VPWR.t2537 253.446
R912 VPWR.n7791 VPWR.t3388 252.006
R913 VPWR.n7691 VPWR.t3584 251.977
R914 VPWR.n6877 VPWR.t3507 251.977
R915 VPWR.n6799 VPWR.t3508 251.946
R916 VPWR.t1757 VPWR.t258 251.768
R917 VPWR.t2081 VPWR.t291 251.768
R918 VPWR.t506 VPWR.t3174 251.768
R919 VPWR.n5870 VPWR.t695 249.885
R920 VPWR.n1440 VPWR.t20 249.885
R921 VPWR.n2128 VPWR.t584 249.885
R922 VPWR.n1679 VPWR.t44 249.826
R923 VPWR.t1486 VPWR.t1488 248.599
R924 VPWR.t2055 VPWR.t2057 248.599
R925 VPWR.t2303 VPWR.t2301 248.599
R926 VPWR.t3243 VPWR.t3241 248.599
R927 VPWR.t844 VPWR.t842 248.599
R928 VPWR.t1266 VPWR.t1268 248.599
R929 VPWR.t3253 VPWR.n2567 248.411
R930 VPWR.n9138 VPWR.t673 246.541
R931 VPWR.n1126 VPWR.t679 246.411
R932 VPWR.n2423 VPWR.t338 246.411
R933 VPWR.t2877 VPWR.t1209 245.054
R934 VPWR.n3032 VPWR.t299 244.537
R935 VPWR.n6292 VPWR.t162 244.537
R936 VPWR.n5637 VPWR.t47 244.537
R937 VPWR.n5866 VPWR.t636 244.496
R938 VPWR.n4067 VPWR.t146 244.482
R939 VPWR.n5869 VPWR.t694 244.482
R940 VPWR.n1383 VPWR.t19 244.482
R941 VPWR.n2126 VPWR.t583 244.482
R942 VPWR.n2130 VPWR.t360 243.636
R943 VPWR.n2795 VPWR.t71 243.636
R944 VPWR.n2997 VPWR.t366 243.065
R945 VPWR.n8374 VPWR.t438 242.889
R946 VPWR.n3037 VPWR.t97 242.709
R947 VPWR.n2989 VPWR.t147 242.571
R948 VPWR.n3067 VPWR.t491 242.552
R949 VPWR.n6157 VPWR.t227 242.552
R950 VPWR.n6949 VPWR.t434 242.135
R951 VPWR.n6951 VPWR.t435 242.135
R952 VPWR.n7041 VPWR.t578 242.135
R953 VPWR.n7381 VPWR.t579 242.135
R954 VPWR.n7288 VPWR.t513 242.135
R955 VPWR.n7293 VPWR.t514 242.135
R956 VPWR.n7044 VPWR.t431 242.135
R957 VPWR.n7283 VPWR.t432 242.135
R958 VPWR.n3053 VPWR.t91 242.135
R959 VPWR.n3047 VPWR.t90 242.135
R960 VPWR.n3251 VPWR.t188 242.135
R961 VPWR.n3241 VPWR.t189 242.135
R962 VPWR.n3958 VPWR.t729 242.135
R963 VPWR.n4024 VPWR.t687 242.135
R964 VPWR.n4016 VPWR.t365 242.135
R965 VPWR.n4106 VPWR.t734 242.135
R966 VPWR.n9195 VPWR.t242 242.135
R967 VPWR.n41 VPWR.t618 242.135
R968 VPWR.n42 VPWR.t619 242.135
R969 VPWR.n43 VPWR.t256 242.135
R970 VPWR.n48 VPWR.t257 242.135
R971 VPWR.n9151 VPWR.t564 242.135
R972 VPWR.n57 VPWR.t565 242.135
R973 VPWR.n62 VPWR.t453 242.135
R974 VPWR.n59 VPWR.t672 242.135
R975 VPWR.n6067 VPWR.t238 242.135
R976 VPWR.n6075 VPWR.t239 242.135
R977 VPWR.n6103 VPWR.t598 242.135
R978 VPWR.n6063 VPWR.t599 242.135
R979 VPWR.n7710 VPWR.t77 242.135
R980 VPWR.n9062 VPWR.t575 242.135
R981 VPWR.n193 VPWR.t576 242.135
R982 VPWR.n283 VPWR.t65 242.135
R983 VPWR.n210 VPWR.t206 242.135
R984 VPWR.n212 VPWR.t207 242.135
R985 VPWR.n7901 VPWR.t536 242.135
R986 VPWR.n6217 VPWR.t573 242.135
R987 VPWR.n8925 VPWR.t562 242.135
R988 VPWR.n8867 VPWR.t410 242.135
R989 VPWR.n8868 VPWR.t411 242.135
R990 VPWR.n6740 VPWR.t263 242.135
R991 VPWR.n8151 VPWR.t67 242.135
R992 VPWR.n8122 VPWR.t68 242.135
R993 VPWR.n5937 VPWR.t499 242.135
R994 VPWR.n5943 VPWR.t500 242.135
R995 VPWR.n5924 VPWR.t115 242.135
R996 VPWR.n5928 VPWR.t194 242.135
R997 VPWR.n5930 VPWR.t195 242.135
R998 VPWR.n8196 VPWR.t371 242.135
R999 VPWR.n8110 VPWR.t372 242.135
R1000 VPWR.n8786 VPWR.t259 242.135
R1001 VPWR.n8732 VPWR.t260 242.135
R1002 VPWR.n8757 VPWR.t689 242.135
R1003 VPWR.n8739 VPWR.t690 242.135
R1004 VPWR.n8629 VPWR.t657 242.135
R1005 VPWR.n8614 VPWR.t650 242.135
R1006 VPWR.n8619 VPWR.t651 242.135
R1007 VPWR.n8467 VPWR.t569 242.135
R1008 VPWR.n8484 VPWR.t570 242.135
R1009 VPWR.n8457 VPWR.t141 242.135
R1010 VPWR.n8499 VPWR.t220 242.135
R1011 VPWR.n8537 VPWR.t221 242.135
R1012 VPWR.n6421 VPWR.t437 242.135
R1013 VPWR.n6357 VPWR.t50 242.135
R1014 VPWR.n6540 VPWR.t707 242.135
R1015 VPWR.n6470 VPWR.t708 242.135
R1016 VPWR.n6501 VPWR.t277 242.135
R1017 VPWR.n6511 VPWR.t278 242.135
R1018 VPWR.n1196 VPWR.t37 242.135
R1019 VPWR.n386 VPWR.t38 242.135
R1020 VPWR.n725 VPWR.t510 242.135
R1021 VPWR.n1132 VPWR.t511 242.135
R1022 VPWR.n1121 VPWR.t678 242.135
R1023 VPWR.n835 VPWR.t596 242.135
R1024 VPWR.n1025 VPWR.t653 242.135
R1025 VPWR.n753 VPWR.t654 242.135
R1026 VPWR.n868 VPWR.t736 242.135
R1027 VPWR.n765 VPWR.t737 242.135
R1028 VPWR.n953 VPWR.t475 242.135
R1029 VPWR.n761 VPWR.t476 242.135
R1030 VPWR.n812 VPWR.t159 242.135
R1031 VPWR.n641 VPWR.t389 242.135
R1032 VPWR.n692 VPWR.t390 242.135
R1033 VPWR.n494 VPWR.t459 242.135
R1034 VPWR.n5458 VPWR.t295 242.135
R1035 VPWR.n5462 VPWR.t296 242.135
R1036 VPWR.n5628 VPWR.t46 242.135
R1037 VPWR.n407 VPWR.t608 242.135
R1038 VPWR.n464 VPWR.t465 242.135
R1039 VPWR.n5467 VPWR.t546 242.135
R1040 VPWR.n490 VPWR.t547 242.135
R1041 VPWR.n1293 VPWR.t604 242.135
R1042 VPWR.n1274 VPWR.t605 242.135
R1043 VPWR.n4772 VPWR.t191 242.135
R1044 VPWR.n4785 VPWR.t192 242.135
R1045 VPWR.n1677 VPWR.t43 242.135
R1046 VPWR.n553 VPWR.t493 242.135
R1047 VPWR.n548 VPWR.t494 242.135
R1048 VPWR.n1591 VPWR.t717 242.135
R1049 VPWR.n2555 VPWR.t413 242.135
R1050 VPWR.n2564 VPWR.t414 242.135
R1051 VPWR.n4912 VPWR.t41 242.135
R1052 VPWR.n4919 VPWR.t404 242.135
R1053 VPWR.n4921 VPWR.t405 242.135
R1054 VPWR.n1897 VPWR.t614 242.135
R1055 VPWR.n5014 VPWR.t401 242.135
R1056 VPWR.n1963 VPWR.t402 242.135
R1057 VPWR.n5131 VPWR.t647 242.135
R1058 VPWR.n1839 VPWR.t648 242.135
R1059 VPWR.n2137 VPWR.t359 242.135
R1060 VPWR.n2473 VPWR.t179 242.135
R1061 VPWR.n2478 VPWR.t180 242.135
R1062 VPWR.n2457 VPWR.t461 242.135
R1063 VPWR.n2460 VPWR.t462 242.135
R1064 VPWR.n2466 VPWR.t337 242.135
R1065 VPWR.n4466 VPWR.t380 242.135
R1066 VPWR.n2004 VPWR.t381 242.135
R1067 VPWR.n2719 VPWR.t610 242.135
R1068 VPWR.n2373 VPWR.t201 242.135
R1069 VPWR.n2058 VPWR.t265 242.135
R1070 VPWR.n2047 VPWR.t266 242.135
R1071 VPWR.n4435 VPWR.t289 242.135
R1072 VPWR.n4451 VPWR.t290 242.135
R1073 VPWR.n4537 VPWR.t314 242.135
R1074 VPWR.n4486 VPWR.t165 242.135
R1075 VPWR.n2932 VPWR.t621 242.135
R1076 VPWR.n3624 VPWR.t507 242.135
R1077 VPWR.n3631 VPWR.t508 242.135
R1078 VPWR.n3584 VPWR.t532 242.135
R1079 VPWR.n3526 VPWR.t533 242.135
R1080 VPWR.n3726 VPWR.t34 242.135
R1081 VPWR.n3504 VPWR.t35 242.135
R1082 VPWR.n3396 VPWR.t419 242.135
R1083 VPWR.n3406 VPWR.t420 242.135
R1084 VPWR.n3419 VPWR.t55 242.135
R1085 VPWR.n3495 VPWR.t56 242.135
R1086 VPWR.n2817 VPWR.t70 242.135
R1087 VPWR.n7218 VPWR.t471 242.135
R1088 VPWR.n7130 VPWR.t470 242.135
R1089 VPWR.n7074 VPWR.t28 242.135
R1090 VPWR.n7050 VPWR.t29 242.135
R1091 VPWR.n2020 VPWR.t611 242.133
R1092 VPWR.n4532 VPWR.t164 242.133
R1093 VPWR.n2886 VPWR.t622 242.133
R1094 VPWR VPWR.t766 240.018
R1095 VPWR.t1740 VPWR 240.018
R1096 VPWR.t1890 VPWR.t104 238.339
R1097 VPWR.t1321 VPWR.t1223 238.339
R1098 VPWR.n3201 VPWR.t3358 236.891
R1099 VPWR.n1684 VPWR.t3433 236.891
R1100 VPWR.n4635 VPWR.t517 236.755
R1101 VPWR.t863 VPWR.t1657 236.661
R1102 VPWR.t1277 VPWR.t1903 234.982
R1103 VPWR.n6109 VPWR.t1555 234.982
R1104 VPWR.t2869 VPWR 234.982
R1105 VPWR.t1389 VPWR.t2570 234.982
R1106 VPWR.n9049 VPWR.t2490 234.982
R1107 VPWR.t1626 VPWR.t1663 234.982
R1108 VPWR.t2487 VPWR.t2206 234.982
R1109 VPWR.n1204 VPWR.t1968 234.982
R1110 VPWR.t2211 VPWR.t1841 234.982
R1111 VPWR.t3286 VPWR.t1048 234.982
R1112 VPWR.n559 VPWR.t1405 234.982
R1113 VPWR.t2595 VPWR.t1153 234.982
R1114 VPWR.t1159 VPWR.t83 234.982
R1115 VPWR.t1821 VPWR.t2263 234.982
R1116 VPWR.t1751 VPWR.t3158 234.982
R1117 VPWR.n3674 VPWR.t2354 234.982
R1118 VPWR.t2280 VPWR.t2358 234.982
R1119 VPWR.n1834 VPWR.t85 234.727
R1120 VPWR.n7159 VPWR.t176 234.554
R1121 VPWR.n7156 VPWR.t177 234.554
R1122 VPWR.n7562 VPWR.t641 234.554
R1123 VPWR.n7527 VPWR.t642 234.554
R1124 VPWR.n7531 VPWR.t719 234.554
R1125 VPWR.n7528 VPWR.t720 234.554
R1126 VPWR.n7299 VPWR.t558 234.554
R1127 VPWR.n7330 VPWR.t559 234.554
R1128 VPWR.n3277 VPWR.t283 234.554
R1129 VPWR.n3233 VPWR.t284 234.554
R1130 VPWR.n7122 VPWR.t13 234.554
R1131 VPWR.n7119 VPWR.t14 234.554
R1132 VPWR.n2992 VPWR.t106 233.311
R1133 VPWR.n3148 VPWR.t589 233.311
R1134 VPWR.n3057 VPWR.t253 233.311
R1135 VPWR.n3029 VPWR.t130 233.311
R1136 VPWR.n4102 VPWR.t702 233.311
R1137 VPWR.n4097 VPWR.t274 233.311
R1138 VPWR.n3247 VPWR.t343 233.311
R1139 VPWR.n3243 VPWR.t155 233.311
R1140 VPWR.n78 VPWR.t700 233.311
R1141 VPWR.n75 VPWR.t229 233.311
R1142 VPWR.n66 VPWR.t423 233.311
R1143 VPWR.n7644 VPWR.t502 233.311
R1144 VPWR.n7641 VPWR.t16 233.311
R1145 VPWR.n7652 VPWR.t2 233.311
R1146 VPWR.n6016 VPWR.t335 233.311
R1147 VPWR.n6275 VPWR.t349 233.311
R1148 VPWR.n6166 VPWR.t553 233.311
R1149 VPWR.n6173 VPWR.t302 233.311
R1150 VPWR.n6169 VPWR.t520 233.311
R1151 VPWR.n221 VPWR.t479 233.311
R1152 VPWR.n218 VPWR.t721 233.311
R1153 VPWR.n8296 VPWR.t524 233.311
R1154 VPWR.n8879 VPWR.t198 233.311
R1155 VPWR.n8876 VPWR.t208 233.311
R1156 VPWR.n6654 VPWR.t131 233.311
R1157 VPWR.n8147 VPWR.t8 233.311
R1158 VPWR.n6593 VPWR.t74 233.311
R1159 VPWR.n6590 VPWR.t78 233.311
R1160 VPWR.n8745 VPWR.t724 233.311
R1161 VPWR.n8741 VPWR.t223 233.311
R1162 VPWR.n5875 VPWR.t233 233.311
R1163 VPWR.n8617 VPWR.t61 233.311
R1164 VPWR.n6497 VPWR.t616 233.311
R1165 VPWR.n6493 VPWR.t87 233.311
R1166 VPWR.n6486 VPWR.t268 233.311
R1167 VPWR.n5790 VPWR.t505 233.311
R1168 VPWR.n5787 VPWR.t738 233.311
R1169 VPWR.n728 VPWR.t185 233.311
R1170 VPWR.n802 VPWR.t250 233.311
R1171 VPWR.n607 VPWR.t384 233.311
R1172 VPWR.n604 VPWR.t623 233.311
R1173 VPWR.n597 VPWR.t316 233.311
R1174 VPWR.n1444 VPWR.t639 233.311
R1175 VPWR.n417 VPWR.t138 233.311
R1176 VPWR.n414 VPWR.t537 233.311
R1177 VPWR.n1281 VPWR.t731 233.311
R1178 VPWR.n1278 VPWR.t416 233.311
R1179 VPWR.n1289 VPWR.t272 233.311
R1180 VPWR.n4799 VPWR.t659 233.311
R1181 VPWR.n4795 VPWR.t325 233.311
R1182 VPWR.n1551 VPWR.t519 233.311
R1183 VPWR.n1547 VPWR.t203 233.311
R1184 VPWR.n531 VPWR.t174 233.311
R1185 VPWR.n1906 VPWR.t697 233.311
R1186 VPWR.n4927 VPWR.t664 233.311
R1187 VPWR.n4923 VPWR.t123 233.311
R1188 VPWR.n1842 VPWR.t485 233.311
R1189 VPWR.n2118 VPWR.t582 233.311
R1190 VPWR.n2438 VPWR.t541 233.311
R1191 VPWR.n2435 VPWR.t725 233.311
R1192 VPWR.n2220 VPWR.t329 233.311
R1193 VPWR.n2216 VPWR.t566 233.311
R1194 VPWR.n2014 VPWR.t630 233.311
R1195 VPWR.n2029 VPWR.t53 233.311
R1196 VPWR.n2025 VPWR.t281 233.311
R1197 VPWR.n2011 VPWR.t526 233.311
R1198 VPWR.n4501 VPWR.t450 233.311
R1199 VPWR.n4498 VPWR.t691 233.311
R1200 VPWR.n2895 VPWR.t218 233.311
R1201 VPWR.n2891 VPWR.t472 233.311
R1202 VPWR.n3376 VPWR.t82 233.311
R1203 VPWR.n3373 VPWR.t350 233.311
R1204 VPWR.n3384 VPWR.t354 233.311
R1205 VPWR.n3511 VPWR.t467 233.311
R1206 VPWR.t597 VPWR.t2850 233.304
R1207 VPWR.t680 VPWR.t1361 233.304
R1208 VPWR.t66 VPWR.t2751 233.304
R1209 VPWR.t409 VPWR.t1367 233.304
R1210 VPWR.t2854 VPWR.t649 233.304
R1211 VPWR.t956 VPWR.t442 233.304
R1212 VPWR VPWR.t2601 233.304
R1213 VPWR.t303 VPWR.t333 231.625
R1214 VPWR.n58 VPWR.t671 231.625
R1215 VPWR.t2800 VPWR 231.625
R1216 VPWR.t905 VPWR.t294 231.625
R1217 VPWR.t836 VPWR.t874 231.625
R1218 VPWR.n7488 VPWR.t3574 230.734
R1219 VPWR.n7600 VPWR.t3580 230.734
R1220 VPWR.n7416 VPWR.t3506 230.734
R1221 VPWR.n3830 VPWR.t3586 230.734
R1222 VPWR.n3191 VPWR.t3397 230.734
R1223 VPWR.n3938 VPWR.t3478 230.734
R1224 VPWR.n3896 VPWR.t3380 230.734
R1225 VPWR.n4040 VPWR.t3535 230.734
R1226 VPWR.n4030 VPWR.t3546 230.734
R1227 VPWR.n4083 VPWR.t3461 230.734
R1228 VPWR.n4082 VPWR.t3521 230.734
R1229 VPWR.n3319 VPWR.t3405 230.734
R1230 VPWR.n7744 VPWR.t3427 230.734
R1231 VPWR.n7666 VPWR.t3499 230.734
R1232 VPWR.n7775 VPWR.t3540 230.734
R1233 VPWR.n7801 VPWR.t3341 230.734
R1234 VPWR.n7830 VPWR.t3536 230.734
R1235 VPWR.n6005 VPWR.t3369 230.734
R1236 VPWR.n6035 VPWR.t3424 230.734
R1237 VPWR.n8027 VPWR.t3404 230.734
R1238 VPWR.n9057 VPWR.t3484 230.734
R1239 VPWR.n8978 VPWR.t3481 230.734
R1240 VPWR.n8997 VPWR.t3333 230.734
R1241 VPWR.n7939 VPWR.t3344 230.734
R1242 VPWR.n6245 VPWR.t3524 230.734
R1243 VPWR.n6281 VPWR.t3434 230.734
R1244 VPWR.n6304 VPWR.t3354 230.734
R1245 VPWR.n8272 VPWR.t3544 230.734
R1246 VPWR.n6714 VPWR.t3501 230.734
R1247 VPWR.n6743 VPWR.t3362 230.734
R1248 VPWR.n6772 VPWR.t3537 230.734
R1249 VPWR.n6626 VPWR.t3459 230.734
R1250 VPWR.n8470 VPWR.t3477 230.734
R1251 VPWR.n6389 VPWR.t3516 230.734
R1252 VPWR.n6416 VPWR.t3350 230.734
R1253 VPWR.n1502 VPWR.t3385 230.734
R1254 VPWR.n5645 VPWR.t3392 230.734
R1255 VPWR.n5622 VPWR.t3370 230.734
R1256 VPWR.n5512 VPWR.t3500 230.734
R1257 VPWR.n5478 VPWR.t3485 230.734
R1258 VPWR.n1475 VPWR.t3416 230.734
R1259 VPWR.n1272 VPWR.t3560 230.734
R1260 VPWR.n4789 VPWR.t3480 230.734
R1261 VPWR.n4782 VPWR.t3355 230.734
R1262 VPWR.n5265 VPWR.t3346 230.734
R1263 VPWR.n1694 VPWR.t3449 230.734
R1264 VPWR.n1650 VPWR.t3342 230.734
R1265 VPWR.n2170 VPWR.t3555 230.734
R1266 VPWR.n2711 VPWR.t3383 230.734
R1267 VPWR.n4362 VPWR.t3363 230.734
R1268 VPWR.n2353 VPWR.t3365 230.734
R1269 VPWR.n4521 VPWR.t3562 230.734
R1270 VPWR.n2912 VPWR.t3389 230.734
R1271 VPWR.n2912 VPWR.t3510 230.734
R1272 VPWR.n4233 VPWR.t3386 230.734
R1273 VPWR.n2846 VPWR.t3582 230.734
R1274 VPWR.n3605 VPWR.t3470 230.734
R1275 VPWR.n3707 VPWR.t3576 230.734
R1276 VPWR.n2810 VPWR.t3407 230.734
R1277 VPWR.n3650 VPWR.t3550 230.734
R1278 VPWR.n2786 VPWR.t3547 230.734
R1279 VPWR.n7090 VPWR.t3437 230.734
R1280 VPWR.t2552 VPWR.t522 228.269
R1281 VPWR.n2692 VPWR.t2331 228.269
R1282 VPWR VPWR.t2385 226.59
R1283 VPWR.n6123 VPWR.t3504 224.883
R1284 VPWR.n6254 VPWR.t3578 224.883
R1285 VPWR.t718 VPWR 221.964
R1286 VPWR.n6943 VPWR 221.964
R1287 VPWR.n7281 VPWR 221.964
R1288 VPWR VPWR.n7280 221.964
R1289 VPWR VPWR.n7279 221.964
R1290 VPWR VPWR.t1807 221.555
R1291 VPWR.t2311 VPWR.t652 221.555
R1292 VPWR VPWR.t1334 219.876
R1293 VPWR VPWR.t1667 219.876
R1294 VPWR.n6955 VPWR 219.004
R1295 VPWR VPWR.t3060 216.519
R1296 VPWR.t1328 VPWR 216.519
R1297 VPWR.t1500 VPWR.t3113 214.841
R1298 VPWR.t2484 VPWR.t1117 213.163
R1299 VPWR.t885 VPWR.t2038 213.084
R1300 VPWR.t3278 VPWR 211.484
R1301 VPWR VPWR.t2293 209.806
R1302 VPWR VPWR.t2822 209.806
R1303 VPWR VPWR.t2858 209.806
R1304 VPWR.t709 VPWR.t2911 209.806
R1305 VPWR.t1313 VPWR 209.806
R1306 VPWR VPWR.t1139 209.806
R1307 VPWR.t2011 VPWR.t24 209.806
R1308 VPWR.n4708 VPWR.t2661 209.107
R1309 VPWR.t2391 VPWR 208.127
R1310 VPWR VPWR.t776 208.127
R1311 VPWR VPWR.t3109 208.127
R1312 VPWR.t3107 VPWR 208.127
R1313 VPWR VPWR.t3111 208.127
R1314 VPWR.n1766 VPWR.t769 207.464
R1315 VPWR VPWR.t3304 206.45
R1316 VPWR VPWR.t2972 206.45
R1317 VPWR VPWR.t1980 206.45
R1318 VPWR VPWR.t2648 206.45
R1319 VPWR.t935 VPWR.t421 206.45
R1320 VPWR VPWR.t2674 206.45
R1321 VPWR VPWR.t1990 206.45
R1322 VPWR VPWR.t63 206.45
R1323 VPWR VPWR.t3042 206.45
R1324 VPWR.t1783 VPWR 206.45
R1325 VPWR VPWR.t921 206.45
R1326 VPWR.t1391 VPWR 206.45
R1327 VPWR VPWR.t3199 206.45
R1328 VPWR.t1119 VPWR 206.45
R1329 VPWR VPWR.t2978 206.45
R1330 VPWR VPWR.t1922 206.45
R1331 VPWR VPWR.t1926 206.45
R1332 VPWR VPWR.t2963 206.45
R1333 VPWR.t954 VPWR 206.45
R1334 VPWR.t1151 VPWR 206.45
R1335 VPWR VPWR.t2694 206.45
R1336 VPWR.t903 VPWR 204.77
R1337 VPWR VPWR.t996 204.77
R1338 VPWR VPWR.t309 203.093
R1339 VPWR VPWR.t330 203.093
R1340 VPWR.t534 VPWR 203.093
R1341 VPWR VPWR.t344 203.093
R1342 VPWR VPWR.t2393 203.093
R1343 VPWR VPWR.t824 203.093
R1344 VPWR.t1165 VPWR 203.093
R1345 VPWR.t178 VPWR 203.093
R1346 VPWR.t1809 VPWR 203.093
R1347 VPWR.t2796 VPWR 203.093
R1348 VPWR.t3082 VPWR.t865 201.413
R1349 VPWR.t1195 VPWR.t1495 201.413
R1350 VPWR.t1655 VPWR.t3225 199.736
R1351 VPWR.n1930 VPWR.t2945 198.577
R1352 VPWR.n7535 VPWR.t2380 197.762
R1353 VPWR.n7372 VPWR.t2271 197.762
R1354 VPWR.n7052 VPWR.t2072 197.762
R1355 VPWR.n6588 VPWR.t3328 197.762
R1356 VPWR.n8608 VPWR.t3098 197.762
R1357 VPWR.n1554 VPWR.t1231 197.762
R1358 VPWR.n2223 VPWR.t2025 197.762
R1359 VPWR.n2035 VPWR.t1570 197.762
R1360 VPWR.n4496 VPWR.t2192 197.762
R1361 VPWR.n7150 VPWR.t1477 197.762
R1362 VPWR.n7155 VPWR.t2477 197.762
R1363 VPWR.n1297 VPWR.t3270 197.391
R1364 VPWR.n3266 VPWR.t3274 197.286
R1365 VPWR.n6054 VPWR.t1356 197.286
R1366 VPWR.n7904 VPWR.t3260 197.286
R1367 VPWR.n8149 VPWR.t2792 197.286
R1368 VPWR.n5952 VPWR.t1176 197.286
R1369 VPWR.n8684 VPWR.t2005 197.286
R1370 VPWR.n5762 VPWR.t2776 197.286
R1371 VPWR.n1138 VPWR.t1539 197.286
R1372 VPWR.n1574 VPWR.t1285 197.286
R1373 VPWR.n2036 VPWR.t3037 197.286
R1374 VPWR.n4456 VPWR.t2964 197.286
R1375 VPWR.n3499 VPWR.t955 197.286
R1376 VPWR.n3539 VPWR.t1140 197.286
R1377 VPWR.n2009 VPWR.t860 196.773
R1378 VPWR VPWR.t742 195.327
R1379 VPWR.t2221 VPWR 195.327
R1380 VPWR.t2291 VPWR 195.327
R1381 VPWR.t3119 VPWR 194.701
R1382 VPWR.n3514 VPWR.t1152 194.159
R1383 VPWR.n7953 VPWR.t2807 194.012
R1384 VPWR.n2833 VPWR.t1255 194.012
R1385 VPWR.n3987 VPWR.t1867 193.945
R1386 VPWR.n3887 VPWR.t1808 193.945
R1387 VPWR.n3250 VPWR.t2736 193.945
R1388 VPWR.n7648 VPWR.t2186 193.945
R1389 VPWR.n6163 VPWR.t2045 193.945
R1390 VPWR.n8738 VPWR.t2344 193.945
R1391 VPWR.n6500 VPWR.t2714 193.945
R1392 VPWR.n5780 VPWR.t1263 193.945
R1393 VPWR.n4792 VPWR.t2563 193.945
R1394 VPWR.n2449 VPWR.t2275 193.945
R1395 VPWR.n3380 VPWR.t3212 193.945
R1396 VPWR.n1137 VPWR.t1074 193.917
R1397 VPWR.n715 VPWR.t3157 193.917
R1398 VPWR.n4749 VPWR.t1060 193.917
R1399 VPWR.n5295 VPWR.t1062 193.917
R1400 VPWR.n9137 VPWR.t2649 193.72
R1401 VPWR.n9194 VPWR.t1556 193.72
R1402 VPWR.n195 VPWR.t2491 193.72
R1403 VPWR.n8968 VPWR.t2109 193.72
R1404 VPWR.n8850 VPWR.t2859 193.72
R1405 VPWR.n6670 VPWR.t1672 193.72
R1406 VPWR.n5934 VPWR.t2553 193.72
R1407 VPWR.n355 VPWR.t1734 193.72
R1408 VPWR.n995 VPWR.t1969 193.72
R1409 VPWR.n970 VPWR.t1855 193.72
R1410 VPWR.n799 VPWR.t3068 193.72
R1411 VPWR.n5684 VPWR.t2892 193.72
R1412 VPWR.n5562 VPWR.t3076 193.72
R1413 VPWR.n1375 VPWR.t904 193.72
R1414 VPWR.n1964 VPWR.t2979 193.72
R1415 VPWR.n2116 VPWR.t3256 193.72
R1416 VPWR.n2235 VPWR.t1648 193.72
R1417 VPWR.n2299 VPWR.t3301 193.72
R1418 VPWR.n3633 VPWR.t1293 193.72
R1419 VPWR.n2785 VPWR.t2695 193.72
R1420 VPWR.t3137 VPWR.t48 193.022
R1421 VPWR VPWR.t939 192.369
R1422 VPWR VPWR.t2820 192.369
R1423 VPWR.t2966 VPWR 192.369
R1424 VPWR.n5136 VPWR.t767 191.8
R1425 VPWR.n5100 VPWR.t1120 190.81
R1426 VPWR.n5100 VPWR.t1491 190.81
R1427 VPWR.n3161 VPWR.t1840 190.284
R1428 VPWR.n6530 VPWR.t3250 190.284
R1429 VPWR.n1849 VPWR.t1949 190.284
R1430 VPWR.n2277 VPWR.t2708 190.284
R1431 VPWR.n2048 VPWR.t1078 190.228
R1432 VPWR.t2038 VPWR 189.409
R1433 VPWR.n5879 VPWR.t2386 189.391
R1434 VPWR.n5141 VPWR.t1160 189.327
R1435 VPWR.t2658 VPWR 187.987
R1436 VPWR.n8444 VPWR.t3043 187.513
R1437 VPWR.n4648 VPWR.t3014 187.513
R1438 VPWR.n5022 VPWR.t1402 187.513
R1439 VPWR.n247 VPWR.t1210 187.083
R1440 VPWR.n2541 VPWR.t2365 187.083
R1441 VPWR.n3450 VPWR.t1925 187.083
R1442 VPWR.t1994 VPWR.t1992 184.63
R1443 VPWR.n8185 VPWR.t2554 184.63
R1444 VPWR.t3048 VPWR.t321 184.63
R1445 VPWR VPWR.t2968 184.63
R1446 VPWR.t3038 VPWR.t1740 184.63
R1447 VPWR VPWR.n3877 182.952
R1448 VPWR VPWR.t252 182.952
R1449 VPWR.t128 VPWR 182.952
R1450 VPWR.t104 VPWR 182.952
R1451 VPWR.n3878 VPWR 182.952
R1452 VPWR.t273 VPWR 182.952
R1453 VPWR.t333 VPWR 182.952
R1454 VPWR.t421 VPWR 182.952
R1455 VPWR.t228 VPWR 182.952
R1456 VPWR.t477 VPWR 182.952
R1457 VPWR.t196 VPWR 182.952
R1458 VPWR VPWR.t267 182.952
R1459 VPWR.t2993 VPWR.t2036 182.952
R1460 VPWR.t1225 VPWR.t1186 182.952
R1461 VPWR.t222 VPWR 182.952
R1462 VPWR.t503 VPWR 182.952
R1463 VPWR VPWR.t637 182.952
R1464 VPWR.n470 VPWR 182.952
R1465 VPWR.t136 VPWR 182.952
R1466 VPWR.t324 VPWR 182.952
R1467 VPWR.t1043 VPWR.t1393 182.952
R1468 VPWR.t122 VPWR 182.952
R1469 VPWR.t279 VPWR 182.952
R1470 VPWR.t628 VPWR 182.952
R1471 VPWR.t448 VPWR 182.952
R1472 VPWR VPWR.t466 182.952
R1473 VPWR.t216 VPWR 182.952
R1474 VPWR.t2077 VPWR.t1179 181.273
R1475 VPWR.t2747 VPWR.t2650 181.273
R1476 VPWR.t2804 VPWR.t1709 181.273
R1477 VPWR.t1359 VPWR.t2492 181.273
R1478 VPWR.t3081 VPWR.t1843 181.273
R1479 VPWR.t1689 VPWR.t1669 181.273
R1480 VPWR.t267 VPWR.t2199 181.273
R1481 VPWR.t2000 VPWR.t2800 181.273
R1482 VPWR VPWR.t2254 181.273
R1483 VPWR.t901 VPWR.t990 181.273
R1484 VPWR.t2828 VPWR.t3077 181.273
R1485 VPWR.t1286 VPWR.t982 181.273
R1486 VPWR.t2895 VPWR.t2165 181.273
R1487 VPWR.t3251 VPWR.t972 181.273
R1488 VPWR.t1115 VPWR.t2010 181.273
R1489 VPWR.t2523 VPWR.t2976 181.273
R1490 VPWR.t958 VPWR.t3302 181.273
R1491 VPWR.t2507 VPWR.t2961 181.273
R1492 VPWR.t952 VPWR.t980 181.273
R1493 VPWR.t966 VPWR.t1137 181.273
R1494 VPWR.t1294 VPWR.t2511 181.273
R1495 VPWR.t2505 VPWR.t2696 181.273
R1496 VPWR.t2527 VPWR.t1256 181.273
R1497 VPWR.n6127 VPWR 179.595
R1498 VPWR VPWR.n6642 179.595
R1499 VPWR.n6447 VPWR 179.595
R1500 VPWR.t231 VPWR 179.595
R1501 VPWR.n471 VPWR 179.595
R1502 VPWR.n5402 VPWR.n5401 179.131
R1503 VPWR.n2549 VPWR.n2189 179.131
R1504 VPWR.n6621 VPWR.n6620 178.359
R1505 VPWR.t3142 VPWR 177.916
R1506 VPWR.t2900 VPWR 177.916
R1507 VPWR.t865 VPWR.t1707 177.916
R1508 VPWR.t3131 VPWR 177.916
R1509 VPWR.t1701 VPWR.t3137 177.916
R1510 VPWR VPWR.t3235 177.916
R1511 VPWR.t1697 VPWR.t1169 177.916
R1512 VPWR.t2948 VPWR 177.916
R1513 VPWR.t1403 VPWR.t2942 177.916
R1514 VPWR.n6489 VPWR.n6488 176.733
R1515 VPWR.t3097 VPWR.t1733 176.238
R1516 VPWR.n3854 VPWR.n3853 175.834
R1517 VPWR.n2563 VPWR.n2187 175.834
R1518 VPWR.n3497 VPWR.n3496 175.834
R1519 VPWR.n1895 VPWR.n1893 175.43
R1520 VPWR.n5434 VPWR.n5433 174.595
R1521 VPWR.n5133 VPWR.n5132 174.595
R1522 VPWR.t929 VPWR 174.559
R1523 VPWR.t1495 VPWR.t1343 174.559
R1524 VPWR.t2020 VPWR 174.559
R1525 VPWR.t2816 VPWR 174.559
R1526 VPWR.n4414 VPWR.n4413 173.754
R1527 VPWR.t427 VPWR.t1866 172.881
R1528 VPWR.t1880 VPWR 172.881
R1529 VPWR VPWR.t2980 172.881
R1530 VPWR.t1353 VPWR 172.881
R1531 VPWR.t2093 VPWR.t2993 172.881
R1532 VPWR VPWR.t3030 172.881
R1533 VPWR.t2018 VPWR 172.881
R1534 VPWR.t1920 VPWR.t2787 172.881
R1535 VPWR.t2317 VPWR 172.881
R1536 VPWR.t925 VPWR 172.881
R1537 VPWR.n1924 VPWR.n1923 171.982
R1538 VPWR.n1919 VPWR.n1918 171.982
R1539 VPWR.n1788 VPWR.n1786 171.674
R1540 VPWR.n8595 VPWR.n8594 170.916
R1541 VPWR.n1428 VPWR.n1427 170.916
R1542 VPWR.n1911 VPWR.n1910 170.862
R1543 VPWR.n1835 VPWR.t3548 170.734
R1544 VPWR.n4643 VPWR.t3441 170.71
R1545 VPWR.n1817 VPWR.n1816 169.934
R1546 VPWR.n2991 VPWR.t3384 169.667
R1547 VPWR.n3147 VPWR.t3522 169.667
R1548 VPWR.n3056 VPWR.t3408 169.667
R1549 VPWR.n3028 VPWR.t3393 169.667
R1550 VPWR.n4096 VPWR.t3415 169.667
R1551 VPWR.n4101 VPWR.t3340 169.667
R1552 VPWR.n3242 VPWR.t3371 169.667
R1553 VPWR.n3246 VPWR.t3476 169.667
R1554 VPWR.n74 VPWR.t3399 169.667
R1555 VPWR.n77 VPWR.t3339 169.667
R1556 VPWR.n65 VPWR.t3495 169.667
R1557 VPWR.n7640 VPWR.t3338 169.667
R1558 VPWR.n7643 VPWR.t3528 169.667
R1559 VPWR.n7651 VPWR.t3360 169.667
R1560 VPWR.n6015 VPWR.t3472 169.667
R1561 VPWR.n6274 VPWR.t3483 169.667
R1562 VPWR.n6165 VPWR.t3542 169.667
R1563 VPWR.n6168 VPWR.t3518 169.667
R1564 VPWR.n6172 VPWR.t3455 169.667
R1565 VPWR.n217 VPWR.t3585 169.667
R1566 VPWR.n220 VPWR.t3520 169.667
R1567 VPWR.n8295 VPWR.t3462 169.667
R1568 VPWR.n8875 VPWR.t3509 169.667
R1569 VPWR.n8878 VPWR.t3345 169.667
R1570 VPWR.n6653 VPWR.t3515 169.667
R1571 VPWR.n8146 VPWR.t3543 169.667
R1572 VPWR.n6589 VPWR.t3444 169.667
R1573 VPWR.n6592 VPWR.t3559 169.667
R1574 VPWR.n8740 VPWR.t3410 169.667
R1575 VPWR.n8744 VPWR.t3469 169.667
R1576 VPWR.n5874 VPWR.t3552 169.667
R1577 VPWR.n8616 VPWR.t3356 169.667
R1578 VPWR.n6492 VPWR.t3366 169.667
R1579 VPWR.n6496 VPWR.t3419 169.667
R1580 VPWR.n6485 VPWR.t3428 169.667
R1581 VPWR.n5786 VPWR.t3533 169.667
R1582 VPWR.n5789 VPWR.t3387 169.667
R1583 VPWR.n727 VPWR.t3336 169.667
R1584 VPWR.n801 VPWR.t3361 169.667
R1585 VPWR.n603 VPWR.t3488 169.667
R1586 VPWR.n606 VPWR.t3348 169.667
R1587 VPWR.n596 VPWR.t3381 169.667
R1588 VPWR.n1443 VPWR.t3572 169.667
R1589 VPWR.n413 VPWR.t3446 169.667
R1590 VPWR.n416 VPWR.t3394 169.667
R1591 VPWR.n1277 VPWR.t3401 169.667
R1592 VPWR.n1280 VPWR.t3352 169.667
R1593 VPWR.n1288 VPWR.t3445 169.667
R1594 VPWR.n4794 VPWR.t3375 169.667
R1595 VPWR.n4798 VPWR.t3571 169.667
R1596 VPWR.n1546 VPWR.t3587 169.667
R1597 VPWR.n1550 VPWR.t3523 169.667
R1598 VPWR.n530 VPWR.t3391 169.667
R1599 VPWR.n1905 VPWR.t3498 169.667
R1600 VPWR.n4922 VPWR.t3563 169.667
R1601 VPWR.n4926 VPWR.t3494 169.667
R1602 VPWR.n1841 VPWR.t3436 169.667
R1603 VPWR.n2117 VPWR.t3465 169.667
R1604 VPWR.n2434 VPWR.t3513 169.667
R1605 VPWR.n2437 VPWR.t3450 169.667
R1606 VPWR.n2215 VPWR.t3517 169.667
R1607 VPWR.n2219 VPWR.t3378 169.667
R1608 VPWR.n2013 VPWR.t3486 169.667
R1609 VPWR.n2028 VPWR.t3539 169.667
R1610 VPWR.n2024 VPWR.t3364 169.667
R1611 VPWR.n2010 VPWR.t3503 169.667
R1612 VPWR.n4497 VPWR.t3568 169.667
R1613 VPWR.n4500 VPWR.t3422 169.667
R1614 VPWR.n2890 VPWR.t3490 169.667
R1615 VPWR.n2894 VPWR.t3349 169.667
R1616 VPWR.n3372 VPWR.t3443 169.667
R1617 VPWR.n3375 VPWR.t3567 169.667
R1618 VPWR.n3383 VPWR.t3398 169.667
R1619 VPWR.n3510 VPWR.t3489 169.667
R1620 VPWR.n5613 VPWR.n459 169.555
R1621 VPWR VPWR.t2163 169.524
R1622 VPWR.t1290 VPWR.t2094 169.524
R1623 VPWR.n4696 VPWR.n4695 169.44
R1624 VPWR.n7680 VPWR.n7678 169.032
R1625 VPWR.n6193 VPWR.n6191 169.032
R1626 VPWR.n986 VPWR.n985 169.028
R1627 VPWR.n545 VPWR.n544 169.028
R1628 VPWR.n543 VPWR.n542 169.028
R1629 VPWR.n6528 VPWR.n6527 169.017
R1630 VPWR.n1380 VPWR.n1379 169.017
R1631 VPWR.n4422 VPWR.n4421 169.017
R1632 VPWR.n719 VPWR.n718 168.91
R1633 VPWR.n1714 VPWR.n556 168.91
R1634 VPWR.n1929 VPWR.n1928 168.91
R1635 VPWR.n2314 VPWR.n2313 168.91
R1636 VPWR.n8049 VPWR.n8048 168.91
R1637 VPWR.n8138 VPWR.n8137 168.91
R1638 VPWR.n2308 VPWR.n2307 168.91
R1639 VPWR.n979 VPWR.n978 168.781
R1640 VPWR.n2043 VPWR.n2042 168.781
R1641 VPWR.n4739 VPWR.n4736 168.374
R1642 VPWR.n8179 VPWR.n8178 167.855
R1643 VPWR.t2204 VPWR.t1934 167.845
R1644 VPWR.t1517 VPWR.t157 167.845
R1645 VPWR.t606 VPWR.t1301 167.845
R1646 VPWR.n8053 VPWR.n8052 167.623
R1647 VPWR.n4680 VPWR.n4677 167.28
R1648 VPWR.n711 VPWR.n710 167.038
R1649 VPWR.n4701 VPWR.n4700 166.692
R1650 VPWR.n600 VPWR.n599 166.619
R1651 VPWR.n8424 VPWR.n5877 166.542
R1652 VPWR.n612 VPWR.n602 166.542
R1653 VPWR.n1892 VPWR.n1891 166.542
R1654 VPWR.n5119 VPWR.n5118 166.542
R1655 VPWR.n1087 VPWR.n1086 166.381
R1656 VPWR.n4361 VPWR.n4360 166.381
R1657 VPWR.n4441 VPWR.n4440 166.381
R1658 VPWR.n9204 VPWR.n30 166.363
R1659 VPWR.n8116 VPWR.n8114 166.363
R1660 VPWR.n7529 VPWR.t3526 166.282
R1661 VPWR.n7561 VPWR.t3497 166.282
R1662 VPWR.n7298 VPWR.t3473 166.282
R1663 VPWR.n3276 VPWR.t3452 166.282
R1664 VPWR.n7121 VPWR.t3545 166.282
R1665 VPWR.n7158 VPWR.t3337 166.282
R1666 VPWR.t3063 VPWR.t2727 166.167
R1667 VPWR.t1174 VPWR.t1205 166.167
R1668 VPWR.t1173 VPWR.t3021 166.167
R1669 VPWR.t774 VPWR.t944 166.167
R1670 VPWR.t1664 VPWR.t1723 166.167
R1671 VPWR.t1663 VPWR.t2053 166.167
R1672 VPWR.t1334 VPWR.t1720 166.167
R1673 VPWR.t1963 VPWR.t1819 166.167
R1674 VPWR.t1962 VPWR.t3308 166.167
R1675 VPWR.t2808 VPWR.t2487 166.167
R1676 VPWR.t1933 VPWR.t998 166.167
R1677 VPWR.t1007 VPWR.t2959 166.167
R1678 VPWR.t2115 VPWR.t2814 166.167
R1679 VPWR.t2112 VPWR.t3181 166.167
R1680 VPWR.t3276 VPWR.t1685 166.167
R1681 VPWR.t1791 VPWR.t1686 166.167
R1682 VPWR.t822 VPWR.t1757 166.167
R1683 VPWR.t951 VPWR.t1517 166.167
R1684 VPWR.t1037 VPWR.t2369 166.167
R1685 VPWR.t1036 VPWR.t1565 166.167
R1686 VPWR.t1816 VPWR.t1002 166.167
R1687 VPWR.t2670 VPWR.t2208 166.167
R1688 VPWR.t2778 VPWR.t2211 166.167
R1689 VPWR.t3044 VPWR.t3005 166.167
R1690 VPWR.t1298 VPWR.t1616 166.167
R1691 VPWR.t1301 VPWR.t2624 166.167
R1692 VPWR.t1748 VPWR.t1328 166.167
R1693 VPWR.t2306 VPWR.t917 166.167
R1694 VPWR.t2260 VPWR.t2081 166.167
R1695 VPWR.t2263 VPWR.t2283 166.167
R1696 VPWR.t1947 VPWR.t1809 166.167
R1697 VPWR.t1944 VPWR.t1506 166.167
R1698 VPWR.t780 VPWR.t1996 166.167
R1699 VPWR VPWR.t2167 166.167
R1700 VPWR.t2567 VPWR.t2531 166.167
R1701 VPWR.t1974 VPWR.t2796 166.167
R1702 VPWR.t1975 VPWR.t2914 166.167
R1703 VPWR.t2384 VPWR.t1449 166.167
R1704 VPWR.n7470 VPWR.n7469 165.767
R1705 VPWR.n6945 VPWR.n6944 165.767
R1706 VPWR.n7558 VPWR.n7557 165.767
R1707 VPWR.n7032 VPWR.n7031 165.767
R1708 VPWR.n7295 VPWR.n7294 165.767
R1709 VPWR.n3042 VPWR.n3041 165.767
R1710 VPWR.n4060 VPWR.n4059 165.767
R1711 VPWR.n4088 VPWR.n4087 165.767
R1712 VPWR.n3261 VPWR.n3260 165.767
R1713 VPWR.n72 VPWR.n71 165.767
R1714 VPWR.n214 VPWR.n213 165.767
R1715 VPWR.n8887 VPWR.n8886 165.767
R1716 VPWR.n8491 VPWR.n8490 165.767
R1717 VPWR.n8493 VPWR.n8492 165.767
R1718 VPWR.n5797 VPWR.n5784 165.767
R1719 VPWR.n411 VPWR.n410 165.767
R1720 VPWR.n403 VPWR.n402 165.767
R1721 VPWR.n5606 VPWR.n460 165.767
R1722 VPWR.n1782 VPWR.n1781 165.767
R1723 VPWR.n1715 VPWR.n555 165.767
R1724 VPWR.n2226 VPWR.n2225 165.767
R1725 VPWR.n2316 VPWR.n2315 165.767
R1726 VPWR.n4495 VPWR.n4494 165.767
R1727 VPWR.n3413 VPWR.n3412 165.767
R1728 VPWR.n7115 VPWR.n7114 165.767
R1729 VPWR.n7191 VPWR.n7190 165.767
R1730 VPWR.n3178 VPWR.n3177 165.72
R1731 VPWR.n54 VPWR.n53 165.72
R1732 VPWR.n6012 VPWR.n6011 165.72
R1733 VPWR.n8324 VPWR.n8323 165.72
R1734 VPWR.n8690 VPWR.n8689 165.72
R1735 VPWR.n8648 VPWR.n8647 165.72
R1736 VPWR.n5647 VPWR.n5646 165.72
R1737 VPWR.n1564 VPWR.n1563 165.72
R1738 VPWR.n5146 VPWR.n5145 165.72
R1739 VPWR.n2114 VPWR.n2113 165.72
R1740 VPWR.n2248 VPWR.n2247 165.72
R1741 VPWR.n3404 VPWR.n3401 165.72
R1742 VPWR.n1815 VPWR.n1814 165.681
R1743 VPWR.n7545 VPWR.n7544 165.369
R1744 VPWR.n7064 VPWR.n7063 165.369
R1745 VPWR.n7287 VPWR.n7286 165.369
R1746 VPWR.n3258 VPWR.n3235 165.369
R1747 VPWR.n6180 VPWR.n6179 165.369
R1748 VPWR.n8736 VPWR.n8735 165.369
R1749 VPWR.n8599 VPWR.n8596 165.369
R1750 VPWR.n2444 VPWR.n2433 165.369
R1751 VPWR.n7183 VPWR.n7182 165.369
R1752 VPWR.n7152 VPWR.n7151 165.369
R1753 VPWR.n8626 VPWR.n8625 165.202
R1754 VPWR.n1141 VPWR.n1140 164.843
R1755 VPWR.n5418 VPWR.n5417 164.843
R1756 VPWR.n4744 VPWR.n4743 164.843
R1757 VPWR.n2055 VPWR.n2053 164.843
R1758 VPWR.n1148 VPWR.n1147 164.596
R1759 VPWR.n9033 VPWR.n9032 164.558
R1760 VPWR.n4951 VPWR.n4950 164.558
R1761 VPWR.n2147 VPWR.n2146 164.558
R1762 VPWR.n3680 VPWR.n3678 164.558
R1763 VPWR.t36 VPWR.t1554 164.488
R1764 VPWR.t312 VPWR.t1945 164.488
R1765 VPWR.n8598 VPWR.n8597 164.215
R1766 VPWR.n1110 VPWR.n732 164.215
R1767 VPWR.n1041 VPWR.n1039 164.215
R1768 VPWR.n1389 VPWR.n1388 164.215
R1769 VPWR.n4662 VPWR.n4661 164.215
R1770 VPWR.n526 VPWR.n525 164.215
R1771 VPWR.n1943 VPWR.n1942 164.215
R1772 VPWR.n1853 VPWR.n1852 164.215
R1773 VPWR.n1832 VPWR.n1831 164.215
R1774 VPWR.n1830 VPWR.n1829 164.215
R1775 VPWR.n207 VPWR.n206 163.44
R1776 VPWR.n6523 VPWR.n6522 163.44
R1777 VPWR.n3418 VPWR.n3417 163.44
R1778 VPWR.n1291 VPWR.n1284 163.369
R1779 VPWR.n3146 VPWR.n3145 163.268
R1780 VPWR.n6733 VPWR.n6732 163.221
R1781 VPWR.n6344 VPWR.n6343 163.221
R1782 VPWR.t1903 VPWR.t964 162.81
R1783 VPWR.t2586 VPWR.t796 162.81
R1784 VPWR.t2850 VPWR.t1880 162.81
R1785 VPWR.t1608 VPWR.t1346 162.81
R1786 VPWR.t2980 VPWR.t1705 162.81
R1787 VPWR.t2842 VPWR.t1389 162.81
R1788 VPWR.t1361 VPWR.t1626 162.81
R1789 VPWR.t1520 VPWR.t1844 162.81
R1790 VPWR.t2717 VPWR.t2680 162.81
R1791 VPWR.t2206 VPWR.t2832 162.81
R1792 VPWR.t2844 VPWR.t1129 162.81
R1793 VPWR.t2751 VPWR.t1353 162.81
R1794 VPWR.t2554 VPWR.t2156 162.81
R1795 VPWR.t1238 VPWR.t2729 162.81
R1796 VPWR.t3030 VPWR.t2854 162.81
R1797 VPWR.t2755 VPWR.t2018 162.81
R1798 VPWR.t594 VPWR.t1936 162.81
R1799 VPWR.t1979 VPWR.t834 162.81
R1800 VPWR.t1940 VPWR.t1699 162.81
R1801 VPWR.t1369 VPWR.t3282 162.81
R1802 VPWR.t1841 VPWR.t956 162.81
R1803 VPWR.t2608 VPWR.t863 162.81
R1804 VPWR.t2838 VPWR.t3286 162.81
R1805 VPWR VPWR.t3313 162.81
R1806 VPWR.t3167 VPWR.t1197 162.81
R1807 VPWR.t2503 VPWR.t3201 162.81
R1808 VPWR.t1183 VPWR.t984 162.81
R1809 VPWR.t1153 VPWR.t978 162.81
R1810 VPWR.t974 VPWR.t1821 162.81
R1811 VPWR.t1203 VPWR.t1399 162.81
R1812 VPWR.t2509 VPWR.t2020 162.81
R1813 VPWR.t3158 VPWR.t968 162.81
R1814 VPWR.t988 VPWR.t1930 162.81
R1815 VPWR.t3231 VPWR.t2519 162.81
R1816 VPWR.t2517 VPWR.t2816 162.81
R1817 VPWR.t2521 VPWR.t925 162.81
R1818 VPWR.n4107 VPWR.n4095 162.47
R1819 VPWR.n3052 VPWR.n3051 162.47
R1820 VPWR.n3158 VPWR.n3157 162.47
R1821 VPWR.n3272 VPWR.n3271 162.47
R1822 VPWR.n9175 VPWR.n9172 162.47
R1823 VPWR.n6039 VPWR.n6038 162.47
R1824 VPWR.n7996 VPWR.n7988 162.47
R1825 VPWR.n6268 VPWR.n6267 162.47
R1826 VPWR.n6412 VPWR.n6352 162.47
R1827 VPWR.n1133 VPWR.n723 162.47
R1828 VPWR.n1123 VPWR.n726 162.47
R1829 VPWR.n1294 VPWR.n1276 162.47
R1830 VPWR.n5486 VPWR.n487 162.47
R1831 VPWR.n1665 VPWR.n1664 162.47
R1832 VPWR.n5308 VPWR.n5307 162.47
R1833 VPWR.n2468 VPWR.n2425 162.47
R1834 VPWR.n2459 VPWR.n2428 162.47
R1835 VPWR.n2430 VPWR.n2429 162.47
R1836 VPWR.n1962 VPWR.n1961 162.47
R1837 VPWR.n5105 VPWR.n5104 162.47
R1838 VPWR.n4488 VPWR.n4487 162.47
R1839 VPWR.n2375 VPWR.n2298 162.47
R1840 VPWR.n4459 VPWR.n4458 162.47
R1841 VPWR.n3392 VPWR.n3389 162.47
R1842 VPWR.n3741 VPWR.n3740 162.47
R1843 VPWR.n4429 VPWR.n2007 161.992
R1844 VPWR.n3998 VPWR.n3997 161.859
R1845 VPWR.n3900 VPWR.n3899 161.859
R1846 VPWR.n7659 VPWR.n7658 161.859
R1847 VPWR.n6607 VPWR.n6606 161.859
R1848 VPWR.n6491 VPWR.n6490 161.859
R1849 VPWR.n5777 VPWR.n5774 161.859
R1850 VPWR.n4813 VPWR.n4812 161.859
R1851 VPWR.n1565 VPWR.n1562 161.859
R1852 VPWR.n2234 VPWR.n2233 161.859
R1853 VPWR.n2682 VPWR.n2681 161.859
R1854 VPWR.n4491 VPWR.n4489 161.859
R1855 VPWR.n3391 VPWR.n3390 161.859
R1856 VPWR.n731 VPWR.n730 161.817
R1857 VPWR.t3073 VPWR.t2733 161.131
R1858 VPWR.t1805 VPWR.t1113 161.131
R1859 VPWR.t1872 VPWR.t2765 161.131
R1860 VPWR.t2014 VPWR.t2179 161.131
R1861 VPWR.t424 VPWR.t3071 161.131
R1862 VPWR.t2987 VPWR.t1823 161.131
R1863 VPWR.t1311 VPWR 161.131
R1864 VPWR.t3269 VPWR.t603 161.131
R1865 VPWR.t2719 VPWR.t2723 161.131
R1866 VPWR.t2412 VPWR.t1542 161.131
R1867 VPWR.t770 VPWR.t2556 161.131
R1868 VPWR.t3329 VPWR.t1401 161.131
R1869 VPWR.t3056 VPWR.t1573 161.131
R1870 VPWR.t1117 VPWR.t1195 161.131
R1871 VPWR.t2335 VPWR.t2193 161.131
R1872 VPWR.n1435 VPWR.n1385 160.918
R1873 VPWR.n1935 VPWR.n1934 160.918
R1874 VPWR.n2699 VPWR.n2698 160.918
R1875 VPWR.n4401 VPWR.n4400 160.918
R1876 VPWR.n4378 VPWR.n4377 160.918
R1877 VPWR.n4432 VPWR.n4430 160.918
R1878 VPWR.n1779 VPWR.n1778 160.649
R1879 VPWR.n1911 VPWR.t1456 160.279
R1880 VPWR.n3159 VPWR.n3156 160.143
R1881 VPWR.n5106 VPWR.n5103 160.143
R1882 VPWR.n2480 VPWR.n2477 160.143
R1883 VPWR.n2263 VPWR.n2262 160.143
R1884 VPWR.n1411 VPWR.t1304 159.46
R1885 VPWR.n2728 VPWR.t1983 159.46
R1886 VPWR.n4446 VPWR.t3120 159.46
R1887 VPWR.n1034 VPWR.t1125 159.46
R1888 VPWR.t1715 VPWR.t1468 159.452
R1889 VPWR VPWR.t1608 159.452
R1890 VPWR.t1466 VPWR.t1282 159.452
R1891 VPWR.t900 VPWR.t2702 159.452
R1892 VPWR.t3129 VPWR.t2482 159.452
R1893 VPWR.t1288 VPWR.t1502 159.452
R1894 VPWR VPWR.t1693 159.452
R1895 VPWR.t758 VPWR.t2525 159.452
R1896 VPWR.t1651 VPWR.t3237 159.452
R1897 VPWR.t3165 VPWR.t2769 159.452
R1898 VPWR.t2120 VPWR.t1395 159.452
R1899 VPWR.t2905 VPWR.t3058 159.452
R1900 VPWR.n5413 VPWR.t2538 158.084
R1901 VPWR.n547 VPWR.t2325 158.06
R1902 VPWR.n3174 VPWR.t831 158.06
R1903 VPWR.n6088 VPWR.t2218 158.06
R1904 VPWR.n6177 VPWR.t819 158.06
R1905 VPWR.n4688 VPWR.t3016 158.06
R1906 VPWR.n3371 VPWR.t942 158.06
R1907 VPWR.t1848 VPWR.t1350 157.774
R1908 VPWR.t2420 VPWR.t3028 157.774
R1909 VPWR.t2159 VPWR.t2428 157.774
R1910 VPWR.t388 VPWR.t1165 157.774
R1911 VPWR.t2414 VPWR.t388 157.774
R1912 VPWR VPWR.t1514 157.774
R1913 VPWR.t2430 VPWR.t1795 157.774
R1914 VPWR.t806 VPWR.t18 157.774
R1915 VPWR.t1901 VPWR.t1339 157.774
R1916 VPWR.t2597 VPWR.t1901 157.774
R1917 VPWR.t2692 VPWR.t199 157.774
R1918 VPWR VPWR.t2399 157.774
R1919 VPWR.n2448 VPWR.t1216 157.145
R1920 VPWR.n1574 VPWR.t1316 156.446
R1921 VPWR.t1441 VPWR.t3273 156.095
R1922 VPWR.t1905 VPWR.t1682 156.095
R1923 VPWR.n3155 VPWR.t829 155.161
R1924 VPWR.n6182 VPWR.t817 155.161
R1925 VPWR.n3055 VPWR.t3208 155.16
R1926 VPWR.n6158 VPWR.t2665 155.16
R1927 VPWR.n1570 VPWR.t1318 155.16
R1928 VPWR.t2925 VPWR.t2819 154.417
R1929 VPWR.n3213 VPWR.t588 154.417
R1930 VPWR.t480 VPWR.t406 154.417
R1931 VPWR.t3220 VPWR.t935 154.417
R1932 VPWR.t1992 VPWR.t2880 154.417
R1933 VPWR.t2673 VPWR.t2079 154.417
R1934 VPWR.t1846 VPWR.t782 154.417
R1935 VPWR.t574 VPWR.t361 154.417
R1936 VPWR.t1787 VPWR.t2420 154.417
R1937 VPWR.t3308 VPWR.t1614 154.417
R1938 VPWR.t907 VPWR.t2808 154.417
R1939 VPWR.t1850 VPWR.t2204 154.417
R1940 VPWR.t3181 VPWR.t2893 154.417
R1941 VPWR.t397 VPWR.t568 154.417
R1942 VPWR.t2426 VPWR.t1783 154.417
R1943 VPWR.t2254 VPWR.t951 154.417
R1944 VPWR.t2238 VPWR.t2177 154.417
R1945 VPWR.n493 VPWR.t905 154.417
R1946 VPWR.t3161 VPWR.t2468 154.417
R1947 VPWR.t2624 VPWR.t1628 154.417
R1948 VPWR.t747 VPWR.t1748 154.417
R1949 VPWR.n4766 VPWR.t515 154.417
R1950 VPWR.t190 VPWR.t21 154.417
R1951 VPWR.t2034 VPWR.t2802 154.417
R1952 VPWR.t2283 VPWR.t1928 154.417
R1953 VPWR.t1922 VPWR.t1337 154.417
R1954 VPWR.t1506 VPWR.t2466 154.417
R1955 VPWR.t2470 VPWR.t1144 154.417
R1956 VPWR.t2531 VPWR.t3223 154.417
R1957 VPWR.t1499 VPWR.t2743 154.417
R1958 VPWR.t2914 VPWR.t1131 154.417
R1959 VPWR.n9047 VPWR.t2423 154.181
R1960 VPWR.n5295 VPWR.t2330 154.118
R1961 VPWR.n2444 VPWR.t1214 153.94
R1962 VPWR.n3413 VPWR.t938 153.726
R1963 VPWR.n4060 VPWR.t1889 153.726
R1964 VPWR.n4088 VPWR.t1955 153.726
R1965 VPWR.n198 VPWR.t2425 153.523
R1966 VPWR.n6186 VPWR.t2663 153.523
R1967 VPWR.n3059 VPWR.t3204 152.879
R1968 VPWR.n2994 VPWR.t1891 152.879
R1969 VPWR.n4089 VPWR.t1959 152.879
R1970 VPWR.n35 VPWR.t2294 152.879
R1971 VPWR.n7638 VPWR.t3072 152.879
R1972 VPWR.n6230 VPWR.t2823 152.879
R1973 VPWR.n8432 VPWR.t2251 152.879
R1974 VPWR.t2202 VPWR 152.739
R1975 VPWR VPWR.t2307 152.739
R1976 VPWR.t838 VPWR.t1695 152.739
R1977 VPWR.t1845 VPWR.t3013 152.739
R1978 VPWR.t2010 VPWR.t1119 152.739
R1979 VPWR.t2351 VPWR 152.739
R1980 VPWR.n6953 VPWR.t2304 151.633
R1981 VPWR.n7033 VPWR.t3244 151.633
R1982 VPWR.n3160 VPWR.t3002 151.633
R1983 VPWR.n73 VPWR.t3246 151.633
R1984 VPWR.n216 VPWR.t2699 151.633
R1985 VPWR.n8874 VPWR.t2481 151.633
R1986 VPWR.n7124 VPWR.t843 151.633
R1987 VPWR.n7147 VPWR.t1269 151.633
R1988 VPWR.n6942 VPWR.t2058 151.633
R1989 VPWR.n7553 VPWR.t1489 151.633
R1990 VPWR.n5785 VPWR.t3240 151.633
R1991 VPWR.n412 VPWR.t2772 151.633
R1992 VPWR.n4454 VPWR.t2908 151.633
R1993 VPWR.n961 VPWR.t919 151.633
R1994 VPWR.n857 VPWR.t2605 151.633
R1995 VPWR.n1850 VPWR.t3279 151.633
R1996 VPWR.n717 VPWR.t761 151.201
R1997 VPWR.t2496 VPWR.t1848 151.06
R1998 VPWR.t3042 VPWR.t139 151.06
R1999 VPWR.t655 VPWR.t2426 151.06
R2000 VPWR.t3075 VPWR.t709 151.06
R2001 VPWR.t24 VPWR.t1292 151.06
R2002 VPWR.n3266 VPWR.t1442 151.016
R2003 VPWR.n36 VPWR.t2296 150.429
R2004 VPWR.n6064 VPWR.t2220 150.429
R2005 VPWR.n6231 VPWR.t2825 150.429
R2006 VPWR.n7665 VPWR.t3070 150.429
R2007 VPWR.n8430 VPWR.t2249 150.429
R2008 VPWR.n4689 VPWR.t3010 150.429
R2009 VPWR.n587 VPWR.t2216 149.696
R2010 VPWR.n861 VPWR.t2173 149.696
R2011 VPWR.n6610 VPWR.t811 149.642
R2012 VPWR.n2694 VPWR.t2760 149.389
R2013 VPWR.t2501 VPWR.t3101 149.382
R2014 VPWR.t921 VPWR.t735 149.382
R2015 VPWR.t1622 VPWR.t1894 149.382
R2016 VPWR.t2236 VPWR.t2763 149.382
R2017 VPWR.t3111 VPWR.t3050 149.382
R2018 VPWR.t2909 VPWR 149.382
R2019 VPWR.n612 VPWR.t3083 149.107
R2020 VPWR.n6537 VPWR.n6536 148.772
R2021 VPWR.n6670 VPWR.t1668 148.364
R2022 VPWR.n2116 VPWR.t3254 148.364
R2023 VPWR.t3304 VPWR.t2957 147.703
R2024 VPWR.t2972 VPWR.t2232 147.703
R2025 VPWR.t3062 VPWR.t2217 147.703
R2026 VPWR.t2674 VPWR.t1817 147.703
R2027 VPWR.t1864 VPWR.t1296 147.703
R2028 VPWR.t1329 VPWR.t3145 147.703
R2029 VPWR.t1443 VPWR.t1643 147.703
R2030 VPWR.t1219 VPWR.t1321 147.703
R2031 VPWR.t1695 VPWR.t3170 147.703
R2032 VPWR.t2721 VPWR.t2032 147.703
R2033 VPWR.t1795 VPWR.t36 147.703
R2034 VPWR.t1207 VPWR.t1391 147.703
R2035 VPWR.t2787 VPWR.t2658 147.703
R2036 VPWR.t2548 VPWR.t2626 147.703
R2037 VPWR.t1405 VPWR.t1512 147.703
R2038 VPWR.t1532 VPWR.t1462 147.703
R2039 VPWR.t2533 VPWR.t1886 147.703
R2040 VPWR.t1759 VPWR.t1313 147.703
R2041 VPWR.t1000 VPWR.t1536 147.703
R2042 VPWR.t2059 VPWR.t2871 147.703
R2043 VPWR.t2903 VPWR.t2692 147.703
R2044 VPWR.t1755 VPWR.t1673 147.703
R2045 VPWR.n4119 VPWR.t3088 147.45
R2046 VPWR.n616 VPWR.t2984 147.45
R2047 VPWR.n5313 VPWR.t2353 147.45
R2048 VPWR.n3079 VPWR.t2392 147.448
R2049 VPWR.n4053 VPWR.t777 147.448
R2050 VPWR.n3214 VPWR.t1718 147.448
R2051 VPWR.n659 VPWR.t2415 147.448
R2052 VPWR.n5124 VPWR.t1714 147.448
R2053 VPWR.n709 VPWR.t2213 146.538
R2054 VPWR.n549 VPWR.t2253 146.538
R2055 VPWR.t2550 VPWR.n5935 146.025
R2056 VPWR.t3113 VPWR.t1175 146.025
R2057 VPWR.t814 VPWR.t1647 146.025
R2058 VPWR.t2440 VPWR.t970 146.025
R2059 VPWR.t2666 VPWR.t2073 146.025
R2060 VPWR.n64 VPWR.t884 145.868
R2061 VPWR.n8870 VPWR.t890 145.868
R2062 VPWR.n1784 VPWR.t2861 145.868
R2063 VPWR.n26 VPWR.t878 145.868
R2064 VPWR.n8109 VPWR.t882 145.868
R2065 VPWR.n8603 VPWR.t1481 145.868
R2066 VPWR.n5804 VPWR.t880 145.868
R2067 VPWR.n1113 VPWR.t2635 145.868
R2068 VPWR.n1947 VPWR.t3299 145.868
R2069 VPWR.n1855 VPWR.t852 145.868
R2070 VPWR.n2008 VPWR.t1243 145.868
R2071 VPWR.n7107 VPWR.t886 145.868
R2072 VPWR.n966 VPWR.t3033 145.81
R2073 VPWR.n536 VPWR.t2643 145.81
R2074 VPWR.n640 VPWR.t1166 145.796
R2075 VPWR.t2731 VPWR.t2737 144.346
R2076 VPWR.t1998 VPWR.t2096 144.346
R2077 VPWR.t1807 VPWR.t1801 144.346
R2078 VPWR.t1801 VPWR.t1803 144.346
R2079 VPWR.t1803 VPWR.t1805 144.346
R2080 VPWR.t1866 VPWR.t1868 144.346
R2081 VPWR.t1868 VPWR.t1870 144.346
R2082 VPWR.t1870 VPWR.t1872 144.346
R2083 VPWR.t2179 VPWR.t2183 144.346
R2084 VPWR.t794 VPWR.t3063 144.346
R2085 VPWR.t1885 VPWR.t2501 144.346
R2086 VPWR.t3024 VPWR.t2899 144.346
R2087 VPWR.t2046 VPWR.t2050 144.346
R2088 VPWR.t3259 VPWR.t943 144.346
R2089 VPWR.t2054 VPWR.t1664 144.346
R2090 VPWR.t3323 VPWR.t3321 144.346
R2091 VPWR.t2486 VPWR.t2809 144.346
R2092 VPWR.t2682 VPWR.t899 144.346
R2093 VPWR.t1932 VPWR.t999 144.346
R2094 VPWR.t1971 VPWR.t1007 144.346
R2095 VPWR.t2709 VPWR.t2715 144.346
R2096 VPWR.t2991 VPWR.t812 144.346
R2097 VPWR.t3095 VPWR.t3097 144.346
R2098 VPWR.t1685 VPWR.t1792 144.346
R2099 VPWR.t2345 VPWR.t2347 144.346
R2100 VPWR.t2347 VPWR.t2341 144.346
R2101 VPWR.t2985 VPWR.t1563 144.346
R2102 VPWR.t735 VPWR.t1636 144.346
R2103 VPWR.t1598 VPWR.t1600 144.346
R2104 VPWR.t1592 VPWR.t1596 144.346
R2105 VPWR.t1596 VPWR.t1577 144.346
R2106 VPWR VPWR.t1583 144.346
R2107 VPWR.t1594 VPWR.t1587 144.346
R2108 VPWR.t1587 VPWR.t1590 144.346
R2109 VPWR.t1566 VPWR.t1037 144.346
R2110 VPWR.t1073 VPWR.t1051 144.346
R2111 VPWR.t1051 VPWR.t1053 144.346
R2112 VPWR.t1095 VPWR.t1097 144.346
R2113 VPWR.t1097 VPWR.t1089 144.346
R2114 VPWR.t1099 VPWR.t1101 144.346
R2115 VPWR.t1107 VPWR.t1111 144.346
R2116 VPWR.t1111 VPWR.t1081 144.346
R2117 VPWR.t2208 VPWR.t2777 144.346
R2118 VPWR.t3160 VPWR.t1045 144.346
R2119 VPWR.t1234 VPWR.t1232 144.346
R2120 VPWR.t1325 VPWR.t1747 144.346
R2121 VPWR.t2136 VPWR.t2146 144.346
R2122 VPWR.t2132 VPWR.t2152 144.346
R2123 VPWR.t2134 VPWR.t2130 144.346
R2124 VPWR.t1067 VPWR.t1059 144.346
R2125 VPWR.t1065 VPWR.t1069 144.346
R2126 VPWR.t1435 VPWR.t1425 144.346
R2127 VPWR.t1411 VPWR.t1407 144.346
R2128 VPWR.t1437 VPWR.t1413 144.346
R2129 VPWR.t1419 VPWR.t1417 144.346
R2130 VPWR.t1427 VPWR.t1423 144.346
R2131 VPWR.t1429 VPWR.t1427 144.346
R2132 VPWR.t2556 VPWR.t2558 144.346
R2133 VPWR.t2558 VPWR.t2560 144.346
R2134 VPWR.t2560 VPWR.t2562 144.346
R2135 VPWR.t2272 VPWR.t2278 144.346
R2136 VPWR.t1897 VPWR.t1526 144.346
R2137 VPWR.t2596 VPWR.t1879 144.346
R2138 VPWR.t1121 VPWR.t1191 144.346
R2139 VPWR.t612 VPWR.t3038 144.346
R2140 VPWR.t1950 VPWR.t2223 144.346
R2141 VPWR.t2022 VPWR.t2028 144.346
R2142 VPWR.t2282 VPWR.t2260 144.346
R2143 VPWR.t1567 VPWR.t1571 144.346
R2144 VPWR.t2434 VPWR.t2444 144.346
R2145 VPWR.t2456 VPWR.t2462 144.346
R2146 VPWR.t2458 VPWR.t2456 144.346
R2147 VPWR.t1071 VPWR.t1079 144.346
R2148 VPWR.t1077 VPWR.t1075 144.346
R2149 VPWR.t1343 VPWR.t1907 144.346
R2150 VPWR.t2195 VPWR.t2189 144.346
R2151 VPWR.t3209 VPWR.t3215 144.346
R2152 VPWR.t1754 VPWR.t1143 144.346
R2153 VPWR.t2399 VPWR.t2741 144.346
R2154 VPWR.t2913 VPWR.t1974 144.346
R2155 VPWR.n6345 VPWR.t2198 143.138
R2156 VPWR.n4731 VPWR.t1678 143.06
R2157 VPWR.t2371 VPWR.t810 142.668
R2158 VPWR.t1604 VPWR 142.668
R2159 VPWR.t1725 VPWR.t2134 142.668
R2160 VPWR.t1431 VPWR.t1942 142.668
R2161 VPWR.t911 VPWR.t867 142.668
R2162 VPWR.t2452 VPWR.t2442 142.668
R2163 VPWR.t2678 VPWR.t2884 142.668
R2164 VPWR.n8734 VPWR.t888 142.571
R2165 VPWR.n456 VPWR.t3049 142.571
R2166 VPWR.n5511 VPWR.t1384 142.571
R2167 VPWR.n1384 VPWR.t807 142.571
R2168 VPWR.n4788 VPWR.t876 142.571
R2169 VPWR.n4693 VPWR.t2863 142.571
R2170 VPWR.n1703 VPWR.t2602 142.571
R2171 VPWR.n5027 VPWR.t1729 142.571
R2172 VPWR.n4406 VPWR.t2583 142.571
R2173 VPWR.n1901 VPWR.t2865 141.75
R2174 VPWR.t1439 VPWR.t1441 140.989
R2175 VPWR.t2818 VPWR.t3271 140.989
R2176 VPWR.t169 VPWR.t1277 140.989
R2177 VPWR.t1020 VPWR.t1274 140.989
R2178 VPWR.t830 VPWR.t828 140.989
R2179 VPWR.t2163 VPWR.t2077 140.989
R2180 VPWR.t2389 VPWR.t2391 140.989
R2181 VPWR.t3071 VPWR.t3069 140.989
R2182 VPWR.t1357 VPWR.t794 140.989
R2183 VPWR.t3060 VPWR.t1835 140.989
R2184 VPWR.t1557 VPWR.t3020 140.989
R2185 VPWR.t1171 VPWR.t1827 140.989
R2186 VPWR.t1630 VPWR.t2747 140.989
R2187 VPWR.t2650 VPWR.t3219 140.989
R2188 VPWR.t3247 VPWR.t3245 140.989
R2189 VPWR.t816 VPWR.t818 140.989
R2190 VPWR.t2662 VPWR.t2664 140.989
R2191 VPWR.t2822 VPWR.t2824 140.989
R2192 VPWR.t1709 VPWR.t2982 140.989
R2193 VPWR.t2879 VPWR.t2804 140.989
R2194 VPWR.t2846 VPWR.t1994 140.989
R2195 VPWR.t2570 VPWR.t166 140.989
R2196 VPWR.t2572 VPWR.t2089 140.989
R2197 VPWR.t1549 VPWR.t2679 140.989
R2198 VPWR.t1551 VPWR.t2498 140.989
R2199 VPWR.t1447 VPWR.t1359 140.989
R2200 VPWR.t2492 VPWR.t2054 140.989
R2201 VPWR.t1665 VPWR.t2102 140.989
R2202 VPWR.t1548 VPWR.t1352 140.989
R2203 VPWR.t2422 VPWR.t2424 140.989
R2204 VPWR.t1964 VPWR.t3117 140.989
R2205 VPWR.t2700 VPWR.t2698 140.989
R2206 VPWR.t2989 VPWR.t3149 140.989
R2207 VPWR.t2995 VPWR.t2989 140.989
R2208 VPWR.t3147 VPWR.t2995 140.989
R2209 VPWR.t891 VPWR.t893 140.989
R2210 VPWR.t1844 VPWR.t3082 140.989
R2211 VPWR.t3079 VPWR.t1914 140.989
R2212 VPWR.t1667 VPWR.t1671 140.989
R2213 VPWR.t1524 VPWR.t1689 140.989
R2214 VPWR.t1669 VPWR.t3309 140.989
R2215 VPWR.t1831 VPWR.t2488 140.989
R2216 VPWR.t999 VPWR.t1177 140.989
R2217 VPWR.t2158 VPWR.t1552 140.989
R2218 VPWR.t1934 VPWR.t2085 140.989
R2219 VPWR.t2789 VPWR.t1971 140.989
R2220 VPWR.t1008 VPWR.t1833 140.989
R2221 VPWR.t1201 VPWR.t1199 140.989
R2222 VPWR.t1199 VPWR.t1701 140.989
R2223 VPWR.t2937 VPWR.t1238 140.989
R2224 VPWR.t2935 VPWR.t1918 140.989
R2225 VPWR.t1544 VPWR.t1546 140.989
R2226 VPWR.t2248 VPWR.t2250 140.989
R2227 VPWR.t1792 VPWR.t1731 140.989
R2228 VPWR.t1797 VPWR.t1553 140.989
R2229 VPWR.t1798 VPWR.t2006 140.989
R2230 VPWR.t2656 VPWR.t2654 140.989
R2231 VPWR.t1561 VPWR.t3084 140.989
R2232 VPWR.t2397 VPWR.t2395 140.989
R2233 VPWR.t2395 VPWR.t1697 140.989
R2234 VPWR.t1936 VPWR.t1979 140.989
R2235 VPWR.t1632 VPWR.t2539 140.989
R2236 VPWR.t790 VPWR.t1837 140.989
R2237 VPWR.t1124 VPWR.t1126 140.989
R2238 VPWR.t2632 VPWR.t2638 140.989
R2239 VPWR.t2630 VPWR.t2634 140.989
R2240 VPWR.t1123 VPWR.t1128 140.989
R2241 VPWR.t1128 VPWR.t3316 140.989
R2242 VPWR.t760 VPWR.t758 140.989
R2243 VPWR.t3267 VPWR.t3269 140.989
R2244 VPWR.t2408 VPWR.t2646 140.989
R2245 VPWR.t990 VPWR.t1270 140.989
R2246 VPWR.t2777 VPWR.t901 140.989
R2247 VPWR.t804 VPWR.t800 140.989
R2248 VPWR.t800 VPWR.t808 140.989
R2249 VPWR.t798 VPWR.t1305 140.989
R2250 VPWR.t2337 VPWR.t2339 140.989
R2251 VPWR.t2911 VPWR.t2828 140.989
R2252 VPWR.t3077 VPWR.t3160 140.989
R2253 VPWR.t1048 VPWR.t463 140.989
R2254 VPWR.t1046 VPWR.t1769 140.989
R2255 VPWR.t2810 VPWR.t2515 140.989
R2256 VPWR.t1315 VPWR.t1317 140.989
R2257 VPWR.t1747 VPWR.t1286 140.989
R2258 VPWR.t1022 VPWR.t1326 140.989
R2259 VPWR.t788 VPWR.t2867 140.989
R2260 VPWR VPWR.t2144 140.989
R2261 VPWR.t2324 VPWR.t2329 140.989
R2262 VPWR.t1612 VPWR.t1610 140.989
R2263 VPWR.t2620 VPWR.t2612 140.989
R2264 VPWR.t1492 VPWR.t2620 140.989
R2265 VPWR.t1490 VPWR.t1492 140.989
R2266 VPWR.t2326 VPWR.t2319 140.989
R2267 VPWR.t3163 VPWR.t3164 140.989
R2268 VPWR.t3009 VPWR.t3015 140.989
R2269 VPWR.t1677 VPWR.t2349 140.989
R2270 VPWR.t972 VPWR.t2366 140.989
R2271 VPWR.t1879 VPWR.t3251 140.989
R2272 VPWR.t1018 VPWR.t2597 140.989
R2273 VPWR.t756 VPWR.t751 140.989
R2274 VPWR.t751 VPWR.t754 140.989
R2275 VPWR.t764 VPWR.t1711 140.989
R2276 VPWR.t1711 VPWR.t1713 140.989
R2277 VPWR.t3011 VPWR.t1510 140.989
R2278 VPWR.t1750 VPWR.t853 140.989
R2279 VPWR.t1749 VPWR.t1750 140.989
R2280 VPWR.t2940 VPWR.t2944 140.989
R2281 VPWR.t1455 VPWR.t1457 140.989
R2282 VPWR.t3290 VPWR.t3296 140.989
R2283 VPWR.t3292 VPWR.t3298 140.989
R2284 VPWR.t2976 VPWR.t1950 140.989
R2285 VPWR.t2225 VPWR.t1763 140.989
R2286 VPWR.t960 VPWR.t2881 140.989
R2287 VPWR.t1026 VPWR.t914 140.989
R2288 VPWR.t3302 VPWR.t2282 140.989
R2289 VPWR.t2261 VPWR.t1024 140.989
R2290 VPWR.t1619 VPWR.t2101 140.989
R2291 VPWR.t1982 VPWR.t1984 140.989
R2292 VPWR.t1984 VPWR.t2576 140.989
R2293 VPWR.t2576 VPWR.t2584 140.989
R2294 VPWR.t2584 VPWR.t2580 140.989
R2295 VPWR.t2574 VPWR.t2578 140.989
R2296 VPWR.t2578 VPWR.t2582 140.989
R2297 VPWR.t859 VPWR.t861 140.989
R2298 VPWR.t1988 VPWR.t3127 140.989
R2299 VPWR.t1240 VPWR.t1246 140.989
R2300 VPWR.t1246 VPWR.t1250 140.989
R2301 VPWR.t1250 VPWR.t1244 140.989
R2302 VPWR.t1244 VPWR.t1248 140.989
R2303 VPWR.t3123 VPWR.t3119 140.989
R2304 VPWR.t2907 VPWR.t2905 140.989
R2305 VPWR.t2961 VPWR.t1507 140.989
R2306 VPWR.t1945 VPWR.t1775 140.989
R2307 VPWR.t125 VPWR.t1751 140.989
R2308 VPWR.t1016 VPWR.t1752 140.989
R2309 VPWR.t2532 VPWR.t1149 140.989
R2310 VPWR.t2951 VPWR.t966 140.989
R2311 VPWR.t2359 VPWR.t1010 140.989
R2312 VPWR.t1014 VPWR.t2400 140.989
R2313 VPWR.t2741 VPWR.t1294 140.989
R2314 VPWR.t2511 VPWR.t2011 140.989
R2315 VPWR.t2696 VPWR.t2913 140.989
R2316 VPWR.t1976 VPWR.t1761 140.989
R2317 VPWR.t2970 VPWR.t2527 140.989
R2318 VPWR.t1256 VPWR.t740 140.989
R2319 VPWR.t2381 VPWR.t1771 140.989
R2320 VPWR.n497 VPWR.t2340 140.417
R2321 VPWR.t3089 VPWR.t1958 139.311
R2322 VPWR.t2113 VPWR.t2480 139.311
R2323 VPWR VPWR.t1280 139.311
R2324 VPWR.t1814 VPWR.t3239 139.311
R2325 VPWR.t1299 VPWR.t2771 139.311
R2326 VPWR.t3017 VPWR.t1063 139.311
R2327 VPWR VPWR.t1433 139.311
R2328 VPWR.t1573 VPWR.t3036 139.311
R2329 VPWR.t264 VPWR.t1071 139.311
R2330 VPWR.n3033 VPWR.t3454 137.977
R2331 VPWR.n6290 VPWR.t3403 137.977
R2332 VPWR.t1978 VPWR 137.633
R2333 VPWR.t2836 VPWR.t1451 137.633
R2334 VPWR VPWR.t1124 137.633
R2335 VPWR.t110 VPWR.t2724 137.633
R2336 VPWR VPWR.t798 137.633
R2337 VPWR.t2535 VPWR.t1303 137.633
R2338 VPWR.t2174 VPWR.t2142 137.633
R2339 VPWR VPWR.t1749 137.633
R2340 VPWR.t2224 VPWR.t2013 137.633
R2341 VPWR VPWR.t1982 137.633
R2342 VPWR.n8571 VPWR.n8567 137.606
R2343 VPWR.n6355 VPWR.n6354 137.606
R2344 VPWR.n5408 VPWR.n5407 137.606
R2345 VPWR.n1901 VPWR.n1900 137.606
R2346 VPWR.t187 VPWR.t2735 135.954
R2347 VPWR VPWR.t2739 135.954
R2348 VPWR VPWR.t1181 135.954
R2349 VPWR VPWR.t840 135.954
R2350 VPWR.t276 VPWR.t2713 135.954
R2351 VPWR.t688 VPWR.t2343 135.954
R2352 VPWR VPWR.t2311 135.954
R2353 VPWR.t2003 VPWR.t1103 135.954
R2354 VPWR.t772 VPWR.t1055 135.954
R2355 VPWR.t1215 VPWR.t2276 135.954
R2356 VPWR.t2864 VPWR.t1497 135.954
R2357 VPWR.n1325 VPWR.n1324 135.371
R2358 VPWR.n6948 VPWR.t3430 134.964
R2359 VPWR.n7043 VPWR.t3429 134.964
R2360 VPWR.n7290 VPWR.t3458 134.964
R2361 VPWR.n4067 VPWR.t3367 134.964
R2362 VPWR.n3237 VPWR.t3414 134.964
R2363 VPWR.n60 VPWR.t3557 134.964
R2364 VPWR.n44 VPWR.t3439 134.964
R2365 VPWR.n40 VPWR.t3569 134.964
R2366 VPWR.n6068 VPWR.t3435 134.964
R2367 VPWR.n8866 VPWR.t3413 134.964
R2368 VPWR.n5939 VPWR.t3451 134.964
R2369 VPWR.n8195 VPWR.t3460 134.964
R2370 VPWR.n8756 VPWR.t3573 134.964
R2371 VPWR.n5869 VPWR.t3575 134.964
R2372 VPWR.n6507 VPWR.t3570 134.964
R2373 VPWR.n6539 VPWR.t3457 134.964
R2374 VPWR.n382 VPWR.t3491 134.964
R2375 VPWR.n724 VPWR.t3390 134.964
R2376 VPWR.n1122 VPWR.t3505 134.964
R2377 VPWR.n750 VPWR.t3496 134.964
R2378 VPWR.n952 VPWR.t3440 134.964
R2379 VPWR.n644 VPWR.t3406 134.964
R2380 VPWR.n5459 VPWR.t3453 134.964
R2381 VPWR.n1383 VPWR.t3529 134.964
R2382 VPWR.n4918 VPWR.t3400 134.964
R2383 VPWR.n2126 VPWR.t3466 134.964
R2384 VPWR.n2188 VPWR.t3402 134.964
R2385 VPWR.n2458 VPWR.t3425 134.964
R2386 VPWR.n2467 VPWR.t3377 134.964
R2387 VPWR.n2474 VPWR.t3577 134.964
R2388 VPWR.n2017 VPWR.t3527 134.964
R2389 VPWR.n2057 VPWR.t3412 134.964
R2390 VPWR.n3501 VPWR.t3553 134.964
R2391 VPWR.n3402 VPWR.t3418 134.964
R2392 VPWR.n3626 VPWR.t3456 134.964
R2393 VPWR.n7073 VPWR.t3551 134.964
R2394 VPWR.n8454 VPWR.n8453 134.528
R2395 VPWR.n8013 VPWR.t2313 134.276
R2396 VPWR.t1938 VPWR.t1515 134.276
R2397 VPWR.t2234 VPWR.t2148 134.276
R2398 VPWR.t3003 VPWR.t795 132.597
R2399 VPWR.t522 VPWR.t1721 132.597
R2400 VPWR VPWR.t2138 132.597
R2401 VPWR.t1031 VPWR.t2327 132.597
R2402 VPWR.t1323 VPWR.t1067 132.597
R2403 VPWR.t1147 VPWR.t1878 132.597
R2404 VPWR.t1339 VPWR.t2106 132.597
R2405 VPWR.t3280 VPWR.t2603 132.597
R2406 VPWR.t2946 VPWR.t2228 132.597
R2407 VPWR.t1145 VPWR.t2024 132.597
R2408 VPWR.t2030 VPWR.t2191 132.597
R2409 VPWR.t2826 VPWR.n3521 132.597
R2410 VPWR.t1105 VPWR.t2875 130.919
R2411 VPWR VPWR.t2838 130.919
R2412 VPWR.t2240 VPWR.t2150 130.919
R2413 VPWR.t1445 VPWR 130.919
R2414 VPWR.n4638 VPWR.t3541 130.833
R2415 VPWR.n1675 VPWR.t3359 130.546
R2416 VPWR.n2694 VPWR.t2332 129.799
R2417 VPWR.n6610 VPWR.t2939 129.708
R2418 VPWR.n1506 VPWR.n1505 129.47
R2419 VPWR VPWR.n6109 129.24
R2420 VPWR.t3021 VPWR.t255 129.24
R2421 VPWR.t1720 VPWR.t205 129.24
R2422 VPWR.t3325 VPWR.t1781 129.24
R2423 VPWR.t1614 VPWR.t193 129.24
R2424 VPWR.t9 VPWR.t907 129.24
R2425 VPWR.t2416 VPWR.t2041 129.24
R2426 VPWR VPWR.n5863 129.24
R2427 VPWR.t637 VPWR 129.24
R2428 VPWR.t893 VPWR.t3081 127.562
R2429 VPWR.t2832 VPWR 127.562
R2430 VPWR.t1937 VPWR.t2397 127.562
R2431 VPWR.t1575 VPWR.t1038 127.562
R2432 VPWR.t1371 VPWR.t3152 127.562
R2433 VPWR.t948 VPWR.t1228 127.562
R2434 VPWR.t154 VPWR 125.883
R2435 VPWR.n3213 VPWR 125.883
R2436 VPWR VPWR.n3879 125.883
R2437 VPWR.t15 VPWR 125.883
R2438 VPWR.n6127 VPWR 125.883
R2439 VPWR VPWR.n6111 125.883
R2440 VPWR VPWR.n58 125.883
R2441 VPWR.t300 VPWR 125.883
R2442 VPWR.n6227 VPWR 125.883
R2443 VPWR.n8012 VPWR 125.883
R2444 VPWR.n9049 VPWR 125.883
R2445 VPWR VPWR.n9048 125.883
R2446 VPWR.t72 VPWR 125.883
R2447 VPWR.n6642 VPWR 125.883
R2448 VPWR.n6658 VPWR 125.883
R2449 VPWR.n8186 VPWR 125.883
R2450 VPWR.t2921 VPWR.t1850 125.883
R2451 VPWR VPWR.n8185 125.883
R2452 VPWR.t86 VPWR 125.883
R2453 VPWR.t3310 VPWR.t1482 125.883
R2454 VPWR.t382 VPWR 125.883
R2455 VPWR VPWR.n1205 125.883
R2456 VPWR VPWR.n1203 125.883
R2457 VPWR.t2362 VPWR.t1107 125.883
R2458 VPWR VPWR.n1202 125.883
R2459 VPWR.t415 VPWR 125.883
R2460 VPWR VPWR.n470 125.883
R2461 VPWR.t202 VPWR 125.883
R2462 VPWR.n559 VPWR 125.883
R2463 VPWR.t2915 VPWR.t2320 125.883
R2464 VPWR.n4766 VPWR 125.883
R2465 VPWR.t539 VPWR 125.883
R2466 VPWR.t2968 VPWR 125.883
R2467 VPWR.n2567 VPWR 125.883
R2468 VPWR.n2568 VPWR 125.883
R2469 VPWR VPWR.n1847 125.883
R2470 VPWR VPWR.n5016 125.883
R2471 VPWR.t327 VPWR 125.883
R2472 VPWR.t976 VPWR 125.883
R2473 VPWR VPWR.n2691 125.883
R2474 VPWR VPWR.n2000 125.883
R2475 VPWR.t80 VPWR 125.883
R2476 VPWR.t931 VPWR 125.883
R2477 VPWR.n4249 VPWR 125.883
R2478 VPWR.n3877 VPWR 124.206
R2479 VPWR.t2343 VPWR 124.206
R2480 VPWR.t1793 VPWR.t3154 124.206
R2481 VPWR.t1373 VPWR.t1093 124.206
R2482 VPWR.t1375 VPWR.t1264 124.206
R2483 VPWR.n1776 VPWR 124.206
R2484 VPWR.n4765 VPWR 124.206
R2485 VPWR.t2562 VPWR 124.206
R2486 VPWR VPWR.t696 124.206
R2487 VPWR.n3521 VPWR 124.206
R2488 VPWR.n8567 VPWR.t1226 123.496
R2489 VPWR.n6354 VPWR.t2994 123.496
R2490 VPWR.n5407 VPWR.t2542 123.496
R2491 VPWR.n1900 VPWR.t1044 123.496
R2492 VPWR.n5429 VPWR.n5428 123.469
R2493 VPWR.t1276 VPWR.t282 122.526
R2494 VPWR.t793 VPWR.t2219 122.526
R2495 VPWR.t945 VPWR.t2846 122.526
R2496 VPWR.t998 VPWR.t2684 122.526
R2497 VPWR.t1691 VPWR.t1656 122.526
R2498 VPWR.t219 VPWR.t1225 122.526
R2499 VPWR.t3282 VPWR.t3284 122.526
R2500 VPWR.t1091 VPWR.t1508 122.526
R2501 VPWR VPWR.t2408 122.526
R2502 VPWR.t2541 VPWR.t2606 122.526
R2503 VPWR.t848 VPWR.t749 122.526
R2504 VPWR.t1193 VPWR.t1040 122.526
R2505 VPWR.t2707 VPWR.t2306 122.526
R2506 VPWR.t796 VPWR.t2100 120.849
R2507 VPWR.t2499 VPWR.t1884 120.849
R2508 VPWR VPWR.t1357 120.849
R2509 VPWR.t1346 VPWR.t3142 120.849
R2510 VPWR.t3026 VPWR.t2900 120.849
R2511 VPWR VPWR.t1464 120.849
R2512 VPWR.t1843 VPWR.t3133 120.849
R2513 VPWR.t2156 VPWR.t3131 120.849
R2514 VPWR.t3275 VPWR.t889 120.849
R2515 VPWR.t2201 VPWR.t2416 120.849
R2516 VPWR.t2094 VPWR.t2197 120.849
R2517 VPWR.t1280 VPWR.t2413 120.849
R2518 VPWR.t3235 VPWR.t3184 120.849
R2519 VPWR.t2214 VPWR.t2410 120.849
R2520 VPWR.t2592 VPWR.t1561 120.849
R2521 VPWR.t2095 VPWR.t2212 120.849
R2522 VPWR.t879 VPWR.t2965 120.849
R2523 VPWR.t2723 VPWR.t1862 120.849
R2524 VPWR.t2644 VPWR.t2412 120.849
R2525 VPWR.t2897 VPWR.t920 120.849
R2526 VPWR.t1190 VPWR.t1383 120.849
R2527 VPWR.t3313 VPWR.t2948 120.849
R2528 VPWR.t1194 VPWR.t3048 120.849
R2529 VPWR VPWR.t3053 120.849
R2530 VPWR.t3053 VPWR.t3167 120.849
R2531 VPWR.t2601 VPWR.t3318 120.849
R2532 VPWR.t2860 VPWR.t773 120.849
R2533 VPWR.t1433 VPWR.t591 120.849
R2534 VPWR.t3162 VPWR.t875 120.849
R2535 VPWR.t846 VPWR.t1905 120.849
R2536 VPWR.t2227 VPWR.t1728 120.849
R2537 VPWR.t2888 VPWR.t2676 120.849
R2538 VPWR.n9048 VPWR.n9047 120.481
R2539 VPWR.n8185 VPWR.n8184 120.481
R2540 VPWR.n8679 VPWR.n8678 120.481
R2541 VPWR.n1202 VPWR.n1201 120.481
R2542 VPWR.n1203 VPWR.n717 120.481
R2543 VPWR.n5018 VPWR.n5017 120.481
R2544 VPWR.n2690 VPWR.n2689 120.481
R2545 VPWR.n4248 VPWR.n4247 120.481
R2546 VPWR.n7280 VPWR.n7046 120.481
R2547 VPWR.n7379 VPWR.n7281 120.481
R2548 VPWR.n7460 VPWR.n6955 120.481
R2549 VPWR.n7513 VPWR.n6943 120.481
R2550 VPWR.n8014 VPWR.n8013 120.481
R2551 VPWR.n6694 VPWR.n6658 120.481
R2552 VPWR.n6449 VPWR.n6448 120.481
R2553 VPWR.n1207 VPWR.n1206 120.481
R2554 VPWR.n2567 VPWR.n2566 120.481
R2555 VPWR.n2691 VPWR.n2009 120.481
R2556 VPWR.n3673 VPWR.n3672 120.481
R2557 VPWR.n7279 VPWR.n7278 120.481
R2558 VPWR.n3279 VPWR.t3272 119.608
R2559 VPWR.n109 VPWR.t2651 119.608
R2560 VPWR.n37 VPWR.t1558 119.608
R2561 VPWR.n6057 VPWR.t1358 119.608
R2562 VPWR.n289 VPWR.t2111 119.608
R2563 VPWR.n8989 VPWR.t2493 119.608
R2564 VPWR.n7905 VPWR.t3258 119.608
R2565 VPWR.n7942 VPWR.t2805 119.608
R2566 VPWR.n8910 VPWR.t2857 119.608
R2567 VPWR.n8124 VPWR.t2790 119.608
R2568 VPWR.n8336 VPWR.t1670 119.608
R2569 VPWR.n5936 VPWR.t2551 119.608
R2570 VPWR.n8202 VPWR.t1178 119.608
R2571 VPWR.n350 VPWR.t2007 119.608
R2572 VPWR.n8673 VPWR.t1732 119.608
R2573 VPWR.n5775 VPWR.t2774 119.608
R2574 VPWR.n1149 VPWR.t1541 119.608
R2575 VPWR.n1005 VPWR.t1967 119.608
R2576 VPWR.n982 VPWR.t1853 119.608
R2577 VPWR.n804 VPWR.t3066 119.608
R2578 VPWR.n444 VPWR.t2890 119.608
R2579 VPWR.n5581 VPWR.t3078 119.608
R2580 VPWR.n1482 VPWR.t902 119.608
R2581 VPWR.n1542 VPWR.t1287 119.608
R2582 VPWR.n4962 VPWR.t2977 119.608
R2583 VPWR.n2175 VPWR.t3252 119.608
R2584 VPWR.n2243 VPWR.t1646 119.608
R2585 VPWR.n2661 VPWR.t3035 119.608
R2586 VPWR.n2303 VPWR.t3303 119.608
R2587 VPWR.n4464 VPWR.t2962 119.608
R2588 VPWR.n2842 VPWR.t1257 119.608
R2589 VPWR.n3533 VPWR.t1138 119.608
R2590 VPWR.n3724 VPWR.t953 119.608
R2591 VPWR.n3515 VPWR.t1150 119.608
R2592 VPWR.n3653 VPWR.t1295 119.608
R2593 VPWR.n4262 VPWR.t2697 119.608
R2594 VPWR.n7759 VPWR.n7758 119.236
R2595 VPWR.n6110 VPWR.t2834 119.171
R2596 VPWR.t6 VPWR.t1365 119.171
R2597 VPWR.t1970 VPWR.t1550 119.171
R2598 VPWR.t2852 VPWR.t60 119.171
R2599 VPWR.t1693 VPWR.t249 119.171
R2600 VPWR VPWR.t947 119.171
R2601 VPWR VPWR.t1680 119.171
R2602 VPWR.t1681 VPWR.t1858 119.171
R2603 VPWR VPWR.t3231 119.171
R2604 VPWR.n5115 VPWR.n1847 119.094
R2605 VPWR.n2695 VPWR.n2694 118.743
R2606 VPWR.n3881 VPWR.n3880 118.513
R2607 VPWR.n4767 VPWR.n4766 117.906
R2608 VPWR.t3271 VPWR 117.492
R2609 VPWR VPWR.t1557 117.492
R2610 VPWR VPWR.t2110 117.492
R2611 VPWR.t2680 VPWR.t1687 117.492
R2612 VPWR VPWR.t2789 117.492
R2613 VPWR VPWR.t2711 117.492
R2614 VPWR.t1731 VPWR 117.492
R2615 VPWR VPWR.t2215 117.492
R2616 VPWR.t474 VPWR.t1604 117.492
R2617 VPWR VPWR.t2889 117.492
R2618 VPWR VPWR.t1612 117.492
R2619 VPWR.t766 VPWR.t646 117.492
R2620 VPWR.t3197 VPWR 117.492
R2621 VPWR.t916 VPWR.t870 117.492
R2622 VPWR.t2580 VPWR.t116 117.492
R2623 VPWR.t3127 VPWR.t1203 117.492
R2624 VPWR.n4661 VPWR.t2231 117.451
R2625 VPWR.n6611 VPWR.n6610 117.132
R2626 VPWR.n3878 VPWR.n2990 116.73
R2627 VPWR.n7809 VPWR.n6111 116.73
R2628 VPWR.n6109 VPWR.n32 116.73
R2629 VPWR.n9144 VPWR.n58 116.73
R2630 VPWR.n6110 VPWR.n6108 116.73
R2631 VPWR.n8012 VPWR.n8011 116.73
R2632 VPWR.n9050 VPWR.n9049 116.73
R2633 VPWR.n6297 VPWR.n6227 116.73
R2634 VPWR.n8187 VPWR.n8186 116.73
R2635 VPWR.n8291 VPWR.n5935 116.73
R2636 VPWR.n6765 VPWR.n6642 116.73
R2637 VPWR.n6447 VPWR.n6446 116.73
R2638 VPWR.n8677 VPWR.n8676 116.73
R2639 VPWR.n8466 VPWR.n5863 116.73
R2640 VPWR.n1205 VPWR.n714 116.73
R2641 VPWR.n1204 VPWR.n716 116.73
R2642 VPWR.n1434 VPWR.n1386 116.73
R2643 VPWR.n470 VPWR.n451 116.73
R2644 VPWR.n5591 VPWR.n471 116.73
R2645 VPWR.n5453 VPWR.n493 116.73
R2646 VPWR.n1776 VPWR.n1775 116.73
R2647 VPWR.n4765 VPWR.n4764 116.73
R2648 VPWR.n5289 VPWR.n1777 116.73
R2649 VPWR.n2569 VPWR.n2568 116.73
R2650 VPWR.n5016 VPWR.n5015 116.73
R2651 VPWR.n4477 VPWR.n2000 116.73
R2652 VPWR.n2693 VPWR.n2692 116.73
R2653 VPWR.n2302 VPWR.n2301 116.73
R2654 VPWR.n3675 VPWR.n3674 116.73
R2655 VPWR.n4250 VPWR.n4249 116.73
R2656 VPWR.n3521 VPWR.n3500 116.73
R2657 VPWR.n3214 VPWR.n3213 116.728
R2658 VPWR.n6128 VPWR.n6127 116.728
R2659 VPWR.n1499 VPWR.n1373 116.728
R2660 VPWR.n1661 VPWR.n559 116.728
R2661 VPWR.n3853 VPWR.t2078 116.322
R2662 VPWR.n6488 VPWR.t2200 116.322
R2663 VPWR.n5401 VPWR.t2178 116.322
R2664 VPWR.n2187 VPWR.t2166 116.322
R2665 VPWR.n2189 VPWR.t1746 116.322
R2666 VPWR.n3496 VPWR.t3194 116.322
R2667 VPWR.t3141 VPWR 115.814
R2668 VPWR.t563 VPWR.t3026 115.814
R2669 VPWR.t2779 VPWR 115.814
R2670 VPWR.t3236 VPWR 115.814
R2671 VPWR.t3227 VPWR.t1655 115.814
R2672 VPWR VPWR.t838 115.814
R2673 VPWR.t1636 VPWR 115.814
R2674 VPWR.t1653 VPWR 115.814
R2675 VPWR.t2599 VPWR.t2128 115.814
R2676 VPWR VPWR.t2610 115.814
R2677 VPWR.t1385 VPWR.t2923 115.814
R2678 VPWR VPWR.t1331 115.814
R2679 VPWR.t3169 VPWR 115.814
R2680 VPWR VPWR.t1737 115.814
R2681 VPWR.t2942 VPWR.t3007 115.814
R2682 VPWR.t1645 VPWR.t857 115.814
R2683 VPWR.t2676 VPWR.t418 115.814
R2684 VPWR.t2402 VPWR 115.814
R2685 VPWR VPWR.t2389 114.135
R2686 VPWR.t778 VPWR 114.135
R2687 VPWR.t1307 VPWR.t3099 114.135
R2688 VPWR VPWR.t2985 114.135
R2689 VPWR.t2387 VPWR 114.135
R2690 VPWR.t744 VPWR.t2405 114.135
R2691 VPWR VPWR.t2324 114.135
R2692 VPWR.t1421 VPWR.t2868 114.135
R2693 VPWR VPWR.t2272 114.135
R2694 VPWR VPWR.t1899 114.135
R2695 VPWR.t851 VPWR.t855 114.135
R2696 VPWR.t3331 VPWR 114.135
R2697 VPWR.t1735 VPWR.t2436 114.135
R2698 VPWR.t828 VPWR 112.457
R2699 VPWR.t1839 VPWR 112.457
R2700 VPWR.t3101 VPWR 112.457
R2701 VPWR.t3245 VPWR 112.457
R2702 VPWR.t2824 VPWR 112.457
R2703 VPWR.t2698 VPWR 112.457
R2704 VPWR.t2753 VPWR.t2161 112.457
R2705 VPWR VPWR.t3249 112.457
R2706 VPWR.n6448 VPWR.t1239 112.457
R2707 VPWR.t1602 VPWR.t923 112.457
R2708 VPWR VPWR.t1581 112.457
R2709 VPWR.t3284 VPWR.t789 112.457
R2710 VPWR VPWR.t3267 112.457
R2711 VPWR VPWR.t2955 112.457
R2712 VPWR.t2116 VPWR 112.457
R2713 VPWR.t1409 VPWR.t1133 112.457
R2714 VPWR.t2169 VPWR 112.457
R2715 VPWR.t3135 VPWR 112.457
R2716 VPWR VPWR.t3290 112.457
R2717 VPWR.t2448 VPWR.t2917 112.457
R2718 VPWR.t2438 VPWR.t2686 112.457
R2719 VPWR.t2765 VPWR 110.778
R2720 VPWR VPWR.t2014 110.778
R2721 VPWR.t1308 VPWR.t883 110.778
R2722 VPWR VPWR.t2286 110.778
R2723 VPWR VPWR.t2371 110.778
R2724 VPWR.t2934 VPWR 110.778
R2725 VPWR.t1966 VPWR.t1726 110.778
R2726 VPWR.t2873 VPWR.t1085 110.778
R2727 VPWR.t1041 VPWR.t3294 110.778
R2728 VPWR.t1136 VPWR.t3292 110.778
R2729 VPWR VPWR.t814 110.778
R2730 VPWR.n5447 VPWR.t2799 110.227
R2731 VPWR VPWR.t1020 109.1
R2732 VPWR.t1468 VPWR 109.1
R2733 VPWR VPWR.t3182 109.1
R2734 VPWR.t2957 VPWR 109.1
R2735 VPWR.t2232 VPWR 109.1
R2736 VPWR.t1817 VPWR 109.1
R2737 VPWR VPWR.t1864 109.1
R2738 VPWR.t2089 VPWR 109.1
R2739 VPWR.t2679 VPWR 109.1
R2740 VPWR.t2498 VPWR 109.1
R2741 VPWR.t2102 VPWR 109.1
R2742 VPWR.t1352 VPWR 109.1
R2743 VPWR.t1916 VPWR 109.1
R2744 VPWR.t498 VPWR.t2486 109.1
R2745 VPWR VPWR.t1831 109.1
R2746 VPWR.t370 VPWR.t1932 109.1
R2747 VPWR.t1833 VPWR 109.1
R2748 VPWR.t1825 VPWR 109.1
R2749 VPWR.t2593 VPWR.t2991 109.1
R2750 VPWR VPWR.t1329 109.1
R2751 VPWR VPWR.t1773 109.1
R2752 VPWR VPWR.t1797 109.1
R2753 VPWR.t2032 VPWR 109.1
R2754 VPWR.t1777 VPWR 109.1
R2755 VPWR.t3052 VPWR 109.1
R2756 VPWR.t1765 VPWR 109.1
R2757 VPWR VPWR.t3172 109.1
R2758 VPWR VPWR.t1207 109.1
R2759 VPWR VPWR.t1912 109.1
R2760 VPWR.t1767 VPWR 109.1
R2761 VPWR.t3306 VPWR.t1234 109.1
R2762 VPWR.t715 VPWR.t1325 109.1
R2763 VPWR VPWR.t1022 109.1
R2764 VPWR.t1512 VPWR 109.1
R2765 VPWR.t2867 VPWR 109.1
R2766 VPWR.t2320 VPWR.n1777 109.1
R2767 VPWR.t3164 VPWR.t243 109.1
R2768 VPWR VPWR.t1675 109.1
R2769 VPWR.t92 VPWR.t2596 109.1
R2770 VPWR VPWR.t869 109.1
R2771 VPWR VPWR.t1679 109.1
R2772 VPWR VPWR.t2008 109.1
R2773 VPWR VPWR.t1986 109.1
R2774 VPWR.t2871 VPWR 109.1
R2775 VPWR.t1763 VPWR 109.1
R2776 VPWR VPWR.t1026 109.1
R2777 VPWR VPWR.t2903 109.1
R2778 VPWR.t2446 VPWR.t3034 109.1
R2779 VPWR.t2688 VPWR.t2458 109.1
R2780 VPWR.t1775 VPWR 109.1
R2781 VPWR.t3176 VPWR 109.1
R2782 VPWR VPWR.t1167 109.1
R2783 VPWR VPWR.t1016 109.1
R2784 VPWR.t1010 VPWR 109.1
R2785 VPWR.t1771 VPWR 109.1
R2786 VPWR.n1314 VPWR.t2788 107.882
R2787 VPWR VPWR.t2731 107.421
R2788 VPWR VPWR.t2315 107.421
R2789 VPWR.t671 VPWR 107.421
R2790 VPWR.t2809 VPWR 107.421
R2791 VPWR VPWR.t2709 107.421
R2792 VPWR VPWR.t1856 107.421
R2793 VPWR.t2369 VPWR.t790 107.421
R2794 VPWR VPWR.t1920 107.421
R2795 VPWR.t2953 VPWR 107.421
R2796 VPWR.t1197 VPWR.t394 107.421
R2797 VPWR.t3318 VPWR 107.421
R2798 VPWR VPWR.t2616 107.421
R2799 VPWR VPWR.t1897 107.421
R2800 VPWR.t1713 VPWR 107.421
R2801 VPWR.t3298 VPWR.t2351 107.421
R2802 VPWR.t1453 VPWR 107.421
R2803 VPWR VPWR.t2588 105.743
R2804 VPWR.t1141 VPWR 105.743
R2805 VPWR VPWR.t89 105.743
R2806 VPWR.t297 VPWR 105.743
R2807 VPWR.t181 VPWR 105.743
R2808 VPWR.t732 VPWR 105.743
R2809 VPWR.t237 VPWR 105.743
R2810 VPWR.t1348 VPWR 105.743
R2811 VPWR.t160 VPWR 105.743
R2812 VPWR.t285 VPWR 105.743
R2813 VPWR VPWR.t2938 105.743
R2814 VPWR.t436 VPWR 105.743
R2815 VPWR.t634 VPWR 105.743
R2816 VPWR.t3091 VPWR.t1478 105.743
R2817 VPWR.t2997 VPWR.t2726 105.743
R2818 VPWR VPWR.t1252 105.743
R2819 VPWR.t677 VPWR 105.743
R2820 VPWR VPWR.t2781 105.743
R2821 VPWR.t2333 VPWR 105.743
R2822 VPWR.t3050 VPWR 105.743
R2823 VPWR.t385 VPWR 105.743
R2824 VPWR VPWR.t2533 105.743
R2825 VPWR VPWR.t460 105.743
R2826 VPWR VPWR.t1730 105.743
R2827 VPWR.t400 VPWR 105.743
R2828 VPWR VPWR.t2949 105.743
R2829 VPWR.t996 VPWR 105.743
R2830 VPWR.t1012 VPWR.t2460 105.743
R2831 VPWR.t101 VPWR 105.743
R2832 VPWR VPWR.t54 105.743
R2833 VPWR.t927 VPWR 105.743
R2834 VPWR.t1341 VPWR.t2564 105.743
R2835 VPWR VPWR.t2403 105.743
R2836 VPWR.t548 VPWR 105.743
R2837 VPWR.t246 VPWR 105.743
R2838 VPWR.n6234 VPWR.n6233 104.809
R2839 VPWR VPWR.t1641 104.064
R2840 VPWR.t1990 VPWR 104.064
R2841 VPWR VPWR.t1447 104.064
R2842 VPWR VPWR.t2568 104.064
R2843 VPWR.t2568 VPWR.t3103 104.064
R2844 VPWR VPWR.t2767 104.064
R2845 VPWR.t1083 VPWR.t1540 104.064
R2846 VPWR.t1188 VPWR.t1105 104.064
R2847 VPWR.t1270 VPWR 104.064
R2848 VPWR VPWR.t1742 104.064
R2849 VPWR.t3199 VPWR 104.064
R2850 VPWR.t2881 VPWR 104.064
R2851 VPWR VPWR.t954 104.064
R2852 VPWR.t2812 VPWR 104.064
R2853 VPWR VPWR.t3178 102.385
R2854 VPWR VPWR.t665 102.385
R2855 VPWR.t1743 VPWR 102.385
R2856 VPWR.t1355 VPWR 102.385
R2857 VPWR.t1185 VPWR 102.385
R2858 VPWR.t240 VPWR 102.385
R2859 VPWR.t1555 VPWR 102.385
R2860 VPWR.t1882 VPWR 102.385
R2861 VPWR.t897 VPWR 102.385
R2862 VPWR VPWR.t1520 102.385
R2863 VPWR.t2791 VPWR 102.385
R2864 VPWR.t560 VPWR 102.385
R2865 VPWR.t1221 VPWR 102.385
R2866 VPWR.t3265 VPWR 102.385
R2867 VPWR.t3093 VPWR.t1480 102.385
R2868 VPWR VPWR.t3107 102.385
R2869 VPWR.t909 VPWR.t2289 102.385
R2870 VPWR VPWR.t1559 102.385
R2871 VPWR VPWR.t2414 102.385
R2872 VPWR.t834 VPWR 102.385
R2873 VPWR VPWR.t1004 102.385
R2874 VPWR VPWR.t806 102.385
R2875 VPWR.t3263 VPWR 102.385
R2876 VPWR.t321 VPWR 102.385
R2877 VPWR.t1460 VPWR 102.385
R2878 VPWR VPWR.t3255 102.385
R2879 VPWR.t2761 VPWR 102.385
R2880 VPWR.t1344 VPWR 102.385
R2881 VPWR.t2016 VPWR 102.385
R2882 VPWR VPWR.t1534 102.385
R2883 VPWR.t1621 VPWR.t986 102.385
R2884 VPWR.t2742 VPWR.n3673 102.385
R2885 VPWR.n4248 VPWR.t741 102.385
R2886 VPWR.n1778 VPWR.t2758 101.465
R2887 VPWR.n1893 VPWR.t1741 101.112
R2888 VPWR.t1717 VPWR 100.707
R2889 VPWR.t776 VPWR 100.707
R2890 VPWR.t3233 VPWR 100.707
R2891 VPWR.t1109 VPWR.t2002 100.707
R2892 VPWR.t1087 VPWR.t2876 100.707
R2893 VPWR VPWR.t2140 100.707
R2894 VPWR VPWR.t2618 100.707
R2895 VPWR VPWR.t1211 100.707
R2896 VPWR.t2949 VPWR.t2034 100.707
R2897 VPWR.t3193 VPWR.t933 100.707
R2898 VPWR.t1888 VPWR 99.0288
R2899 VPWR.t3020 VPWR.t617 99.0288
R2900 VPWR.t3 VPWR.t2879 99.0288
R2901 VPWR.t1177 VPWR.t881 99.0288
R2902 VPWR.t2199 VPWR 99.0288
R2903 VPWR.t3054 VPWR 99.0288
R2904 VPWR.t2768 VPWR.t887 99.0288
R2905 VPWR VPWR.t2118 99.0288
R2906 VPWR.t1600 VPWR 99.0288
R2907 VPWR.t2919 VPWR 99.0288
R2908 VPWR VPWR.t2798 99.0288
R2909 VPWR.t2175 VPWR.t2126 99.0288
R2910 VPWR VPWR.t1057 99.0288
R2911 VPWR.t1217 VPWR.t39 99.0288
R2912 VPWR.t2886 VPWR 99.0288
R2913 VPWR.t1242 VPWR 99.0288
R2914 VPWR.t1507 VPWR.t379 99.0288
R2915 VPWR VPWR.t941 99.0288
R2916 VPWR.t1387 VPWR.t643 99.0288
R2917 VPWR.t740 VPWR.t151 99.0288
R2918 VPWR VPWR.t2181 97.3503
R2919 VPWR.t2727 VPWR.t597 97.3503
R2920 VPWR.t2668 VPWR.t3024 97.3503
R2921 VPWR VPWR.t2048 97.3503
R2922 VPWR.t1723 VPWR.t680 97.3503
R2923 VPWR.t1719 VPWR.t3022 97.3503
R2924 VPWR.t2959 VPWR.t66 97.3503
R2925 VPWR.t2814 VPWR.t409 97.3503
R2926 VPWR.t649 VPWR.t3276 97.3503
R2927 VPWR VPWR.t822 97.3503
R2928 VPWR.t442 VPWR.t2670 97.3503
R2929 VPWR.t1637 VPWR.t3044 97.3503
R2930 VPWR.t1415 VPWR.t1739 97.3503
R2931 VPWR VPWR.t1278 97.3503
R2932 VPWR VPWR.t2026 97.3503
R2933 VPWR VPWR.t3213 97.3503
R2934 VPWR.n3177 VPWR.t797 96.1553
R2935 VPWR.n53 VPWR.t3027 96.1553
R2936 VPWR.n30 VPWR.t1347 96.1553
R2937 VPWR.n6011 VPWR.t2500 96.1553
R2938 VPWR.n8114 VPWR.t2157 96.1553
R2939 VPWR.n8323 VPWR.t2681 96.1553
R2940 VPWR.n6601 VPWR.t1782 96.1553
R2941 VPWR.n8689 VPWR.t1650 96.1553
R2942 VPWR.n8647 VPWR.t3185 96.1553
R2943 VPWR.n6527 VPWR.t2417 96.1553
R2944 VPWR.n599 VPWR.t2411 96.1553
R2945 VPWR.n459 VPWR.t3314 96.1553
R2946 VPWR.n5646 VPWR.t3168 96.1553
R2947 VPWR.n1379 VPWR.t2609 96.1553
R2948 VPWR.n1563 VPWR.t949 96.1553
R2949 VPWR.n4677 VPWR.t2617 96.1553
R2950 VPWR.n5145 VPWR.t2323 96.1553
R2951 VPWR.n2113 VPWR.t847 96.1553
R2952 VPWR.n2247 VPWR.t913 96.1553
R2953 VPWR.n2027 VPWR.t2495 96.1553
R2954 VPWR.n4413 VPWR.t1454 96.1553
R2955 VPWR.n4421 VPWR.t1400 96.1553
R2956 VPWR.n3401 VPWR.t2677 96.1553
R2957 VPWR.t2794 VPWR.t3143 95.6719
R2958 VPWR VPWR.t3207 95.6719
R2959 VPWR.t1309 VPWR 95.6719
R2960 VPWR.t1333 VPWR.t873 95.6719
R2961 VPWR.t1335 VPWR 95.6719
R2962 VPWR.t1960 VPWR 95.6719
R2963 VPWR.t3086 VPWR 95.6719
R2964 VPWR.t820 VPWR 95.6719
R2965 VPWR.t2604 VPWR.t950 95.6719
R2966 VPWR.t2172 VPWR.t3065 95.6719
R2967 VPWR.t1554 VPWR 95.6719
R2968 VPWR.t2625 VPWR.t1811 95.6719
R2969 VPWR.t2660 VPWR.t1415 95.6719
R2970 VPWR VPWR.t1419 95.6719
R2971 VPWR VPWR.t1620 95.6719
R2972 VPWR.t1161 VPWR 95.6719
R2973 VPWR VPWR.t1948 95.6719
R2974 VPWR.t1618 VPWR 95.6719
R2975 VPWR.t994 VPWR.t2434 95.6719
R2976 VPWR.t1137 VPWR.t2565 95.6719
R2977 VPWR.t1498 VPWR.t1028 95.6719
R2978 VPWR VPWR.t1956 94.7045
R2979 VPWR VPWR.t3139 94.7045
R2980 VPWR VPWR.t1307 93.9934
R2981 VPWR.t2571 VPWR 93.9934
R2982 VPWR.t2110 VPWR.t849 93.9934
R2983 VPWR VPWR.t1963 93.9934
R2984 VPWR VPWR.t2115 93.9934
R2985 VPWR.t823 VPWR 93.9934
R2986 VPWR.t1452 VPWR.t3156 93.9934
R2987 VPWR.t172 VPWR.t2136 93.9934
R2988 VPWR.t2866 VPWR 93.9934
R2989 VPWR.t2305 VPWR.t912 93.9934
R2990 VPWR.t1876 VPWR.t2450 93.9934
R2991 VPWR.t2193 VPWR 93.9934
R2992 VPWR VPWR.t780 93.9934
R2993 VPWR.t2167 VPWR.t2061 93.9934
R2994 VPWR.t980 VPWR 93.9934
R2995 VPWR.t2354 VPWR.t2783 93.9934
R2996 VPWR.n3298 VPWR.t1904 93.81
R2997 VPWR.n94 VPWR.t2740 93.81
R2998 VPWR.n9173 VPWR.t3196 93.81
R2999 VPWR.n6059 VPWR.t1881 93.81
R3000 VPWR.n8021 VPWR.t1390 93.81
R3001 VPWR.n243 VPWR.t1182 93.81
R3002 VPWR.n9005 VPWR.t1627 93.81
R3003 VPWR.n7926 VPWR.t2981 93.81
R3004 VPWR.n8897 VPWR.t841 93.81
R3005 VPWR.n8118 VPWR.t1354 93.81
R3006 VPWR.n8319 VPWR.t2703 93.81
R3007 VPWR.n5944 VPWR.t2207 93.81
R3008 VPWR.n8112 VPWR.t1130 93.81
R3009 VPWR.n8777 VPWR.t2019 93.81
R3010 VPWR.n8660 VPWR.t3031 93.81
R3011 VPWR.n5810 VPWR.t1273 93.81
R3012 VPWR.n1169 VPWR.t1189 93.81
R3013 VPWR.n1023 VPWR.t2312 93.81
R3014 VPWR.n996 VPWR.t3283 93.81
R3015 VPWR.n942 VPWR.t924 93.81
R3016 VPWR.n807 VPWR.t1941 93.81
R3017 VPWR.n436 VPWR.t3202 93.81
R3018 VPWR.n468 VPWR.t3287 93.81
R3019 VPWR.n1466 VPWR.t1842 93.81
R3020 VPWR.n1602 VPWR.t1184 93.81
R3021 VPWR.n4946 VPWR.t837 93.81
R3022 VPWR.n1845 VPWR.t1900 93.81
R3023 VPWR.n2159 VPWR.t1154 93.81
R3024 VPWR.n2258 VPWR.t2300 93.81
R3025 VPWR.n2347 VPWR.t1822 93.81
R3026 VPWR.n2090 VPWR.t1736 93.81
R3027 VPWR.n1999 VPWR.t2021 93.81
R3028 VPWR.n2858 VPWR.t926 93.81
R3029 VPWR.n3579 VPWR.t2281 93.81
R3030 VPWR.n3712 VPWR.t3159 93.81
R3031 VPWR.n2790 VPWR.t2817 93.81
R3032 VPWR.n3519 VPWR.t1931 93.81
R3033 VPWR.n3625 VPWR.t3232 93.81
R3034 VPWR.n7989 VPWR.t3519 92.9727
R3035 VPWR.n3062 VPWR.t3357 92.9693
R3036 VPWR.n7636 VPWR.t3347 92.9693
R3037 VPWR.n6156 VPWR.t3530 92.9693
R3038 VPWR.n4093 VPWR.t3579 92.9668
R3039 VPWR.n3065 VPWR.t3525 92.9047
R3040 VPWR.n9201 VPWR.t3438 92.9047
R3041 VPWR.n9133 VPWR.t3512 92.9047
R3042 VPWR.n8966 VPWR.t3374 92.9047
R3043 VPWR.n6159 VPWR.t3431 92.9047
R3044 VPWR.n337 VPWR.t3474 92.9047
R3045 VPWR.n5867 VPWR.t3432 92.9047
R3046 VPWR.n6361 VPWR.t3493 92.9047
R3047 VPWR.n822 VPWR.t3417 92.9047
R3048 VPWR.n495 VPWR.t3514 92.9047
R3049 VPWR.n5003 VPWR.t3538 92.9047
R3050 VPWR.n1902 VPWR.t3475 92.9047
R3051 VPWR.n2296 VPWR.t3334 92.9047
R3052 VPWR.n1995 VPWR.t3373 92.9047
R3053 VPWR.n6666 VPWR.t3534 92.904
R3054 VPWR.n8622 VPWR.t3566 92.904
R3055 VPWR.n813 VPWR.t3583 92.904
R3056 VPWR.n404 VPWR.t3468 92.904
R3057 VPWR.n465 VPWR.t3426 92.904
R3058 VPWR.n1539 VPWR.t3502 92.904
R3059 VPWR.t3018 VPWR.t2295 92.315
R3060 VPWR.t1707 VPWR.t439 92.315
R3061 VPWR.t1006 VPWR 92.315
R3062 VPWR VPWR.t1683 92.315
R3063 VPWR.t1581 VPWR.t1854 92.315
R3064 VPWR.t1407 VPWR.t2614 92.315
R3065 VPWR VPWR.t2595 92.315
R3066 VPWR VPWR.t2494 92.315
R3067 VPWR.t2098 VPWR.t2532 92.315
R3068 VPWR.t2358 VPWR 92.315
R3069 VPWR.t826 VPWR 91.745
R3070 VPWR.t3205 VPWR 91.745
R3071 VPWR VPWR.t1892 91.745
R3072 VPWR VPWR.t2901 91.745
R3073 VPWR.n6704 VPWR.t1708 91.4648
R3074 VPWR.n6646 VPWR.t1704 91.4648
R3075 VPWR.n6358 VPWR.t1702 91.4648
R3076 VPWR.n6347 VPWR.t1692 91.4648
R3077 VPWR.n820 VPWR.t1698 91.4648
R3078 VPWR.n1213 VPWR.t1696 91.4648
R3079 VPWR.n9152 VPWR.t3549 91.34
R3080 VPWR.n209 VPWR.t3423 91.34
R3081 VPWR.n8784 VPWR.t3565 91.34
R3082 VPWR.n870 VPWR.t3479 91.34
R3083 VPWR.n5631 VPWR.t3372 91.34
R3084 VPWR.n551 VPWR.t3511 91.34
R3085 VPWR.n5137 VPWR.t3487 91.34
R3086 VPWR.n4469 VPWR.t3395 91.34
R3087 VPWR.n2822 VPWR.t3558 91.34
R3088 VPWR.n3582 VPWR.t3464 91.34
R3089 VPWR.n9064 VPWR.t3531 91.34
R3090 VPWR.n5927 VPWR.t3421 91.34
R3091 VPWR.n6441 VPWR.t3492 91.34
R3092 VPWR.n1294 VPWR.t3467 91.34
R3093 VPWR.n5013 VPWR.t3396 91.34
R3094 VPWR.n2136 VPWR.t3382 91.34
R3095 VPWR.n3423 VPWR.t3343 91.34
R3096 VPWR.n2934 VPWR.t3532 91.34
R3097 VPWR.n6098 VPWR.t3561 91.2541
R3098 VPWR.n8156 VPWR.t3556 91.2541
R3099 VPWR.n8473 VPWR.t3411 91.2541
R3100 VPWR.n3045 VPWR.t3353 91.2541
R3101 VPWR.n4013 VPWR.t3447 91.2541
R3102 VPWR.n8612 VPWR.t3564 91.2541
R3103 VPWR.n4777 VPWR.t3581 91.2541
R3104 VPWR.n4433 VPWR.t3420 91.2541
R3105 VPWR.n4695 VPWR.t2123 90.683
R3106 VPWR.t2244 VPWR.t3195 90.6365
R3107 VPWR VPWR.t2848 90.6365
R3108 VPWR.t3184 VPWR.t2690 90.6365
R3109 VPWR.t1852 VPWR.t3150 90.6365
R3110 VPWR.t1003 VPWR.t1260 90.6365
R3111 VPWR.t1813 VPWR.t1262 90.6365
R3112 VPWR.t2543 VPWR.t1634 90.6365
R3113 VPWR.t412 VPWR.t3135 90.6365
R3114 VPWR.t483 VPWR.t3011 90.6365
R3115 VPWR.t2063 VPWR.t3288 90.6365
R3116 VPWR.t970 VPWR 90.6365
R3117 VPWR.t2444 VPWR.t2652 90.6365
R3118 VPWR.t2494 VPWR.t51 90.6365
R3119 VPWR VPWR.t2507 90.6365
R3120 VPWR.n4529 VPWR.t3376 89.7
R3121 VPWR.t2899 VPWR.t1363 88.9581
R3122 VPWR VPWR.t2590 88.9581
R3123 VPWR VPWR.t1230 88.9581
R3124 VPWR.t982 VPWR 88.9581
R3125 VPWR.t2152 VPWR.t2352 88.9581
R3126 VPWR VPWR.t958 88.9581
R3127 VPWR.n5472 VPWR.t3448 88.7695
R3128 VPWR.n8440 VPWR.t3379 88.005
R3129 VPWR VPWR.t3327 87.2797
R3130 VPWR.n6658 VPWR.t3079 87.2797
R3131 VPWR.t1126 VPWR.t1034 87.2797
R3132 VPWR.t2628 VPWR.t1779 87.2797
R3133 VPWR.t2773 VPWR.t1258 87.2797
R3134 VPWR.t1799 VPWR.t1272 87.2797
R3135 VPWR.n1386 VPWR.t802 87.2797
R3136 VPWR.t1896 VPWR.t1319 87.2797
R3137 VPWR.t1236 VPWR.t2132 87.2797
R3138 VPWR.t861 VPWR.t525 87.2797
R3139 VPWR.t531 VPWR.t2280 87.2797
R3140 VPWR.n4113 VPWR.t3554 86.9758
R3141 VPWR.n6704 VPWR.t866 86.7743
R3142 VPWR.n5860 VPWR.t1281 86.7743
R3143 VPWR.n6358 VPWR.t3138 86.7743
R3144 VPWR.n6392 VPWR.t1824 86.7743
R3145 VPWR.n820 VPWR.t1170 86.7743
R3146 VPWR.n1409 VPWR.t2898 86.7743
R3147 VPWR.n1305 VPWR.t2659 86.7743
R3148 VPWR.n4678 VPWR.t1386 86.7743
R3149 VPWR.n4678 VPWR.t2237 86.7743
R3150 VPWR.n1938 VPWR.t2064 86.7743
R3151 VPWR.n4010 VPWR.t3335 86.1982
R3152 VPWR.t2181 VPWR.t0 85.6012
R3153 VPWR.t2048 VPWR.t551 85.6012
R3154 VPWR.t1209 VPWR.t2749 85.6012
R3155 VPWR.t3032 VPWR.t1579 85.6012
R3156 VPWR VPWR.t2632 85.6012
R3157 VPWR.t1542 VPWR 85.6012
R3158 VPWR.t3040 VPWR 85.6012
R3159 VPWR.t2124 VPWR.t2642 85.6012
R3160 VPWR.t1571 VPWR.n2690 85.6012
R3161 VPWR.t3125 VPWR.t1459 85.6012
R3162 VPWR.t3213 VPWR.t352 85.6012
R3163 VPWR.t33 VPWR.t952 85.6012
R3164 VPWR.t2638 VPWR 83.9228
R3165 VPWR.t2364 VPWR.t2169 83.9228
R3166 VPWR.t1504 VPWR.t1163 83.9228
R3167 VPWR VPWR.t1135 83.9228
R3168 VPWR.t2704 VPWR.t976 83.9228
R3169 VPWR.t2918 VPWR.t2454 83.9228
R3170 VPWR.t588 VPWR.t1717 82.2443
R3171 VPWR.t2091 VPWR.t3257 82.2443
R3172 VPWR.t881 VPWR.t2830 82.2443
R3173 VPWR.t2893 VPWR 82.2443
R3174 VPWR.t2385 VPWR 82.2443
R3175 VPWR.t2258 VPWR.t1791 82.2443
R3176 VPWR.t918 VPWR.t1585 82.2443
R3177 VPWR.t1837 VPWR.t2840 82.2443
R3178 VPWR.t2083 VPWR 82.2443
R3179 VPWR.n1203 VPWR.t760 82.2443
R3180 VPWR VPWR.t1061 82.2443
R3181 VPWR.t753 VPWR.t1161 82.2443
R3182 VPWR.t2513 VPWR.t1493 82.2443
R3183 VPWR.t2454 VPWR.t2687 82.2443
R3184 VPWR VPWR.t1077 82.2443
R3185 VPWR.t2242 VPWR 80.5659
R3186 VPWR.t2053 VPWR 80.5659
R3187 VPWR.t1914 VPWR 80.5659
R3188 VPWR.t1918 VPWR 80.5659
R3189 VPWR.t1546 VPWR.t231 80.5659
R3190 VPWR.t1649 VPWR.t2745 80.5659
R3191 VPWR.t1910 VPWR 80.5659
R3192 VPWR.t1565 VPWR 80.5659
R3193 VPWR.n1202 VPWR.t2919 80.5659
R3194 VPWR VPWR.t2778 80.5659
R3195 VPWR.t1634 VPWR.t1639 80.5659
R3196 VPWR.t1639 VPWR.t2545 80.5659
R3197 VPWR.t1628 VPWR 80.5659
R3198 VPWR.t3013 VPWR.n4765 80.5659
R3199 VPWR.t3255 VPWR.t580 80.5659
R3200 VPWR.t1493 VPWR.t836 80.5659
R3201 VPWR.t1951 VPWR 80.5659
R3202 VPWR VPWR.t1624 80.5659
R3203 VPWR.t1928 VPWR 80.5659
R3204 VPWR.t2331 VPWR.t279 80.5659
R3205 VPWR.n2691 VPWR.t859 80.5659
R3206 VPWR.t258 VPWR.t2755 78.8874
R3207 VPWR.n1206 VPWR.t3229 78.8874
R3208 VPWR.t2974 VPWR 78.8874
R3209 VPWR.t2407 VPWR 78.8874
R3210 VPWR.t1163 VPWR.t2322 78.8874
R3211 VPWR.t2299 VPWR.t2704 78.8874
R3212 VPWR.t291 VPWR.t974 78.8874
R3213 VPWR.t1149 VPWR.t1621 78.8874
R3214 VPWR.t2519 VPWR.t506 78.8874
R3215 VPWR.n3880 VPWR.t95 77.209
R3216 VPWR.t145 VPWR.n3878 77.209
R3217 VPWR.t347 VPWR.t285 77.209
R3218 VPWR.t391 VPWR.n6447 77.209
R3219 VPWR.n8678 VPWR.t3188 77.209
R3220 VPWR.t1379 VPWR.t1083 77.209
R3221 VPWR.n1373 VPWR.t376 77.209
R3222 VPWR VPWR.t1397 77.209
R3223 VPWR.t1510 VPWR.n1847 77.209
R3224 VPWR.t2432 VPWR 77.209
R3225 VPWR.t288 VPWR.t3123 77.209
R3226 VPWR.t741 VPWR 77.209
R3227 VPWR VPWR.t3319 77.209
R3228 VPWR.n7038 VPWR.n7037 76.0005
R3229 VPWR.n3917 VPWR.n3916 76.0005
R3230 VPWR.n6755 VPWR.n6754 76.0005
R3231 VPWR.n8507 VPWR.n8506 76.0005
R3232 VPWR.n7270 VPWR.n7269 76.0005
R3233 VPWR.t1884 VPWR.t1355 75.5305
R3234 VPWR.t1980 VPWR.t3115 75.5305
R3235 VPWR.t2856 VPWR.t3132 75.5305
R3236 VPWR.t1968 VPWR.t1369 75.5305
R3237 VPWR.t1262 VPWR.t2356 75.5305
R3238 VPWR.t1381 VPWR.t1799 75.5305
R3239 VPWR.t2802 VPWR.t2513 75.5305
R3240 VPWR.t525 VPWR.t1453 75.5305
R3241 VPWR.t992 VPWR.t531 75.5305
R3242 VPWR VPWR.t895 73.8521
R3243 VPWR.n8677 VPWR.t1733 73.8521
R3244 VPWR.n1205 VPWR.t3067 73.8521
R3245 VPWR VPWR.t2083 73.8521
R3246 VPWR.t3316 VPWR.t184 73.8521
R3247 VPWR.t3261 VPWR.t1049 73.8521
R3248 VPWR.t3105 VPWR.t1381 73.8521
R3249 VPWR.t270 VPWR.t1659 73.8521
R3250 VPWR.t3172 VPWR.t270 73.8521
R3251 VPWR.t1657 VPWR 73.8521
R3252 VPWR.t3046 VPWR 73.8521
R3253 VPWR.n1777 VPWR.t2757 73.8521
R3254 VPWR.t1878 VPWR 73.8521
R3255 VPWR.n5017 VPWR.t3329 73.8521
R3256 VPWR VPWR.t2432 73.8521
R3257 VPWR.n2301 VPWR.t3300 73.8521
R3258 VPWR.t1079 VPWR 73.8521
R3259 VPWR.t51 VPWR.t2622 73.8521
R3260 VPWR VPWR.t2484 73.8521
R3261 VPWR.t466 VPWR.t1151 73.8521
R3262 VPWR VPWR.t1499 73.8521
R3263 VPWR.n5427 VPWR.t1638 72.7812
R3264 VPWR.t3115 VPWR.t2244 72.1736
R3265 VPWR.t2690 VPWR.t2258 72.1736
R3266 VPWR.t3315 VPWR.t2209 72.1736
R3267 VPWR.t873 VPWR.t2877 70.4952
R3268 VPWR.t3327 VPWR 70.4952
R3269 VPWR.t1053 VPWR.t3261 70.4952
R3270 VPWR.t2537 VPWR.t2239 70.4952
R3271 VPWR.t2239 VPWR.t2543 70.4952
R3272 VPWR.t1135 VPWR 70.4952
R3273 VPWR VPWR.t2464 70.4952
R3274 VPWR.n2692 VPWR.t2759 70.4952
R3275 VPWR.n1273 VPWR.t3268 69.185
R3276 VPWR.t2161 VPWR.t2856 68.8168
R3277 VPWR.t2418 VPWR.t745 68.8168
R3278 VPWR.n6448 VPWR.t2934 68.8168
R3279 VPWR.t1912 VPWR.t3315 68.8168
R3280 VPWR VPWR.t2120 68.8168
R3281 VPWR.t1899 VPWR.t483 68.8168
R3282 VPWR.n5860 VPWR.t1224 68.0124
R3283 VPWR.n6392 VPWR.t2988 68.0124
R3284 VPWR.n1409 VPWR.t2536 68.0124
R3285 VPWR.n4737 VPWR.t2350 68.0124
R3286 VPWR.n1938 VPWR.t1042 68.0124
R3287 VPWR.n5429 VPWR.n5427 67.1757
R3288 VPWR.t1823 VPWR.t133 67.1383
R3289 VPWR.n8678 VPWR.t3236 67.1383
R3290 VPWR.t157 VPWR.t1940 67.1383
R3291 VPWR.t184 VPWR.t2387 67.1383
R3292 VPWR.t1049 VPWR.t1379 67.1383
R3293 VPWR VPWR.t3040 67.1383
R3294 VPWR.t3201 VPWR.t606 67.1383
R3295 VPWR.n5017 VPWR.t3331 67.1383
R3296 VPWR.n5093 VPWR.n5092 66.8908
R3297 VPWR.n5093 VPWR.n5091 66.8908
R3298 VPWR.n1505 VPWR.t2645 65.9307
R3299 VPWR.n1505 VPWR.t2647 65.9307
R3300 VPWR.n1324 VPWR.t1863 65.8293
R3301 VPWR.n1324 VPWR.t1861 65.8289
R3302 VPWR VPWR.t1173 65.4599
R3303 VPWR.t3149 VPWR 65.4599
R3304 VPWR VPWR.t1962 65.4599
R3305 VPWR.t3132 VPWR.t3180 65.4599
R3306 VPWR.t3249 VPWR.t2201 65.4599
R3307 VPWR.t2590 VPWR 65.4599
R3308 VPWR.t2724 VPWR 65.4599
R3309 VPWR.t857 VPWR.t960 65.4599
R3310 VPWR.t867 VPWR.t2299 65.4599
R3311 VPWR VPWR.t1569 65.4599
R3312 VPWR.n4757 VPWR.n4690 65.3584
R3313 VPWR.n1889 VPWR.n1888 65.3584
R3314 VPWR.n6452 VPWR.t785 64.8416
R3315 VPWR.n1215 VPWR.t839 64.8416
R3316 VPWR.n6453 VPWR.n6452 64.1827
R3317 VPWR.t3143 VPWR.t1439 63.7814
R3318 VPWR VPWR.t962 63.7814
R3319 VPWR.t1377 VPWR 63.7814
R3320 VPWR.t3117 VPWR 63.7814
R3321 VPWR.t1365 VPWR 63.7814
R3322 VPWR VPWR.t2852 63.7814
R3323 VPWR.t2515 VPWR 63.7814
R3324 VPWR.t1248 VPWR.t288 63.7814
R3325 VPWR.n3673 VPWR.t2402 63.7814
R3326 VPWR.t2383 VPWR.n4248 63.7814
R3327 VPWR.n3298 VPWR.t965 63.3219
R3328 VPWR.n3279 VPWR.t963 63.3219
R3329 VPWR.n94 VPWR.t1364 63.3219
R3330 VPWR.n109 VPWR.t2748 63.3219
R3331 VPWR.n9173 VPWR.t3116 63.3219
R3332 VPWR.n37 VPWR.t1378 63.3219
R3333 VPWR.n6057 VPWR.t2835 63.3219
R3334 VPWR.n6059 VPWR.t2851 63.3219
R3335 VPWR.n8021 VPWR.t2843 63.3219
R3336 VPWR.n243 VPWR.t2750 63.3219
R3337 VPWR.n289 VPWR.t3118 63.3219
R3338 VPWR.n8989 VPWR.t1360 63.3219
R3339 VPWR.n9005 VPWR.t1362 63.3219
R3340 VPWR.n7905 VPWR.t2847 63.3219
R3341 VPWR.n7926 VPWR.t1706 63.3219
R3342 VPWR.n7942 VPWR.t1710 63.3219
R3343 VPWR.n8897 VPWR.t1368 63.3219
R3344 VPWR.n8910 VPWR.t2754 63.3219
R3345 VPWR.n8118 VPWR.t2752 63.3219
R3346 VPWR.n8124 VPWR.t1366 63.3219
R3347 VPWR.n8336 VPWR.t1690 63.3219
R3348 VPWR.n8319 VPWR.t1688 63.3219
R3349 VPWR.n5936 VPWR.t2849 63.3219
R3350 VPWR.n5944 VPWR.t2833 63.3219
R3351 VPWR.n8202 VPWR.t2831 63.3219
R3352 VPWR.n8112 VPWR.t2845 63.3219
R3353 VPWR.n6710 VPWR.t894 63.3219
R3354 VPWR.n6710 VPWR.t892 63.3219
R3355 VPWR.n6601 VPWR.t2043 63.3219
R3356 VPWR.n8777 VPWR.t2756 63.3219
R3357 VPWR.n350 VPWR.t2746 63.3219
R3358 VPWR.n8660 VPWR.t2855 63.3219
R3359 VPWR.n8673 VPWR.t2853 63.3219
R3360 VPWR.n6359 VPWR.t1202 63.3219
R3361 VPWR.n6359 VPWR.t1200 63.3219
R3362 VPWR.n5810 VPWR.t1382 63.3219
R3363 VPWR.n5775 VPWR.t1376 63.3219
R3364 VPWR.n1169 VPWR.t1374 63.3219
R3365 VPWR.n1149 VPWR.t1380 63.3219
R3366 VPWR.n819 VPWR.t2398 63.3219
R3367 VPWR.n819 VPWR.t2396 63.3219
R3368 VPWR.n1023 VPWR.t2841 63.3219
R3369 VPWR.n1005 VPWR.t2837 63.3219
R3370 VPWR.n996 VPWR.t1370 63.3219
R3371 VPWR.n982 VPWR.t1372 63.3219
R3372 VPWR.n933 VPWR.t1633 63.3219
R3373 VPWR.n933 VPWR.t2540 63.3219
R3374 VPWR.n807 VPWR.t1700 63.3219
R3375 VPWR.n804 VPWR.t1694 63.3219
R3376 VPWR.n436 VPWR.t2504 63.3219
R3377 VPWR.n444 VPWR.t2516 63.3219
R3378 VPWR.n468 VPWR.t2839 63.3219
R3379 VPWR.n5581 VPWR.t2829 63.3219
R3380 VPWR.n1466 VPWR.t957 63.3219
R3381 VPWR.n1482 VPWR.t991 63.3219
R3382 VPWR.n1314 VPWR.t1921 63.3219
R3383 VPWR.n4731 VPWR.t2615 63.3219
R3384 VPWR.n4737 VPWR.t1943 63.3219
R3385 VPWR.n4692 VPWR.t1396 63.3219
R3386 VPWR.n1542 VPWR.t983 63.3219
R3387 VPWR.n1602 VPWR.t985 63.3219
R3388 VPWR.n4946 VPWR.t2514 63.3219
R3389 VPWR.n4962 VPWR.t2524 63.3219
R3390 VPWR.n1844 VPWR.t1511 63.3219
R3391 VPWR.n1844 VPWR.t3012 63.3219
R3392 VPWR.n2175 VPWR.t973 63.3219
R3393 VPWR.n2159 VPWR.t979 63.3219
R3394 VPWR.n2258 VPWR.t977 63.3219
R3395 VPWR.n2243 VPWR.t961 63.3219
R3396 VPWR.n2661 VPWR.t971 63.3219
R3397 VPWR.n2303 VPWR.t959 63.3219
R3398 VPWR.n2347 VPWR.t975 63.3219
R3399 VPWR.n2090 VPWR.t995 63.3219
R3400 VPWR.n2027 VPWR.t2623 63.3219
R3401 VPWR.n4415 VPWR.t1989 63.3219
R3402 VPWR.n4415 VPWR.t3128 63.3219
R3403 VPWR.n4464 VPWR.t2508 63.3219
R3404 VPWR.n1999 VPWR.t2510 63.3219
R3405 VPWR.n2842 VPWR.t2528 63.3219
R3406 VPWR.n2858 VPWR.t2522 63.3219
R3407 VPWR.n3533 VPWR.t967 63.3219
R3408 VPWR.n3579 VPWR.t993 63.3219
R3409 VPWR.n3712 VPWR.t969 63.3219
R3410 VPWR.n3724 VPWR.t981 63.3219
R3411 VPWR.n2790 VPWR.t2518 63.3219
R3412 VPWR.n3515 VPWR.t987 63.3219
R3413 VPWR.n3519 VPWR.t989 63.3219
R3414 VPWR.n3625 VPWR.t2520 63.3219
R3415 VPWR.n3653 VPWR.t2512 63.3219
R3416 VPWR.n4262 VPWR.t2506 63.3219
R3417 VPWR.n1216 VPWR.n1215 62.7967
R3418 VPWR VPWR.t3062 62.103
R3419 VPWR.t943 VPWR 62.103
R3420 VPWR VPWR.t1006 62.103
R3421 VPWR.t1686 VPWR 62.103
R3422 VPWR VPWR.t823 62.103
R3423 VPWR.t1583 VPWR.t918 62.103
R3424 VPWR VPWR.t1816 62.103
R3425 VPWR.t2322 VPWR.t1157 62.103
R3426 VPWR.t2687 VPWR.t2452 62.103
R3427 VPWR VPWR.t2383 62.103
R3428 VPWR.n6452 VPWR.t3000 60.902
R3429 VPWR.n1215 VPWR.t3171 60.902
R3430 VPWR VPWR.t1276 60.4245
R3431 VPWR.t2834 VPWR 60.4245
R3432 VPWR.t812 VPWR 60.4245
R3433 VPWR VPWR.t1544 60.4245
R3434 VPWR.t2289 VPWR.t1649 60.4245
R3435 VPWR VPWR.t2345 60.4245
R3436 VPWR.t2654 VPWR 60.4245
R3437 VPWR.t2606 VPWR.t2075 60.4245
R3438 VPWR.t2545 VPWR.t1637 60.4245
R3439 VPWR.t1045 VPWR 60.4245
R3440 VPWR.t580 VPWR.t3253 60.4245
R3441 VPWR.t2223 VPWR 60.4245
R3442 VPWR VPWR.t916 60.4245
R3443 VPWR.t2785 VPWR.t3056 60.4245
R3444 VPWR.t2450 VPWR.t2918 60.4245
R3445 VPWR VPWR.t1944 60.4245
R3446 VPWR VPWR.t1754 60.4245
R3447 VPWR.t2783 VPWR.t1341 60.4245
R3448 VPWR.t2361 VPWR 60.4245
R3449 VPWR VPWR.t1975 60.4245
R3450 VPWR.n3879 VPWR.n2998 60.2417
R3451 VPWR.n3877 VPWR.n3876 60.2417
R3452 VPWR.t0 VPWR.t2185 58.7461
R3453 VPWR VPWR.t1309 58.7461
R3454 VPWR.t551 VPWR.t2044 58.7461
R3455 VPWR.t3257 VPWR.t945 58.7461
R3456 VPWR.t2672 VPWR.t2091 58.7461
R3457 VPWR VPWR.t1551 58.7461
R3458 VPWR VPWR.t1335 58.7461
R3459 VPWR.t899 VPWR 58.7461
R3460 VPWR VPWR.t2935 58.7461
R3461 VPWR VPWR.t3086 58.7461
R3462 VPWR.t1683 VPWR 58.7461
R3463 VPWR.t1585 VPWR.t3032 58.7461
R3464 VPWR VPWR.t1046 58.7461
R3465 VPWR.t2642 VPWR.t2154 58.7461
R3466 VPWR.t1157 VPWR.t753 58.7461
R3467 VPWR.t1278 VPWR 58.7461
R3468 VPWR.t1728 VPWR.t2317 58.7461
R3469 VPWR.n2690 VPWR.t1569 58.7461
R3470 VPWR.t3058 VPWR.t1785 58.7461
R3471 VPWR.t352 VPWR.t3211 58.7461
R3472 VPWR.n6732 VPWR.t1467 58.4849
R3473 VPWR.n6343 VPWR.t1289 58.4849
R3474 VPWR.n710 VPWR.t3226 58.4849
R3475 VPWR.n5091 VPWR.t1738 57.7418
R3476 VPWR.n4690 VPWR.t1332 57.7414
R3477 VPWR.n1888 VPWR.t1279 57.7414
R3478 VPWR.n5092 VPWR.t2052 57.7414
R3479 VPWR VPWR.t3247 57.0676
R3480 VPWR VPWR.t2700 57.0676
R3481 VPWR.t2393 VPWR.t498 57.0676
R3482 VPWR.t824 VPWR.t370 57.0676
R3483 VPWR VPWR.t820 57.0676
R3484 VPWR VPWR.t2630 57.0676
R3485 VPWR.t1264 VPWR.t2773 57.0676
R3486 VPWR.t1272 VPWR.t1653 57.0676
R3487 VPWR.t2284 VPWR.t715 57.0676
R3488 VPWR.t2126 VPWR.t1236 57.0676
R3489 VPWR.t1745 VPWR.t2364 57.0676
R3490 VPWR.t2927 VPWR.t92 57.0676
R3491 VPWR.t1530 VPWR.t1504 57.0676
R3492 VPWR VPWR.t1618 57.0676
R3493 VPWR.n5427 VPWR.t3047 57.0216
R3494 VPWR.n4690 VPWR.t1398 56.7568
R3495 VPWR.n1888 VPWR.t2318 56.7568
R3496 VPWR.n5092 VPWR.t2288 56.7568
R3497 VPWR.n5091 VPWR.t1116 56.7564
R3498 VPWR.n7469 VPWR.t827 55.4067
R3499 VPWR.n6944 VPWR.t2821 55.4067
R3500 VPWR.n7557 VPWR.t940 55.4067
R3501 VPWR.n7031 VPWR.t3206 55.4067
R3502 VPWR.n3051 VPWR.t3183 55.4067
R3503 VPWR.n3145 VPWR.t1469 55.4067
R3504 VPWR.n3157 VPWR.t1156 55.4067
R3505 VPWR.n4059 VPWR.t2040 55.4067
R3506 VPWR.n4087 VPWR.t1744 55.4067
R3507 VPWR.n3271 VPWR.t2795 55.4067
R3508 VPWR.n71 VPWR.t1883 55.4067
R3509 VPWR.n213 VPWR.t898 55.4067
R3510 VPWR.n8886 VPWR.t3130 55.4067
R3511 VPWR.n5784 VPWR.t1652 55.4067
R3512 VPWR.n726 VPWR.t2526 55.4067
R3513 VPWR.n410 VPWR.t3166 55.4067
R3514 VPWR.n5104 VPWR.t1987 55.4067
R3515 VPWR.n4458 VPWR.t3059 55.4067
R3516 VPWR.n7114 VPWR.t1893 55.4067
R3517 VPWR.n7190 VPWR.t2902 55.4067
R3518 VPWR.t3273 VPWR 55.3892
R3519 VPWR VPWR.t830 55.3892
R3520 VPWR.t3207 VPWR 55.3892
R3521 VPWR VPWR.t1954 55.3892
R3522 VPWR.t3069 VPWR 55.3892
R3523 VPWR.t451 VPWR.t1630 55.3892
R3524 VPWR.t883 VPWR.t3220 55.3892
R3525 VPWR.t2664 VPWR 55.3892
R3526 VPWR VPWR.t2422 55.3892
R3527 VPWR.t113 VPWR.t1524 55.3892
R3528 VPWR.t3145 VPWR 55.3892
R3529 VPWR VPWR.t2248 55.3892
R3530 VPWR.t887 VPWR.t3221 55.3892
R3531 VPWR.t2726 VPWR.t2592 55.3892
R3532 VPWR.t2636 VPWR 55.3892
R3533 VPWR VPWR.t2430 55.3892
R3534 VPWR VPWR.t2337 55.3892
R3535 VPWR.t1232 VPWR 55.3892
R3536 VPWR.t1317 VPWR 55.3892
R3537 VPWR.t2352 VPWR.t2124 55.3892
R3538 VPWR.t2329 VPWR 55.3892
R3539 VPWR.t1213 VPWR 55.3892
R3540 VPWR VPWR.t1745 55.3892
R3541 VPWR.t1948 VPWR 55.3892
R3542 VPWR VPWR.t871 55.3892
R3543 VPWR.t2759 VPWR 55.3892
R3544 VPWR.t941 VPWR 55.3892
R3545 VPWR.t1143 VPWR.t33 55.3892
R3546 VPWR.n4692 VPWR.t2121 55.1136
R3547 VPWR.t133 VPWR.t1654 53.7107
R3548 VPWR.t2118 VPWR 53.7107
R3549 VPWR.t3152 VPWR.t1852 53.7107
R3550 VPWR.t1034 VPWR.t2628 53.7107
R3551 VPWR.t1779 VPWR.t2636 53.7107
R3552 VPWR VPWR.t2529 53.7107
R3553 VPWR.t1258 VPWR.t1003 53.7107
R3554 VPWR.t1260 VPWR.t1813 53.7107
R3555 VPWR.n1386 VPWR.t804 53.7107
R3556 VPWR VPWR.t770 53.7107
R3557 VPWR.t1211 VPWR 53.7107
R3558 VPWR.t2652 VPWR.t2438 53.7107
R3559 VPWR VPWR.t2335 53.7107
R3560 VPWR VPWR.t1155 52.0323
R3561 VPWR.t1641 VPWR 52.0323
R3562 VPWR VPWR.t1743 52.0323
R3563 VPWR.t3099 VPWR.t2668 52.0323
R3564 VPWR.t2806 VPWR 52.0323
R3565 VPWR.t2042 VPWR 52.0323
R3566 VPWR VPWR.t2552 52.0323
R3567 VPWR VPWR.t1500 52.0323
R3568 VPWR VPWR.t2158 52.0323
R3569 VPWR VPWR.t3190 52.0323
R3570 VPWR VPWR.t3129 52.0323
R3571 VPWR VPWR.t1443 52.0323
R3572 VPWR VPWR.t1221 52.0323
R3573 VPWR.t1559 VPWR 52.0323
R3574 VPWR.t3084 VPWR 52.0323
R3575 VPWR VPWR.t1908 52.0323
R3576 VPWR VPWR.t1632 52.0323
R3577 VPWR.t1854 VPWR.t1594 52.0323
R3578 VPWR VPWR.t1538 52.0323
R3579 VPWR VPWR.t2775 52.0323
R3580 VPWR VPWR.t1651 52.0323
R3581 VPWR VPWR.t2548 52.0323
R3582 VPWR VPWR.t3217 52.0323
R3583 VPWR.t3217 VPWR.t2625 52.0323
R3584 VPWR VPWR.t3165 52.0323
R3585 VPWR VPWR.t1518 52.0323
R3586 VPWR VPWR.t1460 52.0323
R3587 VPWR VPWR.t1532 52.0323
R3588 VPWR.t2612 VPWR 52.0323
R3589 VPWR.t1972 VPWR 52.0323
R3590 VPWR.t2614 VPWR.t1435 52.0323
R3591 VPWR VPWR.t385 52.0323
R3592 VPWR.t1536 VPWR 52.0323
R3593 VPWR VPWR.t3064 52.0323
R3594 VPWR VPWR.t2059 52.0323
R3595 VPWR.t3300 VPWR 52.0323
R3596 VPWR.t2256 VPWR 52.0323
R3597 VPWR.t2622 VPWR 52.0323
R3598 VPWR VPWR.t1988 52.0323
R3599 VPWR VPWR.t1242 52.0323
R3600 VPWR VPWR.t1755 52.0323
R3601 VPWR.t933 VPWR 52.0323
R3602 VPWR.t1906 VPWR 52.0323
R3603 VPWR.t2564 VPWR.t2098 52.0323
R3604 VPWR VPWR.t1014 52.0323
R3605 VPWR VPWR.t1254 52.0323
R3606 VPWR VPWR.t339 52.0323
R3607 VPWR.n2698 VPWR.t1118 51.2205
R3608 VPWR.n7036 VPWR.t3482 50.5057
R3609 VPWR.n3915 VPWR.t3351 50.5057
R3610 VPWR.n6753 VPWR.t3368 50.5057
R3611 VPWR.n8505 VPWR.t3409 50.5057
R3612 VPWR.n7268 VPWR.t3442 50.5057
R3613 VPWR VPWR.t1185 50.3539
R3614 VPWR.t3219 VPWR 50.3539
R3615 VPWR VPWR.t1030 50.3539
R3616 VPWR VPWR.t2672 50.3539
R3617 VPWR VPWR.t1846 50.3539
R3618 VPWR.t3309 VPWR 50.3539
R3619 VPWR.t1819 VPWR.t2717 50.3539
R3620 VPWR.t1721 VPWR 50.3539
R3621 VPWR.t2368 VPWR 50.3539
R3622 VPWR.t3180 VPWR 50.3539
R3623 VPWR VPWR.t3275 50.3539
R3624 VPWR.t3312 VPWR.t219 50.3539
R3625 VPWR VPWR.t3265 50.3539
R3626 VPWR VPWR.t2004 50.3539
R3627 VPWR VPWR.t1227 50.3539
R3628 VPWR.t3150 VPWR.t1452 50.3539
R3629 VPWR.t3156 VPWR.t792 50.3539
R3630 VPWR.t1004 VPWR 50.3539
R3631 VPWR.t920 VPWR 50.3539
R3632 VPWR VPWR.t457 50.3539
R3633 VPWR VPWR.t1190 50.3539
R3634 VPWR VPWR.t1194 50.3539
R3635 VPWR.t2252 VPWR 50.3539
R3636 VPWR.t2138 VPWR.t172 50.3539
R3637 VPWR.t2757 VPWR 50.3539
R3638 VPWR.t773 VPWR 50.3539
R3639 VPWR.t1742 VPWR 50.3539
R3640 VPWR VPWR.t3162 50.3539
R3641 VPWR.t2165 VPWR.t412 50.3539
R3642 VPWR.t1679 VPWR 50.3539
R3643 VPWR VPWR.t1528 50.3539
R3644 VPWR.t1033 VPWR 50.3539
R3645 VPWR.t3294 VPWR.t2063 50.3539
R3646 VPWR VPWR.t2785 50.3539
R3647 VPWR.t2462 VPWR.t1876 50.3539
R3648 VPWR.t1785 VPWR 50.3539
R3649 VPWR VPWR.t2195 50.3539
R3650 VPWR.t2884 VPWR 50.3539
R3651 VPWR VPWR.t2812 50.3539
R3652 VPWR.t665 VPWR 48.6754
R3653 VPWR.t489 VPWR 48.6754
R3654 VPWR.t95 VPWR 48.6754
R3655 VPWR VPWR.t427 48.6754
R3656 VPWR VPWR.t145 48.6754
R3657 VPWR.t75 VPWR 48.6754
R3658 VPWR VPWR.t303 48.6754
R3659 VPWR VPWR.t240 48.6754
R3660 VPWR.t2293 VPWR.t3018 48.6754
R3661 VPWR.t2295 VPWR.t1377 48.6754
R3662 VPWR.t1205 VPWR 48.6754
R3663 VPWR.t571 VPWR 48.6754
R3664 VPWR.t373 VPWR 48.6754
R3665 VPWR.t439 VPWR.t891 48.6754
R3666 VPWR VPWR.t560 48.6754
R3667 VPWR.t706 VPWR 48.6754
R3668 VPWR VPWR.t634 48.6754
R3669 VPWR.t1773 VPWR 48.6754
R3670 VPWR.t1514 VPWR.t2604 48.6754
R3671 VPWR VPWR.t509 48.6754
R3672 VPWR.t603 VPWR 48.6754
R3673 VPWR.t376 VPWR 48.6754
R3674 VPWR.t2209 VPWR.t2608 48.6754
R3675 VPWR.t18 VPWR 48.6754
R3676 VPWR.t1811 VPWR.t1298 48.6754
R3677 VPWR VPWR.t492 48.6754
R3678 VPWR.t1417 VPWR.t2660 48.6754
R3679 VPWR.t1423 VPWR 48.6754
R3680 VPWR.t199 VPWR 48.6754
R3681 VPWR.t2436 VPWR.t994 48.6754
R3682 VPWR VPWR.t101 48.6754
R3683 VPWR.t1028 VPWR.t2361 48.6754
R3684 VPWR VPWR.t548 48.6754
R3685 VPWR.n5448 VPWR.t906 47.7312
R3686 VPWR.t2183 VPWR 46.997
R3687 VPWR.t2246 VPWR.t563 46.997
R3688 VPWR.t2050 VPWR 46.997
R3689 VPWR.t225 VPWR 46.997
R3690 VPWR.t849 VPWR.t1719 46.997
R3691 VPWR.t3022 VPWR.t1333 46.997
R3692 VPWR VPWR.t391 46.997
R3693 VPWR.t3188 VPWR 46.997
R3694 VPWR.t2767 VPWR 46.997
R3695 VPWR.t3229 VPWR 46.997
R3696 VPWR.t1675 VPWR 46.997
R3697 VPWR.t1739 VPWR.t1421 46.997
R3698 VPWR.t1401 VPWR 46.997
R3699 VPWR VPWR.t400 46.997
R3700 VPWR.t2028 VPWR 46.997
R3701 VPWR.t912 VPWR.t1645 46.997
R3702 VPWR.t3215 VPWR 46.997
R3703 VPWR.t418 VPWR.t1789 46.997
R3704 VPWR.t2061 VPWR.t3193 46.997
R3705 VPWR VPWR.t2826 46.997
R3706 VPWR.t2588 VPWR 45.3185
R3707 VPWR.t962 VPWR.t2794 45.3185
R3708 VPWR.t3182 VPWR 45.3185
R3709 VPWR.t3203 VPWR 45.3185
R3710 VPWR VPWR.t2039 45.3185
R3711 VPWR.t617 VPWR.t1174 45.3185
R3712 VPWR VPWR.t2104 45.3185
R3713 VPWR.t944 VPWR.t3 45.3185
R3714 VPWR VPWR.t2087 45.3185
R3715 VPWR.t2938 VPWR 45.3185
R3716 VPWR VPWR.t1916 45.3185
R3717 VPWR VPWR.t2001 45.3185
R3718 VPWR VPWR.t1952 45.3185
R3719 VPWR VPWR.t1829 45.3185
R3720 VPWR.t950 VPWR.t2172 45.3185
R3721 VPWR VPWR.t1592 45.3185
R3722 VPWR VPWR.t3052 45.3185
R3723 VPWR VPWR.t2333 45.3185
R3724 VPWR.t2128 VPWR.t2175 45.3185
R3725 VPWR.t1061 VPWR 45.3185
R3726 VPWR.t869 VPWR 45.3185
R3727 VPWR VPWR.t1159 45.3185
R3728 VPWR.t2008 VPWR 45.3185
R3729 VPWR VPWR.t3121 45.3185
R3730 VPWR VPWR.t2883 45.3185
R3731 VPWR VPWR.t1874 45.3185
R3732 VPWR.t379 VPWR.t1947 45.3185
R3733 VPWR.t1996 VPWR 45.3185
R3734 VPWR.t2565 VPWR.t1498 45.3185
R3735 VPWR.t151 VPWR.t2384 45.3185
R3736 VPWR.n2698 VPWR.t2485 44.3255
R3737 VPWR.n2707 VPWR.t1196 44.3255
R3738 VPWR.n2707 VPWR.t1496 44.3255
R3739 VPWR.t786 VPWR 43.6401
R3740 VPWR.t889 VPWR.t2112 43.6401
R3741 VPWR.t745 VPWR 43.6401
R3742 VPWR VPWR.t1937 43.6401
R3743 VPWR.t2539 VPWR.t1602 43.6401
R3744 VPWR.t1451 VPWR.t1966 43.6401
R3745 VPWR.t2002 VPWR.t1087 43.6401
R3746 VPWR.t2876 VPWR.t1091 43.6401
R3747 VPWR.t2146 VPWR 43.6401
R3748 VPWR.t2122 VPWR 43.6401
R3749 VPWR.n1893 VPWR.t3039 43.5512
R3750 VPWR.n4661 VPWR.t1973 42.3555
R3751 VPWR VPWR.t1890 41.9616
R3752 VPWR VPWR.t2418 41.9616
R3753 VPWR.t1480 VPWR.t3095 41.9616
R3754 VPWR.n1206 VPWR.t1978 41.9616
R3755 VPWR.t2955 VPWR 41.9616
R3756 VPWR.t1331 VPWR 41.9616
R3757 VPWR VPWR.t2931 41.9616
R3758 VPWR.t39 VPWR.t2523 41.9616
R3759 VPWR VPWR.t1240 41.9616
R3760 VPWR.t937 VPWR 41.9616
R3761 VPWR.t643 VPWR.t2505 41.9616
R3762 VPWR.n3218 VPWR.t1275 41.5552
R3763 VPWR.n3218 VPWR.t1021 41.5552
R3764 VPWR.n69 VPWR.t1310 41.5552
R3765 VPWR.n69 VPWR.t2105 41.5552
R3766 VPWR.n49 VPWR.t1172 41.5552
R3767 VPWR.n49 VPWR.t1828 41.5552
R3768 VPWR.n6066 VPWR.t3061 41.5552
R3769 VPWR.n6066 VPWR.t1836 41.5552
R3770 VPWR.n5962 VPWR.t2573 41.5552
R3771 VPWR.n5962 VPWR.t2090 41.5552
R3772 VPWR.n215 VPWR.t1336 41.5552
R3773 VPWR.n215 VPWR.t2088 41.5552
R3774 VPWR.n8976 VPWR.t1666 41.5552
R3775 VPWR.n8976 VPWR.t2103 41.5552
R3776 VPWR.n7907 VPWR.t946 41.5552
R3777 VPWR.n7907 VPWR.t2092 41.5552
R3778 VPWR.n8872 VPWR.t2114 41.5552
R3779 VPWR.n8872 VPWR.t1826 41.5552
R3780 VPWR.n6656 VPWR.t3080 41.5552
R3781 VPWR.n6656 VPWR.t1915 41.5552
R3782 VPWR.n8177 VPWR.t1009 41.5552
R3783 VPWR.n8177 VPWR.t1834 41.5552
R3784 VPWR.n8126 VPWR.t1935 41.5552
R3785 VPWR.n8126 VPWR.t2086 41.5552
R3786 VPWR.n5931 VPWR.t1961 41.5552
R3787 VPWR.n5931 VPWR.t1917 41.5552
R3788 VPWR.n5947 VPWR.t2489 41.5552
R3789 VPWR.n5947 VPWR.t1832 41.5552
R3790 VPWR.n8737 VPWR.t821 41.5552
R3791 VPWR.n8737 VPWR.t1830 41.5552
R3792 VPWR.n8620 VPWR.t1684 41.5552
R3793 VPWR.n8620 VPWR.t1774 41.5552
R3794 VPWR.n6377 VPWR.t2936 41.5552
R3795 VPWR.n6377 VPWR.t1919 41.5552
R3796 VPWR.n5782 VPWR.t1815 41.5552
R3797 VPWR.n5782 VPWR.t1766 41.5552
R3798 VPWR.n720 VPWR.t2874 41.5552
R3799 VPWR.n720 VPWR.t1778 41.5552
R3800 VPWR.n842 VPWR.t1939 41.5552
R3801 VPWR.n842 VPWR.t1911 41.5552
R3802 VPWR.n817 VPWR.t1909 41.5552
R3803 VPWR.n817 VPWR.t1516 41.5552
R3804 VPWR.n1088 VPWR.t1035 41.5552
R3805 VPWR.n1088 VPWR.t1780 41.5552
R3806 VPWR.n1017 VPWR.t791 41.5552
R3807 VPWR.n1017 VPWR.t1838 41.5552
R3808 VPWR.n408 VPWR.t1300 41.5552
R3809 VPWR.n408 VPWR.t1768 41.5552
R3810 VPWR.n463 VPWR.t1047 41.5552
R3811 VPWR.n463 VPWR.t1770 41.5552
R3812 VPWR.n1381 VPWR.t2210 41.5552
R3813 VPWR.n1381 VPWR.t1913 41.5552
R3814 VPWR.n1655 VPWR.t1327 41.5552
R3815 VPWR.n1655 VPWR.t1023 41.5552
R3816 VPWR.n4914 VPWR.t2226 41.5552
R3817 VPWR.n4914 VPWR.t1764 41.5552
R3818 VPWR.n2123 VPWR.t2598 41.5552
R3819 VPWR.n2123 VPWR.t1019 41.5552
R3820 VPWR.n2309 VPWR.t2262 41.5552
R3821 VPWR.n2309 VPWR.t1025 41.5552
R3822 VPWR.n2292 VPWR.t915 41.5552
R3823 VPWR.n2292 VPWR.t1027 41.5552
R3824 VPWR.n2062 VPWR.t2689 41.5552
R3825 VPWR.n2062 VPWR.t1013 41.5552
R3826 VPWR.n4544 VPWR.t1946 41.5552
R3827 VPWR.n4544 VPWR.t1776 41.5552
R3828 VPWR.n4232 VPWR.t2382 41.5552
R3829 VPWR.n4232 VPWR.t1772 41.5552
R3830 VPWR.n3574 VPWR.t2566 41.5552
R3831 VPWR.n3574 VPWR.t1029 41.5552
R3832 VPWR.n3606 VPWR.t2360 41.5552
R3833 VPWR.n3606 VPWR.t1011 41.5552
R3834 VPWR.n3524 VPWR.t1015 41.5552
R3835 VPWR.n3524 VPWR.t2401 41.5552
R3836 VPWR.n3507 VPWR.t1753 41.5552
R3837 VPWR.n3507 VPWR.t1017 41.5552
R3838 VPWR.n2813 VPWR.t1977 41.5552
R3839 VPWR.n2813 VPWR.t1762 41.5552
R3840 VPWR.n6255 VPWR.n6254 41.3997
R3841 VPWR VPWR.t1715 40.2832
R3842 VPWR VPWR.t778 40.2832
R3843 VPWR.t877 VPWR.t1885 40.2832
R3844 VPWR.t1703 VPWR 40.2832
R3845 VPWR.t2745 VPWR.t1798 40.2832
R3846 VPWR.t1540 VPWR.t1109 40.2832
R3847 VPWR.t2610 VPWR 40.2832
R3848 VPWR.t1528 VPWR.t1681 40.2832
R3849 VPWR.n1778 VPWR.t2321 39.8538
R3850 VPWR VPWR.t3141 38.6047
R3851 VPWR.t2830 VPWR.t2368 38.6047
R3852 VPWR.t1656 VPWR.t1290 38.6047
R3853 VPWR VPWR.t2779 38.6047
R3854 VPWR VPWR.t1484 38.6047
R3855 VPWR.t1478 VPWR.t3093 38.6047
R3856 VPWR.t2215 VPWR 38.6047
R3857 VPWR.t1169 VPWR.t594 38.6047
R3858 VPWR.t1093 VPWR.t1188 38.6047
R3859 VPWR.t802 VPWR 38.6047
R3860 VPWR VPWR.t3169 38.6047
R3861 VPWR.t2464 VPWR.t1012 38.6047
R3862 VPWR.t986 VPWR.t1906 38.6047
R3863 VPWR.n4700 VPWR.t2117 38.4155
R3864 VPWR.n4700 VPWR.t1134 38.4155
R3865 VPWR.n7544 VPWR.t2374 37.4305
R3866 VPWR.n7063 VPWR.t2070 37.4305
R3867 VPWR.n7286 VPWR.t2265 37.4305
R3868 VPWR.n3997 VPWR.t1873 37.4305
R3869 VPWR.n3899 VPWR.t1806 37.4305
R3870 VPWR.n3235 VPWR.t2734 37.4305
R3871 VPWR.n7658 VPWR.t2180 37.4305
R3872 VPWR.n6179 VPWR.t2047 37.4305
R3873 VPWR.n6606 VPWR.t3326 37.4305
R3874 VPWR.n8735 VPWR.t2346 37.4305
R3875 VPWR.n8596 VPWR.t3092 37.4305
R3876 VPWR.n6490 VPWR.t2712 37.4305
R3877 VPWR.n5774 VPWR.t1265 37.4305
R3878 VPWR.n5417 VPWR.t2544 37.4305
R3879 VPWR.n4812 VPWR.t2557 37.4305
R3880 VPWR.n1562 VPWR.t1229 37.4305
R3881 VPWR.n1918 VPWR.t1404 37.4305
R3882 VPWR.n1918 VPWR.t2943 37.4305
R3883 VPWR.n1814 VPWR.t1859 37.4305
R3884 VPWR.n2433 VPWR.t2277 37.4305
R3885 VPWR.n2233 VPWR.t2023 37.4305
R3886 VPWR.n2681 VPWR.t1574 37.4305
R3887 VPWR.n4489 VPWR.t2194 37.4305
R3888 VPWR.n3390 VPWR.t3210 37.4305
R3889 VPWR.n7182 VPWR.t1475 37.4305
R3890 VPWR.n7151 VPWR.t2475 37.4305
R3891 VPWR.n7758 VPWR.t3463 36.9896
R3892 VPWR.n6233 VPWR.t3471 36.9896
R3893 VPWR.t2733 VPWR 36.9263
R3894 VPWR.t3103 VPWR.t2753 36.9263
R3895 VPWR.t2711 VPWR 36.9263
R3896 VPWR.t2006 VPWR 36.9263
R3897 VPWR.t2529 VPWR.t1375 36.9263
R3898 VPWR.t2889 VPWR 36.9263
R3899 VPWR VPWR.t3197 36.9263
R3900 VPWR.n6124 VPWR.n6123 36.6122
R3901 VPWR.n5877 VPWR.t1545 36.4455
R3902 VPWR.n602 VPWR.t2655 36.4455
R3903 VPWR.n1891 VPWR.t3332 36.4455
R3904 VPWR.n5118 VPWR.t3198 36.4455
R3905 VPWR.n7294 VPWR.t833 36.1587
R3906 VPWR.n7294 VPWR.t2967 36.1587
R3907 VPWR.n4095 VPWR.t3305 36.1587
R3908 VPWR.n4095 VPWR.t2958 36.1587
R3909 VPWR.n3041 VPWR.t1642 36.1587
R3910 VPWR.n3041 VPWR.t787 36.1587
R3911 VPWR.n3260 VPWR.t3179 36.1587
R3912 VPWR.n3260 VPWR.t2589 36.1587
R3913 VPWR.n9172 VPWR.t1981 36.1587
R3914 VPWR.n9172 VPWR.t2245 36.1587
R3915 VPWR.n6038 VPWR.t2973 36.1587
R3916 VPWR.n6038 VPWR.t2233 36.1587
R3917 VPWR.n7988 VPWR.t1297 36.1587
R3918 VPWR.n7988 VPWR.t1865 36.1587
R3919 VPWR.n6267 VPWR.t2675 36.1587
R3920 VPWR.n6267 VPWR.t1818 36.1587
R3921 VPWR.n6352 VPWR.t1444 36.1587
R3922 VPWR.n6352 VPWR.t1644 36.1587
R3923 VPWR.n8490 VPWR.t1222 36.1587
R3924 VPWR.n8490 VPWR.t1953 36.1587
R3925 VPWR.n8492 VPWR.t1220 36.1587
R3926 VPWR.n8492 VPWR.t1322 36.1587
R3927 VPWR.n6536 VPWR.t3146 36.1587
R3928 VPWR.n6536 VPWR.t1330 36.1587
R3929 VPWR.n723 VPWR.t2722 36.1587
R3930 VPWR.n723 VPWR.t2033 36.1587
R3931 VPWR.n1276 VPWR.t1392 36.1587
R3932 VPWR.n1276 VPWR.t1208 36.1587
R3933 VPWR.n487 VPWR.t2549 36.1587
R3934 VPWR.n487 VPWR.t2627 36.1587
R3935 VPWR.n402 VPWR.t3218 36.1587
R3936 VPWR.n402 VPWR.t1812 36.1587
R3937 VPWR.n460 VPWR.t3264 36.1587
R3938 VPWR.n460 VPWR.t2334 36.1587
R3939 VPWR.n1284 VPWR.t1660 36.1587
R3940 VPWR.n1284 VPWR.t3173 36.1587
R3941 VPWR.n1664 VPWR.t1406 36.1587
R3942 VPWR.n1664 VPWR.t1513 36.1587
R3943 VPWR.n1781 VPWR.t2916 36.1587
R3944 VPWR.n1781 VPWR.t1032 36.1587
R3945 VPWR.n555 VPWR.t1533 36.1587
R3946 VPWR.n555 VPWR.t1463 36.1587
R3947 VPWR.n2425 VPWR.t1537 36.1587
R3948 VPWR.n2425 VPWR.t1001 36.1587
R3949 VPWR.n2428 VPWR.t1314 36.1587
R3950 VPWR.n2428 VPWR.t1760 36.1587
R3951 VPWR.n2429 VPWR.t1887 36.1587
R3952 VPWR.n2429 VPWR.t2534 36.1587
R3953 VPWR.n1961 VPWR.t2060 36.1587
R3954 VPWR.n1961 VPWR.t2872 36.1587
R3955 VPWR.n4487 VPWR.t1756 36.1587
R3956 VPWR.n4487 VPWR.t1674 36.1587
R3957 VPWR.n2298 VPWR.t2693 36.1587
R3958 VPWR.n2298 VPWR.t2904 36.1587
R3959 VPWR.n2225 VPWR.t2310 36.1587
R3960 VPWR.n2225 VPWR.t1146 36.1587
R3961 VPWR.n2315 VPWR.t2017 36.1587
R3962 VPWR.n2315 VPWR.t1875 36.1587
R3963 VPWR.n4494 VPWR.t2031 36.1587
R3964 VPWR.n4494 VPWR.t3177 36.1587
R3965 VPWR.n3389 VPWR.t2074 36.1587
R3966 VPWR.n3389 VPWR.t1168 36.1587
R3967 VPWR.n3740 VPWR.t934 36.1587
R3968 VPWR.n3740 VPWR.t2062 36.1587
R3969 VPWR.n3412 VPWR.t1535 36.1587
R3970 VPWR.n3412 VPWR.t1997 36.1587
R3971 VPWR.n5307 VPWR.t2176 35.4605
R3972 VPWR.t2848 VPWR.n5935 35.2479
R3973 VPWR.t1550 VPWR.t1606 35.2479
R3974 VPWR.t1482 VPWR.t3091 35.2479
R3975 VPWR.t1563 VPWR.t2997 35.2479
R3976 VPWR.t3005 VPWR.t3046 35.2479
R3977 VPWR.t1228 VPWR.t3306 35.2479
R3978 VPWR.t1397 VPWR.t3009 35.2479
R3979 VPWR.t947 VPWR 35.2479
R3980 VPWR.t749 VPWR.t2407 35.2479
R3981 VPWR.t3034 VPWR.t2440 35.2479
R3982 VPWR.t2460 VPWR.t2688 35.2479
R3983 VPWR.t1399 VPWR.t3125 35.2479
R3984 VPWR.n4695 VPWR.t1324 35.1791
R3985 VPWR.n2455 VPWR.n2430 34.6358
R3986 VPWR.n7506 VPWR.n7505 34.6358
R3987 VPWR.n7549 VPWR.n7548 34.6358
R3988 VPWR.n7363 VPWR.n7362 34.6358
R3989 VPWR.n3169 VPWR.n3168 34.6358
R3990 VPWR.n4065 VPWR.n4064 34.6358
R3991 VPWR.n3265 VPWR.n3234 34.6358
R3992 VPWR.n93 VPWR.n63 34.6358
R3993 VPWR.n89 VPWR.n63 34.6358
R3994 VPWR.n9157 VPWR.n9156 34.6358
R3995 VPWR.n8896 VPWR.n8869 34.6358
R3996 VPWR.n8169 VPWR.n8168 34.6358
R3997 VPWR.n8129 VPWR.n8128 34.6358
R3998 VPWR.n8317 VPWR.n8316 34.6358
R3999 VPWR.n6612 VPWR.n6587 34.6358
R4000 VPWR.n8772 VPWR.n8733 34.6358
R4001 VPWR.n8683 VPWR.n352 34.6358
R4002 VPWR.n8497 VPWR.n5861 34.6358
R4003 VPWR.n6534 VPWR.n6484 34.6358
R4004 VPWR.n5827 VPWR.n5826 34.6358
R4005 VPWR.n5435 VPWR.n5432 34.6358
R4006 VPWR.n1434 VPWR.n1387 34.6358
R4007 VPWR.n1450 VPWR.n1449 34.6358
R4008 VPWR.n4756 VPWR.n4691 34.6358
R4009 VPWR.n4752 VPWR.n4691 34.6358
R4010 VPWR.n4764 VPWR.n4647 34.6358
R4011 VPWR.n5290 VPWR.n5289 34.6358
R4012 VPWR.n1916 VPWR.n1915 34.6358
R4013 VPWR.n5089 VPWR.n5088 34.6358
R4014 VPWR.n5088 VPWR.n1851 34.6358
R4015 VPWR.n5155 VPWR.n5154 34.6358
R4016 VPWR.n2573 VPWR.n2572 34.6358
R4017 VPWR.n2260 VPWR.n2257 34.6358
R4018 VPWR.n2323 VPWR.n2322 34.6358
R4019 VPWR.n2368 VPWR.n2302 34.6358
R4020 VPWR.n3736 VPWR.n3498 34.6358
R4021 VPWR.n3537 VPWR.n3536 34.6358
R4022 VPWR.n3676 VPWR.n3675 34.6358
R4023 VPWR.n7113 VPWR.n7048 34.6358
R4024 VPWR.n7173 VPWR.n7172 34.6358
R4025 VPWR.n8048 VPWR.t1847 34.4755
R4026 VPWR.n8052 VPWR.t1849 34.4755
R4027 VPWR.n9032 VPWR.t2421 34.4755
R4028 VPWR.n8178 VPWR.t2429 34.4755
R4029 VPWR.n8137 VPWR.t1851 34.4755
R4030 VPWR.n8625 VPWR.t2427 34.4755
R4031 VPWR.n718 VPWR.t2431 34.4755
R4032 VPWR.n5428 VPWR.t3045 34.4755
R4033 VPWR.n556 VPWR.t2406 34.4755
R4034 VPWR.n1928 VPWR.t2229 34.4755
R4035 VPWR.n4950 VPWR.t2803 34.4755
R4036 VPWR.n2146 VPWR.t1340 34.4755
R4037 VPWR.n2313 VPWR.t1345 34.4755
R4038 VPWR.n2307 VPWR.t1338 34.4755
R4039 VPWR.n3678 VPWR.t1342 34.4755
R4040 VPWR.n7469 VPWR.t2302 34.0906
R4041 VPWR.n6944 VPWR.t2056 34.0906
R4042 VPWR.n7557 VPWR.t1487 34.0906
R4043 VPWR.n7031 VPWR.t3242 34.0906
R4044 VPWR.n3051 VPWR.t2390 34.0906
R4045 VPWR.n3145 VPWR.t1716 34.0906
R4046 VPWR.n3157 VPWR.t3004 34.0906
R4047 VPWR.n4059 VPWR.t779 34.0906
R4048 VPWR.n4087 VPWR.t3090 34.0906
R4049 VPWR.n3271 VPWR.t1440 34.0906
R4050 VPWR.n71 VPWR.t3248 34.0906
R4051 VPWR.n213 VPWR.t2701 34.0906
R4052 VPWR.n8886 VPWR.t2483 34.0906
R4053 VPWR.n5784 VPWR.t3238 34.0906
R4054 VPWR.n726 VPWR.t759 34.0906
R4055 VPWR.n410 VPWR.t2770 34.0906
R4056 VPWR.n5104 VPWR.t3281 34.0906
R4057 VPWR.n4458 VPWR.t2906 34.0906
R4058 VPWR.n7114 VPWR.t845 34.0906
R4059 VPWR.n7190 VPWR.t1267 34.0906
R4060 VPWR.n841 VPWR.n840 33.8829
R4061 VPWR.n4724 VPWR.n4702 33.6462
R4062 VPWR.n5318 VPWR.n5317 33.6462
R4063 VPWR VPWR.t2550 33.5694
R4064 VPWR.t2041 VPWR.t2593 33.5694
R4065 VPWR.t2036 VPWR 33.5694
R4066 VPWR.t1186 VPWR 33.5694
R4067 VPWR.t2634 VPWR.t1123 33.5694
R4068 VPWR.t1081 VPWR.t2873 33.5694
R4069 VPWR.t2075 VPWR 33.5694
R4070 VPWR.t1319 VPWR.t948 33.5694
R4071 VPWR.t1395 VPWR.t2862 33.5694
R4072 VPWR.t1393 VPWR 33.5694
R4073 VPWR.n5428 VPWR.t3006 33.4905
R4074 VPWR.n5417 VPWR.t1640 33.4905
R4075 VPWR.n8304 VPWR.n5934 33.1299
R4076 VPWR.n6646 VPWR.t1465 32.8338
R4077 VPWR.n6347 VPWR.t1291 32.8338
R4078 VPWR.n1213 VPWR.t3228 32.8338
R4079 VPWR.n800 VPWR.n799 32.7534
R4080 VPWR.n5313 VPWR.n5312 32.5491
R4081 VPWR.n5421 VPWR.t1635 32.5055
R4082 VPWR.n5421 VPWR.t2546 32.5055
R4083 VPWR.n8453 VPWR.n8451 32.4088
R4084 VPWR.n8453 VPWR.n8452 32.4084
R4085 VPWR.n5023 VPWR.n5022 32.377
R4086 VPWR.n4937 VPWR.n4936 32.377
R4087 VPWR.n1429 VPWR.n1389 32.0005
R4088 VPWR.n2253 VPWR.n2214 32.0005
R4089 VPWR.t2219 VPWR.t2242 31.891
R4090 VPWR.n8013 VPWR.t2571 31.891
R4091 VPWR.t2684 VPWR.t2921 31.891
R4092 VPWR.t923 VPWR.t1575 31.891
R4093 VPWR.t1579 VPWR 31.891
R4094 VPWR.t792 VPWR 31.891
R4095 VPWR.t243 VPWR.t2326 31.891
R4096 VPWR.t1133 VPWR.t1437 31.891
R4097 VPWR.t1680 VPWR 31.891
R4098 VPWR.t1624 VPWR.t2707 31.891
R4099 VPWR.t2917 VPWR.t2446 31.891
R4100 VPWR.t2686 VPWR.t2448 31.891
R4101 VPWR.n6732 VPWR.t1283 31.6057
R4102 VPWR.n6343 VPWR.t1503 31.6057
R4103 VPWR.n710 VPWR.t930 31.6057
R4104 VPWR.n5286 VPWR.n1779 31.2476
R4105 VPWR.n2450 VPWR.n2449 30.8711
R4106 VPWR.n1436 VPWR.n1435 30.8711
R4107 VPWR.n2577 VPWR.n2576 30.8711
R4108 VPWR.n100 VPWR.t3100 30.5355
R4109 VPWR.n50 VPWR.t3110 30.5355
R4110 VPWR.n9254 VPWR.t3102 30.5355
R4111 VPWR.n8909 VPWR.t3104 30.5355
R4112 VPWR.n5951 VPWR.t3114 30.5355
R4113 VPWR.n353 VPWR.t3108 30.5355
R4114 VPWR.n5809 VPWR.t3106 30.5355
R4115 VPWR.n882 VPWR.t922 30.5355
R4116 VPWR.n4830 VPWR.t3112 30.5355
R4117 VPWR.n1725 VPWR.t1623 30.5355
R4118 VPWR.n5032 VPWR.n5031 30.4946
R4119 VPWR.t2307 VPWR.t315 30.2125
R4120 VPWR.t2212 VPWR.t929 30.2125
R4121 VPWR.t1726 VPWR.t1566 30.2125
R4122 VPWR.t1085 VPWR.t1777 30.2125
R4123 VPWR.t1894 VPWR.t744 30.2125
R4124 VPWR.t2274 VPWR 30.2125
R4125 VPWR.n2568 VPWR.t2909 30.2125
R4126 VPWR.t3296 VPWR.t1041 30.2125
R4127 VPWR.t3288 VPWR.t1136 30.2125
R4128 VPWR.t2442 VPWR.t1735 30.2125
R4129 VPWR.t3223 VPWR.t2951 30.2125
R4130 VPWR.n3690 VPWR.n3516 30.1181
R4131 VPWR.n8290 VPWR.n8289 29.7417
R4132 VPWR.n622 VPWR.n595 29.0829
R4133 VPWR.n8050 VPWR.n8049 28.9887
R4134 VPWR.n8567 VPWR.t1187 28.7575
R4135 VPWR.n6354 VPWR.t2037 28.7575
R4136 VPWR.n5407 VPWR.t2076 28.7575
R4137 VPWR.n1900 VPWR.t1394 28.7575
R4138 VPWR.n8451 VPWR.t2780 28.5655
R4139 VPWR.n9048 VPWR 28.5341
R4140 VPWR.t789 VPWR.t2836 28.5341
R4141 VPWR.t2965 VPWR.t2974 28.5341
R4142 VPWR VPWR.n1776 28.5341
R4143 VPWR.t2130 VPWR.t2599 28.5341
R4144 VPWR.t1610 VPWR.t2860 28.5341
R4145 VPWR.t2923 VPWR.t2230 28.5341
R4146 VPWR.t2868 VPWR.t1409 28.5341
R4147 VPWR VPWR.t2895 28.5341
R4148 VPWR.t1457 VPWR 28.5341
R4149 VPWR.t2013 VPWR.t1951 28.5341
R4150 VPWR VPWR.t931 28.5341
R4151 VPWR.n1845 VPWR.t2009 28.5169
R4152 VPWR.n3853 VPWR.t1180 28.4628
R4153 VPWR.n6488 VPWR.t2706 28.4628
R4154 VPWR.n5401 VPWR.t1523 28.4628
R4155 VPWR.n2187 VPWR.t2896 28.4628
R4156 VPWR.n2189 VPWR.t2969 28.4628
R4157 VPWR.n3496 VPWR.t932 28.4628
R4158 VPWR.n2318 VPWR.n2035 27.8593
R4159 VPWR.n7173 VPWR.n7150 27.8593
R4160 VPWR.n7539 VPWR.t2376 27.5805
R4161 VPWR.n7539 VPWR.t2378 27.5805
R4162 VPWR.n7544 VPWR.t743 27.5805
R4163 VPWR.n7063 VPWR.t2292 27.5805
R4164 VPWR.n7058 VPWR.t2066 27.5805
R4165 VPWR.n7058 VPWR.t2068 27.5805
R4166 VPWR.n7284 VPWR.t2267 27.5805
R4167 VPWR.n7284 VPWR.t2269 27.5805
R4168 VPWR.n7286 VPWR.t2222 27.5805
R4169 VPWR.n3156 VPWR.t1999 27.5805
R4170 VPWR.n3156 VPWR.t2097 27.5805
R4171 VPWR.n3997 VPWR.t2766 27.5805
R4172 VPWR.n3991 VPWR.t1869 27.5805
R4173 VPWR.n3991 VPWR.t1871 27.5805
R4174 VPWR.n3899 VPWR.t1114 27.5805
R4175 VPWR.n3892 VPWR.t1802 27.5805
R4176 VPWR.n3892 VPWR.t1804 27.5805
R4177 VPWR.n3235 VPWR.t3074 27.5805
R4178 VPWR.n3236 VPWR.t2738 27.5805
R4179 VPWR.n3236 VPWR.t2732 27.5805
R4180 VPWR.n100 VPWR.t3025 27.5805
R4181 VPWR.n50 VPWR.t1349 27.5805
R4182 VPWR.n9254 VPWR.t2502 27.5805
R4183 VPWR.n7647 VPWR.t2182 27.5805
R4184 VPWR.n7647 VPWR.t2184 27.5805
R4185 VPWR.n7658 VPWR.t2015 27.5805
R4186 VPWR.n6179 VPWR.t2287 27.5805
R4187 VPWR.n6162 VPWR.t2049 27.5805
R4188 VPWR.n6162 VPWR.t2051 27.5805
R4189 VPWR.n206 VPWR.t850 27.5805
R4190 VPWR.n206 VPWR.t3023 27.5805
R4191 VPWR.n8909 VPWR.t2162 27.5805
R4192 VPWR.n5951 VPWR.t2683 27.5805
R4193 VPWR.n6600 VPWR.t3322 27.5805
R4194 VPWR.n6600 VPWR.t3324 27.5805
R4195 VPWR.n6606 VPWR.t2372 27.5805
R4196 VPWR.n8752 VPWR.t2348 27.5805
R4197 VPWR.n8752 VPWR.t2342 27.5805
R4198 VPWR.n8735 VPWR.t3234 27.5805
R4199 VPWR.n5877 VPWR.t3055 27.5805
R4200 VPWR.n353 VPWR.t3189 27.5805
R4201 VPWR.n8452 VPWR.t2801 27.5805
R4202 VPWR.n8596 VPWR.t3311 27.5805
R4203 VPWR.n8602 VPWR.t3094 27.5805
R4204 VPWR.n8602 VPWR.t3096 27.5805
R4205 VPWR.n6506 VPWR.t2716 27.5805
R4206 VPWR.n6506 VPWR.t2710 27.5805
R4207 VPWR.n6490 VPWR.t746 27.5805
R4208 VPWR.n6522 VPWR.t813 27.5805
R4209 VPWR.n6522 VPWR.t2992 27.5805
R4210 VPWR.n5809 VPWR.t1800 27.5805
R4211 VPWR.n5778 VPWR.t1259 27.5805
R4212 VPWR.n5778 VPWR.t1261 27.5805
R4213 VPWR.n5774 VPWR.t2530 27.5805
R4214 VPWR.n1190 VPWR.t1112 27.5805
R4215 VPWR.n1190 VPWR.t1082 27.5805
R4216 VPWR.n1183 VPWR.t1104 27.5805
R4217 VPWR.n1183 VPWR.t1108 27.5805
R4218 VPWR.n1178 VPWR.t1100 27.5805
R4219 VPWR.n1178 VPWR.t1102 27.5805
R4220 VPWR.n1173 VPWR.t1094 27.5805
R4221 VPWR.n1165 VPWR.t1098 27.5805
R4222 VPWR.n1165 VPWR.t1090 27.5805
R4223 VPWR.n1161 VPWR.t1092 27.5805
R4224 VPWR.n1161 VPWR.t1096 27.5805
R4225 VPWR.n1155 VPWR.t1110 27.5805
R4226 VPWR.n1155 VPWR.t1088 27.5805
R4227 VPWR.n1147 VPWR.t1050 27.5805
R4228 VPWR.n1147 VPWR.t1084 27.5805
R4229 VPWR.n1140 VPWR.t1052 27.5805
R4230 VPWR.n1140 VPWR.t1054 27.5805
R4231 VPWR.n985 VPWR.t3153 27.5805
R4232 VPWR.n985 VPWR.t3151 27.5805
R4233 VPWR.n940 VPWR.t1576 27.5805
R4234 VPWR.n940 VPWR.t1599 27.5805
R4235 VPWR.n978 VPWR.t1591 27.5805
R4236 VPWR.n978 VPWR.t3155 27.5805
R4237 VPWR.n971 VPWR.t1595 27.5805
R4238 VPWR.n971 VPWR.t1588 27.5805
R4239 VPWR.n755 VPWR.t1580 27.5805
R4240 VPWR.n755 VPWR.t1582 27.5805
R4241 VPWR.n757 VPWR.t1584 27.5805
R4242 VPWR.n757 VPWR.t1586 27.5805
R4243 VPWR.n759 VPWR.t1589 27.5805
R4244 VPWR.n948 VPWR.t1597 27.5805
R4245 VPWR.n948 VPWR.t1578 27.5805
R4246 VPWR.n763 VPWR.t1601 27.5805
R4247 VPWR.n763 VPWR.t1593 27.5805
R4248 VPWR.n882 VPWR.t2547 27.5805
R4249 VPWR.n602 VPWR.t2119 27.5805
R4250 VPWR.n592 VPWR.t1564 27.5805
R4251 VPWR.n592 VPWR.t2986 27.5805
R4252 VPWR.n4712 VPWR.t1428 27.5805
R4253 VPWR.n4712 VPWR.t1430 27.5805
R4254 VPWR.n4709 VPWR.t1420 27.5805
R4255 VPWR.n4709 VPWR.t1424 27.5805
R4256 VPWR.n4706 VPWR.t1416 27.5805
R4257 VPWR.n4706 VPWR.t1418 27.5805
R4258 VPWR.n4703 VPWR.t1410 27.5805
R4259 VPWR.n4699 VPWR.t1414 27.5805
R4260 VPWR.n4699 VPWR.t1438 27.5805
R4261 VPWR.n4725 VPWR.t1408 27.5805
R4262 VPWR.n4725 VPWR.t1412 27.5805
R4263 VPWR.n4729 VPWR.t1426 27.5805
R4264 VPWR.n4729 VPWR.t1436 27.5805
R4265 VPWR.n4812 VPWR.t771 27.5805
R4266 VPWR.n4806 VPWR.t2559 27.5805
R4267 VPWR.n4806 VPWR.t2561 27.5805
R4268 VPWR.n4830 VPWR.t3051 27.5805
R4269 VPWR.n1562 VPWR.t1320 27.5805
R4270 VPWR.n1545 VPWR.t1233 27.5805
R4271 VPWR.n1545 VPWR.t1235 27.5805
R4272 VPWR.n4736 VPWR.t1066 27.5805
R4273 VPWR.n4736 VPWR.t1432 27.5805
R4274 VPWR.n4743 VPWR.t1068 27.5805
R4275 VPWR.n4743 VPWR.t1070 27.5805
R4276 VPWR.n544 VPWR.t1056 27.5805
R4277 VPWR.n544 VPWR.t1058 27.5805
R4278 VPWR.n542 VPWR.t2135 27.5805
R4279 VPWR.n542 VPWR.t1064 27.5805
R4280 VPWR.n5303 VPWR.t2129 27.5805
R4281 VPWR.n5303 VPWR.t2131 27.5805
R4282 VPWR.n539 VPWR.t2133 27.5805
R4283 VPWR.n539 VPWR.t2127 27.5805
R4284 VPWR.n537 VPWR.t2125 27.5805
R4285 VPWR.n537 VPWR.t2153 27.5805
R4286 VPWR.n534 VPWR.t2155 27.5805
R4287 VPWR.n529 VPWR.t2137 27.5805
R4288 VPWR.n529 VPWR.t2139 27.5805
R4289 VPWR.n527 VPWR.t2141 27.5805
R4290 VPWR.n527 VPWR.t2147 27.5805
R4291 VPWR.n522 VPWR.t2149 27.5805
R4292 VPWR.n522 VPWR.t2151 27.5805
R4293 VPWR.n1725 VPWR.t1895 27.5805
R4294 VPWR.n1891 VPWR.t3122 27.5805
R4295 VPWR.n5103 VPWR.t1192 27.5805
R4296 VPWR.n5103 VPWR.t1122 27.5805
R4297 VPWR.n5118 VPWR.t2932 27.5805
R4298 VPWR.n2433 VPWR.t1212 27.5805
R4299 VPWR.n2431 VPWR.t2279 27.5805
R4300 VPWR.n2431 VPWR.t2273 27.5805
R4301 VPWR.n2477 VPWR.t1527 27.5805
R4302 VPWR.n2477 VPWR.t1898 27.5805
R4303 VPWR.n2096 VPWR.t2439 27.5805
R4304 VPWR.n2096 VPWR.t2445 27.5805
R4305 VPWR.n2262 VPWR.t2705 27.5805
R4306 VPWR.n2262 VPWR.t868 27.5805
R4307 VPWR.n2233 VPWR.t815 27.5805
R4308 VPWR.n2229 VPWR.t2027 27.5805
R4309 VPWR.n2229 VPWR.t2029 27.5805
R4310 VPWR.n2681 VPWR.t3057 27.5805
R4311 VPWR.n2033 VPWR.t1572 27.5805
R4312 VPWR.n2033 VPWR.t1568 27.5805
R4313 VPWR.n2042 VPWR.t2465 27.5805
R4314 VPWR.n2042 VPWR.t1080 27.5805
R4315 VPWR.n2637 VPWR.t2447 27.5805
R4316 VPWR.n2637 VPWR.t2449 27.5805
R4317 VPWR.n2088 VPWR.t2435 27.5805
R4318 VPWR.n2088 VPWR.t2437 27.5805
R4319 VPWR.n2083 VPWR.t2453 27.5805
R4320 VPWR.n2077 VPWR.t2455 27.5805
R4321 VPWR.n2077 VPWR.t2451 27.5805
R4322 VPWR.n2072 VPWR.t2463 27.5805
R4323 VPWR.n2072 VPWR.t2457 27.5805
R4324 VPWR.n2066 VPWR.t2459 27.5805
R4325 VPWR.n2066 VPWR.t2461 27.5805
R4326 VPWR.n2053 VPWR.t1072 27.5805
R4327 VPWR.n2053 VPWR.t1076 27.5805
R4328 VPWR.n4493 VPWR.t2196 27.5805
R4329 VPWR.n4493 VPWR.t2190 27.5805
R4330 VPWR.n4489 VPWR.t2336 27.5805
R4331 VPWR.n3379 VPWR.t3214 27.5805
R4332 VPWR.n3379 VPWR.t3216 27.5805
R4333 VPWR.n3390 VPWR.t2667 27.5805
R4334 VPWR.n3417 VPWR.t781 27.5805
R4335 VPWR.n3417 VPWR.t2885 27.5805
R4336 VPWR.n7182 VPWR.t1957 27.5805
R4337 VPWR.n7148 VPWR.t1471 27.5805
R4338 VPWR.n7148 VPWR.t1473 27.5805
R4339 VPWR.n7151 VPWR.t3140 27.5805
R4340 VPWR.n7153 VPWR.t2479 27.5805
R4341 VPWR.n7153 VPWR.t2473 27.5805
R4342 VPWR.n6082 VPWR.n6081 27.4829
R4343 VPWR.n8767 VPWR.n8766 27.4829
R4344 VPWR.n7456 VPWR.n7455 27.0566
R4345 VPWR.n6616 VPWR.n6587 27.0566
R4346 VPWR.n5276 VPWR.n5275 27.0566
R4347 VPWR.n2365 VPWR.n2364 27.0566
R4348 VPWR.n4243 VPWR.n2792 27.0566
R4349 VPWR.n2801 VPWR.n2799 27.0566
R4350 VPWR.n942 VPWR.t1039 26.9729
R4351 VPWR.t1363 VPWR 26.8556
R4352 VPWR.t2749 VPWR 26.8556
R4353 VPWR.t1367 VPWR 26.8556
R4354 VPWR.t1577 VPWR.t474 26.8556
R4355 VPWR.t2840 VPWR 26.8556
R4356 VPWR.t1522 VPWR.t2238 26.8556
R4357 VPWR.t2798 VPWR.n493 26.8556
R4358 VPWR VPWR.t1411 26.8556
R4359 VPWR.t853 VPWR.t851 26.8556
R4360 VPWR.t870 VPWR.t2305 26.8556
R4361 VPWR.t917 VPWR.t911 26.8556
R4362 VPWR.n4251 VPWR.n4250 26.7859
R4363 VPWR.n5591 VPWR.n473 26.7859
R4364 VPWR.n7402 VPWR.n7401 26.7859
R4365 VPWR.n6051 VPWR.n6050 26.7859
R4366 VPWR.n8045 VPWR.n8044 26.7859
R4367 VPWR.n7922 VPWR.n7921 26.7859
R4368 VPWR.n8257 VPWR.n8256 26.7859
R4369 VPWR.n2153 VPWR.n2152 26.7859
R4370 VPWR.n1570 VPWR.n1569 26.7299
R4371 VPWR.n8048 VPWR.t1991 26.5955
R4372 VPWR.n8052 VPWR.t783 26.5955
R4373 VPWR.n9032 VPWR.t1788 26.5955
R4374 VPWR.n8178 VPWR.t2933 26.5955
R4375 VPWR.n8137 VPWR.t2205 26.5955
R4376 VPWR.n6620 VPWR.t2990 26.5955
R4377 VPWR.n6620 VPWR.t2996 26.5955
R4378 VPWR.n8625 VPWR.t1784 26.5955
R4379 VPWR.n8594 VPWR.t3266 26.5955
R4380 VPWR.n8594 VPWR.t1485 26.5955
R4381 VPWR.n8597 VPWR.t1483 26.5955
R4382 VPWR.n8597 VPWR.t1479 26.5955
R4383 VPWR.n718 VPWR.t2920 26.5955
R4384 VPWR.n1173 VPWR.t1106 26.5955
R4385 VPWR.n730 VPWR.t3317 26.5955
R4386 VPWR.n730 VPWR.t2388 26.5955
R4387 VPWR.n732 VPWR.t2639 26.5955
R4388 VPWR.n732 VPWR.t2631 26.5955
R4389 VPWR.n1039 VPWR.t2637 26.5955
R4390 VPWR.n1039 VPWR.t2633 26.5955
R4391 VPWR.n1086 VPWR.t1127 26.5955
R4392 VPWR.n1086 VPWR.t2629 26.5955
R4393 VPWR.n759 VPWR.t1605 26.5955
R4394 VPWR.n594 VPWR.t1560 26.5955
R4395 VPWR.n628 VPWR.t1562 26.5955
R4396 VPWR.n5433 VPWR.t3041 26.5955
R4397 VPWR.n5433 VPWR.t2338 26.5955
R4398 VPWR.n1427 VPWR.t799 26.5955
R4399 VPWR.n1427 VPWR.t1306 26.5955
R4400 VPWR.n1388 VPWR.t801 26.5955
R4401 VPWR.n1388 VPWR.t809 26.5955
R4402 VPWR.n1385 VPWR.t803 26.5955
R4403 VPWR.n1385 VPWR.t805 26.5955
R4404 VPWR.n4703 VPWR.t1422 26.5955
R4405 VPWR.n1786 VPWR.t2613 26.5955
R4406 VPWR.n1786 VPWR.t2621 26.5955
R4407 VPWR.n1780 VPWR.t2328 26.5955
R4408 VPWR.n1780 VPWR.t2619 26.5955
R4409 VPWR.n5307 VPWR.t1237 26.5955
R4410 VPWR.n534 VPWR.t2145 26.5955
R4411 VPWR.n525 VPWR.t2235 26.5955
R4412 VPWR.n525 VPWR.t2241 26.5955
R4413 VPWR.n556 VPWR.t1461 26.5955
R4414 VPWR.n1942 VPWR.t3289 26.5955
R4415 VPWR.n1942 VPWR.t3293 26.5955
R4416 VPWR.n1934 VPWR.t3297 26.5955
R4417 VPWR.n1934 VPWR.t3295 26.5955
R4418 VPWR.n1910 VPWR.t1458 26.5955
R4419 VPWR.n1910 VPWR.t3291 26.5955
R4420 VPWR.n1928 VPWR.t2930 26.5955
R4421 VPWR.n1923 VPWR.t2947 26.5955
R4422 VPWR.n1923 VPWR.t2941 26.5955
R4423 VPWR.n1852 VPWR.t856 26.5955
R4424 VPWR.n1852 VPWR.t854 26.5955
R4425 VPWR.n4950 VPWR.t2035 26.5955
R4426 VPWR.n5132 VPWR.t765 26.5955
R4427 VPWR.n5132 VPWR.t1712 26.5955
R4428 VPWR.n1831 VPWR.t1158 26.5955
R4429 VPWR.n1831 VPWR.t1162 26.5955
R4430 VPWR.n5149 VPWR.t1531 26.5955
R4431 VPWR.n5149 VPWR.t1164 26.5955
R4432 VPWR.n1829 VPWR.t755 26.5955
R4433 VPWR.n1829 VPWR.t750 26.5955
R4434 VPWR.n1816 VPWR.t757 26.5955
R4435 VPWR.n1816 VPWR.t752 26.5955
R4436 VPWR.n1814 VPWR.t1529 26.5955
R4437 VPWR.n2146 VPWR.t1148 26.5955
R4438 VPWR.n4400 VPWR.t2575 26.5955
R4439 VPWR.n4400 VPWR.t2579 26.5955
R4440 VPWR.n4377 VPWR.t2585 26.5955
R4441 VPWR.n4377 VPWR.t2581 26.5955
R4442 VPWR.n4360 VPWR.t1985 26.5955
R4443 VPWR.n4360 VPWR.t2577 26.5955
R4444 VPWR.n2313 VPWR.t1927 26.5955
R4445 VPWR.n2307 VPWR.t1923 26.5955
R4446 VPWR.n2083 VPWR.t2443 26.5955
R4447 VPWR.n4440 VPWR.t1249 26.5955
R4448 VPWR.n4440 VPWR.t3124 26.5955
R4449 VPWR.n4430 VPWR.t1251 26.5955
R4450 VPWR.n4430 VPWR.t1245 26.5955
R4451 VPWR.n2007 VPWR.t1241 26.5955
R4452 VPWR.n2007 VPWR.t1247 26.5955
R4453 VPWR.n3678 VPWR.t2355 26.5955
R4454 VPWR.n8608 VPWR.n355 26.3534
R4455 VPWR.n4688 VPWR.n4648 25.977
R4456 VPWR.n3177 VPWR.t2587 25.6105
R4457 VPWR.n53 VPWR.t2247 25.6105
R4458 VPWR.n30 VPWR.t1609 25.6105
R4459 VPWR.n6011 VPWR.t2203 25.6105
R4460 VPWR.n8114 VPWR.t2555 25.6105
R4461 VPWR.n8323 VPWR.t2718 25.6105
R4462 VPWR.n8689 VPWR.t910 25.6105
R4463 VPWR.n8647 VPWR.t2259 25.6105
R4464 VPWR.n6527 VPWR.t2594 25.6105
R4465 VPWR.n599 VPWR.t2308 25.6105
R4466 VPWR.n459 VPWR.t2793 25.6105
R4467 VPWR.n5646 VPWR.t1198 25.6105
R4468 VPWR.n1379 VPWR.t864 25.6105
R4469 VPWR.n1563 VPWR.t3307 25.6105
R4470 VPWR.n4677 VPWR.t2764 25.6105
R4471 VPWR.n5145 VPWR.t1505 25.6105
R4472 VPWR.n2113 VPWR.t2910 25.6105
R4473 VPWR.n2247 VPWR.t858 25.6105
R4474 VPWR.n4413 VPWR.t862 25.6105
R4475 VPWR.n4421 VPWR.t1204 25.6105
R4476 VPWR.n3401 VPWR.t1790 25.6105
R4477 VPWR.n1558 VPWR.n1557 25.6005
R4478 VPWR.n2450 VPWR.n2448 25.6005
R4479 VPWR.n3072 VPWR.n3055 25.224
R4480 VPWR.n3174 VPWR.n3154 25.224
R4481 VPWR.n1571 VPWR.n1570 25.224
R4482 VPWR.n2444 VPWR.n2432 25.224
R4483 VPWR.n3411 VPWR.n3371 25.224
R4484 VPWR.n7184 VPWR.n7183 25.224
R4485 VPWR.n7172 VPWR.n7152 25.224
R4486 VPWR.n8188 VPWR.n8187 25.1912
R4487 VPWR.n1032 VPWR.n754 25.1912
R4488 VPWR.n5453 VPWR.n5446 25.1912
R4489 VPWR.n4956 VPWR.n4955 25.1912
R4490 VPWR.n4477 VPWR.n2005 25.1912
R4491 VPWR.n7505 VPWR.n6950 25.1912
R4492 VPWR.n7564 VPWR.n7563 25.1912
R4493 VPWR.n7362 VPWR.n7289 25.1912
R4494 VPWR.n7356 VPWR.n7355 25.1912
R4495 VPWR.n7351 VPWR.n7350 25.1912
R4496 VPWR.n107 VPWR.n106 25.1912
R4497 VPWR.n9156 VPWR.n52 25.1912
R4498 VPWR.n9162 VPWR.n9161 25.1912
R4499 VPWR.n9168 VPWR.n9167 25.1912
R4500 VPWR.n9193 VPWR.n9192 25.1912
R4501 VPWR.n6081 VPWR.n6065 25.1912
R4502 VPWR.n6074 VPWR.n6071 25.1912
R4503 VPWR.n242 VPWR.n211 25.1912
R4504 VPWR.n8905 VPWR.n8904 25.1912
R4505 VPWR.n8168 VPWR.n8123 25.1912
R4506 VPWR.n8332 VPWR.n8331 25.1912
R4507 VPWR.n8316 VPWR.n5929 25.1912
R4508 VPWR.n8289 VPWR.n5938 25.1912
R4509 VPWR.n8773 VPWR.n8772 25.1912
R4510 VPWR.n8633 VPWR.n8632 25.1912
R4511 VPWR.n8656 VPWR.n8655 25.1912
R4512 VPWR.n867 VPWR.n800 25.1912
R4513 VPWR.n2556 VPWR.n2553 25.1912
R4514 VPWR.n2456 VPWR.n2455 25.1912
R4515 VPWR.n4467 VPWR.n4463 25.1912
R4516 VPWR.n3585 VPWR.n3578 25.1912
R4517 VPWR.n3397 VPWR.n3395 25.1912
R4518 VPWR.n3745 VPWR.n3744 25.1912
R4519 VPWR.n3669 VPWR.n3668 25.1912
R4520 VPWR.n7075 VPWR.n7070 25.1912
R4521 VPWR.t2819 VPWR.t169 25.1772
R4522 VPWR.t255 VPWR.t2869 25.1772
R4523 VPWR.t166 VPWR.t2673 25.1772
R4524 VPWR.t205 VPWR.t2187 25.1772
R4525 VPWR.t2197 VPWR.t1288 25.1772
R4526 VPWR.t463 VPWR.t3161 25.1772
R4527 VPWR.t2763 VPWR.t1385 25.1772
R4528 VPWR.t515 VPWR 25.1772
R4529 VPWR.t83 VPWR 25.1772
R4530 VPWR.t3007 VPWR.t2946 25.1772
R4531 VPWR.t1144 VPWR.t125 25.1772
R4532 VPWR.n7471 VPWR.n7470 24.8476
R4533 VPWR.n7401 VPWR.n7032 24.8476
R4534 VPWR.n4061 VPWR.n4060 24.8476
R4535 VPWR.n6055 VPWR.n6054 24.8476
R4536 VPWR.n8888 VPWR.n8887 24.8476
R4537 VPWR.n5798 VPWR.n5797 24.8476
R4538 VPWR.n425 VPWR.n411 24.8476
R4539 VPWR.n1575 VPWR.n1574 24.8476
R4540 VPWR.n5283 VPWR.n5282 24.8476
R4541 VPWR.n3500 VPWR.n3499 24.8476
R4542 VPWR.n7115 VPWR.n7113 24.8476
R4543 VPWR.n7192 VPWR.n7191 24.8476
R4544 VPWR.n7394 VPWR.n7393 24.7608
R4545 VPWR.n1458 VPWR.n1457 24.5271
R4546 VPWR.n947 VPWR.n946 24.5034
R4547 VPWR.n716 VPWR.n715 24.4711
R4548 VPWR.n8891 VPWR.n8870 24.4711
R4549 VPWR.n5805 VPWR.n5804 24.4711
R4550 VPWR.n4750 VPWR.n4749 24.4711
R4551 VPWR.n5295 VPWR.n546 24.4711
R4552 VPWR.n1947 VPWR.n1899 24.4711
R4553 VPWR.n5101 VPWR.n5100 24.4711
R4554 VPWR.n2231 VPWR.n2230 24.4711
R4555 VPWR.n7463 VPWR.n6953 24.0946
R4556 VPWR.n7553 VPWR.n7552 24.0946
R4557 VPWR.n7394 VPWR.n7033 24.0946
R4558 VPWR.n4073 VPWR.n2990 24.0946
R4559 VPWR.n5413 VPWR.n5412 24.0946
R4560 VPWR.n4685 VPWR.n4647 24.0946
R4561 VPWR.n5276 VPWR.n1785 24.0946
R4562 VPWR.n7184 VPWR.n7147 24.0946
R4563 VPWR.n8676 VPWR.n8675 23.7181
R4564 VPWR.n806 VPWR.n714 23.7181
R4565 VPWR.n2569 VPWR.n2115 23.7181
R4566 VPWR.n2693 VPWR.n2031 23.7181
R4567 VPWR.n7461 VPWR.n7460 23.7181
R4568 VPWR.n7460 VPWR.n6954 23.7181
R4569 VPWR.n7066 VPWR.n7046 23.7181
R4570 VPWR.n3072 VPWR.n3071 23.7181
R4571 VPWR.n3876 VPWR.n3039 23.7181
R4572 VPWR.n3876 VPWR.n3040 23.7181
R4573 VPWR.n8184 VPWR.n8117 23.7181
R4574 VPWR.n8679 VPWR.n352 23.7181
R4575 VPWR.n8423 VPWR.n5879 23.7181
R4576 VPWR.n6449 VPWR.n6349 23.7181
R4577 VPWR.n6450 VPWR.n6449 23.7181
R4578 VPWR.n6517 VPWR.n6489 23.7181
R4579 VPWR.n6521 VPWR.n6489 23.7181
R4580 VPWR.n1207 VPWR.n712 23.7181
R4581 VPWR.n825 VPWR.n712 23.7181
R4582 VPWR.n609 VPWR.n601 23.7181
R4583 VPWR.n639 VPWR.n593 23.7181
R4584 VPWR.n439 VPWR.n438 23.7181
R4585 VPWR.n5593 VPWR.n469 23.7181
R4586 VPWR.n1578 VPWR.n1543 23.7181
R4587 VPWR.n1951 VPWR.n1899 23.7181
R4588 VPWR.n5115 VPWR.n1840 23.7181
R4589 VPWR.n2440 VPWR.n2432 23.7181
R4590 VPWR.n4481 VPWR.n1998 23.7181
R4591 VPWR.n4247 VPWR.n2792 23.7181
R4592 VPWR.n3387 VPWR.n3386 23.7181
R4593 VPWR.n7070 VPWR.n7046 23.7181
R4594 VPWR.n2372 VPWR.n2299 23.6853
R4595 VPWR.n640 VPWR.n639 23.5104
R4596 VPWR.t2100 VPWR 23.4987
R4597 VPWR.t1552 VPWR.t1933 23.4987
R4598 VPWR VPWR.t2214 23.4987
R4599 VPWR.t1303 VPWR.t2897 23.4987
R4600 VPWR VPWR.t1896 23.4987
R4601 VPWR.t591 VPWR.t1429 23.4987
R4602 VPWR.t646 VPWR.t764 23.4987
R4603 VPWR.t116 VPWR.t2574 23.4987
R4604 VPWR.t1459 VPWR 23.4987
R4605 VPWR VPWR.t2888 23.4987
R4606 VPWR VPWR.t2742 23.4987
R4607 VPWR.n5817 VPWR.n5816 23.3417
R4608 VPWR.n993 VPWR.n992 23.3417
R4609 VPWR.n5593 VPWR.n5592 23.3417
R4610 VPWR.n4119 VPWR.n4118 22.9652
R4611 VPWR.n8142 VPWR.n8141 22.9652
R4612 VPWR.n8763 VPWR.n8762 22.9652
R4613 VPWR.n6523 VPWR.n6521 22.9652
R4614 VPWR.n840 VPWR.n818 22.9652
R4615 VPWR.n622 VPWR.n621 22.9652
R4616 VPWR.n1853 VPWR.n1851 22.9652
R4617 VPWR.n3418 VPWR.n3370 22.9652
R4618 VPWR.n6512 VPWR.n6491 22.9323
R4619 VPWR.n4073 VPWR.n2989 22.8518
R4620 VPWR.n616 VPWR.n600 22.5887
R4621 VPWR.n4749 VPWR.n4697 22.5887
R4622 VPWR.n5296 VPWR.n5295 22.5887
R4623 VPWR.n2569 VPWR.n2114 22.5887
R4624 VPWR.n5745 VPWR.n5744 22.5559
R4625 VPWR.n3042 VPWR.n3039 22.2123
R4626 VPWR.n3261 VPWR.n3234 22.2123
R4627 VPWR.n8424 VPWR.n8423 22.2123
R4628 VPWR.n8493 VPWR.n5861 22.2123
R4629 VPWR.n6535 VPWR.n6534 22.2123
R4630 VPWR.n612 VPWR.n601 22.2123
R4631 VPWR.n613 VPWR.n612 22.2123
R4632 VPWR.n443 VPWR.n403 22.2123
R4633 VPWR.n5607 VPWR.n5606 22.2123
R4634 VPWR.n1913 VPWR.n1892 22.2123
R4635 VPWR.n1849 VPWR.n1848 22.2123
R4636 VPWR.n5119 VPWR.n1840 22.2123
R4637 VPWR.n5120 VPWR.n5119 22.2123
R4638 VPWR.n2318 VPWR.n2316 22.2123
R4639 VPWR.n2322 VPWR.n2316 22.2123
R4640 VPWR.n3413 VPWR.n3411 22.2123
R4641 VPWR.n3413 VPWR.n3370 22.2123
R4642 VPWR.n445 VPWR.n443 22.1175
R4643 VPWR.t282 VPWR.t2818 21.8203
R4644 VPWR.t2315 VPWR.n6110 21.8203
R4645 VPWR.t2880 VPWR.t3259 21.8203
R4646 VPWR.t2297 VPWR.t6 21.8203
R4647 VPWR.t3190 VPWR.t1970 21.8203
R4648 VPWR.t1502 VPWR 21.8203
R4649 VPWR.t1223 VPWR 21.8203
R4650 VPWR.t60 VPWR.t1661 21.8203
R4651 VPWR.t1227 VPWR.t2768 21.8203
R4652 VPWR.t3065 VPWR 21.8203
R4653 VPWR.t249 VPWR.t1311 21.8203
R4654 VPWR.t1508 VPWR.t1095 21.8203
R4655 VPWR.t1886 VPWR.t2274 21.8203
R4656 VPWR.t2106 VPWR.t1147 21.8203
R4657 VPWR.t1682 VPWR 21.8203
R4658 VPWR.t1858 VPWR.t756 21.8203
R4659 VPWR.n4418 VPWR.n4414 21.7466
R4660 VPWR.n3266 VPWR.n3265 21.4593
R4661 VPWR.n6108 VPWR.n6010 21.4593
R4662 VPWR.n8305 VPWR.n8304 21.4593
R4663 VPWR.n6602 VPWR.n6599 21.4593
R4664 VPWR.n8684 VPWR.n8683 21.4593
R4665 VPWR.n5434 VPWR.n499 21.4593
R4666 VPWR.n5018 VPWR.n1890 21.4593
R4667 VPWR.n2327 VPWR.n2326 21.4593
R4668 VPWR.n4463 VPWR.n2006 21.4593
R4669 VPWR.n3730 VPWR.n3729 21.4593
R4670 VPWR.n1771 VPWR.n549 21.0829
R4671 VPWR.n2312 VPWR.n2311 21.0829
R4672 VPWR.n4770 VPWR.n4635 20.9962
R4673 VPWR.n3885 VPWR.n3032 20.8852
R4674 VPWR.n6293 VPWR.n6292 20.8852
R4675 VPWR.n5638 VPWR.n5637 20.8852
R4676 VPWR.n2445 VPWR.n2444 20.7064
R4677 VPWR.n8437 VPWR.n5866 20.5266
R4678 VPWR.n3175 VPWR.n3174 20.3859
R4679 VPWR.n9186 VPWR.n9185 20.297
R4680 VPWR.t840 VPWR 20.1418
R4681 VPWR.t1590 VPWR.t1793 20.1418
R4682 VPWR.t1252 VPWR.n1204 20.1418
R4683 VPWR.t1089 VPWR.t1373 20.1418
R4684 VPWR.t2781 VPWR.n471 20.1418
R4685 VPWR VPWR.t1043 20.1418
R4686 VPWR.n3913 VPWR.n3911 20.0749
R4687 VPWR.n6760 VPWR.n6752 20.0749
R4688 VPWR.n6071 VPWR.n26 19.9534
R4689 VPWR.n6599 VPWR.n6588 19.9534
R4690 VPWR.n8608 VPWR.n8607 19.9534
R4691 VPWR.n6517 VPWR.n6516 19.9534
R4692 VPWR.n4685 VPWR.n4684 19.9534
R4693 VPWR.n5142 VPWR.n5141 19.9534
R4694 VPWR.n4428 VPWR.n2008 19.9534
R4695 VPWR.n5317 VPWR.n538 19.7491
R4696 VPWR.n4122 VPWR.n4088 19.577
R4697 VPWR.n83 VPWR.n72 19.577
R4698 VPWR.n9205 VPWR.n9204 19.577
R4699 VPWR.n226 VPWR.n214 19.577
R4700 VPWR.n1201 VPWR.n722 19.577
R4701 VPWR.n4758 VPWR.n4757 19.577
R4702 VPWR.n5028 VPWR.n1889 19.577
R4703 VPWR.n4429 VPWR.n4428 19.5476
R4704 VPWR.n1197 VPWR.n719 19.5441
R4705 VPWR.n2336 VPWR.n2335 19.4073
R4706 VPWR.n6726 VPWR.n6725 19.2067
R4707 VPWR.n6408 VPWR.n6407 19.2067
R4708 VPWR.n4828 VPWR.n4827 19.2067
R4709 VPWR.n7764 VPWR.n7763 19.0176
R4710 VPWR.n6238 VPWR.n6237 19.0176
R4711 VPWR.n6182 VPWR.n6158 18.824
R4712 VPWR.n3741 VPWR.n3497 18.824
R4713 VPWR.n6089 VPWR.n6088 18.7912
R4714 VPWR.n3407 VPWR.n3371 18.7912
R4715 VPWR.n426 VPWR.n425 18.7213
R4716 VPWR.t2217 VPWR.t793 18.4634
R4717 VPWR VPWR.t877 18.4634
R4718 VPWR.t3195 VPWR 18.4634
R4719 VPWR.t818 VPWR.t2046 18.4634
R4720 VPWR.t810 VPWR.t3325 18.4634
R4721 VPWR.t2702 VPWR 18.4634
R4722 VPWR.t1129 VPWR 18.4634
R4723 VPWR.t1103 VPWR.t2362 18.4634
R4724 VPWR.t2177 VPWR.t2541 18.4634
R4725 VPWR VPWR.t1183 18.4634
R4726 VPWR.t754 VPWR.t848 18.4634
R4727 VPWR.t3064 VPWR.t1193 18.4634
R4728 VPWR.t1040 VPWR.t1403 18.4634
R4729 VPWR.n8128 VPWR.n8113 18.4476
R4730 VPWR.n1111 VPWR.n1110 18.4476
R4731 VPWR.n4479 VPWR.n4478 18.4476
R4732 VPWR.n2796 VPWR.n2791 18.4476
R4733 VPWR.n3536 VPWR.n3520 18.4476
R4734 VPWR.n7535 VPWR.n7534 18.4147
R4735 VPWR.n7373 VPWR.n7372 18.4147
R4736 VPWR.n7160 VPWR.n7155 18.4147
R4737 VPWR.n968 VPWR.n967 18.2862
R4738 VPWR.n8888 VPWR.n8871 18.0711
R4739 VPWR.n6612 VPWR.n6611 18.0711
R4740 VPWR.n5798 VPWR.n5781 18.0711
R4741 VPWR.n848 VPWR.n816 18.0711
R4742 VPWR.n1931 VPWR.n1930 17.6946
R4743 VPWR.n7571 VPWR.n7569 17.612
R4744 VPWR.n8283 VPWR.n8282 17.612
R4745 VPWR.n3596 VPWR.n3594 17.612
R4746 VPWR.n3663 VPWR.n3662 17.612
R4747 VPWR.n7082 VPWR.n7080 17.612
R4748 VPWR.n7499 VPWR.n7498 17.612
R4749 VPWR.n3288 VPWR.n3285 17.612
R4750 VPWR.n3720 VPWR.n3719 17.612
R4751 VPWR.n6177 VPWR.n6176 17.3181
R4752 VPWR.n8498 VPWR.n8497 17.3181
R4753 VPWR.n1412 VPWR.n1410 17.3181
R4754 VPWR.n1441 VPWR.n1440 17.3181
R4755 VPWR.n1440 VPWR.n1439 17.3181
R4756 VPWR.n1940 VPWR.n1939 17.3181
R4757 VPWR.n3055 VPWR.n3054 17.2853
R4758 VPWR.n2726 VPWR.n2021 17.2339
R4759 VPWR.n4126 VPWR.n4088 16.9977
R4760 VPWR.n6595 VPWR.n6588 16.9417
R4761 VPWR.n1554 VPWR.n1553 16.9417
R4762 VPWR.n2223 VPWR.n2222 16.9417
R4763 VPWR.n4503 VPWR.n4496 16.9417
R4764 VPWR.t600 VPWR.t1302 16.785
R4765 VPWR VPWR.t1201 16.785
R4766 VPWR.t1038 VPWR.t1598 16.785
R4767 VPWR.t3154 VPWR.t1371 16.785
R4768 VPWR.t2862 VPWR 16.785
R4769 VPWR.t3121 VPWR.t2866 16.785
R4770 VPWR.n8438 VPWR.n8437 16.7729
R4771 VPWR.n4509 VPWR.n4508 16.6212
R4772 VPWR.n7107 VPWR.n7106 16.6212
R4773 VPWR.n1715 VPWR.n1714 16.5652
R4774 VPWR.n1515 VPWR.n1513 16.4701
R4775 VPWR.n5452 VPWR.n5451 16.4179
R4776 VPWR.n9175 VPWR.n9174 16.1887
R4777 VPWR.n8187 VPWR.n8113 16.1887
R4778 VPWR.n1090 VPWR.n1087 16.1887
R4779 VPWR.n998 VPWR.n997 16.1887
R4780 VPWR.n4697 VPWR.n4696 16.1887
R4781 VPWR.n4948 VPWR.n4947 16.1887
R4782 VPWR.n2260 VPWR.n2259 16.1887
R4783 VPWR.n4478 VPWR.n4477 16.1887
R4784 VPWR.n4250 VPWR.n2791 16.1887
R4785 VPWR.n3675 VPWR.n3520 16.1887
R4786 VPWR.n7656 VPWR.n7654 16.139
R4787 VPWR.n8017 VPWR.n8014 16.139
R4788 VPWR.n2183 VPWR.n2120 16.139
R4789 VPWR.n936 VPWR.n934 16.0189
R4790 VPWR.n2922 VPWR.n2921 15.995
R4791 VPWR.n7514 VPWR.n7513 15.8683
R4792 VPWR.n4002 VPWR.n2998 15.8683
R4793 VPWR.n3216 VPWR.n3215 15.8683
R4794 VPWR.n9047 VPWR.n9046 15.8683
R4795 VPWR.n4802 VPWR.n4801 15.8683
R4796 VPWR.n1669 VPWR.n1668 15.8683
R4797 VPWR.n4247 VPWR.n2794 15.8683
R4798 VPWR.n3672 VPWR.n3523 15.8683
R4799 VPWR.n3692 VPWR.n3691 15.8683
R4800 VPWR.n3744 VPWR.n3497 15.8123
R4801 VPWR.n9145 VPWR.n9144 15.7465
R4802 VPWR.n5015 VPWR.n1898 15.7465
R4803 VPWR.n2465 VPWR.n2426 15.7465
R4804 VPWR.n954 VPWR.n947 15.7306
R4805 VPWR.n2092 VPWR.n2091 15.7262
R4806 VPWR.n9137 VPWR.n9136 15.6908
R4807 VPWR.n6670 VPWR.n6669 15.6908
R4808 VPWR.n8679 VPWR.n354 15.4358
R4809 VPWR.n1217 VPWR.n1216 15.4358
R4810 VPWR.n5312 VPWR.n540 15.3605
R4811 VPWR.n8439 VPWR.n5865 15.2281
R4812 VPWR.t2739 VPWR 15.1065
R4813 VPWR.t1181 VPWR 15.1065
R4814 VPWR.t1781 VPWR.t3323 15.1065
R4815 VPWR.t1484 VPWR.t3310 15.1065
R4816 VPWR.t2327 VPWR.t2915 15.1065
R4817 VPWR.t2024 VPWR.t2309 15.1065
R4818 VPWR.t1647 VPWR.t2022 15.1065
R4819 VPWR.t2191 VPWR.t3176 15.1065
R4820 VPWR.t2073 VPWR.t3209 15.1065
R4821 VPWR.t1930 VPWR 15.1065
R4822 VPWR.n5812 VPWR.n5811 15.0593
R4823 VPWR.n5453 VPWR.n5452 15.0593
R4824 VPWR.n4757 VPWR.n4756 15.0593
R4825 VPWR.n5031 VPWR.n1889 15.0593
R4826 VPWR.n8197 VPWR.n8109 15.0265
R4827 VPWR.n967 VPWR.n966 14.9948
R4828 VPWR.n4710 VPWR.n4708 14.9948
R4829 VPWR.n6541 VPWR.n6537 14.7405
R4830 VPWR.n6516 VPWR.n6515 14.6829
R4831 VPWR.n1034 VPWR.n1033 14.6829
R4832 VPWR.n2689 VPWR.n2034 14.6829
R4833 VPWR.n1775 VPWR.n549 14.65
R4834 VPWR.n7124 VPWR.n7123 14.65
R4835 VPWR.n3871 VPWR.n3042 14.6331
R4836 VPWR.n7954 VPWR.n7953 14.6253
R4837 VPWR.n2898 VPWR.n2897 14.5851
R4838 VPWR.n5124 VPWR.n5123 14.4976
R4839 VPWR.n8491 VPWR.n5862 14.3624
R4840 VPWR.n291 VPWR.n290 14.3615
R4841 VPWR.n6186 VPWR.n6158 14.3064
R4842 VPWR.n8599 VPWR.n8595 14.3064
R4843 VPWR.n5282 VPWR.n1783 14.3064
R4844 VPWR.n7380 VPWR.n7379 14.2735
R4845 VPWR.n7379 VPWR.n7045 14.2735
R4846 VPWR.n4105 VPWR.n4104 14.2735
R4847 VPWR.n3252 VPWR.n3249 14.2735
R4848 VPWR.n8748 VPWR.n8747 14.2735
R4849 VPWR.n6502 VPWR.n6499 14.2735
R4850 VPWR.n1120 VPWR.n717 14.2735
R4851 VPWR.n857 VPWR.n856 14.2735
R4852 VPWR.n1292 VPWR.n1291 14.2735
R4853 VPWR.n4930 VPWR.n4929 14.2735
R4854 VPWR.n5007 VPWR.n5006 14.2735
R4855 VPWR.n2566 VPWR.n2565 14.2735
R4856 VPWR.n2049 VPWR.n2031 14.2735
R4857 VPWR.n7278 VPWR.n7047 14.2735
R4858 VPWR.n535 VPWR.n533 14.2634
R4859 VPWR.n533 VPWR.n528 14.2634
R4860 VPWR.n8150 VPWR.n8149 13.9299
R4861 VPWR.n960 VPWR.n959 13.902
R4862 VPWR.n4713 VPWR.n4710 13.8976
R4863 VPWR.n7762 VPWR.n7761 13.8687
R4864 VPWR.n6235 VPWR.n6234 13.8687
R4865 VPWR.n7278 VPWR.n7277 13.8432
R4866 VPWR.n68 VPWR.n64 13.5534
R4867 VPWR.n1113 VPWR.n731 13.5534
R4868 VPWR.n4424 VPWR.n2008 13.5534
R4869 VPWR.n231 VPWR.n230 13.5206
R4870 VPWR.n6376 VPWR.n6375 13.5206
R4871 VPWR.n5605 VPWR.n5604 13.5206
R4872 VPWR.t2428 VPWR.t1008 13.4281
R4873 VPWR.t1239 VPWR 13.4281
R4874 VPWR.t3170 VPWR.t3227 13.4281
R4875 VPWR.t652 VPWR.t1036 13.4281
R4876 VPWR.t2875 VPWR.t1099 13.4281
R4877 VPWR.t2140 VPWR.t2240 13.4281
R4878 VPWR.t2616 VPWR.t2236 13.4281
R4879 VPWR.t1620 VPWR.t1018 13.4281
R4880 VPWR VPWR.t846 13.4281
R4881 VPWR.t696 VPWR.t1455 13.4281
R4882 VPWR.n4068 VPWR.n2989 13.4209
R4883 VPWR.n7513 VPWR.n6942 13.177
R4884 VPWR.n3269 VPWR.n3268 13.177
R4885 VPWR.n80 VPWR.n73 13.177
R4886 VPWR.n6055 VPWR.n6010 13.177
R4887 VPWR.n223 VPWR.n216 13.177
R4888 VPWR.n8881 VPWR.n8874 13.177
R4889 VPWR.n8299 VPWR.n8298 13.177
R4890 VPWR.n8687 VPWR.n8686 13.177
R4891 VPWR.n5792 VPWR.n5785 13.177
R4892 VPWR.n1143 VPWR.n1142 13.177
R4893 VPWR.n419 VPWR.n412 13.177
R4894 VPWR.n1785 VPWR.n1784 13.177
R4895 VPWR.n2684 VPWR.n2683 13.177
R4896 VPWR.n3729 VPWR.n3500 13.177
R4897 VPWR.n2833 VPWR.n2832 13.1523
R4898 VPWR.n2130 VPWR.n2115 12.961
R4899 VPWR.n2832 VPWR.n2795 12.961
R4900 VPWR.n4006 VPWR.n2998 12.8005
R4901 VPWR.n7654 VPWR.n7646 12.8005
R4902 VPWR.n6176 VPWR.n6175 12.8005
R4903 VPWR.n9047 VPWR.n198 12.8005
R4904 VPWR.n6671 VPWR.n6657 12.8005
R4905 VPWR.n8184 VPWR.n8116 12.8005
R4906 VPWR.n8425 VPWR.n5872 12.8005
R4907 VPWR.n6364 VPWR.n6349 12.8005
R4908 VPWR.n731 VPWR.n717 12.8005
R4909 VPWR.n1035 VPWR.n1034 12.8005
R4910 VPWR.n621 VPWR.n600 12.8005
R4911 VPWR.n1412 VPWR.n1411 12.8005
R4912 VPWR.n1291 VPWR.n1283 12.8005
R4913 VPWR.n4767 VPWR.n4642 12.8005
R4914 VPWR.n2566 VPWR.n2120 12.8005
R4915 VPWR.n2016 VPWR.n2009 12.8005
R4916 VPWR.n4414 VPWR.n2009 12.8005
R4917 VPWR.n3386 VPWR.n3378 12.8005
R4918 VPWR.n1307 VPWR.n1306 12.5338
R4919 VPWR.n70 VPWR.n68 12.0476
R4920 VPWR.n6694 VPWR.n6657 12.0476
R4921 VPWR.n8325 VPWR.n8324 12.0476
R4922 VPWR.n6695 VPWR.n6694 12.0476
R4923 VPWR.n8762 VPWR.n8736 12.0476
R4924 VPWR.n8691 VPWR.n8690 12.0476
R4925 VPWR.n8650 VPWR.n8648 12.0476
R4926 VPWR.n5147 VPWR.n5146 12.0476
R4927 VPWR.n2572 VPWR.n2114 12.0476
R4928 VPWR.n2249 VPWR.n2248 12.0476
R4929 VPWR.n3420 VPWR.n3418 12.0147
R4930 VPWR.t2144 VPWR 11.7496
R4931 VPWR.t1069 VPWR.t1323 11.7496
R4932 VPWR.t2026 VPWR.t1145 11.7496
R4933 VPWR.t2189 VPWR.t2030 11.7496
R4934 VPWR.n4060 VPWR.n2995 11.7271
R4935 VPWR.n72 VPWR.n70 11.6711
R4936 VPWR.n35 VPWR.n34 11.6711
R4937 VPWR.n230 VPWR.n214 11.6711
R4938 VPWR.n1716 VPWR.n554 11.6382
R4939 VPWR.n3881 VPWR.n3038 11.4366
R4940 VPWR.n251 VPWR.n250 11.2946
R4941 VPWR.n8328 VPWR.n8327 11.2946
R4942 VPWR.n8425 VPWR.n8424 11.2946
R4943 VPWR.n5818 VPWR.n5817 11.2946
R4944 VPWR.n1015 VPWR.n1014 11.2946
R4945 VPWR.n992 VPWR.n716 11.2946
R4946 VPWR.n5592 VPWR.n5591 11.2946
R4947 VPWR.n5018 VPWR.n1892 11.2946
R4948 VPWR.n4955 VPWR.n4913 11.2946
R4949 VPWR.n3258 VPWR.n3257 11.2618
R4950 VPWR.n8758 VPWR.n8736 11.2618
R4951 VPWR.n3215 VPWR.n3146 11.0456
R4952 VPWR.n973 VPWR.n972 10.9719
R4953 VPWR.n4733 VPWR.n4730 10.9719
R4954 VPWR.n2098 VPWR.n2097 10.9719
R4955 VPWR.n3161 VPWR.n3160 10.9181
R4956 VPWR.n1850 VPWR.n1849 10.9181
R4957 VPWR.n5613 VPWR.n5612 10.9013
R4958 VPWR.n3280 VPWR.n3278 10.8853
R4959 VPWR.n6104 VPWR.n6058 10.8853
R4960 VPWR.n8152 VPWR.n8150 10.8853
R4961 VPWR.n8675 VPWR.n8615 10.8853
R4962 VPWR.n5933 VPWR.n5932 10.6672
R4963 VPWR.n4118 VPWR.n4117 10.5744
R4964 VPWR.n8626 VPWR.n8621 10.5417
R4965 VPWR.n1201 VPWR.n719 10.5417
R4966 VPWR.n627 VPWR.n626 10.4965
R4967 VPWR.n4639 VPWR.n4638 10.2593
R4968 VPWR.n2695 VPWR.n2693 10.2499
R4969 VPWR.n102 VPWR.n101 10.1652
R4970 VPWR.n5419 VPWR.n5418 10.1652
R4971 VPWR.n6380 VPWR.n6378 10.1592
R4972 VPWR.t2096 VPWR.t3003 10.0712
R4973 VPWR.t2039 VPWR.t1888 10.0712
R4974 VPWR VPWR.t2499 10.0712
R4975 VPWR.t1030 VPWR.t1308 10.0712
R4976 VPWR.t2410 VPWR 10.0712
R4977 VPWR.t1284 VPWR.t1315 10.0712
R4978 VPWR.t1326 VPWR.t234 10.0712
R4979 VPWR.t1462 VPWR.t2640 10.0712
R4980 VPWR.t2150 VPWR.t2234 10.0712
R4981 VPWR.t1059 VPWR.t2122 10.0712
R4982 VPWR.t1191 VPWR.t3280 10.0712
R4983 VPWR.t403 VPWR.t2225 10.0712
R4984 VPWR.t1024 VPWR.t2886 10.0712
R4985 VPWR.t1534 VPWR.t937 10.0712
R4986 VPWR.t1139 VPWR.t2567 10.0712
R4987 VPWR.n6652 VPWR.n6650 10.0005
R4988 VPWR.n836 VPWR.n834 10.0005
R4989 VPWR.n9179 VPWR.n9178 9.91684
R4990 VPWR.n4074 VPWR.n4073 9.8812
R4991 VPWR.n5491 VPWR.n5490 9.8812
R4992 VPWR.n4771 VPWR.n4770 9.8812
R4993 VPWR.n8493 VPWR.n8491 9.78874
R4994 VPWR.n1565 VPWR.n1564 9.78874
R4995 VPWR.n1936 VPWR.n1935 9.78874
R4996 VPWR.n5151 VPWR.n5150 9.78874
R4997 VPWR.n3089 VPWR.n3088 9.73273
R4998 VPWR.n3206 VPWR.n3205 9.73273
R4999 VPWR.n7664 VPWR.n7639 9.73273
R5000 VPWR.n7671 VPWR.n7670 9.73273
R5001 VPWR.n7756 VPWR.n6128 9.73273
R5002 VPWR.n9030 VPWR.n9029 9.73273
R5003 VPWR.n9050 VPWR.n196 9.73273
R5004 VPWR.n6272 VPWR.n6271 9.73273
R5005 VPWR.n8261 VPWR.n8260 9.73273
R5006 VPWR.n6765 VPWR.n6643 9.73273
R5007 VPWR.n6634 VPWR.n6586 9.73273
R5008 VPWR.n8466 VPWR.n5864 9.73273
R5009 VPWR.n6385 VPWR.n6384 9.73273
R5010 VPWR.n6412 VPWR.n6411 9.73273
R5011 VPWR.n6446 VPWR.n6351 9.73273
R5012 VPWR.n6446 VPWR.n6445 9.73273
R5013 VPWR.n5642 VPWR.n451 9.73273
R5014 VPWR.n5643 VPWR.n5642 9.73273
R5015 VPWR.n5621 VPWR.n458 9.73273
R5016 VPWR.n5627 VPWR.n457 9.73273
R5017 VPWR.n5495 VPWR.n5494 9.73273
R5018 VPWR.n5486 VPWR.n5485 9.73273
R5019 VPWR.n1500 VPWR.n1499 9.73273
R5020 VPWR.n1499 VPWR.n1374 9.73273
R5021 VPWR.n1495 VPWR.n1494 9.73273
R5022 VPWR.n4824 VPWR.n4823 9.73273
R5023 VPWR.n4823 VPWR.n4790 9.73273
R5024 VPWR.n4819 VPWR.n4818 9.73273
R5025 VPWR.n4818 VPWR.n4791 9.73273
R5026 VPWR.n4814 VPWR.n4791 9.73273
R5027 VPWR.n1661 VPWR.n560 9.73273
R5028 VPWR.n1662 VPWR.n1661 9.73273
R5029 VPWR.n2718 VPWR.n2022 9.73273
R5030 VPWR.n4518 VPWR.n4488 9.73273
R5031 VPWR.n4514 VPWR.n4513 9.73273
R5032 VPWR.n4513 VPWR.n4492 9.73273
R5033 VPWR.n3612 VPWR.n3525 9.73273
R5034 VPWR.n3643 VPWR.n3642 9.73273
R5035 VPWR.n3886 VPWR.n3885 9.65664
R5036 VPWR.n6293 VPWR.n6288 9.65664
R5037 VPWR.n5638 VPWR.n452 9.65664
R5038 VPWR.n5491 VPWR.n486 9.65664
R5039 VPWR.n1321 VPWR.n1320 9.62695
R5040 VPWR.n4116 VPWR.n4115 9.6005
R5041 VPWR.n8261 VPWR.n5948 9.52116
R5042 VPWR.n1316 VPWR.n1315 9.52116
R5043 VPWR.n3613 VPWR.n3612 9.52116
R5044 VPWR.n1138 VPWR.n1137 9.41227
R5045 VPWR.n861 VPWR.n806 9.41227
R5046 VPWR.n2257 VPWR.n2214 9.41227
R5047 VPWR.n3738 VPWR.n3737 9.41227
R5048 VPWR.n5449 VPWR.n5447 9.38145
R5049 VPWR.n1208 VPWR.n1207 9.32328
R5050 VPWR.n196 VPWR.n195 9.30959
R5051 VPWR.n1494 VPWR.n1375 9.30959
R5052 VPWR.n6876 VPWR.n6875 9.3005
R5053 VPWR.n6224 VPWR.n6223 9.3005
R5054 VPWR.n6874 VPWR.n6873 9.3005
R5055 VPWR.n260 VPWR.n259 9.3005
R5056 VPWR.n294 VPWR.n293 9.3005
R5057 VPWR.n271 VPWR.n270 9.3005
R5058 VPWR.n262 VPWR.n261 9.3005
R5059 VPWR.n8069 VPWR.n8068 9.3005
R5060 VPWR.n8067 VPWR.n8066 9.3005
R5061 VPWR.n6798 VPWR.n6797 9.3005
R5062 VPWR.n6826 VPWR.n6825 9.3005
R5063 VPWR.n6807 VPWR.n6806 9.3005
R5064 VPWR.n6796 VPWR.n6795 9.3005
R5065 VPWR.n8847 VPWR.n8846 9.3005
R5066 VPWR.n8922 VPWR.n8921 9.3005
R5067 VPWR.n8837 VPWR.n8836 9.3005
R5068 VPWR.n8839 VPWR.n8838 9.3005
R5069 VPWR.n6472 VPWR.n6471 9.3005
R5070 VPWR.n6480 VPWR.n6479 9.3005
R5071 VPWR.n6469 VPWR.n6468 9.3005
R5072 VPWR.n8712 VPWR.n8711 9.3005
R5073 VPWR.n8793 VPWR.n8792 9.3005
R5074 VPWR.n8795 VPWR.n8794 9.3005
R5075 VPWR.n8715 VPWR.n8714 9.3005
R5076 VPWR.n5833 VPWR.n5832 9.3005
R5077 VPWR.n5835 VPWR.n5834 9.3005
R5078 VPWR.n5748 VPWR.n5747 9.3005
R5079 VPWR.n5750 VPWR.n5749 9.3005
R5080 VPWR.n656 VPWR.n655 9.3005
R5081 VPWR.n699 VPWR.n698 9.3005
R5082 VPWR.n1426 VPWR.n1425 9.3005
R5083 VPWR.n1335 VPWR.n1334 9.3005
R5084 VPWR.n1362 VPWR.n1361 9.3005
R5085 VPWR.n1364 VPWR.n1363 9.3005
R5086 VPWR.n5500 VPWR.n5499 9.3005
R5087 VPWR.n5681 VPWR.n5680 9.3005
R5088 VPWR.n5700 VPWR.n5699 9.3005
R5089 VPWR.n5698 VPWR.n5697 9.3005
R5090 VPWR.n5671 VPWR.n5670 9.3005
R5091 VPWR.n5673 VPWR.n5672 9.3005
R5092 VPWR.n5577 VPWR.n5576 9.3005
R5093 VPWR.n5574 VPWR.n5573 9.3005
R5094 VPWR.n5502 VPWR.n5501 9.3005
R5095 VPWR.n1393 VPWR.n1392 9.3005
R5096 VPWR.n1395 VPWR.n1394 9.3005
R5097 VPWR.n1423 VPWR.n1422 9.3005
R5098 VPWR.n1353 VPWR.n1352 9.3005
R5099 VPWR.n1337 VPWR.n1336 9.3005
R5100 VPWR.n1636 VPWR.n1635 9.3005
R5101 VPWR.n1791 VPWR.n1790 9.3005
R5102 VPWR.n4860 VPWR.n4859 9.3005
R5103 VPWR.n1793 VPWR.n1792 9.3005
R5104 VPWR.n1737 VPWR.n1736 9.3005
R5105 VPWR.n1739 VPWR.n1738 9.3005
R5106 VPWR.n1638 VPWR.n1637 9.3005
R5107 VPWR.n1588 VPWR.n1587 9.3005
R5108 VPWR.n2578 VPWR.n2577 9.3005
R5109 VPWR.n2540 VPWR.n2539 9.3005
R5110 VPWR.n5072 VPWR.n5071 9.3005
R5111 VPWR.n5033 VPWR.n5032 9.3005
R5112 VPWR.n5036 VPWR.n5035 9.3005
R5113 VPWR.n5074 VPWR.n5073 9.3005
R5114 VPWR.n2581 VPWR.n2580 9.3005
R5115 VPWR.n2543 VPWR.n2542 9.3005
R5116 VPWR.n2532 VPWR.n2531 9.3005
R5117 VPWR.n2528 VPWR.n2527 9.3005
R5118 VPWR.n4403 VPWR.n4402 9.3005
R5119 VPWR.n2680 VPWR.n2679 9.3005
R5120 VPWR.n4376 VPWR.n4375 9.3005
R5121 VPWR.n4398 VPWR.n4397 9.3005
R5122 VPWR.n4374 VPWR.n4373 9.3005
R5123 VPWR.n2650 VPWR.n2649 9.3005
R5124 VPWR.n2652 VPWR.n2651 9.3005
R5125 VPWR.n2677 VPWR.n2676 9.3005
R5126 VPWR.n3542 VPWR.n3541 9.3005
R5127 VPWR.n3490 VPWR.n3489 9.3005
R5128 VPWR.n4265 VPWR.n4264 9.3005
R5129 VPWR.n2938 VPWR.n2937 9.3005
R5130 VPWR.n4228 VPWR.n4227 9.3005
R5131 VPWR.n4226 VPWR.n4225 9.3005
R5132 VPWR.n4268 VPWR.n4267 9.3005
R5133 VPWR.n4289 VPWR.n4288 9.3005
R5134 VPWR.n4291 VPWR.n4290 9.3005
R5135 VPWR.n3545 VPWR.n3544 9.3005
R5136 VPWR.n3492 VPWR.n3491 9.3005
R5137 VPWR.n3466 VPWR.n3465 9.3005
R5138 VPWR.n7817 VPWR.n7816 9.3005
R5139 VPWR.n7690 VPWR.n7689 9.3005
R5140 VPWR.n7707 VPWR.n7706 9.3005
R5141 VPWR.n7688 VPWR.n7687 9.3005
R5142 VPWR.n7820 VPWR.n7819 9.3005
R5143 VPWR.n7842 VPWR.n7841 9.3005
R5144 VPWR.n7844 VPWR.n7843 9.3005
R5145 VPWR.n9206 VPWR.n9205 9.3005
R5146 VPWR.n9209 VPWR.n9208 9.3005
R5147 VPWR.n3296 VPWR.n3295 9.3005
R5148 VPWR.n3325 VPWR.n3324 9.3005
R5149 VPWR.n3869 VPWR.n3868 9.3005
R5150 VPWR.n3988 VPWR.n3987 9.3005
R5151 VPWR.n4156 VPWR.n4155 9.3005
R5152 VPWR.n4164 VPWR.n4163 9.3005
R5153 VPWR.n4138 VPWR.n4137 9.3005
R5154 VPWR.n4166 VPWR.n4165 9.3005
R5155 VPWR.n3985 VPWR.n3984 9.3005
R5156 VPWR.n3866 VPWR.n3865 9.3005
R5157 VPWR.n3842 VPWR.n3841 9.3005
R5158 VPWR.n3844 VPWR.n3843 9.3005
R5159 VPWR.n3314 VPWR.n3313 9.3005
R5160 VPWR.n3323 VPWR.n3322 9.3005
R5161 VPWR.n3294 VPWR.n3293 9.3005
R5162 VPWR.n7453 VPWR.n7452 9.3005
R5163 VPWR.n7579 VPWR.n7578 9.3005
R5164 VPWR.n7604 VPWR.n7603 9.3005
R5165 VPWR.n7577 VPWR.n7576 9.3005
R5166 VPWR.n7595 VPWR.n7594 9.3005
R5167 VPWR.n7606 VPWR.n7605 9.3005
R5168 VPWR.n7450 VPWR.n7449 9.3005
R5169 VPWR.n7430 VPWR.n7429 9.3005
R5170 VPWR.n7428 VPWR.n7427 9.3005
R5171 VPWR.n7198 VPWR.n7197 9.3005
R5172 VPWR.n7206 VPWR.n7205 9.3005
R5173 VPWR.n7196 VPWR.n7195 9.3005
R5174 VPWR.n7225 VPWR.n7224 9.3005
R5175 VPWR.n3643 VPWR.n3633 9.20381
R5176 VPWR.n5452 VPWR.n492 9.16726
R5177 VPWR.n4055 VPWR.n4054 9.09802
R5178 VPWR.n8260 VPWR.n5949 9.09802
R5179 VPWR.n6618 VPWR.n6617 9.09802
R5180 VPWR.n8461 VPWR.n5864 9.09802
R5181 VPWR.n6411 VPWR.n6353 9.09802
R5182 VPWR.n4824 VPWR.n4787 9.09802
R5183 VPWR.n1710 VPWR.n1709 9.09802
R5184 VPWR.n5606 VPWR.n5605 9.03579
R5185 VPWR.n1578 VPWR.n1577 9.03579
R5186 VPWR.n1716 VPWR.n1715 9.03579
R5187 VPWR.n2241 VPWR.n2240 9.03579
R5188 VPWR.n2689 VPWR.n2035 9.03579
R5189 VPWR.n3691 VPWR.n3690 9.03579
R5190 VPWR.n8831 VPWR.n8830 9.02415
R5191 VPWR.n6462 VPWR.n6461 9.02415
R5192 VPWR.n5742 VPWR.n5741 9.02415
R5193 VPWR.n1226 VPWR.n1225 9.02415
R5194 VPWR.n5664 VPWR.n5663 9.02415
R5195 VPWR.n1519 VPWR.n1518 9.02415
R5196 VPWR.n4997 VPWR.n4996 9.02415
R5197 VPWR.n3748 VPWR.n3747 9.02415
R5198 VPWR.n7957 VPWR.n7956 9.00388
R5199 VPWR.n6872 VPWR.n6871 9.0005
R5200 VPWR.n6879 VPWR.n6878 9.0005
R5201 VPWR.n6220 VPWR.n6219 9.0005
R5202 VPWR.n8077 VPWR.n8076 9.0005
R5203 VPWR.n8071 VPWR.n8070 9.0005
R5204 VPWR.n8064 VPWR.n8063 9.0005
R5205 VPWR.n200 VPWR.n199 9.0005
R5206 VPWR.n286 VPWR.n285 9.0005
R5207 VPWR.n276 VPWR.n275 9.0005
R5208 VPWR.n265 VPWR.n264 9.0005
R5209 VPWR.n9082 VPWR.n9081 9.0005
R5210 VPWR.n6794 VPWR.n6793 9.0005
R5211 VPWR.n6801 VPWR.n6800 9.0005
R5212 VPWR.n6822 VPWR.n6821 9.0005
R5213 VPWR.n6813 VPWR.n6812 9.0005
R5214 VPWR.n8246 VPWR.n8245 9.0005
R5215 VPWR.n8835 VPWR.n8834 9.0005
R5216 VPWR.n8841 VPWR.n8840 9.0005
R5217 VPWR.n8853 VPWR.n8852 9.0005
R5218 VPWR.n8928 VPWR.n8927 9.0005
R5219 VPWR.n6467 VPWR.n6466 9.0005
R5220 VPWR.n6474 VPWR.n6473 9.0005
R5221 VPWR.n6559 VPWR.n6558 9.0005
R5222 VPWR.n6562 VPWR.n6561 9.0005
R5223 VPWR.n8557 VPWR.n8556 9.0005
R5224 VPWR.n8534 VPWR.n8533 9.0005
R5225 VPWR.n8717 VPWR.n8716 9.0005
R5226 VPWR.n8798 VPWR.n8797 9.0005
R5227 VPWR.n5746 VPWR.n5745 9.0005
R5228 VPWR.n5752 VPWR.n5751 9.0005
R5229 VPWR.n5838 VPWR.n5837 9.0005
R5230 VPWR.n662 VPWR.n661 9.0005
R5231 VPWR.n695 VPWR.n694 9.0005
R5232 VPWR.n1366 VPWR.n1365 9.0005
R5233 VPWR.n1349 VPWR.n1348 9.0005
R5234 VPWR.n1359 VPWR.n1358 9.0005
R5235 VPWR.n5504 VPWR.n5503 9.0005
R5236 VPWR.n5498 VPWR.n5497 9.0005
R5237 VPWR.n5669 VPWR.n5668 9.0005
R5238 VPWR.n5675 VPWR.n5674 9.0005
R5239 VPWR.n5687 VPWR.n5686 9.0005
R5240 VPWR.n5695 VPWR.n5694 9.0005
R5241 VPWR.n5572 VPWR.n5571 9.0005
R5242 VPWR.n1340 VPWR.n1339 9.0005
R5243 VPWR.n1421 VPWR.n1420 9.0005
R5244 VPWR.n1397 VPWR.n1396 9.0005
R5245 VPWR.n1391 VPWR.n1390 9.0005
R5246 VPWR.n1641 VPWR.n1640 9.0005
R5247 VPWR.n1594 VPWR.n1593 9.0005
R5248 VPWR.n1634 VPWR.n1633 9.0005
R5249 VPWR.n1796 VPWR.n1795 9.0005
R5250 VPWR.n4651 VPWR.n4650 9.0005
R5251 VPWR.n4856 VPWR.n4855 9.0005
R5252 VPWR.n1605 VPWR.n1604 9.0005
R5253 VPWR.n1741 VPWR.n1740 9.0005
R5254 VPWR.n1735 VPWR.n1734 9.0005
R5255 VPWR.n2545 VPWR.n2544 9.0005
R5256 VPWR.n5076 VPWR.n5075 9.0005
R5257 VPWR.n5070 VPWR.n5069 9.0005
R5258 VPWR VPWR.n1886 9.0005
R5259 VPWR.n5038 VPWR.n5037 9.0005
R5260 VPWR.n2538 VPWR.n2537 9.0005
R5261 VPWR.n2492 VPWR.n2491 9.0005
R5262 VPWR.n2526 VPWR.n2525 9.0005
R5263 VPWR.n2583 VPWR.n2582 9.0005
R5264 VPWR.n4396 VPWR.n4395 9.0005
R5265 VPWR.n4548 VPWR.n4547 9.0005
R5266 VPWR.n4372 VPWR.n4371 9.0005
R5267 VPWR.n4380 VPWR.n4379 9.0005
R5268 VPWR.n2675 VPWR.n2673 9.0005
R5269 VPWR.n2675 VPWR.n2674 9.0005
R5270 VPWR.n2654 VPWR.n2653 9.0005
R5271 VPWR.n2648 VPWR.n2647 9.0005
R5272 VPWR.n3494 VPWR.n3493 9.0005
R5273 VPWR.n4230 VPWR.n4229 9.0005
R5274 VPWR.n4224 VPWR.n4223 9.0005
R5275 VPWR.n2943 VPWR.n2942 9.0005
R5276 VPWR.n4270 VPWR.n4269 9.0005
R5277 VPWR.n4293 VPWR.n4292 9.0005
R5278 VPWR.n4287 VPWR.n4286 9.0005
R5279 VPWR.n3488 VPWR.n3487 9.0005
R5280 VPWR.n3453 VPWR.n3452 9.0005
R5281 VPWR.n3462 VPWR.n3461 9.0005
R5282 VPWR.n3547 VPWR.n3546 9.0005
R5283 VPWR.n7823 VPWR.n7822 9.0005
R5284 VPWR.n7840 VPWR.n7839 9.0005
R5285 VPWR.n7846 VPWR.n7845 9.0005
R5286 VPWR.n9211 VPWR.n9210 9.0005
R5287 VPWR VPWR.n9218 9.0005
R5288 VPWR.n129 VPWR.n128 9.0005
R5289 VPWR.n120 VPWR.n119 9.0005
R5290 VPWR.n6131 VPWR.n6130 9.0005
R5291 VPWR.n7693 VPWR.n7692 9.0005
R5292 VPWR.n7713 VPWR.n7712 9.0005
R5293 VPWR.n3864 VPWR.n3863 9.0005
R5294 VPWR.n3846 VPWR.n3845 9.0005
R5295 VPWR.n3840 VPWR.n3839 9.0005
R5296 VPWR.n3983 VPWR.n3982 9.0005
R5297 VPWR.n3964 VPWR.n3963 9.0005
R5298 VPWR.n3327 VPWR.n3326 9.0005
R5299 VPWR.n3321 VPWR.n3320 9.0005
R5300 VPWR.n3310 VPWR.n3309 9.0005
R5301 VPWR.n3301 VPWR.n3300 9.0005
R5302 VPWR.n4168 VPWR.n4167 9.0005
R5303 VPWR.n4162 VPWR.n4161 9.0005
R5304 VPWR.n4152 VPWR.n4151 9.0005
R5305 VPWR.n4143 VPWR.n4142 9.0005
R5306 VPWR.n7132 VPWR.n7131 9.0005
R5307 VPWR.n7448 VPWR.n7447 9.0005
R5308 VPWR.n7608 VPWR.n7607 9.0005
R5309 VPWR.n7602 VPWR.n7601 9.0005
R5310 VPWR.n7582 VPWR.n7581 9.0005
R5311 VPWR.n7591 VPWR.n7590 9.0005
R5312 VPWR.n7432 VPWR.n7431 9.0005
R5313 VPWR.n7426 VPWR.n7425 9.0005
R5314 VPWR.n7211 VPWR.n7210 9.0005
R5315 VPWR.n7200 VPWR.n7199 9.0005
R5316 VPWR.n7221 VPWR.n7220 9.0005
R5317 VPWR.n5964 VPWR.n5963 8.88645
R5318 VPWR.n6356 VPWR.n6355 8.88645
R5319 VPWR.n3509 VPWR.n3508 8.88645
R5320 VPWR.n4727 VPWR.n4726 8.77764
R5321 VPWR.n1930 VPWR.n1929 8.65932
R5322 VPWR.n2531 VPWR.n2530 8.65932
R5323 VPWR.n4936 VPWR.n4920 8.62646
R5324 VPWR.n2059 VPWR.n2044 8.62646
R5325 VPWR.n7811 VPWR.n7809 8.49383
R5326 VPWR.n6636 VPWR.n6634 8.49383
R5327 VPWR.n4491 VPWR.n4490 8.46331
R5328 VPWR.n3185 VPWR.n3184 8.44958
R5329 VPWR.n7752 VPWR.n6128 8.44958
R5330 VPWR.n7809 VPWR.n6114 8.44958
R5331 VPWR.n6036 VPWR.n6034 8.44958
R5332 VPWR.n8011 VPWR.n5968 8.44958
R5333 VPWR.n6298 VPWR.n6297 8.44958
R5334 VPWR.n6766 VPWR.n6765 8.44958
R5335 VPWR.n1704 VPWR.n1702 8.44958
R5336 VPWR.n536 VPWR.n535 8.41193
R5337 VPWR.n2074 VPWR.n2073 8.41193
R5338 VPWR.t2737 VPWR.t187 8.39273
R5339 VPWR.t3178 VPWR.t3073 8.39273
R5340 VPWR.t795 VPWR.t3001 8.39273
R5341 VPWR.t2715 VPWR.t276 8.39273
R5342 VPWR.t1856 VPWR.t784 8.39273
R5343 VPWR.t48 VPWR.t2937 8.39273
R5344 VPWR.t2001 VPWR.t3054 8.39273
R5345 VPWR.t1829 VPWR.t3233 8.39273
R5346 VPWR.t2341 VPWR.t688 8.39273
R5347 VPWR.t3225 VPWR.t2095 8.39273
R5348 VPWR.t762 VPWR 8.39273
R5349 VPWR.t1101 VPWR.t2003 8.39273
R5350 VPWR.t1057 VPWR.t772 8.39273
R5351 VPWR.t2618 VPWR.t1031 8.39273
R5352 VPWR.t2278 VPWR.t1215 8.39273
R5353 VPWR.t1526 VPWR.t178 8.39273
R5354 VPWR.t2931 VPWR.t2761 8.39273
R5355 VPWR.t2603 VPWR.t3278 8.39273
R5356 VPWR.t2228 VPWR.t2940 8.39273
R5357 VPWR.t1497 VPWR.t612 8.39273
R5358 VPWR.t3174 VPWR 8.39273
R5359 VPWR.n6346 VPWR.n6344 8.28285
R5360 VPWR.n4053 VPWR.n4052 8.23801
R5361 VPWR.n3870 VPWR.n3869 8.04017
R5362 VPWR.n4028 VPWR.n2997 8.01134
R5363 VPWR.n4739 VPWR.n4738 7.97427
R5364 VPWR.n8887 VPWR.n8873 7.90638
R5365 VPWR.n5797 VPWR.n5783 7.90638
R5366 VPWR.n411 VPWR.n409 7.90638
R5367 VPWR.n3918 VPWR.n3917 7.87742
R5368 VPWR.n6758 VPWR.n6755 7.87742
R5369 VPWR.n4128 VPWR.n4127 7.81487
R5370 VPWR.n3088 VPWR.n3048 7.75995
R5371 VPWR.n9051 VPWR.n9050 7.75995
R5372 VPWR.n8468 VPWR.n8466 7.75995
R5373 VPWR.n6445 VPWR.n6422 7.75995
R5374 VPWR.n5629 VPWR.n5627 7.75995
R5375 VPWR.n5485 VPWR.n491 7.75995
R5376 VPWR.n4836 VPWR.n4835 7.75995
R5377 VPWR.n2720 VPWR.n2718 7.75995
R5378 VPWR.n4519 VPWR.n4518 7.75995
R5379 VPWR.n2819 VPWR.n2818 7.75995
R5380 VPWR.n627 VPWR.n625 7.71815
R5381 VPWR.n1310 VPWR.n1309 7.61703
R5382 VPWR.n4417 VPWR.n4416 7.58569
R5383 VPWR.n3680 VPWR.n3679 7.52991
R5384 VPWR.n8500 VPWR.n8498 7.4432
R5385 VPWR.n8439 VPWR.n8438 7.28326
R5386 VPWR.n3911 VPWR.n3909 7.25383
R5387 VPWR.n7765 VPWR.n7764 7.25383
R5388 VPWR.n6237 VPWR.n6232 7.25383
R5389 VPWR.n6752 VPWR.n6750 7.25383
R5390 VPWR.n7784 VPWR.n7782 7.21067
R5391 VPWR.n6030 VPWR.n6027 7.21067
R5392 VPWR.n6083 VPWR.n6082 7.15344
R5393 VPWR.n7917 VPWR.n7916 7.15344
R5394 VPWR.n8768 VPWR.n8767 7.15344
R5395 VPWR.n8650 VPWR.n8649 7.15344
R5396 VPWR.n1033 VPWR.n1032 7.15344
R5397 VPWR.n1429 VPWR.n1428 7.15344
R5398 VPWR.n1932 VPWR.n1931 7.15344
R5399 VPWR.n2149 VPWR.n2148 7.15344
R5400 VPWR.n8486 VPWR.n8485 7.12524
R5401 VPWR.n7037 VPWR.n7036 7.11866
R5402 VPWR.n3916 VPWR.n3915 7.11866
R5403 VPWR.n6754 VPWR.n6753 7.11866
R5404 VPWR.n8506 VPWR.n8505 7.11866
R5405 VPWR.n7269 VPWR.n7268 7.11866
R5406 VPWR.n2075 VPWR.n2074 6.94907
R5407 VPWR.n7992 VPWR.n7991 6.93383
R5408 VPWR.n4069 VPWR.n4068 6.77697
R5409 VPWR.n5490 VPWR.n5489 6.77075
R5410 VPWR.n3639 VPWR.n3638 6.77075
R5411 VPWR.t2104 VPWR.t1882 6.71428
R5412 VPWR.t2087 VPWR.t897 6.71428
R5413 VPWR.t2085 VPWR.t2791 6.71428
R5414 VPWR.t2999 VPWR.t1691 6.71428
R5415 VPWR.t1952 VPWR.t1219 6.71428
R5416 VPWR.t3186 VPWR.t655 6.71428
R5417 VPWR.t1908 VPWR.t1938 6.71428
R5418 VPWR.t1515 VPWR.t1910 6.71428
R5419 VPWR.t1769 VPWR.t3263 6.71428
R5420 VPWR.t2405 VPWR.t2252 6.71428
R5421 VPWR.t2148 VPWR.t2174 6.71428
R5422 VPWR.t855 VPWR.t1033 6.71428
R5423 VPWR.t1337 VPWR.t2261 6.71428
R5424 VPWR.t1926 VPWR.t1619 6.71428
R5425 VPWR.t2101 VPWR.t1344 6.71428
R5426 VPWR.t2883 VPWR.t2016 6.71428
R5427 VPWR.t54 VPWR.t1924 6.71428
R5428 VPWR.n8431 VPWR.n5866 6.67717
R5429 VPWR.n3888 VPWR.n3886 6.66496
R5430 VPWR.n3904 VPWR.n3903 6.66496
R5431 VPWR.n7673 VPWR.n7637 6.66496
R5432 VPWR.n7757 VPWR.n7756 6.66496
R5433 VPWR.n6044 VPWR.n6014 6.66496
R5434 VPWR.n6045 VPWR.n6044 6.66496
R5435 VPWR.n8011 VPWR.n5969 6.66496
R5436 VPWR.n6265 VPWR.n6264 6.66496
R5437 VPWR.n6288 VPWR.n6287 6.66496
R5438 VPWR.n6297 VPWR.n6228 6.66496
R5439 VPWR.n6644 VPWR.n6643 6.66496
R5440 VPWR.n452 VPWR.n451 6.66496
R5441 VPWR.n5494 VPWR.n486 6.66496
R5442 VPWR.n4408 VPWR.n4407 6.66496
R5443 VPWR.n3635 VPWR.n3634 6.66496
R5444 VPWR.n7816 VPWR.n7815 6.59529
R5445 VPWR.n1185 VPWR.n1184 6.58336
R5446 VPWR.n1151 VPWR.n1148 6.58336
R5447 VPWR.n4640 VPWR.n4639 6.49462
R5448 VPWR.n3909 VPWR.n3908 6.48583
R5449 VPWR.n7766 VPWR.n7765 6.48583
R5450 VPWR.n6263 VPWR.n6232 6.48583
R5451 VPWR.n6750 VPWR.n6645 6.48583
R5452 VPWR.n5637 VPWR.n5636 6.41151
R5453 VPWR.n2549 VPWR.n2548 6.4005
R5454 VPWR.n8898 VPWR.n8896 6.18775
R5455 VPWR.n449 VPWR.n448 6.03025
R5456 VPWR.n5579 VPWR.n5578 6.03025
R5457 VPWR.n4278 VPWR.n4277 6.03025
R5458 VPWR.n95 VPWR.n93 6.02403
R5459 VPWR.n244 VPWR.n242 6.02403
R5460 VPWR.n7916 VPWR.n7915 6.02403
R5461 VPWR.n936 VPWR.n935 6.02403
R5462 VPWR.n2696 VPWR.n2695 5.96824
R5463 VPWR.n1304 VPWR.n1303 5.85939
R5464 VPWR.n4114 VPWR.n4113 5.85546
R5465 VPWR.n4708 VPWR.n4707 5.85193
R5466 VPWR.n4726 VPWR.n4724 5.85193
R5467 VPWR.n2728 VPWR.n2727 5.50133
R5468 VPWR.n4015 VPWR.n4010 5.48841
R5469 VPWR.n4033 VPWR.n4029 5.42606
R5470 VPWR.n4076 VPWR.n4074 5.42606
R5471 VPWR.n5870 VPWR.n5869 5.40233
R5472 VPWR.n1440 VPWR.n1383 5.40233
R5473 VPWR.n1679 VPWR.n1678 5.40233
R5474 VPWR.n2128 VPWR.n2126 5.40233
R5475 VPWR.n8456 VPWR.n8455 5.39479
R5476 VPWR.n3034 VPWR.n3032 5.31652
R5477 VPWR.n6292 VPWR.n6291 5.31652
R5478 VPWR.n3151 VPWR.n3150 5.29281
R5479 VPWR.n4032 VPWR.n4031 5.29281
R5480 VPWR.n6121 VPWR.n6120 5.29281
R5481 VPWR.n6118 VPWR.n6117 5.29281
R5482 VPWR.n6116 VPWR.n6115 5.29281
R5483 VPWR.n6113 VPWR.n6112 5.29281
R5484 VPWR.n6009 VPWR.n6008 5.29281
R5485 VPWR.n6029 VPWR.n6028 5.29281
R5486 VPWR.n5967 VPWR.n5966 5.29281
R5487 VPWR.n1686 VPWR.n1685 5.29281
R5488 VPWR.n2888 VPWR.n2887 5.29281
R5489 VPWR.n4007 VPWR.n4006 5.28746
R5490 VPWR.n5141 VPWR.n1837 5.28746
R5491 VPWR.n722 VPWR.n721 5.27109
R5492 VPWR.n5423 VPWR.n5422 5.27109
R5493 VPWR.n4767 VPWR.n4645 5.25888
R5494 VPWR.n6036 VPWR.n6035 5.18397
R5495 VPWR.n6282 VPWR.n6281 5.18397
R5496 VPWR.n6416 VPWR.n6415 5.18397
R5497 VPWR.n5622 VPWR.n5621 5.18397
R5498 VPWR.n5513 VPWR.n5512 5.18397
R5499 VPWR.n1316 VPWR.n1272 5.18397
R5500 VPWR.n4790 VPWR.n4789 5.18397
R5501 VPWR.n4363 VPWR.n4362 5.18397
R5502 VPWR.n2787 VPWR.n2786 5.18397
R5503 VPWR.n1836 VPWR.n1834 5.05749
R5504 VPWR.t1155 VPWR.t1998 5.03584
R5505 VPWR.t1113 VPWR.t181 5.03584
R5506 VPWR.t3109 VPWR.t1171 5.03584
R5507 VPWR.t3321 VPWR.t2042 5.03584
R5508 VPWR.t1002 VPWR.t879 5.03584
R5509 VPWR.t1055 VPWR.t3017 5.03584
R5510 VPWR.t3015 VPWR.t1845 5.03584
R5511 VPWR.t1413 VPWR.t2116 5.03584
R5512 VPWR.t2276 VPWR.t1213 5.03584
R5513 VPWR.t1986 VPWR.t1121 5.03584
R5514 VPWR.t2944 VPWR.t2929 5.03584
R5515 VPWR.t3036 VPWR.t1567 5.03584
R5516 VPWR.t1075 VPWR.t264 5.03584
R5517 VPWR.t1907 VPWR.t355 5.03584
R5518 VPWR.n3202 VPWR.n3201 5.03171
R5519 VPWR.n1684 VPWR.n1683 5.03171
R5520 VPWR VPWR.n7531 4.9774
R5521 VPWR.n7666 VPWR.n7665 4.9724
R5522 VPWR.n8978 VPWR.n8977 4.9724
R5523 VPWR.n4234 VPWR.n4233 4.9724
R5524 VPWR.n3037 VPWR.n3036 4.93613
R5525 VPWR.n4642 VPWR.n4641 4.91363
R5526 VPWR.n947 VPWR.n762 4.91172
R5527 VPWR.n2085 VPWR.n2084 4.91172
R5528 VPWR.n9187 VPWR.n9186 4.89462
R5529 VPWR.n8291 VPWR.n8290 4.89462
R5530 VPWR.n1217 VPWR.n1214 4.89462
R5531 VPWR.n4680 VPWR.n4679 4.89462
R5532 VPWR.n2245 VPWR.n2244 4.89462
R5533 VPWR.n2664 VPWR.n2663 4.89462
R5534 VPWR.n6394 VPWR.n6393 4.86662
R5535 VPWR.n4009 VPWR.n4008 4.8005
R5536 VPWR.n1680 VPWR.n1679 4.76083
R5537 VPWR.n1151 VPWR.n1150 4.75479
R5538 VPWR.n934 VPWR.n932 4.72311
R5539 VPWR.n4773 VPWR.n4771 4.69218
R5540 VPWR.n6947 VPWR.n6946 4.67352
R5541 VPWR.n7292 VPWR.n7291 4.67352
R5542 VPWR.n3078 VPWR.n3050 4.67352
R5543 VPWR.n4108 VPWR.n4107 4.67352
R5544 VPWR.n3239 VPWR.n3238 4.67352
R5545 VPWR.n9140 VPWR.n61 4.67352
R5546 VPWR.n56 VPWR.n55 4.67352
R5547 VPWR.n46 VPWR.n45 4.67352
R5548 VPWR.n39 VPWR.n38 4.67352
R5549 VPWR.n9200 VPWR.n32 4.67352
R5550 VPWR.n9196 VPWR.n32 4.67352
R5551 VPWR.n209 VPWR.n208 4.67352
R5552 VPWR.n5927 VPWR.n5926 4.67352
R5553 VPWR.n5941 VPWR.n5940 4.67352
R5554 VPWR.n8194 VPWR.n8193 4.67352
R5555 VPWR.n8754 VPWR.n8753 4.67352
R5556 VPWR.n8628 VPWR.n8627 4.67352
R5557 VPWR.n8442 VPWR.n8441 4.67352
R5558 VPWR.n6509 VPWR.n6508 4.67352
R5559 VPWR.n1133 VPWR.n1130 4.67352
R5560 VPWR.n1125 VPWR.n1124 4.67352
R5561 VPWR.n752 VPWR.n751 4.67352
R5562 VPWR.n810 VPWR.n809 4.67352
R5563 VPWR.n5463 VPWR.n5460 4.67352
R5564 VPWR.n5441 VPWR.n5440 4.67352
R5565 VPWR.n5443 VPWR.n5441 4.67352
R5566 VPWR.n1298 VPWR.n1294 4.67352
R5567 VPWR.n1296 VPWR.n1295 4.67352
R5568 VPWR.n1721 VPWR.n551 4.67352
R5569 VPWR.n1722 VPWR.n1721 4.67352
R5570 VPWR.n1723 VPWR.n1722 4.67352
R5571 VPWR.n4917 VPWR.n4916 4.67352
R5572 VPWR.n5013 VPWR.n5012 4.67352
R5573 VPWR.n5012 VPWR.n1959 4.67352
R5574 VPWR.n1962 VPWR.n1959 4.67352
R5575 VPWR.n5135 VPWR.n5134 4.67352
R5576 VPWR.n2131 VPWR.n2129 4.67352
R5577 VPWR.n2562 VPWR.n2561 4.67352
R5578 VPWR.n2461 VPWR.n2459 4.67352
R5579 VPWR.n2469 VPWR.n2468 4.67352
R5580 VPWR.n2376 VPWR.n2375 4.67352
R5581 VPWR.n2375 VPWR.n2374 4.67352
R5582 VPWR.n2002 VPWR.n2001 4.67352
R5583 VPWR.n3582 VPWR.n3581 4.67352
R5584 VPWR.n3503 VPWR.n3502 4.67352
R5585 VPWR.n3629 VPWR.n3628 4.67352
R5586 VPWR.n7072 VPWR.n7071 4.67352
R5587 VPWR.n950 VPWR.n949 4.65505
R5588 VPWR.n1507 VPWR.n1506 4.65505
R5589 VPWR.n6311 VPWR.n6225 4.6505
R5590 VPWR.n6178 VPWR.n6177 4.6505
R5591 VPWR.n6181 VPWR.n6180 4.6505
R5592 VPWR.n6183 VPWR.n6182 4.6505
R5593 VPWR.n6184 VPWR.n6158 4.6505
R5594 VPWR.n6310 VPWR.n6309 4.6505
R5595 VPWR.n6308 VPWR.n6307 4.6505
R5596 VPWR.n6306 VPWR.n6305 4.6505
R5597 VPWR.n6303 VPWR.n6302 4.6505
R5598 VPWR.n6301 VPWR.n6300 4.6505
R5599 VPWR.n6299 VPWR.n6298 4.6505
R5600 VPWR.n6297 VPWR.n6296 4.6505
R5601 VPWR.n6294 VPWR.n6293 4.6505
R5602 VPWR.n6283 VPWR.n6282 4.6505
R5603 VPWR.n6280 VPWR.n6279 4.6505
R5604 VPWR.n6278 VPWR.n6277 4.6505
R5605 VPWR.n6273 VPWR.n6272 4.6505
R5606 VPWR.n6269 VPWR.n6268 4.6505
R5607 VPWR.n6260 VPWR.n6259 4.6505
R5608 VPWR.n6253 VPWR.n6252 4.6505
R5609 VPWR.n6251 VPWR.n6250 4.6505
R5610 VPWR.n6249 VPWR.n6248 4.6505
R5611 VPWR.n6247 VPWR.n6246 4.6505
R5612 VPWR.n6244 VPWR.n6243 4.6505
R5613 VPWR.n6241 VPWR.n5968 4.6505
R5614 VPWR.n8011 VPWR.n8010 4.6505
R5615 VPWR.n8058 VPWR.n8057 4.6505
R5616 VPWR.n8054 VPWR.n8053 4.6505
R5617 VPWR.n8049 VPWR.n8047 4.6505
R5618 VPWR.n8014 VPWR.n5965 4.6505
R5619 VPWR.n7911 VPWR.n7908 4.6505
R5620 VPWR.n7912 VPWR.n7906 4.6505
R5621 VPWR.n7919 VPWR.n7904 4.6505
R5622 VPWR.n7952 VPWR.n7951 4.6505
R5623 VPWR.n8018 VPWR.n8017 4.6505
R5624 VPWR.n8020 VPWR.n8019 4.6505
R5625 VPWR.n8024 VPWR.n8023 4.6505
R5626 VPWR.n8026 VPWR.n8025 4.6505
R5627 VPWR.n8029 VPWR.n8028 4.6505
R5628 VPWR.n8031 VPWR.n8030 4.6505
R5629 VPWR.n8033 VPWR.n8032 4.6505
R5630 VPWR.n8036 VPWR.n8035 4.6505
R5631 VPWR.n8038 VPWR.n8037 4.6505
R5632 VPWR.n8040 VPWR.n8039 4.6505
R5633 VPWR.n8042 VPWR.n8041 4.6505
R5634 VPWR.n8044 VPWR.n8043 4.6505
R5635 VPWR.n9050 VPWR.n194 4.6505
R5636 VPWR.n9047 VPWR.n8974 4.6505
R5637 VPWR.n8972 VPWR.n198 4.6505
R5638 VPWR.n8971 VPWR.n198 4.6505
R5639 VPWR.n255 VPWR.n207 4.6505
R5640 VPWR.n230 VPWR.n229 4.6505
R5641 VPWR.n228 VPWR.n214 4.6505
R5642 VPWR.n225 VPWR.n216 4.6505
R5643 VPWR.n254 VPWR.n253 4.6505
R5644 VPWR.n252 VPWR.n251 4.6505
R5645 VPWR.n249 VPWR.n248 4.6505
R5646 VPWR.n246 VPWR.n245 4.6505
R5647 VPWR.n242 VPWR.n241 4.6505
R5648 VPWR.n240 VPWR.n211 4.6505
R5649 VPWR.n237 VPWR.n236 4.6505
R5650 VPWR.n234 VPWR.n233 4.6505
R5651 VPWR.n232 VPWR.n231 4.6505
R5652 VPWR.n227 VPWR.n226 4.6505
R5653 VPWR.n9065 VPWR.n9064 4.6505
R5654 VPWR.n9059 VPWR.n9058 4.6505
R5655 VPWR.n9056 VPWR.n9055 4.6505
R5656 VPWR.n9054 VPWR.n9053 4.6505
R5657 VPWR.n9052 VPWR.n9051 4.6505
R5658 VPWR.n8980 VPWR.n196 4.6505
R5659 VPWR.n8982 VPWR.n8981 4.6505
R5660 VPWR.n8984 VPWR.n8983 4.6505
R5661 VPWR.n8988 VPWR.n8987 4.6505
R5662 VPWR.n8992 VPWR.n8991 4.6505
R5663 VPWR.n8994 VPWR.n8993 4.6505
R5664 VPWR.n8996 VPWR.n8995 4.6505
R5665 VPWR.n8999 VPWR.n8998 4.6505
R5666 VPWR.n9002 VPWR.n9001 4.6505
R5667 VPWR.n9004 VPWR.n9003 4.6505
R5668 VPWR.n9008 VPWR.n9007 4.6505
R5669 VPWR.n9010 VPWR.n9009 4.6505
R5670 VPWR.n9012 VPWR.n9011 4.6505
R5671 VPWR.n9014 VPWR.n9013 4.6505
R5672 VPWR.n9017 VPWR.n9016 4.6505
R5673 VPWR.n9021 VPWR.n9020 4.6505
R5674 VPWR.n9023 VPWR.n9022 4.6505
R5675 VPWR.n9025 VPWR.n9024 4.6505
R5676 VPWR.n9027 VPWR.n9026 4.6505
R5677 VPWR.n9029 VPWR.n9028 4.6505
R5678 VPWR.n9031 VPWR.n9030 4.6505
R5679 VPWR.n9035 VPWR.n9034 4.6505
R5680 VPWR.n9037 VPWR.n9036 4.6505
R5681 VPWR.n9040 VPWR.n9039 4.6505
R5682 VPWR.n9042 VPWR.n9041 4.6505
R5683 VPWR.n9044 VPWR.n9043 4.6505
R5684 VPWR.n9046 VPWR.n9045 4.6505
R5685 VPWR.n8970 VPWR.n8969 4.6505
R5686 VPWR.n257 VPWR.n256 4.6505
R5687 VPWR.n8056 VPWR.n8055 4.6505
R5688 VPWR.n8051 VPWR.n8050 4.6505
R5689 VPWR.n8046 VPWR.n8045 4.6505
R5690 VPWR.n7910 VPWR.n7909 4.6505
R5691 VPWR.n7914 VPWR.n7913 4.6505
R5692 VPWR.n7918 VPWR.n7917 4.6505
R5693 VPWR.n7921 VPWR.n7920 4.6505
R5694 VPWR.n7923 VPWR.n7922 4.6505
R5695 VPWR.n7925 VPWR.n7924 4.6505
R5696 VPWR.n7929 VPWR.n7928 4.6505
R5697 VPWR.n7931 VPWR.n7930 4.6505
R5698 VPWR.n7934 VPWR.n7933 4.6505
R5699 VPWR.n7936 VPWR.n7935 4.6505
R5700 VPWR.n7938 VPWR.n7937 4.6505
R5701 VPWR.n7941 VPWR.n7940 4.6505
R5702 VPWR.n7945 VPWR.n7944 4.6505
R5703 VPWR.n7947 VPWR.n7946 4.6505
R5704 VPWR.n7950 VPWR.n7949 4.6505
R5705 VPWR.n7955 VPWR.n7954 4.6505
R5706 VPWR.n6266 VPWR.n6265 4.6505
R5707 VPWR.n6285 VPWR.n6284 4.6505
R5708 VPWR.n6287 VPWR.n6286 4.6505
R5709 VPWR.n6194 VPWR.n6193 4.6505
R5710 VPWR.n6199 VPWR.n6198 4.6505
R5711 VPWR.n6779 VPWR.n6640 4.6505
R5712 VPWR.n6694 VPWR.n6693 4.6505
R5713 VPWR.n6597 VPWR.n6588 4.6505
R5714 VPWR.n6603 VPWR.n6602 4.6505
R5715 VPWR.n6778 VPWR.n6777 4.6505
R5716 VPWR.n6776 VPWR.n6775 4.6505
R5717 VPWR.n6774 VPWR.n6773 4.6505
R5718 VPWR.n6771 VPWR.n6770 4.6505
R5719 VPWR.n6769 VPWR.n6768 4.6505
R5720 VPWR.n6767 VPWR.n6766 4.6505
R5721 VPWR.n6765 VPWR.n6764 4.6505
R5722 VPWR.n6761 VPWR.n6760 4.6505
R5723 VPWR.n6747 VPWR.n6746 4.6505
R5724 VPWR.n6745 VPWR.n6744 4.6505
R5725 VPWR.n6742 VPWR.n6741 4.6505
R5726 VPWR.n6727 VPWR.n6726 4.6505
R5727 VPWR.n6723 VPWR.n6722 4.6505
R5728 VPWR.n6697 VPWR.n6696 4.6505
R5729 VPWR.n8199 VPWR.n8109 4.6505
R5730 VPWR.n8187 VPWR.n8111 4.6505
R5731 VPWR.n8134 VPWR.n8133 4.6505
R5732 VPWR.n8136 VPWR.n8135 4.6505
R5733 VPWR.n8139 VPWR.n8138 4.6505
R5734 VPWR.n8143 VPWR.n8142 4.6505
R5735 VPWR.n8172 VPWR.n8171 4.6505
R5736 VPWR.n8174 VPWR.n8173 4.6505
R5737 VPWR.n8180 VPWR.n8179 4.6505
R5738 VPWR.n8893 VPWR.n8870 4.6505
R5739 VPWR.n8890 VPWR.n8871 4.6505
R5740 VPWR.n8887 VPWR.n8885 4.6505
R5741 VPWR.n8883 VPWR.n8874 4.6505
R5742 VPWR.n8914 VPWR.n8913 4.6505
R5743 VPWR.n8908 VPWR.n8907 4.6505
R5744 VPWR.n8906 VPWR.n8905 4.6505
R5745 VPWR.n8904 VPWR.n8903 4.6505
R5746 VPWR.n8900 VPWR.n8899 4.6505
R5747 VPWR.n8896 VPWR.n8895 4.6505
R5748 VPWR.n8894 VPWR.n8869 4.6505
R5749 VPWR.n8892 VPWR.n8891 4.6505
R5750 VPWR.n8889 VPWR.n8888 4.6505
R5751 VPWR.n8916 VPWR.n8915 4.6505
R5752 VPWR.n8198 VPWR.n8197 4.6505
R5753 VPWR.n8189 VPWR.n8188 4.6505
R5754 VPWR.n8128 VPWR.n8127 4.6505
R5755 VPWR.n8130 VPWR.n8129 4.6505
R5756 VPWR.n8132 VPWR.n8131 4.6505
R5757 VPWR.n8141 VPWR.n8140 4.6505
R5758 VPWR.n8153 VPWR.n8152 4.6505
R5759 VPWR.n8155 VPWR.n8154 4.6505
R5760 VPWR.n8158 VPWR.n8157 4.6505
R5761 VPWR.n8161 VPWR.n8160 4.6505
R5762 VPWR.n8163 VPWR.n8162 4.6505
R5763 VPWR.n8166 VPWR.n8123 4.6505
R5764 VPWR.n8168 VPWR.n8167 4.6505
R5765 VPWR.n8170 VPWR.n8169 4.6505
R5766 VPWR.n8176 VPWR.n8175 4.6505
R5767 VPWR.n8181 VPWR.n8117 4.6505
R5768 VPWR.n8184 VPWR.n8183 4.6505
R5769 VPWR.n8833 VPWR.n8832 4.6505
R5770 VPWR.n8342 VPWR.n8341 4.6505
R5771 VPWR.n8339 VPWR.n8338 4.6505
R5772 VPWR.n8335 VPWR.n8334 4.6505
R5773 VPWR.n8333 VPWR.n8332 4.6505
R5774 VPWR.n8331 VPWR.n8330 4.6505
R5775 VPWR.n8329 VPWR.n8328 4.6505
R5776 VPWR.n8326 VPWR.n8325 4.6505
R5777 VPWR.n8322 VPWR.n8321 4.6505
R5778 VPWR.n8318 VPWR.n8317 4.6505
R5779 VPWR.n8316 VPWR.n8315 4.6505
R5780 VPWR.n8314 VPWR.n5929 4.6505
R5781 VPWR.n8311 VPWR.n8310 4.6505
R5782 VPWR.n8309 VPWR.n8308 4.6505
R5783 VPWR.n8307 VPWR.n8306 4.6505
R5784 VPWR.n8304 VPWR.n8303 4.6505
R5785 VPWR.n8302 VPWR.n8301 4.6505
R5786 VPWR.n8300 VPWR.n8299 4.6505
R5787 VPWR.n8294 VPWR.n8293 4.6505
R5788 VPWR.n8292 VPWR.n8291 4.6505
R5789 VPWR.n8289 VPWR.n8288 4.6505
R5790 VPWR.n8287 VPWR.n5938 4.6505
R5791 VPWR.n8284 VPWR.n8283 4.6505
R5792 VPWR.n8282 VPWR.n8281 4.6505
R5793 VPWR.n8280 VPWR.n8279 4.6505
R5794 VPWR.n8278 VPWR.n8277 4.6505
R5795 VPWR.n8276 VPWR.n8275 4.6505
R5796 VPWR.n8274 VPWR.n8273 4.6505
R5797 VPWR.n8271 VPWR.n8270 4.6505
R5798 VPWR.n8268 VPWR.n8267 4.6505
R5799 VPWR.n8266 VPWR.n8265 4.6505
R5800 VPWR.n8264 VPWR.n8263 4.6505
R5801 VPWR.n8262 VPWR.n8261 4.6505
R5802 VPWR.n8260 VPWR.n8259 4.6505
R5803 VPWR.n8258 VPWR.n8257 4.6505
R5804 VPWR.n8256 VPWR.n8255 4.6505
R5805 VPWR.n6691 VPWR.n6657 4.6505
R5806 VPWR.n6699 VPWR.n6698 4.6505
R5807 VPWR.n6701 VPWR.n6700 4.6505
R5808 VPWR.n6703 VPWR.n6702 4.6505
R5809 VPWR.n6707 VPWR.n6706 4.6505
R5810 VPWR.n6709 VPWR.n6708 4.6505
R5811 VPWR.n6713 VPWR.n6712 4.6505
R5812 VPWR.n6716 VPWR.n6715 4.6505
R5813 VPWR.n6718 VPWR.n6717 4.6505
R5814 VPWR.n6720 VPWR.n6719 4.6505
R5815 VPWR.n6725 VPWR.n6724 4.6505
R5816 VPWR.n6729 VPWR.n6728 4.6505
R5817 VPWR.n6731 VPWR.n6730 4.6505
R5818 VPWR.n6735 VPWR.n6734 4.6505
R5819 VPWR.n6737 VPWR.n6736 4.6505
R5820 VPWR.n6739 VPWR.n6738 4.6505
R5821 VPWR.n6763 VPWR.n6643 4.6505
R5822 VPWR.n6599 VPWR.n6598 4.6505
R5823 VPWR.n6605 VPWR.n6604 4.6505
R5824 VPWR.n6609 VPWR.n6608 4.6505
R5825 VPWR.n6613 VPWR.n6612 4.6505
R5826 VPWR.n6614 VPWR.n6587 4.6505
R5827 VPWR.n6616 VPWR.n6615 4.6505
R5828 VPWR.n6619 VPWR.n6618 4.6505
R5829 VPWR.n6623 VPWR.n6622 4.6505
R5830 VPWR.n6625 VPWR.n6624 4.6505
R5831 VPWR.n6629 VPWR.n6628 4.6505
R5832 VPWR.n6631 VPWR.n6630 4.6505
R5833 VPWR.n6632 VPWR.n6586 4.6505
R5834 VPWR.n6634 VPWR.n6633 4.6505
R5835 VPWR.n6637 VPWR.n6636 4.6505
R5836 VPWR.n6639 VPWR.n6638 4.6505
R5837 VPWR.n6460 VPWR.n6346 4.6505
R5838 VPWR.n6455 VPWR.n6348 4.6505
R5839 VPWR.n6449 VPWR.n6350 4.6505
R5840 VPWR.n6446 VPWR.n6420 4.6505
R5841 VPWR.n6524 VPWR.n6523 4.6505
R5842 VPWR.n6529 VPWR.n6528 4.6505
R5843 VPWR.n6531 VPWR.n6530 4.6505
R5844 VPWR.n6368 VPWR.n6367 4.6505
R5845 VPWR.n6370 VPWR.n6369 4.6505
R5846 VPWR.n6373 VPWR.n6372 4.6505
R5847 VPWR.n6375 VPWR.n6374 4.6505
R5848 VPWR.n6382 VPWR.n6381 4.6505
R5849 VPWR.n6384 VPWR.n6383 4.6505
R5850 VPWR.n6386 VPWR.n6385 4.6505
R5851 VPWR.n6388 VPWR.n6387 4.6505
R5852 VPWR.n6391 VPWR.n6390 4.6505
R5853 VPWR.n6395 VPWR.n6394 4.6505
R5854 VPWR.n6397 VPWR.n6396 4.6505
R5855 VPWR.n6399 VPWR.n6398 4.6505
R5856 VPWR.n6401 VPWR.n6400 4.6505
R5857 VPWR.n6403 VPWR.n6402 4.6505
R5858 VPWR.n6405 VPWR.n6404 4.6505
R5859 VPWR.n6407 VPWR.n6406 4.6505
R5860 VPWR.n6409 VPWR.n6408 4.6505
R5861 VPWR.n6411 VPWR.n6410 4.6505
R5862 VPWR.n6413 VPWR.n6412 4.6505
R5863 VPWR.n6415 VPWR.n6414 4.6505
R5864 VPWR.n6418 VPWR.n6417 4.6505
R5865 VPWR.n6419 VPWR.n6351 4.6505
R5866 VPWR.n6445 VPWR.n6444 4.6505
R5867 VPWR.n6443 VPWR.n6422 4.6505
R5868 VPWR.n6442 VPWR.n6441 4.6505
R5869 VPWR.n8423 VPWR 4.6505
R5870 VPWR.n8424 VPWR.n5878 4.6505
R5871 VPWR.n8426 VPWR.n8425 4.6505
R5872 VPWR.n8491 VPWR.n8489 4.6505
R5873 VPWR.n8494 VPWR.n8493 4.6505
R5874 VPWR.n8605 VPWR.n8604 4.6505
R5875 VPWR.n8609 VPWR.n8608 4.6505
R5876 VPWR.n8676 VPWR.n8610 4.6505
R5877 VPWR.n8642 VPWR.n8621 4.6505
R5878 VPWR.n8641 VPWR.n8626 4.6505
R5879 VPWR.n8630 VPWR.n354 4.6505
R5880 VPWR.n8681 VPWR.n352 4.6505
R5881 VPWR.n8685 VPWR.n8684 4.6505
R5882 VPWR.n8760 VPWR.n8736 4.6505
R5883 VPWR.n8762 VPWR.n8761 4.6505
R5884 VPWR.n8785 VPWR.n8784 4.6505
R5885 VPWR.n8782 VPWR.n8781 4.6505
R5886 VPWR.n8780 VPWR.n8779 4.6505
R5887 VPWR.n8776 VPWR.n8775 4.6505
R5888 VPWR.n8774 VPWR.n8773 4.6505
R5889 VPWR.n8769 VPWR.n8768 4.6505
R5890 VPWR.n8749 VPWR.n8748 4.6505
R5891 VPWR.n8759 VPWR.n8758 4.6505
R5892 VPWR.n8764 VPWR.n8763 4.6505
R5893 VPWR.n8766 VPWR.n8765 4.6505
R5894 VPWR.n8770 VPWR.n8733 4.6505
R5895 VPWR.n8772 VPWR.n8771 4.6505
R5896 VPWR.n8788 VPWR.n8787 4.6505
R5897 VPWR.n8607 VPWR.n8606 4.6505
R5898 VPWR.n8671 VPWR.n8615 4.6505
R5899 VPWR.n8668 VPWR.n8667 4.6505
R5900 VPWR.n8665 VPWR.n8664 4.6505
R5901 VPWR.n8663 VPWR.n8662 4.6505
R5902 VPWR.n8659 VPWR.n8658 4.6505
R5903 VPWR.n8657 VPWR.n8656 4.6505
R5904 VPWR.n8655 VPWR.n8654 4.6505
R5905 VPWR.n8653 VPWR.n8652 4.6505
R5906 VPWR.n8651 VPWR.n8650 4.6505
R5907 VPWR.n8646 VPWR.n8645 4.6505
R5908 VPWR.n8644 VPWR.n8643 4.6505
R5909 VPWR.n8639 VPWR.n8638 4.6505
R5910 VPWR.n8634 VPWR.n8633 4.6505
R5911 VPWR.n8632 VPWR.n8631 4.6505
R5912 VPWR.n8680 VPWR.n8679 4.6505
R5913 VPWR.n8683 VPWR.n8682 4.6505
R5914 VPWR.n8688 VPWR.n8687 4.6505
R5915 VPWR.n8692 VPWR.n8691 4.6505
R5916 VPWR.n8600 VPWR.n8599 4.6505
R5917 VPWR.n8429 VPWR.n8428 4.6505
R5918 VPWR.n8434 VPWR.n8433 4.6505
R5919 VPWR.n8437 VPWR.n8436 4.6505
R5920 VPWR.n8446 VPWR.n8445 4.6505
R5921 VPWR.n8450 VPWR.n8449 4.6505
R5922 VPWR.n8460 VPWR.n8459 4.6505
R5923 VPWR.n8463 VPWR.n8462 4.6505
R5924 VPWR.n8464 VPWR.n5864 4.6505
R5925 VPWR.n8466 VPWR.n8465 4.6505
R5926 VPWR.n8469 VPWR.n8468 4.6505
R5927 VPWR.n8472 VPWR.n8471 4.6505
R5928 VPWR.n8475 VPWR.n8474 4.6505
R5929 VPWR.n8477 VPWR.n8476 4.6505
R5930 VPWR.n8479 VPWR.n8478 4.6505
R5931 VPWR.n8487 VPWR.n8486 4.6505
R5932 VPWR.n8488 VPWR.n5862 4.6505
R5933 VPWR.n8495 VPWR.n5861 4.6505
R5934 VPWR.n8497 VPWR.n8496 4.6505
R5935 VPWR.n8501 VPWR.n8500 4.6505
R5936 VPWR.n8504 VPWR.n8503 4.6505
R5937 VPWR.n8509 VPWR.n8508 4.6505
R5938 VPWR.n8512 VPWR.n8511 4.6505
R5939 VPWR.n8514 VPWR.n8513 4.6505
R5940 VPWR.n6365 VPWR.n6349 4.6505
R5941 VPWR.n6451 VPWR.n6450 4.6505
R5942 VPWR.n6457 VPWR.n6456 4.6505
R5943 VPWR.n6459 VPWR.n6458 4.6505
R5944 VPWR.n6503 VPWR.n6502 4.6505
R5945 VPWR.n6513 VPWR.n6512 4.6505
R5946 VPWR.n6515 VPWR.n6514 4.6505
R5947 VPWR.n6518 VPWR.n6517 4.6505
R5948 VPWR.n6521 VPWR.n6520 4.6505
R5949 VPWR.n6526 VPWR.n6525 4.6505
R5950 VPWR.n6532 VPWR.n6484 4.6505
R5951 VPWR.n6534 VPWR.n6533 4.6505
R5952 VPWR.n6543 VPWR.n6542 4.6505
R5953 VPWR.n1224 VPWR.n709 4.6505
R5954 VPWR.n1223 VPWR.n711 4.6505
R5955 VPWR.n1207 VPWR.n713 4.6505
R5956 VPWR.n858 VPWR.n857 4.6505
R5957 VPWR.n862 VPWR.n861 4.6505
R5958 VPWR.n864 VPWR.n714 4.6505
R5959 VPWR.n612 VPWR.n611 4.6505
R5960 VPWR.n621 VPWR.n620 4.6505
R5961 VPWR.n637 VPWR.n593 4.6505
R5962 VPWR.n1218 VPWR.n1217 4.6505
R5963 VPWR.n1212 VPWR.n1211 4.6505
R5964 VPWR.n829 VPWR.n828 4.6505
R5965 VPWR.n831 VPWR.n830 4.6505
R5966 VPWR.n833 VPWR.n832 4.6505
R5967 VPWR.n838 VPWR.n837 4.6505
R5968 VPWR.n845 VPWR.n844 4.6505
R5969 VPWR.n867 VPWR.n866 4.6505
R5970 VPWR.n871 VPWR.n870 4.6505
R5971 VPWR.n984 VPWR.n983 4.6505
R5972 VPWR.n987 VPWR.n986 4.6505
R5973 VPWR.n991 VPWR.n716 4.6505
R5974 VPWR.n1007 VPWR.n1006 4.6505
R5975 VPWR.n1011 VPWR.n1010 4.6505
R5976 VPWR.n1114 VPWR.n1113 4.6505
R5977 VPWR.n1120 VPWR.n1119 4.6505
R5978 VPWR.n1137 VPWR.n1136 4.6505
R5979 VPWR.n1139 VPWR.n1138 4.6505
R5980 VPWR.n1164 VPWR.n1163 4.6505
R5981 VPWR.n1175 VPWR.n1174 4.6505
R5982 VPWR.n1177 VPWR.n1176 4.6505
R5983 VPWR.n1180 VPWR.n1179 4.6505
R5984 VPWR.n1192 VPWR.n1191 4.6505
R5985 VPWR.n1194 VPWR.n722 4.6505
R5986 VPWR.n1199 VPWR.n719 4.6505
R5987 VPWR.n5794 VPWR.n5785 4.6505
R5988 VPWR.n5797 VPWR.n5796 4.6505
R5989 VPWR.n5800 VPWR.n5781 4.6505
R5990 VPWR.n5804 VPWR.n5803 4.6505
R5991 VPWR.n5822 VPWR.n5779 4.6505
R5992 VPWR.n5799 VPWR.n5798 4.6505
R5993 VPWR.n5802 VPWR.n5801 4.6505
R5994 VPWR.n5806 VPWR.n5805 4.6505
R5995 VPWR.n5808 VPWR.n5807 4.6505
R5996 VPWR.n5814 VPWR.n5813 4.6505
R5997 VPWR.n5816 VPWR.n5815 4.6505
R5998 VPWR.n5819 VPWR.n5818 4.6505
R5999 VPWR.n5821 VPWR.n5820 4.6505
R6000 VPWR.n5824 VPWR.n5823 4.6505
R6001 VPWR.n5826 VPWR.n5825 4.6505
R6002 VPWR.n5828 VPWR.n5827 4.6505
R6003 VPWR.n1112 VPWR.n1111 4.6505
R6004 VPWR.n1116 VPWR.n717 4.6505
R6005 VPWR.n1128 VPWR.n1127 4.6505
R6006 VPWR.n1130 VPWR.n1129 4.6505
R6007 VPWR.n1134 VPWR.n1133 4.6505
R6008 VPWR.n1144 VPWR.n1143 4.6505
R6009 VPWR.n1146 VPWR.n1145 4.6505
R6010 VPWR.n1152 VPWR.n1151 4.6505
R6011 VPWR.n1154 VPWR.n1153 4.6505
R6012 VPWR.n1158 VPWR.n1157 4.6505
R6013 VPWR.n1160 VPWR.n1159 4.6505
R6014 VPWR.n1168 VPWR.n1167 4.6505
R6015 VPWR.n1172 VPWR.n1171 4.6505
R6016 VPWR.n1182 VPWR.n1181 4.6505
R6017 VPWR.n1187 VPWR.n1186 4.6505
R6018 VPWR.n1189 VPWR.n1188 4.6505
R6019 VPWR.n1201 VPWR.n1200 4.6505
R6020 VPWR.n1198 VPWR.n1197 4.6505
R6021 VPWR.n5744 VPWR.n5743 4.6505
R6022 VPWR.n939 VPWR.n938 4.6505
R6023 VPWR.n944 VPWR.n943 4.6505
R6024 VPWR.n946 VPWR.n945 4.6505
R6025 VPWR.n955 VPWR.n954 4.6505
R6026 VPWR.n959 VPWR.n958 4.6505
R6027 VPWR.n962 VPWR.n961 4.6505
R6028 VPWR.n965 VPWR.n964 4.6505
R6029 VPWR.n969 VPWR.n968 4.6505
R6030 VPWR.n974 VPWR.n973 4.6505
R6031 VPWR.n977 VPWR.n976 4.6505
R6032 VPWR.n981 VPWR.n980 4.6505
R6033 VPWR.n989 VPWR.n988 4.6505
R6034 VPWR.n994 VPWR.n993 4.6505
R6035 VPWR.n999 VPWR.n998 4.6505
R6036 VPWR.n1002 VPWR.n1001 4.6505
R6037 VPWR.n1004 VPWR.n1003 4.6505
R6038 VPWR.n1009 VPWR.n1008 4.6505
R6039 VPWR.n1013 VPWR.n1012 4.6505
R6040 VPWR.n1016 VPWR.n1015 4.6505
R6041 VPWR.n1020 VPWR.n1019 4.6505
R6042 VPWR.n1022 VPWR.n1021 4.6505
R6043 VPWR.n1027 VPWR.n1026 4.6505
R6044 VPWR.n1030 VPWR.n754 4.6505
R6045 VPWR.n1032 VPWR.n1031 4.6505
R6046 VPWR.n1036 VPWR.n1035 4.6505
R6047 VPWR.n1038 VPWR.n1037 4.6505
R6048 VPWR.n937 VPWR.n936 4.6505
R6049 VPWR.n865 VPWR.n800 4.6505
R6050 VPWR.n860 VPWR.n859 4.6505
R6051 VPWR.n856 VPWR.n855 4.6505
R6052 VPWR.n852 VPWR.n851 4.6505
R6053 VPWR.n849 VPWR.n848 4.6505
R6054 VPWR.n847 VPWR.n846 4.6505
R6055 VPWR.n840 VPWR.n839 4.6505
R6056 VPWR.n826 VPWR.n712 4.6505
R6057 VPWR.n1210 VPWR.n1209 4.6505
R6058 VPWR.n1220 VPWR.n1219 4.6505
R6059 VPWR.n1222 VPWR.n1221 4.6505
R6060 VPWR VPWR.n601 4.6505
R6061 VPWR.n614 VPWR.n613 4.6505
R6062 VPWR.n618 VPWR.n617 4.6505
R6063 VPWR.n623 VPWR.n622 4.6505
R6064 VPWR.n625 VPWR.n624 4.6505
R6065 VPWR.n632 VPWR.n631 4.6505
R6066 VPWR.n634 VPWR.n633 4.6505
R6067 VPWR.n636 VPWR.n635 4.6505
R6068 VPWR.n639 VPWR.n638 4.6505
R6069 VPWR.n643 VPWR.n642 4.6505
R6070 VPWR.n646 VPWR.n645 4.6505
R6071 VPWR.n1517 VPWR.n1371 4.6505
R6072 VPWR.n1457 VPWR.n1456 4.6505
R6073 VPWR.n1453 VPWR.n1380 4.6505
R6074 VPWR.n1452 VPWR.n1382 4.6505
R6075 VPWR.n1431 VPWR.n1389 4.6505
R6076 VPWR.n1508 VPWR.n1507 4.6505
R6077 VPWR.n1501 VPWR.n1500 4.6505
R6078 VPWR.n1499 VPWR.n1498 4.6505
R6079 VPWR.n1492 VPWR.n1491 4.6505
R6080 VPWR.n1449 VPWR.n1448 4.6505
R6081 VPWR.n1447 VPWR.n1446 4.6505
R6082 VPWR.n1442 VPWR.n1441 4.6505
R6083 VPWR.n1439 VPWR.n1438 4.6505
R6084 VPWR.n1434 VPWR.n1433 4.6505
R6085 VPWR.n5414 VPWR.n5413 4.6505
R6086 VPWR.n5430 VPWR.n5429 4.6505
R6087 VPWR.n5605 VPWR.n462 4.6505
R6088 VPWR.n421 VPWR.n412 4.6505
R6089 VPWR.n423 VPWR.n411 4.6505
R6090 VPWR.n441 VPWR.n403 4.6505
R6091 VPWR.n425 VPWR.n424 4.6505
R6092 VPWR.n428 VPWR.n427 4.6505
R6093 VPWR.n430 VPWR.n429 4.6505
R6094 VPWR.n432 VPWR.n431 4.6505
R6095 VPWR.n434 VPWR.n433 4.6505
R6096 VPWR.n440 VPWR.n439 4.6505
R6097 VPWR.n443 VPWR.n442 4.6505
R6098 VPWR.n447 VPWR.n446 4.6505
R6099 VPWR.n450 VPWR.n449 4.6505
R6100 VPWR.n5580 VPWR.n5579 4.6505
R6101 VPWR.n5584 VPWR.n5583 4.6505
R6102 VPWR.n5586 VPWR.n5585 4.6505
R6103 VPWR.n5588 VPWR.n5587 4.6505
R6104 VPWR.n5589 VPWR.n473 4.6505
R6105 VPWR.n5591 VPWR.n5590 4.6505
R6106 VPWR.n5594 VPWR.n5593 4.6505
R6107 VPWR.n5597 VPWR.n5596 4.6505
R6108 VPWR.n5600 VPWR.n5599 4.6505
R6109 VPWR.n5602 VPWR.n5601 4.6505
R6110 VPWR.n5604 VPWR.n5603 4.6505
R6111 VPWR.n5608 VPWR.n5607 4.6505
R6112 VPWR.n5610 VPWR.n5609 4.6505
R6113 VPWR.n5612 VPWR.n5611 4.6505
R6114 VPWR.n5616 VPWR.n5615 4.6505
R6115 VPWR.n5618 VPWR.n5617 4.6505
R6116 VPWR.n5619 VPWR.n458 4.6505
R6117 VPWR.n5621 VPWR.n5620 4.6505
R6118 VPWR.n5624 VPWR.n5623 4.6505
R6119 VPWR.n5625 VPWR.n457 4.6505
R6120 VPWR.n5627 VPWR.n5626 4.6505
R6121 VPWR.n5630 VPWR.n5629 4.6505
R6122 VPWR.n5632 VPWR.n5631 4.6505
R6123 VPWR.n5636 VPWR.n5635 4.6505
R6124 VPWR.n5639 VPWR.n5638 4.6505
R6125 VPWR.n5640 VPWR.n451 4.6505
R6126 VPWR.n5642 VPWR.n5641 4.6505
R6127 VPWR.n5644 VPWR.n5643 4.6505
R6128 VPWR.n5649 VPWR.n5648 4.6505
R6129 VPWR.n5651 VPWR.n5650 4.6505
R6130 VPWR.n5653 VPWR.n5652 4.6505
R6131 VPWR.n5404 VPWR.n5403 4.6505
R6132 VPWR.n5406 VPWR.n5405 4.6505
R6133 VPWR.n5410 VPWR.n5409 4.6505
R6134 VPWR.n5412 VPWR.n5411 4.6505
R6135 VPWR.n5416 VPWR.n5415 4.6505
R6136 VPWR.n5420 VPWR.n5419 4.6505
R6137 VPWR.n5424 VPWR.n5423 4.6505
R6138 VPWR.n5426 VPWR.n5425 4.6505
R6139 VPWR.n5432 VPWR.n5431 4.6505
R6140 VPWR.n5436 VPWR.n5435 4.6505
R6141 VPWR.n5440 VPWR.n5439 4.6505
R6142 VPWR.n5444 VPWR.n5443 4.6505
R6143 VPWR.n5446 VPWR.n5445 4.6505
R6144 VPWR.n5454 VPWR.n5453 4.6505
R6145 VPWR.n5457 VPWR.n5456 4.6505
R6146 VPWR.n5464 VPWR.n5463 4.6505
R6147 VPWR.n5469 VPWR.n5468 4.6505
R6148 VPWR.n5471 VPWR.n5470 4.6505
R6149 VPWR.n5475 VPWR.n5474 4.6505
R6150 VPWR.n5477 VPWR.n5476 4.6505
R6151 VPWR.n5480 VPWR.n5479 4.6505
R6152 VPWR.n5483 VPWR.n491 4.6505
R6153 VPWR.n5485 VPWR.n5484 4.6505
R6154 VPWR.n5487 VPWR.n5486 4.6505
R6155 VPWR.n5489 VPWR.n5488 4.6505
R6156 VPWR.n5492 VPWR.n5491 4.6505
R6157 VPWR.n5494 VPWR.n5493 4.6505
R6158 VPWR.n5496 VPWR.n5495 4.6505
R6159 VPWR.n1430 VPWR.n1429 4.6505
R6160 VPWR.n1432 VPWR.n1387 4.6505
R6161 VPWR.n1437 VPWR.n1436 4.6505
R6162 VPWR.n1451 VPWR.n1450 4.6505
R6163 VPWR.n1455 VPWR.n1454 4.6505
R6164 VPWR.n1459 VPWR.n1458 4.6505
R6165 VPWR.n1461 VPWR.n1460 4.6505
R6166 VPWR.n1463 VPWR.n1462 4.6505
R6167 VPWR.n1465 VPWR.n1464 4.6505
R6168 VPWR.n1469 VPWR.n1468 4.6505
R6169 VPWR.n1471 VPWR.n1470 4.6505
R6170 VPWR.n1474 VPWR.n1473 4.6505
R6171 VPWR.n1477 VPWR.n1476 4.6505
R6172 VPWR.n1479 VPWR.n1478 4.6505
R6173 VPWR.n1481 VPWR.n1480 4.6505
R6174 VPWR.n1485 VPWR.n1484 4.6505
R6175 VPWR.n1487 VPWR.n1486 4.6505
R6176 VPWR.n1490 VPWR.n1489 4.6505
R6177 VPWR.n1494 VPWR.n1493 4.6505
R6178 VPWR.n1496 VPWR.n1495 4.6505
R6179 VPWR.n1497 VPWR.n1374 4.6505
R6180 VPWR.n1504 VPWR.n1503 4.6505
R6181 VPWR.n1510 VPWR.n1509 4.6505
R6182 VPWR.n1512 VPWR.n1511 4.6505
R6183 VPWR.n1516 VPWR.n1515 4.6505
R6184 VPWR.n1299 VPWR.n1298 4.6505
R6185 VPWR.n1303 VPWR.n1302 4.6505
R6186 VPWR.n1308 VPWR.n1307 4.6505
R6187 VPWR.n1311 VPWR.n1310 4.6505
R6188 VPWR.n1313 VPWR.n1312 4.6505
R6189 VPWR.n1317 VPWR.n1316 4.6505
R6190 VPWR.n1319 VPWR.n1318 4.6505
R6191 VPWR.n1322 VPWR.n1321 4.6505
R6192 VPWR.n1644 VPWR.n1643 4.6505
R6193 VPWR.n1714 VPWR.n1713 4.6505
R6194 VPWR.n1717 VPWR.n1716 4.6505
R6195 VPWR.n1773 VPWR.n549 4.6505
R6196 VPWR.n1770 VPWR.n1726 4.6505
R6197 VPWR.n1555 VPWR.n1554 4.6505
R6198 VPWR.n1559 VPWR.n1558 4.6505
R6199 VPWR.n1570 VPWR.n1544 4.6505
R6200 VPWR.n1574 VPWR.n1573 4.6505
R6201 VPWR.n1658 VPWR.n1657 4.6505
R6202 VPWR.n1661 VPWR.n1660 4.6505
R6203 VPWR.n1666 VPWR.n1665 4.6505
R6204 VPWR.n1672 VPWR.n1671 4.6505
R6205 VPWR.n1674 VPWR.n1673 4.6505
R6206 VPWR.n1681 VPWR.n1680 4.6505
R6207 VPWR.n1683 VPWR.n1682 4.6505
R6208 VPWR.n1688 VPWR.n1687 4.6505
R6209 VPWR.n1691 VPWR.n1690 4.6505
R6210 VPWR.n1693 VPWR.n1692 4.6505
R6211 VPWR.n1696 VPWR.n1695 4.6505
R6212 VPWR.n1698 VPWR.n1697 4.6505
R6213 VPWR.n1700 VPWR.n1699 4.6505
R6214 VPWR.n1702 VPWR.n1701 4.6505
R6215 VPWR.n1705 VPWR.n1704 4.6505
R6216 VPWR.n1707 VPWR.n1706 4.6505
R6217 VPWR.n1709 VPWR.n1708 4.6505
R6218 VPWR.n1712 VPWR.n1711 4.6505
R6219 VPWR.n1721 VPWR.n1720 4.6505
R6220 VPWR.n1724 VPWR.n1723 4.6505
R6221 VPWR.n1775 VPWR.n1774 4.6505
R6222 VPWR.n5322 VPWR.n526 4.6505
R6223 VPWR.n5321 VPWR.n528 4.6505
R6224 VPWR.n5302 VPWR.n541 4.6505
R6225 VPWR.n5301 VPWR.n543 4.6505
R6226 VPWR.n5298 VPWR.n545 4.6505
R6227 VPWR.n5295 VPWR.n5294 4.6505
R6228 VPWR.n5292 VPWR.n547 4.6505
R6229 VPWR.n5285 VPWR.n1782 4.6505
R6230 VPWR.n5282 VPWR.n5281 4.6505
R6231 VPWR.n5280 VPWR.n1783 4.6505
R6232 VPWR.n5279 VPWR.n1784 4.6505
R6233 VPWR.n5278 VPWR.n1785 4.6505
R6234 VPWR.n4686 VPWR.n4685 4.6505
R6235 VPWR.n4762 VPWR.n4688 4.6505
R6236 VPWR.n4749 VPWR.n4748 4.6505
R6237 VPWR.n4735 VPWR.n4698 4.6505
R6238 VPWR.n4719 VPWR.n4704 4.6505
R6239 VPWR.n4718 VPWR.n4705 4.6505
R6240 VPWR.n4716 VPWR.n4708 4.6505
R6241 VPWR.n4715 VPWR.n4710 4.6505
R6242 VPWR.n4842 VPWR.n4841 4.6505
R6243 VPWR.n4837 VPWR.n4836 4.6505
R6244 VPWR.n4835 VPWR.n4834 4.6505
R6245 VPWR.n4833 VPWR.n4832 4.6505
R6246 VPWR.n4829 VPWR.n4828 4.6505
R6247 VPWR.n4827 VPWR.n4826 4.6505
R6248 VPWR.n4825 VPWR.n4824 4.6505
R6249 VPWR.n4823 VPWR.n4822 4.6505
R6250 VPWR.n4821 VPWR.n4790 4.6505
R6251 VPWR.n4820 VPWR.n4819 4.6505
R6252 VPWR.n4818 VPWR.n4817 4.6505
R6253 VPWR.n4816 VPWR.n4791 4.6505
R6254 VPWR.n4815 VPWR.n4814 4.6505
R6255 VPWR.n4811 VPWR.n4810 4.6505
R6256 VPWR.n4809 VPWR.n4808 4.6505
R6257 VPWR.n4805 VPWR.n4804 4.6505
R6258 VPWR.n4803 VPWR.n4802 4.6505
R6259 VPWR.n4676 VPWR.n4675 4.6505
R6260 VPWR.n4682 VPWR.n4681 4.6505
R6261 VPWR.n4684 VPWR.n4683 4.6505
R6262 VPWR.n4687 VPWR.n4647 4.6505
R6263 VPWR.n4764 VPWR.n4763 4.6505
R6264 VPWR.n4761 VPWR.n4760 4.6505
R6265 VPWR.n4759 VPWR.n4758 4.6505
R6266 VPWR.n4756 VPWR.n4755 4.6505
R6267 VPWR.n4754 VPWR.n4691 4.6505
R6268 VPWR.n4753 VPWR.n4752 4.6505
R6269 VPWR.n4751 VPWR.n4750 4.6505
R6270 VPWR.n4747 VPWR.n4697 4.6505
R6271 VPWR.n4746 VPWR.n4745 4.6505
R6272 VPWR.n4742 VPWR.n4741 4.6505
R6273 VPWR.n4740 VPWR.n4739 4.6505
R6274 VPWR.n4734 VPWR.n4733 4.6505
R6275 VPWR.n4728 VPWR.n4727 4.6505
R6276 VPWR.n4724 VPWR.n4723 4.6505
R6277 VPWR.n4722 VPWR.n4702 4.6505
R6278 VPWR.n4721 VPWR.n4720 4.6505
R6279 VPWR.n4767 VPWR.n4646 4.6505
R6280 VPWR.n4768 VPWR.n4767 4.6505
R6281 VPWR.n4770 VPWR.n4769 4.6505
R6282 VPWR.n4774 VPWR.n4773 4.6505
R6283 VPWR.n4776 VPWR.n4775 4.6505
R6284 VPWR.n4784 VPWR.n4783 4.6505
R6285 VPWR.n5319 VPWR.n5318 4.6505
R6286 VPWR.n5317 VPWR.n5316 4.6505
R6287 VPWR.n5315 VPWR.n5314 4.6505
R6288 VPWR.n5312 VPWR.n5311 4.6505
R6289 VPWR.n5310 VPWR.n5309 4.6505
R6290 VPWR.n5306 VPWR.n5305 4.6505
R6291 VPWR.n5300 VPWR.n5299 4.6505
R6292 VPWR.n5297 VPWR.n5296 4.6505
R6293 VPWR.n5293 VPWR.n546 4.6505
R6294 VPWR.n5291 VPWR.n5290 4.6505
R6295 VPWR.n5289 VPWR.n5288 4.6505
R6296 VPWR.n5287 VPWR.n5286 4.6505
R6297 VPWR.n5284 VPWR.n5283 4.6505
R6298 VPWR.n5277 VPWR.n5276 4.6505
R6299 VPWR.n5275 VPWR.n5274 4.6505
R6300 VPWR.n5273 VPWR.n5272 4.6505
R6301 VPWR.n5271 VPWR.n5270 4.6505
R6302 VPWR.n5269 VPWR.n5268 4.6505
R6303 VPWR.n5267 VPWR.n5266 4.6505
R6304 VPWR.n5264 VPWR.n5263 4.6505
R6305 VPWR.n5262 VPWR.n5261 4.6505
R6306 VPWR.n5260 VPWR.n5259 4.6505
R6307 VPWR.n5258 VPWR.n5257 4.6505
R6308 VPWR.n5256 VPWR.n5255 4.6505
R6309 VPWR.n1772 VPWR.n1771 4.6505
R6310 VPWR.n1668 VPWR.n1667 4.6505
R6311 VPWR.n1663 VPWR.n1662 4.6505
R6312 VPWR.n1659 VPWR.n560 4.6505
R6313 VPWR.n1654 VPWR.n1653 4.6505
R6314 VPWR.n1652 VPWR.n1651 4.6505
R6315 VPWR.n1649 VPWR.n1648 4.6505
R6316 VPWR.n1646 VPWR.n1645 4.6505
R6317 VPWR.n1557 VPWR.n1556 4.6505
R6318 VPWR.n1561 VPWR.n1560 4.6505
R6319 VPWR.n1567 VPWR.n1566 4.6505
R6320 VPWR.n1569 VPWR.n1568 4.6505
R6321 VPWR.n1572 VPWR.n1571 4.6505
R6322 VPWR.n1576 VPWR.n1575 4.6505
R6323 VPWR.n1579 VPWR.n1578 4.6505
R6324 VPWR.n1583 VPWR.n1582 4.6505
R6325 VPWR.n1586 VPWR.n1585 4.6505
R6326 VPWR.n2548 VPWR.n2547 4.6505
R6327 VPWR.n2566 VPWR.n2186 4.6505
R6328 VPWR.n2143 VPWR.n2122 4.6505
R6329 VPWR.n2142 VPWR.n2124 4.6505
R6330 VPWR.n2125 VPWR.n2115 4.6505
R6331 VPWR.n2570 VPWR.n2569 4.6505
R6332 VPWR.n2444 VPWR.n2443 4.6505
R6333 VPWR.n2448 VPWR.n2447 4.6505
R6334 VPWR.n2557 VPWR.n2556 4.6505
R6335 VPWR.n2561 VPWR.n2560 4.6505
R6336 VPWR.n2184 VPWR.n2183 4.6505
R6337 VPWR.n2180 VPWR.n2179 4.6505
R6338 VPWR.n2178 VPWR.n2177 4.6505
R6339 VPWR.n2174 VPWR.n2173 4.6505
R6340 VPWR.n2172 VPWR.n2171 4.6505
R6341 VPWR.n2169 VPWR.n2168 4.6505
R6342 VPWR.n2167 VPWR.n2166 4.6505
R6343 VPWR.n2164 VPWR.n2163 4.6505
R6344 VPWR.n2162 VPWR.n2161 4.6505
R6345 VPWR.n2158 VPWR.n2157 4.6505
R6346 VPWR.n2156 VPWR.n2155 4.6505
R6347 VPWR.n2154 VPWR.n2153 4.6505
R6348 VPWR.n2136 VPWR.n2135 4.6505
R6349 VPWR.n2132 VPWR.n2131 4.6505
R6350 VPWR.n5157 VPWR.n1830 4.6505
R6351 VPWR.n5144 VPWR.n1832 4.6505
R6352 VPWR.n5139 VPWR.n1833 4.6505
R6353 VPWR.n5123 VPWR.n5122 4.6505
R6354 VPWR.n5119 VPWR.n5117 4.6505
R6355 VPWR.n5113 VPWR.n1848 4.6505
R6356 VPWR.n5112 VPWR.n1849 4.6505
R6357 VPWR.n5111 VPWR.n1850 4.6505
R6358 VPWR.n5100 VPWR.n5099 4.6505
R6359 VPWR.n5085 VPWR.n1853 4.6505
R6360 VPWR.n1912 VPWR.n1892 4.6505
R6361 VPWR.n1920 VPWR.n1919 4.6505
R6362 VPWR.n1922 VPWR.n1921 4.6505
R6363 VPWR.n1925 VPWR.n1924 4.6505
R6364 VPWR.n1930 VPWR.n1927 4.6505
R6365 VPWR.n1931 VPWR.n1909 4.6505
R6366 VPWR.n1944 VPWR.n1943 4.6505
R6367 VPWR.n1948 VPWR.n1947 4.6505
R6368 VPWR.n5015 VPWR.n1958 4.6505
R6369 VPWR.n4936 VPWR.n4935 4.6505
R6370 VPWR.n4953 VPWR.n4952 4.6505
R6371 VPWR.n4949 VPWR.n4948 4.6505
R6372 VPWR.n4945 VPWR.n4944 4.6505
R6373 VPWR.n4942 VPWR.n4941 4.6505
R6374 VPWR.n4940 VPWR.n4939 4.6505
R6375 VPWR.n4938 VPWR.n4937 4.6505
R6376 VPWR.n4934 VPWR.n4920 4.6505
R6377 VPWR.n4931 VPWR.n4930 4.6505
R6378 VPWR.n4965 VPWR.n4964 4.6505
R6379 VPWR.n4961 VPWR.n4960 4.6505
R6380 VPWR.n4959 VPWR.n4958 4.6505
R6381 VPWR.n4957 VPWR.n4956 4.6505
R6382 VPWR.n4955 VPWR.n4954 4.6505
R6383 VPWR.n5031 VPWR.n5030 4.6505
R6384 VPWR.n5029 VPWR.n5028 4.6505
R6385 VPWR.n5026 VPWR.n5025 4.6505
R6386 VPWR.n5024 VPWR.n5023 4.6505
R6387 VPWR.n5021 VPWR.n5020 4.6505
R6388 VPWR.n5019 VPWR.n5018 4.6505
R6389 VPWR VPWR.n1913 4.6505
R6390 VPWR.n1915 VPWR.n1914 4.6505
R6391 VPWR.n1917 VPWR.n1916 4.6505
R6392 VPWR.n1933 VPWR.n1932 4.6505
R6393 VPWR.n1937 VPWR.n1936 4.6505
R6394 VPWR.n1941 VPWR.n1940 4.6505
R6395 VPWR.n1946 VPWR.n1945 4.6505
R6396 VPWR.n1949 VPWR.n1899 4.6505
R6397 VPWR.n1954 VPWR.n1953 4.6505
R6398 VPWR.n1957 VPWR.n1898 4.6505
R6399 VPWR.n5012 VPWR.n5011 4.6505
R6400 VPWR.n5010 VPWR.n1959 4.6505
R6401 VPWR.n5008 VPWR.n5007 4.6505
R6402 VPWR.n5159 VPWR.n5158 4.6505
R6403 VPWR.n5156 VPWR.n5155 4.6505
R6404 VPWR.n5154 VPWR.n5153 4.6505
R6405 VPWR.n5152 VPWR.n5151 4.6505
R6406 VPWR.n5148 VPWR.n5147 4.6505
R6407 VPWR.n5143 VPWR.n5142 4.6505
R6408 VPWR.n5141 VPWR.n1838 4.6505
R6409 VPWR.n5141 VPWR.n5140 4.6505
R6410 VPWR.n5138 VPWR.n5137 4.6505
R6411 VPWR.n5128 VPWR.n5127 4.6505
R6412 VPWR.n5126 VPWR.n5125 4.6505
R6413 VPWR.n5121 VPWR.n5120 4.6505
R6414 VPWR VPWR.n1840 4.6505
R6415 VPWR.n5116 VPWR.n5115 4.6505
R6416 VPWR.n5110 VPWR.n5109 4.6505
R6417 VPWR.n5108 VPWR.n5107 4.6505
R6418 VPWR.n5102 VPWR.n5101 4.6505
R6419 VPWR.n5098 VPWR.n5097 4.6505
R6420 VPWR.n5096 VPWR.n5095 4.6505
R6421 VPWR.n5090 VPWR.n5089 4.6505
R6422 VPWR.n5088 VPWR.n5087 4.6505
R6423 VPWR.n5086 VPWR.n1851 4.6505
R6424 VPWR.n2576 VPWR.n2575 4.6505
R6425 VPWR.n2574 VPWR.n2573 4.6505
R6426 VPWR.n2572 VPWR.n2571 4.6505
R6427 VPWR.n2139 VPWR.n2138 4.6505
R6428 VPWR.n2141 VPWR.n2140 4.6505
R6429 VPWR.n2145 VPWR.n2144 4.6505
R6430 VPWR.n2150 VPWR.n2149 4.6505
R6431 VPWR.n2152 VPWR.n2151 4.6505
R6432 VPWR.n2553 VPWR.n2552 4.6505
R6433 VPWR.n2551 VPWR.n2550 4.6505
R6434 VPWR.n2442 VPWR.n2432 4.6505
R6435 VPWR.n2446 VPWR.n2445 4.6505
R6436 VPWR.n2451 VPWR.n2450 4.6505
R6437 VPWR.n2452 VPWR.n2430 4.6505
R6438 VPWR.n2455 VPWR.n2454 4.6505
R6439 VPWR.n2462 VPWR.n2461 4.6505
R6440 VPWR.n2463 VPWR.n2426 4.6505
R6441 VPWR.n2465 VPWR.n2464 4.6505
R6442 VPWR.n2470 VPWR.n2469 4.6505
R6443 VPWR.n2472 VPWR.n2471 4.6505
R6444 VPWR.n2476 VPWR.n2475 4.6505
R6445 VPWR.n2482 VPWR.n2481 4.6505
R6446 VPWR.n4411 VPWR.n2009 4.6505
R6447 VPWR.n4423 VPWR.n4422 4.6505
R6448 VPWR.n4425 VPWR.n4424 4.6505
R6449 VPWR.n4426 VPWR.n2008 4.6505
R6450 VPWR.n4455 VPWR.n4454 4.6505
R6451 VPWR.n4457 VPWR.n4456 4.6505
R6452 VPWR.n2061 VPWR.n2044 4.6505
R6453 VPWR.n2046 VPWR.n2031 4.6505
R6454 VPWR.n2693 VPWR.n2032 4.6505
R6455 VPWR.n2370 VPWR.n2302 4.6505
R6456 VPWR.n2333 VPWR.n2308 4.6505
R6457 VPWR.n2332 VPWR.n2310 4.6505
R6458 VPWR.n2331 VPWR.n2312 4.6505
R6459 VPWR.n2329 VPWR.n2314 4.6505
R6460 VPWR.n2326 VPWR.n2325 4.6505
R6461 VPWR.n2320 VPWR.n2316 4.6505
R6462 VPWR.n2317 VPWR.n2035 4.6505
R6463 VPWR.n2687 VPWR.n2034 4.6505
R6464 VPWR.n2686 VPWR.n2036 4.6505
R6465 VPWR.n2224 VPWR.n2223 4.6505
R6466 VPWR.n2227 VPWR.n2226 4.6505
R6467 VPWR.n2230 VPWR.n2228 4.6505
R6468 VPWR.n2377 VPWR.n2376 4.6505
R6469 VPWR.n2372 VPWR.n2371 4.6505
R6470 VPWR.n2364 VPWR.n2363 4.6505
R6471 VPWR.n2362 VPWR.n2361 4.6505
R6472 VPWR.n2360 VPWR.n2359 4.6505
R6473 VPWR.n2358 VPWR.n2357 4.6505
R6474 VPWR.n2356 VPWR.n2355 4.6505
R6475 VPWR.n2352 VPWR.n2351 4.6505
R6476 VPWR.n2350 VPWR.n2349 4.6505
R6477 VPWR.n2346 VPWR.n2345 4.6505
R6478 VPWR.n2344 VPWR.n2343 4.6505
R6479 VPWR.n2342 VPWR.n2341 4.6505
R6480 VPWR.n2340 VPWR.n2339 4.6505
R6481 VPWR.n2338 VPWR.n2337 4.6505
R6482 VPWR.n2685 VPWR.n2684 4.6505
R6483 VPWR.n2101 VPWR.n2100 4.6505
R6484 VPWR.n2099 VPWR.n2098 4.6505
R6485 VPWR.n2095 VPWR.n2094 4.6505
R6486 VPWR.n2093 VPWR.n2092 4.6505
R6487 VPWR.n2087 VPWR.n2086 4.6505
R6488 VPWR.n2082 VPWR.n2081 4.6505
R6489 VPWR.n2080 VPWR.n2079 4.6505
R6490 VPWR.n2076 VPWR.n2075 4.6505
R6491 VPWR.n2071 VPWR.n2070 4.6505
R6492 VPWR.n2069 VPWR.n2068 4.6505
R6493 VPWR.n2065 VPWR.n2064 4.6505
R6494 VPWR.n2050 VPWR.n2049 4.6505
R6495 VPWR.n2697 VPWR.n2696 4.6505
R6496 VPWR.n2702 VPWR.n2701 4.6505
R6497 VPWR.n2704 VPWR.n2703 4.6505
R6498 VPWR.n2706 VPWR.n2705 4.6505
R6499 VPWR.n2710 VPWR.n2709 4.6505
R6500 VPWR.n2713 VPWR.n2712 4.6505
R6501 VPWR.n2715 VPWR.n2714 4.6505
R6502 VPWR.n2716 VPWR.n2022 4.6505
R6503 VPWR.n2718 VPWR.n2717 4.6505
R6504 VPWR.n2721 VPWR.n2720 4.6505
R6505 VPWR.n2724 VPWR.n2021 4.6505
R6506 VPWR.n4409 VPWR.n4408 4.6505
R6507 VPWR.n4437 VPWR.n4436 4.6505
R6508 VPWR.n4461 VPWR.n4460 4.6505
R6509 VPWR.n4468 VPWR.n4467 4.6505
R6510 VPWR.n4470 VPWR.n4469 4.6505
R6511 VPWR.n4472 VPWR.n4471 4.6505
R6512 VPWR.n4475 VPWR.n2005 4.6505
R6513 VPWR.n4477 VPWR.n4476 4.6505
R6514 VPWR.n4506 VPWR.n4495 4.6505
R6515 VPWR.n4505 VPWR.n4496 4.6505
R6516 VPWR.n4539 VPWR.n4538 4.6505
R6517 VPWR.n4536 VPWR.n4535 4.6505
R6518 VPWR.n4534 VPWR.n4533 4.6505
R6519 VPWR.n4525 VPWR.n4524 4.6505
R6520 VPWR.n4523 VPWR.n4522 4.6505
R6521 VPWR.n4520 VPWR.n4519 4.6505
R6522 VPWR.n4518 VPWR.n4517 4.6505
R6523 VPWR.n4516 VPWR.n4488 4.6505
R6524 VPWR.n4515 VPWR.n4514 4.6505
R6525 VPWR.n4513 VPWR.n4512 4.6505
R6526 VPWR.n4511 VPWR.n4492 4.6505
R6527 VPWR.n4510 VPWR.n4509 4.6505
R6528 VPWR.n4508 VPWR.n4507 4.6505
R6529 VPWR.n4482 VPWR.n4481 4.6505
R6530 VPWR.n4480 VPWR.n4479 4.6505
R6531 VPWR.n4463 VPWR.n4462 4.6505
R6532 VPWR.n4453 VPWR.n4452 4.6505
R6533 VPWR.n4450 VPWR.n4449 4.6505
R6534 VPWR.n4448 VPWR.n4447 4.6505
R6535 VPWR.n4445 VPWR.n4444 4.6505
R6536 VPWR.n4443 VPWR.n4442 4.6505
R6537 VPWR.n4428 VPWR.n4427 4.6505
R6538 VPWR.n4419 VPWR.n4418 4.6505
R6539 VPWR.n4405 VPWR.n4404 4.6505
R6540 VPWR.n2732 VPWR.n2731 4.6505
R6541 VPWR.n2730 VPWR.n2729 4.6505
R6542 VPWR.n2726 VPWR.n2725 4.6505
R6543 VPWR.n2060 VPWR.n2059 4.6505
R6544 VPWR.n2689 VPWR.n2688 4.6505
R6545 VPWR.n2319 VPWR.n2318 4.6505
R6546 VPWR.n2322 VPWR.n2321 4.6505
R6547 VPWR.n2324 VPWR.n2323 4.6505
R6548 VPWR.n2328 VPWR.n2327 4.6505
R6549 VPWR.n2335 VPWR.n2334 4.6505
R6550 VPWR.n2366 VPWR.n2365 4.6505
R6551 VPWR.n2369 VPWR.n2368 4.6505
R6552 VPWR.n2232 VPWR.n2231 4.6505
R6553 VPWR.n2237 VPWR.n2236 4.6505
R6554 VPWR.n2239 VPWR.n2238 4.6505
R6555 VPWR.n2242 VPWR.n2241 4.6505
R6556 VPWR.n2246 VPWR.n2245 4.6505
R6557 VPWR.n2250 VPWR.n2249 4.6505
R6558 VPWR.n2252 VPWR.n2251 4.6505
R6559 VPWR.n2254 VPWR.n2253 4.6505
R6560 VPWR.n2257 VPWR.n2256 4.6505
R6561 VPWR.n2261 VPWR.n2260 4.6505
R6562 VPWR.n2265 VPWR.n2264 4.6505
R6563 VPWR.n2267 VPWR.n2266 4.6505
R6564 VPWR.n2269 VPWR.n2268 4.6505
R6565 VPWR.n3576 VPWR.n3575 4.6505
R6566 VPWR.n3672 VPWR.n3671 4.6505
R6567 VPWR.n3733 VPWR.n3499 4.6505
R6568 VPWR.n3732 VPWR.n3500 4.6505
R6569 VPWR.n3688 VPWR.n3516 4.6505
R6570 VPWR.n3685 VPWR.n3517 4.6505
R6571 VPWR.n3675 VPWR.n3518 4.6505
R6572 VPWR.n3540 VPWR.n3539 4.6505
R6573 VPWR.n3409 VPWR.n3371 4.6505
R6574 VPWR.n3414 VPWR.n3413 4.6505
R6575 VPWR.n3418 VPWR.n3416 4.6505
R6576 VPWR.n3728 VPWR.n3727 4.6505
R6577 VPWR.n3721 VPWR.n3720 4.6505
R6578 VPWR.n3719 VPWR.n3718 4.6505
R6579 VPWR.n3717 VPWR.n3716 4.6505
R6580 VPWR.n3715 VPWR.n3714 4.6505
R6581 VPWR.n3711 VPWR.n3710 4.6505
R6582 VPWR.n3709 VPWR.n3708 4.6505
R6583 VPWR.n3706 VPWR.n3705 4.6505
R6584 VPWR.n3704 VPWR.n3703 4.6505
R6585 VPWR.n3702 VPWR.n3701 4.6505
R6586 VPWR.n3699 VPWR.n3698 4.6505
R6587 VPWR.n3697 VPWR.n3696 4.6505
R6588 VPWR.n3695 VPWR.n3694 4.6505
R6589 VPWR.n3693 VPWR.n3692 4.6505
R6590 VPWR.n3586 VPWR.n3585 4.6505
R6591 VPWR.n3590 VPWR.n3589 4.6505
R6592 VPWR.n3592 VPWR.n3591 4.6505
R6593 VPWR.n3594 VPWR.n3593 4.6505
R6594 VPWR.n3597 VPWR.n3596 4.6505
R6595 VPWR.n3600 VPWR.n3599 4.6505
R6596 VPWR.n3602 VPWR.n3601 4.6505
R6597 VPWR.n3604 VPWR.n3603 4.6505
R6598 VPWR.n3609 VPWR.n3608 4.6505
R6599 VPWR.n3610 VPWR.n3525 4.6505
R6600 VPWR.n3612 VPWR.n3611 4.6505
R6601 VPWR.n3615 VPWR.n3614 4.6505
R6602 VPWR.n3617 VPWR.n3616 4.6505
R6603 VPWR.n3619 VPWR.n3618 4.6505
R6604 VPWR.n3622 VPWR.n3621 4.6505
R6605 VPWR.n3623 VPWR.n3523 4.6505
R6606 VPWR.n3668 VPWR.n3667 4.6505
R6607 VPWR.n3664 VPWR.n3663 4.6505
R6608 VPWR.n3662 VPWR.n3661 4.6505
R6609 VPWR.n3660 VPWR.n3659 4.6505
R6610 VPWR.n3658 VPWR.n3657 4.6505
R6611 VPWR.n3656 VPWR.n3655 4.6505
R6612 VPWR.n3652 VPWR.n3651 4.6505
R6613 VPWR.n3649 VPWR.n3648 4.6505
R6614 VPWR.n3646 VPWR.n3645 4.6505
R6615 VPWR.n3644 VPWR.n3643 4.6505
R6616 VPWR.n3642 VPWR.n3641 4.6505
R6617 VPWR.n3640 VPWR.n3639 4.6505
R6618 VPWR.n4250 VPWR.n2789 4.6505
R6619 VPWR.n2836 VPWR.n2835 4.6505
R6620 VPWR.n4245 VPWR.n2792 4.6505
R6621 VPWR.n2935 VPWR.n2934 4.6505
R6622 VPWR.n2929 VPWR.n2928 4.6505
R6623 VPWR.n2927 VPWR.n2926 4.6505
R6624 VPWR.n2925 VPWR.n2924 4.6505
R6625 VPWR.n2923 VPWR.n2922 4.6505
R6626 VPWR.n2921 VPWR.n2920 4.6505
R6627 VPWR.n2918 VPWR.n2917 4.6505
R6628 VPWR.n2916 VPWR.n2915 4.6505
R6629 VPWR.n2914 VPWR.n2913 4.6505
R6630 VPWR.n2911 VPWR.n2910 4.6505
R6631 VPWR.n2909 VPWR.n2908 4.6505
R6632 VPWR.n2907 VPWR.n2906 4.6505
R6633 VPWR.n2905 VPWR.n2904 4.6505
R6634 VPWR.n2903 VPWR.n2902 4.6505
R6635 VPWR.n2901 VPWR.n2900 4.6505
R6636 VPWR.n2899 VPWR.n2898 4.6505
R6637 VPWR.n4259 VPWR.n4258 4.6505
R6638 VPWR.n4257 VPWR.n4256 4.6505
R6639 VPWR.n4255 VPWR.n4254 4.6505
R6640 VPWR.n4252 VPWR.n4251 4.6505
R6641 VPWR.n2797 VPWR.n2796 4.6505
R6642 VPWR.n2799 VPWR.n2798 4.6505
R6643 VPWR.n2802 VPWR.n2801 4.6505
R6644 VPWR.n2804 VPWR.n2803 4.6505
R6645 VPWR.n2807 VPWR.n2806 4.6505
R6646 VPWR.n2809 VPWR.n2808 4.6505
R6647 VPWR.n2812 VPWR.n2811 4.6505
R6648 VPWR.n2816 VPWR.n2815 4.6505
R6649 VPWR.n2820 VPWR.n2819 4.6505
R6650 VPWR.n2823 VPWR.n2822 4.6505
R6651 VPWR.n2830 VPWR.n2829 4.6505
R6652 VPWR.n2832 VPWR.n2831 4.6505
R6653 VPWR.n2839 VPWR.n2838 4.6505
R6654 VPWR.n2841 VPWR.n2840 4.6505
R6655 VPWR.n2845 VPWR.n2844 4.6505
R6656 VPWR.n2848 VPWR.n2847 4.6505
R6657 VPWR.n2850 VPWR.n2849 4.6505
R6658 VPWR.n2852 VPWR.n2851 4.6505
R6659 VPWR.n2855 VPWR.n2854 4.6505
R6660 VPWR.n2857 VPWR.n2856 4.6505
R6661 VPWR.n2861 VPWR.n2860 4.6505
R6662 VPWR.n2863 VPWR.n2862 4.6505
R6663 VPWR.n2864 VPWR.n2794 4.6505
R6664 VPWR.n4247 VPWR.n4246 4.6505
R6665 VPWR.n4244 VPWR.n4243 4.6505
R6666 VPWR.n4240 VPWR.n4239 4.6505
R6667 VPWR.n4238 VPWR.n4237 4.6505
R6668 VPWR.n4236 VPWR.n4235 4.6505
R6669 VPWR.n4261 VPWR.n4260 4.6505
R6670 VPWR.n3634 VPWR.n2784 4.6505
R6671 VPWR.n3670 VPWR.n3669 4.6505
R6672 VPWR.n3578 VPWR.n3577 4.6505
R6673 VPWR.n3538 VPWR.n3537 4.6505
R6674 VPWR.n3536 VPWR.n3535 4.6505
R6675 VPWR.n3677 VPWR.n3676 4.6505
R6676 VPWR.n3682 VPWR.n3681 4.6505
R6677 VPWR.n3684 VPWR.n3683 4.6505
R6678 VPWR.n3687 VPWR.n3686 4.6505
R6679 VPWR.n3690 VPWR.n3689 4.6505
R6680 VPWR.n3731 VPWR.n3730 4.6505
R6681 VPWR.n3734 VPWR.n3498 4.6505
R6682 VPWR.n3736 VPWR.n3735 4.6505
R6683 VPWR.n3739 VPWR.n3738 4.6505
R6684 VPWR.n3742 VPWR.n3741 4.6505
R6685 VPWR.n3744 VPWR.n3743 4.6505
R6686 VPWR.n3746 VPWR.n3745 4.6505
R6687 VPWR.n3388 VPWR.n3387 4.6505
R6688 VPWR.n3393 VPWR.n3392 4.6505
R6689 VPWR.n3395 VPWR.n3394 4.6505
R6690 VPWR.n3398 VPWR.n3397 4.6505
R6691 VPWR.n3408 VPWR.n3407 4.6505
R6692 VPWR.n3411 VPWR.n3410 4.6505
R6693 VPWR.n3415 VPWR.n3370 4.6505
R6694 VPWR.n3421 VPWR.n3420 4.6505
R6695 VPWR.n3424 VPWR.n3423 4.6505
R6696 VPWR.n6054 VPWR.n6053 4.6505
R6697 VPWR.n6106 VPWR.n6058 4.6505
R6698 VPWR.n6088 VPWR.n6087 4.6505
R6699 VPWR.n7739 VPWR.n7738 4.6505
R6700 VPWR.n7741 VPWR.n7740 4.6505
R6701 VPWR.n7743 VPWR.n7742 4.6505
R6702 VPWR.n7746 VPWR.n7745 4.6505
R6703 VPWR.n7748 VPWR.n7747 4.6505
R6704 VPWR.n7750 VPWR.n7749 4.6505
R6705 VPWR.n7753 VPWR.n7752 4.6505
R6706 VPWR.n7754 VPWR.n6128 4.6505
R6707 VPWR.n7772 VPWR.n7771 4.6505
R6708 VPWR.n7774 VPWR.n7773 4.6505
R6709 VPWR.n7777 VPWR.n7776 4.6505
R6710 VPWR.n7779 VPWR.n7778 4.6505
R6711 VPWR.n7782 VPWR.n7781 4.6505
R6712 VPWR.n7785 VPWR.n7784 4.6505
R6713 VPWR.n7787 VPWR.n7786 4.6505
R6714 VPWR.n7790 VPWR.n7789 4.6505
R6715 VPWR.n7794 VPWR.n7793 4.6505
R6716 VPWR.n7796 VPWR.n7795 4.6505
R6717 VPWR.n7798 VPWR.n7797 4.6505
R6718 VPWR.n7800 VPWR.n7799 4.6505
R6719 VPWR.n7803 VPWR.n7802 4.6505
R6720 VPWR.n7805 VPWR.n7804 4.6505
R6721 VPWR.n7807 VPWR.n6114 4.6505
R6722 VPWR.n7809 VPWR.n7808 4.6505
R6723 VPWR.n7812 VPWR.n7811 4.6505
R6724 VPWR.n7815 VPWR.n7814 4.6505
R6725 VPWR.n6007 VPWR.n6006 4.6505
R6726 VPWR.n6021 VPWR.n6020 4.6505
R6727 VPWR.n6023 VPWR.n6022 4.6505
R6728 VPWR.n6025 VPWR.n6024 4.6505
R6729 VPWR.n6027 VPWR.n6026 4.6505
R6730 VPWR.n6031 VPWR.n6030 4.6505
R6731 VPWR.n6034 VPWR.n6033 4.6505
R6732 VPWR.n6040 VPWR.n6039 4.6505
R6733 VPWR.n6108 VPWR.n6107 4.6505
R6734 VPWR.n6105 VPWR.n6104 4.6505
R6735 VPWR.n6102 VPWR.n6101 4.6505
R6736 VPWR.n6100 VPWR.n6099 4.6505
R6737 VPWR.n6097 VPWR.n6096 4.6505
R6738 VPWR.n6094 VPWR.n6093 4.6505
R6739 VPWR.n6090 VPWR.n6089 4.6505
R6740 VPWR.n6084 VPWR.n6083 4.6505
R6741 VPWR.n6077 VPWR.n6076 4.6505
R6742 VPWR.n6074 VPWR.n6073 4.6505
R6743 VPWR.n9139 VPWR.n9130 4.6505
R6744 VPWR.n88 VPWR.n64 4.6505
R6745 VPWR.n86 VPWR.n70 4.6505
R6746 VPWR.n85 VPWR.n72 4.6505
R6747 VPWR.n82 VPWR.n73 4.6505
R6748 VPWR.n104 VPWR.n103 4.6505
R6749 VPWR.n99 VPWR.n98 4.6505
R6750 VPWR.n97 VPWR.n96 4.6505
R6751 VPWR.n93 VPWR.n92 4.6505
R6752 VPWR.n91 VPWR.n63 4.6505
R6753 VPWR.n90 VPWR.n89 4.6505
R6754 VPWR.n84 VPWR.n83 4.6505
R6755 VPWR.n113 VPWR.n112 4.6505
R6756 VPWR.n108 VPWR.n107 4.6505
R6757 VPWR.n106 VPWR.n105 4.6505
R6758 VPWR.n9141 VPWR.n9140 4.6505
R6759 VPWR.n9154 VPWR.n52 4.6505
R6760 VPWR.n9153 VPWR.n9152 4.6505
R6761 VPWR.n9150 VPWR.n9149 4.6505
R6762 VPWR.n9146 VPWR.n9145 4.6505
R6763 VPWR.n9144 VPWR.n9143 4.6505
R6764 VPWR.n9156 VPWR.n9155 4.6505
R6765 VPWR.n9158 VPWR.n9157 4.6505
R6766 VPWR.n9159 VPWR.n51 4.6505
R6767 VPWR.n9167 VPWR.n9166 4.6505
R6768 VPWR.n9163 VPWR.n9162 4.6505
R6769 VPWR.n9161 VPWR.n9160 4.6505
R6770 VPWR.n9169 VPWR.n9168 4.6505
R6771 VPWR.n9171 VPWR.n9170 4.6505
R6772 VPWR.n9176 VPWR.n9175 4.6505
R6773 VPWR.n9188 VPWR.n9187 4.6505
R6774 VPWR.n9185 VPWR.n9184 4.6505
R6775 VPWR.n9181 VPWR.n9180 4.6505
R6776 VPWR.n9178 VPWR.n9177 4.6505
R6777 VPWR.n9190 VPWR.n9189 4.6505
R6778 VPWR.n9200 VPWR.n9199 4.6505
R6779 VPWR.n9198 VPWR.n32 4.6505
R6780 VPWR.n9197 VPWR.n9196 4.6505
R6781 VPWR.n9192 VPWR.n9191 4.6505
R6782 VPWR.n6072 VPWR.n6071 4.6505
R6783 VPWR.n6081 VPWR.n6080 4.6505
R6784 VPWR.n6086 VPWR.n6085 4.6505
R6785 VPWR.n6056 VPWR.n6055 4.6505
R6786 VPWR.n6052 VPWR.n6051 4.6505
R6787 VPWR.n6050 VPWR.n6049 4.6505
R6788 VPWR.n6048 VPWR.n6047 4.6505
R6789 VPWR.n6046 VPWR.n6045 4.6505
R6790 VPWR.n6041 VPWR.n6014 4.6505
R6791 VPWR.n6037 VPWR.n6036 4.6505
R6792 VPWR.n7756 VPWR.n7755 4.6505
R6793 VPWR.n7657 VPWR.n7656 4.6505
R6794 VPWR.n7661 VPWR.n7660 4.6505
R6795 VPWR.n7662 VPWR.n7639 4.6505
R6796 VPWR.n7664 VPWR.n7663 4.6505
R6797 VPWR.n7668 VPWR.n7667 4.6505
R6798 VPWR.n7670 VPWR.n7669 4.6505
R6799 VPWR.n7672 VPWR.n7671 4.6505
R6800 VPWR.n7674 VPWR.n7673 4.6505
R6801 VPWR.n7681 VPWR.n7680 4.6505
R6802 VPWR.n7686 VPWR.n7685 4.6505
R6803 VPWR.n3259 VPWR.n3258 4.6505
R6804 VPWR.n3262 VPWR.n3261 4.6505
R6805 VPWR.n3267 VPWR.n3266 4.6505
R6806 VPWR.n3281 VPWR.n3280 4.6505
R6807 VPWR.n3215 VPWR.n3212 4.6505
R6808 VPWR.n3174 VPWR.n3173 4.6505
R6809 VPWR.n3171 VPWR.n3155 4.6505
R6810 VPWR.n3164 VPWR.n3160 4.6505
R6811 VPWR.n3163 VPWR.n3161 4.6505
R6812 VPWR.n3874 VPWR.n3039 4.6505
R6813 VPWR.n3873 VPWR.n3042 4.6505
R6814 VPWR.n3074 VPWR.n3055 4.6505
R6815 VPWR.n4060 VPWR.n4058 4.6505
R6816 VPWR.n4071 VPWR.n2990 4.6505
R6817 VPWR.n4118 VPWR.n4090 4.6505
R6818 VPWR.n4124 VPWR.n4088 4.6505
R6819 VPWR.n4133 VPWR.n4132 4.6505
R6820 VPWR.n4131 VPWR.n4130 4.6505
R6821 VPWR.n4129 VPWR.n4128 4.6505
R6822 VPWR.n4121 VPWR.n4120 4.6505
R6823 VPWR.n4109 VPWR.n4108 4.6505
R6824 VPWR.n4123 VPWR.n4122 4.6505
R6825 VPWR.n4126 VPWR.n4125 4.6505
R6826 VPWR.n3994 VPWR.n3993 4.6505
R6827 VPWR.n3996 VPWR.n3995 4.6505
R6828 VPWR.n4000 VPWR.n3999 4.6505
R6829 VPWR.n4003 VPWR.n4002 4.6505
R6830 VPWR.n4004 VPWR.n2998 4.6505
R6831 VPWR.n4018 VPWR.n4017 4.6505
R6832 VPWR.n4023 VPWR.n4022 4.6505
R6833 VPWR.n4026 VPWR.n4025 4.6505
R6834 VPWR.n4034 VPWR.n4033 4.6505
R6835 VPWR.n4037 VPWR.n4036 4.6505
R6836 VPWR.n4039 VPWR.n4038 4.6505
R6837 VPWR.n4042 VPWR.n4041 4.6505
R6838 VPWR.n4044 VPWR.n4043 4.6505
R6839 VPWR.n4046 VPWR.n4045 4.6505
R6840 VPWR.n4048 VPWR.n4047 4.6505
R6841 VPWR.n4050 VPWR.n4049 4.6505
R6842 VPWR.n4052 VPWR.n4051 4.6505
R6843 VPWR.n4056 VPWR.n4055 4.6505
R6844 VPWR.n4057 VPWR.n2995 4.6505
R6845 VPWR.n4062 VPWR.n4061 4.6505
R6846 VPWR.n4064 VPWR.n4063 4.6505
R6847 VPWR.n4066 VPWR.n4065 4.6505
R6848 VPWR.n4070 VPWR.n4069 4.6505
R6849 VPWR.n4073 VPWR.n4072 4.6505
R6850 VPWR.n4077 VPWR.n4076 4.6505
R6851 VPWR.n4079 VPWR.n4078 4.6505
R6852 VPWR.n4081 VPWR.n4080 4.6505
R6853 VPWR.n4085 VPWR.n4084 4.6505
R6854 VPWR.n4135 VPWR.n4134 4.6505
R6855 VPWR.n3990 VPWR.n3989 4.6505
R6856 VPWR.n3073 VPWR.n3072 4.6505
R6857 VPWR.n3071 VPWR.n3060 4.6505
R6858 VPWR.n3882 VPWR.n3881 4.6505
R6859 VPWR.n3885 VPWR.n3884 4.6505
R6860 VPWR.n3889 VPWR.n3888 4.6505
R6861 VPWR.n3891 VPWR.n3890 4.6505
R6862 VPWR.n3895 VPWR.n3894 4.6505
R6863 VPWR.n3898 VPWR.n3897 4.6505
R6864 VPWR.n3902 VPWR.n3901 4.6505
R6865 VPWR.n3905 VPWR.n3904 4.6505
R6866 VPWR.n3914 VPWR.n3913 4.6505
R6867 VPWR.n3920 VPWR.n3919 4.6505
R6868 VPWR.n3922 VPWR.n3921 4.6505
R6869 VPWR.n3090 VPWR.n3089 4.6505
R6870 VPWR.n3088 VPWR.n3087 4.6505
R6871 VPWR.n3086 VPWR.n3048 4.6505
R6872 VPWR.n3083 VPWR.n3082 4.6505
R6873 VPWR.n3081 VPWR.n3080 4.6505
R6874 VPWR.n3078 VPWR.n3077 4.6505
R6875 VPWR.n3210 VPWR.n3209 4.6505
R6876 VPWR.n3207 VPWR.n3206 4.6505
R6877 VPWR.n3205 VPWR.n3204 4.6505
R6878 VPWR.n3203 VPWR.n3202 4.6505
R6879 VPWR.n3200 VPWR.n3199 4.6505
R6880 VPWR.n3197 VPWR.n3196 4.6505
R6881 VPWR.n3195 VPWR.n3194 4.6505
R6882 VPWR.n3193 VPWR.n3192 4.6505
R6883 VPWR.n3190 VPWR.n3189 4.6505
R6884 VPWR.n3188 VPWR.n3187 4.6505
R6885 VPWR.n3186 VPWR.n3185 4.6505
R6886 VPWR.n3184 VPWR.n3183 4.6505
R6887 VPWR.n3182 VPWR.n3181 4.6505
R6888 VPWR.n3180 VPWR.n3179 4.6505
R6889 VPWR.n3176 VPWR.n3175 4.6505
R6890 VPWR.n3172 VPWR.n3154 4.6505
R6891 VPWR.n3170 VPWR.n3169 4.6505
R6892 VPWR.n3168 VPWR.n3167 4.6505
R6893 VPWR.n3166 VPWR.n3165 4.6505
R6894 VPWR.n3162 VPWR.n3040 4.6505
R6895 VPWR.n3876 VPWR.n3875 4.6505
R6896 VPWR.n3872 VPWR.n3871 4.6505
R6897 VPWR.n3232 VPWR.n3231 4.6505
R6898 VPWR.n3230 VPWR.n3229 4.6505
R6899 VPWR.n3228 VPWR.n3227 4.6505
R6900 VPWR.n3225 VPWR.n3224 4.6505
R6901 VPWR.n3223 VPWR.n3222 4.6505
R6902 VPWR.n3221 VPWR.n3220 4.6505
R6903 VPWR.n3217 VPWR.n3216 4.6505
R6904 VPWR.n3253 VPWR.n3252 4.6505
R6905 VPWR.n3257 VPWR.n3256 4.6505
R6906 VPWR.n3263 VPWR.n3234 4.6505
R6907 VPWR.n3265 VPWR.n3264 4.6505
R6908 VPWR.n3270 VPWR.n3269 4.6505
R6909 VPWR.n3274 VPWR.n3273 4.6505
R6910 VPWR.n3285 VPWR.n3284 4.6505
R6911 VPWR.n3289 VPWR.n3288 4.6505
R6912 VPWR.n3291 VPWR.n3290 4.6505
R6913 VPWR.n7163 VPWR.n7160 4.6505
R6914 VPWR.n7060 VPWR.n7059 4.6505
R6915 VPWR.n7065 VPWR.n7064 4.6505
R6916 VPWR.n7108 VPWR.n7107 4.6505
R6917 VPWR.n7116 VPWR.n7115 4.6505
R6918 VPWR.n7125 VPWR.n7124 4.6505
R6919 VPWR.n7278 VPWR.n7129 4.6505
R6920 VPWR.n7414 VPWR.n7029 4.6505
R6921 VPWR.n7399 VPWR.n7032 4.6505
R6922 VPWR.n7396 VPWR.n7033 4.6505
R6923 VPWR.n7372 VPWR.n7371 4.6505
R6924 VPWR.n7368 VPWR.n7285 4.6505
R6925 VPWR.n7365 VPWR.n7287 4.6505
R6926 VPWR.n7353 VPWR.n7295 4.6505
R6927 VPWR.n7526 VPWR.n6940 4.6505
R6928 VPWR.n7511 VPWR.n6942 4.6505
R6929 VPWR.n7508 VPWR.n6945 4.6505
R6930 VPWR.n7470 VPWR.n7468 4.6505
R6931 VPWR.n7465 VPWR.n6953 4.6505
R6932 VPWR.n7536 VPWR.n7535 4.6505
R6933 VPWR.n7541 VPWR.n7540 4.6505
R6934 VPWR.n7546 VPWR.n7545 4.6505
R6935 VPWR.n7554 VPWR.n7553 4.6505
R6936 VPWR.n7559 VPWR.n7558 4.6505
R6937 VPWR.n7525 VPWR.n7524 4.6505
R6938 VPWR.n7523 VPWR.n7522 4.6505
R6939 VPWR.n7521 VPWR.n7520 4.6505
R6940 VPWR.n7519 VPWR.n7518 4.6505
R6941 VPWR.n7517 VPWR.n7516 4.6505
R6942 VPWR.n7515 VPWR.n7514 4.6505
R6943 VPWR.n7513 VPWR.n7512 4.6505
R6944 VPWR.n7503 VPWR.n6950 4.6505
R6945 VPWR.n7500 VPWR.n7499 4.6505
R6946 VPWR.n7498 VPWR.n7497 4.6505
R6947 VPWR.n7496 VPWR.n7495 4.6505
R6948 VPWR.n7494 VPWR.n7493 4.6505
R6949 VPWR.n7492 VPWR.n7491 4.6505
R6950 VPWR.n7490 VPWR.n7489 4.6505
R6951 VPWR.n7487 VPWR.n7486 4.6505
R6952 VPWR.n7485 VPWR.n7484 4.6505
R6953 VPWR.n7483 VPWR.n7482 4.6505
R6954 VPWR.n7481 VPWR.n7480 4.6505
R6955 VPWR.n7479 VPWR.n7478 4.6505
R6956 VPWR.n7477 VPWR.n7476 4.6505
R6957 VPWR.n7475 VPWR.n7474 4.6505
R6958 VPWR.n7460 VPWR.n7459 4.6505
R6959 VPWR.n7455 VPWR.n7454 4.6505
R6960 VPWR.n7413 VPWR.n7412 4.6505
R6961 VPWR.n7411 VPWR.n7410 4.6505
R6962 VPWR.n7409 VPWR.n7408 4.6505
R6963 VPWR.n7407 VPWR.n7406 4.6505
R6964 VPWR.n7405 VPWR.n7404 4.6505
R6965 VPWR.n7403 VPWR.n7402 4.6505
R6966 VPWR.n7393 VPWR.n7392 4.6505
R6967 VPWR.n7389 VPWR.n7388 4.6505
R6968 VPWR.n7387 VPWR.n7386 4.6505
R6969 VPWR.n7385 VPWR.n7384 4.6505
R6970 VPWR.n7383 VPWR.n7382 4.6505
R6971 VPWR.n7380 VPWR 4.6505
R6972 VPWR.n7379 VPWR.n7378 4.6505
R6973 VPWR.n7374 VPWR.n7373 4.6505
R6974 VPWR.n7360 VPWR.n7289 4.6505
R6975 VPWR.n7357 VPWR.n7356 4.6505
R6976 VPWR.n7068 VPWR.n7046 4.6505
R6977 VPWR.n7076 VPWR.n7075 4.6505
R6978 VPWR.n7080 VPWR.n7079 4.6505
R6979 VPWR.n7083 VPWR.n7082 4.6505
R6980 VPWR.n7085 VPWR.n7084 4.6505
R6981 VPWR.n7087 VPWR.n7086 4.6505
R6982 VPWR.n7089 VPWR.n7088 4.6505
R6983 VPWR.n7092 VPWR.n7091 4.6505
R6984 VPWR.n7094 VPWR.n7093 4.6505
R6985 VPWR.n7096 VPWR.n7095 4.6505
R6986 VPWR.n7098 VPWR.n7097 4.6505
R6987 VPWR.n7100 VPWR.n7099 4.6505
R6988 VPWR.n7102 VPWR.n7101 4.6505
R6989 VPWR.n7104 VPWR.n7103 4.6505
R6990 VPWR.n7106 VPWR.n7105 4.6505
R6991 VPWR.n7128 VPWR.n7047 4.6505
R6992 VPWR.n7264 VPWR.n7263 4.6505
R6993 VPWR.n7267 VPWR.n7266 4.6505
R6994 VPWR.n7272 VPWR.n7271 4.6505
R6995 VPWR.n7275 VPWR.n7274 4.6505
R6996 VPWR.n7277 VPWR.n7276 4.6505
R6997 VPWR.n7118 VPWR.n7117 4.6505
R6998 VPWR.n7113 VPWR.n7112 4.6505
R6999 VPWR.n7110 VPWR.n7109 4.6505
R7000 VPWR.n7070 VPWR.n7069 4.6505
R7001 VPWR.n7067 VPWR.n7066 4.6505
R7002 VPWR.n7062 VPWR.n7061 4.6505
R7003 VPWR.n7057 VPWR.n7056 4.6505
R7004 VPWR.n7352 VPWR.n7351 4.6505
R7005 VPWR.n7355 VPWR.n7354 4.6505
R7006 VPWR.n7362 VPWR.n7361 4.6505
R7007 VPWR.n7364 VPWR.n7363 4.6505
R7008 VPWR.n7367 VPWR.n7366 4.6505
R7009 VPWR.n7370 VPWR.n7369 4.6505
R7010 VPWR.n7395 VPWR.n7394 4.6505
R7011 VPWR.n7398 VPWR.n7397 4.6505
R7012 VPWR.n7401 VPWR.n7400 4.6505
R7013 VPWR.n7457 VPWR.n7456 4.6505
R7014 VPWR.n7458 VPWR.n6954 4.6505
R7015 VPWR.n7462 VPWR.n7461 4.6505
R7016 VPWR.n7464 VPWR.n7463 4.6505
R7017 VPWR.n7467 VPWR.n7466 4.6505
R7018 VPWR.n7472 VPWR.n7471 4.6505
R7019 VPWR.n7505 VPWR.n7504 4.6505
R7020 VPWR.n7507 VPWR.n7506 4.6505
R7021 VPWR.n7510 VPWR.n7509 4.6505
R7022 VPWR.n7534 VPWR.n7533 4.6505
R7023 VPWR.n7538 VPWR.n7537 4.6505
R7024 VPWR.n7543 VPWR.n7542 4.6505
R7025 VPWR.n7548 VPWR.n7547 4.6505
R7026 VPWR.n7550 VPWR.n7549 4.6505
R7027 VPWR.n7552 VPWR.n7551 4.6505
R7028 VPWR.n7556 VPWR.n7555 4.6505
R7029 VPWR.n7565 VPWR.n7564 4.6505
R7030 VPWR.n7569 VPWR.n7568 4.6505
R7031 VPWR.n7572 VPWR.n7571 4.6505
R7032 VPWR.n7574 VPWR.n7573 4.6505
R7033 VPWR.n7193 VPWR.n7192 4.6505
R7034 VPWR.n7191 VPWR.n7189 4.6505
R7035 VPWR.n7188 VPWR.n7187 4.6505
R7036 VPWR.n7186 VPWR.n7147 4.6505
R7037 VPWR.n7185 VPWR.n7184 4.6505
R7038 VPWR.n7183 VPWR.n7181 4.6505
R7039 VPWR.n7180 VPWR.n7179 4.6505
R7040 VPWR.n7178 VPWR.n7149 4.6505
R7041 VPWR.n7177 VPWR.n7176 4.6505
R7042 VPWR.n7175 VPWR.n7150 4.6505
R7043 VPWR.n7174 VPWR.n7173 4.6505
R7044 VPWR.n7172 VPWR.n7171 4.6505
R7045 VPWR.n7170 VPWR.n7152 4.6505
R7046 VPWR.n7169 VPWR.n7168 4.6505
R7047 VPWR.n7167 VPWR.n7154 4.6505
R7048 VPWR.n7166 VPWR.n7165 4.6505
R7049 VPWR.n7164 VPWR.n7155 4.6505
R7050 VPWR.n2278 VPWR.n2277 4.64677
R7051 VPWR.n385 VPWR.n384 4.62272
R7052 VPWR.n4117 VPWR.n4116 4.5918
R7053 VPWR.n2289 VPWR.n2288 4.57445
R7054 VPWR.n9086 VPWR.n9085 4.57427
R7055 VPWR.n8061 VPWR.n8060 4.57427
R7056 VPWR.n7997 VPWR.n7996 4.57427
R7057 VPWR.n7900 VPWR.n7872 4.57427
R7058 VPWR.n8253 VPWR.n5952 4.57427
R7059 VPWR.n8104 VPWR.n8103 4.57427
R7060 VPWR.n8573 VPWR.n8572 4.57427
R7061 VPWR.n8539 VPWR.n8538 4.57427
R7062 VPWR.n8376 VPWR.n8375 4.57427
R7063 VPWR.n1091 VPWR.n1090 4.57427
R7064 VPWR.n1058 VPWR.n1057 4.57427
R7065 VPWR.n932 VPWR.n931 4.57427
R7066 VPWR.n890 VPWR.n889 4.57427
R7067 VPWR.n5514 VPWR.n5513 4.57427
R7068 VPWR.n5564 VPWR.n5563 4.57427
R7069 VPWR.n5399 VPWR.n5398 4.57427
R7070 VPWR.n1413 VPWR.n1412 4.57427
R7071 VPWR.n5253 VPWR.n5252 4.57427
R7072 VPWR.n4663 VPWR.n4662 4.57427
R7073 VPWR.n524 VPWR.n523 4.57427
R7074 VPWR.n1748 VPWR.n1727 4.57427
R7075 VPWR.n5083 VPWR.n1855 4.57427
R7076 VPWR.n1881 VPWR.n1880 4.57427
R7077 VPWR.n5161 VPWR.n1817 4.57427
R7078 VPWR.n1813 VPWR.n1812 4.57427
R7079 VPWR.n4388 VPWR.n4387 4.57427
R7080 VPWR.n4364 VPWR.n4363 4.57427
R7081 VPWR.n2640 VPWR.n2639 4.57427
R7082 VPWR.n2665 VPWR.n2664 4.57427
R7083 VPWR.n4300 VPWR.n2787 4.57427
R7084 VPWR.n4279 VPWR.n4278 4.57427
R7085 VPWR.n3555 VPWR.n3554 4.57427
R7086 VPWR.n3572 VPWR.n3571 4.57427
R7087 VPWR.n9264 VPWR.n26 4.57427
R7088 VPWR.n7832 VPWR.n7831 4.57427
R7089 VPWR.n7854 VPWR.n7853 4.57427
R7090 VPWR.n9222 VPWR.n9221 4.57427
R7091 VPWR.n3940 VPWR.n3939 4.57427
R7092 VPWR.n3960 VPWR.n3959 4.57427
R7093 VPWR.n3832 VPWR.n3831 4.57427
R7094 VPWR.n3856 VPWR.n3855 4.57427
R7095 VPWR.n7440 VPWR.n7439 4.57427
R7096 VPWR.n7418 VPWR.n7417 4.57427
R7097 VPWR.n7350 VPWR.n7349 4.57427
R7098 VPWR.n7332 VPWR.n7331 4.57427
R7099 VPWR.n5763 VPWR.n5762 4.57412
R7100 VPWR.n8204 VPWR.n8203 4.57282
R7101 VPWR.n8595 VPWR.n8593 4.57282
R7102 VPWR.n1110 VPWR.n1109 4.57282
R7103 VPWR.n4672 VPWR.n4671 4.57282
R7104 VPWR.n7053 VPWR.n7052 4.57282
R7105 VPWR.n8006 VPWR.n8005 4.57249
R7106 VPWR.n1767 VPWR.n1766 4.57249
R7107 VPWR.n6076 VPWR.n6070 4.57193
R7108 VPWR.n8433 VPWR.n8430 4.57193
R7109 VPWR.n1298 VPWR.n1297 4.57193
R7110 VPWR.n8243 VPWR.n8242 4.57152
R7111 VPWR.n7489 VPWR.n7488 4.54926
R7112 VPWR.n7417 VPWR.n7416 4.54926
R7113 VPWR.n3831 VPWR.n3830 4.54926
R7114 VPWR.n3897 VPWR.n3896 4.54926
R7115 VPWR.n7667 VPWR.n7666 4.54926
R7116 VPWR.n8023 VPWR.n8022 4.54926
R7117 VPWR.n8028 VPWR.n8027 4.54926
R7118 VPWR.n9029 VPWR.n8978 4.54926
R7119 VPWR.n8998 VPWR.n8997 4.54926
R7120 VPWR.n9007 VPWR.n9006 4.54926
R7121 VPWR.n7940 VPWR.n7939 4.54926
R7122 VPWR.n7928 VPWR.n7927 4.54926
R7123 VPWR.n6281 VPWR.n6280 4.54926
R7124 VPWR.n8273 VPWR.n8272 4.54926
R7125 VPWR.n6715 VPWR.n6714 4.54926
R7126 VPWR.n6390 VPWR.n6389 4.54926
R7127 VPWR.n6417 VPWR.n6416 4.54926
R7128 VPWR.n5648 VPWR.n5645 4.54926
R7129 VPWR.n5623 VPWR.n5622 4.54926
R7130 VPWR.n1476 VPWR.n1475 4.54926
R7131 VPWR.n1468 VPWR.n1467 4.54926
R7132 VPWR.n1503 VPWR.n1502 4.54926
R7133 VPWR.n1319 VPWR.n1272 4.54926
R7134 VPWR.n5266 VPWR.n5265 4.54926
R7135 VPWR.n1651 VPWR.n1650 4.54926
R7136 VPWR.n2171 VPWR.n2170 4.54926
R7137 VPWR.n2161 VPWR.n2160 4.54926
R7138 VPWR.n2712 VPWR.n2711 4.54926
R7139 VPWR.n4363 VPWR.n4361 4.54926
R7140 VPWR.n2355 VPWR.n2353 4.54926
R7141 VPWR.n2349 VPWR.n2348 4.54926
R7142 VPWR.n2847 VPWR.n2846 4.54926
R7143 VPWR.n2860 VPWR.n2859 4.54926
R7144 VPWR.n3608 VPWR.n3605 4.54926
R7145 VPWR.n3714 VPWR.n3713 4.54926
R7146 VPWR.n3708 VPWR.n3707 4.54926
R7147 VPWR.n2811 VPWR.n2810 4.54926
R7148 VPWR.n3651 VPWR.n3650 4.54926
R7149 VPWR.n7091 VPWR.n7090 4.54926
R7150 VPWR.n8422 VPWR.n8421 4.53667
R7151 VPWR.n929 VPWR.n928 4.53667
R7152 VPWR.n1896 VPWR.n1895 4.52113
R7153 VPWR.n653 VPWR.n652 4.50829
R7154 VPWR.n7227 VPWR.n7194 4.50829
R7155 VPWR.n296 VPWR.n258 4.50828
R7156 VPWR.n8918 VPWR.n8917 4.50828
R7157 VPWR.n8790 VPWR.n8789 4.50828
R7158 VPWR.n5830 VPWR.n5829 4.50828
R7159 VPWR.n5757 VPWR.n5756 4.5005
R7160 VPWR.n704 VPWR.n703 4.5005
R7161 VPWR VPWR.n2489 4.5005
R7162 VPWR.n2584 VPWR.n2112 4.5005
R7163 VPWR.n4221 VPWR.n4220 4.5005
R7164 VPWR.n3750 VPWR.n3369 4.5005
R7165 VPWR.n7991 VPWR.n7990 4.49637
R7166 VPWR.n8433 VPWR.n8432 4.47034
R7167 VPWR.n1678 VPWR.n1675 4.46761
R7168 VPWR.n4640 VPWR.n4636 4.46111
R7169 VPWR.n3855 VPWR.n3854 4.44348
R7170 VPWR.n1167 VPWR.n1166 4.38907
R7171 VPWR.n758 VPWR.n756 4.38907
R7172 VPWR.n2092 VPWR.n2089 4.38907
R7173 VPWR.n2079 VPWR.n2078 4.38907
R7174 VPWR.n7531 VPWR.n7530 4.36875
R7175 VPWR.n7560 VPWR.n7527 4.36875
R7176 VPWR.n7382 VPWR.n7381 4.36875
R7177 VPWR.n7283 VPWR.n7282 4.36875
R7178 VPWR.n7293 VPWR.n7292 4.36875
R7179 VPWR.n4107 VPWR.n4106 4.36875
R7180 VPWR.n3275 VPWR.n3233 4.36875
R7181 VPWR.n9152 VPWR.n9151 4.36875
R7182 VPWR.n57 VPWR.n56 4.36875
R7183 VPWR.n9196 VPWR.n9195 4.36875
R7184 VPWR.n6063 VPWR.n6062 4.36875
R7185 VPWR.n6076 VPWR.n6075 4.36875
R7186 VPWR.n210 VPWR.n209 4.36875
R7187 VPWR.n7901 VPWR.n7900 4.36875
R7188 VPWR.n8122 VPWR.n8121 4.36875
R7189 VPWR.n5928 VPWR.n5927 4.36875
R7190 VPWR.n8629 VPWR.n8628 4.36875
R7191 VPWR.n8614 VPWR.n8613 4.36875
R7192 VPWR.n386 VPWR.n385 4.36875
R7193 VPWR.n1133 VPWR.n1132 4.36875
R7194 VPWR.n753 VPWR.n752 4.36875
R7195 VPWR.n870 VPWR.n868 4.36875
R7196 VPWR.n5463 VPWR.n5462 4.36875
R7197 VPWR.n1294 VPWR.n1293 4.36875
R7198 VPWR.n1295 VPWR.n1274 4.36875
R7199 VPWR.n1325 VPWR.n1323 4.36875
R7200 VPWR.n553 VPWR.n551 4.36875
R7201 VPWR.n1723 VPWR.n548 4.36875
R7202 VPWR.n1897 VPWR.n1896 4.36875
R7203 VPWR.n5014 VPWR.n5013 4.36875
R7204 VPWR.n1963 VPWR.n1962 4.36875
R7205 VPWR.n5137 VPWR.n5131 4.36875
R7206 VPWR.n2137 VPWR.n2136 4.36875
R7207 VPWR.n2461 VPWR.n2460 4.36875
R7208 VPWR.n2374 VPWR.n2373 4.36875
R7209 VPWR.n2055 VPWR.n2054 4.36875
R7210 VPWR.n4435 VPWR.n4434 4.36875
R7211 VPWR.n4451 VPWR.n4450 4.36875
R7212 VPWR.n4538 VPWR.n4537 4.36875
R7213 VPWR.n3504 VPWR.n3503 4.36875
R7214 VPWR.n3406 VPWR.n3405 4.36875
R7215 VPWR.n7120 VPWR.n7119 4.36875
R7216 VPWR.n7157 VPWR.n7156 4.36875
R7217 VPWR.n3052 VPWR.n3050 4.31796
R7218 VPWR.n8834 VPWR.n8833 4.31796
R7219 VPWR.n889 VPWR.n885 4.31796
R7220 VPWR.n4644 VPWR.n4643 4.29023
R7221 VPWR.n3241 VPWR.n3240 4.26717
R7222 VPWR.n6511 VPWR.n6510 4.26717
R7223 VPWR.n3080 VPWR.n3079 4.1939
R7224 VPWR.n545 VPWR 4.18512
R7225 VPWR.n870 VPWR.n869 4.16558
R7226 VPWR.n5412 VPWR.n500 4.14168
R7227 VPWR.n3737 VPWR.n3736 4.14168
R7228 VPWR.n3089 VPWR.n3043 4.12612
R7229 VPWR.n3300 VPWR.n3299 4.12612
R7230 VPWR.n7900 VPWR.n7899 4.11479
R7231 VPWR.n7996 VPWR.n7995 4.06399
R7232 VPWR.n8571 VPWR.n8570 4.06399
R7233 VPWR.n889 VPWR.n888 4.06399
R7234 VPWR.n3031 VPWR.n3030 4.02033
R7235 VPWR.n3036 VPWR.n3035 4.02033
R7236 VPWR.n4104 VPWR.n4098 4.02033
R7237 VPWR.n4104 VPWR.n4103 4.02033
R7238 VPWR.n3215 VPWR.n3149 4.02033
R7239 VPWR.n3249 VPWR.n3244 4.02033
R7240 VPWR.n3249 VPWR.n3248 4.02033
R7241 VPWR.n80 VPWR.n76 4.02033
R7242 VPWR.n80 VPWR.n79 4.02033
R7243 VPWR.n68 VPWR.n67 4.02033
R7244 VPWR.n7646 VPWR.n7642 4.02033
R7245 VPWR.n7646 VPWR.n7645 4.02033
R7246 VPWR.n7654 VPWR.n7653 4.02033
R7247 VPWR.n6043 VPWR.n6017 4.02033
R7248 VPWR.n6176 VPWR.n6167 4.02033
R7249 VPWR.n6175 VPWR.n6170 4.02033
R7250 VPWR.n6175 VPWR.n6174 4.02033
R7251 VPWR.n223 VPWR.n219 4.02033
R7252 VPWR.n223 VPWR.n222 4.02033
R7253 VPWR.n7990 VPWR.n5970 4.02033
R7254 VPWR.n6289 VPWR.n6229 4.02033
R7255 VPWR.n8881 VPWR.n8877 4.02033
R7256 VPWR.n8881 VPWR.n8880 4.02033
R7257 VPWR.n6657 VPWR.n6655 4.02033
R7258 VPWR.n8150 VPWR.n8148 4.02033
R7259 VPWR.n6595 VPWR.n6591 4.02033
R7260 VPWR.n6595 VPWR.n6594 4.02033
R7261 VPWR.n8747 VPWR.n8742 4.02033
R7262 VPWR.n8747 VPWR.n8746 4.02033
R7263 VPWR.n8425 VPWR.n5876 4.02033
R7264 VPWR.n8675 VPWR.n8618 4.02033
R7265 VPWR.n6499 VPWR.n6494 4.02033
R7266 VPWR.n6499 VPWR.n6498 4.02033
R7267 VPWR.n6489 VPWR.n6487 4.02033
R7268 VPWR.n5792 VPWR.n5788 4.02033
R7269 VPWR.n5792 VPWR.n5791 4.02033
R7270 VPWR.n731 VPWR.n729 4.02033
R7271 VPWR.n806 VPWR.n803 4.02033
R7272 VPWR.n609 VPWR.n605 4.02033
R7273 VPWR.n609 VPWR.n608 4.02033
R7274 VPWR.n600 VPWR.n598 4.02033
R7275 VPWR.n419 VPWR.n415 4.02033
R7276 VPWR.n419 VPWR.n418 4.02033
R7277 VPWR.n1283 VPWR.n1279 4.02033
R7278 VPWR.n1283 VPWR.n1282 4.02033
R7279 VPWR.n1291 VPWR.n1290 4.02033
R7280 VPWR.n4801 VPWR.n4796 4.02033
R7281 VPWR.n4801 VPWR.n4800 4.02033
R7282 VPWR.n1553 VPWR.n1548 4.02033
R7283 VPWR.n1553 VPWR.n1552 4.02033
R7284 VPWR.n533 VPWR.n532 4.02033
R7285 VPWR.n1931 VPWR.n1907 4.02033
R7286 VPWR.n4929 VPWR.n4924 4.02033
R7287 VPWR.n4929 VPWR.n4928 4.02033
R7288 VPWR.n5115 VPWR.n1843 4.02033
R7289 VPWR.n2120 VPWR.n2119 4.02033
R7290 VPWR.n2440 VPWR.n2436 4.02033
R7291 VPWR.n2440 VPWR.n2439 4.02033
R7292 VPWR.n2222 VPWR.n2217 4.02033
R7293 VPWR.n2222 VPWR.n2221 4.02033
R7294 VPWR.n2016 VPWR.n2015 4.02033
R7295 VPWR.n2031 VPWR.n2030 4.02033
R7296 VPWR.n2696 VPWR.n2026 4.02033
R7297 VPWR.n4414 VPWR.n2012 4.02033
R7298 VPWR.n4503 VPWR.n4499 4.02033
R7299 VPWR.n4503 VPWR.n4502 4.02033
R7300 VPWR.n2897 VPWR.n2892 4.02033
R7301 VPWR.n2897 VPWR.n2896 4.02033
R7302 VPWR.n3378 VPWR.n3374 4.02033
R7303 VPWR.n3378 VPWR.n3377 4.02033
R7304 VPWR.n3386 VPWR.n3385 4.02033
R7305 VPWR.n3691 VPWR.n3512 4.02033
R7306 VPWR.n1585 VPWR.n1584 4.0132
R7307 VPWR.n3423 VPWR.n3422 4.0132
R7308 VPWR.n112 VPWR.n111 3.9624
R7309 VPWR.n4538 VPWR.n4484 3.9624
R7310 VPWR.n5946 VPWR.n5945 3.91455
R7311 VPWR.n4789 VPWR.n4788 3.91455
R7312 VPWR.n4025 VPWR.n2997 3.91379
R7313 VPWR.n2480 VPWR.n2479 3.91161
R7314 VPWR.n1024 VPWR.n1022 3.8558
R7315 VPWR.n765 VPWR.n764 3.81002
R7316 VPWR.n4029 VPWR.n4028 3.78037
R7317 VPWR.n3638 VPWR.n3637 3.78037
R7318 VPWR.n96 VPWR.n95 3.76521
R7319 VPWR.n245 VPWR.n244 3.76521
R7320 VPWR.n8912 VPWR.n8911 3.76521
R7321 VPWR.n8321 VPWR.n8320 3.76521
R7322 VPWR.n5818 VPWR.n5780 3.76521
R7323 VPWR.n1435 VPWR.n1434 3.76521
R7324 VPWR.n4952 VPWR.n4951 3.76521
R7325 VPWR.n2149 VPWR.n2147 3.76521
R7326 VPWR.n2449 VPWR.n2430 3.76521
R7327 VPWR.n3681 VPWR.n3680 3.76521
R7328 VPWR.n6561 VPWR 3.75923
R7329 VPWR.n5136 VPWR.n5135 3.75923
R7330 VPWR.n4068 VPWR.n4067 3.7583
R7331 VPWR.n7330 VPWR.n7329 3.70844
R7332 VPWR.n7949 VPWR.n7948 3.70298
R7333 VPWR.n5252 VPWR.n5251 3.70298
R7334 VPWR.n2838 VPWR.n2837 3.70298
R7335 VPWR.n3648 VPWR.n3647 3.70298
R7336 VPWR.n3637 VPWR.n3635 3.69446
R7337 VPWR.n3908 VPWR.n3027 3.66983
R7338 VPWR.n7766 VPWR.n7757 3.66983
R7339 VPWR.n6264 VPWR.n6263 3.66983
R7340 VPWR.n6645 VPWR.n6644 3.66983
R7341 VPWR.n2131 VPWR.n2130 3.6578
R7342 VPWR.n1171 VPWR.n1170 3.65764
R7343 VPWR.n3034 VPWR.n3033 3.65009
R7344 VPWR.n6291 VPWR.n6290 3.65009
R7345 VPWR.n5451 VPWR.n5450 3.61789
R7346 VPWR.n3903 VPWR.n3027 3.59719
R7347 VPWR.n6706 VPWR.n6705 3.59719
R7348 VPWR.n2729 VPWR.n2728 3.59719
R7349 VPWR.n8987 VPWR.n8985 3.59382
R7350 VPWR.n1488 VPWR.n1487 3.59382
R7351 VPWR.n3068 VPWR.n3067 3.57776
R7352 VPWR.n6189 VPWR.n6157 3.57776
R7353 VPWR.n7530 VPWR.n7529 3.50526
R7354 VPWR.n7561 VPWR.n7560 3.50526
R7355 VPWR.n3276 VPWR.n3275 3.50526
R7356 VPWR.n7121 VPWR.n7120 3.50526
R7357 VPWR.n7158 VPWR.n7157 3.50526
R7358 VPWR.n1126 VPWR.n1125 3.5042
R7359 VPWR.n2469 VPWR.n2423 3.5042
R7360 VPWR.n1837 VPWR.n1836 3.47876
R7361 VPWR.n6757 VPWR.n6756 3.47425
R7362 VPWR.n8483 VPWR.n8482 3.47425
R7363 VPWR.n454 VPWR.n453 3.47425
R7364 VPWR.n489 VPWR.n488 3.47425
R7365 VPWR.n2019 VPWR.n2018 3.47425
R7366 VPWR.n2827 VPWR.n2826 3.47425
R7367 VPWR.n4530 VPWR.n4528 3.43649
R7368 VPWR.n4644 VPWR.n4635 3.42615
R7369 VPWR.n6884 VPWR.n6883 3.4105
R7370 VPWR.n9072 VPWR.n9071 3.4105
R7371 VPWR.n296 VPWR.n295 3.4105
R7372 VPWR.n7961 VPWR.n7960 3.4105
R7373 VPWR.n7967 VPWR.n7966 3.4105
R7374 VPWR.n8208 VPWR.n8207 3.4105
R7375 VPWR.n8236 VPWR.n8235 3.4105
R7376 VPWR.n8102 VPWR.n5955 3.4105
R7377 VPWR.n8919 VPWR.n8918 3.4105
R7378 VPWR.n8588 VPWR.n8587 3.4105
R7379 VPWR.n8525 VPWR.n8524 3.4105
R7380 VPWR.n8541 VPWR.n8540 3.4105
R7381 VPWR VPWR.n8555 3.4105
R7382 VPWR.n8791 VPWR.n8790 3.4105
R7383 VPWR.n8721 VPWR.n8720 3.4105
R7384 VPWR.n8801 VPWR.n8800 3.4105
R7385 VPWR.n6465 VPWR.n6464 3.4105
R7386 VPWR.n6434 VPWR.n6433 3.4105
R7387 VPWR.n8377 VPWR.n8367 3.4105
R7388 VPWR.n701 VPWR.n700 3.4105
R7389 VPWR.n1106 VPWR.n1105 3.4105
R7390 VPWR.n1051 VPWR.n1050 3.4105
R7391 VPWR.n1060 VPWR.n1059 3.4105
R7392 VPWR.n5831 VPWR.n5830 3.4105
R7393 VPWR.n5739 VPWR.n381 3.4105
R7394 VPWR.n1230 VPWR.n1229 3.4105
R7395 VPWR.n911 VPWR.n910 3.4105
R7396 VPWR.n926 VPWR.n766 3.4105
R7397 VPWR.n5392 VPWR.n5391 3.4105
R7398 VPWR.n1629 VPWR.n1628 3.4105
R7399 VPWR.n5245 VPWR.n5244 3.4105
R7400 VPWR.n4653 VPWR.n4652 3.4105
R7401 VPWR.n1763 VPWR.n1762 3.4105
R7402 VPWR.n5041 VPWR.n5040 3.4105
R7403 VPWR.n2488 VPWR.n2485 3.4105
R7404 VPWR.n2590 VPWR.n2589 3.4105
R7405 VPWR.n5177 VPWR.n5176 3.4105
R7406 VPWR.n2400 VPWR.n2399 3.4105
R7407 VPWR.n2671 VPWR.n2670 3.4105
R7408 VPWR.n3483 VPWR.n3482 3.4105
R7409 VPWR.n2958 VPWR.n2957 3.4105
R7410 VPWR.n3752 VPWR.n3751 3.4105
R7411 VPWR.n9214 VPWR.n9213 3.4105
R7412 VPWR.n7705 VPWR.n7704 3.4105
R7413 VPWR.n3980 VPWR.n3979 3.4105
R7414 VPWR.n7227 VPWR.n7226 3.4105
R7415 VPWR.n9289 VPWR.n9288 3.4105
R7416 VPWR.n48 VPWR.n47 3.40367
R7417 VPWR.n5403 VPWR.n5402 3.38874
R7418 VPWR.n5289 VPWR.n1779 3.38874
R7419 VPWR.n2550 VPWR.n2549 3.38874
R7420 VPWR.n3179 VPWR.n3178 3.38562
R7421 VPWR.n5648 VPWR.n5647 3.38562
R7422 VPWR.n3201 VPWR.n3200 3.37141
R7423 VPWR.n1687 VPWR.n1684 3.37141
R7424 VPWR.t1835 VPWR.t237 3.35739
R7425 VPWR.t1827 VPWR.t1348 3.35739
R7426 VPWR.t1296 VPWR.t534 3.35739
R7427 VPWR.t782 VPWR.t2496 3.35739
R7428 VPWR.t1350 VPWR.t1549 3.35739
R7429 VPWR.t344 VPWR.t1787 3.35739
R7430 VPWR.t63 VPWR.t2108 3.35739
R7431 VPWR.t1687 VPWR.t900 3.35739
R7432 VPWR.t1175 VPWR.t2682 3.35739
R7433 VPWR.t2525 VPWR.t677 3.35739
R7434 VPWR.t509 VPWR.t2721 3.35739
R7435 VPWR.t1860 VPWR.t110 3.35739
R7436 VPWR.t808 VPWR 3.35739
R7437 VPWR.t1305 VPWR.t2535 3.35739
R7438 VPWR.t2142 VPWR.t2171 3.35739
R7439 VPWR.t460 VPWR.t1759 3.35739
R7440 VPWR.t336 VPWR.t1000 3.35739
R7441 VPWR.t874 VPWR.t2224 3.35739
R7442 VPWR.t1761 VPWR.t246 3.35739
R7443 VPWR.n1163 VPWR.n1162 3.29193
R7444 VPWR.n2829 VPWR.n2795 3.27977
R7445 VPWR.n3064 VPWR.n3063 3.25799
R7446 VPWR.n7678 VPWR.n7677 3.25799
R7447 VPWR.n6191 VPWR.n6190 3.25799
R7448 VPWR.n3047 VPWR.n3046 3.2477
R7449 VPWR.n8484 VPWR.n8483 3.2477
R7450 VPWR.n455 VPWR.n454 3.2477
R7451 VPWR.n490 VPWR.n489 3.2477
R7452 VPWR.n2020 VPWR.n2019 3.2477
R7453 VPWR.n4532 VPWR.n4531 3.2477
R7454 VPWR.n2828 VPWR.n2827 3.2477
R7455 VPWR.n8443 VPWR.n8440 3.23
R7456 VPWR.n1306 VPWR.n1304 3.21361
R7457 VPWR.n4108 VPWR.n4094 3.2005
R7458 VPWR.n9140 VPWR.n9139 3.2005
R7459 VPWR.n8445 VPWR.n8439 3.2005
R7460 VPWR.n8443 VPWR.n8442 3.2005
R7461 VPWR.n9001 VPWR.n9000 3.17405
R7462 VPWR.n7933 VPWR.n7932 3.17405
R7463 VPWR.n1473 VPWR.n1472 3.17405
R7464 VPWR.n2166 VPWR.n2165 3.17405
R7465 VPWR.n2355 VPWR.n2354 3.17405
R7466 VPWR.n2854 VPWR.n2853 3.17405
R7467 VPWR.n4254 VPWR.n4253 3.17405
R7468 VPWR.n7035 VPWR.n7034 3.16454
R7469 VPWR.n8864 VPWR.n8863 3.14971
R7470 VPWR.n811 VPWR.n810 3.14971
R7471 VPWR.n3583 VPWR.n3582 3.14971
R7472 VPWR.n3630 VPWR.n3629 3.14971
R7473 VPWR.n1836 VPWR.n1835 3.13093
R7474 VPWR.n4065 VPWR.n2993 3.12116
R7475 VPWR.n3059 VPWR.n3058 3.12116
R7476 VPWR.n6277 VPWR.n6276 3.12116
R7477 VPWR.n8299 VPWR.n8297 3.12116
R7478 VPWR.n1446 VPWR.n1445 3.12116
R7479 VPWR.n4640 VPWR.n4637 3.10638
R7480 VPWR.n6441 VPWR.n6440 3.09667
R7481 VPWR.n6696 VPWR.n6695 3.06827
R7482 VPWR.n2182 VPWR.n2181 3.06827
R7483 VPWR.n1078 VPWR.n1041 3.06326
R7484 VPWR.n9064 VPWR.n9063 3.05891
R7485 VPWR.n3404 VPWR.n3403 3.04812
R7486 VPWR.n4031 VPWR.n4030 3.01588
R7487 VPWR.n4084 VPWR.n4083 3.01588
R7488 VPWR.n9092 VPWR.n9091 3.0005
R7489 VPWR.n7983 VPWR.n7982 3.0005
R7490 VPWR.n8935 VPWR.n8934 3.0005
R7491 VPWR.n6564 VPWR.n6563 3.0005
R7492 VPWR.n8554 VPWR.n8515 3.0005
R7493 VPWR.n8394 VPWR.n8393 3.0005
R7494 VPWR.n5845 VPWR.n5844 3.0005
R7495 VPWR.n1075 VPWR.n1074 3.0005
R7496 VPWR.n691 VPWR.n690 3.0005
R7497 VPWR.n900 VPWR.n899 3.0005
R7498 VPWR.n5557 VPWR.n5556 3.0005
R7499 VPWR.n1404 VPWR.n1403 3.0005
R7500 VPWR.n4656 VPWR.n4655 3.0005
R7501 VPWR.n5067 VPWR.n5066 3.0005
R7502 VPWR.n2524 VPWR.n2523 3.0005
R7503 VPWR.n2947 VPWR.n2946 3.0005
R7504 VPWR.n9251 VPWR.n9250 3.0005
R7505 VPWR.n7298 VPWR.n7297 2.99733
R7506 VPWR.n9202 VPWR.n9200 2.99733
R7507 VPWR.n7996 VPWR.n7992 2.99733
R7508 VPWR.n8833 VPWR.n338 2.99733
R7509 VPWR.n8429 VPWR.n5868 2.99733
R7510 VPWR.n5440 VPWR.n496 2.99733
R7511 VPWR.n2376 VPWR.n2297 2.99733
R7512 VPWR.n7685 VPWR.n7684 2.98339
R7513 VPWR.n6198 VPWR.n6197 2.98339
R7514 VPWR.n8373 VPWR.n8372 2.98339
R7515 VPWR.n7601 VPWR.n7600 2.96248
R7516 VPWR.n3320 VPWR.n3319 2.96248
R7517 VPWR.n6381 VPWR.n6376 2.96248
R7518 VPWR.n1671 VPWR.n1669 2.96248
R7519 VPWR.n4841 VPWR.n4840 2.94563
R7520 VPWR.n2934 VPWR.n2933 2.94563
R7521 VPWR.n7760 VPWR.n6126 2.92182
R7522 VPWR.n6240 VPWR.n6239 2.92182
R7523 VPWR.n3068 VPWR.n3064 2.91308
R7524 VPWR.n7677 VPWR.n7676 2.91308
R7525 VPWR.n6190 VPWR.n6189 2.91308
R7526 VPWR.n3071 VPWR.n3061 2.87861
R7527 VPWR.n9139 VPWR.n9135 2.87861
R7528 VPWR.n9204 VPWR.n9203 2.87861
R7529 VPWR.n198 VPWR.n197 2.87861
R7530 VPWR.n6186 VPWR.n6161 2.87861
R7531 VPWR.n8116 VPWR.n8115 2.87861
R7532 VPWR.n6671 VPWR.n6668 2.87861
R7533 VPWR.n8626 VPWR.n8624 2.87861
R7534 VPWR.n5872 VPWR.n5871 2.87861
R7535 VPWR.n6364 VPWR.n6363 2.87861
R7536 VPWR.n825 VPWR.n824 2.87861
R7537 VPWR.n816 VPWR.n815 2.87861
R7538 VPWR.n438 VPWR.n406 2.87861
R7539 VPWR.n469 VPWR.n467 2.87861
R7540 VPWR.n499 VPWR.n498 2.87861
R7541 VPWR.n1543 VPWR.n1541 2.87861
R7542 VPWR.n5006 VPWR.n5005 2.87861
R7543 VPWR.n1951 VPWR.n1904 2.87861
R7544 VPWR.n2295 VPWR.n2293 2.87861
R7545 VPWR.n1998 VPWR.n1997 2.87861
R7546 VPWR.n5943 VPWR.n5942 2.84494
R7547 VPWR.n2004 VPWR.n2003 2.84494
R7548 VPWR.n8968 VPWR.n8967 2.79415
R7549 VPWR.n7039 VPWR.n7038 2.76904
R7550 VPWR.n3958 VPWR.n3957 2.75684
R7551 VPWR.n6013 VPWR.n6012 2.75091
R7552 VPWR.n2993 VPWR.n2992 2.71052
R7553 VPWR.n3149 VPWR.n3148 2.71052
R7554 VPWR.n3058 VPWR.n3057 2.71052
R7555 VPWR.n3030 VPWR.n3029 2.71052
R7556 VPWR.n4098 VPWR.n4097 2.71052
R7557 VPWR.n4103 VPWR.n4102 2.71052
R7558 VPWR.n3244 VPWR.n3243 2.71052
R7559 VPWR.n3248 VPWR.n3247 2.71052
R7560 VPWR.n76 VPWR.n75 2.71052
R7561 VPWR.n79 VPWR.n78 2.71052
R7562 VPWR.n67 VPWR.n66 2.71052
R7563 VPWR.n7642 VPWR.n7641 2.71052
R7564 VPWR.n7645 VPWR.n7644 2.71052
R7565 VPWR.n7653 VPWR.n7652 2.71052
R7566 VPWR.n6017 VPWR.n6016 2.71052
R7567 VPWR.n6276 VPWR.n6275 2.71052
R7568 VPWR.n6167 VPWR.n6166 2.71052
R7569 VPWR.n6170 VPWR.n6169 2.71052
R7570 VPWR.n6174 VPWR.n6173 2.71052
R7571 VPWR.n219 VPWR.n218 2.71052
R7572 VPWR.n222 VPWR.n221 2.71052
R7573 VPWR.n8297 VPWR.n8296 2.71052
R7574 VPWR.n8877 VPWR.n8876 2.71052
R7575 VPWR.n8880 VPWR.n8879 2.71052
R7576 VPWR.n6655 VPWR.n6654 2.71052
R7577 VPWR.n8148 VPWR.n8147 2.71052
R7578 VPWR.n6591 VPWR.n6590 2.71052
R7579 VPWR.n6594 VPWR.n6593 2.71052
R7580 VPWR.n8742 VPWR.n8741 2.71052
R7581 VPWR.n8746 VPWR.n8745 2.71052
R7582 VPWR.n5876 VPWR.n5875 2.71052
R7583 VPWR.n8618 VPWR.n8617 2.71052
R7584 VPWR.n6494 VPWR.n6493 2.71052
R7585 VPWR.n6498 VPWR.n6497 2.71052
R7586 VPWR.n6487 VPWR.n6486 2.71052
R7587 VPWR.n5788 VPWR.n5787 2.71052
R7588 VPWR.n5791 VPWR.n5790 2.71052
R7589 VPWR.n729 VPWR.n728 2.71052
R7590 VPWR.n803 VPWR.n802 2.71052
R7591 VPWR.n605 VPWR.n604 2.71052
R7592 VPWR.n608 VPWR.n607 2.71052
R7593 VPWR.n598 VPWR.n597 2.71052
R7594 VPWR.n1445 VPWR.n1444 2.71052
R7595 VPWR.n415 VPWR.n414 2.71052
R7596 VPWR.n418 VPWR.n417 2.71052
R7597 VPWR.n1279 VPWR.n1278 2.71052
R7598 VPWR.n1282 VPWR.n1281 2.71052
R7599 VPWR.n1290 VPWR.n1289 2.71052
R7600 VPWR.n4796 VPWR.n4795 2.71052
R7601 VPWR.n4800 VPWR.n4799 2.71052
R7602 VPWR.n1548 VPWR.n1547 2.71052
R7603 VPWR.n1552 VPWR.n1551 2.71052
R7604 VPWR.n532 VPWR.n531 2.71052
R7605 VPWR.n1907 VPWR.n1906 2.71052
R7606 VPWR.n4924 VPWR.n4923 2.71052
R7607 VPWR.n4928 VPWR.n4927 2.71052
R7608 VPWR.n1843 VPWR.n1842 2.71052
R7609 VPWR.n2119 VPWR.n2118 2.71052
R7610 VPWR.n2436 VPWR.n2435 2.71052
R7611 VPWR.n2439 VPWR.n2438 2.71052
R7612 VPWR.n2217 VPWR.n2216 2.71052
R7613 VPWR.n2221 VPWR.n2220 2.71052
R7614 VPWR.n2015 VPWR.n2014 2.71052
R7615 VPWR.n2030 VPWR.n2029 2.71052
R7616 VPWR.n2026 VPWR.n2025 2.71052
R7617 VPWR.n2012 VPWR.n2011 2.71052
R7618 VPWR.n4499 VPWR.n4498 2.71052
R7619 VPWR.n4502 VPWR.n4501 2.71052
R7620 VPWR.n2892 VPWR.n2891 2.71052
R7621 VPWR.n2896 VPWR.n2895 2.71052
R7622 VPWR.n3374 VPWR.n3373 2.71052
R7623 VPWR.n3377 VPWR.n3376 2.71052
R7624 VPWR.n3385 VPWR.n3384 2.71052
R7625 VPWR.n3512 VPWR.n3511 2.71052
R7626 VPWR.n7763 VPWR.n7762 2.65275
R7627 VPWR.n6238 VPWR.n6235 2.65275
R7628 VPWR.n3192 VPWR.n3191 2.64665
R7629 VPWR.n4041 VPWR.n4040 2.64665
R7630 VPWR.n4084 VPWR.n4082 2.64665
R7631 VPWR.n7745 VPWR.n7744 2.64665
R7632 VPWR.n7776 VPWR.n7775 2.64665
R7633 VPWR.n7802 VPWR.n7801 2.64665
R7634 VPWR.n7831 VPWR.n7830 2.64665
R7635 VPWR.n6006 VPWR.n6005 2.64665
R7636 VPWR.n6246 VPWR.n6245 2.64665
R7637 VPWR.n6305 VPWR.n6304 2.64665
R7638 VPWR.n6773 VPWR.n6772 2.64665
R7639 VPWR.n1695 VPWR.n1694 2.64665
R7640 VPWR.n2913 VPWR.n2912 2.64665
R7641 VPWR.n6712 VPWR.n6711 2.64513
R7642 VPWR.n6627 VPWR.n6626 2.64513
R7643 VPWR.n3273 VPWR.n3272 2.63579
R7644 VPWR.n5777 VPWR.n5776 2.63579
R7645 VPWR.n4460 VPWR.n4459 2.63579
R7646 VPWR.n3066 VPWR.n3065 2.61352
R7647 VPWR.n9134 VPWR.n9133 2.61352
R7648 VPWR.n9202 VPWR.n9201 2.61352
R7649 VPWR.n8967 VPWR.n8966 2.61352
R7650 VPWR.n6160 VPWR.n6159 2.61352
R7651 VPWR.n338 VPWR.n337 2.61352
R7652 VPWR.n6667 VPWR.n6666 2.61352
R7653 VPWR.n8623 VPWR.n8622 2.61352
R7654 VPWR.n5868 VPWR.n5867 2.61352
R7655 VPWR.n6362 VPWR.n6361 2.61352
R7656 VPWR.n823 VPWR.n822 2.61352
R7657 VPWR.n814 VPWR.n813 2.61352
R7658 VPWR.n405 VPWR.n404 2.61352
R7659 VPWR.n466 VPWR.n465 2.61352
R7660 VPWR.n496 VPWR.n495 2.61352
R7661 VPWR.n1540 VPWR.n1539 2.61352
R7662 VPWR.n5004 VPWR.n5003 2.61352
R7663 VPWR.n1903 VPWR.n1902 2.61352
R7664 VPWR.n2297 VPWR.n2296 2.61352
R7665 VPWR.n1996 VPWR.n1995 2.61352
R7666 VPWR.n2563 VPWR.n2562 2.54018
R7667 VPWR.n3287 VPWR.n3286 2.53934
R7668 VPWR.n8016 VPWR.n8015 2.53934
R7669 VPWR.n2700 VPWR.n2699 2.53934
R7670 VPWR.n3506 VPWR.n3505 2.53934
R7671 VPWR.n4012 VPWR.n4011 2.50603
R7672 VPWR.n6062 VPWR.n6061 2.48939
R7673 VPWR.n8121 VPWR.n8120 2.48939
R7674 VPWR.n8613 VPWR.n8612 2.4386
R7675 VPWR.n4434 VPWR.n4433 2.4386
R7676 VPWR.n2709 VPWR.n2708 2.43356
R7677 VPWR.n5473 VPWR.n5472 2.4268
R7678 VPWR.n1678 VPWR.n1677 2.40784
R7679 VPWR.n5442 VPWR.n494 2.3878
R7680 VPWR.n8985 VPWR.n8984 2.38473
R7681 VPWR.n1489 VPWR.n1488 2.38473
R7682 VPWR.n5449 VPWR.n5448 2.34574
R7683 VPWR.n6948 VPWR.n6947 2.33701
R7684 VPWR.n7043 VPWR.n7042 2.33701
R7685 VPWR.n7291 VPWR.n7290 2.33701
R7686 VPWR.n3238 VPWR.n3237 2.33701
R7687 VPWR.n61 VPWR.n60 2.33701
R7688 VPWR.n45 VPWR.n44 2.33701
R7689 VPWR.n40 VPWR.n39 2.33701
R7690 VPWR.n6069 VPWR.n6068 2.33701
R7691 VPWR.n8866 VPWR.n8865 2.33701
R7692 VPWR.n5940 VPWR.n5939 2.33701
R7693 VPWR.n8195 VPWR.n8194 2.33701
R7694 VPWR.n6508 VPWR.n6507 2.33701
R7695 VPWR.n383 VPWR.n382 2.33701
R7696 VPWR.n1130 VPWR.n724 2.33701
R7697 VPWR.n751 VPWR.n750 2.33701
R7698 VPWR.n645 VPWR.n644 2.33701
R7699 VPWR.n5460 VPWR.n5459 2.33701
R7700 VPWR.n4918 VPWR.n4917 2.33701
R7701 VPWR.n2128 VPWR.n2127 2.33701
R7702 VPWR.n2129 VPWR.n2128 2.33701
R7703 VPWR.n2561 VPWR.n2188 2.33701
R7704 VPWR.n2459 VPWR.n2458 2.33701
R7705 VPWR.n2468 VPWR.n2467 2.33701
R7706 VPWR.n2475 VPWR.n2474 2.33701
R7707 VPWR.n2057 VPWR.n2056 2.33701
R7708 VPWR.n3502 VPWR.n3501 2.33701
R7709 VPWR.n3403 VPWR.n3402 2.33701
R7710 VPWR.n7073 VPWR.n7072 2.33701
R7711 VPWR.n5970 VPWR.n5969 2.32777
R7712 VPWR.n6734 VPWR.n6733 2.32777
R7713 VPWR.n6263 VPWR.n6262 2.29662
R7714 VPWR.n6186 VPWR.n6185 2.29662
R7715 VPWR.n6187 VPWR.n6186 2.29662
R7716 VPWR.n6762 VPWR.n6645 2.29662
R7717 VPWR.n6692 VPWR.n6657 2.29662
R7718 VPWR.n1326 VPWR.n1325 2.29662
R7719 VPWR.n4711 VPWR.n4642 2.29662
R7720 VPWR.n1951 VPWR.n1950 2.29662
R7721 VPWR.n1952 VPWR.n1951 2.29662
R7722 VPWR.n2696 VPWR.n2023 2.29662
R7723 VPWR.n3637 VPWR.n3636 2.29662
R7724 VPWR.n7767 VPWR.n7766 2.29662
R7725 VPWR.n4006 VPWR.n4005 2.29662
R7726 VPWR.n4028 VPWR.n4027 2.29662
R7727 VPWR.n3908 VPWR.n3907 2.29662
R7728 VPWR.n8973 VPWR.n198 2.29643
R7729 VPWR.n6454 VPWR.n6453 2.29643
R7730 VPWR.n8425 VPWR.n5873 2.29643
R7731 VPWR.n4714 VPWR.n4713 2.29643
R7732 VPWR.n5094 VPWR.n5093 2.29643
R7733 VPWR.n1931 VPWR.n1908 2.29643
R7734 VPWR.n2045 VPWR.n2031 2.29643
R7735 VPWR.n3215 VPWR.n3211 2.29643
R7736 VPWR.n4009 VPWR.n4007 2.29615
R7737 VPWR.n2992 VPWR.n2991 2.28969
R7738 VPWR.n3057 VPWR.n3056 2.28969
R7739 VPWR.n3029 VPWR.n3028 2.28969
R7740 VPWR.n4102 VPWR.n4101 2.28969
R7741 VPWR.n4097 VPWR.n4096 2.28969
R7742 VPWR.n3148 VPWR.n3147 2.28969
R7743 VPWR.n3247 VPWR.n3246 2.28969
R7744 VPWR.n3243 VPWR.n3242 2.28969
R7745 VPWR.n78 VPWR.n77 2.28969
R7746 VPWR.n75 VPWR.n74 2.28969
R7747 VPWR.n66 VPWR.n65 2.28969
R7748 VPWR.n7644 VPWR.n7643 2.28969
R7749 VPWR.n7641 VPWR.n7640 2.28969
R7750 VPWR.n7652 VPWR.n7651 2.28969
R7751 VPWR.n6016 VPWR.n6015 2.28969
R7752 VPWR.n6275 VPWR.n6274 2.28969
R7753 VPWR.n6166 VPWR.n6165 2.28969
R7754 VPWR.n6173 VPWR.n6172 2.28969
R7755 VPWR.n6169 VPWR.n6168 2.28969
R7756 VPWR.n221 VPWR.n220 2.28969
R7757 VPWR.n218 VPWR.n217 2.28969
R7758 VPWR.n8296 VPWR.n8295 2.28969
R7759 VPWR.n8879 VPWR.n8878 2.28969
R7760 VPWR.n8876 VPWR.n8875 2.28969
R7761 VPWR.n6654 VPWR.n6653 2.28969
R7762 VPWR.n8147 VPWR.n8146 2.28969
R7763 VPWR.n6593 VPWR.n6592 2.28969
R7764 VPWR.n6590 VPWR.n6589 2.28969
R7765 VPWR.n8745 VPWR.n8744 2.28969
R7766 VPWR.n8741 VPWR.n8740 2.28969
R7767 VPWR.n5875 VPWR.n5874 2.28969
R7768 VPWR.n8617 VPWR.n8616 2.28969
R7769 VPWR.n6497 VPWR.n6496 2.28969
R7770 VPWR.n6493 VPWR.n6492 2.28969
R7771 VPWR.n6486 VPWR.n6485 2.28969
R7772 VPWR.n5790 VPWR.n5789 2.28969
R7773 VPWR.n5787 VPWR.n5786 2.28969
R7774 VPWR.n728 VPWR.n727 2.28969
R7775 VPWR.n802 VPWR.n801 2.28969
R7776 VPWR.n607 VPWR.n606 2.28969
R7777 VPWR.n604 VPWR.n603 2.28969
R7778 VPWR.n597 VPWR.n596 2.28969
R7779 VPWR.n1444 VPWR.n1443 2.28969
R7780 VPWR.n417 VPWR.n416 2.28969
R7781 VPWR.n414 VPWR.n413 2.28969
R7782 VPWR.n1281 VPWR.n1280 2.28969
R7783 VPWR.n1278 VPWR.n1277 2.28969
R7784 VPWR.n1289 VPWR.n1288 2.28969
R7785 VPWR.n4799 VPWR.n4798 2.28969
R7786 VPWR.n4795 VPWR.n4794 2.28969
R7787 VPWR.n1551 VPWR.n1550 2.28969
R7788 VPWR.n1547 VPWR.n1546 2.28969
R7789 VPWR.n531 VPWR.n530 2.28969
R7790 VPWR.n1906 VPWR.n1905 2.28969
R7791 VPWR.n4927 VPWR.n4926 2.28969
R7792 VPWR.n4923 VPWR.n4922 2.28969
R7793 VPWR.n1842 VPWR.n1841 2.28969
R7794 VPWR.n2118 VPWR.n2117 2.28969
R7795 VPWR.n2438 VPWR.n2437 2.28969
R7796 VPWR.n2435 VPWR.n2434 2.28969
R7797 VPWR.n2220 VPWR.n2219 2.28969
R7798 VPWR.n2216 VPWR.n2215 2.28969
R7799 VPWR.n2014 VPWR.n2013 2.28969
R7800 VPWR.n2029 VPWR.n2028 2.28969
R7801 VPWR.n2025 VPWR.n2024 2.28969
R7802 VPWR.n2011 VPWR.n2010 2.28969
R7803 VPWR.n4501 VPWR.n4500 2.28969
R7804 VPWR.n4498 VPWR.n4497 2.28969
R7805 VPWR.n2895 VPWR.n2894 2.28969
R7806 VPWR.n2891 VPWR.n2890 2.28969
R7807 VPWR.n3376 VPWR.n3375 2.28969
R7808 VPWR.n3373 VPWR.n3372 2.28969
R7809 VPWR.n3384 VPWR.n3383 2.28969
R7810 VPWR.n3511 VPWR.n3510 2.28969
R7811 VPWR.n8756 VPWR.n8755 2.28621
R7812 VPWR.n4111 VPWR.n4091 2.28407
R7813 VPWR.n4112 VPWR.n4111 2.28407
R7814 VPWR.n4645 VPWR.n4644 2.28374
R7815 VPWR.n6672 VPWR.n6671 2.28218
R7816 VPWR.n8390 VPWR.n5879 2.28218
R7817 VPWR.n5169 VPWR.n1815 2.28206
R7818 VPWR.n3563 VPWR.n3534 2.28206
R7819 VPWR.n9256 VPWR.n9255 2.28198
R7820 VPWR.n8705 VPWR.n351 2.28171
R7821 VPWR.n5006 VPWR.n5002 2.28171
R7822 VPWR.n707 VPWR.n587 2.28167
R7823 VPWR.n9139 VPWR.n138 2.28159
R7824 VPWR.n3903 VPWR.n3031 2.27488
R7825 VPWR.n6044 VPWR.n6043 2.27488
R7826 VPWR.n6229 VPWR.n6228 2.27488
R7827 VPWR.n4407 VPWR.n2016 2.27488
R7828 VPWR.n6608 VPWR.n6607 2.25932
R7829 VPWR.n8768 VPWR.n8734 2.25932
R7830 VPWR.n6515 VPWR.n6491 2.25932
R7831 VPWR.n5826 VPWR.n5777 2.25932
R7832 VPWR.n1143 VPWR.n1141 2.25932
R7833 VPWR.n5435 VPWR.n5434 2.25932
R7834 VPWR.n1439 VPWR.n1384 2.25932
R7835 VPWR.n1566 VPWR.n1565 2.25932
R7836 VPWR.n4745 VPWR.n4744 2.25932
R7837 VPWR.n4764 VPWR.n4648 2.25932
R7838 VPWR.n5022 VPWR.n5021 2.25932
R7839 VPWR.n5021 VPWR.n1890 2.25932
R7840 VPWR.n5028 VPWR.n5027 2.25932
R7841 VPWR.n2684 VPWR.n2682 2.25932
R7842 VPWR.n3392 VPWR.n3391 2.25932
R7843 VPWR.n6099 VPWR.n6098 2.23542
R7844 VPWR.n8157 VPWR.n8156 2.23542
R7845 VPWR.n8612 VPWR.n8611 2.23542
R7846 VPWR.n1996 VPWR.n1994 2.23542
R7847 VPWR.n5615 VPWR.n5613 2.19165
R7848 VPWR.n6061 VPWR.n6060 2.18463
R7849 VPWR.n8120 VPWR.n8119 2.18463
R7850 VPWR.n8779 VPWR.n8778 2.18463
R7851 VPWR.n8662 VPWR.n8661 2.18463
R7852 VPWR.n809 VPWR.n808 2.18463
R7853 VPWR.n4442 VPWR.n4441 2.18463
R7854 VPWR.n3581 VPWR.n3580 2.18463
R7855 VPWR.n3628 VPWR.n3627 2.18463
R7856 VPWR.n8375 VPWR.n8374 2.18453
R7857 VPWR.n7041 VPWR.n7040 2.1578
R7858 VPWR.n4641 VPWR.n4640 2.13383
R7859 VPWR.n3067 VPWR.n3066 2.12365
R7860 VPWR.n6160 VPWR.n6157 2.12365
R7861 VPWR.n8341 VPWR.n8340 2.08304
R7862 VPWR.n4094 VPWR.n4093 2.07374
R7863 VPWR.n4116 VPWR.n4114 2.07374
R7864 VPWR.n6949 VPWR.n6948 2.03225
R7865 VPWR.n7044 VPWR.n7043 2.03225
R7866 VPWR.n60 VPWR.n59 2.03225
R7867 VPWR.n41 VPWR.n40 2.03225
R7868 VPWR.n6068 VPWR.n6067 2.03225
R7869 VPWR.n8867 VPWR.n8866 2.03225
R7870 VPWR.n8196 VPWR.n8195 2.03225
R7871 VPWR.n8757 VPWR.n8756 2.03225
R7872 VPWR.n6540 VPWR.n6539 2.03225
R7873 VPWR.n725 VPWR.n724 2.03225
R7874 VPWR.n1122 VPWR.n1121 2.03225
R7875 VPWR.n5459 VPWR.n5458 2.03225
R7876 VPWR.n4919 VPWR.n4918 2.03225
R7877 VPWR.n2458 VPWR.n2457 2.03225
R7878 VPWR.n2467 VPWR.n2466 2.03225
R7879 VPWR.n2474 VPWR.n2473 2.03225
R7880 VPWR.n2058 VPWR.n2057 2.03225
R7881 VPWR.n7074 VPWR.n7073 2.03225
R7882 VPWR.n953 VPWR.n952 2.02422
R7883 VPWR.n3227 VPWR.n3226 2.01042
R7884 VPWR.n8035 VPWR.n8034 2.01042
R7885 VPWR.n8270 VPWR.n8269 2.01042
R7886 VPWR.n1648 VPWR.n1647 2.01042
R7887 VPWR.n3599 VPWR.n3598 2.01042
R7888 VPWR.n3621 VPWR.n3620 2.01042
R7889 VPWR.n3701 VPWR.n3700 2.01042
R7890 VPWR.n2806 VPWR.n2805 2.01042
R7891 VPWR.n1677 VPWR.n1676 1.99683
R7892 VPWR.n1123 VPWR.n1122 1.98145
R7893 VPWR.n5443 VPWR.n5442 1.98145
R7894 VPWR.n1604 VPWR.n1603 1.98145
R7895 VPWR.n6206 VPWR.n6205 1.93767
R7896 VPWR.n6828 VPWR.n6827 1.93767
R7897 VPWR.n6550 VPWR.n6549 1.93767
R7898 VPWR.n1333 VPWR.n1332 1.93767
R7899 VPWR.n1610 VPWR.n1609 1.93767
R7900 VPWR.n2497 VPWR.n2496 1.93767
R7901 VPWR.n2276 VPWR.n2275 1.93767
R7902 VPWR.n3446 VPWR.n3445 1.93767
R7903 VPWR.n7725 VPWR.n7724 1.93767
R7904 VPWR.n5702 VPWR.n5701 1.93767
R7905 VPWR.n4985 VPWR.n4984 1.93767
R7906 VPWR.n2967 VPWR.n2966 1.93767
R7907 VPWR.n6628 VPWR.n6627 1.90463
R7908 VPWR.n7791 VPWR.n7790 1.88295
R7909 VPWR.n3159 VPWR.n3158 1.88285
R7910 VPWR.n799 VPWR.n714 1.88285
R7911 VPWR.n617 VPWR.n615 1.88285
R7912 VPWR.n5106 VPWR.n5105 1.88285
R7913 VPWR.n3939 VPWR.n3938 1.85065
R7914 VPWR.n4783 VPWR.n4782 1.85065
R7915 VPWR.n960 VPWR.n758 1.82907
R7916 VPWR.n2564 VPWR.n2563 1.82907
R7917 VPWR.n3046 VPWR.n3045 1.81289
R7918 VPWR.n8254 VPWR.n5950 1.80429
R7919 VPWR.n8575 VPWR.n8574 1.80429
R7920 VPWR.n1093 VPWR.n1092 1.80429
R7921 VPWR.n5516 VPWR.n5515 1.80429
R7922 VPWR.n5254 VPWR.n1789 1.80429
R7923 VPWR.n5084 VPWR.n1854 1.80429
R7924 VPWR.n3934 VPWR.n3933 1.80429
R7925 VPWR.n9266 VPWR.n9265 1.80429
R7926 VPWR.n8059 VPWR.n5960 1.80429
R7927 VPWR.n4359 VPWR.n4358 1.80429
R7928 VPWR.n4302 VPWR.n4301 1.80429
R7929 VPWR.n7325 VPWR.n7324 1.80429
R7930 VPWR.n2636 VPWR.n2635 1.80353
R7931 VPWR.n7856 VPWR.n7855 1.80353
R7932 VPWR.n3573 VPWR.n3532 1.80353
R7933 VPWR.n7415 VPWR.n7028 1.80353
R7934 VPWR.n8344 VPWR.n8343 1.80347
R7935 VPWR.n5400 VPWR.n501 1.80347
R7936 VPWR.n5324 VPWR.n5323 1.80347
R7937 VPWR.n5160 VPWR.n1828 1.80347
R7938 VPWR.n3829 VPWR.n3828 1.80347
R7939 VPWR.n8457 VPWR.n8456 1.77828
R7940 VPWR.n3035 VPWR.n3034 1.74595
R7941 VPWR.n6291 VPWR.n6289 1.74595
R7942 VPWR.n8455 VPWR.n8454 1.73764
R7943 VPWR.n2018 VPWR.n2017 1.73737
R7944 VPWR.n4447 VPWR.n4446 1.72748
R7945 VPWR.n952 VPWR.n951 1.72066
R7946 VPWR.n2337 VPWR.n2336 1.68839
R7947 VPWR.n7676 VPWR.n7637 1.68673
R7948 VPWR.t1954 VPWR.t3089 1.67895
R7949 VPWR.t1958 VPWR.t3087 1.67895
R7950 VPWR.t2286 VPWR.t816 1.67895
R7951 VPWR.n8186 VPWR.t2844 1.67895
R7952 VPWR.t2482 VPWR.t2113 1.67895
R7953 VPWR.t2480 VPWR.t1825 1.67895
R7954 VPWR.t139 VPWR.t2000 1.67895
R7955 VPWR.t1538 VPWR.t1073 1.67895
R7956 VPWR.t3237 VPWR.t1814 1.67895
R7957 VPWR.t3239 VPWR.t1765 1.67895
R7958 VPWR.t2769 VPWR.t1299 1.67895
R7959 VPWR.t2771 VPWR.t1767 1.67895
R7960 VPWR.t768 VPWR.t1622 1.67895
R7961 VPWR.t2154 VPWR 1.67895
R7962 VPWR.t1063 VPWR.t1725 1.67895
R7963 VPWR.t1942 VPWR.t1065 1.67895
R7964 VPWR.t2349 VPWR.t1431 1.67895
R7965 VPWR.t1425 VPWR.t1677 1.67895
R7966 VPWR.t1730 VPWR.t2227 1.67895
R7967 VPWR.t2963 VPWR.t2907 1.67895
R7968 VPWR.n2000 VPWR.t2509 1.67895
R7969 VPWR.t1167 VPWR.t2666 1.67895
R7970 VPWR.n3674 VPWR.t988 1.67895
R7971 VPWR.n4249 VPWR.t2517 1.67895
R7972 VPWR.n6539 VPWR.n6538 1.67669
R7973 VPWR.n2555 VPWR.n2554 1.67669
R7974 VPWR.n3045 VPWR.n3044 1.66186
R7975 VPWR.n8474 VPWR.n8473 1.66186
R7976 VPWR.n4783 VPWR.n4777 1.66186
R7977 VPWR.n6126 VPWR.n6125 1.65335
R7978 VPWR.n6256 VPWR.n6240 1.65335
R7979 VPWR.n4530 VPWR.n4529 1.63881
R7980 VPWR.n55 VPWR.n54 1.6259
R7981 VPWR.n3405 VPWR.n3404 1.6259
R7982 VPWR.n3919 VPWR.n3918 1.6241
R7983 VPWR.n9058 VPWR.n9057 1.6241
R7984 VPWR.n6759 VPWR.n6758 1.6241
R7985 VPWR.n6758 VPWR.n6757 1.6241
R7986 VPWR.n6744 VPWR.n6743 1.6241
R7987 VPWR.n8471 VPWR.n8470 1.6241
R7988 VPWR.n5474 VPWR.n5473 1.6241
R7989 VPWR.n5479 VPWR.n5478 1.6241
R7990 VPWR.n4522 VPWR.n4521 1.6241
R7991 VPWR.n7793 VPWR.n7791 1.62167
R7992 VPWR.n6096 VPWR.n6095 1.52431
R7993 VPWR.n8865 VPWR.n8864 1.52431
R7994 VPWR.n8160 VPWR.n8159 1.52431
R7995 VPWR.n5942 VPWR.n5941 1.52431
R7996 VPWR.n8193 VPWR.n8192 1.52431
R7997 VPWR.n8784 VPWR.n8783 1.52431
R7998 VPWR.n8667 VPWR.n8666 1.52431
R7999 VPWR.n1582 VPWR.n1581 1.52431
R8000 VPWR.n2003 VPWR.n2002 1.52431
R8001 VPWR.n6175 VPWR.n6171 1.50646
R8002 VPWR.n6596 VPWR.n6595 1.50646
R8003 VPWR.n6499 VPWR.n6495 1.50646
R8004 VPWR.n610 VPWR.n609 1.50646
R8005 VPWR.n1286 VPWR.n1283 1.50646
R8006 VPWR.n1553 VPWR.n1549 1.50646
R8007 VPWR.n2441 VPWR.n2440 1.50646
R8008 VPWR.n2222 VPWR.n2218 1.50646
R8009 VPWR.n3381 VPWR.n3378 1.50646
R8010 VPWR.n7649 VPWR.n7646 1.50646
R8011 VPWR.n3249 VPWR.n3245 1.50646
R8012 VPWR.n4120 VPWR.n4089 1.50638
R8013 VPWR.n4064 VPWR.n2994 1.50638
R8014 VPWR.n9192 VPWR.n35 1.50638
R8015 VPWR.n8301 VPWR.n5934 1.50638
R8016 VPWR.n8599 VPWR.n8598 1.50638
R8017 VPWR.n8676 VPWR.n355 1.50638
R8018 VPWR.n998 VPWR.n995 1.50638
R8019 VPWR.n4694 VPWR.n4693 1.50638
R8020 VPWR.n2236 VPWR.n2235 1.50638
R8021 VPWR.n2302 VPWR.n2299 1.50638
R8022 VPWR.n6295 VPWR.n6229 1.49961
R8023 VPWR.n8009 VPWR.n5970 1.49961
R8024 VPWR.n5115 VPWR.n5114 1.49961
R8025 VPWR.n2378 VPWR.n2293 1.49961
R8026 VPWR.n6043 VPWR.n6042 1.49961
R8027 VPWR.n3071 VPWR.n3070 1.49961
R8028 VPWR.n3883 VPWR.n3036 1.49961
R8029 VPWR.n3906 VPWR.n3031 1.49961
R8030 VPWR.n3691 VPWR.n3513 1.49956
R8031 VPWR.n6176 VPWR.n6164 1.49932
R8032 VPWR.n224 VPWR.n223 1.49932
R8033 VPWR.n8150 VPWR.n8145 1.49932
R8034 VPWR.n8882 VPWR.n8881 1.49932
R8035 VPWR.n6519 VPWR.n6489 1.49932
R8036 VPWR.n8675 VPWR.n8672 1.49932
R8037 VPWR.n8640 VPWR.n8626 1.49932
R8038 VPWR.n8747 VPWR.n8743 1.49932
R8039 VPWR.n863 VPWR.n806 1.49932
R8040 VPWR.n619 VPWR.n600 1.49932
R8041 VPWR.n1115 VPWR.n731 1.49932
R8042 VPWR.n5793 VPWR.n5792 1.49932
R8043 VPWR.n1291 VPWR.n1287 1.49932
R8044 VPWR.n420 VPWR.n419 1.49932
R8045 VPWR.n5320 VPWR.n533 1.49932
R8046 VPWR.n4801 VPWR.n4797 1.49932
R8047 VPWR.n2185 VPWR.n2120 1.49932
R8048 VPWR.n4929 VPWR.n4925 1.49932
R8049 VPWR.n4410 VPWR.n2016 1.49932
R8050 VPWR.n4414 VPWR.n4412 1.49932
R8051 VPWR.n4483 VPWR.n1998 1.49932
R8052 VPWR.n4504 VPWR.n4503 1.49932
R8053 VPWR.n3386 VPWR.n3382 1.49932
R8054 VPWR.n2897 VPWR.n2893 1.49932
R8055 VPWR.n7654 VPWR.n7650 1.49932
R8056 VPWR.n87 VPWR.n68 1.49932
R8057 VPWR.n81 VPWR.n80 1.49932
R8058 VPWR.n4104 VPWR.n4100 1.49932
R8059 VPWR.n8306 VPWR.n8305 1.47352
R8060 VPWR.n8459 VPWR.n8458 1.47352
R8061 VPWR.n6542 VPWR.n6535 1.47352
R8062 VPWR.n837 VPWR.n818 1.47352
R8063 VPWR.n5141 VPWR.n1833 1.47352
R8064 VPWR.n1157 VPWR.n1156 1.46336
R8065 VPWR.n973 VPWR.n970 1.46336
R8066 VPWR.n5305 VPWR.n5304 1.46336
R8067 VPWR.n2068 VPWR.n2067 1.46336
R8068 VPWR.n3911 VPWR.n3910 1.45117
R8069 VPWR.n7764 VPWR.n7759 1.45117
R8070 VPWR.n6237 VPWR.n6236 1.45117
R8071 VPWR.n6752 VPWR.n6751 1.45117
R8072 VPWR.n6124 VPWR.n6122 1.4399
R8073 VPWR.n631 VPWR.n630 1.41226
R8074 VPWR.n1026 VPWR.n1024 1.38171
R8075 VPWR.n9019 VPWR.n9018 1.37571
R8076 VPWR.n8991 VPWR.n8990 1.37571
R8077 VPWR.n7944 VPWR.n7943 1.37571
R8078 VPWR.n5583 VPWR.n5582 1.37571
R8079 VPWR.n1484 VPWR.n1483 1.37571
R8080 VPWR.n2177 VPWR.n2176 1.37571
R8081 VPWR.n4379 VPWR.n4378 1.37571
R8082 VPWR.n4242 VPWR.n4241 1.37571
R8083 VPWR.n2844 VPWR.n2843 1.37571
R8084 VPWR.n3655 VPWR.n3654 1.37571
R8085 VPWR.n4782 VPWR.n4781 1.35979
R8086 VPWR.n8703 VPWR.n8702 1.35461
R8087 VPWR.n4870 VPWR.n4869 1.35461
R8088 VPWR.n4231 VPWR.n2865 1.35461
R8089 VPWR.n3329 VPWR.n3328 1.35461
R8090 VPWR.n9128 VPWR.n9127 1.35461
R8091 VPWR.n8965 VPWR.n8964 1.35461
R8092 VPWR.n4567 VPWR.n4566 1.35461
R8093 VPWR.n4170 VPWR.n4169 1.35461
R8094 VPWR.n7262 VPWR.n7261 1.35461
R8095 VPWR.n6869 VPWR.n6868 1.35459
R8096 VPWR.n6791 VPWR.n6790 1.35459
R8097 VPWR.n1642 VPWR.n561 1.35459
R8098 VPWR.n2546 VPWR.n2190 1.35459
R8099 VPWR.n2392 VPWR.n2391 1.35459
R8100 VPWR.n7737 VPWR.n7736 1.35459
R8101 VPWR.n7610 VPWR.n7609 1.35459
R8102 VPWR.n9132 VPWR.n9131 1.32113
R8103 VPWR.n4432 VPWR.n4431 1.32113
R8104 VPWR.n4014 VPWR.n4013 1.30773
R8105 VPWR.n8899 VPWR.n8898 1.30623
R8106 VPWR.n6722 VPWR.n6721 1.26992
R8107 VPWR.n6125 VPWR.n6119 1.26897
R8108 VPWR.n7763 VPWR.n7760 1.26897
R8109 VPWR.n6239 VPWR.n6238 1.26897
R8110 VPWR.n3066 VPWR.n3061 1.2502
R8111 VPWR.n9135 VPWR.n9134 1.2502
R8112 VPWR.n9203 VPWR.n9202 1.2502
R8113 VPWR.n6161 VPWR.n6160 1.2502
R8114 VPWR.n8115 VPWR.n338 1.2502
R8115 VPWR.n6668 VPWR.n6667 1.2502
R8116 VPWR.n8624 VPWR.n8623 1.2502
R8117 VPWR.n5871 VPWR.n5868 1.2502
R8118 VPWR.n6363 VPWR.n6362 1.2502
R8119 VPWR.n824 VPWR.n823 1.2502
R8120 VPWR.n815 VPWR.n814 1.2502
R8121 VPWR.n406 VPWR.n405 1.2502
R8122 VPWR.n467 VPWR.n466 1.2502
R8123 VPWR.n498 VPWR.n496 1.2502
R8124 VPWR.n1541 VPWR.n1540 1.2502
R8125 VPWR.n5005 VPWR.n5004 1.2502
R8126 VPWR.n1904 VPWR.n1903 1.2502
R8127 VPWR.n2297 VPWR.n2295 1.2502
R8128 VPWR.n1997 VPWR.n1996 1.2502
R8129 VPWR.n3938 VPWR.n3937 1.24652
R8130 VPWR.n446 VPWR.n445 1.2395
R8131 VPWR.n812 VPWR.n811 1.21955
R8132 VPWR.n3584 VPWR.n3583 1.21955
R8133 VPWR.n3631 VPWR.n3630 1.21955
R8134 VPWR.n4015 VPWR.n4014 1.1988
R8135 VPWR.n4013 VPWR.n4012 1.1988
R8136 VPWR.n8444 VPWR.n8443 1.16875
R8137 VPWR.n3888 VPWR.n3887 1.16414
R8138 VPWR.n4016 VPWR.n4015 1.14433
R8139 VPWR.n9122 VPWR.n148 1.13896
R8140 VPWR.n8959 VPWR.n299 1.13896
R8141 VPWR.n7894 VPWR.n7893 1.13896
R8142 VPWR.n8348 VPWR.n8347 1.13896
R8143 VPWR.n8416 VPWR.n8415 1.13896
R8144 VPWR.n923 VPWR.n922 1.13896
R8145 VPWR.n5379 VPWR.n5378 1.13896
R8146 VPWR.n5328 VPWR.n5327 1.13896
R8147 VPWR.n1825 VPWR.n1806 1.13896
R8148 VPWR.n4575 VPWR.n1975 1.13896
R8149 VPWR.n2629 VPWR.n2628 1.13896
R8150 VPWR.n4354 VPWR.n4353 1.13896
R8151 VPWR.n2503 VPWR.n2502 1.13896
R8152 VPWR.n1616 VPWR.n1615 1.13896
R8153 VPWR.n1328 VPWR.n1263 1.13896
R8154 VPWR.n648 VPWR.n577 1.13896
R8155 VPWR.n6545 VPWR.n6319 1.13896
R8156 VPWR.n6834 VPWR.n6833 1.13896
R8157 VPWR.n6201 VPWR.n6138 1.13896
R8158 VPWR.n2271 VPWR.n2196 1.13896
R8159 VPWR.n7731 VPWR.n7730 1.13896
R8160 VPWR.n4178 VPWR.n2983 1.13896
R8161 VPWR.n8960 VPWR.n8959 1.13896
R8162 VPWR.n4575 VPWR.n4574 1.13896
R8163 VPWR.n9123 VPWR.n9122 1.13896
R8164 VPWR.n9076 VPWR.n166 1.13885
R8165 VPWR.n8860 VPWR.n316 1.13885
R8166 VPWR.n8212 VPWR.n8211 1.13885
R8167 VPWR.n8729 VPWR.n345 1.13885
R8168 VPWR.n8582 VPWR.n8581 1.13885
R8169 VPWR.n5771 VPWR.n364 1.13885
R8170 VPWR.n1100 VPWR.n1099 1.13885
R8171 VPWR.n5706 VPWR.n5705 1.13885
R8172 VPWR.n5535 VPWR.n5534 1.13885
R8173 VPWR.n4632 VPWR.n4631 1.13885
R8174 VPWR.n5226 VPWR.n5225 1.13885
R8175 VPWR.n4989 VPWR.n4988 1.13885
R8176 VPWR.n5045 VPWR.n5044 1.13885
R8177 VPWR.n5988 VPWR.n5987 1.13885
R8178 VPWR.n3825 VPWR.n3824 1.13885
R8179 VPWR.n7002 VPWR.n7001 1.13885
R8180 VPWR.n3974 VPWR.n3973 1.13885
R8181 VPWR.n9278 VPWR.n9277 1.13885
R8182 VPWR.n6924 VPWR.n6923 1.13885
R8183 VPWR.n3359 VPWR.n3332 1.13885
R8184 VPWR.n4418 VPWR.n4417 1.13828
R8185 VPWR.n147 VPWR.n146 1.13717
R8186 VPWR.n298 VPWR.n297 1.13717
R8187 VPWR.n8079 VPWR.n8078 1.13717
R8188 VPWR.n6867 VPWR.n6866 1.13717
R8189 VPWR.n7891 VPWR.n7890 1.13717
R8190 VPWR.n8827 VPWR.n8826 1.13717
R8191 VPWR.n8090 VPWR.n8089 1.13717
R8192 VPWR.n6789 VPWR.n6788 1.13717
R8193 VPWR.n8358 VPWR.n8357 1.13717
R8194 VPWR.n8701 VPWR.n8700 1.13717
R8195 VPWR.n8579 VPWR.n8578 1.13717
R8196 VPWR.n6341 VPWR.n6340 1.13717
R8197 VPWR.n6432 VPWR.n6431 1.13717
R8198 VPWR.n5738 VPWR.n5737 1.13717
R8199 VPWR.n1097 VPWR.n1096 1.13717
R8200 VPWR.n1232 VPWR.n1231 1.13717
R8201 VPWR.n784 VPWR.n783 1.13717
R8202 VPWR.n5660 VPWR.n5659 1.13717
R8203 VPWR.n5520 VPWR.n5519 1.13717
R8204 VPWR.n1523 VPWR.n1522 1.13717
R8205 VPWR.n5367 VPWR.n5366 1.13717
R8206 VPWR.n4875 VPWR.n4874 1.13717
R8207 VPWR.n5211 VPWR.n5210 1.13717
R8208 VPWR.n1537 VPWR.n1536 1.13717
R8209 VPWR.n1761 VPWR.n1760 1.13717
R8210 VPWR.n4993 VPWR.n4992 1.13717
R8211 VPWR.n1869 VPWR.n1868 1.13717
R8212 VPWR.n2421 VPWR.n2420 1.13717
R8213 VPWR.n2595 VPWR.n2594 1.13717
R8214 VPWR.n2390 VPWR.n2389 1.13717
R8215 VPWR.n4351 VPWR.n4350 1.13717
R8216 VPWR.n2634 VPWR.n2633 1.13717
R8217 VPWR.n7858 VPWR.n7857 1.13717
R8218 VPWR.n2874 VPWR.n2873 1.13717
R8219 VPWR.n3754 VPWR.n3753 1.13717
R8220 VPWR.n3531 VPWR.n3530 1.13717
R8221 VPWR.n3107 VPWR.n3106 1.13717
R8222 VPWR.n7027 VPWR.n7026 1.13717
R8223 VPWR.n6968 VPWR.n6967 1.13717
R8224 VPWR.n6990 VPWR.n6989 1.13717
R8225 VPWR.n3827 VPWR.n3826 1.13717
R8226 VPWR.n3822 VPWR.n3819 1.13717
R8227 VPWR.n3773 VPWR.n3771 1.13717
R8228 VPWR.n3791 VPWR.n3790 1.13717
R8229 VPWR.n5995 VPWR.n5994 1.13717
R8230 VPWR.n7020 VPWR.n7019 1.13717
R8231 VPWR.n1827 VPWR.n1826 1.13717
R8232 VPWR.n5191 VPWR.n5190 1.13717
R8233 VPWR.n5197 VPWR.n5183 1.13717
R8234 VPWR.n5326 VPWR.n5325 1.13717
R8235 VPWR.n5348 VPWR.n5347 1.13717
R8236 VPWR.n5354 VPWR.n5340 1.13717
R8237 VPWR.n5377 VPWR.n5376 1.13717
R8238 VPWR.n5388 VPWR.n5387 1.13717
R8239 VPWR.n5381 VPWR.n511 1.13717
R8240 VPWR.n925 VPWR.n924 1.13717
R8241 VPWR.n914 VPWR.n913 1.13717
R8242 VPWR.n920 VPWR.n794 1.13717
R8243 VPWR.n8418 VPWR.n8417 1.13717
R8244 VPWR.n8407 VPWR.n8406 1.13717
R8245 VPWR.n8413 VPWR.n8399 1.13717
R8246 VPWR.n8346 VPWR.n8345 1.13717
R8247 VPWR.n5908 VPWR.n5907 1.13717
R8248 VPWR.n5914 VPWR.n5900 1.13717
R8249 VPWR.n7896 VPWR.n7895 1.13717
R8250 VPWR.n7970 VPWR.n7969 1.13717
R8251 VPWR.n7977 VPWR.n7976 1.13717
R8252 VPWR.n2608 VPWR.n2607 1.13717
R8253 VPWR.n2624 VPWR.n2623 1.13717
R8254 VPWR.n2627 VPWR.n2040 1.13717
R8255 VPWR.n5986 VPWR.n5984 1.13717
R8256 VPWR.n3119 VPWR.n3118 1.13717
R8257 VPWR.n3803 VPWR.n3802 1.13717
R8258 VPWR.n7000 VPWR.n6998 1.13717
R8259 VPWR.n3932 VPWR.n3931 1.13717
R8260 VPWR.n9285 VPWR.n9284 1.13717
R8261 VPWR.n3976 VPWR.n3975 1.13717
R8262 VPWR.n3971 VPWR.n3968 1.13717
R8263 VPWR.n4306 VPWR.n4305 1.13717
R8264 VPWR.n2757 VPWR.n2756 1.13717
R8265 VPWR.n2763 VPWR.n2749 1.13717
R8266 VPWR.n5061 VPWR.n5060 1.13717
R8267 VPWR.n5054 VPWR.n5053 1.13717
R8268 VPWR.n5043 VPWR.n5042 1.13717
R8269 VPWR.n5242 VPWR.n5241 1.13717
R8270 VPWR.n5235 VPWR.n5234 1.13717
R8271 VPWR.n5224 VPWR.n5223 1.13717
R8272 VPWR.n5551 VPWR.n5550 1.13717
R8273 VPWR.n5544 VPWR.n5543 1.13717
R8274 VPWR.n5533 VPWR.n5532 1.13717
R8275 VPWR.n1069 VPWR.n1068 1.13717
R8276 VPWR.n1062 VPWR.n1061 1.13717
R8277 VPWR.n1102 VPWR.n1101 1.13717
R8278 VPWR.n8550 VPWR.n8549 1.13717
R8279 VPWR.n8543 VPWR.n8542 1.13717
R8280 VPWR.n8584 VPWR.n8583 1.13717
R8281 VPWR.n8225 VPWR.n8224 1.13717
R8282 VPWR.n8232 VPWR.n8231 1.13717
R8283 VPWR.n8210 VPWR.n8209 1.13717
R8284 VPWR.n9097 VPWR.n9096 1.13717
R8285 VPWR.n176 VPWR.n175 1.13717
R8286 VPWR.n9078 VPWR.n9077 1.13717
R8287 VPWR.n4357 VPWR.n4356 1.13717
R8288 VPWR.n4316 VPWR.n4315 1.13717
R8289 VPWR.n2780 VPWR.n2779 1.13717
R8290 VPWR.n4334 VPWR.n4333 1.13717
R8291 VPWR.n3016 VPWR.n3015 1.13717
R8292 VPWR.n9215 VPWR.n24 1.13717
R8293 VPWR.n9237 VPWR.n9236 1.13717
R8294 VPWR.n9245 VPWR.n9244 1.13717
R8295 VPWR.n9276 VPWR.n9272 1.13717
R8296 VPWR.n7735 VPWR.n7734 1.13717
R8297 VPWR.n7612 VPWR.n7611 1.13717
R8298 VPWR.n3477 VPWR.n3476 1.13717
R8299 VPWR.n3438 VPWR.n3437 1.13717
R8300 VPWR.n7702 VPWR.n7701 1.13717
R8301 VPWR.n7634 VPWR.n7628 1.13717
R8302 VPWR.n2511 VPWR.n2510 1.13717
R8303 VPWR.n2518 VPWR.n2517 1.13717
R8304 VPWR.n2501 VPWR.n2499 1.13717
R8305 VPWR.n1625 VPWR.n1624 1.13717
R8306 VPWR.n1618 VPWR.n576 1.13717
R8307 VPWR.n1614 VPWR.n1612 1.13717
R8308 VPWR.n1255 VPWR.n1254 1.13717
R8309 VPWR.n1261 VPWR.n1248 1.13717
R8310 VPWR.n1331 VPWR.n1330 1.13717
R8311 VPWR.n678 VPWR.n591 1.13717
R8312 VPWR.n685 VPWR.n684 1.13717
R8313 VPWR.n651 VPWR.n650 1.13717
R8314 VPWR.n6575 VPWR.n6574 1.13717
R8315 VPWR.n6581 VPWR.n6568 1.13717
R8316 VPWR.n6548 VPWR.n6547 1.13717
R8317 VPWR.n6854 VPWR.n6853 1.13717
R8318 VPWR.n6860 VPWR.n6847 1.13717
R8319 VPWR.n6832 VPWR.n6830 1.13717
R8320 VPWR.n6886 VPWR.n6885 1.13717
R8321 VPWR.n6892 VPWR.n6151 1.13717
R8322 VPWR.n6204 VPWR.n6203 1.13717
R8323 VPWR.n2402 VPWR.n2401 1.13717
R8324 VPWR.n2408 VPWR.n2209 1.13717
R8325 VPWR.n2274 VPWR.n2273 1.13717
R8326 VPWR.n7729 VPWR.n7727 1.13717
R8327 VPWR.n3444 VPWR.n3443 1.13717
R8328 VPWR.n6930 VPWR.n6929 1.13717
R8329 VPWR.n6916 VPWR.n6915 1.13717
R8330 VPWR.n6922 VPWR.n6920 1.13717
R8331 VPWR.n3135 VPWR.n3132 1.13717
R8332 VPWR.n3339 VPWR.n3338 1.13717
R8333 VPWR.n3331 VPWR.n3330 1.13717
R8334 VPWR.n3356 VPWR.n3355 1.13717
R8335 VPWR.n4176 VPWR.n4175 1.13717
R8336 VPWR.n4217 VPWR.n4216 1.13717
R8337 VPWR.n2955 VPWR.n2883 1.13717
R8338 VPWR.n2969 VPWR.n2968 1.13717
R8339 VPWR.n4573 VPWR.n4571 1.13717
R8340 VPWR.n4904 VPWR.n4903 1.13717
R8341 VPWR.n4888 VPWR.n4887 1.13717
R8342 VPWR.n4987 VPWR.n4986 1.13717
R8343 VPWR.n4620 VPWR.n4619 1.13717
R8344 VPWR.n4604 VPWR.n4603 1.13717
R8345 VPWR.n4630 VPWR.n4629 1.13717
R8346 VPWR.n5731 VPWR.n5730 1.13717
R8347 VPWR.n5715 VPWR.n5714 1.13717
R8348 VPWR.n5704 VPWR.n5703 1.13717
R8349 VPWR.n5850 VPWR.n5849 1.13717
R8350 VPWR.n373 VPWR.n372 1.13717
R8351 VPWR.n5773 VPWR.n5772 1.13717
R8352 VPWR.n8820 VPWR.n8819 1.13717
R8353 VPWR.n8804 VPWR.n8803 1.13717
R8354 VPWR.n8731 VPWR.n8730 1.13717
R8355 VPWR.n8940 VPWR.n8939 1.13717
R8356 VPWR.n325 VPWR.n324 1.13717
R8357 VPWR.n8862 VPWR.n8861 1.13717
R8358 VPWR.n8957 VPWR.n8954 1.13717
R8359 VPWR.n314 VPWR.n310 1.13717
R8360 VPWR.n8963 VPWR.n8962 1.13717
R8361 VPWR.n1990 VPWR.n1989 1.13717
R8362 VPWR.n1974 VPWR.n1973 1.13717
R8363 VPWR.n4590 VPWR.n4589 1.13717
R8364 VPWR.n9120 VPWR.n9117 1.13717
R8365 VPWR.n161 VPWR.n160 1.13717
R8366 VPWR.n9126 VPWR.n9125 1.13717
R8367 VPWR.n2982 VPWR.n2981 1.13717
R8368 VPWR.n4204 VPWR.n4201 1.13717
R8369 VPWR.n4185 VPWR.n4184 1.13717
R8370 VPWR.n7241 VPWR.n7240 1.13717
R8371 VPWR.n7229 VPWR.n7228 1.13717
R8372 VPWR.n7255 VPWR.n7254 1.13717
R8373 VPWR.n7260 VPWR.n7259 1.13717
R8374 VPWR.n3823 VPWR.n3822 1.1368
R8375 VPWR.n5198 VPWR.n5197 1.1368
R8376 VPWR.n5355 VPWR.n5354 1.1368
R8377 VPWR.n5381 VPWR.n5380 1.1368
R8378 VPWR.n921 VPWR.n920 1.1368
R8379 VPWR.n8414 VPWR.n8413 1.1368
R8380 VPWR.n5915 VPWR.n5914 1.1368
R8381 VPWR.n7976 VPWR.n7863 1.1368
R8382 VPWR.n2625 VPWR.n2624 1.1368
R8383 VPWR.n7021 VPWR.n7020 1.1368
R8384 VPWR.n6991 VPWR.n6990 1.1368
R8385 VPWR.n3972 VPWR.n3971 1.1368
R8386 VPWR.n2764 VPWR.n2763 1.1368
R8387 VPWR.n7635 VPWR.n7634 1.1368
R8388 VPWR.n2517 VPWR.n2504 1.1368
R8389 VPWR.n1618 VPWR.n1617 1.1368
R8390 VPWR.n1262 VPWR.n1261 1.1368
R8391 VPWR.n684 VPWR.n677 1.1368
R8392 VPWR.n6582 VPWR.n6581 1.1368
R8393 VPWR.n6861 VPWR.n6860 1.1368
R8394 VPWR.n6893 VPWR.n6892 1.1368
R8395 VPWR.n2409 VPWR.n2408 1.1368
R8396 VPWR.n6917 VPWR.n6916 1.1368
R8397 VPWR.n8958 VPWR.n8957 1.1368
R8398 VPWR.n315 VPWR.n314 1.1368
R8399 VPWR.n162 VPWR.n161 1.1368
R8400 VPWR.n9121 VPWR.n9120 1.1368
R8401 VPWR.n4205 VPWR.n4204 1.1368
R8402 VPWR.n7229 VPWR.n7141 1.1368
R8403 VPWR.n2596 VPWR.n2595 1.13669
R8404 VPWR.n1760 VPWR.n514 1.13669
R8405 VPWR.n5368 VPWR.n5367 1.13669
R8406 VPWR.n785 VPWR.n784 1.13669
R8407 VPWR.n6431 VPWR.n5888 1.13669
R8408 VPWR.n8359 VPWR.n8358 1.13669
R8409 VPWR.n7892 VPWR.n7891 1.13669
R8410 VPWR.n2633 VPWR.n2631 1.13669
R8411 VPWR.n7859 VPWR.n7858 1.13669
R8412 VPWR.n3108 VPWR.n3107 1.13669
R8413 VPWR.n7026 VPWR.n7024 1.13669
R8414 VPWR.n4352 VPWR.n4351 1.13669
R8415 VPWR.n1870 VPWR.n1869 1.13669
R8416 VPWR.n5060 VPWR.n5046 1.13669
R8417 VPWR.n5212 VPWR.n5211 1.13669
R8418 VPWR.n5241 VPWR.n5227 1.13669
R8419 VPWR.n5521 VPWR.n5520 1.13669
R8420 VPWR.n5550 VPWR.n5536 1.13669
R8421 VPWR.n1098 VPWR.n1097 1.13669
R8422 VPWR.n1068 VPWR.n746 1.13669
R8423 VPWR.n8580 VPWR.n8579 1.13669
R8424 VPWR.n8549 VPWR.n361 1.13669
R8425 VPWR.n8091 VPWR.n8090 1.13669
R8426 VPWR.n8225 VPWR.n8213 1.13669
R8427 VPWR.n8080 VPWR.n8079 1.13669
R8428 VPWR.n9098 VPWR.n9097 1.13669
R8429 VPWR.n3931 VPWR.n3005 1.13669
R8430 VPWR.n9284 VPWR.n9282 1.13669
R8431 VPWR.n9279 VPWR.n24 1.13669
R8432 VPWR.n9244 VPWR.n25 1.13669
R8433 VPWR.n7734 VPWR.n7732 1.13669
R8434 VPWR.n2422 VPWR.n2421 1.13669
R8435 VPWR.n1538 VPWR.n1537 1.13669
R8436 VPWR.n1524 VPWR.n1523 1.13669
R8437 VPWR.n1233 VPWR.n1232 1.13669
R8438 VPWR.n6340 VPWR.n6338 1.13669
R8439 VPWR.n6788 VPWR.n6585 1.13669
R8440 VPWR.n6866 VPWR.n6864 1.13669
R8441 VPWR.n2389 VPWR.n2387 1.13669
R8442 VPWR.n7613 VPWR.n7612 1.13669
R8443 VPWR.n3360 VPWR.n3135 1.13669
R8444 VPWR.n3358 VPWR.n3356 1.13669
R8445 VPWR.n4992 VPWR.n4990 1.13669
R8446 VPWR.n4905 VPWR.n4904 1.13669
R8447 VPWR.n4876 VPWR.n4875 1.13669
R8448 VPWR.n4621 VPWR.n4620 1.13669
R8449 VPWR.n5659 VPWR.n394 1.13669
R8450 VPWR.n5732 VPWR.n5731 1.13669
R8451 VPWR.n5737 VPWR.n5735 1.13669
R8452 VPWR.n5851 VPWR.n5850 1.13669
R8453 VPWR.n8700 VPWR.n8698 1.13669
R8454 VPWR.n8821 VPWR.n8820 1.13669
R8455 VPWR.n8826 VPWR.n8824 1.13669
R8456 VPWR.n8941 VPWR.n8940 1.13669
R8457 VPWR.n1991 VPWR.n1990 1.13669
R8458 VPWR.n4591 VPWR.n4590 1.13669
R8459 VPWR.n4177 VPWR.n4176 1.13669
R8460 VPWR.n103 VPWR.n102 1.12991
R8461 VPWR.n8913 VPWR.n8912 1.12991
R8462 VPWR.n6346 VPWR.n6345 1.12991
R8463 VPWR.n5813 VPWR.n5812 1.12991
R8464 VPWR.n1041 VPWR.n1040 1.12991
R8465 VPWR.n617 VPWR.n616 1.12991
R8466 VPWR.n4681 VPWR.n4680 1.12991
R8467 VPWR.n2663 VPWR.n2662 1.12991
R8468 VPWR.n6259 VPWR.n6257 1.10819
R8469 VPWR.n5314 VPWR.n5313 1.09764
R8470 VPWR.n6261 VPWR.n6240 1.09272
R8471 VPWR.n6189 VPWR.n6188 1.09272
R8472 VPWR.n6366 VPWR.n6364 1.09272
R8473 VPWR.n8427 VPWR.n5872 1.09272
R8474 VPWR.n1580 VPWR.n1543 1.09272
R8475 VPWR.n7768 VPWR.n6126 1.09272
R8476 VPWR.n7676 VPWR.n7675 1.09272
R8477 VPWR.n3069 VPWR.n3068 1.09272
R8478 VPWR.n8182 VPWR.n8116 1.09216
R8479 VPWR.n827 VPWR.n825 1.09216
R8480 VPWR.n5437 VPWR.n499 1.09216
R8481 VPWR.n5595 VPWR.n469 1.09216
R8482 VPWR.n438 VPWR.n435 1.09216
R8483 VPWR.n9204 VPWR.n31 1.09216
R8484 VPWR.n850 VPWR.n816 1.09203
R8485 VPWR.n1127 VPWR.n1126 1.08641
R8486 VPWR.n2472 VPWR.n2423 1.08641
R8487 VPWR.n9034 VPWR.n9033 1.05835
R8488 VPWR.n5468 VPWR.n5466 1.05773
R8489 VPWR.n4533 VPWR.n4485 1.05773
R8490 VPWR.n4094 VPWR.n4091 0.992049
R8491 VPWR.n4116 VPWR.n4112 0.992049
R8492 VPWR.n47 VPWR.n46 0.965579
R8493 VPWR.n236 VPWR.n235 0.965579
R8494 VPWR.n264 VPWR.n263 0.965579
R8495 VPWR.n5926 VPWR.n5925 0.965579
R8496 VPWR.n5599 VPWR.n5598 0.965579
R8497 VPWR.n5457 VPWR.n492 0.965579
R8498 VPWR.n9180 VPWR.n9179 0.948229
R8499 VPWR.n7040 VPWR.n7039 0.935332
R8500 VPWR.n8503 VPWR.n8502 0.935332
R8501 VPWR.n7274 VPWR.n7273 0.935332
R8502 VPWR.n9134 VPWR.n9132 0.914786
R8503 VPWR.n5137 VPWR.n5136 0.914786
R8504 VPWR.n4433 VPWR.n4432 0.914786
R8505 VPWR.n761 VPWR.n760 0.911172
R8506 VPWR.n3215 VPWR.n3214 0.899674
R8507 VPWR.n7654 VPWR.n7648 0.899674
R8508 VPWR.n6176 VPWR.n6163 0.899674
R8509 VPWR.n2120 VPWR.n2116 0.899674
R8510 VPWR.n3386 VPWR.n3380 0.899674
R8511 VPWR.n7529 VPWR.n7528 0.863992
R8512 VPWR.n7562 VPWR.n7561 0.863992
R8513 VPWR.n7299 VPWR.n7298 0.863992
R8514 VPWR.n3277 VPWR.n3276 0.863992
R8515 VPWR.n7122 VPWR.n7121 0.863992
R8516 VPWR.n7159 VPWR.n7158 0.863992
R8517 VPWR.n4111 VPWR.n4110 0.842756
R8518 VPWR.n3038 VPWR.n3037 0.828042
R8519 VPWR.n427 VPWR.n426 0.813843
R8520 VPWR.n4017 VPWR.n4009 0.790287
R8521 VPWR.n8150 VPWR.n8125 0.769318
R8522 VPWR.n8675 VPWR.n8674 0.769318
R8523 VPWR.n806 VPWR.n805 0.769318
R8524 VPWR.n293 VPWR.n292 0.762405
R8525 VPWR.n1994 VPWR.n1993 0.762405
R8526 VPWR.n3168 VPWR.n3159 0.753441
R8527 VPWR.n4120 VPWR.n4119 0.753441
R8528 VPWR.n9187 VPWR.n36 0.753441
R8529 VPWR.n6083 VPWR.n6064 0.753441
R8530 VPWR.n8242 VPWR.n8241 0.753441
R8531 VPWR.n844 VPWR.n841 0.753441
R8532 VPWR.n844 VPWR.n843 0.753441
R8533 VPWR.n1090 VPWR.n1089 0.753441
R8534 VPWR.n1019 VPWR.n1018 0.753441
R8535 VPWR.n1001 VPWR.n1000 0.753441
R8536 VPWR.n629 VPWR.n627 0.753441
R8537 VPWR.n5409 VPWR.n5408 0.753441
R8538 VPWR.n4750 VPWR.n4694 0.753441
R8539 VPWR.n4758 VPWR.n4689 0.753441
R8540 VPWR.n5107 VPWR.n5106 0.753441
R8541 VPWR.n2264 VPWR.n2263 0.753441
R8542 VPWR.n2240 VPWR.n2239 0.753441
R8543 VPWR.n2235 VPWR.n2234 0.753441
R8544 VPWR.n2368 VPWR.n2367 0.753441
R8545 VPWR.n6648 VPWR.n6647 0.740996
R8546 VPWR.n2305 VPWR.n2304 0.740996
R8547 VPWR.n976 VPWR.n975 0.731929
R8548 VPWR.n4702 VPWR.n4701 0.731929
R8549 VPWR.n4733 VPWR.n4732 0.731929
R8550 VPWR.n6800 VPWR.n6799 0.698804
R8551 VPWR.n8338 VPWR.n8337 0.660817
R8552 VPWR VPWR.n6559 0.660817
R8553 VPWR.n4964 VPWR.n4963 0.660817
R8554 VPWR.n7692 VPWR.n7691 0.656731
R8555 VPWR.n6878 VPWR.n6877 0.656731
R8556 VPWR.n3063 VPWR.n3062 0.651997
R8557 VPWR.n7678 VPWR.n7636 0.651997
R8558 VPWR.n6191 VPWR.n6156 0.651997
R8559 VPWR.n3071 VPWR.n3059 0.644287
R8560 VPWR.n6671 VPWR.n6670 0.644287
R8561 VPWR.n5872 VPWR.n5870 0.644287
R8562 VPWR.n825 VPWR.n821 0.644287
R8563 VPWR.n438 VPWR.n437 0.644287
R8564 VPWR.n499 VPWR.n497 0.644287
R8565 VPWR.n5006 VPWR.n1964 0.644287
R8566 VPWR.n1951 VPWR.n1901 0.644287
R8567 VPWR.n7498 VPWR.n6952 0.635211
R8568 VPWR.n7474 VPWR.n7473 0.635211
R8569 VPWR.n7571 VPWR.n7570 0.635211
R8570 VPWR.n7514 VPWR.n6941 0.635211
R8571 VPWR.n7455 VPWR.n6956 0.635211
R8572 VPWR.n7402 VPWR.n7030 0.635211
R8573 VPWR.n3871 VPWR.n3870 0.635211
R8574 VPWR.n3175 VPWR.n3153 0.635211
R8575 VPWR.n3209 VPWR.n3208 0.635211
R8576 VPWR.n3999 VPWR.n3998 0.635211
R8577 VPWR.n4002 VPWR.n4001 0.635211
R8578 VPWR.n3901 VPWR.n3900 0.635211
R8579 VPWR.n4127 VPWR.n4126 0.635211
R8580 VPWR.n3288 VPWR.n3287 0.635211
R8581 VPWR.n3216 VPWR.n3144 0.635211
R8582 VPWR.n7656 VPWR.n7655 0.635211
R8583 VPWR.n7660 VPWR.n7659 0.635211
R8584 VPWR.n6050 VPWR.n6013 0.635211
R8585 VPWR.n8017 VPWR.n8016 0.635211
R8586 VPWR.n8044 VPWR.n5964 0.635211
R8587 VPWR.n9020 VPWR.n9019 0.635211
R8588 VPWR.n9046 VPWR.n8975 0.635211
R8589 VPWR.n8987 VPWR.n8986 0.635211
R8590 VPWR.n9016 VPWR.n9015 0.635211
R8591 VPWR.n8984 VPWR.n8979 0.635211
R8592 VPWR.n7952 VPWR.n7902 0.635211
R8593 VPWR.n7922 VPWR.n7903 0.635211
R8594 VPWR.n8282 VPWR.n5946 0.635211
R8595 VPWR.n8257 VPWR.n5949 0.635211
R8596 VPWR.n6725 VPWR.n6649 0.635211
R8597 VPWR.n6726 VPWR.n6648 0.635211
R8598 VPWR.n6617 VPWR.n6616 0.635211
R8599 VPWR.n8462 VPWR.n8461 0.635211
R8600 VPWR.n8485 VPWR.n5862 0.635211
R8601 VPWR.n6407 VPWR.n6356 0.635211
R8602 VPWR.n6408 VPWR.n6353 0.635211
R8603 VPWR.n446 VPWR.n401 0.635211
R8604 VPWR.n5615 VPWR.n5614 0.635211
R8605 VPWR.n457 VPWR.n456 0.635211
R8606 VPWR.n5513 VPWR.n5511 0.635211
R8607 VPWR.n473 VPWR.n472 0.635211
R8608 VPWR.n1487 VPWR.n1377 0.635211
R8609 VPWR.n1458 VPWR.n1378 0.635211
R8610 VPWR.n1489 VPWR.n1376 0.635211
R8611 VPWR.n1515 VPWR.n1514 0.635211
R8612 VPWR.n1371 VPWR.n1370 0.635211
R8613 VPWR.n4827 VPWR.n4787 0.635211
R8614 VPWR.n4814 VPWR.n4813 0.635211
R8615 VPWR.n4802 VPWR.n4793 0.635211
R8616 VPWR.n4828 VPWR.n4786 0.635211
R8617 VPWR.n1704 VPWR.n1703 0.635211
R8618 VPWR.n1711 VPWR.n1710 0.635211
R8619 VPWR.n1671 VPWR.n1670 0.635211
R8620 VPWR.n1668 VPWR.n558 0.635211
R8621 VPWR.n2183 VPWR.n2182 0.635211
R8622 VPWR.n2153 VPWR.n2121 0.635211
R8623 VPWR.n2701 VPWR.n2700 0.635211
R8624 VPWR.n2727 VPWR.n2726 0.635211
R8625 VPWR.n4408 VPWR.n4406 0.635211
R8626 VPWR.n2364 VPWR.n2305 0.635211
R8627 VPWR.n2337 VPWR.n2306 0.635211
R8628 VPWR.n4492 VPWR.n4491 0.635211
R8629 VPWR.n4243 VPWR.n4242 0.635211
R8630 VPWR.n2835 VPWR.n2834 0.635211
R8631 VPWR.n2794 VPWR.n2793 0.635211
R8632 VPWR.n3596 VPWR.n3595 0.635211
R8633 VPWR.n3523 VPWR.n3522 0.635211
R8634 VPWR.n3719 VPWR.n3506 0.635211
R8635 VPWR.n3692 VPWR.n3509 0.635211
R8636 VPWR.n2801 VPWR.n2800 0.635211
R8637 VPWR.n3662 VPWR.n3632 0.635211
R8638 VPWR.n4251 VPWR.n2788 0.635211
R8639 VPWR.n7082 VPWR.n7081 0.635211
R8640 VPWR.n7106 VPWR.n7049 0.635211
R8641 VPWR.n6257 VPWR.n6256 0.615885
R8642 VPWR.n7991 VPWR.n7989 0.61457
R8643 VPWR.n951 VPWR.n950 0.607615
R8644 VPWR.n6895 VPWR.n164 0.546928
R8645 VPWR.n675 VPWR.n363 0.546928
R8646 VPWR.n5201 VPWR.n1805 0.546928
R8647 VPWR.n7038 VPWR.n7035 0.539826
R8648 VPWR.n8508 VPWR.n8507 0.539826
R8649 VPWR.n7271 VPWR.n7270 0.539826
R8650 VPWR.n4840 VPWR.n4839 0.529114
R8651 VPWR.n3209 VPWR.n3146 0.509294
R8652 VPWR.n7297 VPWR.n7296 0.508436
R8653 VPWR.n7329 VPWR.n7328 0.508436
R8654 VPWR.n7995 VPWR.n7994 0.508436
R8655 VPWR.n8570 VPWR.n8569 0.508436
R8656 VPWR.n888 VPWR.n887 0.508436
R8657 VPWR.n5134 VPWR.n5133 0.508436
R8658 VPWR.n9138 VPWR.n9137 0.491807
R8659 VPWR.n7684 VPWR.n7683 0.491355
R8660 VPWR.n6197 VPWR.n6196 0.491355
R8661 VPWR.n6256 VPWR.n6255 0.488391
R8662 VPWR.n3691 VPWR.n3514 0.440094
R8663 VPWR.n1513 VPWR.n1371 0.428356
R8664 VPWR.n8921 VPWR.n8920 0.426482
R8665 VPWR.n7670 VPWR.n7638 0.42364
R8666 VPWR.n6287 VPWR.n6230 0.42364
R8667 VPWR.n6381 VPWR.n6380 0.42364
R8668 VPWR.n5685 VPWR.n5684 0.42364
R8669 VPWR.n5563 VPWR.n5562 0.42364
R8670 VPWR.n4793 VPWR.n4792 0.42364
R8671 VPWR.n1788 VPWR.n1787 0.42364
R8672 VPWR.n1795 VPWR.n1794 0.42364
R8673 VPWR.n2787 VPWR.n2785 0.42364
R8674 VPWR.n6364 VPWR.n6360 0.411567
R8675 VPWR.n3774 VPWR.n3120 0.3805
R8676 VPWR.n3937 VPWR.n3936 0.378081
R8677 VPWR.n248 VPWR.n247 0.376971
R8678 VPWR.n8604 VPWR.n8603 0.376971
R8679 VPWR.n4944 VPWR.n4943 0.376971
R8680 VPWR.n2542 VPWR.n2541 0.376971
R8681 VPWR.n3200 VPWR.n3151 0.369731
R8682 VPWR.n3185 VPWR.n3152 0.369731
R8683 VPWR.n4033 VPWR.n4032 0.369731
R8684 VPWR.n4052 VPWR.n2996 0.369731
R8685 VPWR.n4076 VPWR.n4075 0.369731
R8686 VPWR.n4128 VPWR.n4086 0.369731
R8687 VPWR.n7752 VPWR.n7751 0.369731
R8688 VPWR.n6122 VPWR.n6121 0.369731
R8689 VPWR.n7782 VPWR.n6118 0.369731
R8690 VPWR.n7784 VPWR.n7783 0.369731
R8691 VPWR.n7790 VPWR.n6116 0.369731
R8692 VPWR.n7793 VPWR.n7792 0.369731
R8693 VPWR.n6114 VPWR.n6113 0.369731
R8694 VPWR.n7811 VPWR.n7810 0.369731
R8695 VPWR.n7815 VPWR.n6009 0.369731
R8696 VPWR.n6027 VPWR.n6019 0.369731
R8697 VPWR.n6030 VPWR.n6029 0.369731
R8698 VPWR.n6034 VPWR.n6018 0.369731
R8699 VPWR.n6259 VPWR.n6258 0.369731
R8700 VPWR.n5968 VPWR.n5967 0.369731
R8701 VPWR.n6298 VPWR.n6226 0.369731
R8702 VPWR.n6636 VPWR.n6635 0.369731
R8703 VPWR.n6766 VPWR.n6641 0.369731
R8704 VPWR.n1687 VPWR.n1686 0.369731
R8705 VPWR.n1702 VPWR.n557 0.369731
R8706 VPWR.n2921 VPWR.n2888 0.369731
R8707 VPWR.n2898 VPWR.n2889 0.369731
R8708 VPWR.n1186 VPWR.n1185 0.366214
R8709 VPWR.n966 VPWR.n965 0.366214
R8710 VPWR.n5309 VPWR.n5308 0.366214
R8711 VPWR.n5318 VPWR.n536 0.366214
R8712 VPWR.n4436 VPWR.n4429 0.358558
R8713 VPWR.n9101 VPWR.n164 0.356928
R8714 VPWR.n9102 VPWR.n9101 0.356928
R8715 VPWR.n5855 VPWR.n363 0.356928
R8716 VPWR.n5855 VPWR.n5854 0.356928
R8717 VPWR.n5203 VPWR.n5201 0.356928
R8718 VPWR.n5203 VPWR.n5202 0.356928
R8719 VPWR.n1124 VPWR.n1123 0.356056
R8720 VPWR.n2554 VPWR.n2188 0.356056
R8721 VPWR.n2479 VPWR.n2478 0.356056
R8722 VPWR.n4466 VPWR.n4465 0.356056
R8723 VPWR.n3726 VPWR.n3725 0.356056
R8724 VPWR.n3759 VPWR.n3758 0.352216
R8725 VPWR.n1209 VPWR.n1208 0.349591
R8726 VPWR.n3124 VPWR.n2782 0.347759
R8727 VPWR.n2975 VPWR.n2974 0.34507
R8728 VPWR.n3792 VPWR.n3791 0.342503
R8729 VPWR.n3774 VPWR.n3773 0.3424
R8730 VPWR.n4210 VPWR.n2883 0.3424
R8731 VPWR.n3774 VPWR.n3123 0.341811
R8732 VPWR.n4319 VPWR.n4308 0.341811
R8733 VPWR.n4319 VPWR.n4318 0.341811
R8734 VPWR.n3756 VPWR.n3755 0.341811
R8735 VPWR.n4210 VPWR.n2972 0.341811
R8736 VPWR.n7953 VPWR.n7952 0.322528
R8737 VPWR.n2835 VPWR.n2833 0.322528
R8738 VPWR.n8066 VPWR.n8065 0.317855
R8739 VPWR.n6652 VPWR.n6651 0.317855
R8740 VPWR.n6696 VPWR.n6652 0.317855
R8741 VPWR.n4832 VPWR.n4831 0.317855
R8742 VPWR.n3438 VPWR.n3128 0.31175
R8743 VPWR.n2781 VPWR.n2780 0.311379
R8744 VPWR.n4335 VPWR.n4334 0.311379
R8745 VPWR.n4216 VPWR.n4211 0.311379
R8746 VPWR.n3476 VPWR.n3364 0.311321
R8747 VPWR.n6812 VPWR.n6810 0.308192
R8748 VPWR.n6950 VPWR.n6949 0.305262
R8749 VPWR.n7499 VPWR.n6951 0.305262
R8750 VPWR.n7534 VPWR.n7528 0.305262
R8751 VPWR.n7563 VPWR.n7562 0.305262
R8752 VPWR.n7569 VPWR.n7527 0.305262
R8753 VPWR.n7381 VPWR.n7380 0.305262
R8754 VPWR.n7045 VPWR.n7044 0.305262
R8755 VPWR.n7373 VPWR.n7283 0.305262
R8756 VPWR.n7289 VPWR.n7288 0.305262
R8757 VPWR.n7356 VPWR.n7293 0.305262
R8758 VPWR.n7350 VPWR.n7299 0.305262
R8759 VPWR.n7331 VPWR.n7330 0.305262
R8760 VPWR.n3054 VPWR.n3053 0.305262
R8761 VPWR.n4106 VPWR.n4105 0.305262
R8762 VPWR.n3278 VPWR.n3277 0.305262
R8763 VPWR.n3285 VPWR.n3233 0.305262
R8764 VPWR.n3252 VPWR.n3251 0.305262
R8765 VPWR.n3257 VPWR.n3241 0.305262
R8766 VPWR.n107 VPWR.n62 0.305262
R8767 VPWR.n9144 VPWR.n59 0.305262
R8768 VPWR.n9151 VPWR.n52 0.305262
R8769 VPWR.n9145 VPWR.n57 0.305262
R8770 VPWR.n9167 VPWR.n43 0.305262
R8771 VPWR.n9162 VPWR.n48 0.305262
R8772 VPWR.n9185 VPWR.n41 0.305262
R8773 VPWR.n9180 VPWR.n42 0.305262
R8774 VPWR.n6104 VPWR.n6103 0.305262
R8775 VPWR.n6089 VPWR.n6063 0.305262
R8776 VPWR.n6067 VPWR.n6065 0.305262
R8777 VPWR.n6075 VPWR.n6074 0.305262
R8778 VPWR.n211 VPWR.n210 0.305262
R8779 VPWR.n231 VPWR.n212 0.305262
R8780 VPWR.n7954 VPWR.n7901 0.305262
R8781 VPWR.n8904 VPWR.n8867 0.305262
R8782 VPWR.n8899 VPWR.n8868 0.305262
R8783 VPWR.n8152 VPWR.n8151 0.305262
R8784 VPWR.n8123 VPWR.n8122 0.305262
R8785 VPWR.n8332 VPWR.n5924 0.305262
R8786 VPWR.n5929 VPWR.n5928 0.305262
R8787 VPWR.n5938 VPWR.n5937 0.305262
R8788 VPWR.n8283 VPWR.n5943 0.305262
R8789 VPWR.n8197 VPWR.n8196 0.305262
R8790 VPWR.n8188 VPWR.n8110 0.305262
R8791 VPWR.n8758 VPWR.n8757 0.305262
R8792 VPWR.n8748 VPWR.n8739 0.305262
R8793 VPWR.n8787 VPWR.n8786 0.305262
R8794 VPWR.n8773 VPWR.n8732 0.305262
R8795 VPWR.n8633 VPWR.n8629 0.305262
R8796 VPWR.n8615 VPWR.n8614 0.305262
R8797 VPWR.n8656 VPWR.n8619 0.305262
R8798 VPWR.n8445 VPWR.n8444 0.305262
R8799 VPWR.n8459 VPWR.n8457 0.305262
R8800 VPWR.n8538 VPWR.n8537 0.305262
R8801 VPWR.n6375 VPWR.n6357 0.305262
R8802 VPWR.n6502 VPWR.n6501 0.305262
R8803 VPWR.n6512 VPWR.n6511 0.305262
R8804 VPWR.n1197 VPWR.n1196 0.305262
R8805 VPWR.n5744 VPWR.n386 0.305262
R8806 VPWR.n1127 VPWR.n725 0.305262
R8807 VPWR.n1132 VPWR.n1131 0.305262
R8808 VPWR.n1121 VPWR.n1120 0.305262
R8809 VPWR.n1026 VPWR.n1025 0.305262
R8810 VPWR.n754 VPWR.n753 0.305262
R8811 VPWR.n868 VPWR.n867 0.305262
R8812 VPWR.n932 VPWR.n765 0.305262
R8813 VPWR.n856 VPWR.n812 0.305262
R8814 VPWR.n642 VPWR.n641 0.305262
R8815 VPWR.n427 VPWR.n407 0.305262
R8816 VPWR.n5604 VPWR.n464 0.305262
R8817 VPWR.n5458 VPWR.n5457 0.305262
R8818 VPWR.n5462 VPWR.n5461 0.305262
R8819 VPWR.n5446 VPWR.n494 0.305262
R8820 VPWR.n1293 VPWR.n1292 0.305262
R8821 VPWR.n1303 VPWR.n1274 0.305262
R8822 VPWR.n554 VPWR.n553 0.305262
R8823 VPWR.n1775 VPWR.n548 0.305262
R8824 VPWR.n4920 VPWR.n4919 0.305262
R8825 VPWR.n4930 VPWR.n4921 0.305262
R8826 VPWR.n4956 VPWR.n4912 0.305262
R8827 VPWR.n1898 VPWR.n1897 0.305262
R8828 VPWR.n5015 VPWR.n5014 0.305262
R8829 VPWR.n5007 VPWR.n1963 0.305262
R8830 VPWR.n5131 VPWR.n1833 0.305262
R8831 VPWR.n5125 VPWR.n1839 0.305262
R8832 VPWR.n2138 VPWR.n2137 0.305262
R8833 VPWR.n2556 VPWR.n2555 0.305262
R8834 VPWR.n2565 VPWR.n2564 0.305262
R8835 VPWR.n2457 VPWR.n2456 0.305262
R8836 VPWR.n2460 VPWR.n2426 0.305262
R8837 VPWR.n2466 VPWR.n2465 0.305262
R8838 VPWR.n2473 VPWR.n2472 0.305262
R8839 VPWR.n2373 VPWR.n2372 0.305262
R8840 VPWR.n2059 VPWR.n2058 0.305262
R8841 VPWR.n2056 VPWR.n2055 0.305262
R8842 VPWR.n4436 VPWR.n4435 0.305262
R8843 VPWR.n4452 VPWR.n4451 0.305262
R8844 VPWR.n4467 VPWR.n4466 0.305262
R8845 VPWR.n2005 VPWR.n2004 0.305262
R8846 VPWR.n4537 VPWR.n4536 0.305262
R8847 VPWR.n3585 VPWR.n3584 0.305262
R8848 VPWR.n3594 VPWR.n3526 0.305262
R8849 VPWR.n3727 VPWR.n3726 0.305262
R8850 VPWR.n3720 VPWR.n3504 0.305262
R8851 VPWR.n3397 VPWR.n3396 0.305262
R8852 VPWR.n3407 VPWR.n3406 0.305262
R8853 VPWR.n3420 VPWR.n3419 0.305262
R8854 VPWR.n3745 VPWR.n3495 0.305262
R8855 VPWR.n3668 VPWR.n3624 0.305262
R8856 VPWR.n3663 VPWR.n3631 0.305262
R8857 VPWR.n7075 VPWR.n7074 0.305262
R8858 VPWR.n7080 VPWR.n7050 0.305262
R8859 VPWR.n7123 VPWR.n7122 0.305262
R8860 VPWR.n7119 VPWR.n7047 0.305262
R8861 VPWR.n7160 VPWR.n7159 0.305262
R8862 VPWR.n954 VPWR.n953 0.304057
R8863 VPWR.n959 VPWR.n761 0.304057
R8864 VPWR.n4780 VPWR.n4779 0.302565
R8865 VPWR.n4779 VPWR.n4778 0.302565
R8866 VPWR.n2933 VPWR.n2932 0.302565
R8867 VPWR.n852 VPWR.n850 0.295115
R8868 VPWR.n6368 VPWR.n6366 0.294492
R8869 VPWR.n1583 VPWR.n1580 0.294492
R8870 VPWR.n829 VPWR.n827 0.294041
R8871 VPWR.n5597 VPWR.n5595 0.294041
R8872 VPWR.n435 VPWR.n434 0.294041
R8873 VPWR.n4110 VPWR 0.290856
R8874 VPWR.n6125 VPWR.n6124 0.282625
R8875 VPWR VPWR.n6261 0.274365
R8876 VPWR.n7768 VPWR 0.274365
R8877 VPWR.n5115 VPWR.n1846 0.272556
R8878 VPWR.n8372 VPWR.n8371 0.264807
R8879 VPWR.n4781 VPWR.n4780 0.264807
R8880 VPWR.n3251 VPWR.n3250 0.254468
R8881 VPWR.n293 VPWR.n291 0.254468
R8882 VPWR.n5933 VPWR.n5930 0.254468
R8883 VPWR.n6501 VPWR.n6500 0.254468
R8884 VPWR.n694 VPWR.n692 0.254468
R8885 VPWR.n1593 VPWR.n1591 0.254468
R8886 VPWR.n943 VPWR.n941 0.25148
R8887 VPWR.n2639 VPWR.n2638 0.25148
R8888 VPWR.n4110 VPWR 0.250033
R8889 VPWR.n6821 VPWR.n6820 0.246654
R8890 VPWR.n980 VPWR.n979 0.246654
R8891 VPWR.n961 VPWR.n960 0.246654
R8892 VPWR.n2044 VPWR.n2043 0.246654
R8893 VPWR.n4714 VPWR.n4711 0.240185
R8894 VPWR.n8640 VPWR.n8639 0.23824
R8895 VPWR.n6188 VPWR 0.236604
R8896 VPWR.n6366 VPWR 0.236604
R8897 VPWR.n8427 VPWR 0.236604
R8898 VPWR.n1580 VPWR 0.236604
R8899 VPWR.n7675 VPWR 0.236604
R8900 VPWR VPWR.n3069 0.236604
R8901 VPWR.n850 VPWR 0.234963
R8902 VPWR VPWR.n8182 0.234145
R8903 VPWR.n827 VPWR 0.234145
R8904 VPWR.n5437 VPWR 0.234145
R8905 VPWR.n5595 VPWR 0.234145
R8906 VPWR.n435 VPWR 0.234145
R8907 VPWR.n31 VPWR 0.234145
R8908 VPWR.n3048 VPWR.n3047 0.227049
R8909 VPWR.n3080 VPWR.n3049 0.227049
R8910 VPWR.n3913 VPWR.n3912 0.227049
R8911 VPWR.n3959 VPWR.n3958 0.227049
R8912 VPWR.n7680 VPWR.n7679 0.227049
R8913 VPWR.n9061 VPWR.n9060 0.227049
R8914 VPWR.n9062 VPWR.n9061 0.227049
R8915 VPWR.n9051 VPWR.n193 0.227049
R8916 VPWR.n6193 VPWR.n6192 0.227049
R8917 VPWR.n6760 VPWR.n6759 0.227049
R8918 VPWR.n6741 VPWR.n6740 0.227049
R8919 VPWR.n8468 VPWR.n8467 0.227049
R8920 VPWR.n8486 VPWR.n8484 0.227049
R8921 VPWR.n6422 VPWR.n6421 0.227049
R8922 VPWR.n8375 VPWR.n8373 0.227049
R8923 VPWR.n5629 VPWR.n5628 0.227049
R8924 VPWR.n5636 VPWR.n455 0.227049
R8925 VPWR.n5468 VPWR.n5467 0.227049
R8926 VPWR.n491 VPWR.n490 0.227049
R8927 VPWR.n4773 VPWR.n4772 0.227049
R8928 VPWR.n4836 VPWR.n4785 0.227049
R8929 VPWR.n2720 VPWR.n2719 0.227049
R8930 VPWR.n2021 VPWR.n2020 0.227049
R8931 VPWR.n4533 VPWR.n4532 0.227049
R8932 VPWR.n4519 VPWR.n4486 0.227049
R8933 VPWR.n2932 VPWR.n2931 0.227049
R8934 VPWR.n2922 VPWR.n2886 0.227049
R8935 VPWR.n2818 VPWR.n2817 0.227049
R8936 VPWR.n2829 VPWR.n2828 0.227049
R8937 VPWR.n7393 VPWR.n7041 0.21623
R8938 VPWR.n8500 VPWR.n8499 0.21623
R8939 VPWR.n7277 VPWR.n7130 0.21623
R8940 VPWR.n2893 VPWR 0.215749
R8941 VPWR.n3993 VPWR.n3992 0.21207
R8942 VPWR.n3894 VPWR.n3893 0.21207
R8943 VPWR.n4055 VPWR.n4053 0.21207
R8944 VPWR.n3220 VPWR.n3219 0.21207
R8945 VPWR.n7665 VPWR.n7664 0.21207
R8946 VPWR.n6282 VPWR.n6231 0.21207
R8947 VPWR.n6622 VPWR.n6621 0.21207
R8948 VPWR.n6380 VPWR.n6379 0.21207
R8949 VPWR.n5686 VPWR.n5685 0.21207
R8950 VPWR.n1361 VPWR.n1360 0.21207
R8951 VPWR.n5275 VPWR.n1788 0.21207
R8952 VPWR.n1640 VPWR.n1639 0.21207
R8953 VPWR.n1657 VPWR.n1656 0.21207
R8954 VPWR.n4235 VPWR.n4234 0.21207
R8955 VPWR.n2942 VPWR.n2941 0.21207
R8956 VPWR.n3608 VPWR.n3607 0.21207
R8957 VPWR.n3614 VPWR.n3613 0.21207
R8958 VPWR.n2815 VPWR.n2814 0.21207
R8959 VPWR.n4264 VPWR.n4263 0.21207
R8960 VPWR.n2392 VPWR.n2378 0.205072
R8961 VPWR.n4566 VPWR.n4483 0.204272
R8962 VPWR.n9194 VPWR.n9193 0.203675
R8963 VPWR.n8969 VPWR.n8968 0.203675
R8964 VPWR.n8851 VPWR.n8850 0.203675
R8965 VPWR.n8739 VPWR.n8738 0.203675
R8966 VPWR.n8432 VPWR.n8431 0.203675
R8967 VPWR.n6541 VPWR.n6540 0.203675
R8968 VPWR.n6559 VPWR.n6483 0.203675
R8969 VPWR.n885 VPWR.n884 0.203675
R8970 VPWR.n661 VPWR.n660 0.203675
R8971 VPWR.n1604 VPWR.n1601 0.203675
R8972 VPWR.n2491 VPWR.n2490 0.203675
R8973 VPWR.n2048 VPWR.n2047 0.203675
R8974 VPWR.n3452 VPWR.n3451 0.203675
R8975 VPWR.n6261 VPWR 0.196835
R8976 VPWR.n6188 VPWR 0.196835
R8977 VPWR VPWR.n8427 0.196835
R8978 VPWR VPWR.n7768 0.196835
R8979 VPWR.n7675 VPWR 0.196835
R8980 VPWR.n3069 VPWR 0.196835
R8981 VPWR.n8182 VPWR 0.196385
R8982 VPWR VPWR.n31 0.196385
R8983 VPWR VPWR.n5437 0.195082
R8984 VPWR.n2064 VPWR.n2063 0.194439
R8985 VPWR.n5201 VPWR.n5200 0.1905
R8986 VPWR.n786 VPWR.n363 0.1905
R8987 VPWR.n7861 VPWR.n164 0.1905
R8988 VPWR.n5204 VPWR.n5203 0.1905
R8989 VPWR.n5856 VPWR.n5855 0.1905
R8990 VPWR.n9101 VPWR.n9100 0.1905
R8991 VPWR.n5854 VPWR.n5853 0.1905
R8992 VPWR.n9103 VPWR.n9102 0.1905
R8993 VPWR.n7712 VPWR.n7710 0.189291
R8994 VPWR.n9063 VPWR.n9062 0.189291
R8995 VPWR.n6219 VPWR.n6217 0.189291
R8996 VPWR.n625 VPWR.n595 0.188735
R8997 VPWR.n631 VPWR.n629 0.188735
R8998 VPWR.n4142 VPWR.n4141 0.185115
R8999 VPWR.n9102 VPWR 0.183019
R9000 VPWR.n5854 VPWR 0.183019
R9001 VPWR.n5202 VPWR 0.183019
R9002 VPWR.n1326 VPWR.n1322 0.180551
R9003 VPWR.n1954 VPWR.n1952 0.180294
R9004 VPWR.n6455 VPWR.n6454 0.179926
R9005 VPWR.n6454 VPWR.n6451 0.179926
R9006 VPWR.n5096 VPWR.n5094 0.179926
R9007 VPWR.n5094 VPWR.n5090 0.179926
R9008 VPWR VPWR.n6295 0.179673
R9009 VPWR VPWR.n8009 0.179673
R9010 VPWR.n5114 VPWR 0.179673
R9011 VPWR.n6042 VPWR 0.179673
R9012 VPWR.n3070 VPWR 0.179673
R9013 VPWR.n3883 VPWR 0.179673
R9014 VPWR.n3906 VPWR 0.179673
R9015 VPWR.n3513 VPWR 0.179498
R9016 VPWR.n2977 VPWR 0.179389
R9017 VPWR.n8743 VPWR 0.178345
R9018 VPWR VPWR.n5793 0.178345
R9019 VPWR VPWR.n420 0.178345
R9020 VPWR.n4100 VPWR 0.178345
R9021 VPWR VPWR.n6164 0.177989
R9022 VPWR VPWR.n224 0.177989
R9023 VPWR.n8145 VPWR 0.177989
R9024 VPWR VPWR.n8882 0.177989
R9025 VPWR.n6519 VPWR 0.177989
R9026 VPWR.n8672 VPWR 0.177989
R9027 VPWR VPWR.n8640 0.177989
R9028 VPWR.n619 VPWR 0.177989
R9029 VPWR.n863 VPWR 0.177989
R9030 VPWR.n1115 VPWR 0.177989
R9031 VPWR.n1287 VPWR 0.177989
R9032 VPWR VPWR.n5320 0.177989
R9033 VPWR.n4797 VPWR 0.177989
R9034 VPWR VPWR.n2185 0.177989
R9035 VPWR.n4925 VPWR 0.177989
R9036 VPWR.n4410 VPWR 0.177989
R9037 VPWR.n4412 VPWR 0.177989
R9038 VPWR.n4483 VPWR 0.177989
R9039 VPWR VPWR.n4504 0.177989
R9040 VPWR.n3382 VPWR 0.177989
R9041 VPWR.n7650 VPWR 0.177989
R9042 VPWR VPWR.n87 0.177989
R9043 VPWR VPWR.n81 0.177989
R9044 VPWR.n642 VPWR.n640 0.172155
R9045 VPWR.n6171 VPWR 0.171212
R9046 VPWR VPWR.n6596 0.171212
R9047 VPWR.n6495 VPWR 0.171212
R9048 VPWR VPWR.n610 0.171212
R9049 VPWR VPWR.n1286 0.171212
R9050 VPWR.n1549 VPWR 0.171212
R9051 VPWR VPWR.n2441 0.171212
R9052 VPWR.n2218 VPWR 0.171212
R9053 VPWR VPWR.n3381 0.171212
R9054 VPWR VPWR.n7649 0.171212
R9055 VPWR.n3245 VPWR 0.171212
R9056 VPWR.n4017 VPWR.n4016 0.163904
R9057 VPWR.n4025 VPWR.n4024 0.163904
R9058 VPWR VPWR.n2045 0.15779
R9059 VPWR VPWR.n1908 0.156488
R9060 VPWR.n119 VPWR.n118 0.152881
R9061 VPWR.n285 VPWR.n283 0.152881
R9062 VPWR.n285 VPWR.n284 0.152881
R9063 VPWR.n8927 VPWR.n8925 0.152881
R9064 VPWR.n8927 VPWR.n8926 0.152881
R9065 VPWR.n8569 VPWR.n8568 0.152881
R9066 VPWR.n836 VPWR.n835 0.152881
R9067 VPWR.n837 VPWR.n836 0.152881
R9068 VPWR.n884 VPWR.n883 0.152881
R9069 VPWR.n660 VPWR.n659 0.152881
R9070 VPWR.n1895 VPWR.n1894 0.152881
R9071 VPWR.n5125 VPWR.n5124 0.152881
R9072 VPWR.n4547 VPWR.n4546 0.152881
R9073 VPWR.n3627 VPWR.n3626 0.152881
R9074 VPWR.n7220 VPWR.n7218 0.152881
R9075 VPWR.n7220 VPWR.n7219 0.152881
R9076 VPWR.n7683 VPWR.n7682 0.151532
R9077 VPWR.n6196 VPWR.n6195 0.151532
R9078 VPWR.n7023 VPWR.n7022 0.151488
R9079 VPWR.n7881 VPWR.n7880 0.151488
R9080 VPWR.n8361 VPWR.n8360 0.151488
R9081 VPWR.n774 VPWR.n512 0.151488
R9082 VPWR.n5357 VPWR.n5356 0.151488
R9083 VPWR.n2598 VPWR.n2597 0.151488
R9084 VPWR.n9281 VPWR.n9280 0.151488
R9085 VPWR.n8082 VPWR.n8081 0.151488
R9086 VPWR.n8084 VPWR.n8083 0.151488
R9087 VPWR.n747 VPWR.n482 0.151488
R9088 VPWR.n1803 VPWR.n483 0.151488
R9089 VPWR.n2736 VPWR.n2735 0.151488
R9090 VPWR.n7615 VPWR.n7614 0.151488
R9091 VPWR.n6863 VPWR.n6862 0.151488
R9092 VPWR.n6584 VPWR.n6583 0.151488
R9093 VPWR.n1235 VPWR.n1234 0.151488
R9094 VPWR.n1526 VPWR.n1525 0.151488
R9095 VPWR.n2411 VPWR.n2410 0.151488
R9096 VPWR.n7138 VPWR.n7137 0.151488
R9097 VPWR.n8943 VPWR.n8942 0.151488
R9098 VPWR.n8823 VPWR.n8822 0.151488
R9099 VPWR.n5734 VPWR.n5733 0.151488
R9100 VPWR.n4595 VPWR.n4594 0.151488
R9101 VPWR.n4593 VPWR.n4592 0.151488
R9102 VPWR.n4338 VPWR.n4337 0.149872
R9103 VPWR.n9129 VPWR.n9128 0.145957
R9104 VPWR.n8511 VPWR.n8510 0.14432
R9105 VPWR.n7266 VPWR.n7265 0.14432
R9106 VPWR.n3795 VPWR.n3794 0.143372
R9107 VPWR.n3008 VPWR.n3007 0.143372
R9108 VPWR.n3362 VPWR.n3361 0.143372
R9109 VPWR.n4207 VPWR.n4206 0.143372
R9110 VPWR VPWR.n3513 0.141026
R9111 VPWR.n6295 VPWR 0.140863
R9112 VPWR.n8009 VPWR 0.140863
R9113 VPWR.n5114 VPWR 0.140863
R9114 VPWR.n2378 VPWR 0.140863
R9115 VPWR.n6042 VPWR 0.140863
R9116 VPWR.n3070 VPWR 0.140863
R9117 VPWR VPWR.n3883 0.140863
R9118 VPWR VPWR.n3906 0.140863
R9119 VPWR.n6164 VPWR 0.140584
R9120 VPWR.n224 VPWR 0.140584
R9121 VPWR.n8145 VPWR 0.140584
R9122 VPWR.n8882 VPWR 0.140584
R9123 VPWR VPWR.n6519 0.140584
R9124 VPWR.n8672 VPWR 0.140584
R9125 VPWR VPWR.n619 0.140584
R9126 VPWR VPWR.n863 0.140584
R9127 VPWR.n1287 VPWR 0.140584
R9128 VPWR.n5320 VPWR 0.140584
R9129 VPWR.n4797 VPWR 0.140584
R9130 VPWR.n2185 VPWR 0.140584
R9131 VPWR.n4925 VPWR 0.140584
R9132 VPWR VPWR.n4410 0.140584
R9133 VPWR.n4412 VPWR 0.140584
R9134 VPWR.n4504 VPWR 0.140584
R9135 VPWR.n3382 VPWR 0.140584
R9136 VPWR.n2893 VPWR 0.140584
R9137 VPWR.n7650 VPWR 0.140584
R9138 VPWR.n87 VPWR 0.140584
R9139 VPWR.n81 VPWR 0.140584
R9140 VPWR.n8743 VPWR 0.140228
R9141 VPWR.n5793 VPWR 0.140228
R9142 VPWR.n420 VPWR 0.140228
R9143 VPWR.n4100 VPWR 0.140228
R9144 VPWR VPWR.n1115 0.139282
R9145 VPWR.n9139 VPWR.n9138 0.138115
R9146 VPWR.n5200 VPWR.n5199 0.125931
R9147 VPWR.n5204 VPWR.n1804 0.125931
R9148 VPWR.n2195 VPWR.n1805 0.125931
R9149 VPWR.n4879 VPWR.n4878 0.125931
R9150 VPWR.n4151 VPWR.n4150 0.123577
R9151 VPWR.n6130 VPWR.n6129 0.123577
R9152 VPWR.n6871 VPWR.n6870 0.123577
R9153 VPWR.n6793 VPWR.n6792 0.123577
R9154 VPWR.n6262 VPWR 0.120655
R9155 VPWR.n6185 VPWR 0.120655
R9156 VPWR.n6187 VPWR 0.120655
R9157 VPWR VPWR.n6762 0.120655
R9158 VPWR VPWR.n6692 0.120655
R9159 VPWR.n1950 VPWR 0.120655
R9160 VPWR.n1952 VPWR 0.120655
R9161 VPWR VPWR.n2023 0.120655
R9162 VPWR.n3636 VPWR 0.120655
R9163 VPWR.n7767 VPWR 0.120655
R9164 VPWR.n4005 VPWR 0.120655
R9165 VPWR.n4027 VPWR 0.120655
R9166 VPWR.n3907 VPWR 0.120655
R9167 VPWR.n6185 VPWR 0.120399
R9168 VPWR.n2023 VPWR 0.120399
R9169 VPWR.n6181 VPWR.n6178 0.120292
R9170 VPWR.n6183 VPWR.n6181 0.120292
R9171 VPWR.n6199 VPWR.n6194 0.120292
R9172 VPWR.n6311 VPWR.n6310 0.120292
R9173 VPWR.n6310 VPWR.n6308 0.120292
R9174 VPWR.n6308 VPWR.n6306 0.120292
R9175 VPWR.n6306 VPWR.n6303 0.120292
R9176 VPWR.n6303 VPWR.n6301 0.120292
R9177 VPWR.n6301 VPWR.n6299 0.120292
R9178 VPWR.n6286 VPWR.n6285 0.120292
R9179 VPWR.n6285 VPWR.n6283 0.120292
R9180 VPWR.n6279 VPWR.n6278 0.120292
R9181 VPWR.n6278 VPWR.n6273 0.120292
R9182 VPWR.n6270 VPWR.n6269 0.120292
R9183 VPWR.n6269 VPWR.n6266 0.120292
R9184 VPWR.n6260 VPWR.n6253 0.120292
R9185 VPWR.n6253 VPWR.n6251 0.120292
R9186 VPWR.n6251 VPWR.n6249 0.120292
R9187 VPWR.n6249 VPWR.n6247 0.120292
R9188 VPWR.n6247 VPWR.n6244 0.120292
R9189 VPWR.n6244 VPWR.n6242 0.120292
R9190 VPWR.n6242 VPWR.n6241 0.120292
R9191 VPWR.n7951 VPWR.n7950 0.120292
R9192 VPWR.n7950 VPWR.n7947 0.120292
R9193 VPWR.n7947 VPWR.n7945 0.120292
R9194 VPWR.n7945 VPWR.n7941 0.120292
R9195 VPWR.n7941 VPWR.n7938 0.120292
R9196 VPWR.n7938 VPWR.n7936 0.120292
R9197 VPWR.n7936 VPWR.n7934 0.120292
R9198 VPWR.n7934 VPWR.n7931 0.120292
R9199 VPWR.n7931 VPWR.n7929 0.120292
R9200 VPWR.n7929 VPWR.n7925 0.120292
R9201 VPWR.n7925 VPWR.n7923 0.120292
R9202 VPWR.n7920 VPWR.n7919 0.120292
R9203 VPWR.n7919 VPWR.n7918 0.120292
R9204 VPWR.n7918 VPWR.n7914 0.120292
R9205 VPWR.n7914 VPWR.n7912 0.120292
R9206 VPWR.n7912 VPWR.n7911 0.120292
R9207 VPWR.n7911 VPWR.n7910 0.120292
R9208 VPWR.n8020 VPWR.n8018 0.120292
R9209 VPWR.n8024 VPWR.n8020 0.120292
R9210 VPWR.n8026 VPWR.n8024 0.120292
R9211 VPWR.n8029 VPWR.n8026 0.120292
R9212 VPWR.n8031 VPWR.n8029 0.120292
R9213 VPWR.n8033 VPWR.n8031 0.120292
R9214 VPWR.n8036 VPWR.n8033 0.120292
R9215 VPWR.n8038 VPWR.n8036 0.120292
R9216 VPWR.n8040 VPWR.n8038 0.120292
R9217 VPWR.n8042 VPWR.n8040 0.120292
R9218 VPWR.n8043 VPWR.n8042 0.120292
R9219 VPWR.n8047 VPWR.n8046 0.120292
R9220 VPWR.n8054 VPWR.n8051 0.120292
R9221 VPWR.n8056 VPWR.n8054 0.120292
R9222 VPWR.n8058 VPWR.n8056 0.120292
R9223 VPWR.n9065 VPWR.n9059 0.120292
R9224 VPWR.n9059 VPWR.n9056 0.120292
R9225 VPWR.n9056 VPWR.n9054 0.120292
R9226 VPWR.n9054 VPWR.n9052 0.120292
R9227 VPWR.n8982 VPWR.n8980 0.120292
R9228 VPWR.n8983 VPWR.n8982 0.120292
R9229 VPWR.n8992 VPWR.n8988 0.120292
R9230 VPWR.n8994 VPWR.n8992 0.120292
R9231 VPWR.n8996 VPWR.n8994 0.120292
R9232 VPWR.n8999 VPWR.n8996 0.120292
R9233 VPWR.n9002 VPWR.n8999 0.120292
R9234 VPWR.n9004 VPWR.n9002 0.120292
R9235 VPWR.n9008 VPWR.n9004 0.120292
R9236 VPWR.n9010 VPWR.n9008 0.120292
R9237 VPWR.n9012 VPWR.n9010 0.120292
R9238 VPWR.n9014 VPWR.n9012 0.120292
R9239 VPWR.n9017 VPWR.n9014 0.120292
R9240 VPWR.n9023 VPWR.n9021 0.120292
R9241 VPWR.n9025 VPWR.n9023 0.120292
R9242 VPWR.n9027 VPWR.n9025 0.120292
R9243 VPWR.n9028 VPWR.n9027 0.120292
R9244 VPWR.n9035 VPWR.n9031 0.120292
R9245 VPWR.n9037 VPWR.n9035 0.120292
R9246 VPWR.n9040 VPWR.n9037 0.120292
R9247 VPWR.n9042 VPWR.n9040 0.120292
R9248 VPWR.n9044 VPWR.n9042 0.120292
R9249 VPWR.n9045 VPWR.n9044 0.120292
R9250 VPWR.n8971 VPWR.n8970 0.120292
R9251 VPWR.n257 VPWR.n255 0.120292
R9252 VPWR.n255 VPWR.n254 0.120292
R9253 VPWR.n254 VPWR.n252 0.120292
R9254 VPWR.n252 VPWR.n249 0.120292
R9255 VPWR.n249 VPWR.n246 0.120292
R9256 VPWR.n240 VPWR.n239 0.120292
R9257 VPWR.n239 VPWR.n238 0.120292
R9258 VPWR.n238 VPWR.n237 0.120292
R9259 VPWR.n237 VPWR.n234 0.120292
R9260 VPWR.n234 VPWR.n232 0.120292
R9261 VPWR.n227 VPWR.n225 0.120292
R9262 VPWR.n6605 VPWR.n6603 0.120292
R9263 VPWR.n6609 VPWR.n6605 0.120292
R9264 VPWR.n6613 VPWR.n6609 0.120292
R9265 VPWR.n6623 VPWR.n6619 0.120292
R9266 VPWR.n6625 VPWR.n6623 0.120292
R9267 VPWR.n6629 VPWR.n6625 0.120292
R9268 VPWR.n6631 VPWR.n6629 0.120292
R9269 VPWR.n6632 VPWR.n6631 0.120292
R9270 VPWR.n6639 VPWR.n6637 0.120292
R9271 VPWR.n6779 VPWR.n6778 0.120292
R9272 VPWR.n6778 VPWR.n6776 0.120292
R9273 VPWR.n6776 VPWR.n6774 0.120292
R9274 VPWR.n6774 VPWR.n6771 0.120292
R9275 VPWR.n6771 VPWR.n6769 0.120292
R9276 VPWR.n6769 VPWR.n6767 0.120292
R9277 VPWR.n6761 VPWR.n6749 0.120292
R9278 VPWR.n6749 VPWR.n6748 0.120292
R9279 VPWR.n6748 VPWR.n6747 0.120292
R9280 VPWR.n6747 VPWR.n6745 0.120292
R9281 VPWR.n6745 VPWR.n6742 0.120292
R9282 VPWR.n6739 VPWR.n6737 0.120292
R9283 VPWR.n6737 VPWR.n6735 0.120292
R9284 VPWR.n6735 VPWR.n6731 0.120292
R9285 VPWR.n6731 VPWR.n6729 0.120292
R9286 VPWR.n6729 VPWR.n6727 0.120292
R9287 VPWR.n6724 VPWR.n6723 0.120292
R9288 VPWR.n6723 VPWR.n6720 0.120292
R9289 VPWR.n6720 VPWR.n6718 0.120292
R9290 VPWR.n6718 VPWR.n6716 0.120292
R9291 VPWR.n6716 VPWR.n6713 0.120292
R9292 VPWR.n6713 VPWR.n6709 0.120292
R9293 VPWR.n6709 VPWR.n6707 0.120292
R9294 VPWR.n6707 VPWR.n6703 0.120292
R9295 VPWR.n6703 VPWR.n6701 0.120292
R9296 VPWR.n6701 VPWR.n6699 0.120292
R9297 VPWR.n6699 VPWR.n6697 0.120292
R9298 VPWR.n8342 VPWR.n8339 0.120292
R9299 VPWR.n8339 VPWR.n8335 0.120292
R9300 VPWR.n8335 VPWR.n8333 0.120292
R9301 VPWR.n8330 VPWR.n8329 0.120292
R9302 VPWR.n8329 VPWR.n8326 0.120292
R9303 VPWR.n8326 VPWR.n8322 0.120292
R9304 VPWR.n8322 VPWR.n8318 0.120292
R9305 VPWR.n8314 VPWR.n8313 0.120292
R9306 VPWR.n8313 VPWR.n8312 0.120292
R9307 VPWR.n8312 VPWR.n8311 0.120292
R9308 VPWR.n8311 VPWR.n8309 0.120292
R9309 VPWR.n8309 VPWR.n8307 0.120292
R9310 VPWR.n8302 VPWR.n8300 0.120292
R9311 VPWR.n8300 VPWR.n8294 0.120292
R9312 VPWR.n8287 VPWR.n8286 0.120292
R9313 VPWR.n8286 VPWR.n8285 0.120292
R9314 VPWR.n8285 VPWR.n8284 0.120292
R9315 VPWR.n8281 VPWR.n8280 0.120292
R9316 VPWR.n8280 VPWR.n8278 0.120292
R9317 VPWR.n8278 VPWR.n8276 0.120292
R9318 VPWR.n8276 VPWR.n8274 0.120292
R9319 VPWR.n8274 VPWR.n8271 0.120292
R9320 VPWR.n8271 VPWR.n8268 0.120292
R9321 VPWR.n8268 VPWR.n8266 0.120292
R9322 VPWR.n8266 VPWR.n8264 0.120292
R9323 VPWR.n8264 VPWR.n8262 0.120292
R9324 VPWR.n8198 VPWR.n8191 0.120292
R9325 VPWR.n8191 VPWR.n8190 0.120292
R9326 VPWR.n8190 VPWR.n8189 0.120292
R9327 VPWR.n8132 VPWR.n8130 0.120292
R9328 VPWR.n8134 VPWR.n8132 0.120292
R9329 VPWR.n8136 VPWR.n8134 0.120292
R9330 VPWR.n8139 VPWR.n8136 0.120292
R9331 VPWR.n8140 VPWR.n8139 0.120292
R9332 VPWR.n8144 VPWR.n8143 0.120292
R9333 VPWR.n8155 VPWR.n8153 0.120292
R9334 VPWR.n8158 VPWR.n8155 0.120292
R9335 VPWR.n8161 VPWR.n8158 0.120292
R9336 VPWR.n8163 VPWR.n8161 0.120292
R9337 VPWR.n8164 VPWR.n8163 0.120292
R9338 VPWR.n8165 VPWR.n8164 0.120292
R9339 VPWR.n8166 VPWR.n8165 0.120292
R9340 VPWR.n8172 VPWR.n8170 0.120292
R9341 VPWR.n8174 VPWR.n8172 0.120292
R9342 VPWR.n8176 VPWR.n8174 0.120292
R9343 VPWR.n8180 VPWR.n8176 0.120292
R9344 VPWR.n8181 VPWR.n8180 0.120292
R9345 VPWR.n8916 VPWR.n8914 0.120292
R9346 VPWR.n8914 VPWR.n8908 0.120292
R9347 VPWR.n8908 VPWR.n8906 0.120292
R9348 VPWR.n8903 VPWR.n8902 0.120292
R9349 VPWR.n8902 VPWR.n8901 0.120292
R9350 VPWR.n8901 VPWR.n8900 0.120292
R9351 VPWR.n8894 VPWR.n8893 0.120292
R9352 VPWR.n8892 VPWR.n8890 0.120292
R9353 VPWR.n8885 VPWR.n8884 0.120292
R9354 VPWR.n8884 VPWR.n8883 0.120292
R9355 VPWR.n6504 VPWR.n6503 0.120292
R9356 VPWR.n6505 VPWR.n6504 0.120292
R9357 VPWR.n6513 VPWR.n6505 0.120292
R9358 VPWR.n6526 VPWR.n6524 0.120292
R9359 VPWR.n6529 VPWR.n6526 0.120292
R9360 VPWR.n6531 VPWR.n6529 0.120292
R9361 VPWR.n6532 VPWR.n6531 0.120292
R9362 VPWR.n6460 VPWR.n6459 0.120292
R9363 VPWR.n6459 VPWR.n6457 0.120292
R9364 VPWR.n6457 VPWR.n6455 0.120292
R9365 VPWR.n6370 VPWR.n6368 0.120292
R9366 VPWR.n6373 VPWR.n6370 0.120292
R9367 VPWR.n6374 VPWR.n6373 0.120292
R9368 VPWR.n6383 VPWR.n6382 0.120292
R9369 VPWR.n6391 VPWR.n6388 0.120292
R9370 VPWR.n6395 VPWR.n6391 0.120292
R9371 VPWR.n6397 VPWR.n6395 0.120292
R9372 VPWR.n6399 VPWR.n6397 0.120292
R9373 VPWR.n6401 VPWR.n6399 0.120292
R9374 VPWR.n6403 VPWR.n6401 0.120292
R9375 VPWR.n6405 VPWR.n6403 0.120292
R9376 VPWR.n6406 VPWR.n6405 0.120292
R9377 VPWR.n6414 VPWR.n6413 0.120292
R9378 VPWR.n6419 VPWR.n6418 0.120292
R9379 VPWR.n6443 VPWR.n6442 0.120292
R9380 VPWR.n8435 VPWR.n8434 0.120292
R9381 VPWR.n8447 VPWR.n8446 0.120292
R9382 VPWR.n8448 VPWR.n8447 0.120292
R9383 VPWR.n8450 VPWR.n8448 0.120292
R9384 VPWR.n8460 VPWR.n8450 0.120292
R9385 VPWR.n8472 VPWR.n8469 0.120292
R9386 VPWR.n8475 VPWR.n8472 0.120292
R9387 VPWR.n8477 VPWR.n8475 0.120292
R9388 VPWR.n8479 VPWR.n8477 0.120292
R9389 VPWR.n8480 VPWR.n8479 0.120292
R9390 VPWR.n8481 VPWR.n8480 0.120292
R9391 VPWR.n8487 VPWR.n8481 0.120292
R9392 VPWR.n8504 VPWR.n8501 0.120292
R9393 VPWR.n8509 VPWR.n8504 0.120292
R9394 VPWR.n8512 VPWR.n8509 0.120292
R9395 VPWR.n8514 VPWR.n8512 0.120292
R9396 VPWR.n8601 VPWR.n8600 0.120292
R9397 VPWR.n8605 VPWR.n8601 0.120292
R9398 VPWR.n8606 VPWR.n8605 0.120292
R9399 VPWR.n8671 VPWR.n8670 0.120292
R9400 VPWR.n8670 VPWR.n8669 0.120292
R9401 VPWR.n8669 VPWR.n8668 0.120292
R9402 VPWR.n8668 VPWR.n8665 0.120292
R9403 VPWR.n8665 VPWR.n8663 0.120292
R9404 VPWR.n8663 VPWR.n8659 0.120292
R9405 VPWR.n8659 VPWR.n8657 0.120292
R9406 VPWR.n8654 VPWR.n8653 0.120292
R9407 VPWR.n8653 VPWR.n8651 0.120292
R9408 VPWR.n8651 VPWR.n8646 0.120292
R9409 VPWR.n8646 VPWR.n8644 0.120292
R9410 VPWR.n8639 VPWR.n8636 0.120292
R9411 VPWR.n8636 VPWR.n8635 0.120292
R9412 VPWR.n8635 VPWR.n8634 0.120292
R9413 VPWR.n8631 VPWR.n8630 0.120292
R9414 VPWR.n8688 VPWR.n8685 0.120292
R9415 VPWR.n8692 VPWR.n8688 0.120292
R9416 VPWR.n8788 VPWR.n8785 0.120292
R9417 VPWR.n8785 VPWR.n8782 0.120292
R9418 VPWR.n8782 VPWR.n8780 0.120292
R9419 VPWR.n8780 VPWR.n8776 0.120292
R9420 VPWR.n8776 VPWR.n8774 0.120292
R9421 VPWR.n8770 VPWR.n8769 0.120292
R9422 VPWR.n8765 VPWR.n8764 0.120292
R9423 VPWR.n8759 VPWR.n8751 0.120292
R9424 VPWR.n8751 VPWR.n8750 0.120292
R9425 VPWR.n8750 VPWR.n8749 0.120292
R9426 VPWR.n618 VPWR.n614 0.120292
R9427 VPWR.n634 VPWR.n632 0.120292
R9428 VPWR.n636 VPWR.n634 0.120292
R9429 VPWR.n637 VPWR.n636 0.120292
R9430 VPWR.n646 VPWR.n643 0.120292
R9431 VPWR.n1224 VPWR.n1223 0.120292
R9432 VPWR.n1223 VPWR.n1222 0.120292
R9433 VPWR.n1222 VPWR.n1220 0.120292
R9434 VPWR.n1220 VPWR.n1218 0.120292
R9435 VPWR.n1218 VPWR.n1212 0.120292
R9436 VPWR.n1212 VPWR.n1210 0.120292
R9437 VPWR.n831 VPWR.n829 0.120292
R9438 VPWR.n833 VPWR.n831 0.120292
R9439 VPWR.n838 VPWR.n833 0.120292
R9440 VPWR.n847 VPWR.n845 0.120292
R9441 VPWR.n853 VPWR.n852 0.120292
R9442 VPWR.n854 VPWR.n853 0.120292
R9443 VPWR.n855 VPWR.n854 0.120292
R9444 VPWR.n860 VPWR.n858 0.120292
R9445 VPWR.n862 VPWR.n860 0.120292
R9446 VPWR.n939 VPWR.n937 0.120292
R9447 VPWR.n944 VPWR.n939 0.120292
R9448 VPWR.n945 VPWR.n944 0.120292
R9449 VPWR.n956 VPWR.n955 0.120292
R9450 VPWR.n957 VPWR.n956 0.120292
R9451 VPWR.n958 VPWR.n957 0.120292
R9452 VPWR.n963 VPWR.n962 0.120292
R9453 VPWR.n964 VPWR.n963 0.120292
R9454 VPWR.n974 VPWR.n969 0.120292
R9455 VPWR.n977 VPWR.n974 0.120292
R9456 VPWR.n981 VPWR.n977 0.120292
R9457 VPWR.n984 VPWR.n981 0.120292
R9458 VPWR.n987 VPWR.n984 0.120292
R9459 VPWR.n989 VPWR.n987 0.120292
R9460 VPWR.n990 VPWR.n989 0.120292
R9461 VPWR.n999 VPWR.n994 0.120292
R9462 VPWR.n1002 VPWR.n999 0.120292
R9463 VPWR.n1004 VPWR.n1002 0.120292
R9464 VPWR.n1007 VPWR.n1004 0.120292
R9465 VPWR.n1009 VPWR.n1007 0.120292
R9466 VPWR.n1011 VPWR.n1009 0.120292
R9467 VPWR.n1013 VPWR.n1011 0.120292
R9468 VPWR.n1016 VPWR.n1013 0.120292
R9469 VPWR.n1020 VPWR.n1016 0.120292
R9470 VPWR.n1021 VPWR.n1020 0.120292
R9471 VPWR.n1028 VPWR.n1027 0.120292
R9472 VPWR.n1029 VPWR.n1028 0.120292
R9473 VPWR.n1030 VPWR.n1029 0.120292
R9474 VPWR.n1038 VPWR.n1036 0.120292
R9475 VPWR.n1114 VPWR.n1112 0.120292
R9476 VPWR.n1119 VPWR.n1118 0.120292
R9477 VPWR.n1118 VPWR.n1117 0.120292
R9478 VPWR.n1135 VPWR.n1134 0.120292
R9479 VPWR.n1144 VPWR.n1139 0.120292
R9480 VPWR.n1146 VPWR.n1144 0.120292
R9481 VPWR.n1152 VPWR.n1146 0.120292
R9482 VPWR.n1154 VPWR.n1152 0.120292
R9483 VPWR.n1158 VPWR.n1154 0.120292
R9484 VPWR.n1160 VPWR.n1158 0.120292
R9485 VPWR.n1164 VPWR.n1160 0.120292
R9486 VPWR.n1168 VPWR.n1164 0.120292
R9487 VPWR.n1172 VPWR.n1168 0.120292
R9488 VPWR.n1175 VPWR.n1172 0.120292
R9489 VPWR.n1177 VPWR.n1175 0.120292
R9490 VPWR.n1180 VPWR.n1177 0.120292
R9491 VPWR.n1182 VPWR.n1180 0.120292
R9492 VPWR.n1187 VPWR.n1182 0.120292
R9493 VPWR.n1189 VPWR.n1187 0.120292
R9494 VPWR.n1192 VPWR.n1189 0.120292
R9495 VPWR.n1193 VPWR.n1192 0.120292
R9496 VPWR.n1194 VPWR.n1193 0.120292
R9497 VPWR.n1198 VPWR.n1195 0.120292
R9498 VPWR.n1195 VPWR.n387 0.120292
R9499 VPWR.n5743 VPWR.n387 0.120292
R9500 VPWR.n5825 VPWR.n5824 0.120292
R9501 VPWR.n5824 VPWR.n5822 0.120292
R9502 VPWR.n5822 VPWR.n5821 0.120292
R9503 VPWR.n5821 VPWR.n5819 0.120292
R9504 VPWR.n5815 VPWR.n5814 0.120292
R9505 VPWR.n5814 VPWR.n5808 0.120292
R9506 VPWR.n5808 VPWR.n5806 0.120292
R9507 VPWR.n5803 VPWR.n5802 0.120292
R9508 VPWR.n5802 VPWR.n5800 0.120292
R9509 VPWR.n5796 VPWR.n5795 0.120292
R9510 VPWR.n5795 VPWR.n5794 0.120292
R9511 VPWR.n1285 VPWR.n1275 0.120292
R9512 VPWR.n1299 VPWR.n1275 0.120292
R9513 VPWR.n1301 VPWR.n1300 0.120292
R9514 VPWR.n1302 VPWR.n1301 0.120292
R9515 VPWR.n1311 VPWR.n1308 0.120292
R9516 VPWR.n1313 VPWR.n1311 0.120292
R9517 VPWR.n1317 VPWR.n1313 0.120292
R9518 VPWR.n1516 VPWR.n1512 0.120292
R9519 VPWR.n1512 VPWR.n1510 0.120292
R9520 VPWR.n1510 VPWR.n1508 0.120292
R9521 VPWR.n1508 VPWR.n1504 0.120292
R9522 VPWR.n1504 VPWR.n1501 0.120292
R9523 VPWR.n1497 VPWR.n1496 0.120292
R9524 VPWR.n1493 VPWR.n1492 0.120292
R9525 VPWR.n1492 VPWR.n1490 0.120292
R9526 VPWR.n1486 VPWR.n1485 0.120292
R9527 VPWR.n1485 VPWR.n1481 0.120292
R9528 VPWR.n1481 VPWR.n1479 0.120292
R9529 VPWR.n1479 VPWR.n1477 0.120292
R9530 VPWR.n1477 VPWR.n1474 0.120292
R9531 VPWR.n1474 VPWR.n1471 0.120292
R9532 VPWR.n1471 VPWR.n1469 0.120292
R9533 VPWR.n1469 VPWR.n1465 0.120292
R9534 VPWR.n1465 VPWR.n1463 0.120292
R9535 VPWR.n1463 VPWR.n1461 0.120292
R9536 VPWR.n1461 VPWR.n1459 0.120292
R9537 VPWR.n1456 VPWR.n1455 0.120292
R9538 VPWR.n1455 VPWR.n1453 0.120292
R9539 VPWR.n1453 VPWR.n1452 0.120292
R9540 VPWR.n1452 VPWR.n1451 0.120292
R9541 VPWR.n1447 VPWR.n1442 0.120292
R9542 VPWR.n1438 VPWR.n1437 0.120292
R9543 VPWR.n1432 VPWR.n1431 0.120292
R9544 VPWR.n5406 VPWR.n5404 0.120292
R9545 VPWR.n5410 VPWR.n5406 0.120292
R9546 VPWR.n5411 VPWR.n5410 0.120292
R9547 VPWR.n5416 VPWR.n5414 0.120292
R9548 VPWR.n5420 VPWR.n5416 0.120292
R9549 VPWR.n5424 VPWR.n5420 0.120292
R9550 VPWR.n5426 VPWR.n5424 0.120292
R9551 VPWR.n5430 VPWR.n5426 0.120292
R9552 VPWR.n5431 VPWR.n5430 0.120292
R9553 VPWR.n5439 VPWR.n5438 0.120292
R9554 VPWR.n5456 VPWR.n5455 0.120292
R9555 VPWR.n5465 VPWR.n5464 0.120292
R9556 VPWR.n5471 VPWR.n5469 0.120292
R9557 VPWR.n5475 VPWR.n5471 0.120292
R9558 VPWR.n5477 VPWR.n5475 0.120292
R9559 VPWR.n5480 VPWR.n5477 0.120292
R9560 VPWR.n5481 VPWR.n5480 0.120292
R9561 VPWR.n5482 VPWR.n5481 0.120292
R9562 VPWR.n5483 VPWR.n5482 0.120292
R9563 VPWR.n5488 VPWR.n5487 0.120292
R9564 VPWR.n5584 VPWR.n5580 0.120292
R9565 VPWR.n5586 VPWR.n5584 0.120292
R9566 VPWR.n5588 VPWR.n5586 0.120292
R9567 VPWR.n5589 VPWR.n5588 0.120292
R9568 VPWR.n5600 VPWR.n5597 0.120292
R9569 VPWR.n5602 VPWR.n5600 0.120292
R9570 VPWR.n5603 VPWR.n5602 0.120292
R9571 VPWR.n462 VPWR.n461 0.120292
R9572 VPWR.n5611 VPWR.n5610 0.120292
R9573 VPWR.n5618 VPWR.n5616 0.120292
R9574 VPWR.n5619 VPWR.n5618 0.120292
R9575 VPWR.n5625 VPWR.n5624 0.120292
R9576 VPWR.n5632 VPWR.n5630 0.120292
R9577 VPWR.n5633 VPWR.n5632 0.120292
R9578 VPWR.n5634 VPWR.n5633 0.120292
R9579 VPWR.n5635 VPWR.n5634 0.120292
R9580 VPWR.n5649 VPWR.n5644 0.120292
R9581 VPWR.n5651 VPWR.n5649 0.120292
R9582 VPWR.n5653 VPWR.n5651 0.120292
R9583 VPWR.n450 VPWR.n447 0.120292
R9584 VPWR.n441 VPWR.n440 0.120292
R9585 VPWR.n434 VPWR.n432 0.120292
R9586 VPWR.n432 VPWR.n430 0.120292
R9587 VPWR.n430 VPWR.n428 0.120292
R9588 VPWR.n423 VPWR.n422 0.120292
R9589 VPWR.n422 VPWR.n421 0.120292
R9590 VPWR.n1556 VPWR.n1555 0.120292
R9591 VPWR.n1561 VPWR.n1559 0.120292
R9592 VPWR.n1567 VPWR.n1561 0.120292
R9593 VPWR.n1568 VPWR.n1567 0.120292
R9594 VPWR.n1573 VPWR.n1572 0.120292
R9595 VPWR.n1579 VPWR.n1576 0.120292
R9596 VPWR.n1586 VPWR.n1583 0.120292
R9597 VPWR.n1646 VPWR.n1644 0.120292
R9598 VPWR.n1649 VPWR.n1646 0.120292
R9599 VPWR.n1652 VPWR.n1649 0.120292
R9600 VPWR.n1654 VPWR.n1652 0.120292
R9601 VPWR.n1658 VPWR.n1654 0.120292
R9602 VPWR.n1659 VPWR.n1658 0.120292
R9603 VPWR.n1666 VPWR.n1663 0.120292
R9604 VPWR.n1667 VPWR.n1666 0.120292
R9605 VPWR.n1674 VPWR.n1672 0.120292
R9606 VPWR.n1681 VPWR.n1674 0.120292
R9607 VPWR.n1682 VPWR.n1681 0.120292
R9608 VPWR.n1689 VPWR.n1688 0.120292
R9609 VPWR.n1691 VPWR.n1689 0.120292
R9610 VPWR.n1693 VPWR.n1691 0.120292
R9611 VPWR.n1696 VPWR.n1693 0.120292
R9612 VPWR.n1698 VPWR.n1696 0.120292
R9613 VPWR.n1700 VPWR.n1698 0.120292
R9614 VPWR.n1701 VPWR.n1700 0.120292
R9615 VPWR.n1707 VPWR.n1705 0.120292
R9616 VPWR.n1708 VPWR.n1707 0.120292
R9617 VPWR.n1717 VPWR.n552 0.120292
R9618 VPWR.n1719 VPWR.n1718 0.120292
R9619 VPWR.n1720 VPWR.n1719 0.120292
R9620 VPWR.n1724 VPWR.n550 0.120292
R9621 VPWR.n1772 VPWR.n1770 0.120292
R9622 VPWR.n5322 VPWR.n5321 0.120292
R9623 VPWR.n5316 VPWR.n5315 0.120292
R9624 VPWR.n5311 VPWR.n5310 0.120292
R9625 VPWR.n5310 VPWR.n5306 0.120292
R9626 VPWR.n5306 VPWR.n5302 0.120292
R9627 VPWR.n5302 VPWR.n5301 0.120292
R9628 VPWR.n5301 VPWR.n5300 0.120292
R9629 VPWR.n5300 VPWR.n5298 0.120292
R9630 VPWR.n5298 VPWR.n5297 0.120292
R9631 VPWR.n5293 VPWR.n5292 0.120292
R9632 VPWR.n5287 VPWR.n5285 0.120292
R9633 VPWR.n5285 VPWR.n5284 0.120292
R9634 VPWR.n5280 VPWR.n5279 0.120292
R9635 VPWR.n5274 VPWR.n5273 0.120292
R9636 VPWR.n5273 VPWR.n5271 0.120292
R9637 VPWR.n5271 VPWR.n5269 0.120292
R9638 VPWR.n5269 VPWR.n5267 0.120292
R9639 VPWR.n5267 VPWR.n5264 0.120292
R9640 VPWR.n5264 VPWR.n5262 0.120292
R9641 VPWR.n5262 VPWR.n5260 0.120292
R9642 VPWR.n5260 VPWR.n5258 0.120292
R9643 VPWR.n5258 VPWR.n5256 0.120292
R9644 VPWR.n4682 VPWR.n4676 0.120292
R9645 VPWR.n4683 VPWR.n4682 0.120292
R9646 VPWR.n4762 VPWR.n4761 0.120292
R9647 VPWR.n4761 VPWR.n4759 0.120292
R9648 VPWR.n4747 VPWR.n4746 0.120292
R9649 VPWR.n4746 VPWR.n4742 0.120292
R9650 VPWR.n4742 VPWR.n4740 0.120292
R9651 VPWR.n4740 VPWR.n4735 0.120292
R9652 VPWR.n4735 VPWR.n4734 0.120292
R9653 VPWR.n4734 VPWR.n4728 0.120292
R9654 VPWR.n4722 VPWR.n4721 0.120292
R9655 VPWR.n4721 VPWR.n4719 0.120292
R9656 VPWR.n4719 VPWR.n4718 0.120292
R9657 VPWR.n4718 VPWR.n4717 0.120292
R9658 VPWR.n4717 VPWR.n4716 0.120292
R9659 VPWR.n4776 VPWR.n4774 0.120292
R9660 VPWR.n4784 VPWR.n4776 0.120292
R9661 VPWR.n4842 VPWR.n4837 0.120292
R9662 VPWR.n4834 VPWR.n4833 0.120292
R9663 VPWR.n4833 VPWR.n4829 0.120292
R9664 VPWR.n4821 VPWR.n4820 0.120292
R9665 VPWR.n4815 VPWR.n4811 0.120292
R9666 VPWR.n4811 VPWR.n4809 0.120292
R9667 VPWR.n4809 VPWR.n4805 0.120292
R9668 VPWR.n4805 VPWR.n4803 0.120292
R9669 VPWR.n2447 VPWR.n2446 0.120292
R9670 VPWR.n2453 VPWR.n2427 0.120292
R9671 VPWR.n2462 VPWR.n2427 0.120292
R9672 VPWR.n2470 VPWR.n2424 0.120292
R9673 VPWR.n2482 VPWR.n2476 0.120292
R9674 VPWR.n2552 VPWR.n2551 0.120292
R9675 VPWR.n2560 VPWR.n2559 0.120292
R9676 VPWR.n2559 VPWR.n2558 0.120292
R9677 VPWR.n2184 VPWR.n2180 0.120292
R9678 VPWR.n2180 VPWR.n2178 0.120292
R9679 VPWR.n2178 VPWR.n2174 0.120292
R9680 VPWR.n2174 VPWR.n2172 0.120292
R9681 VPWR.n2172 VPWR.n2169 0.120292
R9682 VPWR.n2169 VPWR.n2167 0.120292
R9683 VPWR.n2167 VPWR.n2164 0.120292
R9684 VPWR.n2164 VPWR.n2162 0.120292
R9685 VPWR.n2162 VPWR.n2158 0.120292
R9686 VPWR.n2158 VPWR.n2156 0.120292
R9687 VPWR.n2156 VPWR.n2154 0.120292
R9688 VPWR.n2151 VPWR.n2150 0.120292
R9689 VPWR.n2150 VPWR.n2145 0.120292
R9690 VPWR.n2145 VPWR.n2143 0.120292
R9691 VPWR.n2143 VPWR.n2142 0.120292
R9692 VPWR.n2142 VPWR.n2141 0.120292
R9693 VPWR.n2135 VPWR.n2134 0.120292
R9694 VPWR.n2134 VPWR.n2133 0.120292
R9695 VPWR.n2133 VPWR.n2132 0.120292
R9696 VPWR.n2575 VPWR.n2574 0.120292
R9697 VPWR.n5159 VPWR.n5157 0.120292
R9698 VPWR.n5157 VPWR.n5156 0.120292
R9699 VPWR.n5153 VPWR.n5152 0.120292
R9700 VPWR.n5152 VPWR.n5148 0.120292
R9701 VPWR.n5148 VPWR.n5144 0.120292
R9702 VPWR.n5144 VPWR.n5143 0.120292
R9703 VPWR.n5138 VPWR.n5130 0.120292
R9704 VPWR.n5130 VPWR.n5129 0.120292
R9705 VPWR.n5129 VPWR.n5128 0.120292
R9706 VPWR.n5128 VPWR.n5126 0.120292
R9707 VPWR.n5122 VPWR.n5121 0.120292
R9708 VPWR.n5111 VPWR.n5110 0.120292
R9709 VPWR.n5110 VPWR.n5108 0.120292
R9710 VPWR.n5108 VPWR.n5102 0.120292
R9711 VPWR.n5099 VPWR.n5098 0.120292
R9712 VPWR.n5098 VPWR.n5096 0.120292
R9713 VPWR.n5029 VPWR.n5026 0.120292
R9714 VPWR.n5026 VPWR.n5024 0.120292
R9715 VPWR.n1920 VPWR.n1917 0.120292
R9716 VPWR.n1922 VPWR.n1920 0.120292
R9717 VPWR.n1925 VPWR.n1922 0.120292
R9718 VPWR.n1926 VPWR.n1925 0.120292
R9719 VPWR.n1927 VPWR.n1926 0.120292
R9720 VPWR.n1937 VPWR.n1933 0.120292
R9721 VPWR.n1941 VPWR.n1937 0.120292
R9722 VPWR.n1944 VPWR.n1941 0.120292
R9723 VPWR.n1946 VPWR.n1944 0.120292
R9724 VPWR.n1948 VPWR.n1946 0.120292
R9725 VPWR.n1955 VPWR.n1954 0.120292
R9726 VPWR.n1956 VPWR.n1955 0.120292
R9727 VPWR.n1957 VPWR.n1956 0.120292
R9728 VPWR.n5011 VPWR.n1960 0.120292
R9729 VPWR.n5009 VPWR.n5008 0.120292
R9730 VPWR.n4966 VPWR.n4965 0.120292
R9731 VPWR.n4965 VPWR.n4961 0.120292
R9732 VPWR.n4961 VPWR.n4959 0.120292
R9733 VPWR.n4959 VPWR.n4957 0.120292
R9734 VPWR.n4954 VPWR.n4953 0.120292
R9735 VPWR.n4953 VPWR.n4949 0.120292
R9736 VPWR.n4949 VPWR.n4945 0.120292
R9737 VPWR.n4945 VPWR.n4942 0.120292
R9738 VPWR.n4942 VPWR.n4940 0.120292
R9739 VPWR.n4940 VPWR.n4938 0.120292
R9740 VPWR.n4934 VPWR.n4933 0.120292
R9741 VPWR.n4933 VPWR.n4932 0.120292
R9742 VPWR.n4932 VPWR.n4931 0.120292
R9743 VPWR.n2227 VPWR.n2224 0.120292
R9744 VPWR.n2228 VPWR.n2227 0.120292
R9745 VPWR.n2237 VPWR.n2232 0.120292
R9746 VPWR.n2238 VPWR.n2237 0.120292
R9747 VPWR.n2246 VPWR.n2242 0.120292
R9748 VPWR.n2250 VPWR.n2246 0.120292
R9749 VPWR.n2252 VPWR.n2250 0.120292
R9750 VPWR.n2254 VPWR.n2252 0.120292
R9751 VPWR.n2256 VPWR.n2255 0.120292
R9752 VPWR.n2265 VPWR.n2261 0.120292
R9753 VPWR.n2267 VPWR.n2265 0.120292
R9754 VPWR.n2269 VPWR.n2267 0.120292
R9755 VPWR.n2377 VPWR.n2294 0.120292
R9756 VPWR.n2300 VPWR.n2294 0.120292
R9757 VPWR.n2369 VPWR.n2366 0.120292
R9758 VPWR.n2363 VPWR.n2362 0.120292
R9759 VPWR.n2362 VPWR.n2360 0.120292
R9760 VPWR.n2360 VPWR.n2358 0.120292
R9761 VPWR.n2358 VPWR.n2356 0.120292
R9762 VPWR.n2356 VPWR.n2352 0.120292
R9763 VPWR.n2352 VPWR.n2350 0.120292
R9764 VPWR.n2350 VPWR.n2346 0.120292
R9765 VPWR.n2346 VPWR.n2344 0.120292
R9766 VPWR.n2344 VPWR.n2342 0.120292
R9767 VPWR.n2342 VPWR.n2340 0.120292
R9768 VPWR.n2340 VPWR.n2338 0.120292
R9769 VPWR.n2334 VPWR.n2333 0.120292
R9770 VPWR.n2333 VPWR.n2332 0.120292
R9771 VPWR.n2332 VPWR.n2331 0.120292
R9772 VPWR.n2330 VPWR.n2329 0.120292
R9773 VPWR.n2329 VPWR.n2328 0.120292
R9774 VPWR.n2325 VPWR.n2324 0.120292
R9775 VPWR.n2687 VPWR.n2686 0.120292
R9776 VPWR.n2686 VPWR.n2685 0.120292
R9777 VPWR.n2101 VPWR.n2099 0.120292
R9778 VPWR.n2099 VPWR.n2095 0.120292
R9779 VPWR.n2095 VPWR.n2093 0.120292
R9780 VPWR.n2093 VPWR.n2087 0.120292
R9781 VPWR.n2087 VPWR.n2085 0.120292
R9782 VPWR.n2085 VPWR.n2082 0.120292
R9783 VPWR.n2082 VPWR.n2080 0.120292
R9784 VPWR.n2080 VPWR.n2076 0.120292
R9785 VPWR.n2076 VPWR.n2071 0.120292
R9786 VPWR.n2071 VPWR.n2069 0.120292
R9787 VPWR.n2069 VPWR.n2065 0.120292
R9788 VPWR.n2065 VPWR.n2061 0.120292
R9789 VPWR.n2060 VPWR.n2052 0.120292
R9790 VPWR.n2052 VPWR.n2051 0.120292
R9791 VPWR.n2051 VPWR.n2050 0.120292
R9792 VPWR.n2704 VPWR.n2702 0.120292
R9793 VPWR.n2706 VPWR.n2704 0.120292
R9794 VPWR.n2710 VPWR.n2706 0.120292
R9795 VPWR.n2713 VPWR.n2710 0.120292
R9796 VPWR.n2715 VPWR.n2713 0.120292
R9797 VPWR.n2716 VPWR.n2715 0.120292
R9798 VPWR.n2722 VPWR.n2721 0.120292
R9799 VPWR.n2723 VPWR.n2722 0.120292
R9800 VPWR.n2724 VPWR.n2723 0.120292
R9801 VPWR.n2732 VPWR.n2730 0.120292
R9802 VPWR.n4409 VPWR.n4405 0.120292
R9803 VPWR.n4420 VPWR.n4419 0.120292
R9804 VPWR.n4423 VPWR.n4420 0.120292
R9805 VPWR.n4425 VPWR.n4423 0.120292
R9806 VPWR.n4438 VPWR.n4437 0.120292
R9807 VPWR.n4439 VPWR.n4438 0.120292
R9808 VPWR.n4443 VPWR.n4439 0.120292
R9809 VPWR.n4445 VPWR.n4443 0.120292
R9810 VPWR.n4448 VPWR.n4445 0.120292
R9811 VPWR.n4449 VPWR.n4448 0.120292
R9812 VPWR.n4457 VPWR.n4455 0.120292
R9813 VPWR.n4461 VPWR.n4457 0.120292
R9814 VPWR.n4462 VPWR.n4461 0.120292
R9815 VPWR.n4470 VPWR.n4468 0.120292
R9816 VPWR.n4472 VPWR.n4470 0.120292
R9817 VPWR.n4473 VPWR.n4472 0.120292
R9818 VPWR.n4474 VPWR.n4473 0.120292
R9819 VPWR.n4475 VPWR.n4474 0.120292
R9820 VPWR.n4482 VPWR.n4480 0.120292
R9821 VPWR.n4534 VPWR.n4527 0.120292
R9822 VPWR.n4527 VPWR.n4526 0.120292
R9823 VPWR.n4526 VPWR.n4525 0.120292
R9824 VPWR.n4525 VPWR.n4523 0.120292
R9825 VPWR.n4523 VPWR.n4520 0.120292
R9826 VPWR.n4516 VPWR.n4515 0.120292
R9827 VPWR.n4511 VPWR.n4510 0.120292
R9828 VPWR.n4507 VPWR.n4506 0.120292
R9829 VPWR.n4506 VPWR.n4505 0.120292
R9830 VPWR.n3393 VPWR.n3388 0.120292
R9831 VPWR.n3394 VPWR.n3393 0.120292
R9832 VPWR.n3399 VPWR.n3398 0.120292
R9833 VPWR.n3400 VPWR.n3399 0.120292
R9834 VPWR.n3408 VPWR.n3400 0.120292
R9835 VPWR.n3424 VPWR.n3421 0.120292
R9836 VPWR.n3742 VPWR.n3739 0.120292
R9837 VPWR.n3734 VPWR.n3733 0.120292
R9838 VPWR.n3728 VPWR.n3723 0.120292
R9839 VPWR.n3723 VPWR.n3722 0.120292
R9840 VPWR.n3722 VPWR.n3721 0.120292
R9841 VPWR.n3718 VPWR.n3717 0.120292
R9842 VPWR.n3717 VPWR.n3715 0.120292
R9843 VPWR.n3715 VPWR.n3711 0.120292
R9844 VPWR.n3711 VPWR.n3709 0.120292
R9845 VPWR.n3709 VPWR.n3706 0.120292
R9846 VPWR.n3706 VPWR.n3704 0.120292
R9847 VPWR.n3704 VPWR.n3702 0.120292
R9848 VPWR.n3702 VPWR.n3699 0.120292
R9849 VPWR.n3699 VPWR.n3697 0.120292
R9850 VPWR.n3697 VPWR.n3695 0.120292
R9851 VPWR.n3695 VPWR.n3693 0.120292
R9852 VPWR.n3688 VPWR.n3687 0.120292
R9853 VPWR.n3687 VPWR.n3685 0.120292
R9854 VPWR.n3685 VPWR.n3684 0.120292
R9855 VPWR.n3684 VPWR.n3682 0.120292
R9856 VPWR.n3682 VPWR.n3677 0.120292
R9857 VPWR.n3540 VPWR.n3538 0.120292
R9858 VPWR.n3577 VPWR.n3576 0.120292
R9859 VPWR.n3587 VPWR.n3586 0.120292
R9860 VPWR.n3588 VPWR.n3587 0.120292
R9861 VPWR.n3590 VPWR.n3588 0.120292
R9862 VPWR.n3592 VPWR.n3590 0.120292
R9863 VPWR.n3593 VPWR.n3592 0.120292
R9864 VPWR.n3600 VPWR.n3597 0.120292
R9865 VPWR.n3602 VPWR.n3600 0.120292
R9866 VPWR.n3604 VPWR.n3602 0.120292
R9867 VPWR.n3609 VPWR.n3604 0.120292
R9868 VPWR.n3610 VPWR.n3609 0.120292
R9869 VPWR.n3617 VPWR.n3615 0.120292
R9870 VPWR.n3619 VPWR.n3617 0.120292
R9871 VPWR.n3622 VPWR.n3619 0.120292
R9872 VPWR.n3623 VPWR.n3622 0.120292
R9873 VPWR.n3667 VPWR.n3666 0.120292
R9874 VPWR.n3666 VPWR.n3665 0.120292
R9875 VPWR.n3665 VPWR.n3664 0.120292
R9876 VPWR.n3661 VPWR.n3660 0.120292
R9877 VPWR.n3660 VPWR.n3658 0.120292
R9878 VPWR.n3658 VPWR.n3656 0.120292
R9879 VPWR.n3656 VPWR.n3652 0.120292
R9880 VPWR.n3652 VPWR.n3649 0.120292
R9881 VPWR.n3649 VPWR.n3646 0.120292
R9882 VPWR.n3646 VPWR.n3644 0.120292
R9883 VPWR.n3641 VPWR.n3640 0.120292
R9884 VPWR.n4261 VPWR.n4259 0.120292
R9885 VPWR.n4259 VPWR.n4257 0.120292
R9886 VPWR.n4257 VPWR.n4255 0.120292
R9887 VPWR.n4255 VPWR.n4252 0.120292
R9888 VPWR.n2798 VPWR.n2797 0.120292
R9889 VPWR.n2804 VPWR.n2802 0.120292
R9890 VPWR.n2807 VPWR.n2804 0.120292
R9891 VPWR.n2809 VPWR.n2807 0.120292
R9892 VPWR.n2812 VPWR.n2809 0.120292
R9893 VPWR.n2816 VPWR.n2812 0.120292
R9894 VPWR.n2820 VPWR.n2816 0.120292
R9895 VPWR.n2823 VPWR.n2821 0.120292
R9896 VPWR.n2824 VPWR.n2823 0.120292
R9897 VPWR.n2825 VPWR.n2824 0.120292
R9898 VPWR.n2830 VPWR.n2825 0.120292
R9899 VPWR.n2839 VPWR.n2836 0.120292
R9900 VPWR.n2841 VPWR.n2839 0.120292
R9901 VPWR.n2845 VPWR.n2841 0.120292
R9902 VPWR.n2848 VPWR.n2845 0.120292
R9903 VPWR.n2850 VPWR.n2848 0.120292
R9904 VPWR.n2852 VPWR.n2850 0.120292
R9905 VPWR.n2855 VPWR.n2852 0.120292
R9906 VPWR.n2857 VPWR.n2855 0.120292
R9907 VPWR.n2861 VPWR.n2857 0.120292
R9908 VPWR.n2863 VPWR.n2861 0.120292
R9909 VPWR.n2864 VPWR.n2863 0.120292
R9910 VPWR.n4244 VPWR.n4240 0.120292
R9911 VPWR.n4240 VPWR.n4238 0.120292
R9912 VPWR.n4238 VPWR.n4236 0.120292
R9913 VPWR.n2935 VPWR.n2929 0.120292
R9914 VPWR.n2929 VPWR.n2927 0.120292
R9915 VPWR.n2927 VPWR.n2925 0.120292
R9916 VPWR.n2925 VPWR.n2923 0.120292
R9917 VPWR.n2920 VPWR.n2919 0.120292
R9918 VPWR.n2919 VPWR.n2918 0.120292
R9919 VPWR.n2918 VPWR.n2916 0.120292
R9920 VPWR.n2916 VPWR.n2914 0.120292
R9921 VPWR.n2914 VPWR.n2911 0.120292
R9922 VPWR.n2911 VPWR.n2909 0.120292
R9923 VPWR.n2909 VPWR.n2907 0.120292
R9924 VPWR.n2907 VPWR.n2905 0.120292
R9925 VPWR.n2905 VPWR.n2903 0.120292
R9926 VPWR.n2903 VPWR.n2901 0.120292
R9927 VPWR.n2901 VPWR.n2899 0.120292
R9928 VPWR.n7661 VPWR.n7657 0.120292
R9929 VPWR.n7662 VPWR.n7661 0.120292
R9930 VPWR.n7669 VPWR.n7668 0.120292
R9931 VPWR.n7674 VPWR.n7672 0.120292
R9932 VPWR.n7686 VPWR.n7681 0.120292
R9933 VPWR.n7741 VPWR.n7739 0.120292
R9934 VPWR.n7743 VPWR.n7741 0.120292
R9935 VPWR.n7746 VPWR.n7743 0.120292
R9936 VPWR.n7748 VPWR.n7746 0.120292
R9937 VPWR.n7750 VPWR.n7748 0.120292
R9938 VPWR.n7753 VPWR.n7750 0.120292
R9939 VPWR.n7770 VPWR.n7769 0.120292
R9940 VPWR.n7772 VPWR.n7770 0.120292
R9941 VPWR.n7774 VPWR.n7772 0.120292
R9942 VPWR.n7777 VPWR.n7774 0.120292
R9943 VPWR.n7779 VPWR.n7777 0.120292
R9944 VPWR.n7780 VPWR.n7779 0.120292
R9945 VPWR.n7781 VPWR.n7780 0.120292
R9946 VPWR.n7787 VPWR.n7785 0.120292
R9947 VPWR.n7788 VPWR.n7787 0.120292
R9948 VPWR.n7789 VPWR.n7788 0.120292
R9949 VPWR.n7796 VPWR.n7794 0.120292
R9950 VPWR.n7798 VPWR.n7796 0.120292
R9951 VPWR.n7800 VPWR.n7798 0.120292
R9952 VPWR.n7803 VPWR.n7800 0.120292
R9953 VPWR.n7805 VPWR.n7803 0.120292
R9954 VPWR.n7806 VPWR.n7805 0.120292
R9955 VPWR.n7807 VPWR.n7806 0.120292
R9956 VPWR.n7813 VPWR.n7812 0.120292
R9957 VPWR.n7814 VPWR.n7813 0.120292
R9958 VPWR.n6021 VPWR.n6007 0.120292
R9959 VPWR.n6023 VPWR.n6021 0.120292
R9960 VPWR.n6025 VPWR.n6023 0.120292
R9961 VPWR.n6026 VPWR.n6025 0.120292
R9962 VPWR.n6032 VPWR.n6031 0.120292
R9963 VPWR.n6033 VPWR.n6032 0.120292
R9964 VPWR.n6040 VPWR.n6037 0.120292
R9965 VPWR.n6041 VPWR.n6040 0.120292
R9966 VPWR.n6048 VPWR.n6046 0.120292
R9967 VPWR.n6049 VPWR.n6048 0.120292
R9968 VPWR.n6053 VPWR.n6052 0.120292
R9969 VPWR.n6105 VPWR.n6102 0.120292
R9970 VPWR.n6102 VPWR.n6100 0.120292
R9971 VPWR.n6100 VPWR.n6097 0.120292
R9972 VPWR.n6097 VPWR.n6094 0.120292
R9973 VPWR.n6094 VPWR.n6092 0.120292
R9974 VPWR.n6092 VPWR.n6091 0.120292
R9975 VPWR.n6091 VPWR.n6090 0.120292
R9976 VPWR.n6087 VPWR.n6086 0.120292
R9977 VPWR.n6086 VPWR.n6084 0.120292
R9978 VPWR.n6079 VPWR.n6078 0.120292
R9979 VPWR.n6078 VPWR.n6077 0.120292
R9980 VPWR.n9197 VPWR.n33 0.120292
R9981 VPWR.n9191 VPWR.n9190 0.120292
R9982 VPWR.n9190 VPWR.n9188 0.120292
R9983 VPWR.n9184 VPWR.n9183 0.120292
R9984 VPWR.n9183 VPWR.n9182 0.120292
R9985 VPWR.n9182 VPWR.n9181 0.120292
R9986 VPWR.n9177 VPWR.n9176 0.120292
R9987 VPWR.n9176 VPWR.n9171 0.120292
R9988 VPWR.n9166 VPWR.n9165 0.120292
R9989 VPWR.n9165 VPWR.n9164 0.120292
R9990 VPWR.n9164 VPWR.n9163 0.120292
R9991 VPWR.n9160 VPWR.n9159 0.120292
R9992 VPWR.n9159 VPWR.n9158 0.120292
R9993 VPWR.n9153 VPWR.n9150 0.120292
R9994 VPWR.n9150 VPWR.n9148 0.120292
R9995 VPWR.n9148 VPWR.n9147 0.120292
R9996 VPWR.n9147 VPWR.n9146 0.120292
R9997 VPWR.n9142 VPWR.n9141 0.120292
R9998 VPWR.n113 VPWR.n108 0.120292
R9999 VPWR.n105 VPWR.n104 0.120292
R10000 VPWR.n104 VPWR.n99 0.120292
R10001 VPWR.n99 VPWR.n97 0.120292
R10002 VPWR.n90 VPWR.n88 0.120292
R10003 VPWR.n84 VPWR.n82 0.120292
R10004 VPWR.n3254 VPWR.n3253 0.120292
R10005 VPWR.n3255 VPWR.n3254 0.120292
R10006 VPWR.n3256 VPWR.n3255 0.120292
R10007 VPWR.n3262 VPWR.n3259 0.120292
R10008 VPWR.n3270 VPWR.n3267 0.120292
R10009 VPWR.n3274 VPWR.n3270 0.120292
R10010 VPWR.n3281 VPWR.n3274 0.120292
R10011 VPWR.n3283 VPWR.n3282 0.120292
R10012 VPWR.n3284 VPWR.n3283 0.120292
R10013 VPWR.n3291 VPWR.n3289 0.120292
R10014 VPWR.n3232 VPWR.n3230 0.120292
R10015 VPWR.n3230 VPWR.n3228 0.120292
R10016 VPWR.n3228 VPWR.n3225 0.120292
R10017 VPWR.n3225 VPWR.n3223 0.120292
R10018 VPWR.n3223 VPWR.n3221 0.120292
R10019 VPWR.n3221 VPWR.n3217 0.120292
R10020 VPWR.n3210 VPWR.n3207 0.120292
R10021 VPWR.n3204 VPWR.n3203 0.120292
R10022 VPWR.n3199 VPWR.n3198 0.120292
R10023 VPWR.n3198 VPWR.n3197 0.120292
R10024 VPWR.n3197 VPWR.n3195 0.120292
R10025 VPWR.n3195 VPWR.n3193 0.120292
R10026 VPWR.n3193 VPWR.n3190 0.120292
R10027 VPWR.n3190 VPWR.n3188 0.120292
R10028 VPWR.n3188 VPWR.n3186 0.120292
R10029 VPWR.n3183 VPWR.n3182 0.120292
R10030 VPWR.n3182 VPWR.n3180 0.120292
R10031 VPWR.n3180 VPWR.n3176 0.120292
R10032 VPWR.n3172 VPWR.n3171 0.120292
R10033 VPWR.n3167 VPWR.n3166 0.120292
R10034 VPWR.n3166 VPWR.n3164 0.120292
R10035 VPWR.n3163 VPWR.n3162 0.120292
R10036 VPWR.n3086 VPWR.n3085 0.120292
R10037 VPWR.n3085 VPWR.n3084 0.120292
R10038 VPWR.n3084 VPWR.n3083 0.120292
R10039 VPWR.n3083 VPWR.n3081 0.120292
R10040 VPWR.n3077 VPWR.n3076 0.120292
R10041 VPWR.n3076 VPWR.n3075 0.120292
R10042 VPWR.n3891 VPWR.n3889 0.120292
R10043 VPWR.n3895 VPWR.n3891 0.120292
R10044 VPWR.n3898 VPWR.n3895 0.120292
R10045 VPWR.n3902 VPWR.n3898 0.120292
R10046 VPWR.n3905 VPWR.n3902 0.120292
R10047 VPWR.n3920 VPWR.n3914 0.120292
R10048 VPWR.n3922 VPWR.n3920 0.120292
R10049 VPWR.n3994 VPWR.n3990 0.120292
R10050 VPWR.n3996 VPWR.n3994 0.120292
R10051 VPWR.n4000 VPWR.n3996 0.120292
R10052 VPWR.n4003 VPWR.n4000 0.120292
R10053 VPWR.n4019 VPWR.n4018 0.120292
R10054 VPWR.n4020 VPWR.n4019 0.120292
R10055 VPWR.n4021 VPWR.n4020 0.120292
R10056 VPWR.n4023 VPWR.n4021 0.120292
R10057 VPWR.n4026 VPWR.n4023 0.120292
R10058 VPWR.n4035 VPWR.n4034 0.120292
R10059 VPWR.n4037 VPWR.n4035 0.120292
R10060 VPWR.n4039 VPWR.n4037 0.120292
R10061 VPWR.n4042 VPWR.n4039 0.120292
R10062 VPWR.n4044 VPWR.n4042 0.120292
R10063 VPWR.n4046 VPWR.n4044 0.120292
R10064 VPWR.n4048 VPWR.n4046 0.120292
R10065 VPWR.n4050 VPWR.n4048 0.120292
R10066 VPWR.n4051 VPWR.n4050 0.120292
R10067 VPWR.n4057 VPWR.n4056 0.120292
R10068 VPWR.n4070 VPWR.n4066 0.120292
R10069 VPWR.n4079 VPWR.n4077 0.120292
R10070 VPWR.n4081 VPWR.n4079 0.120292
R10071 VPWR.n4085 VPWR.n4081 0.120292
R10072 VPWR.n4135 VPWR.n4133 0.120292
R10073 VPWR.n4133 VPWR.n4131 0.120292
R10074 VPWR.n4131 VPWR.n4129 0.120292
R10075 VPWR.n4123 VPWR.n4121 0.120292
R10076 VPWR.n4109 VPWR.n4092 0.120292
R10077 VPWR.n4099 VPWR.n4092 0.120292
R10078 VPWR.n7533 VPWR.n7532 0.120292
R10079 VPWR.n7538 VPWR.n7536 0.120292
R10080 VPWR.n7541 VPWR.n7538 0.120292
R10081 VPWR.n7543 VPWR.n7541 0.120292
R10082 VPWR.n7546 VPWR.n7543 0.120292
R10083 VPWR.n7547 VPWR.n7546 0.120292
R10084 VPWR.n7551 VPWR.n7550 0.120292
R10085 VPWR.n7556 VPWR.n7554 0.120292
R10086 VPWR.n7559 VPWR.n7556 0.120292
R10087 VPWR.n7565 VPWR.n7559 0.120292
R10088 VPWR.n7567 VPWR.n7566 0.120292
R10089 VPWR.n7568 VPWR.n7567 0.120292
R10090 VPWR.n7574 VPWR.n7572 0.120292
R10091 VPWR.n7526 VPWR.n7525 0.120292
R10092 VPWR.n7525 VPWR.n7523 0.120292
R10093 VPWR.n7523 VPWR.n7521 0.120292
R10094 VPWR.n7521 VPWR.n7519 0.120292
R10095 VPWR.n7519 VPWR.n7517 0.120292
R10096 VPWR.n7517 VPWR.n7515 0.120292
R10097 VPWR.n7511 VPWR.n7510 0.120292
R10098 VPWR.n7510 VPWR.n7508 0.120292
R10099 VPWR.n7508 VPWR.n7507 0.120292
R10100 VPWR.n7503 VPWR.n7502 0.120292
R10101 VPWR.n7502 VPWR.n7501 0.120292
R10102 VPWR.n7501 VPWR.n7500 0.120292
R10103 VPWR.n7497 VPWR.n7496 0.120292
R10104 VPWR.n7496 VPWR.n7494 0.120292
R10105 VPWR.n7494 VPWR.n7492 0.120292
R10106 VPWR.n7492 VPWR.n7490 0.120292
R10107 VPWR.n7490 VPWR.n7487 0.120292
R10108 VPWR.n7487 VPWR.n7485 0.120292
R10109 VPWR.n7485 VPWR.n7483 0.120292
R10110 VPWR.n7483 VPWR.n7481 0.120292
R10111 VPWR.n7481 VPWR.n7479 0.120292
R10112 VPWR.n7479 VPWR.n7477 0.120292
R10113 VPWR.n7477 VPWR.n7475 0.120292
R10114 VPWR.n7468 VPWR.n7467 0.120292
R10115 VPWR.n7467 VPWR.n7465 0.120292
R10116 VPWR.n7464 VPWR.n7462 0.120292
R10117 VPWR.n7458 VPWR.n7457 0.120292
R10118 VPWR.n7414 VPWR.n7413 0.120292
R10119 VPWR.n7413 VPWR.n7411 0.120292
R10120 VPWR.n7411 VPWR.n7409 0.120292
R10121 VPWR.n7409 VPWR.n7407 0.120292
R10122 VPWR.n7407 VPWR.n7405 0.120292
R10123 VPWR.n7405 VPWR.n7403 0.120292
R10124 VPWR.n7399 VPWR.n7398 0.120292
R10125 VPWR.n7398 VPWR.n7396 0.120292
R10126 VPWR.n7392 VPWR.n7391 0.120292
R10127 VPWR.n7391 VPWR.n7390 0.120292
R10128 VPWR.n7390 VPWR.n7389 0.120292
R10129 VPWR.n7389 VPWR.n7387 0.120292
R10130 VPWR.n7387 VPWR.n7385 0.120292
R10131 VPWR.n7385 VPWR.n7383 0.120292
R10132 VPWR.n7383 VPWR 0.120292
R10133 VPWR.n7377 VPWR.n7376 0.120292
R10134 VPWR.n7376 VPWR.n7375 0.120292
R10135 VPWR.n7375 VPWR.n7374 0.120292
R10136 VPWR.n7371 VPWR.n7370 0.120292
R10137 VPWR.n7370 VPWR.n7368 0.120292
R10138 VPWR.n7368 VPWR.n7367 0.120292
R10139 VPWR.n7367 VPWR.n7365 0.120292
R10140 VPWR.n7365 VPWR.n7364 0.120292
R10141 VPWR.n7360 VPWR.n7359 0.120292
R10142 VPWR.n7359 VPWR.n7358 0.120292
R10143 VPWR.n7358 VPWR.n7357 0.120292
R10144 VPWR.n7354 VPWR.n7353 0.120292
R10145 VPWR.n7353 VPWR.n7352 0.120292
R10146 VPWR.n7060 VPWR.n7057 0.120292
R10147 VPWR.n7062 VPWR.n7060 0.120292
R10148 VPWR.n7065 VPWR.n7062 0.120292
R10149 VPWR.n7067 VPWR.n7065 0.120292
R10150 VPWR.n7077 VPWR.n7076 0.120292
R10151 VPWR.n7078 VPWR.n7077 0.120292
R10152 VPWR.n7079 VPWR.n7078 0.120292
R10153 VPWR.n7085 VPWR.n7083 0.120292
R10154 VPWR.n7087 VPWR.n7085 0.120292
R10155 VPWR.n7089 VPWR.n7087 0.120292
R10156 VPWR.n7092 VPWR.n7089 0.120292
R10157 VPWR.n7094 VPWR.n7092 0.120292
R10158 VPWR.n7096 VPWR.n7094 0.120292
R10159 VPWR.n7098 VPWR.n7096 0.120292
R10160 VPWR.n7100 VPWR.n7098 0.120292
R10161 VPWR.n7102 VPWR.n7100 0.120292
R10162 VPWR.n7104 VPWR.n7102 0.120292
R10163 VPWR.n7105 VPWR.n7104 0.120292
R10164 VPWR.n7110 VPWR.n7108 0.120292
R10165 VPWR.n7111 VPWR.n7110 0.120292
R10166 VPWR.n7118 VPWR.n7116 0.120292
R10167 VPWR.n7125 VPWR.n7118 0.120292
R10168 VPWR.n7127 VPWR.n7126 0.120292
R10169 VPWR.n7128 VPWR.n7127 0.120292
R10170 VPWR.n7276 VPWR.n7275 0.120292
R10171 VPWR.n7275 VPWR.n7272 0.120292
R10172 VPWR.n7272 VPWR.n7267 0.120292
R10173 VPWR.n7267 VPWR.n7264 0.120292
R10174 VPWR.n7189 VPWR.n7188 0.120292
R10175 VPWR.n7188 VPWR.n7186 0.120292
R10176 VPWR.n7181 VPWR.n7180 0.120292
R10177 VPWR.n7180 VPWR.n7178 0.120292
R10178 VPWR.n7178 VPWR.n7177 0.120292
R10179 VPWR.n7177 VPWR.n7175 0.120292
R10180 VPWR.n7170 VPWR.n7169 0.120292
R10181 VPWR.n7169 VPWR.n7167 0.120292
R10182 VPWR.n7167 VPWR.n7166 0.120292
R10183 VPWR.n7166 VPWR.n7164 0.120292
R10184 VPWR.n7163 VPWR.n7162 0.120292
R10185 VPWR.n7162 VPWR.n7161 0.120292
R10186 VPWR VPWR.n8973 0.12003
R10187 VPWR.n8973 VPWR 0.12003
R10188 VPWR VPWR.n5873 0.12003
R10189 VPWR.n5873 VPWR 0.12003
R10190 VPWR VPWR.n4714 0.12003
R10191 VPWR VPWR.n9129 0.12003
R10192 VPWR VPWR.n3211 0.12003
R10193 VPWR.n1333 VPWR.n1326 0.116104
R10194 VPWR.n3936 VPWR.n3935 0.113774
R10195 VPWR.n4839 VPWR.n4838 0.113774
R10196 VPWR.n2931 VPWR.n2930 0.113774
R10197 VPWR.n8059 VPWR.n8058 0.109682
R10198 VPWR.n8255 VPWR.n8254 0.109682
R10199 VPWR.n8574 VPWR.n8514 0.109682
R10200 VPWR.n1092 VPWR.n1038 0.109682
R10201 VPWR.n5515 VPWR.n5496 0.109682
R10202 VPWR.n5256 VPWR.n5254 0.109682
R10203 VPWR.n5085 VPWR.n5084 0.109682
R10204 VPWR.n4359 VPWR.n2732 0.109682
R10205 VPWR.n4301 VPWR.n2784 0.109682
R10206 VPWR.n3934 VPWR.n3922 0.109682
R10207 VPWR.n2636 VPWR.n2101 0.109342
R10208 VPWR.n3576 VPWR.n3573 0.109342
R10209 VPWR.n7855 VPWR.n6007 0.109342
R10210 VPWR.n7415 VPWR.n7414 0.109342
R10211 VPWR.n8343 VPWR.n8342 0.108642
R10212 VPWR.n5404 VPWR.n5400 0.108642
R10213 VPWR.n5323 VPWR.n5322 0.108642
R10214 VPWR.n5160 VPWR.n5159 0.108642
R10215 VPWR.n3829 VPWR.n3090 0.108642
R10216 VPWR.n6442 VPWR.n6439 0.107271
R10217 VPWR.n872 VPWR.n871 0.107271
R10218 VPWR.n1430 VPWR.n1426 0.107271
R10219 VPWR.n1770 VPWR.n1769 0.107271
R10220 VPWR.n2685 VPWR.n2680 0.107271
R10221 VPWR.n3542 VPWR.n3540 0.107271
R10222 VPWR.n7454 VPWR.n7453 0.107271
R10223 VPWR.n7590 VPWR.n7589 0.106285
R10224 VPWR.n3309 VPWR.n3308 0.106285
R10225 VPWR.n9039 VPWR.n9038 0.106285
R10226 VPWR.n1500 VPWR.n1372 0.106285
R10227 VPWR.n1320 VPWR.n1319 0.106285
R10228 VPWR.n1348 VPWR.n1347 0.106285
R10229 VPWR.n4808 VPWR.n4807 0.106285
R10230 VPWR.n4402 VPWR.n4401 0.106285
R10231 VPWR.n9066 VPWR.n9065 0.105969
R10232 VPWR.n8200 VPWR.n8199 0.105969
R10233 VPWR.n5580 VPWR.n5577 0.105969
R10234 VPWR.n4676 VPWR.n4674 0.105969
R10235 VPWR.n4405 VPWR.n4403 0.105969
R10236 VPWR.n4265 VPWR.n4261 0.105969
R10237 VPWR.n3990 VPWR.n3988 0.105969
R10238 VPWR.n7057 VPWR.n7055 0.105969
R10239 VPWR.n787 VPWR.n786 0.105956
R10240 VPWR.n5856 VPWR.n362 0.105956
R10241 VPWR.n676 VPWR.n675 0.105956
R10242 VPWR.n5853 VPWR.n5852 0.105956
R10243 VPWR.n6171 VPWR 0.104136
R10244 VPWR.n6596 VPWR 0.104136
R10245 VPWR.n6495 VPWR 0.104136
R10246 VPWR.n610 VPWR 0.104136
R10247 VPWR.n1286 VPWR 0.104136
R10248 VPWR.n1549 VPWR 0.104136
R10249 VPWR.n2441 VPWR 0.104136
R10250 VPWR.n2218 VPWR 0.104136
R10251 VPWR.n3381 VPWR 0.104136
R10252 VPWR.n7649 VPWR 0.104136
R10253 VPWR.n3245 VPWR 0.104136
R10254 VPWR.n3079 VPWR.n3078 0.102087
R10255 VPWR.n3240 VPWR.n3239 0.102087
R10256 VPWR.n128 VPWR.n127 0.102087
R10257 VPWR.n9195 VPWR.n9194 0.102087
R10258 VPWR.n6070 VPWR.n6069 0.102087
R10259 VPWR.n275 VPWR.n274 0.102087
R10260 VPWR.n7994 VPWR.n7993 0.102087
R10261 VPWR.n8852 VPWR.n8851 0.102087
R10262 VPWR.n8430 VPWR.n8429 0.102087
R10263 VPWR.n8572 VPWR.n8571 0.102087
R10264 VPWR.n6372 VPWR.n6371 0.102087
R10265 VPWR.n6510 VPWR.n6509 0.102087
R10266 VPWR.n6542 VPWR.n6541 0.102087
R10267 VPWR.n887 VPWR.n886 0.102087
R10268 VPWR.n1297 VPWR.n1296 0.102087
R10269 VPWR.n4916 VPWR.n4915 0.102087
R10270 VPWR.n2481 VPWR.n2480 0.102087
R10271 VPWR.n2049 VPWR.n2048 0.102087
R10272 VPWR.n1993 VPWR.n1992 0.102087
R10273 VPWR.n4546 VPWR.n4545 0.102087
R10274 VPWR.n7210 VPWR.n7209 0.102087
R10275 VPWR.n614 VPWR 0.0994583
R10276 VPWR.n5316 VPWR 0.0994583
R10277 VPWR.n6296 VPWR 0.0981562
R10278 VPWR VPWR.n6294 0.0981562
R10279 VPWR.n8010 VPWR 0.0981562
R10280 VPWR.n7920 VPWR 0.0981562
R10281 VPWR.n8988 VPWR 0.0981562
R10282 VPWR.n9021 VPWR 0.0981562
R10283 VPWR VPWR.n228 0.0981562
R10284 VPWR.n6603 VPWR 0.0981562
R10285 VPWR.n6619 VPWR 0.0981562
R10286 VPWR.n6764 VPWR 0.0981562
R10287 VPWR VPWR.n6761 0.0981562
R10288 VPWR.n6724 VPWR 0.0981562
R10289 VPWR.n6693 VPWR 0.0981562
R10290 VPWR.n8255 VPWR 0.0981562
R10291 VPWR.n8130 VPWR 0.0981562
R10292 VPWR.n8170 VPWR 0.0981562
R10293 VPWR.n8885 VPWR 0.0981562
R10294 VPWR.n6518 VPWR 0.0981562
R10295 VPWR.n6413 VPWR 0.0981562
R10296 VPWR VPWR.n5878 0.0981562
R10297 VPWR.n8434 VPWR 0.0981562
R10298 VPWR.n8489 VPWR 0.0981562
R10299 VPWR.n8494 VPWR 0.0981562
R10300 VPWR.n8600 VPWR 0.0981562
R10301 VPWR VPWR.n8760 0.0981562
R10302 VPWR.n623 VPWR 0.0981562
R10303 VPWR.n632 VPWR 0.0981562
R10304 VPWR.n845 VPWR 0.0981562
R10305 VPWR.n1134 VPWR 0.0981562
R10306 VPWR.n1139 VPWR 0.0981562
R10307 VPWR.n5825 VPWR 0.0981562
R10308 VPWR.n5796 VPWR 0.0981562
R10309 VPWR.n1322 VPWR 0.0981562
R10310 VPWR VPWR.n1516 0.0981562
R10311 VPWR.n1486 VPWR 0.0981562
R10312 VPWR.n1456 VPWR 0.0981562
R10313 VPWR.n5445 VPWR 0.0981562
R10314 VPWR.n5487 VPWR 0.0981562
R10315 VPWR.n5493 VPWR 0.0981562
R10316 VPWR.n5590 VPWR 0.0981562
R10317 VPWR.n5639 VPWR 0.0981562
R10318 VPWR.n5644 VPWR 0.0981562
R10319 VPWR.n442 VPWR 0.0981562
R10320 VPWR VPWR.n441 0.0981562
R10321 VPWR VPWR.n423 0.0981562
R10322 VPWR.n1705 VPWR 0.0981562
R10323 VPWR.n1713 VPWR 0.0981562
R10324 VPWR VPWR.n552 0.0981562
R10325 VPWR VPWR.n4747 0.0981562
R10326 VPWR VPWR.n4722 0.0981562
R10327 VPWR.n4826 VPWR 0.0981562
R10328 VPWR VPWR.n4815 0.0981562
R10329 VPWR.n2446 VPWR 0.0981562
R10330 VPWR.n2452 VPWR 0.0981562
R10331 VPWR VPWR.n2424 0.0981562
R10332 VPWR.n2560 VPWR 0.0981562
R10333 VPWR.n2151 VPWR 0.0981562
R10334 VPWR.n5030 VPWR 0.0981562
R10335 VPWR.n1917 VPWR 0.0981562
R10336 VPWR VPWR.n5009 0.0981562
R10337 VPWR.n2334 VPWR 0.0981562
R10338 VPWR VPWR.n2320 0.0981562
R10339 VPWR VPWR.n4516 0.0981562
R10340 VPWR VPWR.n4511 0.0981562
R10341 VPWR.n4507 VPWR 0.0981562
R10342 VPWR.n3414 VPWR 0.0981562
R10343 VPWR VPWR.n3742 0.0981562
R10344 VPWR VPWR.n3688 0.0981562
R10345 VPWR.n3615 VPWR 0.0981562
R10346 VPWR.n3671 VPWR 0.0981562
R10347 VPWR VPWR.n2784 0.0981562
R10348 VPWR.n2789 VPWR 0.0981562
R10349 VPWR.n2831 VPWR 0.0981562
R10350 VPWR.n4246 VPWR 0.0981562
R10351 VPWR.n7668 VPWR 0.0981562
R10352 VPWR.n7681 VPWR 0.0981562
R10353 VPWR.n7754 VPWR 0.0981562
R10354 VPWR.n7785 VPWR 0.0981562
R10355 VPWR.n7794 VPWR 0.0981562
R10356 VPWR.n7808 VPWR 0.0981562
R10357 VPWR.n6031 VPWR 0.0981562
R10358 VPWR.n6037 VPWR 0.0981562
R10359 VPWR.n6052 VPWR 0.0981562
R10360 VPWR VPWR.n85 0.0981562
R10361 VPWR.n3183 VPWR 0.0981562
R10362 VPWR.n3173 VPWR 0.0981562
R10363 VPWR.n3167 VPWR 0.0981562
R10364 VPWR VPWR.n3873 0.0981562
R10365 VPWR.n3077 VPWR 0.0981562
R10366 VPWR.n3914 VPWR 0.0981562
R10367 VPWR.n4056 VPWR 0.0981562
R10368 VPWR.n4058 VPWR 0.0981562
R10369 VPWR.n4062 VPWR 0.0981562
R10370 VPWR.n4125 VPWR 0.0981562
R10371 VPWR VPWR.n4124 0.0981562
R10372 VPWR VPWR.n4123 0.0981562
R10373 VPWR.n7532 VPWR 0.0981562
R10374 VPWR.n7512 VPWR 0.0981562
R10375 VPWR VPWR.n7472 0.0981562
R10376 VPWR.n7468 VPWR 0.0981562
R10377 VPWR.n7400 VPWR 0.0981562
R10378 VPWR VPWR.n7399 0.0981562
R10379 VPWR.n7108 VPWR 0.0981562
R10380 VPWR.n7116 VPWR 0.0981562
R10381 VPWR.n7189 VPWR 0.0981562
R10382 VPWR.n7181 VPWR 0.0981562
R10383 VPWR VPWR.n7170 0.0981562
R10384 VPWR VPWR.n8894 0.0968542
R10385 VPWR VPWR.n8770 0.0968542
R10386 VPWR.n1036 VPWR 0.0968542
R10387 VPWR.n5496 VPWR 0.0968542
R10388 VPWR.n5624 VPWR 0.0968542
R10389 VPWR VPWR.n1772 0.0968542
R10390 VPWR VPWR.n5280 0.0968542
R10391 VPWR VPWR.n4751 0.0968542
R10392 VPWR VPWR.n4821 0.0968542
R10393 VPWR VPWR.n5085 0.0968542
R10394 VPWR.n2730 VPWR 0.0968542
R10395 VPWR VPWR.n90 0.0968542
R10396 VPWR.n3774 VPWR.n3759 0.0942472
R10397 VPWR.n4319 VPWR.n2782 0.0942472
R10398 VPWR.n4210 VPWR.n2977 0.0940635
R10399 VPWR VPWR.n6187 0.0930549
R10400 VPWR.n4005 VPWR 0.0930549
R10401 VPWR.n9265 VPWR 0.0875462
R10402 VPWR.n8970 VPWR.n8965 0.0863232
R10403 VPWR.n8703 VPWR.n8692 0.0863232
R10404 VPWR.n4869 VPWR.n4784 0.0863232
R10405 VPWR.n4236 VPWR.n4231 0.0863232
R10406 VPWR.n4169 VPWR.n4085 0.0863232
R10407 VPWR.n7264 VPWR.n7262 0.0863232
R10408 VPWR.n7862 VPWR.n7861 0.0859812
R10409 VPWR.n9100 VPWR.n9099 0.0859812
R10410 VPWR.n6895 VPWR.n6894 0.0859812
R10411 VPWR.n9103 VPWR.n163 0.0859812
R10412 VPWR.n6869 VPWR.n6311 0.0857946
R10413 VPWR.n6791 VPWR.n6779 0.0857946
R10414 VPWR.n1644 VPWR.n1642 0.0857946
R10415 VPWR.n2547 VPWR.n2546 0.0857946
R10416 VPWR.n7739 VPWR.n7737 0.0857946
R10417 VPWR.n7609 VPWR.n7526 0.0857946
R10418 VPWR VPWR.n8008 0.0851354
R10419 VPWR.n7817 VPWR 0.0851354
R10420 VPWR.n3328 VPWR.n3232 0.0850212
R10421 VPWR.n3094 VPWR 0.0830437
R10422 VPWR.n3004 VPWR 0.0830437
R10423 VPWR.n3357 VPWR 0.0830437
R10424 VPWR.n2984 VPWR 0.0830437
R10425 VPWR.n6262 VPWR 0.0826382
R10426 VPWR.n6762 VPWR 0.0826382
R10427 VPWR.n6692 VPWR 0.0826382
R10428 VPWR.n4711 VPWR 0.0826382
R10429 VPWR.n3636 VPWR 0.0826382
R10430 VPWR VPWR.n7767 0.0826382
R10431 VPWR.n3907 VPWR 0.0826382
R10432 VPWR.n4027 VPWR 0.0826382
R10433 VPWR.n1908 VPWR 0.0822696
R10434 VPWR.n2045 VPWR 0.0822696
R10435 VPWR.n3211 VPWR 0.0822696
R10436 VPWR.n1950 VPWR 0.0813361
R10437 VPWR.n1931 VPWR.n1911 0.0800618
R10438 VPWR.n4855 VPWR.n4854 0.0760162
R10439 VPWR.n7861 VPWR.n7860 0.0660062
R10440 VPWR.n9100 VPWR.n165 0.0660062
R10441 VPWR.n6896 VPWR.n6895 0.0660062
R10442 VPWR.n9104 VPWR.n9103 0.0660062
R10443 VPWR.n7822 VPWR.n7821 0.0620385
R10444 VPWR.n6812 VPWR.n6811 0.0620385
R10445 VPWR.n6178 VPWR 0.0603958
R10446 VPWR.n6184 VPWR 0.0603958
R10447 VPWR.n6194 VPWR 0.0603958
R10448 VPWR.n6286 VPWR 0.0603958
R10449 VPWR.n6279 VPWR 0.0603958
R10450 VPWR VPWR.n6270 0.0603958
R10451 VPWR VPWR.n6260 0.0603958
R10452 VPWR VPWR.n7955 0.0603958
R10453 VPWR.n7951 VPWR 0.0603958
R10454 VPWR VPWR.n5965 0.0603958
R10455 VPWR.n8018 VPWR 0.0603958
R10456 VPWR.n8046 VPWR 0.0603958
R10457 VPWR.n8051 VPWR 0.0603958
R10458 VPWR.n194 VPWR 0.0603958
R10459 VPWR.n8980 VPWR 0.0603958
R10460 VPWR.n9031 VPWR 0.0603958
R10461 VPWR VPWR.n8974 0.0603958
R10462 VPWR VPWR.n8972 0.0603958
R10463 VPWR VPWR.n8971 0.0603958
R10464 VPWR.n241 VPWR 0.0603958
R10465 VPWR VPWR.n240 0.0603958
R10466 VPWR.n229 VPWR 0.0603958
R10467 VPWR VPWR.n227 0.0603958
R10468 VPWR.n6597 VPWR 0.0603958
R10469 VPWR.n6598 VPWR 0.0603958
R10470 VPWR.n6614 VPWR 0.0603958
R10471 VPWR.n6615 VPWR 0.0603958
R10472 VPWR VPWR.n6632 0.0603958
R10473 VPWR.n6633 VPWR 0.0603958
R10474 VPWR.n6637 VPWR 0.0603958
R10475 VPWR VPWR.n6763 0.0603958
R10476 VPWR VPWR.n6739 0.0603958
R10477 VPWR VPWR.n6691 0.0603958
R10478 VPWR.n8330 VPWR 0.0603958
R10479 VPWR.n8315 VPWR 0.0603958
R10480 VPWR VPWR.n8314 0.0603958
R10481 VPWR.n8303 VPWR 0.0603958
R10482 VPWR VPWR.n8302 0.0603958
R10483 VPWR VPWR.n8292 0.0603958
R10484 VPWR.n8288 VPWR 0.0603958
R10485 VPWR VPWR.n8287 0.0603958
R10486 VPWR.n8281 VPWR 0.0603958
R10487 VPWR.n8259 VPWR 0.0603958
R10488 VPWR VPWR.n8258 0.0603958
R10489 VPWR.n8199 VPWR 0.0603958
R10490 VPWR VPWR.n8198 0.0603958
R10491 VPWR.n8111 VPWR 0.0603958
R10492 VPWR.n8127 VPWR 0.0603958
R10493 VPWR.n8140 VPWR 0.0603958
R10494 VPWR.n8143 VPWR 0.0603958
R10495 VPWR.n8153 VPWR 0.0603958
R10496 VPWR.n8167 VPWR 0.0603958
R10497 VPWR.n8183 VPWR 0.0603958
R10498 VPWR.n8832 VPWR 0.0603958
R10499 VPWR.n8903 VPWR 0.0603958
R10500 VPWR.n8895 VPWR 0.0603958
R10501 VPWR.n8893 VPWR 0.0603958
R10502 VPWR VPWR.n8892 0.0603958
R10503 VPWR VPWR.n8889 0.0603958
R10504 VPWR.n6503 VPWR 0.0603958
R10505 VPWR.n6514 VPWR 0.0603958
R10506 VPWR.n6520 VPWR 0.0603958
R10507 VPWR.n6524 VPWR 0.0603958
R10508 VPWR.n6533 VPWR 0.0603958
R10509 VPWR.n6543 VPWR 0.0603958
R10510 VPWR.n6350 VPWR 0.0603958
R10511 VPWR.n6365 VPWR 0.0603958
R10512 VPWR.n6382 VPWR 0.0603958
R10513 VPWR.n6386 VPWR 0.0603958
R10514 VPWR.n6388 VPWR 0.0603958
R10515 VPWR.n6409 VPWR 0.0603958
R10516 VPWR.n6410 VPWR 0.0603958
R10517 VPWR.n6414 VPWR 0.0603958
R10518 VPWR.n6418 VPWR 0.0603958
R10519 VPWR.n6420 VPWR 0.0603958
R10520 VPWR.n6444 VPWR 0.0603958
R10521 VPWR VPWR.n6443 0.0603958
R10522 VPWR.n8426 VPWR 0.0603958
R10523 VPWR.n8428 VPWR 0.0603958
R10524 VPWR VPWR.n8435 0.0603958
R10525 VPWR.n8436 VPWR 0.0603958
R10526 VPWR.n8446 VPWR 0.0603958
R10527 VPWR.n8463 VPWR 0.0603958
R10528 VPWR.n8464 VPWR 0.0603958
R10529 VPWR.n8465 VPWR 0.0603958
R10530 VPWR.n8469 VPWR 0.0603958
R10531 VPWR.n8488 VPWR 0.0603958
R10532 VPWR VPWR.n8494 0.0603958
R10533 VPWR.n8495 VPWR 0.0603958
R10534 VPWR VPWR.n8495 0.0603958
R10535 VPWR.n8496 VPWR 0.0603958
R10536 VPWR.n8501 VPWR 0.0603958
R10537 VPWR.n8606 VPWR 0.0603958
R10538 VPWR.n8609 VPWR 0.0603958
R10539 VPWR VPWR.n8609 0.0603958
R10540 VPWR.n8610 VPWR 0.0603958
R10541 VPWR VPWR.n8671 0.0603958
R10542 VPWR.n8654 VPWR 0.0603958
R10543 VPWR VPWR.n8642 0.0603958
R10544 VPWR VPWR.n8641 0.0603958
R10545 VPWR.n8631 VPWR 0.0603958
R10546 VPWR.n8680 VPWR 0.0603958
R10547 VPWR.n8681 VPWR 0.0603958
R10548 VPWR.n8682 VPWR 0.0603958
R10549 VPWR.n8685 VPWR 0.0603958
R10550 VPWR.n8771 VPWR 0.0603958
R10551 VPWR.n8769 VPWR 0.0603958
R10552 VPWR.n8765 VPWR 0.0603958
R10553 VPWR.n8761 VPWR 0.0603958
R10554 VPWR VPWR.n8759 0.0603958
R10555 VPWR.n611 VPWR 0.0603958
R10556 VPWR VPWR.n618 0.0603958
R10557 VPWR.n620 VPWR 0.0603958
R10558 VPWR.n624 VPWR 0.0603958
R10559 VPWR VPWR.n637 0.0603958
R10560 VPWR.n638 VPWR 0.0603958
R10561 VPWR.n643 VPWR 0.0603958
R10562 VPWR.n713 VPWR 0.0603958
R10563 VPWR.n826 VPWR 0.0603958
R10564 VPWR.n839 VPWR 0.0603958
R10565 VPWR.n849 VPWR 0.0603958
R10566 VPWR.n858 VPWR 0.0603958
R10567 VPWR.n864 VPWR 0.0603958
R10568 VPWR.n865 VPWR 0.0603958
R10569 VPWR VPWR.n865 0.0603958
R10570 VPWR.n866 VPWR 0.0603958
R10571 VPWR.n871 VPWR 0.0603958
R10572 VPWR.n937 VPWR 0.0603958
R10573 VPWR.n945 VPWR 0.0603958
R10574 VPWR VPWR.n762 0.0603958
R10575 VPWR.n955 VPWR 0.0603958
R10576 VPWR.n962 VPWR 0.0603958
R10577 VPWR.n969 VPWR 0.0603958
R10578 VPWR.n991 VPWR 0.0603958
R10579 VPWR.n994 VPWR 0.0603958
R10580 VPWR.n1027 VPWR 0.0603958
R10581 VPWR.n1031 VPWR 0.0603958
R10582 VPWR.n1112 VPWR 0.0603958
R10583 VPWR VPWR.n1114 0.0603958
R10584 VPWR.n1116 VPWR 0.0603958
R10585 VPWR.n1119 VPWR 0.0603958
R10586 VPWR.n1128 VPWR 0.0603958
R10587 VPWR.n1129 VPWR 0.0603958
R10588 VPWR.n1136 VPWR 0.0603958
R10589 VPWR.n1200 VPWR 0.0603958
R10590 VPWR VPWR.n1199 0.0603958
R10591 VPWR VPWR.n1198 0.0603958
R10592 VPWR.n5819 VPWR 0.0603958
R10593 VPWR.n5815 VPWR 0.0603958
R10594 VPWR.n5803 VPWR 0.0603958
R10595 VPWR VPWR.n5799 0.0603958
R10596 VPWR VPWR.n1285 0.0603958
R10597 VPWR.n1300 VPWR 0.0603958
R10598 VPWR.n1308 VPWR 0.0603958
R10599 VPWR.n1318 VPWR 0.0603958
R10600 VPWR.n1498 VPWR 0.0603958
R10601 VPWR VPWR.n1497 0.0603958
R10602 VPWR.n1493 VPWR 0.0603958
R10603 VPWR.n1448 VPWR 0.0603958
R10604 VPWR VPWR.n1447 0.0603958
R10605 VPWR.n1438 VPWR 0.0603958
R10606 VPWR.n1433 VPWR 0.0603958
R10607 VPWR VPWR.n1432 0.0603958
R10608 VPWR VPWR.n1430 0.0603958
R10609 VPWR.n5414 VPWR 0.0603958
R10610 VPWR.n5436 VPWR 0.0603958
R10611 VPWR.n5439 VPWR 0.0603958
R10612 VPWR.n5444 VPWR 0.0603958
R10613 VPWR.n5454 VPWR 0.0603958
R10614 VPWR.n5456 VPWR 0.0603958
R10615 VPWR.n5455 VPWR 0.0603958
R10616 VPWR.n5464 VPWR 0.0603958
R10617 VPWR.n5469 VPWR 0.0603958
R10618 VPWR.n5484 VPWR 0.0603958
R10619 VPWR.n5488 VPWR 0.0603958
R10620 VPWR.n5492 VPWR 0.0603958
R10621 VPWR.n5594 VPWR 0.0603958
R10622 VPWR VPWR.n462 0.0603958
R10623 VPWR.n5608 VPWR 0.0603958
R10624 VPWR.n5610 VPWR 0.0603958
R10625 VPWR.n5616 VPWR 0.0603958
R10626 VPWR.n5620 VPWR 0.0603958
R10627 VPWR VPWR.n5625 0.0603958
R10628 VPWR.n5626 VPWR 0.0603958
R10629 VPWR.n5630 VPWR 0.0603958
R10630 VPWR.n5640 VPWR 0.0603958
R10631 VPWR.n5641 VPWR 0.0603958
R10632 VPWR.n440 VPWR 0.0603958
R10633 VPWR.n424 VPWR 0.0603958
R10634 VPWR.n1555 VPWR 0.0603958
R10635 VPWR.n1559 VPWR 0.0603958
R10636 VPWR VPWR.n1544 0.0603958
R10637 VPWR.n1572 VPWR 0.0603958
R10638 VPWR.n1573 VPWR 0.0603958
R10639 VPWR.n1576 VPWR 0.0603958
R10640 VPWR.n1660 VPWR 0.0603958
R10641 VPWR.n1663 VPWR 0.0603958
R10642 VPWR.n1672 VPWR 0.0603958
R10643 VPWR.n1688 VPWR 0.0603958
R10644 VPWR.n1712 VPWR 0.0603958
R10645 VPWR VPWR.n1717 0.0603958
R10646 VPWR.n1718 VPWR 0.0603958
R10647 VPWR VPWR.n550 0.0603958
R10648 VPWR.n1774 VPWR 0.0603958
R10649 VPWR VPWR.n1773 0.0603958
R10650 VPWR VPWR.n5319 0.0603958
R10651 VPWR.n5315 VPWR 0.0603958
R10652 VPWR.n5311 VPWR 0.0603958
R10653 VPWR.n5294 VPWR 0.0603958
R10654 VPWR VPWR.n5293 0.0603958
R10655 VPWR VPWR.n5291 0.0603958
R10656 VPWR.n5288 VPWR 0.0603958
R10657 VPWR VPWR.n5287 0.0603958
R10658 VPWR.n5281 VPWR 0.0603958
R10659 VPWR.n5279 VPWR 0.0603958
R10660 VPWR VPWR.n5278 0.0603958
R10661 VPWR VPWR.n5277 0.0603958
R10662 VPWR.n5274 VPWR 0.0603958
R10663 VPWR.n4686 VPWR 0.0603958
R10664 VPWR.n4687 VPWR 0.0603958
R10665 VPWR.n4763 VPWR 0.0603958
R10666 VPWR VPWR.n4762 0.0603958
R10667 VPWR.n4755 VPWR 0.0603958
R10668 VPWR VPWR.n4754 0.0603958
R10669 VPWR VPWR.n4753 0.0603958
R10670 VPWR.n4751 VPWR 0.0603958
R10671 VPWR.n4748 VPWR 0.0603958
R10672 VPWR.n4728 VPWR 0.0603958
R10673 VPWR.n4723 VPWR 0.0603958
R10674 VPWR.n4716 VPWR 0.0603958
R10675 VPWR VPWR.n4715 0.0603958
R10676 VPWR VPWR.n4646 0.0603958
R10677 VPWR.n4768 VPWR 0.0603958
R10678 VPWR.n4769 VPWR 0.0603958
R10679 VPWR.n4774 VPWR 0.0603958
R10680 VPWR.n4834 VPWR 0.0603958
R10681 VPWR VPWR.n4825 0.0603958
R10682 VPWR.n4822 VPWR 0.0603958
R10683 VPWR.n4820 VPWR 0.0603958
R10684 VPWR.n4817 VPWR 0.0603958
R10685 VPWR VPWR.n4816 0.0603958
R10686 VPWR.n2442 VPWR 0.0603958
R10687 VPWR.n2443 VPWR 0.0603958
R10688 VPWR.n2447 VPWR 0.0603958
R10689 VPWR.n2451 VPWR 0.0603958
R10690 VPWR VPWR.n2452 0.0603958
R10691 VPWR.n2454 VPWR 0.0603958
R10692 VPWR VPWR.n2453 0.0603958
R10693 VPWR.n2463 VPWR 0.0603958
R10694 VPWR.n2464 VPWR 0.0603958
R10695 VPWR VPWR.n2470 0.0603958
R10696 VPWR.n2471 VPWR 0.0603958
R10697 VPWR.n2476 VPWR 0.0603958
R10698 VPWR.n2551 VPWR 0.0603958
R10699 VPWR.n2557 VPWR 0.0603958
R10700 VPWR VPWR.n2186 0.0603958
R10701 VPWR VPWR.n2184 0.0603958
R10702 VPWR VPWR.n2139 0.0603958
R10703 VPWR.n2135 VPWR 0.0603958
R10704 VPWR VPWR.n2125 0.0603958
R10705 VPWR.n2570 VPWR 0.0603958
R10706 VPWR.n2571 VPWR 0.0603958
R10707 VPWR.n2574 VPWR 0.0603958
R10708 VPWR.n5153 VPWR 0.0603958
R10709 VPWR.n1838 VPWR 0.0603958
R10710 VPWR VPWR.n1838 0.0603958
R10711 VPWR.n5140 VPWR 0.0603958
R10712 VPWR VPWR.n5139 0.0603958
R10713 VPWR VPWR.n5138 0.0603958
R10714 VPWR.n5122 VPWR 0.0603958
R10715 VPWR.n5117 VPWR 0.0603958
R10716 VPWR VPWR.n5116 0.0603958
R10717 VPWR VPWR.n5113 0.0603958
R10718 VPWR VPWR.n5112 0.0603958
R10719 VPWR VPWR.n5111 0.0603958
R10720 VPWR.n5099 VPWR 0.0603958
R10721 VPWR.n5087 VPWR 0.0603958
R10722 VPWR VPWR.n5086 0.0603958
R10723 VPWR VPWR.n5029 0.0603958
R10724 VPWR.n5020 VPWR 0.0603958
R10725 VPWR.n5020 VPWR 0.0603958
R10726 VPWR VPWR.n5019 0.0603958
R10727 VPWR.n1912 VPWR 0.0603958
R10728 VPWR.n1914 VPWR 0.0603958
R10729 VPWR.n1927 VPWR 0.0603958
R10730 VPWR VPWR.n1909 0.0603958
R10731 VPWR.n1933 VPWR 0.0603958
R10732 VPWR VPWR.n1948 0.0603958
R10733 VPWR.n1949 VPWR 0.0603958
R10734 VPWR.n1958 VPWR 0.0603958
R10735 VPWR.n1960 VPWR 0.0603958
R10736 VPWR VPWR.n5010 0.0603958
R10737 VPWR.n4954 VPWR 0.0603958
R10738 VPWR.n4935 VPWR 0.0603958
R10739 VPWR VPWR.n4934 0.0603958
R10740 VPWR.n2224 VPWR 0.0603958
R10741 VPWR.n2232 VPWR 0.0603958
R10742 VPWR.n2242 VPWR 0.0603958
R10743 VPWR.n2255 VPWR 0.0603958
R10744 VPWR.n2261 VPWR 0.0603958
R10745 VPWR VPWR.n2377 0.0603958
R10746 VPWR.n2371 VPWR 0.0603958
R10747 VPWR VPWR.n2370 0.0603958
R10748 VPWR VPWR.n2369 0.0603958
R10749 VPWR.n2363 VPWR 0.0603958
R10750 VPWR VPWR.n2330 0.0603958
R10751 VPWR.n2325 VPWR 0.0603958
R10752 VPWR.n2321 VPWR 0.0603958
R10753 VPWR VPWR.n2319 0.0603958
R10754 VPWR.n2319 VPWR 0.0603958
R10755 VPWR VPWR.n2317 0.0603958
R10756 VPWR.n2688 VPWR 0.0603958
R10757 VPWR VPWR.n2687 0.0603958
R10758 VPWR VPWR.n2060 0.0603958
R10759 VPWR VPWR.n2046 0.0603958
R10760 VPWR VPWR.n2032 0.0603958
R10761 VPWR.n2697 VPWR 0.0603958
R10762 VPWR.n2702 VPWR 0.0603958
R10763 VPWR VPWR.n2716 0.0603958
R10764 VPWR.n2717 VPWR 0.0603958
R10765 VPWR.n2721 VPWR 0.0603958
R10766 VPWR.n2725 VPWR 0.0603958
R10767 VPWR VPWR.n4409 0.0603958
R10768 VPWR.n4411 VPWR 0.0603958
R10769 VPWR.n4419 VPWR 0.0603958
R10770 VPWR.n4426 VPWR 0.0603958
R10771 VPWR.n4427 VPWR 0.0603958
R10772 VPWR.n4437 VPWR 0.0603958
R10773 VPWR.n4453 VPWR 0.0603958
R10774 VPWR.n4455 VPWR 0.0603958
R10775 VPWR.n4468 VPWR 0.0603958
R10776 VPWR.n4476 VPWR 0.0603958
R10777 VPWR.n4480 VPWR 0.0603958
R10778 VPWR.n4535 VPWR 0.0603958
R10779 VPWR VPWR.n4534 0.0603958
R10780 VPWR.n4517 VPWR 0.0603958
R10781 VPWR.n4515 VPWR 0.0603958
R10782 VPWR.n4512 VPWR 0.0603958
R10783 VPWR.n3388 VPWR 0.0603958
R10784 VPWR.n3398 VPWR 0.0603958
R10785 VPWR.n3409 VPWR 0.0603958
R10786 VPWR.n3410 VPWR 0.0603958
R10787 VPWR.n3415 VPWR 0.0603958
R10788 VPWR VPWR.n3415 0.0603958
R10789 VPWR.n3416 VPWR 0.0603958
R10790 VPWR.n3421 VPWR 0.0603958
R10791 VPWR.n3743 VPWR 0.0603958
R10792 VPWR.n3739 VPWR 0.0603958
R10793 VPWR.n3735 VPWR 0.0603958
R10794 VPWR VPWR.n3734 0.0603958
R10795 VPWR VPWR.n3732 0.0603958
R10796 VPWR VPWR.n3731 0.0603958
R10797 VPWR VPWR.n3728 0.0603958
R10798 VPWR.n3718 VPWR 0.0603958
R10799 VPWR.n3689 VPWR 0.0603958
R10800 VPWR.n3677 VPWR 0.0603958
R10801 VPWR.n3518 VPWR 0.0603958
R10802 VPWR.n3535 VPWR 0.0603958
R10803 VPWR.n3538 VPWR 0.0603958
R10804 VPWR.n3586 VPWR 0.0603958
R10805 VPWR.n3597 VPWR 0.0603958
R10806 VPWR.n3611 VPWR 0.0603958
R10807 VPWR VPWR.n3670 0.0603958
R10808 VPWR.n3667 VPWR 0.0603958
R10809 VPWR.n3661 VPWR 0.0603958
R10810 VPWR.n3644 VPWR 0.0603958
R10811 VPWR.n3641 VPWR 0.0603958
R10812 VPWR.n2797 VPWR 0.0603958
R10813 VPWR.n2802 VPWR 0.0603958
R10814 VPWR.n2821 VPWR 0.0603958
R10815 VPWR.n2836 VPWR 0.0603958
R10816 VPWR VPWR.n4245 0.0603958
R10817 VPWR VPWR.n4244 0.0603958
R10818 VPWR.n2920 VPWR 0.0603958
R10819 VPWR.n7657 VPWR 0.0603958
R10820 VPWR.n7663 VPWR 0.0603958
R10821 VPWR.n7669 VPWR 0.0603958
R10822 VPWR.n7672 VPWR 0.0603958
R10823 VPWR.n7755 VPWR 0.0603958
R10824 VPWR.n7769 VPWR 0.0603958
R10825 VPWR.n7812 VPWR 0.0603958
R10826 VPWR.n6046 VPWR 0.0603958
R10827 VPWR.n6056 VPWR 0.0603958
R10828 VPWR.n6107 VPWR 0.0603958
R10829 VPWR VPWR.n6106 0.0603958
R10830 VPWR VPWR.n6105 0.0603958
R10831 VPWR.n6087 VPWR 0.0603958
R10832 VPWR.n6080 VPWR 0.0603958
R10833 VPWR VPWR.n6079 0.0603958
R10834 VPWR.n6073 VPWR 0.0603958
R10835 VPWR VPWR.n6072 0.0603958
R10836 VPWR.n9199 VPWR 0.0603958
R10837 VPWR VPWR.n9198 0.0603958
R10838 VPWR VPWR.n9197 0.0603958
R10839 VPWR.n9191 VPWR 0.0603958
R10840 VPWR.n9184 VPWR 0.0603958
R10841 VPWR.n9177 VPWR 0.0603958
R10842 VPWR VPWR.n9169 0.0603958
R10843 VPWR.n9166 VPWR 0.0603958
R10844 VPWR.n9160 VPWR 0.0603958
R10845 VPWR.n9155 VPWR 0.0603958
R10846 VPWR VPWR.n9154 0.0603958
R10847 VPWR VPWR.n9153 0.0603958
R10848 VPWR.n9143 VPWR 0.0603958
R10849 VPWR VPWR.n9142 0.0603958
R10850 VPWR.n9130 VPWR 0.0603958
R10851 VPWR.n105 VPWR 0.0603958
R10852 VPWR.n92 VPWR 0.0603958
R10853 VPWR VPWR.n91 0.0603958
R10854 VPWR.n88 VPWR 0.0603958
R10855 VPWR VPWR.n86 0.0603958
R10856 VPWR VPWR.n84 0.0603958
R10857 VPWR.n3253 VPWR 0.0603958
R10858 VPWR.n3259 VPWR 0.0603958
R10859 VPWR.n3263 VPWR 0.0603958
R10860 VPWR.n3264 VPWR 0.0603958
R10861 VPWR.n3267 VPWR 0.0603958
R10862 VPWR.n3282 VPWR 0.0603958
R10863 VPWR.n3289 VPWR 0.0603958
R10864 VPWR.n3212 VPWR 0.0603958
R10865 VPWR VPWR.n3210 0.0603958
R10866 VPWR.n3204 VPWR 0.0603958
R10867 VPWR.n3199 VPWR 0.0603958
R10868 VPWR VPWR.n3172 0.0603958
R10869 VPWR VPWR.n3170 0.0603958
R10870 VPWR.n3164 VPWR 0.0603958
R10871 VPWR VPWR.n3163 0.0603958
R10872 VPWR.n3875 VPWR 0.0603958
R10873 VPWR VPWR.n3874 0.0603958
R10874 VPWR VPWR.n3872 0.0603958
R10875 VPWR.n3872 VPWR 0.0603958
R10876 VPWR.n3087 VPWR 0.0603958
R10877 VPWR VPWR.n3086 0.0603958
R10878 VPWR VPWR.n3074 0.0603958
R10879 VPWR VPWR.n3073 0.0603958
R10880 VPWR.n3060 VPWR 0.0603958
R10881 VPWR VPWR.n3060 0.0603958
R10882 VPWR.n3882 VPWR 0.0603958
R10883 VPWR.n3884 VPWR 0.0603958
R10884 VPWR.n3889 VPWR 0.0603958
R10885 VPWR.n4004 VPWR 0.0603958
R10886 VPWR.n4018 VPWR 0.0603958
R10887 VPWR.n4034 VPWR 0.0603958
R10888 VPWR.n4063 VPWR 0.0603958
R10889 VPWR.n4063 VPWR 0.0603958
R10890 VPWR.n4066 VPWR 0.0603958
R10891 VPWR.n4071 VPWR 0.0603958
R10892 VPWR.n4072 VPWR 0.0603958
R10893 VPWR.n4077 VPWR 0.0603958
R10894 VPWR.n4121 VPWR 0.0603958
R10895 VPWR.n4090 VPWR 0.0603958
R10896 VPWR VPWR.n4109 0.0603958
R10897 VPWR.n7533 VPWR 0.0603958
R10898 VPWR.n7536 VPWR 0.0603958
R10899 VPWR.n7550 VPWR 0.0603958
R10900 VPWR.n7554 VPWR 0.0603958
R10901 VPWR.n7566 VPWR 0.0603958
R10902 VPWR.n7572 VPWR 0.0603958
R10903 VPWR VPWR.n7511 0.0603958
R10904 VPWR.n7504 VPWR 0.0603958
R10905 VPWR VPWR.n7503 0.0603958
R10906 VPWR.n7497 VPWR 0.0603958
R10907 VPWR.n7465 VPWR 0.0603958
R10908 VPWR VPWR.n7464 0.0603958
R10909 VPWR.n7459 VPWR 0.0603958
R10910 VPWR VPWR.n7458 0.0603958
R10911 VPWR.n7454 VPWR 0.0603958
R10912 VPWR.n7396 VPWR 0.0603958
R10913 VPWR VPWR.n7395 0.0603958
R10914 VPWR.n7392 VPWR 0.0603958
R10915 VPWR.n7378 VPWR 0.0603958
R10916 VPWR VPWR.n7377 0.0603958
R10917 VPWR.n7371 VPWR 0.0603958
R10918 VPWR.n7361 VPWR 0.0603958
R10919 VPWR VPWR.n7360 0.0603958
R10920 VPWR.n7354 VPWR 0.0603958
R10921 VPWR.n7068 VPWR 0.0603958
R10922 VPWR.n7069 VPWR 0.0603958
R10923 VPWR.n7076 VPWR 0.0603958
R10924 VPWR.n7083 VPWR 0.0603958
R10925 VPWR.n7112 VPWR 0.0603958
R10926 VPWR VPWR.n7125 0.0603958
R10927 VPWR.n7126 VPWR 0.0603958
R10928 VPWR.n7129 VPWR 0.0603958
R10929 VPWR.n7276 VPWR 0.0603958
R10930 VPWR.n7186 VPWR 0.0603958
R10931 VPWR VPWR.n7185 0.0603958
R10932 VPWR.n7175 VPWR 0.0603958
R10933 VPWR VPWR.n7174 0.0603958
R10934 VPWR.n7171 VPWR 0.0603958
R10935 VPWR.n7164 VPWR 0.0603958
R10936 VPWR VPWR.n7163 0.0603958
R10937 VPWR.n4984 VPWR.n4983 0.059272
R10938 VPWR.n5664 VPWR.n5653 0.0590938
R10939 VPWR.n2278 VPWR.n2276 0.0586222
R10940 VPWR.n6461 VPWR.n6460 0.0577917
R10941 VPWR.n1226 VPWR.n1224 0.0577917
R10942 VPWR.n1518 VPWR.n1517 0.0577917
R10943 VPWR.n3748 VPWR.n3746 0.0577917
R10944 VPWR.n6206 VPWR.n6199 0.0561015
R10945 VPWR.n6827 VPWR.n6639 0.0561015
R10946 VPWR.n6550 VPWR.n6543 0.0561015
R10947 VPWR.n1609 VPWR.n1586 0.0561015
R10948 VPWR.n2496 VPWR.n2482 0.0561015
R10949 VPWR.n2276 VPWR.n2269 0.0561015
R10950 VPWR.n3446 VPWR.n3424 0.0561015
R10951 VPWR.n3292 VPWR.n3291 0.0561015
R10952 VPWR.n7575 VPWR.n7574 0.0561015
R10953 VPWR.n7724 VPWR.n7686 0.0561015
R10954 VPWR.n3758 VPWR.n3756 0.0548679
R10955 VPWR.n114 VPWR.n113 0.0547995
R10956 VPWR.n5701 VPWR.n450 0.0547995
R10957 VPWR.n4843 VPWR.n4842 0.0547995
R10958 VPWR.n4984 VPWR.n4966 0.0547995
R10959 VPWR.n4540 VPWR.n4539 0.0547995
R10960 VPWR.n2966 VPWR.n2935 0.0547995
R10961 VPWR.n4136 VPWR.n4135 0.0547995
R10962 VPWR.n3053 VPWR.n3052 0.0512937
R10963 VPWR.n111 VPWR.n110 0.0512937
R10964 VPWR.n8306 VPWR.n5933 0.0512937
R10965 VPWR.n8755 VPWR.n8754 0.0512937
R10966 VPWR.n8638 VPWR.n8637 0.0512937
R10967 VPWR.n6561 VPWR.n6560 0.0512937
R10968 VPWR.n6471 VPWR.n6470 0.0512937
R10969 VPWR.n384 VPWR.n383 0.0512937
R10970 VPWR.n694 VPWR.n693 0.0512937
R10971 VPWR.n1593 VPWR.n1592 0.0512937
R10972 VPWR.n3451 VPWR.n3450 0.0512937
R10973 VPWR.n3461 VPWR.n3460 0.0512937
R10974 VPWR.n7325 VPWR 0.0497858
R10975 VPWR.n6207 VPWR.n6206 0.0496664
R10976 VPWR.n6827 VPWR.n6826 0.0496664
R10977 VPWR.n6551 VPWR.n6550 0.0496664
R10978 VPWR.n1335 VPWR.n1333 0.0496664
R10979 VPWR.n5701 VPWR.n5700 0.0496664
R10980 VPWR.n1609 VPWR.n1608 0.0496664
R10981 VPWR.n4844 VPWR.n4843 0.0496664
R10982 VPWR.n2496 VPWR.n2495 0.0496664
R10983 VPWR.n4541 VPWR.n4540 0.0496664
R10984 VPWR.n3447 VPWR.n3446 0.0496664
R10985 VPWR.n2966 VPWR.n2965 0.0496664
R10986 VPWR.n7724 VPWR.n7723 0.0496664
R10987 VPWR.n115 VPWR.n114 0.0496664
R10988 VPWR.n3294 VPWR.n3292 0.0496664
R10989 VPWR.n4138 VPWR.n4136 0.0496664
R10990 VPWR.n7577 VPWR.n7575 0.0496664
R10991 VPWR VPWR.n6690 0.047375
R10992 VPWR.n2578 VPWR 0.047375
R10993 VPWR.n3868 VPWR 0.047375
R10994 VPWR.n8001 VPWR.n8000 0.0460729
R10995 VPWR.n6684 VPWR.n6683 0.0460729
R10996 VPWR.n8108 VPWR.n8107 0.0460729
R10997 VPWR.n879 VPWR.n878 0.0460729
R10998 VPWR.n738 VPWR.n737 0.0460729
R10999 VPWR.n1417 VPWR.n1416 0.0460729
R11000 VPWR.n5568 VPWR.n5567 0.0460729
R11001 VPWR.n4667 VPWR.n4666 0.0460729
R11002 VPWR.n4392 VPWR.n4391 0.0460729
R11003 VPWR.n3551 VPWR.n3550 0.0460729
R11004 VPWR.n4274 VPWR.n4273 0.0460729
R11005 VPWR.n7827 VPWR.n7826 0.0460729
R11006 VPWR.n3860 VPWR.n3859 0.0460729
R11007 VPWR.n7444 VPWR.n7443 0.0460729
R11008 VPWR.n5857 VPWR.n5856 0.0460313
R11009 VPWR.n653 VPWR.n646 0.0446272
R11010 VPWR.n7194 VPWR.n7193 0.0433251
R11011 VPWR.n258 VPWR.n257 0.0433251
R11012 VPWR.n8917 VPWR.n8916 0.0433251
R11013 VPWR.n8789 VPWR.n8788 0.0433251
R11014 VPWR.n5829 VPWR.n5828 0.0433251
R11015 VPWR.n6214 VPWR.n6213 0.0421667
R11016 VPWR.n280 VPWR.n279 0.0421667
R11017 VPWR.n6817 VPWR.n6816 0.0421667
R11018 VPWR.n8932 VPWR.n8931 0.0421667
R11019 VPWR.n666 VPWR.n665 0.0421667
R11020 VPWR.n5842 VPWR.n5841 0.0421667
R11021 VPWR.n1344 VPWR.n1343 0.0421667
R11022 VPWR.n5691 VPWR.n5690 0.0421667
R11023 VPWR.n1598 VPWR.n1597 0.0421667
R11024 VPWR.n4851 VPWR.n4850 0.0421667
R11025 VPWR.n4978 VPWR.n4977 0.0421667
R11026 VPWR.n2284 VPWR.n2283 0.0421667
R11027 VPWR.n4552 VPWR.n4551 0.0421667
R11028 VPWR.n3457 VPWR.n3456 0.0421667
R11029 VPWR.n7717 VPWR.n7716 0.0421667
R11030 VPWR.n124 VPWR.n123 0.0421667
R11031 VPWR.n3305 VPWR.n3304 0.0421667
R11032 VPWR.n4147 VPWR.n4146 0.0421667
R11033 VPWR.n7586 VPWR.n7585 0.0421667
R11034 VPWR.n7215 VPWR.n7214 0.0421667
R11035 VPWR.n656 VPWR.n654 0.0408646
R11036 VPWR.n3132 VPWR.n3131 0.0393514
R11037 VPWR.n146 VPWR.n144 0.0393514
R11038 VPWR.n297 VPWR.n205 0.0393514
R11039 VPWR.n6204 VPWR.n6200 0.0393514
R11040 VPWR.n8862 VPWR.n8856 0.0393514
R11041 VPWR.n6830 VPWR.n6829 0.0393514
R11042 VPWR.n8731 VPWR.n8725 0.0393514
R11043 VPWR.n6548 VPWR.n6544 0.0393514
R11044 VPWR.n5773 VPWR.n5767 0.0393514
R11045 VPWR.n651 VPWR.n647 0.0393514
R11046 VPWR.n5703 VPWR.n400 0.0393514
R11047 VPWR.n1331 VPWR.n1327 0.0393514
R11048 VPWR.n4629 VPWR.n4627 0.0393514
R11049 VPWR.n1612 VPWR.n1611 0.0393514
R11050 VPWR.n4986 VPWR.n4911 0.0393514
R11051 VPWR.n2499 VPWR.n2498 0.0393514
R11052 VPWR.n2274 VPWR.n2270 0.0393514
R11053 VPWR.n1973 VPWR.n1971 0.0393514
R11054 VPWR.n2968 VPWR.n2885 0.0393514
R11055 VPWR.n7727 VPWR.n7726 0.0393514
R11056 VPWR.n6920 VPWR.n6919 0.0393514
R11057 VPWR.n2981 VPWR.n2979 0.0393514
R11058 VPWR.n7228 VPWR.n7146 0.0393514
R11059 VPWR.n7712 VPWR.n7711 0.0382581
R11060 VPWR.n6219 VPWR.n6218 0.0382581
R11061 VPWR.n4531 VPWR.n4530 0.0382581
R11062 VPWR.n295 VPWR 0.0369583
R11063 VPWR VPWR.n8919 0.0369583
R11064 VPWR VPWR.n5742 0.0369583
R11065 VPWR.n4997 VPWR 0.0369583
R11066 VPWR.n7226 VPWR 0.0369583
R11067 VPWR.n7958 VPWR.n7957 0.035973
R11068 VPWR.n6661 VPWR.n6660 0.0356562
R11069 VPWR.n8251 VPWR.n8250 0.0356562
R11070 VPWR.n8385 VPWR.n8384 0.0356562
R11071 VPWR.n8565 VPWR.n8564 0.0356562
R11072 VPWR.n1084 VPWR.n1083 0.0356562
R11073 VPWR.n1730 VPWR.n1729 0.0356562
R11074 VPWR.n5164 VPWR.n5163 0.0356562
R11075 VPWR.n2643 VPWR.n2642 0.0356562
R11076 VPWR.n4367 VPWR.n4366 0.0356562
R11077 VPWR.n3569 VPWR.n3568 0.0356562
R11078 VPWR.n4298 VPWR.n4297 0.0356562
R11079 VPWR.n7851 VPWR.n7850 0.0356562
R11080 VPWR.n3835 VPWR.n3834 0.0356562
R11081 VPWR.n3943 VPWR.n3942 0.0356562
R11082 VPWR.n7421 VPWR.n7420 0.0356562
R11083 VPWR.n7347 VPWR.n7346 0.0356562
R11084 VPWR VPWR.n7962 0.0343542
R11085 VPWR.n271 VPWR.n269 0.0343542
R11086 VPWR.n8847 VPWR.n8845 0.0343542
R11087 VPWR.n6480 VPWR.n6478 0.0343542
R11088 VPWR.n8712 VPWR.n8710 0.0343542
R11089 VPWR VPWR.n906 0.0343542
R11090 VPWR.n5760 VPWR.n5759 0.0343542
R11091 VPWR.n1354 VPWR.n1353 0.0343542
R11092 VPWR.n5396 VPWR 0.0343542
R11093 VPWR.n5681 VPWR.n5679 0.0343542
R11094 VPWR.n4861 VPWR.n4860 0.0343542
R11095 VPWR.n4971 VPWR.n4970 0.0343542
R11096 VPWR.n4559 VPWR.n4558 0.0343542
R11097 VPWR.n2938 VPWR.n2936 0.0343542
R11098 VPWR.n133 VPWR.n132 0.0343542
R11099 VPWR.n3315 VPWR.n3314 0.0343542
R11100 VPWR.n4157 VPWR.n4156 0.0343542
R11101 VPWR.n7596 VPWR.n7595 0.0343542
R11102 VPWR.n7206 VPWR.n7204 0.0343542
R11103 VPWR.n9217 VPWR.n9216 0.0342838
R11104 VPWR.n9080 VPWR.n9079 0.0342838
R11105 VPWR.n7889 VPWR.n7888 0.0342838
R11106 VPWR.n8098 VPWR.n8097 0.0342838
R11107 VPWR.n8356 VPWR.n8355 0.0342838
R11108 VPWR.n8532 VPWR.n357 0.0342838
R11109 VPWR.n6428 VPWR.n6427 0.0342838
R11110 VPWR.n742 VPWR.n741 0.0342838
R11111 VPWR.n782 VPWR.n781 0.0342838
R11112 VPWR.n5528 VPWR.n5527 0.0342838
R11113 VPWR.n5365 VPWR.n5364 0.0342838
R11114 VPWR.n5219 VPWR.n5218 0.0342838
R11115 VPWR.n1757 VPWR.n1756 0.0342838
R11116 VPWR.n1885 VPWR.n1874 0.0342838
R11117 VPWR.n2593 VPWR.n2592 0.0342838
R11118 VPWR.n4346 VPWR.n4345 0.0342838
R11119 VPWR.n2039 VPWR.n2038 0.0342838
R11120 VPWR.n5983 VPWR.n5982 0.0342838
R11121 VPWR.n4311 VPWR.n4310 0.0342838
R11122 VPWR.n3117 VPWR.n3116 0.0342838
R11123 VPWR.n3105 VPWR.n3104 0.0342838
R11124 VPWR.n6997 VPWR.n6996 0.0342838
R11125 VPWR.n3002 VPWR.n3001 0.0342838
R11126 VPWR.n7300 VPWR.n2 0.0342838
R11127 VPWR.n6883 VPWR 0.0330521
R11128 VPWR.n8047 VPWR 0.0330521
R11129 VPWR.n8076 VPWR 0.0330521
R11130 VPWR.n225 VPWR 0.0330521
R11131 VPWR VPWR.n6805 0.0330521
R11132 VPWR.n8890 VPWR 0.0330521
R11133 VPWR VPWR.n6419 0.0330521
R11134 VPWR.n8630 VPWR 0.0330521
R11135 VPWR.n8682 VPWR 0.0330521
R11136 VPWR.n8764 VPWR 0.0330521
R11137 VPWR.n700 VPWR 0.0330521
R11138 VPWR.n866 VPWR 0.0330521
R11139 VPWR.n1496 VPWR 0.0330521
R11140 VPWR.n1431 VPWR 0.0330521
R11141 VPWR.n5438 VPWR 0.0330521
R11142 VPWR.n5509 VPWR 0.0330521
R11143 VPWR.n5611 VPWR 0.0330521
R11144 VPWR.n1556 VPWR 0.0330521
R11145 VPWR VPWR.n1579 0.0330521
R11146 VPWR.n1629 VPWR 0.0330521
R11147 VPWR VPWR.n1724 0.0330521
R11148 VPWR.n5292 VPWR 0.0330521
R11149 VPWR.n5249 VPWR 0.0330521
R11150 VPWR.n2533 VPWR 0.0330521
R11151 VPWR.n2552 VPWR 0.0330521
R11152 VPWR.n5121 VPWR 0.0330521
R11153 VPWR.n5081 VPWR 0.0330521
R11154 VPWR.n5030 VPWR 0.0330521
R11155 VPWR.n5011 VPWR 0.0330521
R11156 VPWR.n2256 VPWR 0.0330521
R11157 VPWR.n2399 VPWR 0.0330521
R11158 VPWR.n2366 VPWR 0.0330521
R11159 VPWR.n2324 VPWR 0.0330521
R11160 VPWR.n2317 VPWR 0.0330521
R11161 VPWR VPWR.n4482 0.0330521
R11162 VPWR.n3483 VPWR 0.0330521
R11163 VPWR.n3733 VPWR 0.0330521
R11164 VPWR.n3640 VPWR 0.0330521
R11165 VPWR.n2798 VPWR 0.0330521
R11166 VPWR VPWR.n7674 0.0330521
R11167 VPWR VPWR.n7705 0.0330521
R11168 VPWR.n9262 VPWR 0.0330521
R11169 VPWR.n9154 VPWR 0.0330521
R11170 VPWR.n9141 VPWR 0.0330521
R11171 VPWR.n82 VPWR 0.0330521
R11172 VPWR.n3203 VPWR 0.0330521
R11173 VPWR.n3873 VPWR 0.0330521
R11174 VPWR.n7551 VPWR 0.0330521
R11175 VPWR.n7462 VPWR 0.0330521
R11176 VPWR.n7457 VPWR 0.0330521
R11177 VPWR.n9093 VPWR.n9092 0.0325946
R11178 VPWR.n8221 VPWR.n8220 0.0325946
R11179 VPWR.n8555 VPWR.n8554 0.0325946
R11180 VPWR.n1074 VPWR.n1072 0.0325946
R11181 VPWR.n5556 VPWR.n5554 0.0325946
R11182 VPWR.n4655 VPWR.n4653 0.0325946
R11183 VPWR.n5066 VPWR.n5064 0.0325946
R11184 VPWR.n2746 VPWR.n2745 0.0325946
R11185 VPWR.n3811 VPWR.n3810 0.0325946
R11186 VPWR.n7312 VPWR.n7311 0.0325946
R11187 VPWR.n6296 VPWR 0.03175
R11188 VPWR.n8010 VPWR 0.03175
R11189 VPWR.n5965 VPWR 0.03175
R11190 VPWR VPWR.n194 0.03175
R11191 VPWR.n8972 VPWR 0.03175
R11192 VPWR.n241 VPWR 0.03175
R11193 VPWR VPWR.n6597 0.03175
R11194 VPWR VPWR.n6614 0.03175
R11195 VPWR.n6633 VPWR 0.03175
R11196 VPWR.n6764 VPWR 0.03175
R11197 VPWR.n6763 VPWR 0.03175
R11198 VPWR.n6693 VPWR 0.03175
R11199 VPWR.n8315 VPWR 0.03175
R11200 VPWR.n8292 VPWR 0.03175
R11201 VPWR.n8288 VPWR 0.03175
R11202 VPWR.n8259 VPWR 0.03175
R11203 VPWR VPWR.n8111 0.03175
R11204 VPWR.n8183 VPWR 0.03175
R11205 VPWR.n8832 VPWR 0.03175
R11206 VPWR.n6520 VPWR 0.03175
R11207 VPWR.n6533 VPWR 0.03175
R11208 VPWR VPWR.n6350 0.03175
R11209 VPWR VPWR.n6365 0.03175
R11210 VPWR VPWR.n6386 0.03175
R11211 VPWR VPWR.n6409 0.03175
R11212 VPWR VPWR.n6420 0.03175
R11213 VPWR.n6444 VPWR 0.03175
R11214 VPWR VPWR.n8464 0.03175
R11215 VPWR.n8465 VPWR 0.03175
R11216 VPWR.n8496 VPWR 0.03175
R11217 VPWR VPWR.n8610 0.03175
R11218 VPWR.n8642 VPWR 0.03175
R11219 VPWR VPWR.n8680 0.03175
R11220 VPWR.n638 VPWR 0.03175
R11221 VPWR VPWR.n713 0.03175
R11222 VPWR VPWR.n826 0.03175
R11223 VPWR VPWR.n849 0.03175
R11224 VPWR VPWR.n864 0.03175
R11225 VPWR.n762 VPWR 0.03175
R11226 VPWR VPWR.n991 0.03175
R11227 VPWR VPWR.n1116 0.03175
R11228 VPWR.n1200 VPWR 0.03175
R11229 VPWR.n1199 VPWR 0.03175
R11230 VPWR.n1498 VPWR 0.03175
R11231 VPWR.n1448 VPWR 0.03175
R11232 VPWR.n1433 VPWR 0.03175
R11233 VPWR VPWR.n5436 0.03175
R11234 VPWR VPWR.n5454 0.03175
R11235 VPWR.n5590 VPWR 0.03175
R11236 VPWR VPWR.n5594 0.03175
R11237 VPWR.n5626 VPWR 0.03175
R11238 VPWR VPWR.n5640 0.03175
R11239 VPWR.n1660 VPWR 0.03175
R11240 VPWR.n5288 VPWR 0.03175
R11241 VPWR.n5278 VPWR 0.03175
R11242 VPWR VPWR.n4687 0.03175
R11243 VPWR.n4763 VPWR 0.03175
R11244 VPWR.n4755 VPWR 0.03175
R11245 VPWR.n4715 VPWR 0.03175
R11246 VPWR.n4646 VPWR 0.03175
R11247 VPWR VPWR.n4768 0.03175
R11248 VPWR.n4825 VPWR 0.03175
R11249 VPWR.n4817 VPWR 0.03175
R11250 VPWR.n2454 VPWR 0.03175
R11251 VPWR.n2186 VPWR 0.03175
R11252 VPWR VPWR.n2570 0.03175
R11253 VPWR.n2571 VPWR 0.03175
R11254 VPWR.n5140 VPWR 0.03175
R11255 VPWR.n5116 VPWR 0.03175
R11256 VPWR.n5112 VPWR 0.03175
R11257 VPWR.n5087 VPWR 0.03175
R11258 VPWR.n5019 VPWR 0.03175
R11259 VPWR VPWR.n1949 0.03175
R11260 VPWR VPWR.n1958 0.03175
R11261 VPWR.n4935 VPWR 0.03175
R11262 VPWR.n2370 VPWR 0.03175
R11263 VPWR.n2688 VPWR 0.03175
R11264 VPWR.n2032 VPWR 0.03175
R11265 VPWR.n2717 VPWR 0.03175
R11266 VPWR VPWR.n4411 0.03175
R11267 VPWR.n4427 VPWR 0.03175
R11268 VPWR.n4476 VPWR 0.03175
R11269 VPWR.n3416 VPWR 0.03175
R11270 VPWR.n3732 VPWR 0.03175
R11271 VPWR.n3731 VPWR 0.03175
R11272 VPWR VPWR.n3518 0.03175
R11273 VPWR.n3535 VPWR 0.03175
R11274 VPWR.n3671 VPWR 0.03175
R11275 VPWR.n3670 VPWR 0.03175
R11276 VPWR VPWR.n2789 0.03175
R11277 VPWR.n4246 VPWR 0.03175
R11278 VPWR.n4245 VPWR 0.03175
R11279 VPWR VPWR.n7754 0.03175
R11280 VPWR.n7755 VPWR 0.03175
R11281 VPWR.n7808 VPWR 0.03175
R11282 VPWR VPWR.n6056 0.03175
R11283 VPWR.n6107 VPWR 0.03175
R11284 VPWR.n6106 VPWR 0.03175
R11285 VPWR.n6080 VPWR 0.03175
R11286 VPWR.n9199 VPWR 0.03175
R11287 VPWR.n9198 VPWR 0.03175
R11288 VPWR.n9169 VPWR 0.03175
R11289 VPWR.n9143 VPWR 0.03175
R11290 VPWR.n92 VPWR 0.03175
R11291 VPWR.n3264 VPWR 0.03175
R11292 VPWR.n3212 VPWR 0.03175
R11293 VPWR.n3875 VPWR 0.03175
R11294 VPWR.n3087 VPWR 0.03175
R11295 VPWR.n3073 VPWR 0.03175
R11296 VPWR VPWR.n3882 0.03175
R11297 VPWR VPWR.n4004 0.03175
R11298 VPWR VPWR.n4071 0.03175
R11299 VPWR VPWR.n4090 0.03175
R11300 VPWR.n7512 VPWR 0.03175
R11301 VPWR.n7504 VPWR 0.03175
R11302 VPWR.n7459 VPWR 0.03175
R11303 VPWR.n7395 VPWR 0.03175
R11304 VPWR.n7378 VPWR 0.03175
R11305 VPWR.n7361 VPWR 0.03175
R11306 VPWR VPWR.n7068 0.03175
R11307 VPWR.n7069 VPWR 0.03175
R11308 VPWR VPWR.n7129 0.03175
R11309 VPWR.n7174 VPWR 0.03175
R11310 VPWR.n9270 VPWR.n9269 0.0309054
R11311 VPWR.n7875 VPWR.n7874 0.0309054
R11312 VPWR.n8856 VPWR.n8855 0.0309054
R11313 VPWR.n5921 VPWR.n5920 0.0309054
R11314 VPWR.n8725 VPWR.n8724 0.0309054
R11315 VPWR.n5882 VPWR.n5881 0.0309054
R11316 VPWR.n5767 VPWR.n5766 0.0309054
R11317 VPWR.n769 VPWR.n768 0.0309054
R11318 VPWR.n400 VPWR.n399 0.0309054
R11319 VPWR.n5374 VPWR.n5373 0.0309054
R11320 VPWR.n4627 VPWR.n4626 0.0309054
R11321 VPWR.n520 VPWR.n519 0.0309054
R11322 VPWR.n4911 VPWR.n4910 0.0309054
R11323 VPWR.n1820 VPWR.n1819 0.0309054
R11324 VPWR.n2104 VPWR.n2103 0.0309054
R11325 VPWR.n6003 VPWR.n6002 0.0309054
R11326 VPWR.n3429 VPWR.n3428 0.0309054
R11327 VPWR.n6960 VPWR.n6959 0.0309054
R11328 VPWR.n3925 VPWR.n3924 0.0309054
R11329 VPWR.n7321 VPWR.n7320 0.0309054
R11330 VPWR.n7146 VPWR.n7145 0.0309054
R11331 VPWR VPWR.n8422 0.0296459
R11332 VPWR.n929 VPWR 0.0296459
R11333 VPWR VPWR.n1751 0.0291458
R11334 VPWR VPWR.n2587 0.0291458
R11335 VPWR VPWR.n2668 0.0291458
R11336 VPWR.n6872 VPWR.n6869 0.0284688
R11337 VPWR.n6794 VPWR.n6791 0.0284688
R11338 VPWR.n1642 VPWR.n1641 0.0284688
R11339 VPWR.n2546 VPWR.n2545 0.0284688
R11340 VPWR.n2393 VPWR.n2392 0.0284688
R11341 VPWR.n7737 VPWR.n6131 0.0284688
R11342 VPWR.n7609 VPWR.n7608 0.0284688
R11343 VPWR.n8965 VPWR.n200 0.0282455
R11344 VPWR.n8704 VPWR.n8703 0.0282455
R11345 VPWR.n4869 VPWR.n4868 0.0282455
R11346 VPWR.n4566 VPWR.n4565 0.0282455
R11347 VPWR.n4231 VPWR.n4230 0.0282455
R11348 VPWR.n9128 VPWR.n139 0.0282455
R11349 VPWR.n3328 VPWR.n3327 0.0282455
R11350 VPWR.n7262 VPWR.n7132 0.0282455
R11351 VPWR.n4169 VPWR.n4168 0.0282455
R11352 VPWR.n7898 VPWR.n7897 0.0278438
R11353 VPWR.n7956 VPWR 0.0278438
R11354 VPWR.n9082 VPWR 0.0278438
R11355 VPWR VPWR.n8831 0.0278438
R11356 VPWR.n8534 VPWR 0.0278438
R11357 VPWR VPWR.n8791 0.0278438
R11358 VPWR.n3962 VPWR 0.0278438
R11359 VPWR VPWR.n0 0.0278438
R11360 VPWR.n3352 VPWR.n3351 0.027527
R11361 VPWR.n9109 VPWR.n9108 0.027527
R11362 VPWR.n6148 VPWR.n6147 0.027527
R11363 VPWR.n8935 VPWR.n335 0.027527
R11364 VPWR.n6844 VPWR.n6843 0.027527
R11365 VPWR.n8815 VPWR.n8814 0.027527
R11366 VPWR.n6565 VPWR.n6564 0.027527
R11367 VPWR.n5845 VPWR.n380 0.027527
R11368 VPWR.n690 VPWR.n688 0.027527
R11369 VPWR.n5726 VPWR.n5725 0.027527
R11370 VPWR.n1245 VPWR.n1244 0.027527
R11371 VPWR.n4615 VPWR.n4614 0.027527
R11372 VPWR.n573 VPWR.n572 0.027527
R11373 VPWR.n4899 VPWR.n4898 0.027527
R11374 VPWR.n2523 VPWR.n2521 0.027527
R11375 VPWR.n2206 VPWR.n2205 0.027527
R11376 VPWR.n7625 VPWR.n7624 0.027527
R11377 VPWR.n6912 VPWR.n6911 0.027527
R11378 VPWR.n4193 VPWR.n4192 0.027527
R11379 VPWR.n7235 VPWR.n7234 0.027527
R11380 VPWR.n7986 VPWR.n7985 0.0265417
R11381 VPWR.n9089 VPWR.n9088 0.0265417
R11382 VPWR.n6678 VPWR.n6677 0.0265417
R11383 VPWR.n8379 VPWR.n8378 0.0265417
R11384 VPWR.n893 VPWR.n892 0.0265417
R11385 VPWR VPWR.n5831 0.0265417
R11386 VPWR.n1407 VPWR.n1406 0.0265417
R11387 VPWR.n5560 VPWR.n5559 0.0265417
R11388 VPWR.n1746 VPWR.n1745 0.0265417
R11389 VPWR.n4659 VPWR.n4658 0.0265417
R11390 VPWR.n5175 VPWR.n5174 0.0265417
R11391 VPWR.n1878 VPWR.n1877 0.0265417
R11392 VPWR.n2659 VPWR.n2658 0.0265417
R11393 VPWR.n4385 VPWR.n4384 0.0265417
R11394 VPWR.n3558 VPWR.n3557 0.0265417
R11395 VPWR.n4282 VPWR.n4281 0.0265417
R11396 VPWR.n7835 VPWR.n7834 0.0265417
R11397 VPWR.n9225 VPWR.n9224 0.0265417
R11398 VPWR.n3851 VPWR.n3850 0.0265417
R11399 VPWR.n3955 VPWR.n3954 0.0265417
R11400 VPWR.n7437 VPWR.n7436 0.0265417
R11401 VPWR.n7335 VPWR.n7334 0.0265417
R11402 VPWR.n5205 VPWR.n5204 0.0260562
R11403 VPWR.n4878 VPWR.n4877 0.0260562
R11404 VPWR.n3140 VPWR.n3139 0.0258378
R11405 VPWR.n154 VPWR.n153 0.0258378
R11406 VPWR.n9249 VPWR.n9248 0.0258378
R11407 VPWR.n9228 VPWR.n9227 0.0258378
R11408 VPWR.n9218 VPWR.n9217 0.0258378
R11409 VPWR.n28 VPWR.n27 0.0258378
R11410 VPWR.n303 VPWR.n302 0.0258378
R11411 VPWR.n9081 VPWR.n9080 0.0258378
R11412 VPWR.n191 VPWR.n190 0.0258378
R11413 VPWR.n7885 VPWR.n7884 0.0258378
R11414 VPWR.n7888 VPWR.n7887 0.0258378
R11415 VPWR.n5973 VPWR.n5972 0.0258378
R11416 VPWR.n7981 VPWR.n7980 0.0258378
R11417 VPWR.n332 VPWR.n331 0.0258378
R11418 VPWR.n8097 VPWR.n8096 0.0258378
R11419 VPWR.n8100 VPWR.n8099 0.0258378
R11420 VPWR.n8352 VPWR.n8351 0.0258378
R11421 VPWR.n8355 VPWR.n8354 0.0258378
R11422 VPWR.n5892 VPWR.n5891 0.0258378
R11423 VPWR.n5897 VPWR.n5896 0.0258378
R11424 VPWR.n8811 VPWR.n8810 0.0258378
R11425 VPWR.n8533 VPWR.n8532 0.0258378
R11426 VPWR.n8586 VPWR.n8585 0.0258378
R11427 VPWR.n6425 VPWR.n6424 0.0258378
R11428 VPWR.n6427 VPWR.n6426 0.0258378
R11429 VPWR.n8365 VPWR.n8364 0.0258378
R11430 VPWR.n8396 VPWR.n8395 0.0258378
R11431 VPWR.n5756 VPWR.n5754 0.0258378
R11432 VPWR.n741 VPWR.n740 0.0258378
R11433 VPWR.n1104 VPWR.n1103 0.0258378
R11434 VPWR.n778 VPWR.n777 0.0258378
R11435 VPWR.n781 VPWR.n780 0.0258378
R11436 VPWR.n791 VPWR.n790 0.0258378
R11437 VPWR.n898 VPWR.n897 0.0258378
R11438 VPWR.n5722 VPWR.n5721 0.0258378
R11439 VPWR.n5527 VPWR.n5526 0.0258378
R11440 VPWR.n5530 VPWR.n5529 0.0258378
R11441 VPWR.n5361 VPWR.n5360 0.0258378
R11442 VPWR.n5364 VPWR.n5363 0.0258378
R11443 VPWR.n508 VPWR.n507 0.0258378
R11444 VPWR.n1402 VPWR.n1401 0.0258378
R11445 VPWR.n4611 VPWR.n4610 0.0258378
R11446 VPWR.n5218 VPWR.n5217 0.0258378
R11447 VPWR.n5221 VPWR.n5220 0.0258378
R11448 VPWR.n1754 VPWR.n1753 0.0258378
R11449 VPWR.n1756 VPWR.n1755 0.0258378
R11450 VPWR.n5332 VPWR.n5331 0.0258378
R11451 VPWR.n5337 VPWR.n5336 0.0258378
R11452 VPWR.n4895 VPWR.n4894 0.0258378
R11453 VPWR.n1886 VPWR.n1885 0.0258378
R11454 VPWR.n1876 VPWR.n1875 0.0258378
R11455 VPWR.n2112 VPWR.n2111 0.0258378
R11456 VPWR.n2592 VPWR.n2591 0.0258378
R11457 VPWR.n1810 VPWR.n1809 0.0258378
R11458 VPWR.n5180 VPWR.n5179 0.0258378
R11459 VPWR.n4345 VPWR.n4344 0.0258378
R11460 VPWR.n4348 VPWR.n4347 0.0258378
R11461 VPWR.n4582 VPWR.n4581 0.0258378
R11462 VPWR.n2673 VPWR.n2672 0.0258378
R11463 VPWR.n2038 VPWR.n2037 0.0258378
R11464 VPWR.n2615 VPWR.n2614 0.0258378
R11465 VPWR.n2620 VPWR.n2619 0.0258378
R11466 VPWR.n5979 VPWR.n5978 0.0258378
R11467 VPWR.n5982 VPWR.n5981 0.0258378
R11468 VPWR.n7011 VPWR.n7010 0.0258378
R11469 VPWR.n7016 VPWR.n7015 0.0258378
R11470 VPWR.n4220 VPWR.n2868 0.0258378
R11471 VPWR.n3480 VPWR.n3479 0.0258378
R11472 VPWR.n2771 VPWR.n2770 0.0258378
R11473 VPWR.n2776 VPWR.n2775 0.0258378
R11474 VPWR.n4313 VPWR.n4312 0.0258378
R11475 VPWR.n3114 VPWR.n3113 0.0258378
R11476 VPWR.n3782 VPWR.n3781 0.0258378
R11477 VPWR.n3787 VPWR.n3786 0.0258378
R11478 VPWR.n3100 VPWR.n3099 0.0258378
R11479 VPWR.n3104 VPWR.n3103 0.0258378
R11480 VPWR.n6993 VPWR.n6992 0.0258378
R11481 VPWR.n6996 VPWR.n6995 0.0258378
R11482 VPWR.n6981 VPWR.n6980 0.0258378
R11483 VPWR.n6986 VPWR.n6985 0.0258378
R11484 VPWR.n3024 VPWR.n3023 0.0258378
R11485 VPWR.n3965 VPWR.n3964 0.0258378
R11486 VPWR.n3001 VPWR.n3000 0.0258378
R11487 VPWR.n3978 VPWR.n3977 0.0258378
R11488 VPWR.n7310 VPWR.n7309 0.0258378
R11489 VPWR.n7303 VPWR.n7302 0.0258378
R11490 VPWR.n7301 VPWR.n7300 0.0258378
R11491 VPWR.n9287 VPWR.n9286 0.0258378
R11492 VPWR.n6133 VPWR.n6132 0.0258378
R11493 VPWR.n6936 VPWR.n6935 0.0258378
R11494 VPWR.n7249 VPWR.n7248 0.0258378
R11495 VPWR.n7983 VPWR.n5971 0.0252396
R11496 VPWR.n7962 VPWR.n7961 0.0252396
R11497 VPWR.n9091 VPWR.n188 0.0252396
R11498 VPWR.n6675 VPWR.n6674 0.0252396
R11499 VPWR.n6660 VPWR.n6659 0.0252396
R11500 VPWR.n8252 VPWR.n8251 0.0252396
R11501 VPWR.n8239 VPWR.n8238 0.0252396
R11502 VPWR.n8393 VPWR.n8392 0.0252396
R11503 VPWR.n8384 VPWR.n8383 0.0252396
R11504 VPWR.n8566 VPWR.n8565 0.0252396
R11505 VPWR VPWR.n8515 0.0252396
R11506 VPWR.n901 VPWR.n900 0.0252396
R11507 VPWR.n906 VPWR.n766 0.0252396
R11508 VPWR.n1085 VPWR.n1084 0.0252396
R11509 VPWR.n1404 VPWR.n1398 0.0252396
R11510 VPWR.n5397 VPWR.n5396 0.0252396
R11511 VPWR.n5510 VPWR.n5509 0.0252396
R11512 VPWR.n5557 VPWR.n474 0.0252396
R11513 VPWR.n1743 VPWR.n1742 0.0252396
R11514 VPWR.n1729 VPWR.n1728 0.0252396
R11515 VPWR.n5250 VPWR.n5249 0.0252396
R11516 VPWR.n5172 VPWR.n5171 0.0252396
R11517 VPWR.n5163 VPWR.n5162 0.0252396
R11518 VPWR.n5082 VPWR.n5081 0.0252396
R11519 VPWR.n5068 VPWR.n5067 0.0252396
R11520 VPWR.n2656 VPWR.n2655 0.0252396
R11521 VPWR.n2642 VPWR.n2641 0.0252396
R11522 VPWR.n4366 VPWR.n4365 0.0252396
R11523 VPWR.n4382 VPWR.n4381 0.0252396
R11524 VPWR.n3561 VPWR.n3560 0.0252396
R11525 VPWR.n3570 VPWR.n3569 0.0252396
R11526 VPWR.n4299 VPWR.n4298 0.0252396
R11527 VPWR.n4285 VPWR.n4284 0.0252396
R11528 VPWR.n7838 VPWR.n7837 0.0252396
R11529 VPWR.n7852 VPWR.n7851 0.0252396
R11530 VPWR.n9263 VPWR.n9262 0.0252396
R11531 VPWR.n9252 VPWR.n9251 0.0252396
R11532 VPWR.n3848 VPWR.n3847 0.0252396
R11533 VPWR.n3834 VPWR.n3833 0.0252396
R11534 VPWR.n3942 VPWR.n3941 0.0252396
R11535 VPWR.n3952 VPWR.n3951 0.0252396
R11536 VPWR.n7434 VPWR.n7433 0.0252396
R11537 VPWR.n7420 VPWR.n7419 0.0252396
R11538 VPWR.n7348 VPWR.n7347 0.0252396
R11539 VPWR.n7338 VPWR.n7337 0.0252396
R11540 VPWR.n3143 VPWR.n3142 0.0241486
R11541 VPWR.n142 VPWR.n141 0.0241486
R11542 VPWR.n9272 VPWR.n9271 0.0241486
R11543 VPWR.n203 VPWR.n202 0.0241486
R11544 VPWR.n8078 VPWR.n8077 0.0241486
R11545 VPWR.n6315 VPWR.n6314 0.0241486
R11546 VPWR.n7896 VPWR.n7876 0.0241486
R11547 VPWR.n343 VPWR.n342 0.0241486
R11548 VPWR.n8089 VPWR.n8088 0.0241486
R11549 VPWR.n6783 VPWR.n6782 0.0241486
R11550 VPWR.n8345 VPWR.n5922 0.0241486
R11551 VPWR.n8695 VPWR.n8694 0.0241486
R11552 VPWR.n8578 VPWR.n8577 0.0241486
R11553 VPWR.n6333 VPWR.n6332 0.0241486
R11554 VPWR.n8418 VPWR.n5883 0.0241486
R11555 VPWR.n392 VPWR.n391 0.0241486
R11556 VPWR.n1096 VPWR.n1095 0.0241486
R11557 VPWR.n585 VPWR.n584 0.0241486
R11558 VPWR.n925 VPWR.n770 0.0241486
R11559 VPWR.n5656 VPWR.n5655 0.0241486
R11560 VPWR.n5519 VPWR.n5518 0.0241486
R11561 VPWR.n1271 VPWR.n1270 0.0241486
R11562 VPWR.n5376 VPWR.n5375 0.0241486
R11563 VPWR.n4873 VPWR.n4872 0.0241486
R11564 VPWR.n5210 VPWR.n5209 0.0241486
R11565 VPWR.n1535 VPWR.n1534 0.0241486
R11566 VPWR.n5325 VPWR.n521 0.0241486
R11567 VPWR.n1968 VPWR.n1967 0.0241486
R11568 VPWR.n1868 VPWR.n1867 0.0241486
R11569 VPWR.n2419 VPWR.n2418 0.0241486
R11570 VPWR.n1827 VPWR.n1821 0.0241486
R11571 VPWR.n2382 VPWR.n2381 0.0241486
R11572 VPWR.n4357 VPWR.n2734 0.0241486
R11573 VPWR.n4570 VPWR.n4569 0.0241486
R11574 VPWR.n2634 VPWR.n2105 0.0241486
R11575 VPWR.n7857 VPWR.n6004 0.0241486
R11576 VPWR.n2872 VPWR.n2871 0.0241486
R11577 VPWR.n3368 VPWR.n3367 0.0241486
R11578 VPWR.n4305 VPWR.n4304 0.0241486
R11579 VPWR.n3531 VPWR.n3528 0.0241486
R11580 VPWR.n3827 VPWR.n3092 0.0241486
R11581 VPWR.n7027 VPWR.n6961 0.0241486
R11582 VPWR.n3932 VPWR.n3926 0.0241486
R11583 VPWR.n7323 VPWR.n7322 0.0241486
R11584 VPWR.n6136 VPWR.n6135 0.0241486
R11585 VPWR.n6939 VPWR.n6938 0.0241486
R11586 VPWR.n4174 VPWR.n4173 0.0241486
R11587 VPWR.n7134 VPWR.n7133 0.0241486
R11588 VPWR.n8895 VPWR 0.0239375
R11589 VPWR.n8771 VPWR 0.0239375
R11590 VPWR VPWR.n862 0.0239375
R11591 VPWR.n964 VPWR 0.0239375
R11592 VPWR.n1031 VPWR 0.0239375
R11593 VPWR VPWR.n1075 0.0239375
R11594 VPWR.n5493 VPWR 0.0239375
R11595 VPWR.n5620 VPWR 0.0239375
R11596 VPWR.n5291 VPWR 0.0239375
R11597 VPWR.n5281 VPWR 0.0239375
R11598 VPWR.n4656 VPWR 0.0239375
R11599 VPWR.n4753 VPWR 0.0239375
R11600 VPWR.n4822 VPWR 0.0239375
R11601 VPWR.n5117 VPWR 0.0239375
R11602 VPWR.n5086 VPWR 0.0239375
R11603 VPWR.n1909 VPWR 0.0239375
R11604 VPWR.n2725 VPWR 0.0239375
R11605 VPWR.n91 VPWR 0.0239375
R11606 VPWR VPWR.n6183 0.0226354
R11607 VPWR VPWR.n6184 0.0226354
R11608 VPWR.n6299 VPWR 0.0226354
R11609 VPWR.n6294 VPWR 0.0226354
R11610 VPWR.n6283 VPWR 0.0226354
R11611 VPWR.n6273 VPWR 0.0226354
R11612 VPWR.n6266 VPWR 0.0226354
R11613 VPWR.n6241 VPWR 0.0226354
R11614 VPWR.n7955 VPWR 0.0226354
R11615 VPWR.n7923 VPWR 0.0226354
R11616 VPWR.n7910 VPWR 0.0226354
R11617 VPWR.n8043 VPWR 0.0226354
R11618 VPWR.n9052 VPWR 0.0226354
R11619 VPWR.n8983 VPWR 0.0226354
R11620 VPWR VPWR.n9017 0.0226354
R11621 VPWR.n9028 VPWR 0.0226354
R11622 VPWR.n9045 VPWR 0.0226354
R11623 VPWR.n8974 VPWR 0.0226354
R11624 VPWR.n246 VPWR 0.0226354
R11625 VPWR.n232 VPWR 0.0226354
R11626 VPWR.n229 VPWR 0.0226354
R11627 VPWR.n228 VPWR 0.0226354
R11628 VPWR.n6598 VPWR 0.0226354
R11629 VPWR VPWR.n6613 0.0226354
R11630 VPWR.n6615 VPWR 0.0226354
R11631 VPWR.n6767 VPWR 0.0226354
R11632 VPWR.n6742 VPWR 0.0226354
R11633 VPWR.n6727 VPWR 0.0226354
R11634 VPWR.n6697 VPWR 0.0226354
R11635 VPWR.n6691 VPWR 0.0226354
R11636 VPWR.n8333 VPWR 0.0226354
R11637 VPWR.n8318 VPWR 0.0226354
R11638 VPWR.n8307 VPWR 0.0226354
R11639 VPWR.n8303 VPWR 0.0226354
R11640 VPWR.n8294 VPWR 0.0226354
R11641 VPWR.n8284 VPWR 0.0226354
R11642 VPWR.n8262 VPWR 0.0226354
R11643 VPWR.n8258 VPWR 0.0226354
R11644 VPWR.n8189 VPWR 0.0226354
R11645 VPWR.n8127 VPWR 0.0226354
R11646 VPWR VPWR.n8144 0.0226354
R11647 VPWR VPWR.n8166 0.0226354
R11648 VPWR.n8167 VPWR 0.0226354
R11649 VPWR VPWR.n8181 0.0226354
R11650 VPWR.n8906 VPWR 0.0226354
R11651 VPWR.n8900 VPWR 0.0226354
R11652 VPWR.n8889 VPWR 0.0226354
R11653 VPWR.n8883 VPWR 0.0226354
R11654 VPWR VPWR.n6513 0.0226354
R11655 VPWR.n6514 VPWR 0.0226354
R11656 VPWR VPWR.n6518 0.0226354
R11657 VPWR VPWR.n6532 0.0226354
R11658 VPWR.n6451 VPWR 0.0226354
R11659 VPWR.n6374 VPWR 0.0226354
R11660 VPWR.n6383 VPWR 0.0226354
R11661 VPWR.n6410 VPWR 0.0226354
R11662 VPWR VPWR.n8426 0.0226354
R11663 VPWR.n8428 VPWR 0.0226354
R11664 VPWR.n8436 VPWR 0.0226354
R11665 VPWR VPWR.n8460 0.0226354
R11666 VPWR VPWR.n8463 0.0226354
R11667 VPWR VPWR.n8487 0.0226354
R11668 VPWR VPWR.n8488 0.0226354
R11669 VPWR.n8489 VPWR 0.0226354
R11670 VPWR.n8657 VPWR 0.0226354
R11671 VPWR.n8644 VPWR 0.0226354
R11672 VPWR.n8641 VPWR 0.0226354
R11673 VPWR.n8634 VPWR 0.0226354
R11674 VPWR VPWR.n8681 0.0226354
R11675 VPWR.n8722 VPWR 0.0226354
R11676 VPWR.n8774 VPWR 0.0226354
R11677 VPWR.n8761 VPWR 0.0226354
R11678 VPWR.n8760 VPWR 0.0226354
R11679 VPWR.n8749 VPWR 0.0226354
R11680 VPWR.n620 VPWR 0.0226354
R11681 VPWR VPWR.n623 0.0226354
R11682 VPWR.n624 VPWR 0.0226354
R11683 VPWR.n1210 VPWR 0.0226354
R11684 VPWR VPWR.n838 0.0226354
R11685 VPWR.n839 VPWR 0.0226354
R11686 VPWR VPWR.n847 0.0226354
R11687 VPWR.n855 VPWR 0.0226354
R11688 VPWR.n958 VPWR 0.0226354
R11689 VPWR VPWR.n990 0.0226354
R11690 VPWR.n1021 VPWR 0.0226354
R11691 VPWR VPWR.n1030 0.0226354
R11692 VPWR.n1117 VPWR 0.0226354
R11693 VPWR VPWR.n1128 0.0226354
R11694 VPWR.n1129 VPWR 0.0226354
R11695 VPWR VPWR.n1135 0.0226354
R11696 VPWR.n1136 VPWR 0.0226354
R11697 VPWR VPWR.n1194 0.0226354
R11698 VPWR.n5743 VPWR 0.0226354
R11699 VPWR.n5828 VPWR 0.0226354
R11700 VPWR.n5806 VPWR 0.0226354
R11701 VPWR.n5799 VPWR 0.0226354
R11702 VPWR.n5794 VPWR 0.0226354
R11703 VPWR VPWR.n1299 0.0226354
R11704 VPWR.n1302 VPWR 0.0226354
R11705 VPWR.n1318 VPWR 0.0226354
R11706 VPWR.n1517 VPWR 0.0226354
R11707 VPWR.n1501 VPWR 0.0226354
R11708 VPWR.n1490 VPWR 0.0226354
R11709 VPWR.n1459 VPWR 0.0226354
R11710 VPWR.n1451 VPWR 0.0226354
R11711 VPWR.n1442 VPWR 0.0226354
R11712 VPWR.n1437 VPWR 0.0226354
R11713 VPWR VPWR.n5444 0.0226354
R11714 VPWR.n5445 VPWR 0.0226354
R11715 VPWR VPWR.n5465 0.0226354
R11716 VPWR VPWR.n5483 0.0226354
R11717 VPWR.n5484 VPWR 0.0226354
R11718 VPWR VPWR.n5492 0.0226354
R11719 VPWR VPWR.n5589 0.0226354
R11720 VPWR.n5603 VPWR 0.0226354
R11721 VPWR.n461 VPWR 0.0226354
R11722 VPWR VPWR.n5608 0.0226354
R11723 VPWR VPWR.n5619 0.0226354
R11724 VPWR.n5635 VPWR 0.0226354
R11725 VPWR VPWR.n5639 0.0226354
R11726 VPWR.n5641 VPWR 0.0226354
R11727 VPWR.n447 VPWR 0.0226354
R11728 VPWR.n442 VPWR 0.0226354
R11729 VPWR.n428 VPWR 0.0226354
R11730 VPWR.n424 VPWR 0.0226354
R11731 VPWR.n421 VPWR 0.0226354
R11732 VPWR.n1568 VPWR 0.0226354
R11733 VPWR.n1544 VPWR 0.0226354
R11734 VPWR VPWR.n1659 0.0226354
R11735 VPWR.n1667 VPWR 0.0226354
R11736 VPWR.n1682 VPWR 0.0226354
R11737 VPWR.n1701 VPWR 0.0226354
R11738 VPWR VPWR.n1712 0.0226354
R11739 VPWR.n1713 VPWR 0.0226354
R11740 VPWR.n1720 VPWR 0.0226354
R11741 VPWR.n1774 VPWR 0.0226354
R11742 VPWR.n1773 VPWR 0.0226354
R11743 VPWR.n5294 VPWR 0.0226354
R11744 VPWR.n5284 VPWR 0.0226354
R11745 VPWR.n5277 VPWR 0.0226354
R11746 VPWR VPWR.n4686 0.0226354
R11747 VPWR.n4759 VPWR 0.0226354
R11748 VPWR.n4754 VPWR 0.0226354
R11749 VPWR.n4748 VPWR 0.0226354
R11750 VPWR.n4723 VPWR 0.0226354
R11751 VPWR.n4769 VPWR 0.0226354
R11752 VPWR.n4837 VPWR 0.0226354
R11753 VPWR.n4829 VPWR 0.0226354
R11754 VPWR.n4826 VPWR 0.0226354
R11755 VPWR.n4816 VPWR 0.0226354
R11756 VPWR.n4803 VPWR 0.0226354
R11757 VPWR VPWR.n2442 0.0226354
R11758 VPWR.n2443 VPWR 0.0226354
R11759 VPWR VPWR.n2451 0.0226354
R11760 VPWR VPWR.n2462 0.0226354
R11761 VPWR VPWR.n2463 0.0226354
R11762 VPWR.n2464 VPWR 0.0226354
R11763 VPWR.n2471 VPWR 0.0226354
R11764 VPWR.n2547 VPWR 0.0226354
R11765 VPWR VPWR.n2557 0.0226354
R11766 VPWR.n2558 VPWR 0.0226354
R11767 VPWR.n2154 VPWR 0.0226354
R11768 VPWR.n2141 VPWR 0.0226354
R11769 VPWR.n2139 VPWR 0.0226354
R11770 VPWR.n2132 VPWR 0.0226354
R11771 VPWR.n2125 VPWR 0.0226354
R11772 VPWR.n2575 VPWR 0.0226354
R11773 VPWR.n5143 VPWR 0.0226354
R11774 VPWR.n5139 VPWR 0.0226354
R11775 VPWR.n5113 VPWR 0.0226354
R11776 VPWR.n5102 VPWR 0.0226354
R11777 VPWR.n5090 VPWR 0.0226354
R11778 VPWR.n1914 VPWR 0.0226354
R11779 VPWR VPWR.n1957 0.0226354
R11780 VPWR.n5010 VPWR 0.0226354
R11781 VPWR.n5008 VPWR 0.0226354
R11782 VPWR.n4957 VPWR 0.0226354
R11783 VPWR.n4938 VPWR 0.0226354
R11784 VPWR.n4931 VPWR 0.0226354
R11785 VPWR.n2228 VPWR 0.0226354
R11786 VPWR.n2238 VPWR 0.0226354
R11787 VPWR VPWR.n2254 0.0226354
R11788 VPWR VPWR.n2300 0.0226354
R11789 VPWR.n2371 VPWR 0.0226354
R11790 VPWR.n2338 VPWR 0.0226354
R11791 VPWR.n2331 VPWR 0.0226354
R11792 VPWR.n2328 VPWR 0.0226354
R11793 VPWR.n2321 VPWR 0.0226354
R11794 VPWR.n2320 VPWR 0.0226354
R11795 VPWR.n2061 VPWR 0.0226354
R11796 VPWR.n2050 VPWR 0.0226354
R11797 VPWR.n2046 VPWR 0.0226354
R11798 VPWR VPWR.n2697 0.0226354
R11799 VPWR VPWR.n2724 0.0226354
R11800 VPWR VPWR.n4425 0.0226354
R11801 VPWR VPWR.n4426 0.0226354
R11802 VPWR VPWR.n4453 0.0226354
R11803 VPWR.n4462 VPWR 0.0226354
R11804 VPWR VPWR.n4475 0.0226354
R11805 VPWR.n4539 VPWR 0.0226354
R11806 VPWR.n4535 VPWR 0.0226354
R11807 VPWR.n4520 VPWR 0.0226354
R11808 VPWR.n4517 VPWR 0.0226354
R11809 VPWR.n4512 VPWR 0.0226354
R11810 VPWR.n4510 VPWR 0.0226354
R11811 VPWR.n4505 VPWR 0.0226354
R11812 VPWR.n3394 VPWR 0.0226354
R11813 VPWR VPWR.n3408 0.0226354
R11814 VPWR VPWR.n3409 0.0226354
R11815 VPWR.n3410 VPWR 0.0226354
R11816 VPWR VPWR.n3414 0.0226354
R11817 VPWR.n3746 VPWR 0.0226354
R11818 VPWR.n3743 VPWR 0.0226354
R11819 VPWR.n3735 VPWR 0.0226354
R11820 VPWR.n3721 VPWR 0.0226354
R11821 VPWR.n3693 VPWR 0.0226354
R11822 VPWR.n3689 VPWR 0.0226354
R11823 VPWR.n3577 VPWR 0.0226354
R11824 VPWR.n3593 VPWR 0.0226354
R11825 VPWR VPWR.n3610 0.0226354
R11826 VPWR.n3611 VPWR 0.0226354
R11827 VPWR VPWR.n3623 0.0226354
R11828 VPWR.n3664 VPWR 0.0226354
R11829 VPWR.n4252 VPWR 0.0226354
R11830 VPWR VPWR.n2820 0.0226354
R11831 VPWR VPWR.n2830 0.0226354
R11832 VPWR.n2831 VPWR 0.0226354
R11833 VPWR VPWR.n2864 0.0226354
R11834 VPWR.n2959 VPWR 0.0226354
R11835 VPWR.n2923 VPWR 0.0226354
R11836 VPWR.n2899 VPWR 0.0226354
R11837 VPWR VPWR.n7662 0.0226354
R11838 VPWR.n7663 VPWR 0.0226354
R11839 VPWR VPWR.n7753 0.0226354
R11840 VPWR.n7781 VPWR 0.0226354
R11841 VPWR.n7789 VPWR 0.0226354
R11842 VPWR VPWR.n7807 0.0226354
R11843 VPWR.n7814 VPWR 0.0226354
R11844 VPWR.n6026 VPWR 0.0226354
R11845 VPWR.n6033 VPWR 0.0226354
R11846 VPWR VPWR.n6041 0.0226354
R11847 VPWR.n6049 VPWR 0.0226354
R11848 VPWR.n6053 VPWR 0.0226354
R11849 VPWR.n6090 VPWR 0.0226354
R11850 VPWR.n6084 VPWR 0.0226354
R11851 VPWR.n6077 VPWR 0.0226354
R11852 VPWR.n6073 VPWR 0.0226354
R11853 VPWR.n6072 VPWR 0.0226354
R11854 VPWR VPWR.n33 0.0226354
R11855 VPWR.n9188 VPWR 0.0226354
R11856 VPWR.n9181 VPWR 0.0226354
R11857 VPWR.n9171 VPWR 0.0226354
R11858 VPWR.n9163 VPWR 0.0226354
R11859 VPWR.n9158 VPWR 0.0226354
R11860 VPWR.n9155 VPWR 0.0226354
R11861 VPWR.n9146 VPWR 0.0226354
R11862 VPWR.n9130 VPWR 0.0226354
R11863 VPWR.n108 VPWR 0.0226354
R11864 VPWR.n97 VPWR 0.0226354
R11865 VPWR.n86 VPWR 0.0226354
R11866 VPWR.n85 VPWR 0.0226354
R11867 VPWR.n3256 VPWR 0.0226354
R11868 VPWR VPWR.n3262 0.0226354
R11869 VPWR VPWR.n3263 0.0226354
R11870 VPWR VPWR.n3281 0.0226354
R11871 VPWR.n3284 VPWR 0.0226354
R11872 VPWR.n3217 VPWR 0.0226354
R11873 VPWR.n3207 VPWR 0.0226354
R11874 VPWR.n3186 VPWR 0.0226354
R11875 VPWR.n3176 VPWR 0.0226354
R11876 VPWR.n3173 VPWR 0.0226354
R11877 VPWR.n3171 VPWR 0.0226354
R11878 VPWR.n3170 VPWR 0.0226354
R11879 VPWR.n3162 VPWR 0.0226354
R11880 VPWR.n3874 VPWR 0.0226354
R11881 VPWR.n3090 VPWR 0.0226354
R11882 VPWR.n3081 VPWR 0.0226354
R11883 VPWR.n3075 VPWR 0.0226354
R11884 VPWR.n3074 VPWR 0.0226354
R11885 VPWR.n3884 VPWR 0.0226354
R11886 VPWR VPWR.n3905 0.0226354
R11887 VPWR VPWR.n4003 0.0226354
R11888 VPWR VPWR.n4026 0.0226354
R11889 VPWR.n4051 VPWR 0.0226354
R11890 VPWR VPWR.n4057 0.0226354
R11891 VPWR.n4058 VPWR 0.0226354
R11892 VPWR VPWR.n4062 0.0226354
R11893 VPWR VPWR.n4070 0.0226354
R11894 VPWR.n4072 VPWR 0.0226354
R11895 VPWR.n4129 VPWR 0.0226354
R11896 VPWR.n4125 VPWR 0.0226354
R11897 VPWR.n4124 VPWR 0.0226354
R11898 VPWR VPWR.n4099 0.0226354
R11899 VPWR.n7547 VPWR 0.0226354
R11900 VPWR VPWR.n7565 0.0226354
R11901 VPWR.n7568 VPWR 0.0226354
R11902 VPWR.n7515 VPWR 0.0226354
R11903 VPWR.n7507 VPWR 0.0226354
R11904 VPWR.n7500 VPWR 0.0226354
R11905 VPWR.n7475 VPWR 0.0226354
R11906 VPWR.n7472 VPWR 0.0226354
R11907 VPWR.n7403 VPWR 0.0226354
R11908 VPWR.n7400 VPWR 0.0226354
R11909 VPWR.n7374 VPWR 0.0226354
R11910 VPWR.n7364 VPWR 0.0226354
R11911 VPWR.n7357 VPWR 0.0226354
R11912 VPWR.n7352 VPWR 0.0226354
R11913 VPWR VPWR.n7067 0.0226354
R11914 VPWR.n7079 VPWR 0.0226354
R11915 VPWR.n7105 VPWR 0.0226354
R11916 VPWR.n7112 VPWR 0.0226354
R11917 VPWR VPWR.n7128 0.0226354
R11918 VPWR.n7193 VPWR 0.0226354
R11919 VPWR.n7185 VPWR 0.0226354
R11920 VPWR.n7171 VPWR 0.0226354
R11921 VPWR.n7161 VPWR 0.0226354
R11922 VPWR.n3347 VPWR.n3346 0.0224595
R11923 VPWR.n3354 VPWR.n3353 0.0224595
R11924 VPWR.n3335 VPWR.n3334 0.0224595
R11925 VPWR.n3338 VPWR.n3337 0.0224595
R11926 VPWR.n160 VPWR.n156 0.0224595
R11927 VPWR.n159 VPWR.n158 0.0224595
R11928 VPWR.n9111 VPWR.n9110 0.0224595
R11929 VPWR.n9114 VPWR.n9113 0.0224595
R11930 VPWR.n9248 VPWR.n9247 0.0224595
R11931 VPWR.n9245 VPWR.n9230 0.0224595
R11932 VPWR.n310 VPWR.n305 0.0224595
R11933 VPWR.n309 VPWR.n308 0.0224595
R11934 VPWR.n8948 VPWR.n8947 0.0224595
R11935 VPWR.n8951 VPWR.n8950 0.0224595
R11936 VPWR.n170 VPWR.n169 0.0224595
R11937 VPWR.n175 VPWR.n174 0.0224595
R11938 VPWR.n6143 VPWR.n6142 0.0224595
R11939 VPWR.n6150 VPWR.n6149 0.0224595
R11940 VPWR.n6153 VPWR.n6152 0.0224595
R11941 VPWR.n6885 VPWR.n6884 0.0224595
R11942 VPWR.n7977 VPWR.n5975 0.0224595
R11943 VPWR.n7980 VPWR.n7979 0.0224595
R11944 VPWR.n8939 VPWR.n334 0.0224595
R11945 VPWR.n8938 VPWR.n8937 0.0224595
R11946 VPWR.n320 VPWR.n319 0.0224595
R11947 VPWR.n8235 VPWR.n8234 0.0224595
R11948 VPWR.n8232 VPWR.n5955 0.0224595
R11949 VPWR.n6839 VPWR.n6838 0.0224595
R11950 VPWR.n6846 VPWR.n6845 0.0224595
R11951 VPWR.n6849 VPWR.n6848 0.0224595
R11952 VPWR.n6853 VPWR.n6852 0.0224595
R11953 VPWR.n5900 VPWR.n5894 0.0224595
R11954 VPWR.n5898 VPWR.n5897 0.0224595
R11955 VPWR.n8819 VPWR.n8813 0.0224595
R11956 VPWR.n8818 VPWR.n8817 0.0224595
R11957 VPWR.n8720 VPWR.n348 0.0224595
R11958 VPWR.n8526 VPWR.n8525 0.0224595
R11959 VPWR.n8542 VPWR.n8541 0.0224595
R11960 VPWR.n6324 VPWR.n6323 0.0224595
R11961 VPWR.n6567 VPWR.n6566 0.0224595
R11962 VPWR.n6570 VPWR.n6569 0.0224595
R11963 VPWR.n6574 VPWR.n6573 0.0224595
R11964 VPWR.n8399 VPWR.n8367 0.0224595
R11965 VPWR.n8397 VPWR.n8396 0.0224595
R11966 VPWR.n5849 VPWR.n379 0.0224595
R11967 VPWR.n5848 VPWR.n5847 0.0224595
R11968 VPWR.n368 VPWR.n367 0.0224595
R11969 VPWR.n1052 VPWR.n1051 0.0224595
R11970 VPWR.n1061 VPWR.n1060 0.0224595
R11971 VPWR.n670 VPWR.n669 0.0224595
R11972 VPWR.n687 VPWR.n686 0.0224595
R11973 VPWR.n590 VPWR.n589 0.0224595
R11974 VPWR.n701 VPWR.n591 0.0224595
R11975 VPWR.n794 VPWR.n793 0.0224595
R11976 VPWR.n897 VPWR.n896 0.0224595
R11977 VPWR.n5730 VPWR.n5724 0.0224595
R11978 VPWR.n5729 VPWR.n5728 0.0224595
R11979 VPWR.n5710 VPWR.n5709 0.0224595
R11980 VPWR.n5538 VPWR.n5537 0.0224595
R11981 VPWR.n5543 VPWR.n5542 0.0224595
R11982 VPWR.n1240 VPWR.n1239 0.0224595
R11983 VPWR.n1247 VPWR.n1246 0.0224595
R11984 VPWR.n1250 VPWR.n1249 0.0224595
R11985 VPWR.n1254 VPWR.n1253 0.0224595
R11986 VPWR.n511 VPWR.n510 0.0224595
R11987 VPWR.n1401 VPWR.n1400 0.0224595
R11988 VPWR.n4619 VPWR.n4613 0.0224595
R11989 VPWR.n4618 VPWR.n4617 0.0224595
R11990 VPWR.n4599 VPWR.n4598 0.0224595
R11991 VPWR.n5229 VPWR.n5228 0.0224595
R11992 VPWR.n5234 VPWR.n5233 0.0224595
R11993 VPWR.n568 VPWR.n567 0.0224595
R11994 VPWR.n575 VPWR.n574 0.0224595
R11995 VPWR.n563 VPWR.n562 0.0224595
R11996 VPWR.n1628 VPWR.n1625 0.0224595
R11997 VPWR.n5340 VPWR.n5334 0.0224595
R11998 VPWR.n5338 VPWR.n5337 0.0224595
R11999 VPWR.n4903 VPWR.n4897 0.0224595
R12000 VPWR.n4902 VPWR.n4901 0.0224595
R12001 VPWR.n4883 VPWR.n4882 0.0224595
R12002 VPWR.n5048 VPWR.n5047 0.0224595
R12003 VPWR.n5053 VPWR.n5052 0.0224595
R12004 VPWR.n2489 VPWR.n2487 0.0224595
R12005 VPWR.n2520 VPWR.n2519 0.0224595
R12006 VPWR.n2506 VPWR.n2505 0.0224595
R12007 VPWR.n2510 VPWR.n2509 0.0224595
R12008 VPWR.n5183 VPWR.n5177 0.0224595
R12009 VPWR.n5181 VPWR.n5180 0.0224595
R12010 VPWR.n2201 VPWR.n2200 0.0224595
R12011 VPWR.n2208 VPWR.n2207 0.0224595
R12012 VPWR.n2211 VPWR.n2210 0.0224595
R12013 VPWR.n2401 VPWR.n2400 0.0224595
R12014 VPWR.n2751 VPWR.n2750 0.0224595
R12015 VPWR.n2756 VPWR.n2755 0.0224595
R12016 VPWR.n4589 VPWR.n4584 0.0224595
R12017 VPWR.n4588 VPWR.n4587 0.0224595
R12018 VPWR.n1983 VPWR.n1982 0.0224595
R12019 VPWR.n1986 VPWR.n1985 0.0224595
R12020 VPWR.n2623 VPWR.n2617 0.0224595
R12021 VPWR.n2621 VPWR.n2620 0.0224595
R12022 VPWR.n7019 VPWR.n7013 0.0224595
R12023 VPWR.n7017 VPWR.n7016 0.0224595
R12024 VPWR.n4218 VPWR.n4217 0.0224595
R12025 VPWR.n2944 VPWR.n2869 0.0224595
R12026 VPWR.n2957 VPWR.n2956 0.0224595
R12027 VPWR.n2952 VPWR.n2951 0.0224595
R12028 VPWR.n3431 VPWR.n3430 0.0224595
R12029 VPWR.n3436 VPWR.n3435 0.0224595
R12030 VPWR.n3470 VPWR.n3469 0.0224595
R12031 VPWR.n3482 VPWR.n3477 0.0224595
R12032 VPWR.n2772 VPWR.n2771 0.0224595
R12033 VPWR.n2779 VPWR.n2778 0.0224595
R12034 VPWR.n3790 VPWR.n3784 0.0224595
R12035 VPWR.n3788 VPWR.n3787 0.0224595
R12036 VPWR.n3802 VPWR.n3798 0.0224595
R12037 VPWR.n3800 VPWR.n3799 0.0224595
R12038 VPWR.n6989 VPWR.n6983 0.0224595
R12039 VPWR.n6987 VPWR.n6986 0.0224595
R12040 VPWR.n3025 VPWR.n3024 0.0224595
R12041 VPWR.n3968 VPWR.n3967 0.0224595
R12042 VPWR.n7309 VPWR.n7308 0.0224595
R12043 VPWR.n7306 VPWR.n7305 0.0224595
R12044 VPWR.n7620 VPWR.n7619 0.0224595
R12045 VPWR.n7627 VPWR.n7626 0.0224595
R12046 VPWR.n7698 VPWR.n7697 0.0224595
R12047 VPWR.n7704 VPWR.n7702 0.0224595
R12048 VPWR.n6907 VPWR.n6906 0.0224595
R12049 VPWR.n6914 VPWR.n6913 0.0224595
R12050 VPWR.n6926 VPWR.n6925 0.0224595
R12051 VPWR.n6929 VPWR.n6928 0.0224595
R12052 VPWR.n4184 VPWR.n4181 0.0224595
R12053 VPWR.n4183 VPWR.n4182 0.0224595
R12054 VPWR.n4195 VPWR.n4194 0.0224595
R12055 VPWR.n4198 VPWR.n4197 0.0224595
R12056 VPWR.n7254 VPWR.n7251 0.0224595
R12057 VPWR.n7253 VPWR.n7252 0.0224595
R12058 VPWR.n7237 VPWR.n7236 0.0224595
R12059 VPWR.n7144 VPWR.n7143 0.0224595
R12060 VPWR.n1079 VPWR.n1078 0.0217384
R12061 VPWR.n6216 VPWR.n6215 0.0213333
R12062 VPWR.n278 VPWR.n277 0.0213333
R12063 VPWR.n6815 VPWR.n6814 0.0213333
R12064 VPWR.n8934 VPWR.n8933 0.0213333
R12065 VPWR.n6555 VPWR 0.0213333
R12066 VPWR VPWR.n6554 0.0213333
R12067 VPWR.n6563 VPWR.n6328 0.0213333
R12068 VPWR.n6406 VPWR 0.0213333
R12069 VPWR.n5878 VPWR 0.0213333
R12070 VPWR.n611 VPWR 0.0213333
R12071 VPWR.n691 VPWR.n667 0.0213333
R12072 VPWR.n5844 VPWR.n5843 0.0213333
R12073 VPWR.n5800 VPWR 0.0213333
R12074 VPWR VPWR.n1317 0.0213333
R12075 VPWR.n1346 VPWR.n1345 0.0213333
R12076 VPWR.n5411 VPWR 0.0213333
R12077 VPWR.n5431 VPWR 0.0213333
R12078 VPWR.n5689 VPWR.n5688 0.0213333
R12079 VPWR.n1596 VPWR.n1595 0.0213333
R12080 VPWR.n1708 VPWR 0.0213333
R12081 VPWR.n5321 VPWR 0.0213333
R12082 VPWR.n5319 VPWR 0.0213333
R12083 VPWR.n5297 VPWR 0.0213333
R12084 VPWR.n4683 VPWR 0.0213333
R12085 VPWR.n4853 VPWR.n4852 0.0213333
R12086 VPWR.n2484 VPWR 0.0213333
R12087 VPWR VPWR.n2483 0.0213333
R12088 VPWR.n2524 VPWR.n2191 0.0213333
R12089 VPWR.n5156 VPWR 0.0213333
R12090 VPWR.n5126 VPWR 0.0213333
R12091 VPWR.n5024 VPWR 0.0213333
R12092 VPWR VPWR.n1912 0.0213333
R12093 VPWR.n4976 VPWR.n4975 0.0213333
R12094 VPWR.n2286 VPWR.n2285 0.0213333
R12095 VPWR.n4449 VPWR 0.0213333
R12096 VPWR.n4554 VPWR.n4553 0.0213333
R12097 VPWR.n3459 VPWR.n3458 0.0213333
R12098 VPWR.n7715 VPWR.n7714 0.0213333
R12099 VPWR.n126 VPWR.n125 0.0213333
R12100 VPWR.n3307 VPWR.n3306 0.0213333
R12101 VPWR.n4149 VPWR.n4148 0.0213333
R12102 VPWR.n7588 VPWR.n7587 0.0213333
R12103 VPWR VPWR.n7111 0.0213333
R12104 VPWR.n7213 VPWR.n7212 0.0213333
R12105 VPWR.n150 VPWR.n149 0.0202124
R12106 VPWR.n9119 VPWR.n9118 0.0202124
R12107 VPWR.n301 VPWR.n300 0.0202124
R12108 VPWR.n8956 VPWR.n8955 0.0202124
R12109 VPWR.n168 VPWR.n167 0.0202124
R12110 VPWR.n9074 VPWR.n9073 0.0202124
R12111 VPWR.n6140 VPWR.n6139 0.0202124
R12112 VPWR.n6317 VPWR.n6316 0.0202124
R12113 VPWR.n5977 VPWR.n5976 0.0202124
R12114 VPWR.n7878 VPWR.n7877 0.0202124
R12115 VPWR.n318 VPWR.n317 0.0202124
R12116 VPWR.n8858 VPWR.n8857 0.0202124
R12117 VPWR.n5957 VPWR.n5956 0.0202124
R12118 VPWR.n8093 VPWR.n8092 0.0202124
R12119 VPWR.n6836 VPWR.n6835 0.0202124
R12120 VPWR.n6785 VPWR.n6784 0.0202124
R12121 VPWR.n5890 VPWR.n5889 0.0202124
R12122 VPWR.n5917 VPWR.n5916 0.0202124
R12123 VPWR.n347 VPWR.n346 0.0202124
R12124 VPWR.n8727 VPWR.n8726 0.0202124
R12125 VPWR.n8522 VPWR.n8521 0.0202124
R12126 VPWR.n359 VPWR.n358 0.0202124
R12127 VPWR.n6321 VPWR.n6320 0.0202124
R12128 VPWR.n6335 VPWR.n6334 0.0202124
R12129 VPWR.n8363 VPWR.n8362 0.0202124
R12130 VPWR.n5885 VPWR.n5884 0.0202124
R12131 VPWR.n366 VPWR.n365 0.0202124
R12132 VPWR.n5769 VPWR.n5768 0.0202124
R12133 VPWR.n1049 VPWR.n1048 0.0202124
R12134 VPWR.n744 VPWR.n743 0.0202124
R12135 VPWR.n674 VPWR.n673 0.0202124
R12136 VPWR.n579 VPWR.n578 0.0202124
R12137 VPWR.n789 VPWR.n788 0.0202124
R12138 VPWR.n772 VPWR.n771 0.0202124
R12139 VPWR.n5708 VPWR.n5707 0.0202124
R12140 VPWR.n396 VPWR.n395 0.0202124
R12141 VPWR.n481 VPWR.n480 0.0202124
R12142 VPWR.n5523 VPWR.n5522 0.0202124
R12143 VPWR.n1237 VPWR.n1236 0.0202124
R12144 VPWR.n1265 VPWR.n1264 0.0202124
R12145 VPWR.n506 VPWR.n505 0.0202124
R12146 VPWR.n5370 VPWR.n5369 0.0202124
R12147 VPWR.n4597 VPWR.n4596 0.0202124
R12148 VPWR.n4623 VPWR.n4622 0.0202124
R12149 VPWR.n1802 VPWR.n1801 0.0202124
R12150 VPWR.n5214 VPWR.n5213 0.0202124
R12151 VPWR.n565 VPWR.n564 0.0202124
R12152 VPWR.n1529 VPWR.n1528 0.0202124
R12153 VPWR.n5330 VPWR.n5329 0.0202124
R12154 VPWR.n516 VPWR.n515 0.0202124
R12155 VPWR.n4881 VPWR.n4880 0.0202124
R12156 VPWR.n4907 VPWR.n4906 0.0202124
R12157 VPWR.n1863 VPWR.n1862 0.0202124
R12158 VPWR.n1872 VPWR.n1871 0.0202124
R12159 VPWR.n2194 VPWR.n2193 0.0202124
R12160 VPWR.n2413 VPWR.n2412 0.0202124
R12161 VPWR.n1808 VPWR.n1807 0.0202124
R12162 VPWR.n1823 VPWR.n1822 0.0202124
R12163 VPWR.n2198 VPWR.n2197 0.0202124
R12164 VPWR.n2384 VPWR.n2383 0.0202124
R12165 VPWR.n2738 VPWR.n2737 0.0202124
R12166 VPWR.n4340 VPWR.n4339 0.0202124
R12167 VPWR.n4577 VPWR.n4576 0.0202124
R12168 VPWR.n1980 VPWR.n1979 0.0202124
R12169 VPWR.n2600 VPWR.n2599 0.0202124
R12170 VPWR.n2107 VPWR.n2106 0.0202124
R12171 VPWR.n7004 VPWR.n7003 0.0202124
R12172 VPWR.n5997 VPWR.n5996 0.0202124
R12173 VPWR.n2878 VPWR.n2877 0.0202124
R12174 VPWR.n3440 VPWR.n3439 0.0202124
R12175 VPWR.n3475 VPWR.n3474 0.0202124
R12176 VPWR.n4321 VPWR.n4320 0.0202124
R12177 VPWR.n2768 VPWR.n2767 0.0202124
R12178 VPWR.n3777 VPWR.n3776 0.0202124
R12179 VPWR.n3097 VPWR.n3096 0.0202124
R12180 VPWR.n3821 VPWR.n3820 0.0202124
R12181 VPWR.n6974 VPWR.n6973 0.0202124
R12182 VPWR.n6970 VPWR.n6969 0.0202124
R12183 VPWR.n3929 VPWR.n3928 0.0202124
R12184 VPWR.n3970 VPWR.n3969 0.0202124
R12185 VPWR.n7 VPWR.n6 0.0202124
R12186 VPWR.n16 VPWR.n15 0.0202124
R12187 VPWR.n9274 VPWR.n9273 0.0202124
R12188 VPWR.n7617 VPWR.n7616 0.0202124
R12189 VPWR.n7700 VPWR.n7699 0.0202124
R12190 VPWR.n6899 VPWR.n6898 0.0202124
R12191 VPWR.n6932 VPWR.n6931 0.0202124
R12192 VPWR.n3137 VPWR.n3136 0.0202124
R12193 VPWR.n2987 VPWR.n2986 0.0202124
R12194 VPWR.n4203 VPWR.n4202 0.0202124
R12195 VPWR.n7257 VPWR.n7256 0.0202124
R12196 VPWR.n7232 VPWR.n7231 0.0202124
R12197 VPWR.n6881 VPWR.n6880 0.0200312
R12198 VPWR.n8004 VPWR.n8003 0.0200312
R12199 VPWR.n7999 VPWR.n7998 0.0200312
R12200 VPWR.n7985 VPWR.n7984 0.0200312
R12201 VPWR VPWR.n8062 0.0200312
R12202 VPWR.n9090 VPWR.n9089 0.0200312
R12203 VPWR.n9070 VPWR.n9069 0.0200312
R12204 VPWR.n267 VPWR.n266 0.0200312
R12205 VPWR.n6803 VPWR.n6802 0.0200312
R12206 VPWR.n6687 VPWR.n6686 0.0200312
R12207 VPWR.n6682 VPWR.n6681 0.0200312
R12208 VPWR.n6677 VPWR.n6676 0.0200312
R12209 VPWR.n8206 VPWR.n8205 0.0200312
R12210 VPWR.n8843 VPWR.n8842 0.0200312
R12211 VPWR.n6476 VPWR.n6475 0.0200312
R12212 VPWR.n6436 VPWR.n6435 0.0200312
R12213 VPWR.n8370 VPWR.n8369 0.0200312
R12214 VPWR.n8380 VPWR.n8379 0.0200312
R12215 VPWR.n8381 VPWR 0.0200312
R12216 VPWR.n8590 VPWR.n8589 0.0200312
R12217 VPWR.n8708 VPWR.n8707 0.0200312
R12218 VPWR VPWR.n8721 0.0200312
R12219 VPWR.n705 VPWR.n704 0.0200312
R12220 VPWR.n876 VPWR.n875 0.0200312
R12221 VPWR.n881 VPWR.n880 0.0200312
R12222 VPWR.n894 VPWR.n893 0.0200312
R12223 VPWR.n930 VPWR 0.0200312
R12224 VPWR.n736 VPWR.n735 0.0200312
R12225 VPWR.n1108 VPWR.n1107 0.0200312
R12226 VPWR.n5757 VPWR.n5753 0.0200312
R12227 VPWR.n1357 VPWR.n1356 0.0200312
R12228 VPWR.n1421 VPWR.n1419 0.0200312
R12229 VPWR.n1415 VPWR.n1414 0.0200312
R12230 VPWR.n1406 VPWR.n1405 0.0200312
R12231 VPWR.n5559 VPWR.n5558 0.0200312
R12232 VPWR.n5566 VPWR.n5565 0.0200312
R12233 VPWR.n5572 VPWR.n5570 0.0200312
R12234 VPWR.n5677 VPWR.n5676 0.0200312
R12235 VPWR.n1632 VPWR.n1631 0.0200312
R12236 VPWR.n1765 VPWR.n1764 0.0200312
R12237 VPWR.n1750 VPWR.n1749 0.0200312
R12238 VPWR.n1745 VPWR.n1744 0.0200312
R12239 VPWR.n4658 VPWR.n4657 0.0200312
R12240 VPWR.n4665 VPWR.n4664 0.0200312
R12241 VPWR.n4670 VPWR.n4669 0.0200312
R12242 VPWR.n4864 VPWR.n4863 0.0200312
R12243 VPWR.n2536 VPWR.n2535 0.0200312
R12244 VPWR.n2584 VPWR.n2583 0.0200312
R12245 VPWR.n2586 VPWR.n2585 0.0200312
R12246 VPWR.n5174 VPWR.n5173 0.0200312
R12247 VPWR.n1877 VPWR.n1856 0.0200312
R12248 VPWR.n1883 VPWR.n1882 0.0200312
R12249 VPWR.n5039 VPWR.n5038 0.0200312
R12250 VPWR.n4968 VPWR.n4967 0.0200312
R12251 VPWR.n2397 VPWR.n2396 0.0200312
R12252 VPWR.n2667 VPWR.n2666 0.0200312
R12253 VPWR.n2658 VPWR.n2657 0.0200312
R12254 VPWR.n4384 VPWR.n4383 0.0200312
R12255 VPWR.n4390 VPWR.n4389 0.0200312
R12256 VPWR.n4396 VPWR.n4394 0.0200312
R12257 VPWR.n4562 VPWR.n4561 0.0200312
R12258 VPWR.n3486 VPWR.n3485 0.0200312
R12259 VPWR.n3548 VPWR.n3547 0.0200312
R12260 VPWR.n3553 VPWR.n3552 0.0200312
R12261 VPWR.n3559 VPWR.n3558 0.0200312
R12262 VPWR.n4283 VPWR.n4282 0.0200312
R12263 VPWR.n4276 VPWR.n4275 0.0200312
R12264 VPWR.n4271 VPWR.n4270 0.0200312
R12265 VPWR.n4222 VPWR.n4221 0.0200312
R12266 VPWR VPWR.n2958 0.0200312
R12267 VPWR.n7695 VPWR.n7694 0.0200312
R12268 VPWR.n7824 VPWR.n7823 0.0200312
R12269 VPWR.n7829 VPWR.n7828 0.0200312
R12270 VPWR.n7836 VPWR.n7835 0.0200312
R12271 VPWR.n9226 VPWR.n9225 0.0200312
R12272 VPWR.n9220 VPWR.n9219 0.0200312
R12273 VPWR.n9212 VPWR.n9211 0.0200312
R12274 VPWR.n136 VPWR.n135 0.0200312
R12275 VPWR.n3318 VPWR.n3317 0.0200312
R12276 VPWR.n3864 VPWR.n3862 0.0200312
R12277 VPWR.n3858 VPWR.n3857 0.0200312
R12278 VPWR.n3850 VPWR.n3849 0.0200312
R12279 VPWR.n3954 VPWR.n3953 0.0200312
R12280 VPWR.n3983 VPWR.n3981 0.0200312
R12281 VPWR.n4160 VPWR.n4159 0.0200312
R12282 VPWR.n7599 VPWR.n7598 0.0200312
R12283 VPWR.n7448 VPWR.n7446 0.0200312
R12284 VPWR.n7442 VPWR.n7441 0.0200312
R12285 VPWR.n7436 VPWR.n7435 0.0200312
R12286 VPWR.n7336 VPWR.n7335 0.0200312
R12287 VPWR.n7051 VPWR.n1 0.0200312
R12288 VPWR.n7202 VPWR.n7201 0.0200312
R12289 VPWR.n3348 VPWR.n3347 0.0190811
R12290 VPWR.n3355 VPWR.n3349 0.0190811
R12291 VPWR.n9117 VPWR.n9116 0.0190811
R12292 VPWR.n9115 VPWR.n9114 0.0190811
R12293 VPWR.n8954 VPWR.n8953 0.0190811
R12294 VPWR.n8952 VPWR.n8951 0.0190811
R12295 VPWR.n185 VPWR.n184 0.0190811
R12296 VPWR.n6144 VPWR.n6143 0.0190811
R12297 VPWR.n6151 VPWR.n6145 0.0190811
R12298 VPWR.n7967 VPWR.n7867 0.0190811
R12299 VPWR.n324 VPWR.n323 0.0190811
R12300 VPWR.n322 VPWR.n321 0.0190811
R12301 VPWR.n8217 VPWR.n8216 0.0190811
R12302 VPWR.n6840 VPWR.n6839 0.0190811
R12303 VPWR.n6847 VPWR.n6841 0.0190811
R12304 VPWR.n5905 VPWR.n5904 0.0190811
R12305 VPWR.n8803 VPWR.n8802 0.0190811
R12306 VPWR.n8801 VPWR.n349 0.0190811
R12307 VPWR.n8519 VPWR.n8518 0.0190811
R12308 VPWR.n6325 VPWR.n6324 0.0190811
R12309 VPWR.n6568 VPWR.n6326 0.0190811
R12310 VPWR.n8404 VPWR.n8403 0.0190811
R12311 VPWR.n372 VPWR.n371 0.0190811
R12312 VPWR.n370 VPWR.n369 0.0190811
R12313 VPWR.n1046 VPWR.n1045 0.0190811
R12314 VPWR.n671 VPWR.n670 0.0190811
R12315 VPWR.n685 VPWR.n672 0.0190811
R12316 VPWR.n911 VPWR.n798 0.0190811
R12317 VPWR.n5714 VPWR.n5713 0.0190811
R12318 VPWR.n5712 VPWR.n5711 0.0190811
R12319 VPWR.n478 VPWR.n477 0.0190811
R12320 VPWR.n1241 VPWR.n1240 0.0190811
R12321 VPWR.n1248 VPWR.n1242 0.0190811
R12322 VPWR.n5391 VPWR.n5390 0.0190811
R12323 VPWR.n4603 VPWR.n4602 0.0190811
R12324 VPWR.n4601 VPWR.n4600 0.0190811
R12325 VPWR.n5244 VPWR.n1799 0.0190811
R12326 VPWR.n569 VPWR.n568 0.0190811
R12327 VPWR.n576 VPWR.n570 0.0190811
R12328 VPWR.n5345 VPWR.n5344 0.0190811
R12329 VPWR.n4887 VPWR.n4886 0.0190811
R12330 VPWR.n4885 VPWR.n4884 0.0190811
R12331 VPWR.n1860 VPWR.n1859 0.0190811
R12332 VPWR.n2489 VPWR.n2488 0.0190811
R12333 VPWR.n2518 VPWR.n2192 0.0190811
R12334 VPWR.n5188 VPWR.n5187 0.0190811
R12335 VPWR.n2202 VPWR.n2201 0.0190811
R12336 VPWR.n2209 VPWR.n2203 0.0190811
R12337 VPWR.n2742 VPWR.n2741 0.0190811
R12338 VPWR.n1989 VPWR.n1988 0.0190811
R12339 VPWR.n1987 VPWR.n1986 0.0190811
R12340 VPWR.n2605 VPWR.n2604 0.0190811
R12341 VPWR.n2955 VPWR.n2954 0.0190811
R12342 VPWR.n2953 VPWR.n2952 0.0190811
R12343 VPWR.n3432 VPWR.n3431 0.0190811
R12344 VPWR.n3437 VPWR.n3433 0.0190811
R12345 VPWR.n4328 VPWR.n4327 0.0190811
R12346 VPWR.n3769 VPWR.n3768 0.0190811
R12347 VPWR.n3817 VPWR.n3816 0.0190811
R12348 VPWR.n3010 VPWR.n3009 0.0190811
R12349 VPWR.n7318 VPWR.n7317 0.0190811
R12350 VPWR.n7621 VPWR.n7620 0.0190811
R12351 VPWR.n7628 VPWR.n7622 0.0190811
R12352 VPWR.n6908 VPWR.n6907 0.0190811
R12353 VPWR.n6915 VPWR.n6909 0.0190811
R12354 VPWR.n4201 VPWR.n4200 0.0190811
R12355 VPWR.n4199 VPWR.n4198 0.0190811
R12356 VPWR.n7240 VPWR.n7239 0.0190811
R12357 VPWR.n7987 VPWR.n7986 0.0187292
R12358 VPWR.n9088 VPWR.n9087 0.0187292
R12359 VPWR.n192 VPWR 0.0187292
R12360 VPWR.n294 VPWR.n288 0.0187292
R12361 VPWR.n6679 VPWR.n6678 0.0187292
R12362 VPWR.n8102 VPWR.n8101 0.0187292
R12363 VPWR.n8835 VPWR.n336 0.0187292
R12364 VPWR.n8923 VPWR.n8922 0.0187292
R12365 VPWR.n8540 VPWR.n8530 0.0187292
R12366 VPWR VPWR.n356 0.0187292
R12367 VPWR.n8795 VPWR.n8793 0.0187292
R12368 VPWR.n892 VPWR.n891 0.0187292
R12369 VPWR.n1059 VPWR.n1056 0.0187292
R12370 VPWR.n733 VPWR 0.0187292
R12371 VPWR.n5746 VPWR.n381 0.0187292
R12372 VPWR.n5835 VPWR.n5833 0.0187292
R12373 VPWR.n1367 VPWR.n1366 0.0187292
R12374 VPWR.n1408 VPWR.n1407 0.0187292
R12375 VPWR.n5561 VPWR.n5560 0.0187292
R12376 VPWR.n5669 VPWR.n5667 0.0187292
R12377 VPWR.n5700 VPWR.n5698 0.0187292
R12378 VPWR.n1747 VPWR.n1746 0.0187292
R12379 VPWR.n4660 VPWR.n4659 0.0187292
R12380 VPWR.n4845 VPWR.n4844 0.0187292
R12381 VPWR.n1879 VPWR.n1878 0.0187292
R12382 VPWR.n1887 VPWR 0.0187292
R12383 VPWR.n5001 VPWR.n5000 0.0187292
R12384 VPWR.n2660 VPWR.n2659 0.0187292
R12385 VPWR.n4386 VPWR.n4385 0.0187292
R12386 VPWR.n4542 VPWR.n4541 0.0187292
R12387 VPWR.n3751 VPWR.n3494 0.0187292
R12388 VPWR.n3557 VPWR.n3556 0.0187292
R12389 VPWR.n4281 VPWR.n4280 0.0187292
R12390 VPWR.n2965 VPWR.n2964 0.0187292
R12391 VPWR.n7834 VPWR.n7833 0.0187292
R12392 VPWR.n9224 VPWR.n9223 0.0187292
R12393 VPWR.n29 VPWR 0.0187292
R12394 VPWR.n116 VPWR.n115 0.0187292
R12395 VPWR.n3852 VPWR.n3851 0.0187292
R12396 VPWR.n3956 VPWR.n3955 0.0187292
R12397 VPWR VPWR.n2999 0.0187292
R12398 VPWR.n4139 VPWR.n4138 0.0187292
R12399 VPWR.n7438 VPWR.n7437 0.0187292
R12400 VPWR.n7334 VPWR.n7333 0.0187292
R12401 VPWR VPWR.n9290 0.0187292
R12402 VPWR.n7225 VPWR.n7223 0.0187292
R12403 VPWR VPWR.n7194 0.0185211
R12404 VPWR VPWR.n258 0.0185211
R12405 VPWR.n8917 VPWR 0.0185211
R12406 VPWR.n8789 VPWR 0.0185211
R12407 VPWR.n5829 VPWR 0.0185211
R12408 VPWR.n6208 VPWR.n6207 0.0174271
R12409 VPWR.n6211 VPWR.n6210 0.0174271
R12410 VPWR.n286 VPWR.n282 0.0174271
R12411 VPWR.n6826 VPWR.n6824 0.0174271
R12412 VPWR.n6822 VPWR.n6819 0.0174271
R12413 VPWR VPWR.n340 0.0174271
R12414 VPWR.n8929 VPWR.n8928 0.0174271
R12415 VPWR.n6552 VPWR.n6551 0.0174271
R12416 VPWR.n6558 VPWR.n6557 0.0174271
R12417 VPWR.n8799 VPWR.n8798 0.0174271
R12418 VPWR.n657 VPWR.n656 0.0174271
R12419 VPWR.n663 VPWR.n662 0.0174271
R12420 VPWR VPWR.n389 0.0174271
R12421 VPWR.n5839 VPWR.n5838 0.0174271
R12422 VPWR.n1337 VPWR.n1335 0.0174271
R12423 VPWR.n1341 VPWR.n1340 0.0174271
R12424 VPWR.n5665 VPWR 0.0174271
R12425 VPWR.n5695 VPWR.n5693 0.0174271
R12426 VPWR.n1608 VPWR.n1607 0.0174271
R12427 VPWR.n1605 VPWR.n1600 0.0174271
R12428 VPWR.n1752 VPWR 0.0174271
R12429 VPWR.n4848 VPWR.n4847 0.0174271
R12430 VPWR.n2495 VPWR.n2494 0.0174271
R12431 VPWR.n2492 VPWR 0.0174271
R12432 VPWR.n2588 VPWR 0.0174271
R12433 VPWR.n5176 VPWR 0.0174271
R12434 VPWR.n4998 VPWR 0.0174271
R12435 VPWR.n4981 VPWR.n4980 0.0174271
R12436 VPWR.n2281 VPWR.n2280 0.0174271
R12437 VPWR.n2669 VPWR 0.0174271
R12438 VPWR.n4549 VPWR.n4548 0.0174271
R12439 VPWR.n3448 VPWR.n3447 0.0174271
R12440 VPWR.n3454 VPWR.n3453 0.0174271
R12441 VPWR.n2962 VPWR.n2961 0.0174271
R12442 VPWR.n7723 VPWR.n7722 0.0174271
R12443 VPWR.n7720 VPWR.n7719 0.0174271
R12444 VPWR.n9206 VPWR 0.0174271
R12445 VPWR.n121 VPWR.n120 0.0174271
R12446 VPWR.n3296 VPWR.n3294 0.0174271
R12447 VPWR.n3302 VPWR.n3301 0.0174271
R12448 VPWR.n4144 VPWR.n4143 0.0174271
R12449 VPWR.n7579 VPWR.n7577 0.0174271
R12450 VPWR.n7583 VPWR.n7582 0.0174271
R12451 VPWR.n7221 VPWR.n7217 0.0174271
R12452 VPWR.n6672 VPWR.n6665 0.0173937
R12453 VPWR.n8390 VPWR.n8389 0.0173937
R12454 VPWR.n3351 VPWR.n3350 0.0173919
R12455 VPWR.n9235 VPWR.n9234 0.0173919
R12456 VPWR.n307 VPWR.n306 0.0173919
R12457 VPWR.n9095 VPWR.n9094 0.0173919
R12458 VPWR.n6147 VPWR.n6146 0.0173919
R12459 VPWR.n7866 VPWR.n7865 0.0173919
R12460 VPWR.n8936 VPWR.n8935 0.0173919
R12461 VPWR.n8223 VPWR.n8222 0.0173919
R12462 VPWR.n6843 VPWR.n6842 0.0173919
R12463 VPWR.n5903 VPWR.n5902 0.0173919
R12464 VPWR.n8816 VPWR.n8815 0.0173919
R12465 VPWR.n8552 VPWR.n8551 0.0173919
R12466 VPWR.n6564 VPWR.n6327 0.0173919
R12467 VPWR.n8402 VPWR.n8401 0.0173919
R12468 VPWR.n5846 VPWR.n5845 0.0173919
R12469 VPWR.n1071 VPWR.n1070 0.0173919
R12470 VPWR.n690 VPWR.n689 0.0173919
R12471 VPWR.n797 VPWR.n796 0.0173919
R12472 VPWR.n5727 VPWR.n5726 0.0173919
R12473 VPWR.n5553 VPWR.n5552 0.0173919
R12474 VPWR.n1244 VPWR.n1243 0.0173919
R12475 VPWR.n504 VPWR.n503 0.0173919
R12476 VPWR.n4616 VPWR.n4615 0.0173919
R12477 VPWR.n4649 VPWR.n1800 0.0173919
R12478 VPWR.n572 VPWR.n571 0.0173919
R12479 VPWR.n5343 VPWR.n5342 0.0173919
R12480 VPWR.n4900 VPWR.n4899 0.0173919
R12481 VPWR.n5063 VPWR.n5062 0.0173919
R12482 VPWR.n2523 VPWR.n2522 0.0173919
R12483 VPWR.n5186 VPWR.n5185 0.0173919
R12484 VPWR.n2205 VPWR.n2204 0.0173919
R12485 VPWR.n2748 VPWR.n2747 0.0173919
R12486 VPWR.n4586 VPWR.n4585 0.0173919
R12487 VPWR.n2603 VPWR.n2602 0.0173919
R12488 VPWR.n5991 VPWR.n5990 0.0173919
R12489 VPWR.n2946 VPWR.n2945 0.0173919
R12490 VPWR.n3468 VPWR.n3467 0.0173919
R12491 VPWR.n4332 VPWR.n4331 0.0173919
R12492 VPWR.n3765 VPWR.n3764 0.0173919
R12493 VPWR.n3813 VPWR.n3812 0.0173919
R12494 VPWR.n6964 VPWR.n6963 0.0173919
R12495 VPWR.n3014 VPWR.n3013 0.0173919
R12496 VPWR.n7314 VPWR.n7313 0.0173919
R12497 VPWR.n7624 VPWR.n7623 0.0173919
R12498 VPWR.n6911 VPWR.n6910 0.0173919
R12499 VPWR.n4192 VPWR.n4191 0.0173919
R12500 VPWR.n7234 VPWR.n7233 0.0173919
R12501 VPWR.n5169 VPWR.n5168 0.0172664
R12502 VPWR.n3564 VPWR.n3563 0.0172664
R12503 VPWR.n4564 VPWR.n4563 0.0172634
R12504 VPWR.n138 VPWR.n137 0.0172634
R12505 VPWR VPWR.n653 0.017219
R12506 VPWR.n8706 VPWR.n8705 0.017135
R12507 VPWR.n5002 VPWR.n1965 0.017135
R12508 VPWR.n9257 VPWR.n9256 0.0169468
R12509 VPWR.n9256 VPWR.n9253 0.0169468
R12510 VPWR.n2394 VPWR.n2393 0.0169447
R12511 VPWR.n2395 VPWR.n2394 0.0169447
R12512 VPWR.n707 VPWR.n706 0.0169447
R12513 VPWR.n708 VPWR.n707 0.0169447
R12514 VPWR.n9125 VPWR.n9124 0.0168788
R12515 VPWR.n147 VPWR.n143 0.0168788
R12516 VPWR.n8962 VPWR.n8961 0.0168788
R12517 VPWR.n298 VPWR.n204 0.0168788
R12518 VPWR.n8079 VPWR.n5959 0.0168788
R12519 VPWR.n9077 VPWR.n9075 0.0168788
R12520 VPWR.n6203 VPWR.n6202 0.0168788
R12521 VPWR.n6866 VPWR.n6318 0.0168788
R12522 VPWR.n7891 VPWR.n7883 0.0168788
R12523 VPWR.n7895 VPWR.n7879 0.0168788
R12524 VPWR.n8826 VPWR.n8825 0.0168788
R12525 VPWR.n8861 VPWR.n8859 0.0168788
R12526 VPWR.n8090 VPWR.n8086 0.0168788
R12527 VPWR.n8210 VPWR.n8094 0.0168788
R12528 VPWR.n6832 VPWR.n6831 0.0168788
R12529 VPWR.n6788 VPWR.n6786 0.0168788
R12530 VPWR.n8358 VPWR.n8350 0.0168788
R12531 VPWR.n8346 VPWR.n5918 0.0168788
R12532 VPWR.n8700 VPWR.n8699 0.0168788
R12533 VPWR.n8730 VPWR.n8728 0.0168788
R12534 VPWR.n8579 VPWR.n5859 0.0168788
R12535 VPWR.n8583 VPWR.n360 0.0168788
R12536 VPWR.n6547 VPWR.n6546 0.0168788
R12537 VPWR.n6340 VPWR.n6336 0.0168788
R12538 VPWR.n6431 VPWR.n6430 0.0168788
R12539 VPWR.n8417 VPWR.n5886 0.0168788
R12540 VPWR.n5737 VPWR.n5736 0.0168788
R12541 VPWR.n5772 VPWR.n5770 0.0168788
R12542 VPWR.n1097 VPWR.n749 0.0168788
R12543 VPWR.n1101 VPWR.n745 0.0168788
R12544 VPWR.n650 VPWR.n649 0.0168788
R12545 VPWR.n1232 VPWR.n580 0.0168788
R12546 VPWR.n784 VPWR.n776 0.0168788
R12547 VPWR.n924 VPWR.n773 0.0168788
R12548 VPWR.n5659 VPWR.n5658 0.0168788
R12549 VPWR.n5704 VPWR.n397 0.0168788
R12550 VPWR.n5520 VPWR.n485 0.0168788
R12551 VPWR.n5533 VPWR.n5524 0.0168788
R12552 VPWR.n1330 VPWR.n1329 0.0168788
R12553 VPWR.n1523 VPWR.n1266 0.0168788
R12554 VPWR.n5367 VPWR.n5359 0.0168788
R12555 VPWR.n5377 VPWR.n5371 0.0168788
R12556 VPWR.n4875 VPWR.n4634 0.0168788
R12557 VPWR.n4630 VPWR.n4624 0.0168788
R12558 VPWR.n5211 VPWR.n5207 0.0168788
R12559 VPWR.n5224 VPWR.n5215 0.0168788
R12560 VPWR.n1614 VPWR.n1613 0.0168788
R12561 VPWR.n1537 VPWR.n1530 0.0168788
R12562 VPWR.n1760 VPWR.n1759 0.0168788
R12563 VPWR.n5326 VPWR.n517 0.0168788
R12564 VPWR.n4992 VPWR.n4991 0.0168788
R12565 VPWR.n4987 VPWR.n4908 0.0168788
R12566 VPWR.n1869 VPWR.n1865 0.0168788
R12567 VPWR.n5043 VPWR.n1873 0.0168788
R12568 VPWR.n2501 VPWR.n2500 0.0168788
R12569 VPWR.n2421 VPWR.n2414 0.0168788
R12570 VPWR.n2595 VPWR.n2110 0.0168788
R12571 VPWR.n1826 VPWR.n1824 0.0168788
R12572 VPWR.n2273 VPWR.n2272 0.0168788
R12573 VPWR.n2389 VPWR.n2385 0.0168788
R12574 VPWR.n4356 VPWR.n4355 0.0168788
R12575 VPWR.n4351 VPWR.n4341 0.0168788
R12576 VPWR.n4573 VPWR.n4572 0.0168788
R12577 VPWR.n1974 VPWR.n1970 0.0168788
R12578 VPWR.n2627 VPWR.n2626 0.0168788
R12579 VPWR.n2633 VPWR.n2108 0.0168788
R12580 VPWR.n5986 VPWR.n5985 0.0168788
R12581 VPWR.n7858 VPWR.n5998 0.0168788
R12582 VPWR.n3107 VPWR.n3098 0.0168788
R12583 VPWR.n3826 VPWR.n3093 0.0168788
R12584 VPWR.n7000 VPWR.n6999 0.0168788
R12585 VPWR.n7026 VPWR.n6971 0.0168788
R12586 VPWR.n3931 VPWR.n3930 0.0168788
R12587 VPWR.n3975 VPWR.n3003 0.0168788
R12588 VPWR.n5 VPWR.n4 0.0168788
R12589 VPWR.n9284 VPWR.n17 0.0168788
R12590 VPWR.n9276 VPWR.n9275 0.0168788
R12591 VPWR.n24 VPWR.n22 0.0168788
R12592 VPWR.n7729 VPWR.n7728 0.0168788
R12593 VPWR.n7734 VPWR.n6137 0.0168788
R12594 VPWR.n6922 VPWR.n6921 0.0168788
R12595 VPWR.n7612 VPWR.n6933 0.0168788
R12596 VPWR.n3135 VPWR.n3134 0.0168788
R12597 VPWR.n3331 VPWR.n3138 0.0168788
R12598 VPWR.n4176 VPWR.n2988 0.0168788
R12599 VPWR.n2982 VPWR.n2978 0.0168788
R12600 VPWR.n7259 VPWR.n7258 0.0168788
R12601 VPWR.n7230 VPWR.n7229 0.0168788
R12602 VPWR.n8705 VPWR.n8704 0.0167522
R12603 VPWR.n5002 VPWR.n5001 0.0167522
R12604 VPWR.n5170 VPWR.n5169 0.0166276
R12605 VPWR.n3563 VPWR.n3562 0.0166276
R12606 VPWR.n4565 VPWR.n4564 0.0166244
R12607 VPWR.n139 VPWR.n138 0.0166244
R12608 VPWR.n6673 VPWR.n6672 0.016499
R12609 VPWR.n8391 VPWR.n8390 0.016499
R12610 VPWR VPWR.n6342 0.016125
R12611 VPWR VPWR.n8377 0.016125
R12612 VPWR.n1227 VPWR 0.016125
R12613 VPWR VPWR.n1369 0.016125
R12614 VPWR.n3749 VPWR 0.016125
R12615 VPWR VPWR.n2947 0.016125
R12616 VPWR.n3337 VPWR.n3336 0.0157027
R12617 VPWR.n3141 VPWR.n3140 0.0157027
R12618 VPWR.n3142 VPWR.n3141 0.0157027
R12619 VPWR.n3330 VPWR.n3143 0.0157027
R12620 VPWR.n9126 VPWR.n142 0.0157027
R12621 VPWR.n141 VPWR.n140 0.0157027
R12622 VPWR.n156 VPWR.n155 0.0157027
R12623 VPWR.n158 VPWR.n157 0.0157027
R12624 VPWR.n9271 VPWR.n9270 0.0157027
R12625 VPWR.n8963 VPWR.n203 0.0157027
R12626 VPWR.n202 VPWR.n201 0.0157027
R12627 VPWR.n305 VPWR.n304 0.0157027
R12628 VPWR.n308 VPWR.n307 0.0157027
R12629 VPWR.n8077 VPWR.n5961 0.0157027
R12630 VPWR.n6884 VPWR.n6155 0.0157027
R12631 VPWR.n6313 VPWR.n6312 0.0157027
R12632 VPWR.n6314 VPWR.n6313 0.0157027
R12633 VPWR.n6867 VPWR.n6315 0.0157027
R12634 VPWR.n7876 VPWR.n7875 0.0157027
R12635 VPWR.n8830 VPWR.n8829 0.0157027
R12636 VPWR.n8827 VPWR.n343 0.0157027
R12637 VPWR.n342 VPWR.n341 0.0157027
R12638 VPWR.n334 VPWR.n333 0.0157027
R12639 VPWR.n8937 VPWR.n8936 0.0157027
R12640 VPWR.n8088 VPWR.n8087 0.0157027
R12641 VPWR.n6852 VPWR.n6851 0.0157027
R12642 VPWR.n6781 VPWR.n6780 0.0157027
R12643 VPWR.n6782 VPWR.n6781 0.0157027
R12644 VPWR.n6789 VPWR.n6783 0.0157027
R12645 VPWR.n5922 VPWR.n5921 0.0157027
R12646 VPWR.n8701 VPWR.n8695 0.0157027
R12647 VPWR.n8694 VPWR.n8693 0.0157027
R12648 VPWR.n8813 VPWR.n8812 0.0157027
R12649 VPWR.n8817 VPWR.n8816 0.0157027
R12650 VPWR.n8577 VPWR.n8576 0.0157027
R12651 VPWR.n6573 VPWR.n6572 0.0157027
R12652 VPWR.n6331 VPWR.n6330 0.0157027
R12653 VPWR.n6332 VPWR.n6331 0.0157027
R12654 VPWR.n6341 VPWR.n6333 0.0157027
R12655 VPWR.n6463 VPWR.n6462 0.0157027
R12656 VPWR.n5883 VPWR.n5882 0.0157027
R12657 VPWR.n5741 VPWR.n5740 0.0157027
R12658 VPWR.n5738 VPWR.n392 0.0157027
R12659 VPWR.n391 VPWR.n390 0.0157027
R12660 VPWR.n5755 VPWR.n379 0.0157027
R12661 VPWR.n5847 VPWR.n5846 0.0157027
R12662 VPWR.n1095 VPWR.n1094 0.0157027
R12663 VPWR.n702 VPWR.n701 0.0157027
R12664 VPWR.n583 VPWR.n582 0.0157027
R12665 VPWR.n584 VPWR.n583 0.0157027
R12666 VPWR.n1231 VPWR.n585 0.0157027
R12667 VPWR.n1225 VPWR.n586 0.0157027
R12668 VPWR.n770 VPWR.n769 0.0157027
R12669 VPWR.n5663 VPWR.n5662 0.0157027
R12670 VPWR.n5660 VPWR.n5656 0.0157027
R12671 VPWR.n5655 VPWR.n5654 0.0157027
R12672 VPWR.n5724 VPWR.n5723 0.0157027
R12673 VPWR.n5728 VPWR.n5727 0.0157027
R12674 VPWR.n5518 VPWR.n5517 0.0157027
R12675 VPWR.n1253 VPWR.n1252 0.0157027
R12676 VPWR.n1269 VPWR.n1268 0.0157027
R12677 VPWR.n1270 VPWR.n1269 0.0157027
R12678 VPWR.n1522 VPWR.n1271 0.0157027
R12679 VPWR.n1520 VPWR.n1519 0.0157027
R12680 VPWR.n5375 VPWR.n5374 0.0157027
R12681 VPWR.n4874 VPWR.n4873 0.0157027
R12682 VPWR.n4872 VPWR.n4871 0.0157027
R12683 VPWR.n4613 VPWR.n4612 0.0157027
R12684 VPWR.n4617 VPWR.n4616 0.0157027
R12685 VPWR.n5209 VPWR.n5208 0.0157027
R12686 VPWR.n1628 VPWR.n1627 0.0157027
R12687 VPWR.n1533 VPWR.n1532 0.0157027
R12688 VPWR.n1534 VPWR.n1533 0.0157027
R12689 VPWR.n1536 VPWR.n1535 0.0157027
R12690 VPWR.n521 VPWR.n520 0.0157027
R12691 VPWR.n4996 VPWR.n4995 0.0157027
R12692 VPWR.n4993 VPWR.n1968 0.0157027
R12693 VPWR.n1967 VPWR.n1966 0.0157027
R12694 VPWR.n4897 VPWR.n4896 0.0157027
R12695 VPWR.n4901 VPWR.n4900 0.0157027
R12696 VPWR.n1867 VPWR.n1866 0.0157027
R12697 VPWR.n2509 VPWR.n2508 0.0157027
R12698 VPWR.n2417 VPWR.n2416 0.0157027
R12699 VPWR.n2418 VPWR.n2417 0.0157027
R12700 VPWR.n2420 VPWR.n2419 0.0157027
R12701 VPWR.n1821 VPWR.n1820 0.0157027
R12702 VPWR.n2400 VPWR.n2213 0.0157027
R12703 VPWR.n2380 VPWR.n2379 0.0157027
R12704 VPWR.n2381 VPWR.n2380 0.0157027
R12705 VPWR.n2390 VPWR.n2382 0.0157027
R12706 VPWR.n2734 VPWR.n2733 0.0157027
R12707 VPWR.n4571 VPWR.n4570 0.0157027
R12708 VPWR.n4569 VPWR.n4568 0.0157027
R12709 VPWR.n4584 VPWR.n4583 0.0157027
R12710 VPWR.n4587 VPWR.n4586 0.0157027
R12711 VPWR.n2105 VPWR.n2104 0.0157027
R12712 VPWR.n6004 VPWR.n6003 0.0157027
R12713 VPWR.n2873 VPWR.n2872 0.0157027
R12714 VPWR.n2868 VPWR.n2867 0.0157027
R12715 VPWR.n4219 VPWR.n4218 0.0157027
R12716 VPWR.n2945 VPWR.n2944 0.0157027
R12717 VPWR.n3469 VPWR.n3468 0.0157027
R12718 VPWR.n3482 VPWR.n3481 0.0157027
R12719 VPWR.n3479 VPWR.n3478 0.0157027
R12720 VPWR.n3753 VPWR.n3368 0.0157027
R12721 VPWR.n3747 VPWR.n3369 0.0157027
R12722 VPWR.n4304 VPWR.n4303 0.0157027
R12723 VPWR.n3528 VPWR.n3527 0.0157027
R12724 VPWR.n3092 VPWR.n3091 0.0157027
R12725 VPWR.n6961 VPWR.n6960 0.0157027
R12726 VPWR.n3926 VPWR.n3925 0.0157027
R12727 VPWR.n7322 VPWR.n7321 0.0157027
R12728 VPWR.n7704 VPWR.n7703 0.0157027
R12729 VPWR.n6134 VPWR.n6133 0.0157027
R12730 VPWR.n6135 VPWR.n6134 0.0157027
R12731 VPWR.n7735 VPWR.n6136 0.0157027
R12732 VPWR.n6928 VPWR.n6927 0.0157027
R12733 VPWR.n6937 VPWR.n6936 0.0157027
R12734 VPWR.n6938 VPWR.n6937 0.0157027
R12735 VPWR.n7611 VPWR.n6939 0.0157027
R12736 VPWR.n4175 VPWR.n4174 0.0157027
R12737 VPWR.n4173 VPWR.n4172 0.0157027
R12738 VPWR.n4172 VPWR.n4171 0.0157027
R12739 VPWR.n4181 VPWR.n4180 0.0157027
R12740 VPWR.n7260 VPWR.n7134 0.0157027
R12741 VPWR.n7248 VPWR.n7247 0.0157027
R12742 VPWR.n7251 VPWR.n7250 0.0157027
R12743 VPWR.n2640 VPWR.n2636 0.0153255
R12744 VPWR.n3573 VPWR.n3572 0.0153255
R12745 VPWR.n7855 VPWR.n7854 0.0153255
R12746 VPWR.n7418 VPWR.n7415 0.0153255
R12747 VPWR.n8343 VPWR.n5923 0.0150286
R12748 VPWR.n5400 VPWR.n5399 0.0150286
R12749 VPWR.n5323 VPWR.n524 0.0150286
R12750 VPWR.n5161 VPWR.n5160 0.0150286
R12751 VPWR.n3832 VPWR.n3829 0.0150286
R12752 VPWR.n6212 VPWR.n6211 0.0148229
R12753 VPWR.n7871 VPWR.n7870 0.0148229
R12754 VPWR.n7966 VPWR.n7965 0.0148229
R12755 VPWR.n8073 VPWR.n8072 0.0148229
R12756 VPWR.n282 VPWR.n281 0.0148229
R12757 VPWR.n6819 VPWR.n6818 0.0148229
R12758 VPWR.n6664 VPWR.n6663 0.0148229
R12759 VPWR.n8248 VPWR.n8247 0.0148229
R12760 VPWR VPWR.n8105 0.0148229
R12761 VPWR.n8930 VPWR.n8929 0.0148229
R12762 VPWR.n6557 VPWR.n6556 0.0148229
R12763 VPWR.n8388 VPWR.n8387 0.0148229
R12764 VPWR.n8562 VPWR.n8561 0.0148229
R12765 VPWR.n8719 VPWR 0.0148229
R12766 VPWR.n8800 VPWR.n8799 0.0148229
R12767 VPWR.n664 VPWR.n663 0.0148229
R12768 VPWR.n905 VPWR.n904 0.0148229
R12769 VPWR.n910 VPWR.n909 0.0148229
R12770 VPWR.n1081 VPWR.n1080 0.0148229
R12771 VPWR.n5840 VPWR.n5839 0.0148229
R12772 VPWR.n5833 VPWR 0.0148229
R12773 VPWR.n1342 VPWR.n1341 0.0148229
R12774 VPWR.n1393 VPWR.n1391 0.0148229
R12775 VPWR.n5393 VPWR.n5392 0.0148229
R12776 VPWR.n5506 VPWR.n5505 0.0148229
R12777 VPWR.n5693 VPWR.n5692 0.0148229
R12778 VPWR.n1600 VPWR.n1599 0.0148229
R12779 VPWR.n1737 VPWR.n1735 0.0148229
R12780 VPWR.n1733 VPWR.n1732 0.0148229
R12781 VPWR.n5246 VPWR.n5245 0.0148229
R12782 VPWR.n4849 VPWR.n4848 0.0148229
R12783 VPWR VPWR.n2485 0.0148229
R12784 VPWR.n5167 VPWR.n5166 0.0148229
R12785 VPWR.n5078 VPWR.n5077 0.0148229
R12786 VPWR.n4980 VPWR.n4979 0.0148229
R12787 VPWR.n2282 VPWR.n2281 0.0148229
R12788 VPWR.n2650 VPWR.n2648 0.0148229
R12789 VPWR.n2646 VPWR.n2645 0.0148229
R12790 VPWR.n4370 VPWR.n4369 0.0148229
R12791 VPWR.n4550 VPWR.n4549 0.0148229
R12792 VPWR.n3455 VPWR.n3454 0.0148229
R12793 VPWR.n3566 VPWR.n3565 0.0148229
R12794 VPWR.n4295 VPWR.n4294 0.0148229
R12795 VPWR.n2961 VPWR.n2960 0.0148229
R12796 VPWR.n7719 VPWR.n7718 0.0148229
R12797 VPWR.n7846 VPWR.n7844 0.0148229
R12798 VPWR.n7848 VPWR.n7847 0.0148229
R12799 VPWR.n9259 VPWR.n9258 0.0148229
R12800 VPWR.n122 VPWR.n121 0.0148229
R12801 VPWR.n3303 VPWR.n3302 0.0148229
R12802 VPWR.n3842 VPWR.n3840 0.0148229
R12803 VPWR.n3838 VPWR.n3837 0.0148229
R12804 VPWR.n3946 VPWR.n3945 0.0148229
R12805 VPWR.n4145 VPWR.n4144 0.0148229
R12806 VPWR.n7584 VPWR.n7583 0.0148229
R12807 VPWR.n7428 VPWR.n7426 0.0148229
R12808 VPWR.n7424 VPWR.n7423 0.0148229
R12809 VPWR.n7344 VPWR.n7343 0.0148229
R12810 VPWR.n7217 VPWR.n7216 0.0148229
R12811 VPWR.n9106 VPWR.n9105 0.0145155
R12812 VPWR.n312 VPWR.n311 0.0145155
R12813 VPWR.n180 VPWR.n179 0.0145155
R12814 VPWR.n179 VPWR.n178 0.0145155
R12815 VPWR.n6890 VPWR.n6889 0.0145155
R12816 VPWR.n6889 VPWR.n6888 0.0145155
R12817 VPWR.n7974 VPWR.n7973 0.0145155
R12818 VPWR.n7973 VPWR.n7972 0.0145155
R12819 VPWR.n329 VPWR.n328 0.0145155
R12820 VPWR.n328 VPWR.n327 0.0145155
R12821 VPWR.n8228 VPWR.n8227 0.0145155
R12822 VPWR.n8229 VPWR.n8228 0.0145155
R12823 VPWR.n6858 VPWR.n6857 0.0145155
R12824 VPWR.n6857 VPWR.n6856 0.0145155
R12825 VPWR.n5912 VPWR.n5911 0.0145155
R12826 VPWR.n5911 VPWR.n5910 0.0145155
R12827 VPWR.n8808 VPWR.n8807 0.0145155
R12828 VPWR.n8807 VPWR.n8806 0.0145155
R12829 VPWR.n8547 VPWR.n8546 0.0145155
R12830 VPWR.n8546 VPWR.n8545 0.0145155
R12831 VPWR.n6579 VPWR.n6578 0.0145155
R12832 VPWR.n6578 VPWR.n6577 0.0145155
R12833 VPWR.n8411 VPWR.n8410 0.0145155
R12834 VPWR.n8410 VPWR.n8409 0.0145155
R12835 VPWR.n377 VPWR.n376 0.0145155
R12836 VPWR.n376 VPWR.n375 0.0145155
R12837 VPWR.n1066 VPWR.n1065 0.0145155
R12838 VPWR.n1065 VPWR.n1064 0.0145155
R12839 VPWR.n682 VPWR.n681 0.0145155
R12840 VPWR.n681 VPWR.n680 0.0145155
R12841 VPWR.n918 VPWR.n917 0.0145155
R12842 VPWR.n917 VPWR.n916 0.0145155
R12843 VPWR.n5719 VPWR.n5718 0.0145155
R12844 VPWR.n5718 VPWR.n5717 0.0145155
R12845 VPWR.n5548 VPWR.n5547 0.0145155
R12846 VPWR.n5547 VPWR.n5546 0.0145155
R12847 VPWR.n1259 VPWR.n1258 0.0145155
R12848 VPWR.n1258 VPWR.n1257 0.0145155
R12849 VPWR.n5384 VPWR.n5383 0.0145155
R12850 VPWR.n5385 VPWR.n5384 0.0145155
R12851 VPWR.n4608 VPWR.n4607 0.0145155
R12852 VPWR.n4607 VPWR.n4606 0.0145155
R12853 VPWR.n5239 VPWR.n5238 0.0145155
R12854 VPWR.n5238 VPWR.n5237 0.0145155
R12855 VPWR.n1621 VPWR.n1620 0.0145155
R12856 VPWR.n1622 VPWR.n1621 0.0145155
R12857 VPWR.n5352 VPWR.n5351 0.0145155
R12858 VPWR.n5351 VPWR.n5350 0.0145155
R12859 VPWR.n4892 VPWR.n4891 0.0145155
R12860 VPWR.n4891 VPWR.n4890 0.0145155
R12861 VPWR.n5058 VPWR.n5057 0.0145155
R12862 VPWR.n5057 VPWR.n5056 0.0145155
R12863 VPWR.n2515 VPWR.n2514 0.0145155
R12864 VPWR.n2514 VPWR.n2513 0.0145155
R12865 VPWR.n5195 VPWR.n5194 0.0145155
R12866 VPWR.n5194 VPWR.n5193 0.0145155
R12867 VPWR.n2406 VPWR.n2405 0.0145155
R12868 VPWR.n2405 VPWR.n2404 0.0145155
R12869 VPWR.n2761 VPWR.n2760 0.0145155
R12870 VPWR.n2760 VPWR.n2759 0.0145155
R12871 VPWR.n4579 VPWR.n4578 0.0145155
R12872 VPWR.n2612 VPWR.n2611 0.0145155
R12873 VPWR.n2611 VPWR.n2610 0.0145155
R12874 VPWR.n7008 VPWR.n7007 0.0145155
R12875 VPWR.n7007 VPWR.n7006 0.0145155
R12876 VPWR.n4214 VPWR.n4213 0.0145155
R12877 VPWR.n4213 VPWR.n4212 0.0145155
R12878 VPWR.n3472 VPWR.n3471 0.0145155
R12879 VPWR.n4323 VPWR.n4322 0.0145155
R12880 VPWR.n3761 VPWR.n3760 0.0145155
R12881 VPWR.n3806 VPWR.n3805 0.0145155
R12882 VPWR.n3807 VPWR.n3806 0.0145155
R12883 VPWR.n6978 VPWR.n6977 0.0145155
R12884 VPWR.n6977 VPWR.n6976 0.0145155
R12885 VPWR.n3019 VPWR.n3018 0.0145155
R12886 VPWR.n3020 VPWR.n3019 0.0145155
R12887 VPWR.n11 VPWR.n10 0.0145155
R12888 VPWR.n12 VPWR.n11 0.0145155
R12889 VPWR.n9240 VPWR.n9239 0.0145155
R12890 VPWR.n9241 VPWR.n9240 0.0145155
R12891 VPWR.n7632 VPWR.n7631 0.0145155
R12892 VPWR.n7631 VPWR.n7630 0.0145155
R12893 VPWR.n6903 VPWR.n6902 0.0145155
R12894 VPWR.n6902 VPWR.n6901 0.0145155
R12895 VPWR.n3343 VPWR.n3342 0.0145155
R12896 VPWR.n3342 VPWR.n3341 0.0145155
R12897 VPWR.n4188 VPWR.n4187 0.0145155
R12898 VPWR.n4189 VPWR.n4188 0.0145155
R12899 VPWR.n7245 VPWR.n7244 0.0145155
R12900 VPWR.n7244 VPWR.n7243 0.0145155
R12901 VPWR.n3355 VPWR.n3354 0.0140135
R12902 VPWR.n3338 VPWR.n3335 0.0140135
R12903 VPWR.n160 VPWR.n159 0.0140135
R12904 VPWR.n9117 VPWR.n9111 0.0140135
R12905 VPWR.n9269 VPWR.n9268 0.0140135
R12906 VPWR.n9232 VPWR.n9231 0.0140135
R12907 VPWR.n9236 VPWR.n9235 0.0140135
R12908 VPWR.n310 VPWR.n309 0.0140135
R12909 VPWR.n8954 VPWR.n8948 0.0140135
R12910 VPWR.n183 VPWR.n182 0.0140135
R12911 VPWR.n186 VPWR.n185 0.0140135
R12912 VPWR.n9096 VPWR.n9095 0.0140135
R12913 VPWR.n6151 VPWR.n6150 0.0140135
R12914 VPWR.n6885 VPWR.n6153 0.0140135
R12915 VPWR.n7969 VPWR.n7866 0.0140135
R12916 VPWR.n7968 VPWR.n7967 0.0140135
R12917 VPWR.n7874 VPWR.n7873 0.0140135
R12918 VPWR.n8939 VPWR.n8938 0.0140135
R12919 VPWR.n324 VPWR.n320 0.0140135
R12920 VPWR.n8215 VPWR.n8214 0.0140135
R12921 VPWR.n8218 VPWR.n8217 0.0140135
R12922 VPWR.n8224 VPWR.n8223 0.0140135
R12923 VPWR.n6847 VPWR.n6846 0.0140135
R12924 VPWR.n6853 VPWR.n6849 0.0140135
R12925 VPWR.n5907 VPWR.n5903 0.0140135
R12926 VPWR.n5906 VPWR.n5905 0.0140135
R12927 VPWR.n5920 VPWR.n5919 0.0140135
R12928 VPWR.n8819 VPWR.n8818 0.0140135
R12929 VPWR.n8803 VPWR.n348 0.0140135
R12930 VPWR.n8517 VPWR.n8516 0.0140135
R12931 VPWR.n8520 VPWR.n8519 0.0140135
R12932 VPWR.n8551 VPWR.n8550 0.0140135
R12933 VPWR.n6568 VPWR.n6567 0.0140135
R12934 VPWR.n6574 VPWR.n6570 0.0140135
R12935 VPWR.n8406 VPWR.n8402 0.0140135
R12936 VPWR.n8405 VPWR.n8404 0.0140135
R12937 VPWR.n5881 VPWR.n5880 0.0140135
R12938 VPWR.n5849 VPWR.n5848 0.0140135
R12939 VPWR.n372 VPWR.n368 0.0140135
R12940 VPWR.n1044 VPWR.n1043 0.0140135
R12941 VPWR.n1047 VPWR.n1046 0.0140135
R12942 VPWR.n1070 VPWR.n1069 0.0140135
R12943 VPWR.n686 VPWR.n685 0.0140135
R12944 VPWR.n591 VPWR.n590 0.0140135
R12945 VPWR.n913 VPWR.n797 0.0140135
R12946 VPWR.n912 VPWR.n911 0.0140135
R12947 VPWR.n768 VPWR.n767 0.0140135
R12948 VPWR.n5730 VPWR.n5729 0.0140135
R12949 VPWR.n5714 VPWR.n5710 0.0140135
R12950 VPWR.n476 VPWR.n475 0.0140135
R12951 VPWR.n479 VPWR.n478 0.0140135
R12952 VPWR.n5552 VPWR.n5551 0.0140135
R12953 VPWR.n1248 VPWR.n1247 0.0140135
R12954 VPWR.n1254 VPWR.n1250 0.0140135
R12955 VPWR.n5388 VPWR.n504 0.0140135
R12956 VPWR.n5391 VPWR.n5389 0.0140135
R12957 VPWR.n5373 VPWR.n5372 0.0140135
R12958 VPWR.n4619 VPWR.n4618 0.0140135
R12959 VPWR.n4603 VPWR.n4599 0.0140135
R12960 VPWR.n1798 VPWR.n1797 0.0140135
R12961 VPWR.n5244 VPWR.n5243 0.0140135
R12962 VPWR.n5242 VPWR.n1800 0.0140135
R12963 VPWR.n576 VPWR.n575 0.0140135
R12964 VPWR.n1625 VPWR.n563 0.0140135
R12965 VPWR.n5347 VPWR.n5343 0.0140135
R12966 VPWR.n5346 VPWR.n5345 0.0140135
R12967 VPWR.n519 VPWR.n518 0.0140135
R12968 VPWR.n4903 VPWR.n4902 0.0140135
R12969 VPWR.n4887 VPWR.n4883 0.0140135
R12970 VPWR.n1858 VPWR.n1857 0.0140135
R12971 VPWR.n1861 VPWR.n1860 0.0140135
R12972 VPWR.n5062 VPWR.n5061 0.0140135
R12973 VPWR.n2519 VPWR.n2518 0.0140135
R12974 VPWR.n2510 VPWR.n2506 0.0140135
R12975 VPWR.n5190 VPWR.n5186 0.0140135
R12976 VPWR.n5189 VPWR.n5188 0.0140135
R12977 VPWR.n1819 VPWR.n1818 0.0140135
R12978 VPWR.n2209 VPWR.n2208 0.0140135
R12979 VPWR.n2401 VPWR.n2211 0.0140135
R12980 VPWR.n2740 VPWR.n2739 0.0140135
R12981 VPWR.n2743 VPWR.n2742 0.0140135
R12982 VPWR.n2749 VPWR.n2748 0.0140135
R12983 VPWR.n4589 VPWR.n4588 0.0140135
R12984 VPWR.n1989 VPWR.n1983 0.0140135
R12985 VPWR.n2607 VPWR.n2603 0.0140135
R12986 VPWR.n2606 VPWR.n2605 0.0140135
R12987 VPWR.n2103 VPWR.n2102 0.0140135
R12988 VPWR.n5994 VPWR.n5991 0.0140135
R12989 VPWR.n5993 VPWR.n5992 0.0140135
R12990 VPWR.n6002 VPWR.n6001 0.0140135
R12991 VPWR.n4217 VPWR.n2869 0.0140135
R12992 VPWR.n2956 VPWR.n2955 0.0140135
R12993 VPWR.n3437 VPWR.n3436 0.0140135
R12994 VPWR.n3477 VPWR.n3470 0.0140135
R12995 VPWR.n4326 VPWR.n4325 0.0140135
R12996 VPWR.n4329 VPWR.n4328 0.0140135
R12997 VPWR.n4333 VPWR.n4332 0.0140135
R12998 VPWR.n3771 VPWR.n3765 0.0140135
R12999 VPWR.n3770 VPWR.n3769 0.0140135
R13000 VPWR.n3767 VPWR.n3766 0.0140135
R13001 VPWR.n3819 VPWR.n3813 0.0140135
R13002 VPWR.n3818 VPWR.n3817 0.0140135
R13003 VPWR.n3815 VPWR.n3814 0.0140135
R13004 VPWR.n6967 VPWR.n6964 0.0140135
R13005 VPWR.n6966 VPWR.n6965 0.0140135
R13006 VPWR.n6959 VPWR.n6958 0.0140135
R13007 VPWR.n3924 VPWR.n3923 0.0140135
R13008 VPWR.n3011 VPWR.n3010 0.0140135
R13009 VPWR.n3015 VPWR.n3014 0.0140135
R13010 VPWR.n7320 VPWR.n7319 0.0140135
R13011 VPWR.n7317 VPWR.n7316 0.0140135
R13012 VPWR.n7315 VPWR.n7314 0.0140135
R13013 VPWR.n7628 VPWR.n7627 0.0140135
R13014 VPWR.n7702 VPWR.n7698 0.0140135
R13015 VPWR.n6915 VPWR.n6914 0.0140135
R13016 VPWR.n6929 VPWR.n6926 0.0140135
R13017 VPWR.n4184 VPWR.n4183 0.0140135
R13018 VPWR.n4201 VPWR.n4195 0.0140135
R13019 VPWR.n7254 VPWR.n7253 0.0140135
R13020 VPWR.n7240 VPWR.n7237 0.0140135
R13021 VPWR.n8254 VPWR.n8253 0.0139925
R13022 VPWR.n8574 VPWR.n8573 0.0139925
R13023 VPWR.n1092 VPWR.n1091 0.0139925
R13024 VPWR.n5515 VPWR.n5514 0.0139925
R13025 VPWR.n5254 VPWR.n5253 0.0139925
R13026 VPWR.n5084 VPWR.n5083 0.0139925
R13027 VPWR.n3940 VPWR.n3934 0.0139925
R13028 VPWR.n8061 VPWR.n8059 0.0139925
R13029 VPWR.n4364 VPWR.n4359 0.0139925
R13030 VPWR.n4301 VPWR.n4300 0.0139925
R13031 VPWR.n9265 VPWR.n9264 0.0139925
R13032 VPWR.n7349 VPWR.n7325 0.0139925
R13033 VPWR.n6220 VPWR.n6216 0.0135208
R13034 VPWR.n7869 VPWR.n7868 0.0135208
R13035 VPWR.n8071 VPWR.n8069 0.0135208
R13036 VPWR.n8067 VPWR.n8064 0.0135208
R13037 VPWR.n9084 VPWR 0.0135208
R13038 VPWR.n277 VPWR.n276 0.0135208
R13039 VPWR.n6814 VPWR.n6813 0.0135208
R13040 VPWR.n8246 VPWR.n8244 0.0135208
R13041 VPWR.n8934 VPWR.n8853 0.0135208
R13042 VPWR.n6563 VPWR.n6562 0.0135208
R13043 VPWR.n8560 VPWR.n8559 0.0135208
R13044 VPWR.n8558 VPWR.n8557 0.0135208
R13045 VPWR.n8536 VPWR 0.0135208
R13046 VPWR.n8718 VPWR.n8717 0.0135208
R13047 VPWR.n8793 VPWR 0.0135208
R13048 VPWR.n695 VPWR.n691 0.0135208
R13049 VPWR VPWR.n708 0.0135208
R13050 VPWR.n903 VPWR.n902 0.0135208
R13051 VPWR.n5844 VPWR.n5764 0.0135208
R13052 VPWR.n1349 VPWR.n1346 0.0135208
R13053 VPWR.n1397 VPWR.n1395 0.0135208
R13054 VPWR.n5504 VPWR.n5502 0.0135208
R13055 VPWR.n5500 VPWR.n5498 0.0135208
R13056 VPWR.n5688 VPWR.n5687 0.0135208
R13057 VPWR.n1595 VPWR.n1594 0.0135208
R13058 VPWR.n1741 VPWR.n1739 0.0135208
R13059 VPWR.n1796 VPWR.n1793 0.0135208
R13060 VPWR.n4856 VPWR.n4853 0.0135208
R13061 VPWR.n2526 VPWR.n2524 0.0135208
R13062 VPWR.n5076 VPWR.n5074 0.0135208
R13063 VPWR.n5072 VPWR.n5070 0.0135208
R13064 VPWR.n4975 VPWR.n4974 0.0135208
R13065 VPWR.n2287 VPWR.n2286 0.0135208
R13066 VPWR.n2675 VPWR 0.0135208
R13067 VPWR.n2654 VPWR.n2652 0.0135208
R13068 VPWR.n4374 VPWR.n4372 0.0135208
R13069 VPWR.n4380 VPWR.n4376 0.0135208
R13070 VPWR.n4555 VPWR.n4554 0.0135208
R13071 VPWR.n3462 VPWR.n3459 0.0135208
R13072 VPWR.n4293 VPWR.n4291 0.0135208
R13073 VPWR.n4289 VPWR.n4287 0.0135208
R13074 VPWR.n2947 VPWR.n2943 0.0135208
R13075 VPWR.n7714 VPWR.n7713 0.0135208
R13076 VPWR.n7842 VPWR.n7840 0.0135208
R13077 VPWR.n129 VPWR.n126 0.0135208
R13078 VPWR.n3310 VPWR.n3307 0.0135208
R13079 VPWR.n3846 VPWR.n3844 0.0135208
R13080 VPWR.n3948 VPWR.n3947 0.0135208
R13081 VPWR.n3950 VPWR.n3949 0.0135208
R13082 VPWR VPWR.n3961 0.0135208
R13083 VPWR.n4152 VPWR.n4149 0.0135208
R13084 VPWR.n7591 VPWR.n7588 0.0135208
R13085 VPWR.n7432 VPWR.n7430 0.0135208
R13086 VPWR.n7342 VPWR.n7341 0.0135208
R13087 VPWR.n7340 VPWR.n7339 0.0135208
R13088 VPWR.n7327 VPWR 0.0135208
R13089 VPWR.n7212 VPWR.n7211 0.0135208
R13090 VPWR.n9075 VPWR.n9074 0.0130912
R13091 VPWR.n6318 VPWR.n6317 0.0130912
R13092 VPWR.n7879 VPWR.n7878 0.0130912
R13093 VPWR.n8859 VPWR.n8858 0.0130912
R13094 VPWR.n8094 VPWR.n8093 0.0130912
R13095 VPWR.n6786 VPWR.n6785 0.0130912
R13096 VPWR.n5918 VPWR.n5917 0.0130912
R13097 VPWR.n8728 VPWR.n8727 0.0130912
R13098 VPWR.n360 VPWR.n359 0.0130912
R13099 VPWR.n6336 VPWR.n6335 0.0130912
R13100 VPWR.n5886 VPWR.n5885 0.0130912
R13101 VPWR.n5770 VPWR.n5769 0.0130912
R13102 VPWR.n745 VPWR.n744 0.0130912
R13103 VPWR.n580 VPWR.n579 0.0130912
R13104 VPWR.n773 VPWR.n772 0.0130912
R13105 VPWR.n397 VPWR.n396 0.0130912
R13106 VPWR.n5524 VPWR.n5523 0.0130912
R13107 VPWR.n1266 VPWR.n1265 0.0130912
R13108 VPWR.n5371 VPWR.n5370 0.0130912
R13109 VPWR.n4624 VPWR.n4623 0.0130912
R13110 VPWR.n5215 VPWR.n5214 0.0130912
R13111 VPWR.n1530 VPWR.n1529 0.0130912
R13112 VPWR.n517 VPWR.n516 0.0130912
R13113 VPWR.n4908 VPWR.n4907 0.0130912
R13114 VPWR.n1873 VPWR.n1872 0.0130912
R13115 VPWR.n2414 VPWR.n2413 0.0130912
R13116 VPWR.n1824 VPWR.n1823 0.0130912
R13117 VPWR.n2385 VPWR.n2384 0.0130912
R13118 VPWR.n4341 VPWR.n4340 0.0130912
R13119 VPWR.n2108 VPWR.n2107 0.0130912
R13120 VPWR.n5998 VPWR.n5997 0.0130912
R13121 VPWR.n2877 VPWR.n2876 0.0130912
R13122 VPWR.n2971 VPWR.n2970 0.0130912
R13123 VPWR.n3441 VPWR.n3440 0.0130912
R13124 VPWR.n3776 VPWR.n3775 0.0130912
R13125 VPWR.n3122 VPWR.n3121 0.0130912
R13126 VPWR.n3098 VPWR.n3097 0.0130912
R13127 VPWR.n6971 VPWR.n6970 0.0130912
R13128 VPWR.n3930 VPWR.n3929 0.0130912
R13129 VPWR.n6 VPWR.n5 0.0130912
R13130 VPWR.n17 VPWR.n16 0.0130912
R13131 VPWR.n9275 VPWR.n9274 0.0130912
R13132 VPWR.n22 VPWR.n21 0.0130912
R13133 VPWR.n7699 VPWR.n6137 0.0130912
R13134 VPWR.n6933 VPWR.n6932 0.0130912
R13135 VPWR.n3134 VPWR.n3133 0.0130912
R13136 VPWR.n3138 VPWR.n3137 0.0130912
R13137 VPWR.n2988 VPWR.n2987 0.0130912
R13138 VPWR.n7258 VPWR.n7257 0.0130912
R13139 VPWR.n7231 VPWR.n7230 0.0130912
R13140 VPWR.n2875 VPWR.n2874 0.0126061
R13141 VPWR.n3443 VPWR.n3442 0.0126061
R13142 VPWR.n3120 VPWR.n3119 0.0126061
R13143 VPWR.n9268 VPWR.n9267 0.0123243
R13144 VPWR.n9247 VPWR.n9246 0.0123243
R13145 VPWR.n9229 VPWR.n9228 0.0123243
R13146 VPWR.n184 VPWR.n183 0.0123243
R13147 VPWR.n171 VPWR.n170 0.0123243
R13148 VPWR.n173 VPWR.n172 0.0123243
R13149 VPWR.n7979 VPWR.n7978 0.0123243
R13150 VPWR.n8216 VPWR.n8215 0.0123243
R13151 VPWR.n8234 VPWR.n8233 0.0123243
R13152 VPWR.n5954 VPWR.n5953 0.0123243
R13153 VPWR.n5899 VPWR.n5898 0.0123243
R13154 VPWR.n8518 VPWR.n8517 0.0123243
R13155 VPWR.n8527 VPWR.n8526 0.0123243
R13156 VPWR.n8529 VPWR.n8528 0.0123243
R13157 VPWR.n8398 VPWR.n8397 0.0123243
R13158 VPWR.n1045 VPWR.n1044 0.0123243
R13159 VPWR.n1053 VPWR.n1052 0.0123243
R13160 VPWR.n1055 VPWR.n1054 0.0123243
R13161 VPWR.n896 VPWR.n895 0.0123243
R13162 VPWR.n477 VPWR.n476 0.0123243
R13163 VPWR.n5539 VPWR.n5538 0.0123243
R13164 VPWR.n5541 VPWR.n5540 0.0123243
R13165 VPWR.n1400 VPWR.n1399 0.0123243
R13166 VPWR.n1799 VPWR.n1798 0.0123243
R13167 VPWR.n5230 VPWR.n5229 0.0123243
R13168 VPWR.n5232 VPWR.n5231 0.0123243
R13169 VPWR.n5339 VPWR.n5338 0.0123243
R13170 VPWR.n1859 VPWR.n1858 0.0123243
R13171 VPWR.n5049 VPWR.n5048 0.0123243
R13172 VPWR.n5051 VPWR.n5050 0.0123243
R13173 VPWR.n5182 VPWR.n5181 0.0123243
R13174 VPWR.n2741 VPWR.n2740 0.0123243
R13175 VPWR.n2752 VPWR.n2751 0.0123243
R13176 VPWR.n2754 VPWR.n2753 0.0123243
R13177 VPWR.n2622 VPWR.n2621 0.0123243
R13178 VPWR.n7018 VPWR.n7017 0.0123243
R13179 VPWR.n6001 VPWR.n6000 0.0123243
R13180 VPWR.n4327 VPWR.n4326 0.0123243
R13181 VPWR.n2773 VPWR.n2772 0.0123243
R13182 VPWR.n2777 VPWR.n2776 0.0123243
R13183 VPWR.n3789 VPWR.n3788 0.0123243
R13184 VPWR.n3768 VPWR.n3767 0.0123243
R13185 VPWR.n3801 VPWR.n3800 0.0123243
R13186 VPWR.n3816 VPWR.n3815 0.0123243
R13187 VPWR.n6988 VPWR.n6987 0.0123243
R13188 VPWR.n6958 VPWR.n6957 0.0123243
R13189 VPWR.n3026 VPWR.n3025 0.0123243
R13190 VPWR.n3966 VPWR.n3965 0.0123243
R13191 VPWR.n7319 VPWR.n7318 0.0123243
R13192 VPWR.n7308 VPWR.n7307 0.0123243
R13193 VPWR.n7304 VPWR.n7303 0.0123243
R13194 VPWR.n6880 VPWR.n6879 0.0122188
R13195 VPWR.n8008 VPWR.n8007 0.0122188
R13196 VPWR.n9067 VPWR.n9066 0.0122188
R13197 VPWR.n266 VPWR.n265 0.0122188
R13198 VPWR.n269 VPWR.n268 0.0122188
R13199 VPWR.n6805 VPWR.n6804 0.0122188
R13200 VPWR.n6802 VPWR.n6801 0.0122188
R13201 VPWR.n6690 VPWR.n6689 0.0122188
R13202 VPWR.n8201 VPWR.n8200 0.0122188
R13203 VPWR.n340 VPWR.n339 0.0122188
R13204 VPWR.n8842 VPWR.n8841 0.0122188
R13205 VPWR.n8845 VPWR.n8844 0.0122188
R13206 VPWR.n6478 VPWR.n6477 0.0122188
R13207 VPWR.n6475 VPWR.n6474 0.0122188
R13208 VPWR.n6467 VPWR 0.0122188
R13209 VPWR.n6342 VPWR.n6329 0.0122188
R13210 VPWR.n6439 VPWR.n6438 0.0122188
R13211 VPWR.n8592 VPWR.n8591 0.0122188
R13212 VPWR.n8707 VPWR.n8706 0.0122188
R13213 VPWR.n8710 VPWR.n8709 0.0122188
R13214 VPWR.n706 VPWR.n705 0.0122188
R13215 VPWR.n1228 VPWR.n1227 0.0122188
R13216 VPWR.n873 VPWR.n872 0.0122188
R13217 VPWR.n734 VPWR.n733 0.0122188
R13218 VPWR.n389 VPWR.n388 0.0122188
R13219 VPWR.n1355 VPWR.n1354 0.0122188
R13220 VPWR.n1359 VPWR.n1357 0.0122188
R13221 VPWR.n1369 VPWR.n1368 0.0122188
R13222 VPWR.n1426 VPWR.n1424 0.0122188
R13223 VPWR.n5577 VPWR.n5575 0.0122188
R13224 VPWR.n5666 VPWR.n5665 0.0122188
R13225 VPWR.n5676 VPWR.n5675 0.0122188
R13226 VPWR.n5679 VPWR.n5678 0.0122188
R13227 VPWR.n1634 VPWR.n1632 0.0122188
R13228 VPWR.n1769 VPWR.n1768 0.0122188
R13229 VPWR.n4674 VPWR.n4673 0.0122188
R13230 VPWR.n4865 VPWR.n4864 0.0122188
R13231 VPWR.n4862 VPWR.n4861 0.0122188
R13232 VPWR.n2534 VPWR.n2533 0.0122188
R13233 VPWR.n2538 VPWR.n2536 0.0122188
R13234 VPWR.n2579 VPWR.n2578 0.0122188
R13235 VPWR.n5034 VPWR.n5033 0.0122188
R13236 VPWR.n4999 VPWR.n4998 0.0122188
R13237 VPWR.n4967 VPWR.n1965 0.0122188
R13238 VPWR.n4970 VPWR.n4969 0.0122188
R13239 VPWR.n2396 VPWR.n2395 0.0122188
R13240 VPWR.n2680 VPWR.n2678 0.0122188
R13241 VPWR.n4403 VPWR.n4399 0.0122188
R13242 VPWR.n4563 VPWR.n4562 0.0122188
R13243 VPWR.n4560 VPWR.n4559 0.0122188
R13244 VPWR.n3488 VPWR.n3486 0.0122188
R13245 VPWR.n3750 VPWR.n3749 0.0122188
R13246 VPWR.n3543 VPWR.n3542 0.0122188
R13247 VPWR.n4266 VPWR.n4265 0.0122188
R13248 VPWR.n7694 VPWR.n7693 0.0122188
R13249 VPWR.n7818 VPWR.n7817 0.0122188
R13250 VPWR.n9207 VPWR.n9206 0.0122188
R13251 VPWR.n137 VPWR.n136 0.0122188
R13252 VPWR.n134 VPWR.n133 0.0122188
R13253 VPWR.n3316 VPWR.n3315 0.0122188
R13254 VPWR.n3321 VPWR.n3318 0.0122188
R13255 VPWR.n3868 VPWR.n3867 0.0122188
R13256 VPWR.n3988 VPWR.n3986 0.0122188
R13257 VPWR.n4162 VPWR.n4160 0.0122188
R13258 VPWR.n4158 VPWR.n4157 0.0122188
R13259 VPWR.n7597 VPWR.n7596 0.0122188
R13260 VPWR.n7602 VPWR.n7599 0.0122188
R13261 VPWR.n7453 VPWR.n7451 0.0122188
R13262 VPWR.n7055 VPWR.n7054 0.0122188
R13263 VPWR.n7201 VPWR.n7200 0.0122188
R13264 VPWR.n7204 VPWR.n7203 0.0122188
R13265 VPWR.n2290 VPWR.n2289 0.0120783
R13266 VPWR.n2279 VPWR.n2278 0.01206
R13267 VPWR.n3755 VPWR.n3754 0.0118576
R13268 VPWR.n3530 VPWR.n3123 0.0118576
R13269 VPWR.n4308 VPWR.n4306 0.0118576
R13270 VPWR.n4318 VPWR.n4316 0.0118576
R13271 VPWR.n2972 VPWR.n2969 0.0118576
R13272 VPWR.n8244 VPWR.n8243 0.0115187
R13273 VPWR.n5763 VPWR.n5761 0.0114378
R13274 VPWR.n4973 VPWR.n4972 0.0114378
R13275 VPWR.n4983 VPWR.n4982 0.0114077
R13276 VPWR.n1078 VPWR.n1077 0.0111911
R13277 VPWR.n6222 VPWR.n6221 0.0109167
R13278 VPWR.n6224 VPWR.n6222 0.0109167
R13279 VPWR.n6879 VPWR.n6876 0.0109167
R13280 VPWR.n6874 VPWR.n6872 0.0109167
R13281 VPWR.n8002 VPWR.n8001 0.0109167
R13282 VPWR.n7964 VPWR.n7963 0.0109167
R13283 VPWR.n8075 VPWR.n8074 0.0109167
R13284 VPWR.n8072 VPWR.n8071 0.0109167
R13285 VPWR.n9071 VPWR.n192 0.0109167
R13286 VPWR.n262 VPWR.n260 0.0109167
R13287 VPWR.n265 VPWR.n262 0.0109167
R13288 VPWR.n272 VPWR.n271 0.0109167
R13289 VPWR.n6809 VPWR.n6808 0.0109167
R13290 VPWR.n6808 VPWR.n6807 0.0109167
R13291 VPWR.n6801 VPWR.n6798 0.0109167
R13292 VPWR.n6796 VPWR.n6794 0.0109167
R13293 VPWR.n6685 VPWR.n6684 0.0109167
R13294 VPWR.n6665 VPWR.n6664 0.0109167
R13295 VPWR.n6662 VPWR.n6661 0.0109167
R13296 VPWR.n8250 VPWR.n8249 0.0109167
R13297 VPWR.n8247 VPWR.n8246 0.0109167
R13298 VPWR VPWR.n8236 0.0109167
R13299 VPWR.n8207 VPWR.n8108 0.0109167
R13300 VPWR.n8839 VPWR.n8837 0.0109167
R13301 VPWR.n8841 VPWR.n8839 0.0109167
R13302 VPWR.n8848 VPWR.n8847 0.0109167
R13303 VPWR.n6482 VPWR.n6481 0.0109167
R13304 VPWR.n6481 VPWR.n6480 0.0109167
R13305 VPWR.n6474 VPWR.n6472 0.0109167
R13306 VPWR.n6469 VPWR.n6467 0.0109167
R13307 VPWR.n6434 VPWR.n6423 0.0109167
R13308 VPWR.n8389 VPWR.n8388 0.0109167
R13309 VPWR.n8386 VPWR.n8385 0.0109167
R13310 VPWR.n8564 VPWR.n8563 0.0109167
R13311 VPWR.n8561 VPWR.n8560 0.0109167
R13312 VPWR.n8524 VPWR 0.0109167
R13313 VPWR.n8588 VPWR.n356 0.0109167
R13314 VPWR.n8713 VPWR.n8712 0.0109167
R13315 VPWR.n697 VPWR.n696 0.0109167
R13316 VPWR.n699 VPWR.n697 0.0109167
R13317 VPWR.n878 VPWR.n877 0.0109167
R13318 VPWR.n908 VPWR.n907 0.0109167
R13319 VPWR.n1083 VPWR.n1082 0.0109167
R13320 VPWR.n1080 VPWR.n1079 0.0109167
R13321 VPWR.n1050 VPWR 0.0109167
R13322 VPWR.n1106 VPWR.n738 0.0109167
R13323 VPWR.n5750 VPWR.n5748 0.0109167
R13324 VPWR.n5752 VPWR.n5750 0.0109167
R13325 VPWR.n5753 VPWR 0.0109167
R13326 VPWR.n5761 VPWR.n5760 0.0109167
R13327 VPWR.n1351 VPWR.n1350 0.0109167
R13328 VPWR.n1353 VPWR.n1351 0.0109167
R13329 VPWR.n1362 VPWR.n1359 0.0109167
R13330 VPWR.n1366 VPWR.n1364 0.0109167
R13331 VPWR.n1418 VPWR.n1417 0.0109167
R13332 VPWR.n5395 VPWR.n5394 0.0109167
R13333 VPWR.n5508 VPWR.n5507 0.0109167
R13334 VPWR.n5505 VPWR.n5504 0.0109167
R13335 VPWR.n5569 VPWR.n5568 0.0109167
R13336 VPWR.n5673 VPWR.n5671 0.0109167
R13337 VPWR.n5675 VPWR.n5673 0.0109167
R13338 VPWR.n5682 VPWR.n5681 0.0109167
R13339 VPWR.n1590 VPWR.n1589 0.0109167
R13340 VPWR.n1589 VPWR.n1588 0.0109167
R13341 VPWR.n1636 VPWR.n1634 0.0109167
R13342 VPWR.n1641 VPWR.n1638 0.0109167
R13343 VPWR.n1763 VPWR.n1752 0.0109167
R13344 VPWR.n1735 VPWR.n1733 0.0109167
R13345 VPWR.n1731 VPWR.n1730 0.0109167
R13346 VPWR.n5248 VPWR.n5247 0.0109167
R13347 VPWR.n5245 VPWR.n1796 0.0109167
R13348 VPWR.n4668 VPWR.n4667 0.0109167
R13349 VPWR.n4867 VPWR.n4866 0.0109167
R13350 VPWR.n4866 VPWR.n4865 0.0109167
R13351 VPWR.n4860 VPWR.n4858 0.0109167
R13352 VPWR.n2529 VPWR.n2528 0.0109167
R13353 VPWR.n2532 VPWR.n2529 0.0109167
R13354 VPWR.n2540 VPWR.n2538 0.0109167
R13355 VPWR.n2545 VPWR.n2543 0.0109167
R13356 VPWR.n2589 VPWR.n2588 0.0109167
R13357 VPWR.n5168 VPWR.n5167 0.0109167
R13358 VPWR.n5165 VPWR.n5164 0.0109167
R13359 VPWR.n5080 VPWR.n5079 0.0109167
R13360 VPWR.n5077 VPWR.n5076 0.0109167
R13361 VPWR.n5040 VPWR.n1887 0.0109167
R13362 VPWR.n4972 VPWR.n4971 0.0109167
R13363 VPWR.n2291 VPWR.n2290 0.0109167
R13364 VPWR.n2670 VPWR.n2669 0.0109167
R13365 VPWR.n2648 VPWR.n2646 0.0109167
R13366 VPWR.n2644 VPWR.n2643 0.0109167
R13367 VPWR.n4368 VPWR.n4367 0.0109167
R13368 VPWR.n4372 VPWR.n4370 0.0109167
R13369 VPWR.n4393 VPWR.n4392 0.0109167
R13370 VPWR.n4558 VPWR.n4557 0.0109167
R13371 VPWR.n3464 VPWR.n3463 0.0109167
R13372 VPWR.n3466 VPWR.n3464 0.0109167
R13373 VPWR.n3490 VPWR.n3488 0.0109167
R13374 VPWR.n3494 VPWR.n3492 0.0109167
R13375 VPWR.n3550 VPWR.n3549 0.0109167
R13376 VPWR.n3565 VPWR.n3564 0.0109167
R13377 VPWR.n3568 VPWR.n3567 0.0109167
R13378 VPWR.n4297 VPWR.n4296 0.0109167
R13379 VPWR.n4294 VPWR.n4293 0.0109167
R13380 VPWR.n4273 VPWR.n4272 0.0109167
R13381 VPWR.n4228 VPWR.n4226 0.0109167
R13382 VPWR.n4226 VPWR.n4224 0.0109167
R13383 VPWR VPWR.n4222 0.0109167
R13384 VPWR.n2939 VPWR.n2938 0.0109167
R13385 VPWR.n7709 VPWR.n7708 0.0109167
R13386 VPWR.n7708 VPWR.n7707 0.0109167
R13387 VPWR.n7693 VPWR.n7690 0.0109167
R13388 VPWR.n7688 VPWR.n6131 0.0109167
R13389 VPWR.n7826 VPWR.n7825 0.0109167
R13390 VPWR.n7847 VPWR.n7846 0.0109167
R13391 VPWR.n7850 VPWR.n7849 0.0109167
R13392 VPWR.n9261 VPWR.n9260 0.0109167
R13393 VPWR.n9258 VPWR.n9257 0.0109167
R13394 VPWR.n9213 VPWR.n29 0.0109167
R13395 VPWR.n132 VPWR.n131 0.0109167
R13396 VPWR.n3312 VPWR.n3311 0.0109167
R13397 VPWR.n3314 VPWR.n3312 0.0109167
R13398 VPWR.n3323 VPWR.n3321 0.0109167
R13399 VPWR.n3327 VPWR.n3325 0.0109167
R13400 VPWR.n3861 VPWR.n3860 0.0109167
R13401 VPWR.n3840 VPWR.n3838 0.0109167
R13402 VPWR.n3836 VPWR.n3835 0.0109167
R13403 VPWR.n3944 VPWR.n3943 0.0109167
R13404 VPWR.n3947 VPWR.n3946 0.0109167
R13405 VPWR.n3980 VPWR.n2999 0.0109167
R13406 VPWR.n4166 VPWR.n4164 0.0109167
R13407 VPWR.n4164 VPWR.n4162 0.0109167
R13408 VPWR.n4156 VPWR.n4154 0.0109167
R13409 VPWR.n7593 VPWR.n7592 0.0109167
R13410 VPWR.n7595 VPWR.n7593 0.0109167
R13411 VPWR.n7604 VPWR.n7602 0.0109167
R13412 VPWR.n7608 VPWR.n7606 0.0109167
R13413 VPWR.n7445 VPWR.n7444 0.0109167
R13414 VPWR.n7426 VPWR.n7424 0.0109167
R13415 VPWR.n7422 VPWR.n7421 0.0109167
R13416 VPWR.n7346 VPWR.n7345 0.0109167
R13417 VPWR.n7343 VPWR.n7342 0.0109167
R13418 VPWR.n9290 VPWR.n9289 0.0109167
R13419 VPWR.n7198 VPWR.n7196 0.0109167
R13420 VPWR.n7200 VPWR.n7198 0.0109167
R13421 VPWR.n7207 VPWR.n7206 0.0109167
R13422 VPWR.n5974 VPWR.n5973 0.0106351
R13423 VPWR.n5893 VPWR.n5892 0.0106351
R13424 VPWR.n8366 VPWR.n8365 0.0106351
R13425 VPWR.n792 VPWR.n791 0.0106351
R13426 VPWR.n509 VPWR.n508 0.0106351
R13427 VPWR.n5333 VPWR.n5332 0.0106351
R13428 VPWR.n1811 VPWR.n1810 0.0106351
R13429 VPWR.n2616 VPWR.n2615 0.0106351
R13430 VPWR.n7012 VPWR.n7011 0.0106351
R13431 VPWR.n3783 VPWR.n3782 0.0106351
R13432 VPWR.n3797 VPWR.n3796 0.0106351
R13433 VPWR.n6982 VPWR.n6981 0.0106351
R13434 VPWR.n8422 VPWR 0.0101142
R13435 VPWR VPWR.n929 0.0101142
R13436 VPWR.n161 VPWR.n150 0.00975758
R13437 VPWR.n152 VPWR.n151 0.00975758
R13438 VPWR.n9107 VPWR.n9106 0.00975758
R13439 VPWR.n9120 VPWR.n9119 0.00975758
R13440 VPWR.n314 VPWR.n301 0.00975758
R13441 VPWR.n313 VPWR.n312 0.00975758
R13442 VPWR.n8945 VPWR.n8944 0.00975758
R13443 VPWR.n8957 VPWR.n8956 0.00975758
R13444 VPWR.n9097 VPWR.n168 0.00975758
R13445 VPWR.n181 VPWR.n180 0.00975758
R13446 VPWR.n178 VPWR.n177 0.00975758
R13447 VPWR.n6892 VPWR.n6140 0.00975758
R13448 VPWR.n6891 VPWR.n6890 0.00975758
R13449 VPWR.n6888 VPWR.n6887 0.00975758
R13450 VPWR.n7976 VPWR.n5977 0.00975758
R13451 VPWR.n7975 VPWR.n7974 0.00975758
R13452 VPWR.n7972 VPWR.n7971 0.00975758
R13453 VPWR.n8940 VPWR.n318 0.00975758
R13454 VPWR.n330 VPWR.n329 0.00975758
R13455 VPWR.n327 VPWR.n326 0.00975758
R13456 VPWR.n8225 VPWR.n5957 0.00975758
R13457 VPWR.n8227 VPWR.n8226 0.00975758
R13458 VPWR.n8230 VPWR.n8229 0.00975758
R13459 VPWR.n6860 VPWR.n6836 0.00975758
R13460 VPWR.n6859 VPWR.n6858 0.00975758
R13461 VPWR.n6856 VPWR.n6855 0.00975758
R13462 VPWR.n5914 VPWR.n5890 0.00975758
R13463 VPWR.n5913 VPWR.n5912 0.00975758
R13464 VPWR.n5910 VPWR.n5909 0.00975758
R13465 VPWR.n8820 VPWR.n347 0.00975758
R13466 VPWR.n8809 VPWR.n8808 0.00975758
R13467 VPWR.n8806 VPWR.n8805 0.00975758
R13468 VPWR.n8549 VPWR.n8522 0.00975758
R13469 VPWR.n8548 VPWR.n8547 0.00975758
R13470 VPWR.n8545 VPWR.n8544 0.00975758
R13471 VPWR.n6581 VPWR.n6321 0.00975758
R13472 VPWR.n6580 VPWR.n6579 0.00975758
R13473 VPWR.n6577 VPWR.n6576 0.00975758
R13474 VPWR.n8413 VPWR.n8363 0.00975758
R13475 VPWR.n8412 VPWR.n8411 0.00975758
R13476 VPWR.n8409 VPWR.n8408 0.00975758
R13477 VPWR.n5850 VPWR.n366 0.00975758
R13478 VPWR.n378 VPWR.n377 0.00975758
R13479 VPWR.n375 VPWR.n374 0.00975758
R13480 VPWR.n1068 VPWR.n1049 0.00975758
R13481 VPWR.n1067 VPWR.n1066 0.00975758
R13482 VPWR.n1064 VPWR.n1063 0.00975758
R13483 VPWR.n684 VPWR.n674 0.00975758
R13484 VPWR.n683 VPWR.n682 0.00975758
R13485 VPWR.n680 VPWR.n679 0.00975758
R13486 VPWR.n920 VPWR.n789 0.00975758
R13487 VPWR.n919 VPWR.n918 0.00975758
R13488 VPWR.n916 VPWR.n915 0.00975758
R13489 VPWR.n5731 VPWR.n5708 0.00975758
R13490 VPWR.n5720 VPWR.n5719 0.00975758
R13491 VPWR.n5717 VPWR.n5716 0.00975758
R13492 VPWR.n5550 VPWR.n481 0.00975758
R13493 VPWR.n5549 VPWR.n5548 0.00975758
R13494 VPWR.n5546 VPWR.n5545 0.00975758
R13495 VPWR.n1261 VPWR.n1237 0.00975758
R13496 VPWR.n1260 VPWR.n1259 0.00975758
R13497 VPWR.n1257 VPWR.n1256 0.00975758
R13498 VPWR.n5381 VPWR.n506 0.00975758
R13499 VPWR.n5383 VPWR.n5382 0.00975758
R13500 VPWR.n5386 VPWR.n5385 0.00975758
R13501 VPWR.n4620 VPWR.n4597 0.00975758
R13502 VPWR.n4609 VPWR.n4608 0.00975758
R13503 VPWR.n4606 VPWR.n4605 0.00975758
R13504 VPWR.n5241 VPWR.n1802 0.00975758
R13505 VPWR.n5240 VPWR.n5239 0.00975758
R13506 VPWR.n5237 VPWR.n5236 0.00975758
R13507 VPWR.n1618 VPWR.n565 0.00975758
R13508 VPWR.n1620 VPWR.n1619 0.00975758
R13509 VPWR.n1623 VPWR.n1622 0.00975758
R13510 VPWR.n5354 VPWR.n5330 0.00975758
R13511 VPWR.n5353 VPWR.n5352 0.00975758
R13512 VPWR.n5350 VPWR.n5349 0.00975758
R13513 VPWR.n4904 VPWR.n4881 0.00975758
R13514 VPWR.n4893 VPWR.n4892 0.00975758
R13515 VPWR.n4890 VPWR.n4889 0.00975758
R13516 VPWR.n5060 VPWR.n1863 0.00975758
R13517 VPWR.n5059 VPWR.n5058 0.00975758
R13518 VPWR.n5056 VPWR.n5055 0.00975758
R13519 VPWR.n2517 VPWR.n2194 0.00975758
R13520 VPWR.n2516 VPWR.n2515 0.00975758
R13521 VPWR.n2513 VPWR.n2512 0.00975758
R13522 VPWR.n5197 VPWR.n1808 0.00975758
R13523 VPWR.n5196 VPWR.n5195 0.00975758
R13524 VPWR.n5193 VPWR.n5192 0.00975758
R13525 VPWR.n2408 VPWR.n2198 0.00975758
R13526 VPWR.n2407 VPWR.n2406 0.00975758
R13527 VPWR.n2404 VPWR.n2403 0.00975758
R13528 VPWR.n2763 VPWR.n2738 0.00975758
R13529 VPWR.n2762 VPWR.n2761 0.00975758
R13530 VPWR.n2759 VPWR.n2758 0.00975758
R13531 VPWR.n4590 VPWR.n4577 0.00975758
R13532 VPWR.n4580 VPWR.n4579 0.00975758
R13533 VPWR.n1978 VPWR.n1977 0.00975758
R13534 VPWR.n1990 VPWR.n1980 0.00975758
R13535 VPWR.n2624 VPWR.n2600 0.00975758
R13536 VPWR.n2613 VPWR.n2612 0.00975758
R13537 VPWR.n2610 VPWR.n2609 0.00975758
R13538 VPWR.n7020 VPWR.n7004 0.00975758
R13539 VPWR.n7009 VPWR.n7008 0.00975758
R13540 VPWR.n7006 VPWR.n7005 0.00975758
R13541 VPWR.n5996 VPWR.n5995 0.00975758
R13542 VPWR.n4216 VPWR.n2878 0.00975758
R13543 VPWR.n4215 VPWR.n4214 0.00975758
R13544 VPWR.n2883 VPWR.n2882 0.00975758
R13545 VPWR.n3439 VPWR.n3438 0.00975758
R13546 VPWR.n3427 VPWR.n3426 0.00975758
R13547 VPWR.n3473 VPWR.n3472 0.00975758
R13548 VPWR.n3476 VPWR.n3475 0.00975758
R13549 VPWR.n4334 VPWR.n4321 0.00975758
R13550 VPWR.n4324 VPWR.n4323 0.00975758
R13551 VPWR.n2766 VPWR.n2765 0.00975758
R13552 VPWR.n2780 VPWR.n2768 0.00975758
R13553 VPWR.n3791 VPWR.n3777 0.00975758
R13554 VPWR.n3779 VPWR.n3778 0.00975758
R13555 VPWR.n3762 VPWR.n3761 0.00975758
R13556 VPWR.n3773 VPWR.n3772 0.00975758
R13557 VPWR.n3805 VPWR.n3804 0.00975758
R13558 VPWR.n3808 VPWR.n3807 0.00975758
R13559 VPWR.n3822 VPWR.n3821 0.00975758
R13560 VPWR.n6990 VPWR.n6974 0.00975758
R13561 VPWR.n6979 VPWR.n6978 0.00975758
R13562 VPWR.n6976 VPWR.n6975 0.00975758
R13563 VPWR.n6969 VPWR.n6968 0.00975758
R13564 VPWR.n3018 VPWR.n3017 0.00975758
R13565 VPWR.n3021 VPWR.n3020 0.00975758
R13566 VPWR.n3971 VPWR.n3970 0.00975758
R13567 VPWR.n8 VPWR.n7 0.00975758
R13568 VPWR.n10 VPWR.n9 0.00975758
R13569 VPWR.n13 VPWR.n12 0.00975758
R13570 VPWR.n15 VPWR.n14 0.00975758
R13571 VPWR.n9239 VPWR.n9238 0.00975758
R13572 VPWR.n9242 VPWR.n9241 0.00975758
R13573 VPWR.n9244 VPWR.n9243 0.00975758
R13574 VPWR.n7634 VPWR.n7617 0.00975758
R13575 VPWR.n7633 VPWR.n7632 0.00975758
R13576 VPWR.n7630 VPWR.n7629 0.00975758
R13577 VPWR.n7701 VPWR.n7700 0.00975758
R13578 VPWR.n6916 VPWR.n6899 0.00975758
R13579 VPWR.n6904 VPWR.n6903 0.00975758
R13580 VPWR.n6901 VPWR.n6900 0.00975758
R13581 VPWR.n6931 VPWR.n6930 0.00975758
R13582 VPWR.n3356 VPWR.n3333 0.00975758
R13583 VPWR.n3344 VPWR.n3343 0.00975758
R13584 VPWR.n3341 VPWR.n3340 0.00975758
R13585 VPWR.n4187 VPWR.n4186 0.00975758
R13586 VPWR.n4190 VPWR.n4189 0.00975758
R13587 VPWR.n4204 VPWR.n4203 0.00975758
R13588 VPWR.n7256 VPWR.n7255 0.00975758
R13589 VPWR.n7246 VPWR.n7245 0.00975758
R13590 VPWR.n7243 VPWR.n7242 0.00975758
R13591 VPWR.n7241 VPWR.n7232 0.00975758
R13592 VPWR.n6876 VPWR.n6874 0.00961458
R13593 VPWR.n7965 VPWR.n7964 0.00961458
R13594 VPWR.n8074 VPWR.n8073 0.00961458
R13595 VPWR.n9086 VPWR.n9084 0.00961458
R13596 VPWR.n260 VPWR.n200 0.00961458
R13597 VPWR.n273 VPWR.n272 0.00961458
R13598 VPWR.n6798 VPWR.n6796 0.00961458
R13599 VPWR.n6663 VPWR.n6662 0.00961458
R13600 VPWR.n8249 VPWR.n8248 0.00961458
R13601 VPWR.n8237 VPWR 0.00961458
R13602 VPWR.n8105 VPWR.n8104 0.00961458
R13603 VPWR.n8837 VPWR.n8835 0.00961458
R13604 VPWR.n8849 VPWR.n8848 0.00961458
R13605 VPWR.n6472 VPWR.n6469 0.00961458
R13606 VPWR.n6437 VPWR.n6436 0.00961458
R13607 VPWR.n8387 VPWR.n8386 0.00961458
R13608 VPWR.n8563 VPWR.n8562 0.00961458
R13609 VPWR VPWR.n8523 0.00961458
R13610 VPWR.n8539 VPWR.n8536 0.00961458
R13611 VPWR.n8715 VPWR.n8713 0.00961458
R13612 VPWR.n875 VPWR.n874 0.00961458
R13613 VPWR.n909 VPWR.n908 0.00961458
R13614 VPWR.n1082 VPWR.n1081 0.00961458
R13615 VPWR VPWR.n1042 0.00961458
R13616 VPWR.n5748 VPWR.n5746 0.00961458
R13617 VPWR.n1364 VPWR.n1362 0.00961458
R13618 VPWR.n1423 VPWR.n1421 0.00961458
R13619 VPWR.n5394 VPWR.n5393 0.00961458
R13620 VPWR.n5507 VPWR.n5506 0.00961458
R13621 VPWR.n5565 VPWR.n5564 0.00961458
R13622 VPWR.n5671 VPWR.n5669 0.00961458
R13623 VPWR.n5683 VPWR.n5682 0.00961458
R13624 VPWR.n1638 VPWR.n1636 0.00961458
R13625 VPWR.n1732 VPWR.n1731 0.00961458
R13626 VPWR.n5247 VPWR.n5246 0.00961458
R13627 VPWR.n4664 VPWR.n4663 0.00961458
R13628 VPWR.n4868 VPWR.n4867 0.00961458
R13629 VPWR.n4858 VPWR.n4857 0.00961458
R13630 VPWR.n2543 VPWR.n2540 0.00961458
R13631 VPWR.n2583 VPWR.n2581 0.00961458
R13632 VPWR.n5166 VPWR.n5165 0.00961458
R13633 VPWR.n5079 VPWR.n5078 0.00961458
R13634 VPWR.n1882 VPWR.n1881 0.00961458
R13635 VPWR.n2677 VPWR.n2675 0.00961458
R13636 VPWR.n2645 VPWR.n2644 0.00961458
R13637 VPWR.n4369 VPWR.n4368 0.00961458
R13638 VPWR.n4389 VPWR.n4388 0.00961458
R13639 VPWR.n4557 VPWR.n4556 0.00961458
R13640 VPWR.n3492 VPWR.n3490 0.00961458
R13641 VPWR.n3547 VPWR.n3545 0.00961458
R13642 VPWR.n3567 VPWR.n3566 0.00961458
R13643 VPWR.n4296 VPWR.n4295 0.00961458
R13644 VPWR.n4279 VPWR.n4276 0.00961458
R13645 VPWR.n4230 VPWR.n4228 0.00961458
R13646 VPWR.n2940 VPWR.n2939 0.00961458
R13647 VPWR.n7690 VPWR.n7688 0.00961458
R13648 VPWR.n7823 VPWR.n7820 0.00961458
R13649 VPWR.n7849 VPWR.n7848 0.00961458
R13650 VPWR.n9260 VPWR.n9259 0.00961458
R13651 VPWR.n9222 VPWR.n9220 0.00961458
R13652 VPWR.n131 VPWR.n130 0.00961458
R13653 VPWR.n3325 VPWR.n3323 0.00961458
R13654 VPWR.n3866 VPWR.n3864 0.00961458
R13655 VPWR.n3837 VPWR.n3836 0.00961458
R13656 VPWR.n3945 VPWR.n3944 0.00961458
R13657 VPWR.n3961 VPWR.n3960 0.00961458
R13658 VPWR.n4168 VPWR.n4166 0.00961458
R13659 VPWR.n4154 VPWR.n4153 0.00961458
R13660 VPWR.n7606 VPWR.n7604 0.00961458
R13661 VPWR.n7450 VPWR.n7448 0.00961458
R13662 VPWR.n7423 VPWR.n7422 0.00961458
R13663 VPWR.n7345 VPWR.n7344 0.00961458
R13664 VPWR.n7332 VPWR.n7327 0.00961458
R13665 VPWR.n7196 VPWR.n7132 0.00961458
R13666 VPWR.n7208 VPWR.n7207 0.00961458
R13667 VPWR.n3794 VPWR.n3793 0.00956852
R13668 VPWR.n3007 VPWR.n3006 0.00956852
R13669 VPWR.n3363 VPWR.n3362 0.00956852
R13670 VPWR.n4208 VPWR.n4207 0.00956852
R13671 VPWR.n3132 VPWR.n3130 0.00894595
R13672 VPWR.n3330 VPWR.n3329 0.00894595
R13673 VPWR.n9127 VPWR.n9126 0.00894595
R13674 VPWR.n146 VPWR.n145 0.00894595
R13675 VPWR.n9272 VPWR.n9266 0.00894595
R13676 VPWR.n9236 VPWR.n9232 0.00894595
R13677 VPWR.n9215 VPWR.n9214 0.00894595
R13678 VPWR.n8964 VPWR.n8963 0.00894595
R13679 VPWR.n297 VPWR.n296 0.00894595
R13680 VPWR.n8078 VPWR.n5960 0.00894595
R13681 VPWR.n9096 VPWR.n186 0.00894595
R13682 VPWR.n9078 VPWR.n9072 0.00894595
R13683 VPWR.n6205 VPWR.n6204 0.00894595
R13684 VPWR.n6868 VPWR.n6867 0.00894595
R13685 VPWR.n7890 VPWR.n7886 0.00894595
R13686 VPWR.n5975 VPWR.n5974 0.00894595
R13687 VPWR.n7969 VPWR.n7968 0.00894595
R13688 VPWR.n7960 VPWR.n7896 0.00894595
R13689 VPWR.n8828 VPWR.n8827 0.00894595
R13690 VPWR.n8918 VPWR.n8862 0.00894595
R13691 VPWR.n8089 VPWR.n5950 0.00894595
R13692 VPWR.n8224 VPWR.n8218 0.00894595
R13693 VPWR.n8209 VPWR.n8208 0.00894595
R13694 VPWR.n6830 VPWR.n6828 0.00894595
R13695 VPWR.n6790 VPWR.n6789 0.00894595
R13696 VPWR.n8357 VPWR.n8353 0.00894595
R13697 VPWR.n5894 VPWR.n5893 0.00894595
R13698 VPWR.n5907 VPWR.n5906 0.00894595
R13699 VPWR.n8345 VPWR.n8344 0.00894595
R13700 VPWR.n8702 VPWR.n8701 0.00894595
R13701 VPWR.n8790 VPWR.n8731 0.00894595
R13702 VPWR.n8578 VPWR.n8575 0.00894595
R13703 VPWR.n8550 VPWR.n8520 0.00894595
R13704 VPWR.n8587 VPWR.n8584 0.00894595
R13705 VPWR.n6549 VPWR.n6548 0.00894595
R13706 VPWR.n6464 VPWR.n6341 0.00894595
R13707 VPWR.n6433 VPWR.n6432 0.00894595
R13708 VPWR.n8367 VPWR.n8366 0.00894595
R13709 VPWR.n8406 VPWR.n8405 0.00894595
R13710 VPWR.n8419 VPWR.n8418 0.00894595
R13711 VPWR.n5739 VPWR.n5738 0.00894595
R13712 VPWR.n5830 VPWR.n5773 0.00894595
R13713 VPWR.n1096 VPWR.n1093 0.00894595
R13714 VPWR.n1069 VPWR.n1047 0.00894595
R13715 VPWR.n1105 VPWR.n1102 0.00894595
R13716 VPWR.n652 VPWR.n651 0.00894595
R13717 VPWR.n1231 VPWR.n1230 0.00894595
R13718 VPWR.n783 VPWR.n779 0.00894595
R13719 VPWR.n793 VPWR.n792 0.00894595
R13720 VPWR.n913 VPWR.n912 0.00894595
R13721 VPWR.n926 VPWR.n925 0.00894595
R13722 VPWR.n5661 VPWR.n5660 0.00894595
R13723 VPWR.n5703 VPWR.n5702 0.00894595
R13724 VPWR.n5519 VPWR.n5516 0.00894595
R13725 VPWR.n5551 VPWR.n479 0.00894595
R13726 VPWR.n5532 VPWR.n5531 0.00894595
R13727 VPWR.n1332 VPWR.n1331 0.00894595
R13728 VPWR.n1522 VPWR.n1521 0.00894595
R13729 VPWR.n5366 VPWR.n5362 0.00894595
R13730 VPWR.n510 VPWR.n509 0.00894595
R13731 VPWR.n5389 VPWR.n5388 0.00894595
R13732 VPWR.n5376 VPWR.n501 0.00894595
R13733 VPWR.n4874 VPWR.n4870 0.00894595
R13734 VPWR.n4629 VPWR.n4628 0.00894595
R13735 VPWR.n5210 VPWR.n1789 0.00894595
R13736 VPWR.n5243 VPWR.n5242 0.00894595
R13737 VPWR.n5223 VPWR.n5222 0.00894595
R13738 VPWR.n1612 VPWR.n1610 0.00894595
R13739 VPWR.n1536 VPWR.n561 0.00894595
R13740 VPWR.n1762 VPWR.n1761 0.00894595
R13741 VPWR.n5334 VPWR.n5333 0.00894595
R13742 VPWR.n5347 VPWR.n5346 0.00894595
R13743 VPWR.n5325 VPWR.n5324 0.00894595
R13744 VPWR.n4994 VPWR.n4993 0.00894595
R13745 VPWR.n4986 VPWR.n4985 0.00894595
R13746 VPWR.n1868 VPWR.n1854 0.00894595
R13747 VPWR.n5061 VPWR.n1861 0.00894595
R13748 VPWR.n5042 VPWR.n5041 0.00894595
R13749 VPWR.n2499 VPWR.n2497 0.00894595
R13750 VPWR.n2420 VPWR.n2190 0.00894595
R13751 VPWR.n2594 VPWR.n2590 0.00894595
R13752 VPWR.n5177 VPWR.n1811 0.00894595
R13753 VPWR.n5190 VPWR.n5189 0.00894595
R13754 VPWR.n1828 VPWR.n1827 0.00894595
R13755 VPWR.n2275 VPWR.n2274 0.00894595
R13756 VPWR.n2391 VPWR.n2390 0.00894595
R13757 VPWR.n4358 VPWR.n4357 0.00894595
R13758 VPWR.n2749 VPWR.n2743 0.00894595
R13759 VPWR.n4350 VPWR.n4349 0.00894595
R13760 VPWR.n4571 VPWR.n4567 0.00894595
R13761 VPWR.n1973 VPWR.n1972 0.00894595
R13762 VPWR.n2671 VPWR.n2040 0.00894595
R13763 VPWR.n2617 VPWR.n2616 0.00894595
R13764 VPWR.n2607 VPWR.n2606 0.00894595
R13765 VPWR.n2635 VPWR.n2634 0.00894595
R13766 VPWR.n5984 VPWR.n5980 0.00894595
R13767 VPWR.n7013 VPWR.n7012 0.00894595
R13768 VPWR.n5994 VPWR.n5993 0.00894595
R13769 VPWR.n7857 VPWR.n7856 0.00894595
R13770 VPWR.n2873 VPWR.n2865 0.00894595
R13771 VPWR.n2968 VPWR.n2967 0.00894595
R13772 VPWR.n3445 VPWR.n3444 0.00894595
R13773 VPWR.n3753 VPWR.n3752 0.00894595
R13774 VPWR.n4305 VPWR.n4302 0.00894595
R13775 VPWR.n4333 VPWR.n4329 0.00894595
R13776 VPWR.n4315 VPWR.n4314 0.00894595
R13777 VPWR.n3118 VPWR.n3115 0.00894595
R13778 VPWR.n3784 VPWR.n3783 0.00894595
R13779 VPWR.n3771 VPWR.n3770 0.00894595
R13780 VPWR.n3532 VPWR.n3531 0.00894595
R13781 VPWR.n3106 VPWR.n3101 0.00894595
R13782 VPWR.n3798 VPWR.n3797 0.00894595
R13783 VPWR.n3819 VPWR.n3818 0.00894595
R13784 VPWR.n3828 VPWR.n3827 0.00894595
R13785 VPWR.n6998 VPWR.n6994 0.00894595
R13786 VPWR.n6983 VPWR.n6982 0.00894595
R13787 VPWR.n6967 VPWR.n6966 0.00894595
R13788 VPWR.n7028 VPWR.n7027 0.00894595
R13789 VPWR.n3933 VPWR.n3932 0.00894595
R13790 VPWR.n3015 VPWR.n3011 0.00894595
R13791 VPWR.n3979 VPWR.n3976 0.00894595
R13792 VPWR.n7324 VPWR.n7323 0.00894595
R13793 VPWR.n7316 VPWR.n7315 0.00894595
R13794 VPWR.n9288 VPWR.n9285 0.00894595
R13795 VPWR.n7727 VPWR.n7725 0.00894595
R13796 VPWR.n7736 VPWR.n7735 0.00894595
R13797 VPWR.n6920 VPWR.n6918 0.00894595
R13798 VPWR.n7611 VPWR.n7610 0.00894595
R13799 VPWR.n4175 VPWR.n4170 0.00894595
R13800 VPWR.n2981 VPWR.n2980 0.00894595
R13801 VPWR.n7261 VPWR.n7260 0.00894595
R13802 VPWR.n7228 VPWR.n7227 0.00894595
R13803 VPWR.n3125 VPWR.n3124 0.00837842
R13804 VPWR.n2974 VPWR.n2973 0.00837842
R13805 VPWR.n2976 VPWR.n2975 0.00837842
R13806 VPWR.n7998 VPWR.n7997 0.0083125
R13807 VPWR VPWR.n7871 0.0083125
R13808 VPWR.n9069 VPWR.n9068 0.0083125
R13809 VPWR.n6681 VPWR.n6680 0.0083125
R13810 VPWR.n8376 VPWR.n8370 0.0083125
R13811 VPWR.n8591 VPWR 0.0083125
R13812 VPWR.n890 VPWR.n881 0.0083125
R13813 VPWR VPWR.n905 0.0083125
R13814 VPWR.n1414 VPWR.n1413 0.0083125
R13815 VPWR.n5574 VPWR.n5572 0.0083125
R13816 VPWR.n1749 VPWR.n1748 0.0083125
R13817 VPWR.n2585 VPWR.n1813 0.0083125
R13818 VPWR.n5038 VPWR.n5036 0.0083125
R13819 VPWR.n5033 VPWR 0.0083125
R13820 VPWR.n2666 VPWR.n2665 0.0083125
R13821 VPWR.n4398 VPWR.n4396 0.0083125
R13822 VPWR.n3555 VPWR.n3553 0.0083125
R13823 VPWR.n4270 VPWR.n4268 0.0083125
R13824 VPWR.n7832 VPWR.n7829 0.0083125
R13825 VPWR.n9211 VPWR.n9209 0.0083125
R13826 VPWR.n3857 VPWR.n3856 0.0083125
R13827 VPWR.n3985 VPWR.n3983 0.0083125
R13828 VPWR.n7441 VPWR.n7440 0.0083125
R13829 VPWR.n8204 VPWR.n8201 0.00757276
R13830 VPWR.n8593 VPWR.n8592 0.00757276
R13831 VPWR.n1109 VPWR.n734 0.00757276
R13832 VPWR.n4673 VPWR.n4672 0.00757276
R13833 VPWR.n7054 VPWR.n7053 0.00757276
R13834 VPWR.n8243 VPWR.n8240 0.00739914
R13835 VPWR.n9250 VPWR.n9249 0.00725676
R13836 VPWR.n9230 VPWR.n9229 0.00725676
R13837 VPWR.n9092 VPWR.n187 0.00725676
R13838 VPWR.n174 VPWR.n173 0.00725676
R13839 VPWR.n7982 VPWR.n7981 0.00725676
R13840 VPWR.n8220 VPWR.n8219 0.00725676
R13841 VPWR.n5955 VPWR.n5954 0.00725676
R13842 VPWR.n5896 VPWR.n5895 0.00725676
R13843 VPWR.n8554 VPWR.n8553 0.00725676
R13844 VPWR.n8541 VPWR.n8529 0.00725676
R13845 VPWR.n8395 VPWR.n8394 0.00725676
R13846 VPWR.n1074 VPWR.n1073 0.00725676
R13847 VPWR.n1060 VPWR.n1055 0.00725676
R13848 VPWR.n899 VPWR.n898 0.00725676
R13849 VPWR.n5556 VPWR.n5555 0.00725676
R13850 VPWR.n5542 VPWR.n5541 0.00725676
R13851 VPWR.n1403 VPWR.n1402 0.00725676
R13852 VPWR.n4655 VPWR.n4654 0.00725676
R13853 VPWR.n5233 VPWR.n5232 0.00725676
R13854 VPWR.n5336 VPWR.n5335 0.00725676
R13855 VPWR.n5066 VPWR.n5065 0.00725676
R13856 VPWR.n5052 VPWR.n5051 0.00725676
R13857 VPWR.n5179 VPWR.n5178 0.00725676
R13858 VPWR.n2745 VPWR.n2744 0.00725676
R13859 VPWR.n2755 VPWR.n2754 0.00725676
R13860 VPWR.n2619 VPWR.n2618 0.00725676
R13861 VPWR.n7015 VPWR.n7014 0.00725676
R13862 VPWR.n2770 VPWR.n2769 0.00725676
R13863 VPWR.n2778 VPWR.n2777 0.00725676
R13864 VPWR.n3786 VPWR.n3785 0.00725676
R13865 VPWR.n3810 VPWR.n3809 0.00725676
R13866 VPWR.n6985 VPWR.n6984 0.00725676
R13867 VPWR.n3023 VPWR.n3022 0.00725676
R13868 VPWR.n3967 VPWR.n3966 0.00725676
R13869 VPWR.n7311 VPWR.n7310 0.00725676
R13870 VPWR.n7305 VPWR.n7304 0.00725676
R13871 VPWR VPWR.n6882 0.00701042
R13872 VPWR.n7997 VPWR.n7987 0.00701042
R13873 VPWR VPWR.n9083 0.00701042
R13874 VPWR.n6680 VPWR.n6679 0.00701042
R13875 VPWR VPWR.n6465 0.00701042
R13876 VPWR.n8377 VPWR.n8376 0.00701042
R13877 VPWR VPWR.n8718 0.00701042
R13878 VPWR VPWR.n588 0.00701042
R13879 VPWR.n891 VPWR.n890 0.00701042
R13880 VPWR.n5759 VPWR 0.00701042
R13881 VPWR.n1413 VPWR.n1408 0.00701042
R13882 VPWR.n1391 VPWR 0.00701042
R13883 VPWR.n1630 VPWR 0.00701042
R13884 VPWR.n1748 VPWR.n1747 0.00701042
R13885 VPWR.n5176 VPWR.n1813 0.00701042
R13886 VPWR VPWR.n2398 0.00701042
R13887 VPWR.n2041 VPWR 0.00701042
R13888 VPWR.n2665 VPWR.n2660 0.00701042
R13889 VPWR.n3484 VPWR 0.00701042
R13890 VPWR.n3556 VPWR.n3555 0.00701042
R13891 VPWR.n2936 VPWR 0.00701042
R13892 VPWR VPWR.n7696 0.00701042
R13893 VPWR.n7833 VPWR.n7832 0.00701042
R13894 VPWR.n3856 VPWR.n3852 0.00701042
R13895 VPWR.n3963 VPWR 0.00701042
R13896 VPWR.n7440 VPWR.n7438 0.00701042
R13897 VPWR VPWR.n7326 0.00701042
R13898 VPWR.n2977 VPWR.n2976 0.00696227
R13899 VPWR.n8007 VPWR.n8006 0.00693178
R13900 VPWR.n6689 VPWR.n6688 0.00693178
R13901 VPWR.n1768 VPWR.n1767 0.00693178
R13902 VPWR.n3759 VPWR.n3125 0.00657697
R13903 VPWR.n2973 VPWR.n2782 0.00657697
R13904 VPWR.n2972 VPWR.n2971 0.00648266
R13905 VPWR.n3755 VPWR.n3365 0.00648266
R13906 VPWR.n4308 VPWR.n4307 0.00648266
R13907 VPWR.n4318 VPWR.n4317 0.00648266
R13908 VPWR.n3123 VPWR.n3122 0.00648266
R13909 VPWR.n161 VPWR.n152 0.00619697
R13910 VPWR.n9120 VPWR.n9107 0.00619697
R13911 VPWR.n314 VPWR.n313 0.00619697
R13912 VPWR.n8957 VPWR.n8945 0.00619697
R13913 VPWR.n9097 VPWR.n181 0.00619697
R13914 VPWR.n177 VPWR.n176 0.00619697
R13915 VPWR.n6892 VPWR.n6891 0.00619697
R13916 VPWR.n6887 VPWR.n6886 0.00619697
R13917 VPWR.n7976 VPWR.n7975 0.00619697
R13918 VPWR.n7971 VPWR.n7970 0.00619697
R13919 VPWR.n8940 VPWR.n330 0.00619697
R13920 VPWR.n326 VPWR.n325 0.00619697
R13921 VPWR.n8226 VPWR.n8225 0.00619697
R13922 VPWR.n8231 VPWR.n8230 0.00619697
R13923 VPWR.n6860 VPWR.n6859 0.00619697
R13924 VPWR.n6855 VPWR.n6854 0.00619697
R13925 VPWR.n5914 VPWR.n5913 0.00619697
R13926 VPWR.n5909 VPWR.n5908 0.00619697
R13927 VPWR.n8820 VPWR.n8809 0.00619697
R13928 VPWR.n8805 VPWR.n8804 0.00619697
R13929 VPWR.n8549 VPWR.n8548 0.00619697
R13930 VPWR.n8544 VPWR.n8543 0.00619697
R13931 VPWR.n6581 VPWR.n6580 0.00619697
R13932 VPWR.n6576 VPWR.n6575 0.00619697
R13933 VPWR.n8413 VPWR.n8412 0.00619697
R13934 VPWR.n8408 VPWR.n8407 0.00619697
R13935 VPWR.n5850 VPWR.n378 0.00619697
R13936 VPWR.n374 VPWR.n373 0.00619697
R13937 VPWR.n1068 VPWR.n1067 0.00619697
R13938 VPWR.n1063 VPWR.n1062 0.00619697
R13939 VPWR.n684 VPWR.n683 0.00619697
R13940 VPWR.n679 VPWR.n678 0.00619697
R13941 VPWR.n920 VPWR.n919 0.00619697
R13942 VPWR.n915 VPWR.n914 0.00619697
R13943 VPWR.n5731 VPWR.n5720 0.00619697
R13944 VPWR.n5716 VPWR.n5715 0.00619697
R13945 VPWR.n5550 VPWR.n5549 0.00619697
R13946 VPWR.n5545 VPWR.n5544 0.00619697
R13947 VPWR.n1261 VPWR.n1260 0.00619697
R13948 VPWR.n1256 VPWR.n1255 0.00619697
R13949 VPWR.n5382 VPWR.n5381 0.00619697
R13950 VPWR.n5387 VPWR.n5386 0.00619697
R13951 VPWR.n4620 VPWR.n4609 0.00619697
R13952 VPWR.n4605 VPWR.n4604 0.00619697
R13953 VPWR.n5241 VPWR.n5240 0.00619697
R13954 VPWR.n5236 VPWR.n5235 0.00619697
R13955 VPWR.n1619 VPWR.n1618 0.00619697
R13956 VPWR.n1624 VPWR.n1623 0.00619697
R13957 VPWR.n5354 VPWR.n5353 0.00619697
R13958 VPWR.n5349 VPWR.n5348 0.00619697
R13959 VPWR.n4904 VPWR.n4893 0.00619697
R13960 VPWR.n4889 VPWR.n4888 0.00619697
R13961 VPWR.n5060 VPWR.n5059 0.00619697
R13962 VPWR.n5055 VPWR.n5054 0.00619697
R13963 VPWR.n2517 VPWR.n2516 0.00619697
R13964 VPWR.n2512 VPWR.n2511 0.00619697
R13965 VPWR.n5197 VPWR.n5196 0.00619697
R13966 VPWR.n5192 VPWR.n5191 0.00619697
R13967 VPWR.n2408 VPWR.n2407 0.00619697
R13968 VPWR.n2403 VPWR.n2402 0.00619697
R13969 VPWR.n2763 VPWR.n2762 0.00619697
R13970 VPWR.n2758 VPWR.n2757 0.00619697
R13971 VPWR.n4590 VPWR.n4580 0.00619697
R13972 VPWR.n1990 VPWR.n1978 0.00619697
R13973 VPWR.n2624 VPWR.n2613 0.00619697
R13974 VPWR.n2609 VPWR.n2608 0.00619697
R13975 VPWR.n7020 VPWR.n7009 0.00619697
R13976 VPWR.n4216 VPWR.n4215 0.00619697
R13977 VPWR.n2883 VPWR.n2881 0.00619697
R13978 VPWR.n3438 VPWR.n3427 0.00619697
R13979 VPWR.n3476 VPWR.n3473 0.00619697
R13980 VPWR.n4334 VPWR.n4324 0.00619697
R13981 VPWR.n2780 VPWR.n2766 0.00619697
R13982 VPWR.n3791 VPWR.n3779 0.00619697
R13983 VPWR.n3773 VPWR.n3762 0.00619697
R13984 VPWR.n3804 VPWR.n3803 0.00619697
R13985 VPWR.n3822 VPWR.n3808 0.00619697
R13986 VPWR.n6990 VPWR.n6979 0.00619697
R13987 VPWR.n3017 VPWR.n3016 0.00619697
R13988 VPWR.n3971 VPWR.n3021 0.00619697
R13989 VPWR.n9 VPWR.n8 0.00619697
R13990 VPWR.n14 VPWR.n13 0.00619697
R13991 VPWR.n9238 VPWR.n9237 0.00619697
R13992 VPWR.n9244 VPWR.n9242 0.00619697
R13993 VPWR.n7634 VPWR.n7633 0.00619697
R13994 VPWR.n6916 VPWR.n6904 0.00619697
R13995 VPWR.n3356 VPWR.n3344 0.00619697
R13996 VPWR.n3340 VPWR.n3339 0.00619697
R13997 VPWR.n4186 VPWR.n4185 0.00619697
R13998 VPWR.n4204 VPWR.n4190 0.00619697
R13999 VPWR.n7255 VPWR.n7246 0.00619697
R14000 VPWR.n7242 VPWR.n7241 0.00619697
R14001 VPWR.n3364 VPWR.n3363 0.00590801
R14002 VPWR.n6883 VPWR 0.00570833
R14003 VPWR.n7984 VPWR.n7983 0.00570833
R14004 VPWR.n8076 VPWR 0.00570833
R14005 VPWR.n9091 VPWR.n9090 0.00570833
R14006 VPWR.n9087 VPWR.n9086 0.00570833
R14007 VPWR.n6676 VPWR.n6675 0.00570833
R14008 VPWR.n8238 VPWR.n8237 0.00570833
R14009 VPWR.n8104 VPWR.n8102 0.00570833
R14010 VPWR.n8106 VPWR 0.00570833
R14011 VPWR.n8393 VPWR.n8380 0.00570833
R14012 VPWR.n8523 VPWR.n8515 0.00570833
R14013 VPWR.n8540 VPWR.n8539 0.00570833
R14014 VPWR VPWR.n8535 0.00570833
R14015 VPWR.n700 VPWR 0.00570833
R14016 VPWR.n1229 VPWR 0.00570833
R14017 VPWR.n900 VPWR.n894 0.00570833
R14018 VPWR.n1075 VPWR.n1042 0.00570833
R14019 VPWR.n1059 VPWR.n1058 0.00570833
R14020 VPWR VPWR.n5758 0.00570833
R14021 VPWR.n1405 VPWR.n1404 0.00570833
R14022 VPWR.n5558 VPWR.n5557 0.00570833
R14023 VPWR.n5564 VPWR.n5561 0.00570833
R14024 VPWR VPWR.n1629 0.00570833
R14025 VPWR.n1744 VPWR.n1743 0.00570833
R14026 VPWR.n4657 VPWR.n4656 0.00570833
R14027 VPWR.n4663 VPWR.n4660 0.00570833
R14028 VPWR.n5173 VPWR.n5172 0.00570833
R14029 VPWR.n5067 VPWR.n1856 0.00570833
R14030 VPWR.n1881 VPWR.n1879 0.00570833
R14031 VPWR.n2399 VPWR 0.00570833
R14032 VPWR.n2657 VPWR.n2656 0.00570833
R14033 VPWR.n4383 VPWR.n4382 0.00570833
R14034 VPWR.n4388 VPWR.n4386 0.00570833
R14035 VPWR VPWR.n3483 0.00570833
R14036 VPWR.n3560 VPWR.n3559 0.00570833
R14037 VPWR.n4284 VPWR.n4283 0.00570833
R14038 VPWR.n4280 VPWR.n4279 0.00570833
R14039 VPWR VPWR.n2866 0.00570833
R14040 VPWR.n2948 VPWR 0.00570833
R14041 VPWR.n7705 VPWR 0.00570833
R14042 VPWR.n7837 VPWR.n7836 0.00570833
R14043 VPWR.n9251 VPWR.n9226 0.00570833
R14044 VPWR.n9223 VPWR.n9222 0.00570833
R14045 VPWR.n3849 VPWR.n3848 0.00570833
R14046 VPWR.n3953 VPWR.n3952 0.00570833
R14047 VPWR.n3960 VPWR.n3956 0.00570833
R14048 VPWR.n7435 VPWR.n7434 0.00570833
R14049 VPWR.n7337 VPWR.n7336 0.00570833
R14050 VPWR.n7333 VPWR.n7332 0.00570833
R14051 VPWR.n3758 VPWR.n3757 0.005649
R14052 VPWR.n3353 VPWR.n3352 0.00556757
R14053 VPWR.n9110 VPWR.n9109 0.00556757
R14054 VPWR.n9234 VPWR.n9233 0.00556757
R14055 VPWR.n9216 VPWR.n9215 0.00556757
R14056 VPWR.n9214 VPWR.n28 0.00556757
R14057 VPWR.n8947 VPWR.n8946 0.00556757
R14058 VPWR.n9094 VPWR.n9093 0.00556757
R14059 VPWR.n9081 VPWR.n189 0.00556757
R14060 VPWR.n9079 VPWR.n9078 0.00556757
R14061 VPWR.n9072 VPWR.n191 0.00556757
R14062 VPWR.n6149 VPWR.n6148 0.00556757
R14063 VPWR.n7886 VPWR.n7885 0.00556757
R14064 VPWR.n7890 VPWR.n7889 0.00556757
R14065 VPWR.n7865 VPWR.n7864 0.00556757
R14066 VPWR.n8829 VPWR.n8828 0.00556757
R14067 VPWR.n8222 VPWR.n8221 0.00556757
R14068 VPWR.n8096 VPWR.n8095 0.00556757
R14069 VPWR.n8209 VPWR.n8098 0.00556757
R14070 VPWR.n8208 VPWR.n8100 0.00556757
R14071 VPWR.n6845 VPWR.n6844 0.00556757
R14072 VPWR.n8353 VPWR.n8352 0.00556757
R14073 VPWR.n8357 VPWR.n8356 0.00556757
R14074 VPWR.n5902 VPWR.n5901 0.00556757
R14075 VPWR.n8555 VPWR.n8552 0.00556757
R14076 VPWR.n8533 VPWR.n8531 0.00556757
R14077 VPWR.n8584 VPWR.n357 0.00556757
R14078 VPWR.n8587 VPWR.n8586 0.00556757
R14079 VPWR.n6566 VPWR.n6565 0.00556757
R14080 VPWR.n6464 VPWR.n6463 0.00556757
R14081 VPWR.n6433 VPWR.n6425 0.00556757
R14082 VPWR.n6432 VPWR.n6428 0.00556757
R14083 VPWR.n8401 VPWR.n8400 0.00556757
R14084 VPWR.n5740 VPWR.n5739 0.00556757
R14085 VPWR.n1072 VPWR.n1071 0.00556757
R14086 VPWR.n740 VPWR.n739 0.00556757
R14087 VPWR.n1102 VPWR.n742 0.00556757
R14088 VPWR.n1105 VPWR.n1104 0.00556757
R14089 VPWR.n688 VPWR.n687 0.00556757
R14090 VPWR.n1230 VPWR.n586 0.00556757
R14091 VPWR.n779 VPWR.n778 0.00556757
R14092 VPWR.n783 VPWR.n782 0.00556757
R14093 VPWR.n796 VPWR.n795 0.00556757
R14094 VPWR.n5662 VPWR.n5661 0.00556757
R14095 VPWR.n5554 VPWR.n5553 0.00556757
R14096 VPWR.n5526 VPWR.n5525 0.00556757
R14097 VPWR.n5532 VPWR.n5528 0.00556757
R14098 VPWR.n5531 VPWR.n5530 0.00556757
R14099 VPWR.n1246 VPWR.n1245 0.00556757
R14100 VPWR.n1521 VPWR.n1520 0.00556757
R14101 VPWR.n5362 VPWR.n5361 0.00556757
R14102 VPWR.n5366 VPWR.n5365 0.00556757
R14103 VPWR.n503 VPWR.n502 0.00556757
R14104 VPWR.n4653 VPWR.n4649 0.00556757
R14105 VPWR.n5217 VPWR.n5216 0.00556757
R14106 VPWR.n5223 VPWR.n5219 0.00556757
R14107 VPWR.n5222 VPWR.n5221 0.00556757
R14108 VPWR.n574 VPWR.n573 0.00556757
R14109 VPWR.n1762 VPWR.n1754 0.00556757
R14110 VPWR.n1761 VPWR.n1757 0.00556757
R14111 VPWR.n5342 VPWR.n5341 0.00556757
R14112 VPWR.n4995 VPWR.n4994 0.00556757
R14113 VPWR.n5064 VPWR.n5063 0.00556757
R14114 VPWR.n1886 VPWR.n1884 0.00556757
R14115 VPWR.n5042 VPWR.n1874 0.00556757
R14116 VPWR.n5041 VPWR.n1876 0.00556757
R14117 VPWR.n2521 VPWR.n2520 0.00556757
R14118 VPWR.n2590 VPWR.n2112 0.00556757
R14119 VPWR.n2594 VPWR.n2593 0.00556757
R14120 VPWR.n5185 VPWR.n5184 0.00556757
R14121 VPWR.n2207 VPWR.n2206 0.00556757
R14122 VPWR.n2747 VPWR.n2746 0.00556757
R14123 VPWR.n4344 VPWR.n4343 0.00556757
R14124 VPWR.n4350 VPWR.n4346 0.00556757
R14125 VPWR.n4349 VPWR.n4348 0.00556757
R14126 VPWR.n1982 VPWR.n1981 0.00556757
R14127 VPWR.n2672 VPWR.n2671 0.00556757
R14128 VPWR.n2040 VPWR.n2039 0.00556757
R14129 VPWR.n2602 VPWR.n2601 0.00556757
R14130 VPWR.n5980 VPWR.n5979 0.00556757
R14131 VPWR.n5984 VPWR.n5983 0.00556757
R14132 VPWR.n5990 VPWR.n5989 0.00556757
R14133 VPWR.n2957 VPWR.n2949 0.00556757
R14134 VPWR.n3435 VPWR.n3434 0.00556757
R14135 VPWR.n3752 VPWR.n3369 0.00556757
R14136 VPWR.n4331 VPWR.n4330 0.00556757
R14137 VPWR.n2775 VPWR.n2774 0.00556757
R14138 VPWR.n4315 VPWR.n4311 0.00556757
R14139 VPWR.n4314 VPWR.n4313 0.00556757
R14140 VPWR.n3115 VPWR.n3114 0.00556757
R14141 VPWR.n3118 VPWR.n3117 0.00556757
R14142 VPWR.n3781 VPWR.n3780 0.00556757
R14143 VPWR.n3764 VPWR.n3763 0.00556757
R14144 VPWR.n3101 VPWR.n3100 0.00556757
R14145 VPWR.n3106 VPWR.n3105 0.00556757
R14146 VPWR.n3103 VPWR.n3102 0.00556757
R14147 VPWR.n3812 VPWR.n3811 0.00556757
R14148 VPWR.n6994 VPWR.n6993 0.00556757
R14149 VPWR.n6998 VPWR.n6997 0.00556757
R14150 VPWR.n6963 VPWR.n6962 0.00556757
R14151 VPWR.n3013 VPWR.n3012 0.00556757
R14152 VPWR.n3976 VPWR.n3002 0.00556757
R14153 VPWR.n3979 VPWR.n3978 0.00556757
R14154 VPWR.n7313 VPWR.n7312 0.00556757
R14155 VPWR.n7302 VPWR.n7301 0.00556757
R14156 VPWR.n9285 VPWR.n2 0.00556757
R14157 VPWR.n9288 VPWR.n9287 0.00556757
R14158 VPWR.n7626 VPWR.n7625 0.00556757
R14159 VPWR.n6913 VPWR.n6912 0.00556757
R14160 VPWR.n4194 VPWR.n4193 0.00556757
R14161 VPWR.n7236 VPWR.n7235 0.00556757
R14162 VPWR.n3128 VPWR.n3127 0.00554564
R14163 VPWR.n8006 VPWR.n8004 0.00548035
R14164 VPWR.n6688 VPWR.n6687 0.00548035
R14165 VPWR.n1767 VPWR.n1765 0.00548035
R14166 VPWR.n3006 VPWR.n2781 0.00500002
R14167 VPWR.n4336 VPWR.n4335 0.00500002
R14168 VPWR.n4211 VPWR.n2880 0.00500002
R14169 VPWR.n3793 VPWR.n3792 0.00495986
R14170 VPWR.n8205 VPWR.n8204 0.00484057
R14171 VPWR.n8593 VPWR.n8590 0.00484057
R14172 VPWR.n1109 VPWR.n1108 0.00484057
R14173 VPWR.n4672 VPWR.n4670 0.00484057
R14174 VPWR.n7053 VPWR.n7051 0.00484057
R14175 VPWR.n2876 VPWR.n2875 0.00477273
R14176 VPWR.n3442 VPWR.n3441 0.00477273
R14177 VPWR.n6991 VPWR.n6972 0.00460158
R14178 VPWR.n7022 VPWR.n7021 0.00460158
R14179 VPWR.n7863 VPWR.n7862 0.00460158
R14180 VPWR.n7880 VPWR.n5915 0.00460158
R14181 VPWR.n8414 VPWR.n8361 0.00460158
R14182 VPWR.n921 VPWR.n787 0.00460158
R14183 VPWR.n5380 VPWR.n512 0.00460158
R14184 VPWR.n5356 VPWR.n5355 0.00460158
R14185 VPWR.n5199 VPWR.n5198 0.00460158
R14186 VPWR.n2625 VPWR.n2598 0.00460158
R14187 VPWR.n3823 VPWR.n3795 0.00460158
R14188 VPWR.n19 VPWR.n18 0.00460158
R14189 VPWR.n2764 VPWR.n2736 0.00460158
R14190 VPWR.n3972 VPWR.n3008 0.00460158
R14191 VPWR.n6917 VPWR.n6897 0.00460158
R14192 VPWR.n7635 VPWR.n7615 0.00460158
R14193 VPWR.n6894 VPWR.n6893 0.00460158
R14194 VPWR.n6862 VPWR.n6861 0.00460158
R14195 VPWR.n6583 VPWR.n6582 0.00460158
R14196 VPWR.n677 VPWR.n676 0.00460158
R14197 VPWR.n1262 VPWR.n1235 0.00460158
R14198 VPWR.n1617 VPWR.n1526 0.00460158
R14199 VPWR.n2504 VPWR.n2195 0.00460158
R14200 VPWR.n2410 VPWR.n2409 0.00460158
R14201 VPWR.n7141 VPWR.n7136 0.00460158
R14202 VPWR.n7137 VPWR.n162 0.00460158
R14203 VPWR.n315 VPWR.n163 0.00460158
R14204 VPWR.n4206 VPWR.n4205 0.00460158
R14205 VPWR.n8958 VPWR.n8943 0.00460158
R14206 VPWR.n9121 VPWR.n9104 0.00460158
R14207 VPWR.n6215 VPWR.n6214 0.00440625
R14208 VPWR.n8003 VPWR.n8002 0.00440625
R14209 VPWR.n8000 VPWR.n7999 0.00440625
R14210 VPWR.n7868 VPWR.n5971 0.00440625
R14211 VPWR.n8069 VPWR.n8067 0.00440625
R14212 VPWR.n8064 VPWR.n188 0.00440625
R14213 VPWR.n9083 VPWR.n9082 0.00440625
R14214 VPWR.n9071 VPWR.n9070 0.00440625
R14215 VPWR.n279 VPWR.n278 0.00440625
R14216 VPWR VPWR.n294 0.00440625
R14217 VPWR.n6816 VPWR.n6815 0.00440625
R14218 VPWR.n6686 VPWR.n6685 0.00440625
R14219 VPWR.n6683 VPWR.n6682 0.00440625
R14220 VPWR.n6674 VPWR.n6673 0.00440625
R14221 VPWR.n8240 VPWR.n8239 0.00440625
R14222 VPWR.n8107 VPWR.n8106 0.00440625
R14223 VPWR.n8207 VPWR.n8206 0.00440625
R14224 VPWR.n339 VPWR.n336 0.00440625
R14225 VPWR.n8933 VPWR.n8932 0.00440625
R14226 VPWR.n8922 VPWR 0.00440625
R14227 VPWR.n6554 VPWR.n6328 0.00440625
R14228 VPWR.n6465 VPWR.n6329 0.00440625
R14229 VPWR.n6435 VPWR.n6434 0.00440625
R14230 VPWR.n8369 VPWR.n8368 0.00440625
R14231 VPWR.n8392 VPWR.n8391 0.00440625
R14232 VPWR.n8559 VPWR.n8558 0.00440625
R14233 VPWR.n8557 VPWR 0.00440625
R14234 VPWR.n8535 VPWR.n8534 0.00440625
R14235 VPWR.n8589 VPWR.n8588 0.00440625
R14236 VPWR.n8721 VPWR.n8719 0.00440625
R14237 VPWR.n667 VPWR.n666 0.00440625
R14238 VPWR.n1229 VPWR.n1228 0.00440625
R14239 VPWR.n877 VPWR.n876 0.00440625
R14240 VPWR.n880 VPWR.n879 0.00440625
R14241 VPWR.n902 VPWR.n901 0.00440625
R14242 VPWR.n1077 VPWR.n1076 0.00440625
R14243 VPWR.n737 VPWR.n736 0.00440625
R14244 VPWR.n1107 VPWR.n1106 0.00440625
R14245 VPWR.n388 VPWR.n381 0.00440625
R14246 VPWR.n5843 VPWR.n5842 0.00440625
R14247 VPWR.n1345 VPWR.n1344 0.00440625
R14248 VPWR.n1368 VPWR.n1367 0.00440625
R14249 VPWR.n1419 VPWR.n1418 0.00440625
R14250 VPWR.n1416 VPWR.n1415 0.00440625
R14251 VPWR.n1398 VPWR.n1397 0.00440625
R14252 VPWR.n5392 VPWR 0.00440625
R14253 VPWR.n5502 VPWR.n5500 0.00440625
R14254 VPWR.n5498 VPWR.n474 0.00440625
R14255 VPWR.n5567 VPWR.n5566 0.00440625
R14256 VPWR.n5570 VPWR.n5569 0.00440625
R14257 VPWR.n5667 VPWR.n5666 0.00440625
R14258 VPWR.n5690 VPWR.n5689 0.00440625
R14259 VPWR.n1597 VPWR.n1596 0.00440625
R14260 VPWR.n1764 VPWR.n1763 0.00440625
R14261 VPWR.n1751 VPWR.n1750 0.00440625
R14262 VPWR.n1742 VPWR.n1741 0.00440625
R14263 VPWR.n1793 VPWR.n1791 0.00440625
R14264 VPWR.n4652 VPWR.n4651 0.00440625
R14265 VPWR.n4666 VPWR.n4665 0.00440625
R14266 VPWR.n4669 VPWR.n4668 0.00440625
R14267 VPWR.n4852 VPWR.n4851 0.00440625
R14268 VPWR.n2483 VPWR.n2191 0.00440625
R14269 VPWR.n2587 VPWR.n2586 0.00440625
R14270 VPWR.n5171 VPWR.n5170 0.00440625
R14271 VPWR.n5074 VPWR.n5072 0.00440625
R14272 VPWR.n5070 VPWR.n5068 0.00440625
R14273 VPWR VPWR.n1883 0.00440625
R14274 VPWR.n5040 VPWR.n5039 0.00440625
R14275 VPWR.n5000 VPWR.n4999 0.00440625
R14276 VPWR.n4977 VPWR.n4976 0.00440625
R14277 VPWR.n2285 VPWR.n2284 0.00440625
R14278 VPWR.n2670 VPWR.n2041 0.00440625
R14279 VPWR.n2668 VPWR.n2667 0.00440625
R14280 VPWR.n2655 VPWR.n2654 0.00440625
R14281 VPWR.n4376 VPWR.n4374 0.00440625
R14282 VPWR.n4381 VPWR.n4380 0.00440625
R14283 VPWR.n4391 VPWR.n4390 0.00440625
R14284 VPWR.n4394 VPWR.n4393 0.00440625
R14285 VPWR.n4553 VPWR.n4552 0.00440625
R14286 VPWR.n3458 VPWR.n3457 0.00440625
R14287 VPWR.n3549 VPWR.n3548 0.00440625
R14288 VPWR.n3552 VPWR.n3551 0.00440625
R14289 VPWR.n3562 VPWR.n3561 0.00440625
R14290 VPWR.n4291 VPWR.n4289 0.00440625
R14291 VPWR.n4287 VPWR.n4285 0.00440625
R14292 VPWR.n4275 VPWR.n4274 0.00440625
R14293 VPWR.n4272 VPWR.n4271 0.00440625
R14294 VPWR.n2958 VPWR.n2948 0.00440625
R14295 VPWR.n7716 VPWR.n7715 0.00440625
R14296 VPWR.n7825 VPWR.n7824 0.00440625
R14297 VPWR.n7828 VPWR.n7827 0.00440625
R14298 VPWR.n7840 VPWR.n7838 0.00440625
R14299 VPWR.n9253 VPWR.n9252 0.00440625
R14300 VPWR.n9219 VPWR 0.00440625
R14301 VPWR.n9213 VPWR.n9212 0.00440625
R14302 VPWR.n125 VPWR.n124 0.00440625
R14303 VPWR.n3306 VPWR.n3305 0.00440625
R14304 VPWR.n3862 VPWR.n3861 0.00440625
R14305 VPWR.n3859 VPWR.n3858 0.00440625
R14306 VPWR.n3847 VPWR.n3846 0.00440625
R14307 VPWR.n3949 VPWR.n3948 0.00440625
R14308 VPWR.n3951 VPWR.n3950 0.00440625
R14309 VPWR.n3963 VPWR.n3962 0.00440625
R14310 VPWR.n3981 VPWR.n3980 0.00440625
R14311 VPWR.n4148 VPWR.n4147 0.00440625
R14312 VPWR.n7587 VPWR.n7586 0.00440625
R14313 VPWR.n7446 VPWR.n7445 0.00440625
R14314 VPWR.n7443 VPWR.n7442 0.00440625
R14315 VPWR.n7433 VPWR.n7432 0.00440625
R14316 VPWR.n7341 VPWR.n7340 0.00440625
R14317 VPWR.n7339 VPWR.n7338 0.00440625
R14318 VPWR.n7326 VPWR.n0 0.00440625
R14319 VPWR.n9289 VPWR.n1 0.00440625
R14320 VPWR.n7214 VPWR.n7213 0.00440625
R14321 VPWR VPWR.n7225 0.00440625
R14322 VPWR.n8079 VPWR.n5958 0.00406061
R14323 VPWR.n6866 VPWR.n6865 0.00406061
R14324 VPWR.n7891 VPWR.n7882 0.00406061
R14325 VPWR.n8826 VPWR.n344 0.00406061
R14326 VPWR.n8090 VPWR.n8085 0.00406061
R14327 VPWR.n6788 VPWR.n6787 0.00406061
R14328 VPWR.n8358 VPWR.n8349 0.00406061
R14329 VPWR.n8700 VPWR.n8696 0.00406061
R14330 VPWR.n8579 VPWR.n5858 0.00406061
R14331 VPWR.n6340 VPWR.n6339 0.00406061
R14332 VPWR.n6431 VPWR.n6429 0.00406061
R14333 VPWR.n5737 VPWR.n393 0.00406061
R14334 VPWR.n1097 VPWR.n748 0.00406061
R14335 VPWR.n1232 VPWR.n581 0.00406061
R14336 VPWR.n784 VPWR.n775 0.00406061
R14337 VPWR.n5659 VPWR.n5657 0.00406061
R14338 VPWR.n5520 VPWR.n484 0.00406061
R14339 VPWR.n1523 VPWR.n1267 0.00406061
R14340 VPWR.n5367 VPWR.n5358 0.00406061
R14341 VPWR.n4875 VPWR.n4633 0.00406061
R14342 VPWR.n5211 VPWR.n5206 0.00406061
R14343 VPWR.n1537 VPWR.n1531 0.00406061
R14344 VPWR.n1760 VPWR.n1758 0.00406061
R14345 VPWR.n4992 VPWR.n1969 0.00406061
R14346 VPWR.n1869 VPWR.n1864 0.00406061
R14347 VPWR.n2421 VPWR.n2415 0.00406061
R14348 VPWR.n2595 VPWR.n2109 0.00406061
R14349 VPWR.n2389 VPWR.n2388 0.00406061
R14350 VPWR.n4351 VPWR.n4342 0.00406061
R14351 VPWR.n2633 VPWR.n2632 0.00406061
R14352 VPWR.n7858 VPWR.n5999 0.00406061
R14353 VPWR.n2874 VPWR.n2870 0.00406061
R14354 VPWR.n2969 VPWR.n2884 0.00406061
R14355 VPWR.n3754 VPWR.n3366 0.00406061
R14356 VPWR.n4306 VPWR.n2783 0.00406061
R14357 VPWR.n4316 VPWR.n4309 0.00406061
R14358 VPWR.n3530 VPWR.n3529 0.00406061
R14359 VPWR.n3107 VPWR.n3095 0.00406061
R14360 VPWR.n7026 VPWR.n7025 0.00406061
R14361 VPWR.n3931 VPWR.n3927 0.00406061
R14362 VPWR.n9284 VPWR.n9283 0.00406061
R14363 VPWR.n24 VPWR.n23 0.00406061
R14364 VPWR.n7734 VPWR.n7733 0.00406061
R14365 VPWR.n7612 VPWR.n6934 0.00406061
R14366 VPWR.n3135 VPWR.n3129 0.00406061
R14367 VPWR.n4176 VPWR.n2985 0.00406061
R14368 VPWR.n7229 VPWR.n7142 0.00406061
R14369 VPWR.n7892 VPWR.n7881 0.00393497
R14370 VPWR.n8360 VPWR.n8359 0.00393497
R14371 VPWR.n5888 VPWR.n5887 0.00393497
R14372 VPWR.n785 VPWR.n774 0.00393497
R14373 VPWR.n5368 VPWR.n5357 0.00393497
R14374 VPWR.n514 VPWR.n513 0.00393497
R14375 VPWR.n2597 VPWR.n2596 0.00393497
R14376 VPWR.n7024 VPWR.n7023 0.00393497
R14377 VPWR.n3108 VPWR.n3094 0.00393497
R14378 VPWR.n7860 VPWR.n7859 0.00393497
R14379 VPWR.n2631 VPWR.n2630 0.00393497
R14380 VPWR.n165 VPWR.n25 0.00393497
R14381 VPWR.n9099 VPWR.n9098 0.00393497
R14382 VPWR.n8081 VPWR.n8080 0.00393497
R14383 VPWR.n8213 VPWR.n8082 0.00393497
R14384 VPWR.n8091 VPWR.n8084 0.00393497
R14385 VPWR.n8083 VPWR.n361 0.00393497
R14386 VPWR.n8580 VPWR.n5857 0.00393497
R14387 VPWR.n746 VPWR.n362 0.00393497
R14388 VPWR.n1098 VPWR.n747 0.00393497
R14389 VPWR.n5536 VPWR.n482 0.00393497
R14390 VPWR.n5521 VPWR.n483 0.00393497
R14391 VPWR.n5227 VPWR.n1803 0.00393497
R14392 VPWR.n5212 VPWR.n5205 0.00393497
R14393 VPWR.n5046 VPWR.n1804 0.00393497
R14394 VPWR.n2735 VPWR.n1870 0.00393497
R14395 VPWR.n4352 VPWR.n4338 0.00393497
R14396 VPWR.n9282 VPWR.n9281 0.00393497
R14397 VPWR.n3005 VPWR.n3004 0.00393497
R14398 VPWR.n9280 VPWR.n9279 0.00393497
R14399 VPWR.n7732 VPWR.n6896 0.00393497
R14400 VPWR.n6864 VPWR.n6863 0.00393497
R14401 VPWR.n6585 VPWR.n6584 0.00393497
R14402 VPWR.n6338 VPWR.n6337 0.00393497
R14403 VPWR.n1234 VPWR.n1233 0.00393497
R14404 VPWR.n1525 VPWR.n1524 0.00393497
R14405 VPWR.n1538 VPWR.n1527 0.00393497
R14406 VPWR.n2422 VPWR.n2411 0.00393497
R14407 VPWR.n2387 VPWR.n2386 0.00393497
R14408 VPWR.n3358 VPWR.n3357 0.00393497
R14409 VPWR.n7614 VPWR.n7613 0.00393497
R14410 VPWR.n3361 VPWR.n3360 0.00393497
R14411 VPWR.n8942 VPWR.n8941 0.00393497
R14412 VPWR.n8824 VPWR.n8823 0.00393497
R14413 VPWR.n8822 VPWR.n8821 0.00393497
R14414 VPWR.n8698 VPWR.n8697 0.00393497
R14415 VPWR.n5852 VPWR.n5851 0.00393497
R14416 VPWR.n5735 VPWR.n5734 0.00393497
R14417 VPWR.n5733 VPWR.n5732 0.00393497
R14418 VPWR.n4594 VPWR.n394 0.00393497
R14419 VPWR.n4621 VPWR.n4595 0.00393497
R14420 VPWR.n4877 VPWR.n4876 0.00393497
R14421 VPWR.n4905 VPWR.n4879 0.00393497
R14422 VPWR.n4990 VPWR.n4593 0.00393497
R14423 VPWR.n1991 VPWR.n1976 0.00393497
R14424 VPWR.n4177 VPWR.n2984 0.00393497
R14425 VPWR.n4592 VPWR.n4591 0.00393497
R14426 VPWR.n3346 VPWR.n3345 0.00387838
R14427 VPWR.n3349 VPWR.n3348 0.00387838
R14428 VPWR.n155 VPWR.n154 0.00387838
R14429 VPWR.n9116 VPWR.n9115 0.00387838
R14430 VPWR.n9113 VPWR.n9112 0.00387838
R14431 VPWR.n304 VPWR.n303 0.00387838
R14432 VPWR.n8953 VPWR.n8952 0.00387838
R14433 VPWR.n8950 VPWR.n8949 0.00387838
R14434 VPWR.n6142 VPWR.n6141 0.00387838
R14435 VPWR.n6145 VPWR.n6144 0.00387838
R14436 VPWR.n6155 VPWR.n6154 0.00387838
R14437 VPWR.n7959 VPWR.n7958 0.00387838
R14438 VPWR.n333 VPWR.n332 0.00387838
R14439 VPWR.n323 VPWR.n322 0.00387838
R14440 VPWR.n8855 VPWR.n8854 0.00387838
R14441 VPWR.n6838 VPWR.n6837 0.00387838
R14442 VPWR.n6841 VPWR.n6840 0.00387838
R14443 VPWR.n6851 VPWR.n6850 0.00387838
R14444 VPWR.n8812 VPWR.n8811 0.00387838
R14445 VPWR.n8802 VPWR.n8801 0.00387838
R14446 VPWR.n8724 VPWR.n8723 0.00387838
R14447 VPWR.n6323 VPWR.n6322 0.00387838
R14448 VPWR.n6326 VPWR.n6325 0.00387838
R14449 VPWR.n6572 VPWR.n6571 0.00387838
R14450 VPWR.n8421 VPWR.n8420 0.00387838
R14451 VPWR.n5756 VPWR.n5755 0.00387838
R14452 VPWR.n371 VPWR.n370 0.00387838
R14453 VPWR.n5766 VPWR.n5765 0.00387838
R14454 VPWR.n669 VPWR.n668 0.00387838
R14455 VPWR.n672 VPWR.n671 0.00387838
R14456 VPWR.n703 VPWR.n702 0.00387838
R14457 VPWR.n928 VPWR.n927 0.00387838
R14458 VPWR.n5723 VPWR.n5722 0.00387838
R14459 VPWR.n5713 VPWR.n5712 0.00387838
R14460 VPWR.n399 VPWR.n398 0.00387838
R14461 VPWR.n1239 VPWR.n1238 0.00387838
R14462 VPWR.n1242 VPWR.n1241 0.00387838
R14463 VPWR.n1252 VPWR.n1251 0.00387838
R14464 VPWR.n4612 VPWR.n4611 0.00387838
R14465 VPWR.n4602 VPWR.n4601 0.00387838
R14466 VPWR.n4626 VPWR.n4625 0.00387838
R14467 VPWR.n567 VPWR.n566 0.00387838
R14468 VPWR.n570 VPWR.n569 0.00387838
R14469 VPWR.n1627 VPWR.n1626 0.00387838
R14470 VPWR.n4896 VPWR.n4895 0.00387838
R14471 VPWR.n4886 VPWR.n4885 0.00387838
R14472 VPWR.n4910 VPWR.n4909 0.00387838
R14473 VPWR.n2487 VPWR.n2486 0.00387838
R14474 VPWR.n2488 VPWR.n2192 0.00387838
R14475 VPWR.n2508 VPWR.n2507 0.00387838
R14476 VPWR.n2200 VPWR.n2199 0.00387838
R14477 VPWR.n2203 VPWR.n2202 0.00387838
R14478 VPWR.n2213 VPWR.n2212 0.00387838
R14479 VPWR.n4583 VPWR.n4582 0.00387838
R14480 VPWR.n1988 VPWR.n1987 0.00387838
R14481 VPWR.n1985 VPWR.n1984 0.00387838
R14482 VPWR.n4220 VPWR.n4219 0.00387838
R14483 VPWR.n2954 VPWR.n2953 0.00387838
R14484 VPWR.n2951 VPWR.n2950 0.00387838
R14485 VPWR.n3430 VPWR.n3429 0.00387838
R14486 VPWR.n3433 VPWR.n3432 0.00387838
R14487 VPWR.n3481 VPWR.n3480 0.00387838
R14488 VPWR.n7619 VPWR.n7618 0.00387838
R14489 VPWR.n7622 VPWR.n7621 0.00387838
R14490 VPWR.n6906 VPWR.n6905 0.00387838
R14491 VPWR.n6909 VPWR.n6908 0.00387838
R14492 VPWR.n4180 VPWR.n4179 0.00387838
R14493 VPWR.n4200 VPWR.n4199 0.00387838
R14494 VPWR.n4197 VPWR.n4196 0.00387838
R14495 VPWR.n7250 VPWR.n7249 0.00387838
R14496 VPWR.n7239 VPWR.n7238 0.00387838
R14497 VPWR.n7145 VPWR.n7144 0.00387838
R14498 VPWR.n3443 VPWR.n3425 0.0033671
R14499 VPWR.n3119 VPWR.n3112 0.0033671
R14500 VPWR.n3774 VPWR.n3111 0.0032017
R14501 VPWR.n3111 VPWR.n3110 0.0032017
R14502 VPWR.n7139 VPWR.n7138 0.0032017
R14503 VPWR.n4210 VPWR.n4209 0.0032017
R14504 VPWR.n4209 VPWR.n4208 0.0032017
R14505 VPWR.n7140 VPWR.n7139 0.0032017
R14506 VPWR.n6209 VPWR.n6208 0.00310417
R14507 VPWR.n6210 VPWR.n6209 0.00310417
R14508 VPWR.n6213 VPWR.n6212 0.00310417
R14509 VPWR.n6882 VPWR.n6881 0.00310417
R14510 VPWR.n7870 VPWR.n7869 0.00310417
R14511 VPWR.n7966 VPWR 0.00310417
R14512 VPWR.n7897 VPWR.n7872 0.00310417
R14513 VPWR.n8062 VPWR.n8061 0.00310417
R14514 VPWR VPWR.n8075 0.00310417
R14515 VPWR.n9068 VPWR.n9067 0.00310417
R14516 VPWR.n268 VPWR.n267 0.00310417
R14517 VPWR.n276 VPWR.n273 0.00310417
R14518 VPWR.n281 VPWR.n280 0.00310417
R14519 VPWR.n287 VPWR.n286 0.00310417
R14520 VPWR.n6824 VPWR.n6823 0.00310417
R14521 VPWR.n6823 VPWR.n6822 0.00310417
R14522 VPWR.n6818 VPWR.n6817 0.00310417
R14523 VPWR.n6804 VPWR.n6803 0.00310417
R14524 VPWR.n8253 VPWR.n8252 0.00310417
R14525 VPWR.n8844 VPWR.n8843 0.00310417
R14526 VPWR.n8853 VPWR.n8849 0.00310417
R14527 VPWR.n8931 VPWR.n8930 0.00310417
R14528 VPWR.n8928 VPWR.n8924 0.00310417
R14529 VPWR.n6553 VPWR.n6552 0.00310417
R14530 VPWR.n6558 VPWR.n6553 0.00310417
R14531 VPWR.n6556 VPWR.n6555 0.00310417
R14532 VPWR.n6477 VPWR.n6476 0.00310417
R14533 VPWR.n6461 VPWR 0.00310417
R14534 VPWR.n8378 VPWR 0.00310417
R14535 VPWR.n8382 VPWR.n8381 0.00310417
R14536 VPWR.n8573 VPWR.n8566 0.00310417
R14537 VPWR.n8709 VPWR.n8708 0.00310417
R14538 VPWR.n8717 VPWR.n8715 0.00310417
R14539 VPWR.n8800 VPWR.n8722 0.00310417
R14540 VPWR.n8798 VPWR.n8796 0.00310417
R14541 VPWR.n654 VPWR 0.00310417
R14542 VPWR.n658 VPWR.n657 0.00310417
R14543 VPWR.n662 VPWR.n658 0.00310417
R14544 VPWR.n665 VPWR.n664 0.00310417
R14545 VPWR.n704 VPWR.n588 0.00310417
R14546 VPWR VPWR.n1226 0.00310417
R14547 VPWR.n904 VPWR.n903 0.00310417
R14548 VPWR.n910 VPWR 0.00310417
R14549 VPWR.n931 VPWR.n930 0.00310417
R14550 VPWR.n1091 VPWR.n1085 0.00310417
R14551 VPWR.n5758 VPWR.n5757 0.00310417
R14552 VPWR.n5841 VPWR.n5840 0.00310417
R14553 VPWR.n5838 VPWR.n5836 0.00310417
R14554 VPWR.n1338 VPWR.n1337 0.00310417
R14555 VPWR.n1340 VPWR.n1338 0.00310417
R14556 VPWR.n1343 VPWR.n1342 0.00310417
R14557 VPWR.n1356 VPWR.n1355 0.00310417
R14558 VPWR.n1518 VPWR 0.00310417
R14559 VPWR.n1395 VPWR.n1393 0.00310417
R14560 VPWR.n5514 VPWR.n5510 0.00310417
R14561 VPWR VPWR.n5508 0.00310417
R14562 VPWR.n5575 VPWR.n5574 0.00310417
R14563 VPWR.n5678 VPWR.n5677 0.00310417
R14564 VPWR.n5687 VPWR.n5683 0.00310417
R14565 VPWR.n5692 VPWR.n5691 0.00310417
R14566 VPWR.n5696 VPWR.n5695 0.00310417
R14567 VPWR.n1607 VPWR.n1606 0.00310417
R14568 VPWR.n1606 VPWR.n1605 0.00310417
R14569 VPWR.n1599 VPWR.n1598 0.00310417
R14570 VPWR.n1631 VPWR.n1630 0.00310417
R14571 VPWR.n1739 VPWR.n1737 0.00310417
R14572 VPWR.n5253 VPWR.n5250 0.00310417
R14573 VPWR VPWR.n5248 0.00310417
R14574 VPWR.n4863 VPWR.n4862 0.00310417
R14575 VPWR.n4857 VPWR.n4856 0.00310417
R14576 VPWR.n4850 VPWR.n4849 0.00310417
R14577 VPWR.n4847 VPWR.n4846 0.00310417
R14578 VPWR.n2494 VPWR.n2493 0.00310417
R14579 VPWR.n2493 VPWR.n2492 0.00310417
R14580 VPWR.n2485 VPWR.n2484 0.00310417
R14581 VPWR.n2535 VPWR.n2534 0.00310417
R14582 VPWR VPWR.n2584 0.00310417
R14583 VPWR.n5083 VPWR.n5082 0.00310417
R14584 VPWR VPWR.n5080 0.00310417
R14585 VPWR.n5036 VPWR.n5034 0.00310417
R14586 VPWR.n4969 VPWR.n4968 0.00310417
R14587 VPWR.n4979 VPWR.n4978 0.00310417
R14588 VPWR.n4982 VPWR.n4981 0.00310417
R14589 VPWR.n2280 VPWR.n2279 0.00310417
R14590 VPWR.n2283 VPWR.n2282 0.00310417
R14591 VPWR.n2398 VPWR.n2397 0.00310417
R14592 VPWR.n2652 VPWR.n2650 0.00310417
R14593 VPWR.n4365 VPWR.n4364 0.00310417
R14594 VPWR.n4399 VPWR.n4398 0.00310417
R14595 VPWR.n4561 VPWR.n4560 0.00310417
R14596 VPWR.n4556 VPWR.n4555 0.00310417
R14597 VPWR.n4551 VPWR.n4550 0.00310417
R14598 VPWR.n4548 VPWR.n4543 0.00310417
R14599 VPWR.n3449 VPWR.n3448 0.00310417
R14600 VPWR.n3453 VPWR.n3449 0.00310417
R14601 VPWR.n3456 VPWR.n3455 0.00310417
R14602 VPWR.n3485 VPWR.n3484 0.00310417
R14603 VPWR.n3751 VPWR 0.00310417
R14604 VPWR VPWR.n3748 0.00310417
R14605 VPWR.n4300 VPWR.n4299 0.00310417
R14606 VPWR.n4268 VPWR.n4266 0.00310417
R14607 VPWR.n4221 VPWR.n2866 0.00310417
R14608 VPWR.n2943 VPWR.n2940 0.00310417
R14609 VPWR.n2960 VPWR.n2959 0.00310417
R14610 VPWR.n2963 VPWR.n2962 0.00310417
R14611 VPWR.n7722 VPWR.n7721 0.00310417
R14612 VPWR.n7721 VPWR.n7720 0.00310417
R14613 VPWR.n7718 VPWR.n7717 0.00310417
R14614 VPWR.n7696 VPWR.n7695 0.00310417
R14615 VPWR.n7844 VPWR.n7842 0.00310417
R14616 VPWR.n9264 VPWR.n9263 0.00310417
R14617 VPWR VPWR.n9261 0.00310417
R14618 VPWR.n9209 VPWR.n9207 0.00310417
R14619 VPWR.n135 VPWR.n134 0.00310417
R14620 VPWR.n130 VPWR.n129 0.00310417
R14621 VPWR.n123 VPWR.n122 0.00310417
R14622 VPWR.n120 VPWR.n117 0.00310417
R14623 VPWR.n3297 VPWR.n3296 0.00310417
R14624 VPWR.n3301 VPWR.n3297 0.00310417
R14625 VPWR.n3304 VPWR.n3303 0.00310417
R14626 VPWR.n3317 VPWR.n3316 0.00310417
R14627 VPWR.n3844 VPWR.n3842 0.00310417
R14628 VPWR.n3941 VPWR.n3940 0.00310417
R14629 VPWR.n3986 VPWR.n3985 0.00310417
R14630 VPWR.n4159 VPWR.n4158 0.00310417
R14631 VPWR.n4153 VPWR.n4152 0.00310417
R14632 VPWR.n4146 VPWR.n4145 0.00310417
R14633 VPWR.n4143 VPWR.n4140 0.00310417
R14634 VPWR.n7580 VPWR.n7579 0.00310417
R14635 VPWR.n7582 VPWR.n7580 0.00310417
R14636 VPWR.n7585 VPWR.n7584 0.00310417
R14637 VPWR.n7598 VPWR.n7597 0.00310417
R14638 VPWR.n7430 VPWR.n7428 0.00310417
R14639 VPWR.n7349 VPWR.n7348 0.00310417
R14640 VPWR.n7203 VPWR.n7202 0.00310417
R14641 VPWR.n7211 VPWR.n7208 0.00310417
R14642 VPWR.n7216 VPWR.n7215 0.00310417
R14643 VPWR.n7222 VPWR.n7221 0.00310417
R14644 VPWR.n7002 VPWR.n6991 0.0028004
R14645 VPWR.n3824 VPWR.n3823 0.0028004
R14646 VPWR.n7021 VPWR.n5988 0.0028004
R14647 VPWR.n5198 VPWR.n1806 0.0028004
R14648 VPWR.n5355 VPWR.n5328 0.0028004
R14649 VPWR.n5380 VPWR.n5379 0.0028004
R14650 VPWR.n922 VPWR.n921 0.0028004
R14651 VPWR.n8415 VPWR.n8414 0.0028004
R14652 VPWR.n8348 VPWR.n5915 0.0028004
R14653 VPWR.n7893 VPWR.n7863 0.0028004
R14654 VPWR.n2629 VPWR.n2625 0.0028004
R14655 VPWR.n20 VPWR.n19 0.0028004
R14656 VPWR.n3973 VPWR.n3972 0.0028004
R14657 VPWR.n4353 VPWR.n2764 0.0028004
R14658 VPWR.n7731 VPWR.n7635 0.0028004
R14659 VPWR.n6893 VPWR.n6138 0.0028004
R14660 VPWR.n6861 VPWR.n6834 0.0028004
R14661 VPWR.n6582 VPWR.n6319 0.0028004
R14662 VPWR.n677 VPWR.n577 0.0028004
R14663 VPWR.n1263 VPWR.n1262 0.0028004
R14664 VPWR.n1617 VPWR.n1616 0.0028004
R14665 VPWR.n2504 VPWR.n2503 0.0028004
R14666 VPWR.n2409 VPWR.n2196 0.0028004
R14667 VPWR.n6924 VPWR.n6917 0.0028004
R14668 VPWR.n8959 VPWR.n8958 0.0028004
R14669 VPWR.n8959 VPWR.n315 0.0028004
R14670 VPWR.n9122 VPWR.n162 0.0028004
R14671 VPWR.n9122 VPWR.n9121 0.0028004
R14672 VPWR.n4205 VPWR.n4178 0.0028004
R14673 VPWR.n7141 VPWR.n7140 0.0028004
R14674 VPWR.n7259 VPWR.n7135 0.00277474
R14675 VPWR.n9125 VPWR.n9123 0.00251462
R14676 VPWR.n8962 VPWR.n8960 0.00251462
R14677 VPWR.n6203 VPWR.n6201 0.00251462
R14678 VPWR.n6833 VPWR.n6832 0.00251462
R14679 VPWR.n6547 VPWR.n6545 0.00251462
R14680 VPWR.n650 VPWR.n648 0.00251462
R14681 VPWR.n1330 VPWR.n1328 0.00251462
R14682 VPWR.n1615 VPWR.n1614 0.00251462
R14683 VPWR.n2502 VPWR.n2501 0.00251462
R14684 VPWR.n2273 VPWR.n2271 0.00251462
R14685 VPWR.n4356 VPWR.n4354 0.00251462
R14686 VPWR.n4574 VPWR.n4573 0.00251462
R14687 VPWR.n2628 VPWR.n2627 0.00251462
R14688 VPWR.n1826 VPWR.n1825 0.00251462
R14689 VPWR.n5327 VPWR.n5326 0.00251462
R14690 VPWR.n5378 VPWR.n5377 0.00251462
R14691 VPWR.n924 VPWR.n923 0.00251462
R14692 VPWR.n8417 VPWR.n8416 0.00251462
R14693 VPWR.n8347 VPWR.n8346 0.00251462
R14694 VPWR.n7895 VPWR.n7894 0.00251462
R14695 VPWR.n7730 VPWR.n7729 0.00251462
R14696 VPWR.n299 VPWR.n298 0.00251462
R14697 VPWR.n1975 VPWR.n1974 0.00251462
R14698 VPWR.n148 VPWR.n147 0.00251462
R14699 VPWR.n2983 VPWR.n2982 0.00251462
R14700 VPWR.n7024 VPWR.n7002 0.00246749
R14701 VPWR.n7859 VPWR.n5988 0.00246749
R14702 VPWR.n2631 VPWR.n2629 0.00246749
R14703 VPWR.n3824 VPWR.n3108 0.00246749
R14704 VPWR.n2596 VPWR.n1806 0.00246749
R14705 VPWR.n5328 VPWR.n514 0.00246749
R14706 VPWR.n5379 VPWR.n5368 0.00246749
R14707 VPWR.n922 VPWR.n785 0.00246749
R14708 VPWR.n8415 VPWR.n5888 0.00246749
R14709 VPWR.n8359 VPWR.n8348 0.00246749
R14710 VPWR.n7893 VPWR.n7892 0.00246749
R14711 VPWR.n9282 VPWR.n20 0.00246749
R14712 VPWR.n9279 VPWR.n9278 0.00246749
R14713 VPWR.n3973 VPWR.n3005 0.00246749
R14714 VPWR.n4353 VPWR.n4352 0.00246749
R14715 VPWR.n5045 VPWR.n1870 0.00246749
R14716 VPWR.n5226 VPWR.n5212 0.00246749
R14717 VPWR.n5535 VPWR.n5521 0.00246749
R14718 VPWR.n1099 VPWR.n1098 0.00246749
R14719 VPWR.n8581 VPWR.n8580 0.00246749
R14720 VPWR.n8212 VPWR.n8091 0.00246749
R14721 VPWR.n8080 VPWR.n166 0.00246749
R14722 VPWR.n5046 VPWR.n5045 0.00246749
R14723 VPWR.n5227 VPWR.n5226 0.00246749
R14724 VPWR.n5536 VPWR.n5535 0.00246749
R14725 VPWR.n1099 VPWR.n746 0.00246749
R14726 VPWR.n8581 VPWR.n361 0.00246749
R14727 VPWR.n8213 VPWR.n8212 0.00246749
R14728 VPWR.n9098 VPWR.n166 0.00246749
R14729 VPWR.n9278 VPWR.n25 0.00246749
R14730 VPWR.n7613 VPWR.n6924 0.00246749
R14731 VPWR.n3360 VPWR.n3359 0.00246749
R14732 VPWR.n7732 VPWR.n7731 0.00246749
R14733 VPWR.n6864 VPWR.n6138 0.00246749
R14734 VPWR.n6834 VPWR.n6585 0.00246749
R14735 VPWR.n6338 VPWR.n6319 0.00246749
R14736 VPWR.n1233 VPWR.n577 0.00246749
R14737 VPWR.n1524 VPWR.n1263 0.00246749
R14738 VPWR.n1616 VPWR.n1538 0.00246749
R14739 VPWR.n2503 VPWR.n2422 0.00246749
R14740 VPWR.n2387 VPWR.n2196 0.00246749
R14741 VPWR.n3359 VPWR.n3358 0.00246749
R14742 VPWR.n4591 VPWR.n4575 0.00246749
R14743 VPWR.n4178 VPWR.n4177 0.00246749
R14744 VPWR.n8824 VPWR.n316 0.00246749
R14745 VPWR.n8698 VPWR.n345 0.00246749
R14746 VPWR.n5735 VPWR.n364 0.00246749
R14747 VPWR.n5706 VPWR.n394 0.00246749
R14748 VPWR.n4876 VPWR.n4632 0.00246749
R14749 VPWR.n4990 VPWR.n4989 0.00246749
R14750 VPWR.n4989 VPWR.n4905 0.00246749
R14751 VPWR.n4632 VPWR.n4621 0.00246749
R14752 VPWR.n5732 VPWR.n5706 0.00246749
R14753 VPWR.n5851 VPWR.n364 0.00246749
R14754 VPWR.n8821 VPWR.n345 0.00246749
R14755 VPWR.n8941 VPWR.n316 0.00246749
R14756 VPWR.n4575 VPWR.n1991 0.00246749
R14757 VPWR.n5764 VPWR.n5763 0.00228056
R14758 VPWR.n4974 VPWR.n4973 0.00228056
R14759 VPWR.n9246 VPWR.n9245 0.00218919
R14760 VPWR.n175 VPWR.n171 0.00218919
R14761 VPWR.n7978 VPWR.n7977 0.00218919
R14762 VPWR.n7960 VPWR.n7959 0.00218919
R14763 VPWR.n8233 VPWR.n8232 0.00218919
R14764 VPWR.n5900 VPWR.n5899 0.00218919
R14765 VPWR.n8542 VPWR.n8527 0.00218919
R14766 VPWR.n8399 VPWR.n8398 0.00218919
R14767 VPWR.n8420 VPWR.n8419 0.00218919
R14768 VPWR.n1061 VPWR.n1053 0.00218919
R14769 VPWR.n895 VPWR.n794 0.00218919
R14770 VPWR.n927 VPWR.n926 0.00218919
R14771 VPWR.n5543 VPWR.n5539 0.00218919
R14772 VPWR.n1399 VPWR.n511 0.00218919
R14773 VPWR.n5234 VPWR.n5230 0.00218919
R14774 VPWR.n5340 VPWR.n5339 0.00218919
R14775 VPWR.n5053 VPWR.n5049 0.00218919
R14776 VPWR.n5183 VPWR.n5182 0.00218919
R14777 VPWR.n2756 VPWR.n2752 0.00218919
R14778 VPWR.n2623 VPWR.n2622 0.00218919
R14779 VPWR.n7019 VPWR.n7018 0.00218919
R14780 VPWR.n2779 VPWR.n2773 0.00218919
R14781 VPWR.n3790 VPWR.n3789 0.00218919
R14782 VPWR.n3802 VPWR.n3801 0.00218919
R14783 VPWR.n6989 VPWR.n6988 0.00218919
R14784 VPWR.n3968 VPWR.n3026 0.00218919
R14785 VPWR.n7307 VPWR.n7306 0.00218919
R14786 VPWR.n5987 VPWR.n5986 0.00218193
R14787 VPWR.n3826 VPWR.n3825 0.00218193
R14788 VPWR.n7001 VPWR.n7000 0.00218193
R14789 VPWR.n3975 VPWR.n3974 0.00218193
R14790 VPWR.n4 VPWR.n3 0.00218193
R14791 VPWR.n5044 VPWR.n5043 0.00218193
R14792 VPWR.n5225 VPWR.n5224 0.00218193
R14793 VPWR.n5534 VPWR.n5533 0.00218193
R14794 VPWR.n1101 VPWR.n1100 0.00218193
R14795 VPWR.n8583 VPWR.n8582 0.00218193
R14796 VPWR.n8211 VPWR.n8210 0.00218193
R14797 VPWR.n9077 VPWR.n9076 0.00218193
R14798 VPWR.n9277 VPWR.n9276 0.00218193
R14799 VPWR.n6923 VPWR.n6922 0.00218193
R14800 VPWR.n3332 VPWR.n3331 0.00218193
R14801 VPWR.n4988 VPWR.n4987 0.00218193
R14802 VPWR.n4631 VPWR.n4630 0.00218193
R14803 VPWR.n5705 VPWR.n5704 0.00218193
R14804 VPWR.n5772 VPWR.n5771 0.00218193
R14805 VPWR.n8730 VPWR.n8729 0.00218193
R14806 VPWR.n8861 VPWR.n8860 0.00218193
R14807 VPWR.n3110 VPWR.n3109 0.00211562
R14808 VPWR.n4337 VPWR.n4336 0.00211562
R14809 VPWR.n3127 VPWR.n3126 0.00211562
R14810 VPWR.n2880 VPWR.n2879 0.00211562
R14811 VPWR.n3756 VPWR.n3128 0.00185526
R14812 VPWR.n6221 VPWR.n6220 0.00180208
R14813 VPWR VPWR.n6224 0.00180208
R14814 VPWR.n7963 VPWR 0.00180208
R14815 VPWR.n7961 VPWR.n7872 0.00180208
R14816 VPWR VPWR.n7898 0.00180208
R14817 VPWR.n7956 VPWR 0.00180208
R14818 VPWR.n288 VPWR.n287 0.00180208
R14819 VPWR.n295 VPWR 0.00180208
R14820 VPWR.n6813 VPWR.n6809 0.00180208
R14821 VPWR.n6807 VPWR 0.00180208
R14822 VPWR.n6659 VPWR.n5923 0.00180208
R14823 VPWR.n8831 VPWR 0.00180208
R14824 VPWR.n8924 VPWR.n8923 0.00180208
R14825 VPWR.n8919 VPWR 0.00180208
R14826 VPWR.n6562 VPWR.n6482 0.00180208
R14827 VPWR.n6438 VPWR.n6437 0.00180208
R14828 VPWR.n8383 VPWR.n8382 0.00180208
R14829 VPWR.n8796 VPWR.n8795 0.00180208
R14830 VPWR.n8791 VPWR 0.00180208
R14831 VPWR.n696 VPWR.n695 0.00180208
R14832 VPWR VPWR.n699 0.00180208
R14833 VPWR.n874 VPWR.n873 0.00180208
R14834 VPWR.n907 VPWR 0.00180208
R14835 VPWR.n931 VPWR.n766 0.00180208
R14836 VPWR.n1076 VPWR 0.00180208
R14837 VPWR.n5742 VPWR 0.00180208
R14838 VPWR VPWR.n5752 0.00180208
R14839 VPWR.n5836 VPWR.n5835 0.00180208
R14840 VPWR.n5831 VPWR 0.00180208
R14841 VPWR.n1350 VPWR.n1349 0.00180208
R14842 VPWR.n1424 VPWR.n1423 0.00180208
R14843 VPWR VPWR.n5395 0.00180208
R14844 VPWR.n5399 VPWR.n5397 0.00180208
R14845 VPWR VPWR.n5664 0.00180208
R14846 VPWR.n5698 VPWR.n5696 0.00180208
R14847 VPWR.n1594 VPWR.n1590 0.00180208
R14848 VPWR.n1588 VPWR 0.00180208
R14849 VPWR.n1728 VPWR.n524 0.00180208
R14850 VPWR.n4652 VPWR 0.00180208
R14851 VPWR.n4846 VPWR.n4845 0.00180208
R14852 VPWR.n2528 VPWR.n2526 0.00180208
R14853 VPWR VPWR.n2532 0.00180208
R14854 VPWR.n2581 VPWR.n2579 0.00180208
R14855 VPWR.n2589 VPWR 0.00180208
R14856 VPWR VPWR.n5175 0.00180208
R14857 VPWR.n5162 VPWR.n5161 0.00180208
R14858 VPWR VPWR.n4997 0.00180208
R14859 VPWR VPWR.n2291 0.00180208
R14860 VPWR.n2678 VPWR.n2677 0.00180208
R14861 VPWR.n2641 VPWR.n2640 0.00180208
R14862 VPWR.n4543 VPWR.n4542 0.00180208
R14863 VPWR.n3463 VPWR.n3462 0.00180208
R14864 VPWR VPWR.n3466 0.00180208
R14865 VPWR VPWR.n3750 0.00180208
R14866 VPWR.n3545 VPWR.n3543 0.00180208
R14867 VPWR.n3572 VPWR.n3570 0.00180208
R14868 VPWR.n4224 VPWR 0.00180208
R14869 VPWR.n2964 VPWR.n2963 0.00180208
R14870 VPWR.n7713 VPWR.n7709 0.00180208
R14871 VPWR.n7707 VPWR 0.00180208
R14872 VPWR.n7820 VPWR.n7818 0.00180208
R14873 VPWR.n7854 VPWR.n7852 0.00180208
R14874 VPWR.n117 VPWR.n116 0.00180208
R14875 VPWR.n3311 VPWR.n3310 0.00180208
R14876 VPWR.n3867 VPWR.n3866 0.00180208
R14877 VPWR.n3833 VPWR.n3832 0.00180208
R14878 VPWR.n4140 VPWR.n4139 0.00180208
R14879 VPWR.n7592 VPWR.n7591 0.00180208
R14880 VPWR.n7451 VPWR.n7450 0.00180208
R14881 VPWR.n7419 VPWR.n7418 0.00180208
R14882 VPWR.n7223 VPWR.n7222 0.00180208
R14883 VPWR.n7226 VPWR 0.00180208
R14884 VPWR.n2289 VPWR.n2287 0.00164032
R14885 VPWR.n3756 VPWR.n3364 0.0014919
R14886 VPWR.n3792 VPWR.n3774 0.00144128
R14887 VPWR.n4335 VPWR.n4319 0.00140106
R14888 VPWR.n4319 VPWR.n2781 0.00140106
R14889 VPWR.n4211 VPWR.n4210 0.00140106
R14890 VGND.n3205 VGND.n3204 113628
R14891 VGND VGND.n1475 46632.3
R14892 VGND.n6977 VGND.n1475 46118.5
R14893 VGND.n6978 VGND.n1474 46118.5
R14894 VGND.n6978 VGND.n6977 46118.5
R14895 VGND.n8336 VGND.n308 46118.5
R14896 VGND.n1474 VGND.n308 46118.5
R14897 VGND.n8337 VGND.n307 46118.5
R14898 VGND.n8337 VGND.n8336 46118.5
R14899 VGND.n3206 VGND.n3202 46118.5
R14900 VGND.n3202 VGND.n307 46118.5
R14901 VGND.n3206 VGND.n3205 46118.5
R14902 VGND VGND.n5106 18975.6
R14903 VGND.n5105 VGND.n5104 18046.4
R14904 VGND.n5106 VGND.n5105 18046.4
R14905 VGND.n5103 VGND.n3984 18046.4
R14906 VGND.n5104 VGND.n5103 18046.4
R14907 VGND.n3983 VGND.n3982 18046.4
R14908 VGND.n3984 VGND.n3983 18046.4
R14909 VGND.n3981 VGND.n1862 18046.4
R14910 VGND.n3982 VGND.n3981 18046.4
R14911 VGND.n3204 VGND.n3203 18046.4
R14912 VGND.n3203 VGND.n1862 18046.4
R14913 VGND VGND.t1220 4888.89
R14914 VGND.t1220 VGND 4408.43
R14915 VGND.t1093 VGND 4408.43
R14916 VGND.t887 VGND 4408.43
R14917 VGND.t1003 VGND.t863 3877.39
R14918 VGND.t1554 VGND.t1484 3877.39
R14919 VGND VGND.t1000 3363.22
R14920 VGND.t1454 VGND 3346.36
R14921 VGND VGND.t1306 3337.93
R14922 VGND VGND.t1158 3337.93
R14923 VGND.n5811 VGND.t1045 3268.57
R14924 VGND.t1406 VGND 3186.58
R14925 VGND VGND.t851 3186.58
R14926 VGND.t1382 VGND 3175.65
R14927 VGND VGND.t970 3175.65
R14928 VGND.t1149 VGND.t1549 3101.92
R14929 VGND.t1084 VGND.t997 3101.92
R14930 VGND.t1036 VGND.t1102 3101.92
R14931 VGND.t857 VGND.t1528 3101.92
R14932 VGND.t988 VGND.t1297 3101.92
R14933 VGND.t1563 VGND.t875 3101.92
R14934 VGND.t869 VGND.t1318 3101.92
R14935 VGND VGND.t1382 2858.63
R14936 VGND VGND.t1406 2858.63
R14937 VGND.t851 VGND 2858.63
R14938 VGND.t970 VGND 2858.63
R14939 VGND.t1045 VGND 2858.63
R14940 VGND VGND.t958 2857.47
R14941 VGND.t872 VGND 2857.47
R14942 VGND VGND.t1346 2857.47
R14943 VGND VGND.t860 2857.47
R14944 VGND.t1018 VGND 2857.47
R14945 VGND VGND.t1051 2857.47
R14946 VGND.t1546 VGND 2857.47
R14947 VGND.t1087 VGND 2857.47
R14948 VGND.t1516 VGND 2570.88
R14949 VGND.t922 VGND 2570.88
R14950 VGND VGND.t1211 2562.45
R14951 VGND VGND.n2662 2469.73
R14952 VGND.t1152 VGND.t140 2377.01
R14953 VGND.t708 VGND.t1448 2343.29
R14954 VGND.t881 VGND.t1516 2326.44
R14955 VGND.t1429 VGND.t922 2326.44
R14956 VGND.n5812 VGND.t1578 2262.86
R14957 VGND VGND.t1536 2169.94
R14958 VGND VGND.t1033 2164.47
R14959 VGND.t2433 VGND.t1918 2149.43
R14960 VGND.t2399 VGND.t2198 2149.43
R14961 VGND.t297 VGND.t2056 2149.43
R14962 VGND.t2334 VGND.t2830 2149.43
R14963 VGND.t1587 VGND.t267 2149.43
R14964 VGND.t1868 VGND 2115.71
R14965 VGND.t2936 VGND.t2278 2107.28
R14966 VGND.t2229 VGND.t1349 2098.85
R14967 VGND.t1457 VGND.t1599 2098.85
R14968 VGND.t917 VGND.t2876 2098.85
R14969 VGND.t458 VGND.t866 2090.42
R14970 VGND.t2274 VGND 2090.42
R14971 VGND VGND.t881 2081.99
R14972 VGND.t934 VGND 2081.99
R14973 VGND.t552 VGND 2081.99
R14974 VGND VGND.t1012 2081.99
R14975 VGND VGND.t1429 2081.99
R14976 VGND.t1409 VGND 2081.99
R14977 VGND VGND.t1191 2081.99
R14978 VGND VGND.t1214 2081.99
R14979 VGND.t3025 VGND.t946 2027.83
R14980 VGND.t908 VGND.t2687 2022.99
R14981 VGND.t1270 VGND.t1994 2022.99
R14982 VGND.t848 VGND.t490 2022.99
R14983 VGND.t1237 VGND.t3244 2022.99
R14984 VGND.t1024 VGND.t2022 2022.99
R14985 VGND.t1030 VGND.t2154 2022.99
R14986 VGND.t3161 VGND.t1009 1963.98
R14987 VGND.t2538 VGND.t1146 1955.56
R14988 VGND.t1388 VGND.n8908 1938.7
R14989 VGND.t2350 VGND 1862.84
R14990 VGND.t2081 VGND 1854.41
R14991 VGND.t1033 VGND 1852.92
R14992 VGND.t1536 VGND 1852.92
R14993 VGND.t1578 VGND 1852.92
R14994 VGND VGND.t934 1795.4
R14995 VGND VGND.t1321 1795.4
R14996 VGND VGND.t1084 1795.4
R14997 VGND.t1102 VGND 1795.4
R14998 VGND VGND.t857 1795.4
R14999 VGND.t1297 VGND 1795.4
R15000 VGND.t875 VGND 1795.4
R15001 VGND VGND.t869 1795.4
R15002 VGND VGND.t1076 1786.97
R15003 VGND VGND.t1149 1786.97
R15004 VGND.t1131 VGND 1786.97
R15005 VGND.t1059 VGND 1786.97
R15006 VGND VGND.t1279 1786.97
R15007 VGND.t1173 VGND 1786.97
R15008 VGND VGND.t1015 1786.97
R15009 VGND VGND.t1309 1786.97
R15010 VGND.t1355 VGND.t1176 1760
R15011 VGND.t636 VGND.t2648 1753.26
R15012 VGND.t1984 VGND.t552 1753.26
R15013 VGND.t530 VGND.t165 1753.26
R15014 VGND.t2843 VGND.t2767 1753.26
R15015 VGND.t3205 VGND.t1940 1753.26
R15016 VGND.t266 VGND.t2732 1753.26
R15017 VGND.t748 VGND.t437 1753.26
R15018 VGND.t2763 VGND.t2935 1753.26
R15019 VGND.t1614 VGND.t2605 1753.26
R15020 VGND.t2673 VGND.t786 1719.54
R15021 VGND VGND.t1056 1702.68
R15022 VGND.t1394 VGND 1702.68
R15023 VGND.t931 VGND 1702.68
R15024 VGND.t1039 VGND 1694.25
R15025 VGND.t1140 VGND 1694.25
R15026 VGND VGND.n806 1677.39
R15027 VGND.n7812 VGND 1677.39
R15028 VGND VGND.t749 1677.39
R15029 VGND.n9181 VGND 1677.39
R15030 VGND.t3061 VGND.t3057 1618.39
R15031 VGND.t115 VGND.t1944 1618.39
R15032 VGND.t3133 VGND.t1194 1584.67
R15033 VGND.t175 VGND.t2661 1584.67
R15034 VGND.t2095 VGND.t580 1584.67
R15035 VGND.t1836 VGND.t2676 1584.67
R15036 VGND.t2383 VGND.t2598 1584.67
R15037 VGND.t428 VGND.t2378 1584.67
R15038 VGND.t3101 VGND.t99 1584.67
R15039 VGND.t2133 VGND.t791 1584.67
R15040 VGND.t2178 VGND.t2746 1584.67
R15041 VGND.t2363 VGND 1576.25
R15042 VGND.t2548 VGND 1559.39
R15043 VGND VGND.t117 1559.39
R15044 VGND.t958 VGND.t1454 1550.96
R15045 VGND.t1076 VGND.t872 1550.96
R15046 VGND.t1143 VGND.t1361 1550.96
R15047 VGND.t860 VGND.t1059 1550.96
R15048 VGND.t1306 VGND.t1225 1550.96
R15049 VGND.n8909 VGND.t1062 1550.96
R15050 VGND.t1015 VGND.t1285 1550.96
R15051 VGND.t1000 VGND.t1087 1550.96
R15052 VGND.t3011 VGND.t2878 1542.53
R15053 VGND.t1182 VGND.t1978 1534.1
R15054 VGND.t2085 VGND.t1070 1534.1
R15055 VGND.t798 VGND.t955 1534.1
R15056 VGND.t1081 VGND.t546 1475.1
R15057 VGND VGND.t2509 1441.38
R15058 VGND.n5106 VGND 1432.95
R15059 VGND.n5105 VGND 1432.95
R15060 VGND.n5104 VGND 1432.95
R15061 VGND.n5103 VGND 1432.95
R15062 VGND.n3984 VGND 1432.95
R15063 VGND.n3983 VGND 1432.95
R15064 VGND.n3982 VGND 1432.95
R15065 VGND.n3981 VGND 1432.95
R15066 VGND.n1862 VGND 1432.95
R15067 VGND.n3203 VGND 1432.95
R15068 VGND.n3204 VGND 1432.95
R15069 VGND.t482 VGND 1424.52
R15070 VGND.t1188 VGND 1424.52
R15071 VGND VGND.t854 1424.52
R15072 VGND.t1400 VGND 1424.52
R15073 VGND VGND.t1352 1407.66
R15074 VGND.t991 VGND 1407.66
R15075 VGND.t1134 VGND 1407.66
R15076 VGND VGND.t905 1407.66
R15077 VGND VGND.t896 1407.66
R15078 VGND VGND.t1415 1407.66
R15079 VGND.t1262 VGND 1407.66
R15080 VGND.t979 VGND 1407.66
R15081 VGND.t1367 VGND 1407.66
R15082 VGND.t1155 VGND 1407.66
R15083 VGND.t1048 VGND 1407.66
R15084 VGND VGND.t1114 1407.66
R15085 VGND.t408 VGND.t3086 1399.23
R15086 VGND.t1801 VGND.t2255 1399.23
R15087 VGND.t98 VGND.t1923 1399.23
R15088 VGND.t1507 VGND 1399.23
R15089 VGND.t2765 VGND.t2180 1399.23
R15090 VGND.t608 VGND.t1943 1399.23
R15091 VGND.t3125 VGND.t2968 1399.23
R15092 VGND.t1598 VGND 1390.8
R15093 VGND.n4661 VGND.t2231 1382.38
R15094 VGND.n7943 VGND.t1642 1382.38
R15095 VGND.t805 VGND.t2555 1365.52
R15096 VGND.t633 VGND 1357.09
R15097 VGND VGND.t2950 1355.53
R15098 VGND.t946 VGND 1350.06
R15099 VGND.t1927 VGND 1348.66
R15100 VGND VGND.t3039 1340.23
R15101 VGND.t2695 VGND.t1498 1331.8
R15102 VGND.t394 VGND.t1259 1323.37
R15103 VGND.t2217 VGND.t1228 1323.37
R15104 VGND.t1581 VGND 1314.94
R15105 VGND VGND.t976 1314.94
R15106 VGND VGND.t949 1306.51
R15107 VGND.t1531 VGND 1306.51
R15108 VGND VGND.t1234 1306.51
R15109 VGND.t1073 VGND 1306.51
R15110 VGND.t1549 VGND 1306.51
R15111 VGND.t3007 VGND 1306.51
R15112 VGND.t1321 VGND 1306.51
R15113 VGND.t1279 VGND 1306.51
R15114 VGND VGND.t1173 1306.51
R15115 VGND.t1225 VGND 1306.51
R15116 VGND.t997 VGND 1306.51
R15117 VGND VGND.t1036 1306.51
R15118 VGND VGND.t1152 1306.51
R15119 VGND.t1528 VGND 1306.51
R15120 VGND VGND.t988 1306.51
R15121 VGND VGND.t1563 1306.51
R15122 VGND.t1318 VGND 1306.51
R15123 VGND.t1309 VGND 1306.51
R15124 VGND VGND.t937 1306.51
R15125 VGND.t2176 VGND.t3183 1298.08
R15126 VGND.t3194 VGND 1289.66
R15127 VGND.t1501 VGND 1289.66
R15128 VGND.t2683 VGND 1289.66
R15129 VGND.t710 VGND.t2939 1289.66
R15130 VGND VGND.t1647 1289.66
R15131 VGND VGND.t2809 1289.66
R15132 VGND.t1108 VGND 1289.66
R15133 VGND.t609 VGND 1289.66
R15134 VGND.n5813 VGND.t1240 1257.14
R15135 VGND.t2650 VGND.t2476 1255.94
R15136 VGND.t550 VGND.t2492 1255.94
R15137 VGND.t1625 VGND.t242 1255.94
R15138 VGND.t2490 VGND.t2917 1255.94
R15139 VGND.t234 VGND.t542 1255.94
R15140 VGND.t2468 VGND.t2932 1255.94
R15141 VGND.t163 VGND.t254 1255.94
R15142 VGND.t1692 VGND.t3009 1255.94
R15143 VGND.t1938 VGND.t2805 1255.94
R15144 VGND.t627 VGND.t1829 1255.94
R15145 VGND.t1976 VGND.t2710 1255.94
R15146 VGND.t631 VGND.t2748 1255.94
R15147 VGND.t617 VGND.t2083 1255.94
R15148 VGND.t2797 VGND.t611 1255.94
R15149 VGND.t2768 VGND 1239.08
R15150 VGND VGND.t2338 1239.08
R15151 VGND.t878 VGND.t2271 1230.65
R15152 VGND VGND.t1768 1230.65
R15153 VGND.t449 VGND.t1481 1230.65
R15154 VGND.t1364 VGND.t3204 1230.65
R15155 VGND.t1777 VGND.t171 1230.65
R15156 VGND.t1358 VGND.t1990 1230.65
R15157 VGND.t2934 VGND.t1335 1230.65
R15158 VGND.t1330 VGND.t101 1230.65
R15159 VGND.t637 VGND.t925 1230.65
R15160 VGND.t133 VGND.t1185 1213.79
R15161 VGND.t444 VGND.t2336 1196.93
R15162 VGND.t389 VGND 1188.51
R15163 VGND.n9182 VGND.t2030 1188.51
R15164 VGND.n5102 VGND.t651 1180.08
R15165 VGND.t2893 VGND.t1315 1180.08
R15166 VGND.n3208 VGND.t2457 1180.08
R15167 VGND.n9178 VGND.t937 1163.22
R15168 VGND VGND.t1606 1137.93
R15169 VGND.t49 VGND 1137.93
R15170 VGND.t405 VGND.t222 1112.64
R15171 VGND.t226 VGND.t188 1112.64
R15172 VGND.t2054 VGND.t236 1112.64
R15173 VGND.t2609 VGND.t218 1112.64
R15174 VGND.t2881 VGND.t232 1112.64
R15175 VGND.t2615 VGND.t2817 1112.64
R15176 VGND.t2905 VGND.t2474 1112.64
R15177 VGND.t230 VGND.t2625 1112.64
R15178 VGND.t2795 VGND.t2341 1112.64
R15179 VGND.t755 VGND.t623 1112.64
R15180 VGND.t2702 VGND.t2328 1112.64
R15181 VGND.t2716 VGND.t512 1112.64
R15182 VGND.t2781 VGND.t2361 1112.64
R15183 VGND.t2913 VGND.t2712 1112.64
R15184 VGND.t2283 VGND.t2787 1112.64
R15185 VGND.t465 VGND.t629 1112.64
R15186 VGND.t1686 VGND.t2671 1104.21
R15187 VGND VGND.t2044 1104.21
R15188 VGND.t220 VGND 1095.79
R15189 VGND.t2789 VGND 1095.79
R15190 VGND.n5814 VGND 1087.7
R15191 VGND.t1851 VGND 1087.36
R15192 VGND VGND.t1710 1087.36
R15193 VGND VGND.t2437 1078.93
R15194 VGND.t1137 VGND.t2838 1078.93
R15195 VGND.t1904 VGND 1078.93
R15196 VGND VGND.t1706 1078.93
R15197 VGND.t2515 VGND.n78 1078.93
R15198 VGND VGND.t169 1078.93
R15199 VGND.t2052 VGND 1078.93
R15200 VGND.t155 VGND 1078.93
R15201 VGND.t2825 VGND 1078.93
R15202 VGND.t1913 VGND 1070.5
R15203 VGND VGND.t135 1070.5
R15204 VGND VGND.t2640 1062.07
R15205 VGND VGND.t496 1062.07
R15206 VGND.t2573 VGND.t2036 1062.07
R15207 VGND VGND.t181 1062.07
R15208 VGND.t2778 VGND 1053.64
R15209 VGND VGND.t2193 1053.64
R15210 VGND VGND.t2266 1053.64
R15211 VGND.t706 VGND 1045.21
R15212 VGND.t1167 VGND.t2851 1045.21
R15213 VGND.t538 VGND.t1117 1045.21
R15214 VGND.t546 VGND.t1688 1045.21
R15215 VGND.t712 VGND.t1678 1045.21
R15216 VGND VGND.t3037 1045.21
R15217 VGND.t2648 VGND 1036.78
R15218 VGND.t1898 VGND 1036.78
R15219 VGND.t2000 VGND 1036.78
R15220 VGND.t2646 VGND 1036.78
R15221 VGND VGND.t411 1036.78
R15222 VGND VGND.t2930 1036.78
R15223 VGND.t62 VGND 1036.78
R15224 VGND VGND.t782 1036.78
R15225 VGND VGND.t3186 1036.78
R15226 VGND.t2732 VGND 1036.78
R15227 VGND.t2566 VGND 1036.78
R15228 VGND.t1978 VGND 1036.78
R15229 VGND.t2629 VGND 1036.78
R15230 VGND VGND.t554 1036.78
R15231 VGND VGND.t2513 1036.78
R15232 VGND.t1961 VGND 1036.78
R15233 VGND.t2926 VGND 1036.78
R15234 VGND VGND.t1294 1036.78
R15235 VGND VGND.t609 1036.78
R15236 VGND VGND.t214 1028.35
R15237 VGND VGND.t544 1028.35
R15238 VGND VGND.t3079 1028.35
R15239 VGND.t2809 VGND 1028.35
R15240 VGND VGND.t2085 1028.35
R15241 VGND.t949 VGND 1019.92
R15242 VGND VGND.t1003 1019.92
R15243 VGND VGND.t1376 1019.92
R15244 VGND VGND.t1886 1019.92
R15245 VGND.t1105 VGND 1019.92
R15246 VGND.t2949 VGND.t1682 1019.92
R15247 VGND.t1191 VGND 1019.92
R15248 VGND.t1214 VGND 1019.92
R15249 VGND.t1051 VGND 1019.92
R15250 VGND.t1484 VGND 1019.92
R15251 VGND.t1273 VGND 1019.92
R15252 VGND VGND.t1343 1011.49
R15253 VGND VGND.t1409 1011.49
R15254 VGND.t3021 VGND.t2679 1011.49
R15255 VGND VGND.t1379 1011.49
R15256 VGND VGND.t301 1011.49
R15257 VGND.t1128 VGND 1011.49
R15258 VGND.n222 VGND.t86 1011.49
R15259 VGND.n3691 VGND.n3689 1010.52
R15260 VGND.t1525 VGND.t477 994.636
R15261 VGND.t137 VGND.t2582 994.636
R15262 VGND.t1584 VGND.t2270 994.636
R15263 VGND.t187 VGND 986.207
R15264 VGND VGND.t1818 986.207
R15265 VGND.t2771 VGND 969.35
R15266 VGND.t1991 VGND 969.35
R15267 VGND.t432 VGND.t1672 960.92
R15268 VGND.t1674 VGND.t3070 960.92
R15269 VGND.t216 VGND 952.49
R15270 VGND.t1253 VGND.t1854 944.062
R15271 VGND.t264 VGND.t1199 944.062
R15272 VGND VGND.t3221 935.633
R15273 VGND.t2435 VGND 935.633
R15274 VGND VGND.t2845 935.633
R15275 VGND VGND.t784 935.633
R15276 VGND VGND.t2636 935.633
R15277 VGND VGND.t2459 935.633
R15278 VGND.t2160 VGND.t1120 935.633
R15279 VGND VGND.t800 935.633
R15280 VGND VGND.n1624 927.203
R15281 VGND.t1733 VGND.t1501 927.203
R15282 VGND.n5098 VGND 927.203
R15283 VGND VGND.n7684 927.203
R15284 VGND VGND.n8335 927.203
R15285 VGND.t1911 VGND.t1951 927.203
R15286 VGND VGND.n181 927.203
R15287 VGND.t2517 VGND.n3201 927.203
R15288 VGND VGND.n2107 927.203
R15289 VGND.n9179 VGND 927.203
R15290 VGND VGND.t1566 923.727
R15291 VGND.t2497 VGND.t2527 918.774
R15292 VGND.t1373 VGND 918.774
R15293 VGND.t2869 VGND.t1947 918.774
R15294 VGND.n5337 VGND 918.774
R15295 VGND.t1352 VGND 918.774
R15296 VGND.t407 VGND.t1738 918.774
R15297 VGND.t2694 VGND.t2368 918.774
R15298 VGND.t1146 VGND 918.774
R15299 VGND.t2349 VGND.t1 918.774
R15300 VGND VGND.t1134 918.774
R15301 VGND.t2237 VGND.t2256 918.774
R15302 VGND.t2642 VGND.t2873 918.774
R15303 VGND.t1291 VGND 918.774
R15304 VGND.t1920 VGND.t754 918.774
R15305 VGND.t905 VGND 918.774
R15306 VGND.t2560 VGND.t1853 918.774
R15307 VGND.t1424 VGND 918.774
R15308 VGND.t896 VGND 918.774
R15309 VGND.t1415 VGND 918.774
R15310 VGND.t2832 VGND.t1975 918.774
R15311 VGND VGND.t1262 918.774
R15312 VGND VGND.t1507 918.774
R15313 VGND.t952 VGND 918.774
R15314 VGND VGND.t1575 918.774
R15315 VGND.t1009 VGND 918.774
R15316 VGND.t2943 VGND.t2006 918.774
R15317 VGND VGND.t1217 918.774
R15318 VGND VGND.t1367 918.774
R15319 VGND.t1062 VGND 918.774
R15320 VGND.t2766 VGND.t2456 918.774
R15321 VGND.n3032 VGND 918.774
R15322 VGND VGND.t1048 918.774
R15323 VGND.t1120 VGND 918.774
R15324 VGND.t854 VGND 918.774
R15325 VGND.t1114 VGND 918.774
R15326 VGND.t435 VGND.t2967 918.774
R15327 VGND VGND.t1400 918.774
R15328 VGND.t1246 VGND 912.795
R15329 VGND VGND.t1418 912.795
R15330 VGND VGND.t1442 912.795
R15331 VGND.t441 VGND.t2050 910.346
R15332 VGND.t2091 VGND.t396 910.346
R15333 VGND.t1243 VGND.t2572 901.917
R15334 VGND.t1185 VGND 901.917
R15335 VGND.t635 VGND.t2214 893.487
R15336 VGND.t961 VGND.t797 893.487
R15337 VGND.t265 VGND.t1791 885.058
R15338 VGND VGND.t190 885.058
R15339 VGND.t809 VGND.t2326 876.629
R15340 VGND.t2569 VGND.t30 876.629
R15341 VGND.t83 VGND.t144 876.629
R15342 VGND VGND.t3104 868.199
R15343 VGND.t2737 VGND.t1300 868.199
R15344 VGND.t902 VGND.t2026 868.199
R15345 VGND.t560 VGND.t3173 859.77
R15346 VGND.t2138 VGND 851.341
R15347 VGND.t2821 VGND.t3202 851.341
R15348 VGND.t3049 VGND.t82 851.341
R15349 VGND.t590 VGND.t3043 851.341
R15350 VGND VGND.t1355 847.206
R15351 VGND.t1240 VGND 847.206
R15352 VGND VGND.t3021 842.913
R15353 VGND.t2070 VGND.t1636 842.913
R15354 VGND.t2068 VGND.t1637 842.913
R15355 VGND.t1522 VGND.t393 842.913
R15356 VGND.t2636 VGND.t1823 842.913
R15357 VGND.t2393 VGND.t2970 842.913
R15358 VGND.t2754 VGND.t2869 834.484
R15359 VGND.t1966 VGND.t2657 834.484
R15360 VGND.t188 VGND.t407 834.484
R15361 VGND.t3104 VGND.t2694 834.484
R15362 VGND.t1 VGND.t694 834.484
R15363 VGND.t2256 VGND.t2054 834.484
R15364 VGND.t754 VGND.t1789 834.484
R15365 VGND.t1853 VGND.t2881 834.484
R15366 VGND.t1924 VGND.t2905 834.484
R15367 VGND.t2625 VGND.t2737 834.484
R15368 VGND.t2937 VGND.t928 834.484
R15369 VGND.t2341 VGND.t807 834.484
R15370 VGND.t1975 VGND.t755 834.484
R15371 VGND.t2328 VGND.t265 834.484
R15372 VGND.t1773 VGND.t3198 834.484
R15373 VGND.t1799 VGND.t3227 834.484
R15374 VGND.t2361 VGND.t2766 834.484
R15375 VGND.t1942 VGND.t2913 834.484
R15376 VGND.t1591 VGND.t734 834.484
R15377 VGND.t2967 VGND.t465 834.484
R15378 VGND.t2623 VGND.t3144 834.484
R15379 VGND.t1259 VGND.t1948 826.054
R15380 VGND.t1627 VGND.t471 826.054
R15381 VGND.t3121 VGND.t2306 826.054
R15382 VGND.t2299 VGND.t1027 826.054
R15383 VGND.t2981 VGND.t985 826.054
R15384 VGND.t576 VGND.t2616 826.054
R15385 VGND VGND.t186 826.054
R15386 VGND.t1256 VGND.t300 826.054
R15387 VGND.t1228 VGND.t3001 826.054
R15388 VGND.t1992 VGND.t80 817.625
R15389 VGND.t117 VGND.t173 817.625
R15390 VGND.t2865 VGND.t106 817.625
R15391 VGND.t1882 VGND.t381 817.625
R15392 VGND.t463 VGND.t647 817.625
R15393 VGND.t3097 VGND.t458 817.625
R15394 VGND.t2562 VGND.t123 817.625
R15395 VGND.t2486 VGND.t522 817.625
R15396 VGND.t3117 VGND.t2232 817.625
R15397 VGND.t2135 VGND.t2517 817.625
R15398 VGND.t2016 VGND.t2259 817.625
R15399 VGND.t2156 VGND.t2 817.625
R15400 VGND.t2242 VGND.t2191 817.625
R15401 VGND.t2221 VGND.t2971 817.625
R15402 VGND.t3192 VGND.t535 809.196
R15403 VGND.t2772 VGND.t532 809.196
R15404 VGND.t2496 VGND.t2530 809.196
R15405 VGND.t1947 VGND.t2650 809.196
R15406 VGND.t2868 VGND.t1946 809.196
R15407 VGND.t1738 VGND.t216 809.196
R15408 VGND.t1737 VGND.t408 809.196
R15409 VGND.t2368 VGND.t550 809.196
R15410 VGND.t179 VGND.t2277 809.196
R15411 VGND.t3221 VGND.t2237 809.196
R15412 VGND.t2255 VGND.t2236 809.196
R15413 VGND.t3211 VGND.t2915 809.196
R15414 VGND.t3177 VGND.t2560 809.196
R15415 VGND.t1854 VGND.t2557 809.196
R15416 VGND.t2209 VGND.t4 809.196
R15417 VGND.t2932 VGND.t2200 809.196
R15418 VGND.t2181 VGND.t163 809.196
R15419 VGND.t3013 VGND.t309 809.196
R15420 VGND.t213 VGND.t761 809.196
R15421 VGND.t2851 VGND.t2211 809.196
R15422 VGND.t300 VGND.t1938 809.196
R15423 VGND.t1974 VGND.t2829 809.196
R15424 VGND.t1796 VGND.t264 809.196
R15425 VGND.t50 VGND.t697 809.196
R15426 VGND.t3070 VGND.t499 809.196
R15427 VGND.t85 VGND.t2726 809.196
R15428 VGND.t2836 VGND.t207 809.196
R15429 VGND.t2513 VGND.t205 809.196
R15430 VGND.t2456 VGND.t2515 809.196
R15431 VGND.t2455 VGND.t2765 809.196
R15432 VGND.t2748 VGND.t270 809.196
R15433 VGND.t2089 VGND.t3111 809.196
R15434 VGND.t2618 VGND.t1108 809.196
R15435 VGND.t2628 VGND.t2535 809.196
R15436 VGND.t2459 VGND.t1643 809.196
R15437 VGND.t2027 VGND.t1646 809.196
R15438 VGND.t800 VGND.t435 809.196
R15439 VGND.t2968 VGND.t436 809.196
R15440 VGND.t2530 VGND.t3147 800.766
R15441 VGND.t1946 VGND.t394 800.766
R15442 VGND.t2437 VGND.t1737 800.766
R15443 VGND.t3240 VGND.t2352 800.766
R15444 VGND.t2236 VGND.t1904 800.766
R15445 VGND.t3250 VGND.t3053 800.766
R15446 VGND.t583 VGND.t8 800.766
R15447 VGND.t2557 VGND.t2081 800.766
R15448 VGND.t2197 VGND.t2399 800.766
R15449 VGND.t761 VGND.t2229 800.766
R15450 VGND.t2056 VGND.t299 800.766
R15451 VGND.t22 VGND.t2494 800.766
R15452 VGND.t2829 VGND.t2334 800.766
R15453 VGND.t2928 VGND.t1796 800.766
R15454 VGND.t2730 VGND.t3095 800.766
R15455 VGND.t96 VGND.t1911 800.766
R15456 VGND.t1706 VGND.t50 800.766
R15457 VGND.t749 VGND.t548 800.766
R15458 VGND VGND.t462 800.766
R15459 VGND.t2892 VGND.t2683 800.766
R15460 VGND.t3016 VGND.t765 800.766
R15461 VGND.t1599 VGND.t1933 800.766
R15462 VGND.t2876 VGND.t1907 800.766
R15463 VGND.t207 VGND.t1963 800.766
R15464 VGND.t169 VGND.t2455 800.766
R15465 VGND.t269 VGND.t1587 800.766
R15466 VGND.t2847 VGND.t2089 800.766
R15467 VGND.t2654 VGND.t159 800.766
R15468 VGND.t2535 VGND.t2052 800.766
R15469 VGND.t589 VGND.t2160 800.766
R15470 VGND.t92 VGND.t2272 800.766
R15471 VGND.t3135 VGND.t3165 800.766
R15472 VGND.t3167 VGND.t1327 800.766
R15473 VGND.t436 VGND.t2825 800.766
R15474 VGND.t196 VGND.t568 800.766
R15475 VGND.t566 VGND.t3074 800.766
R15476 VGND VGND.n1475 792.337
R15477 VGND.t128 VGND 792.337
R15478 VGND.n6977 VGND 792.337
R15479 VGND.t1880 VGND 792.337
R15480 VGND.t108 VGND.t2376 792.337
R15481 VGND.t1465 VGND.t2004 792.337
R15482 VGND VGND.n6978 792.337
R15483 VGND.t1870 VGND 792.337
R15484 VGND VGND.n1474 792.337
R15485 VGND VGND.n308 792.337
R15486 VGND.t2189 VGND 792.337
R15487 VGND.n8336 VGND 792.337
R15488 VGND.t2172 VGND 792.337
R15489 VGND.t1303 VGND.t183 792.337
R15490 VGND VGND.n8337 792.337
R15491 VGND.t437 VGND.t1370 792.337
R15492 VGND VGND.t3159 792.337
R15493 VGND.n307 VGND 792.337
R15494 VGND.t1006 VGND.t2763 792.337
R15495 VGND VGND.t3066 792.337
R15496 VGND.t2090 VGND.t142 792.337
R15497 VGND.t469 VGND.t2090 792.337
R15498 VGND.n3202 VGND 792.337
R15499 VGND VGND.t1860 792.337
R15500 VGND VGND.n3206 792.337
R15501 VGND.t2855 VGND 792.337
R15502 VGND.n3205 VGND 792.337
R15503 VGND.t460 VGND 783.909
R15504 VGND.t1623 VGND.t3016 783.909
R15505 VGND.t2232 VGND 783.909
R15506 VGND.t1042 VGND.n6629 775.48
R15507 VGND.t1211 VGND.t1531 775.48
R15508 VGND.t2326 VGND.t597 775.48
R15509 VGND.t1902 VGND.t593 775.48
R15510 VGND.t1982 VGND.t2299 775.48
R15511 VGND.t2004 VGND.t2759 775.48
R15512 VGND.t1448 VGND.t1073 775.48
R15513 VGND.t2291 VGND.t380 775.48
R15514 VGND.t744 VGND.t2981 775.48
R15515 VGND.t2374 VGND.t706 775.48
R15516 VGND.n7311 VGND.t1276 775.48
R15517 VGND.t167 VGND.n8253 775.48
R15518 VGND.t1421 VGND.t1131 775.48
R15519 VGND.t1379 VGND.t1231 775.48
R15520 VGND.t1831 VGND.t2986 775.48
R15521 VGND.t2874 VGND.t2389 775.48
R15522 VGND.t2887 VGND.t2387 775.48
R15523 VGND.t1823 VGND.t2178 775.48
R15524 VGND.t43 VGND.t1827 775.48
R15525 VGND.t1769 VGND.t2393 775.48
R15526 VGND.t1699 VGND.n5107 770.683
R15527 VGND VGND.t2548 767.051
R15528 VGND.t224 VGND.t2780 767.051
R15529 VGND.t242 VGND.t2837 767.051
R15530 VGND.t1768 VGND.t2490 767.051
R15531 VGND.t477 VGND.t2468 767.051
R15532 VGND.t254 VGND.t530 767.051
R15533 VGND.t2767 VGND.t2480 767.051
R15534 VGND.t2706 VGND.t266 767.051
R15535 VGND.t1487 VGND.t2892 767.051
R15536 VGND.t2710 VGND.t2263 767.051
R15537 VGND.t2270 VGND.t631 767.051
R15538 VGND.t1937 VGND.t617 767.051
R15539 VGND.t54 VGND.t2240 767.051
R15540 VGND.t2966 VGND.t615 767.051
R15541 VGND.t625 VGND.t1614 767.051
R15542 VGND VGND.t691 758.621
R15543 VGND.t378 VGND.t452 758.621
R15544 VGND.t1027 VGND.t2024 758.621
R15545 VGND.t751 VGND 758.621
R15546 VGND.t985 VGND.t1721 758.621
R15547 VGND.t2930 VGND.t1525 758.621
R15548 VGND.t928 VGND.t428 758.621
R15549 VGND.t890 VGND.t3062 758.621
R15550 VGND.t2746 VGND.t1584 758.621
R15551 VGND VGND.t570 750.192
R15552 VGND.t2093 VGND.t899 750.192
R15553 VGND.t181 VGND.t2504 750.192
R15554 VGND.t3114 VGND.t3051 750.192
R15555 VGND.t1621 VGND.t47 741.763
R15556 VGND.t194 VGND.t2034 741.763
R15557 VGND.t597 VGND.t1988 741.763
R15558 VGND.t3106 VGND.t2000 741.763
R15559 VGND.t2498 VGND.t1862 741.763
R15560 VGND.t2859 VGND.t2646 741.763
R15561 VGND.t1739 VGND.t1653 741.763
R15562 VGND.t544 VGND.t1743 741.763
R15563 VGND.t2674 VGND.t2002 741.763
R15564 VGND.t3079 VGND.t585 741.763
R15565 VGND.t1934 VGND.t789 741.763
R15566 VGND.t578 VGND.t478 741.763
R15567 VGND.t1797 VGND.t2629 741.763
R15568 VGND.t554 VGND.t1840 741.763
R15569 VGND.t2207 VGND.t2926 741.763
R15570 VGND.t2046 VGND.t1593 733.333
R15571 VGND.t2995 VGND.t403 733.333
R15572 VGND.t2861 VGND.t514 733.333
R15573 VGND.t2576 VGND.t2885 733.333
R15574 VGND.t380 VGND.t2293 733.333
R15575 VGND.t638 VGND.t572 733.333
R15576 VGND.t2691 VGND.t2685 724.904
R15577 VGND.t41 VGND.t2842 724.904
R15578 VGND.t1994 VGND.t1996 724.904
R15579 VGND.t1996 VGND.t1998 724.904
R15580 VGND.t1998 VGND.t1992 724.904
R15581 VGND.t813 VGND.t815 724.904
R15582 VGND.t2421 VGND.t2907 724.904
R15583 VGND.t2425 VGND.t2419 724.904
R15584 VGND.t2403 VGND.t2401 724.904
R15585 VGND.t2407 VGND.t2405 724.904
R15586 VGND.t2409 VGND.t2407 724.904
R15587 VGND.t180 VGND.t1324 724.904
R15588 VGND.t457 VGND.t383 724.904
R15589 VGND.t1179 VGND.t1920 724.904
R15590 VGND.t2166 VGND.t2168 724.904
R15591 VGND.t2168 VGND.t2162 724.904
R15592 VGND.t2250 VGND.t2252 724.904
R15593 VGND.t1462 VGND.t584 724.904
R15594 VGND.t1729 VGND.t772 724.904
R15595 VGND.t494 VGND.t488 724.904
R15596 VGND.t2111 VGND.t2113 724.904
R15597 VGND.t2101 VGND.t2107 724.904
R15598 VGND.t2129 VGND.t340 724.904
R15599 VGND.t340 VGND.t328 724.904
R15600 VGND.t328 VGND.t332 724.904
R15601 VGND.t332 VGND.t338 724.904
R15602 VGND.t334 VGND.t314 724.904
R15603 VGND.t659 VGND.t653 724.904
R15604 VGND.t653 VGND.t663 724.904
R15605 VGND.t681 VGND.t675 724.904
R15606 VGND.t677 VGND.t679 724.904
R15607 VGND.t679 VGND.t683 724.904
R15608 VGND.t683 VGND.t655 724.904
R15609 VGND.t657 VGND.t661 724.904
R15610 VGND.t2990 VGND.t3099 724.904
R15611 VGND VGND.t2484 724.904
R15612 VGND.t2523 VGND.t2525 724.904
R15613 VGND.t2525 VGND.t2519 724.904
R15614 VGND.t804 VGND.t2937 724.904
R15615 VGND VGND.t838 724.904
R15616 VGND.t838 VGND.t831 724.904
R15617 VGND.t827 VGND.t821 724.904
R15618 VGND.t833 VGND.t825 724.904
R15619 VGND.t2304 VGND.t2302 724.904
R15620 VGND.t342 VGND.t330 724.904
R15621 VGND.t344 VGND.t348 724.904
R15622 VGND.t348 VGND.t352 724.904
R15623 VGND.t356 VGND.t358 724.904
R15624 VGND.t358 VGND.t360 724.904
R15625 VGND.t360 VGND.t364 724.904
R15626 VGND.t370 VGND.t374 724.904
R15627 VGND.t524 VGND.t518 724.904
R15628 VGND.t518 VGND.t520 724.904
R15629 VGND.t1778 VGND.t1631 724.904
R15630 VGND.t1629 VGND.t2314 724.904
R15631 VGND.t2663 VGND.t2665 724.904
R15632 VGND.t2665 VGND.t2667 724.904
R15633 VGND.t2012 VGND.t560 724.904
R15634 VGND.t3031 VGND.t3035 724.904
R15635 VGND.t3242 VGND.t3246 724.904
R15636 VGND VGND.t1690 724.904
R15637 VGND.t2698 VGND 724.904
R15638 VGND.t2020 VGND.t2016 724.904
R15639 VGND.t1858 VGND.t2464 724.904
R15640 VGND.t2154 VGND.t2158 724.904
R15641 VGND.t2158 VGND.t2152 724.904
R15642 VGND.t2152 VGND.t2156 724.904
R15643 VGND.t1312 VGND.t3004 724.904
R15644 VGND.t718 VGND.t716 724.904
R15645 VGND.t2445 VGND.t2441 724.904
R15646 VGND.t56 VGND.t2078 716.476
R15647 VGND.t130 VGND.t175 716.476
R15648 VGND.t2382 VGND 716.476
R15649 VGND.t2107 VGND.t2117 716.476
R15650 VGND.t2945 VGND.t2012 716.476
R15651 VGND VGND.t1781 716.025
R15652 VGND VGND.t1846 716.025
R15653 VGND.t3123 VGND.t2138 708.047
R15654 VGND.t533 VGND.t279 708.047
R15655 VGND.t2074 VGND.t58 708.047
R15656 VGND.t2050 VGND.t2141 708.047
R15657 VGND.t3131 VGND.t3133 708.047
R15658 VGND.t1948 VGND.t1745 708.047
R15659 VGND.t1864 VGND.t1868 708.047
R15660 VGND.t1929 VGND.t1927 708.047
R15661 VGND.t173 VGND.t128 708.047
R15662 VGND.t271 VGND.t1735 708.047
R15663 VGND.t1959 VGND.t1956 708.047
R15664 VGND.t1956 VGND.t2544 708.047
R15665 VGND.t2544 VGND.t2540 708.047
R15666 VGND.t2540 VGND.t2536 708.047
R15667 VGND.t2542 VGND.t2546 708.047
R15668 VGND.t2546 VGND.t2538 708.047
R15669 VGND.t121 VGND.t119 708.047
R15670 VGND.t506 VGND.t504 708.047
R15671 VGND.t504 VGND.t510 708.047
R15672 VGND.t510 VGND.t502 708.047
R15673 VGND.t502 VGND.t508 708.047
R15674 VGND.t508 VGND.t500 708.047
R15675 VGND.t500 VGND.t3055 708.047
R15676 VGND.t1751 VGND.t2350 708.047
R15677 VGND.t1727 VGND.t2137 708.047
R15678 VGND.t2234 VGND.t275 708.047
R15679 VGND.t1874 VGND.t1902 708.047
R15680 VGND.t422 VGND.t424 708.047
R15681 VGND.t2640 VGND.t285 708.047
R15682 VGND.t111 VGND.t113 708.047
R15683 VGND.t113 VGND.t1731 708.047
R15684 VGND.t1731 VGND.t1733 708.047
R15685 VGND.t1710 VGND.t2203 708.047
R15686 VGND.t704 VGND.t698 708.047
R15687 VGND.t698 VGND.t3215 708.047
R15688 VGND.t3209 VGND.t3207 708.047
R15689 VGND.t3207 VGND.t3213 708.047
R15690 VGND.t3213 VGND.t3217 708.047
R15691 VGND.t1918 VGND.t1755 708.047
R15692 VGND.t1664 VGND.t1662 708.047
R15693 VGND.t30 VGND.t29 708.047
R15694 VGND.t1695 VGND.t31 708.047
R15695 VGND.t2580 VGND.t737 708.047
R15696 VGND.t2293 VGND.t2261 708.047
R15697 VGND.t3091 VGND.t3093 708.047
R15698 VGND.t2325 VGND.t1655 708.047
R15699 VGND.t398 VGND.t450 708.047
R15700 VGND.t2897 VGND.t2899 708.047
R15701 VGND.t2322 VGND.t1656 708.047
R15702 VGND.t2198 VGND.t1759 708.047
R15703 VGND.t574 VGND.t576 708.047
R15704 VGND.t2616 VGND.t2745 708.047
R15705 VGND.t1838 VGND.t1836 708.047
R15706 VGND.t786 VGND.t2383 708.047
R15707 VGND.t2598 VGND.t2602 708.047
R15708 VGND.t1884 VGND.t2182 708.047
R15709 VGND.t562 VGND.t564 708.047
R15710 VGND.t2295 VGND.t2286 708.047
R15711 VGND.t2575 VGND.t1597 708.047
R15712 VGND.t1597 VGND.t1598 708.047
R15713 VGND.t455 VGND.t633 708.047
R15714 VGND.t2385 VGND.t2189 708.047
R15715 VGND.t2679 VGND.t804 708.047
R15716 VGND.t2378 VGND.t2187 708.047
R15717 VGND.t2185 VGND.t2070 708.047
R15718 VGND.t1636 VGND.t3101 708.047
R15719 VGND.t762 VGND.t1896 708.047
R15720 VGND.t1763 VGND.t297 708.047
R15721 VGND.t385 VGND.t389 708.047
R15722 VGND.t2353 VGND.t385 708.047
R15723 VGND.t3235 VGND.t2353 708.047
R15724 VGND.t1795 VGND.t3141 708.047
R15725 VGND.t2613 VGND.t2611 708.047
R15726 VGND.t1894 VGND.t1913 708.047
R15727 VGND.t2146 VGND.t2566 708.047
R15728 VGND.t183 VGND.t2975 708.047
R15729 VGND.t2986 VGND.t1970 708.047
R15730 VGND.t1925 VGND.t51 708.047
R15731 VGND.t2596 VGND.t2588 708.047
R15732 VGND.t724 VGND.t730 708.047
R15733 VGND.t522 VGND.t914 708.047
R15734 VGND.t2946 VGND.t2941 708.047
R15735 VGND.t2889 VGND.t1892 708.047
R15736 VGND.t1647 VGND.t1649 708.047
R15737 VGND.t1890 VGND.t1935 708.047
R15738 VGND.t2066 VGND.t1909 708.047
R15739 VGND.t3159 VGND.t3117 708.047
R15740 VGND.t144 VGND.t3196 708.047
R15741 VGND.t1814 VGND.t83 708.047
R15742 VGND.t2447 VGND.t2449 708.047
R15743 VGND.t78 VGND.t76 708.047
R15744 VGND.t2774 VGND.t2778 708.047
R15745 VGND.t205 VGND.t1808 708.047
R15746 VGND.t2058 VGND.t2453 708.047
R15747 VGND.t140 VGND.t2339 708.047
R15748 VGND.t267 VGND.t2079 708.047
R15749 VGND.t3066 VGND.t2135 708.047
R15750 VGND.t2620 VGND.t2618 708.047
R15751 VGND.t1644 VGND.t1810 708.047
R15752 VGND.t2395 VGND.t2397 708.047
R15753 VGND.t3171 VGND.t3169 708.047
R15754 VGND.t734 VGND.t732 708.047
R15755 VGND.t2030 VGND.t2028 708.047
R15756 VGND.t2272 VGND.t2274 708.047
R15757 VGND.t3165 VGND.t3167 708.047
R15758 VGND.t135 VGND.t2008 708.047
R15759 VGND.t104 VGND.t102 708.047
R15760 VGND.t569 VGND.t2853 708.047
R15761 VGND.t528 VGND.t526 708.047
R15762 VGND.t2366 VGND.t320 699.617
R15763 VGND.t661 VGND 699.617
R15764 VGND.t3041 VGND.t558 699.617
R15765 VGND VGND.t213 699.617
R15766 VGND.t1915 VGND 699.617
R15767 VGND.t2728 VGND.t1793 699.617
R15768 VGND.t3047 VGND.t150 699.617
R15769 VGND.t2811 VGND.t2973 699.617
R15770 VGND.t2652 VGND.t2087 699.617
R15771 VGND VGND.t1959 691.188
R15772 VGND VGND.t704 691.188
R15773 VGND.t1397 VGND.t2164 691.188
R15774 VGND.t2097 VGND.t2895 691.188
R15775 VGND.t1916 VGND 691.188
R15776 VGND.t387 VGND 691.188
R15777 VGND.t3015 VGND.t1635 691.188
R15778 VGND.t2533 VGND.t2195 691.188
R15779 VGND.t2970 VGND.t961 691.188
R15780 VGND.t1812 VGND.t2443 691.188
R15781 VGND.t90 VGND 683.231
R15782 VGND.t2427 VGND.t244 682.76
R15783 VGND.t702 VGND.t1958 682.76
R15784 VGND.t2286 VGND.t1243 682.76
R15785 VGND.t2750 VGND.t667 682.76
R15786 VGND.t1637 VGND.t3151 682.76
R15787 VGND.t374 VGND 682.76
R15788 VGND.t2134 VGND.t2727 682.76
R15789 VGND.t1702 VGND.t2969 682.76
R15790 VGND VGND.t2357 677.764
R15791 VGND VGND.t39 677.764
R15792 VGND.t770 VGND.t2979 674.331
R15793 VGND.t3175 VGND.t758 674.331
R15794 VGND.t540 VGND 674.331
R15795 VGND.t3108 VGND 672.298
R15796 VGND.t687 VGND 672.298
R15797 VGND VGND.t3223 672.298
R15798 VGND.n1483 VGND.n1482 667.915
R15799 VGND.t1834 VGND.t2642 665.9
R15800 VGND.t2819 VGND.t644 665.9
R15801 VGND.t312 VGND 665.9
R15802 VGND.t3229 VGND.t24 665.9
R15803 VGND.t439 VGND.t3233 665.9
R15804 VGND.t2761 VGND.t2634 665.9
R15805 VGND.t2333 VGND.t2429 657.471
R15806 VGND.t2872 VGND.t420 657.471
R15807 VGND.t307 VGND.t463 657.471
R15808 VGND.t536 VGND.t635 657.471
R15809 VGND.t2564 VGND.t2736 657.471
R15810 VGND.t2740 VGND.t2961 657.471
R15811 VGND.t1476 VGND.t657 657.471
R15812 VGND.t1765 VGND.t74 657.471
R15813 VGND.t1908 VGND.t3033 657.471
R15814 VGND.t2681 VGND.t2244 657.471
R15815 VGND.t415 VGND.t1968 649.043
R15816 VGND.t1816 VGND.t2497 649.043
R15817 VGND VGND.n4660 649.043
R15818 VGND.t450 VGND.t587 649.043
R15819 VGND.t60 VGND 649.043
R15820 VGND.t2215 VGND.t2119 649.043
R15821 VGND.t310 VGND.t318 649.043
R15822 VGND.t2174 VGND.t3149 649.043
R15823 VGND.n8338 VGND 649.043
R15824 VGND.t3163 VGND.t2316 649.043
R15825 VGND VGND.n158 649.043
R15826 VGND.t796 VGND 649.043
R15827 VGND.t1607 VGND.t1878 640.614
R15828 VGND.t1603 VGND.t131 640.614
R15829 VGND.t1606 VGND.t2839 640.614
R15830 VGND.t1716 VGND.t422 640.614
R15831 VGND.t3005 VGND.t307 640.614
R15832 VGND.t139 VGND.t1985 640.614
R15833 VGND.t1662 VGND.t2142 640.614
R15834 VGND.t1658 VGND.t2148 640.614
R15835 VGND.t16 VGND.t2212 640.614
R15836 VGND.t12 VGND.t2227 640.614
R15837 VGND VGND.t1424 640.614
R15838 VGND.t1656 VGND.t303 640.614
R15839 VGND.t556 VGND.t2521 640.614
R15840 VGND.t844 VGND.t2048 640.614
R15841 VGND.t1451 VGND.t2170 640.614
R15842 VGND.t1575 VGND.t724 640.614
R15843 VGND.t1688 VGND.t1833 640.614
R15844 VGND.t2891 VGND 640.614
R15845 VGND.t1651 VGND.t787 640.614
R15846 VGND.t791 VGND.t3115 640.614
R15847 VGND.t2638 VGND.t792 640.614
R15848 VGND.t2131 VGND.t796 640.614
R15849 VGND.t1704 VGND.t1952 640.614
R15850 VGND.t797 VGND.t604 640.614
R15851 VGND VGND.t908 632.184
R15852 VGND.n6629 VGND 632.184
R15853 VGND.n6630 VGND 632.184
R15854 VGND.n5338 VGND 632.184
R15855 VGND VGND.t1270 632.184
R15856 VGND.n6337 VGND 632.184
R15857 VGND VGND.t1607 632.184
R15858 VGND VGND.n1590 632.184
R15859 VGND.t1056 VGND 632.184
R15860 VGND.t2567 VGND.t736 632.184
R15861 VGND.n6979 VGND 632.184
R15862 VGND VGND.t1039 632.184
R15863 VGND VGND.n5102 632.184
R15864 VGND VGND.n5101 632.184
R15865 VGND VGND.n5098 632.184
R15866 VGND VGND.t848 632.184
R15867 VGND VGND.n806 632.184
R15868 VGND VGND.n7311 632.184
R15869 VGND VGND.t1394 632.184
R15870 VGND.n7685 VGND 632.184
R15871 VGND.n8254 VGND 632.184
R15872 VGND.n8335 VGND 632.184
R15873 VGND VGND.t1140 632.184
R15874 VGND VGND.t2659 632.184
R15875 VGND.t1714 VGND 632.184
R15876 VGND VGND.t931 632.184
R15877 VGND.t1217 VGND 632.184
R15878 VGND.n181 VGND 632.184
R15879 VGND VGND.t1237 632.184
R15880 VGND.n8908 VGND 632.184
R15881 VGND.n8909 VGND 632.184
R15882 VGND.n3032 VGND 632.184
R15883 VGND.n3201 VGND 632.184
R15884 VGND VGND.t1024 632.184
R15885 VGND VGND.n2107 632.184
R15886 VGND.n2662 VGND 632.184
R15887 VGND.t794 VGND.t3045 632.184
R15888 VGND VGND.n3208 632.184
R15889 VGND VGND.n3207 632.184
R15890 VGND VGND.t1030 632.184
R15891 VGND.n9182 VGND 632.184
R15892 VGND VGND.n9181 632.184
R15893 VGND VGND.n9178 632.184
R15894 VGND.t248 VGND.t2417 623.755
R15895 VGND.t2696 VGND.t2411 623.755
R15896 VGND.t694 VGND.t1412 623.755
R15897 VGND VGND.n5100 623.755
R15898 VGND VGND.n5099 623.755
R15899 VGND.t564 VGND.t2105 623.755
R15900 VGND VGND.t212 623.755
R15901 VGND.t884 VGND.t1799 623.755
R15902 VGND VGND.t3181 623.755
R15903 VGND VGND.n9179 623.755
R15904 VGND.t2773 VGND.t2631 615.327
R15905 VGND.t192 VGND.t2879 615.327
R15906 VGND.t2164 VGND 615.327
R15907 VGND.t2246 VGND.t210 615.327
R15908 VGND.t2257 VGND.t1876 615.327
R15909 VGND.t2099 VGND 615.327
R15910 VGND.t1612 VGND.t2523 615.327
R15911 VGND.t1951 VGND.t1125 615.327
R15912 VGND.t520 VGND 615.327
R15913 VGND.t72 VGND.t3083 615.327
R15914 VGND.t787 VGND.t1676 615.327
R15915 VGND VGND.t2133 615.327
R15916 VGND VGND.t1976 615.327
R15917 VGND.t2083 VGND 615.327
R15918 VGND.n5099 VGND.n1335 613.249
R15919 VGND.n4660 VGND.n4168 613.249
R15920 VGND.n4658 VGND.n4657 613.249
R15921 VGND.n8784 VGND.n158 613.249
R15922 VGND.n8255 VGND.n8254 613.249
R15923 VGND.n7312 VGND.n887 613.249
R15924 VGND.n6857 VGND.n1590 613.249
R15925 VGND.n6455 VGND.n6338 613.249
R15926 VGND.n5815 VGND.n5814 613.249
R15927 VGND.n5812 VGND.n5125 613.249
R15928 VGND.n5811 VGND.n5810 613.249
R15929 VGND.n5813 VGND.n5124 613.249
R15930 VGND.n5940 VGND.n5107 613.249
R15931 VGND.n6337 VGND.n6336 613.249
R15932 VGND.n6384 VGND.n6354 613.249
R15933 VGND.n6976 VGND.n6975 613.249
R15934 VGND.n4659 VGND.n4169 613.249
R15935 VGND.n5102 VGND.n3985 613.249
R15936 VGND.n5100 VGND.n5087 613.249
R15937 VGND.n7811 VGND.n7810 613.249
R15938 VGND.n7942 VGND.n7941 613.249
R15939 VGND.n8339 VGND.n8338 613.249
R15940 VGND.n3980 VGND.n3979 613.249
R15941 VGND.n306 VGND.n305 613.249
R15942 VGND.n8979 VGND.n78 613.249
R15943 VGND.n3201 VGND.n3200 613.249
R15944 VGND.n3264 VGND.n3209 613.249
R15945 VGND.n3207 VGND.n2664 613.249
R15946 VGND.n9180 VGND.n19 613.249
R15947 VGND.n5101 VGND.n3986 611.862
R15948 VGND.n9178 VGND.n9177 611.862
R15949 VGND.n2662 VGND.n2644 611.225
R15950 VGND.n8910 VGND.n8909 611.225
R15951 VGND.n8908 VGND.n8907 611.225
R15952 VGND.n5337 VGND.n5336 610.679
R15953 VGND.n9183 VGND.n9182 609.497
R15954 VGND.n5402 VGND.n5338 609.497
R15955 VGND.n6631 VGND.n6630 609.497
R15956 VGND.n3208 VGND.n2663 609.497
R15957 VGND.n3069 VGND.n3032 609.497
R15958 VGND.n8623 VGND.n222 609.497
R15959 VGND.n8040 VGND.n7943 609.497
R15960 VGND.n7813 VGND.n7812 609.497
R15961 VGND.n7687 VGND.n7685 609.497
R15962 VGND.n7315 VGND.n7314 609.497
R15963 VGND.n6629 VGND.n6628 609.497
R15964 VGND.n6696 VGND.n1624 609.497
R15965 VGND.n4662 VGND.n4661 609.497
R15966 VGND.n6980 VGND.n6979 609.497
R15967 VGND.n5098 VGND.n5097 609.497
R15968 VGND.n7393 VGND.n806 609.497
R15969 VGND.n7311 VGND.n7310 609.497
R15970 VGND.n7313 VGND.n886 609.497
R15971 VGND.n7684 VGND.n7683 609.497
R15972 VGND.n8253 VGND.n8252 609.497
R15973 VGND.n8335 VGND.n8334 609.497
R15974 VGND.n8735 VGND.n181 609.497
R15975 VGND.n3427 VGND.n2107 609.497
R15976 VGND.t1968 VGND.t250 606.898
R15977 VGND.t228 VGND.t1906 606.898
R15978 VGND.t2470 VGND.t2771 606.898
R15979 VGND.t2780 VGND.n6337 606.898
R15980 VGND.t3154 VGND.t2488 606.898
R15981 VGND.t1958 VGND.t3061 606.898
R15982 VGND.t2482 VGND.t187 606.898
R15983 VGND.t262 VGND.t258 606.898
R15984 VGND.t2271 VGND.t246 606.898
R15985 VGND.t599 VGND.t1882 606.898
R15986 VGND.t2472 VGND.t1991 606.898
R15987 VGND.t232 VGND.t417 606.898
R15988 VGND.t29 VGND.t2959 606.898
R15989 VGND.t757 VGND.t2963 606.898
R15990 VGND.t2474 VGND.t98 606.898
R15991 VGND.t1923 VGND.t1164 606.898
R15992 VGND.t1818 VGND.t230 606.898
R15993 VGND.t2903 VGND.t673 606.898
R15994 VGND.t1684 VGND.t1915 606.898
R15995 VGND.t2282 VGND.t2795 606.898
R15996 VGND.t623 VGND.t449 606.898
R15997 VGND.t531 VGND.t2702 606.898
R15998 VGND.t2552 VGND.t802 606.898
R15999 VGND.t2364 VGND.t1950 606.898
R16000 VGND.t1672 VGND.t2363 606.898
R16001 VGND.t3204 VGND.t2716 606.898
R16002 VGND.t728 VGND.t2590 606.898
R16003 VGND.t726 VGND.t2594 606.898
R16004 VGND.t730 VGND.t2586 606.898
R16005 VGND.t362 VGND.t2391 606.898
R16006 VGND.t1833 VGND.t2891 606.898
R16007 VGND.t462 VGND.t1674 606.898
R16008 VGND.t1820 VGND.t152 606.898
R16009 VGND.t154 VGND.t1670 606.898
R16010 VGND.t2656 VGND.t1680 606.898
R16011 VGND.t393 VGND.t2783 606.898
R16012 VGND.t1690 VGND.t2934 606.898
R16013 VGND.t2712 VGND.t608 606.898
R16014 VGND.t1943 VGND.t1161 606.898
R16015 VGND.t101 VGND.t2698 606.898
R16016 VGND.t2787 VGND.t637 606.898
R16017 VGND.t2415 VGND.t746 598.467
R16018 VGND.t2331 VGND.t2409 598.467
R16019 VGND.t1208 VGND.t240 598.467
R16020 VGND.t2956 VGND.t700 598.467
R16021 VGND.t2248 VGND.t1870 598.467
R16022 VGND.t784 VGND 598.467
R16023 VGND.t2553 VGND.t2379 598.467
R16024 VGND.t2948 VGND.t2172 598.467
R16025 VGND.t689 VGND.t1819 598.467
R16026 VGND.t3029 VGND.t261 598.467
R16027 VGND.t109 VGND.t2531 598.467
R16028 VGND.n9180 VGND.t2797 598.467
R16029 VGND.t2042 VGND 598.467
R16030 VGND VGND.t2445 598.467
R16031 VGND VGND.t1246 595.777
R16032 VGND.t1418 VGND 595.777
R16033 VGND.t1442 VGND 595.777
R16034 VGND.t1566 VGND 595.777
R16035 VGND.t3078 VGND.t198 590.038
R16036 VGND.n6354 VGND.t2369 590.038
R16037 VGND.t2536 VGND.t967 590.038
R16038 VGND.t2352 VGND.n6976 590.038
R16039 VGND.t2678 VGND.t1099 590.038
R16040 VGND.t1560 VGND.t2382 590.038
R16041 VGND.t3237 VGND.t671 590.038
R16042 VGND.t2187 VGND 590.038
R16043 VGND.t2584 VGND.t808 590.038
R16044 VGND VGND.t2146 590.038
R16045 VGND.t2975 VGND 590.038
R16046 VGND.t53 VGND 590.038
R16047 VGND.t795 VGND.t368 590.038
R16048 VGND VGND.t1934 590.038
R16049 VGND.t283 VGND.t2413 581.61
R16050 VGND.t2925 VGND.t2863 581.61
R16051 VGND VGND.t180 581.61
R16052 VGND.t584 VGND 581.61
R16053 VGND.t400 VGND.t2815 581.61
R16054 VGND.t305 VGND.t1719 581.61
R16055 VGND.t2200 VGND 581.61
R16056 VGND.t1202 VGND.t2385 581.61
R16057 VGND.t1617 VGND 581.61
R16058 VGND.t391 VGND.t2377 581.61
R16059 VGND.t1631 VGND 581.61
R16060 VGND VGND.t3157 581.61
R16061 VGND.t270 VGND 581.61
R16062 VGND.t3076 VGND 581.61
R16063 VGND.t3004 VGND 581.61
R16064 VGND.t2971 VGND.t973 581.61
R16065 VGND.t401 VGND.t2427 573.181
R16066 VGND.t177 VGND.t1727 573.181
R16067 VGND.t10 VGND 573.181
R16068 VGND.t2297 VGND 573.181
R16069 VGND.t3200 VGND 573.181
R16070 VGND.t742 VGND.t740 573.181
R16071 VGND VGND.t3235 573.181
R16072 VGND.t3023 VGND.t2508 573.181
R16073 VGND.t2223 VGND.t3228 573.181
R16074 VGND.t3064 VGND.t1741 573.181
R16075 VGND.t1646 VGND.t1282 573.181
R16076 VGND.t2833 VGND.t2857 573.181
R16077 VGND.t2028 VGND 573.181
R16078 VGND.t200 VGND 564.751
R16079 VGND.t119 VGND 564.751
R16080 VGND VGND.t3059 564.751
R16081 VGND.t2137 VGND 564.751
R16082 VGND VGND.t3069 564.751
R16083 VGND.t2745 VGND 564.751
R16084 VGND.t1620 VGND.t2115 564.751
R16085 VGND.t309 VGND 564.751
R16086 VGND VGND.t2381 564.751
R16087 VGND.t1682 VGND.t45 564.751
R16088 VGND.t3173 VGND 564.751
R16089 VGND.t1802 VGND.t3068 564.751
R16090 VGND.t1990 VGND 564.751
R16091 VGND VGND.t2774 564.751
R16092 VGND.t204 VGND.t161 564.751
R16093 VGND VGND.t443 564.751
R16094 VGND.t102 VGND.t2221 564.751
R16095 VGND.t1170 VGND.t636 556.322
R16096 VGND.t80 VGND 556.322
R16097 VGND VGND.t2995 556.322
R16098 VGND.t1445 VGND.t1984 556.322
R16099 VGND.t2643 VGND.t426 556.322
R16100 VGND.t2885 VGND 556.322
R16101 VGND.t2883 VGND 556.322
R16102 VGND.t1917 VGND.t2827 556.322
R16103 VGND.t2338 VGND.t1513 556.322
R16104 VGND.t1980 VGND 556.322
R16105 VGND.t645 VGND 556.322
R16106 VGND.t2355 VGND.t2184 556.322
R16107 VGND.t570 VGND.t1021 556.322
R16108 VGND.t1642 VGND.t1090 556.322
R16109 VGND.t6 VGND 556.322
R16110 VGND.t260 VGND.t1522 556.322
R16111 VGND VGND.t2447 556.322
R16112 VGND.t2343 VGND 556.322
R16113 VGND.t2973 VGND.t2708 556.322
R16114 VGND.t2259 VGND 556.322
R16115 VGND.t1701 VGND.t146 556.322
R16116 VGND.t2 VGND 556.322
R16117 VGND.t732 VGND 556.322
R16118 VGND.t2264 VGND 556.322
R16119 VGND.t287 VGND 547.894
R16120 VGND.t1745 VGND 547.894
R16121 VGND VGND.t2076 547.894
R16122 VGND.t2330 VGND.t2431 547.894
R16123 VGND.t3057 VGND 547.894
R16124 VGND.t2997 VGND 547.894
R16125 VGND VGND.t1751 547.894
R16126 VGND VGND.t3106 547.894
R16127 VGND VGND.t281 547.894
R16128 VGND.t285 VGND 547.894
R16129 VGND.t2024 VGND 547.894
R16130 VGND.t2205 VGND 547.894
R16131 VGND.t1755 VGND 547.894
R16132 VGND.t1985 VGND 547.894
R16133 VGND.t2288 VGND 547.894
R16134 VGND.t293 VGND 547.894
R16135 VGND.t1717 VGND 547.894
R16136 VGND VGND.t2321 547.894
R16137 VGND.t1721 VGND 547.894
R16138 VGND.t1759 VGND 547.894
R16139 VGND.t2676 VGND 547.894
R16140 VGND VGND.t2813 547.894
R16141 VGND.n7313 VGND.t2295 547.894
R16142 VGND.t2785 VGND.t2578 547.894
R16143 VGND.t1753 VGND 547.894
R16144 VGND.t1747 VGND 547.894
R16145 VGND.t99 VGND 547.894
R16146 VGND VGND.t1763 547.894
R16147 VGND.t2494 VGND 547.894
R16148 VGND.t1761 VGND 547.894
R16149 VGND VGND.t1749 547.894
R16150 VGND.t2611 VGND 547.894
R16151 VGND.t2738 VGND 547.894
R16152 VGND VGND.t1925 547.894
R16153 VGND.t3239 VGND 547.894
R16154 VGND.t350 VGND.t1766 547.894
R16155 VGND.t1779 VGND 547.894
R16156 VGND VGND.t1890 547.894
R16157 VGND VGND.t2066 547.894
R16158 VGND.t2079 VGND 547.894
R16159 VGND VGND.t2062 547.894
R16160 VGND.t1806 VGND 547.894
R16161 VGND.t2466 VGND 547.894
R16162 VGND.t604 VGND 547.894
R16163 VGND.t2397 VGND 547.894
R16164 VGND.t202 VGND 547.894
R16165 VGND.t2776 VGND 547.894
R16166 VGND.t2064 VGND 547.894
R16167 VGND.t2038 VGND.t602 547.894
R16168 VGND VGND.t1473 539.465
R16169 VGND.t218 VGND.t776 539.465
R16170 VGND.t2203 VGND 539.465
R16171 VGND.t994 VGND 539.465
R16172 VGND.t31 VGND 539.465
R16173 VGND.t2870 VGND.t1872 539.465
R16174 VGND.t1886 VGND 539.465
R16175 VGND.t2578 VGND 539.465
R16176 VGND.n7312 VGND.t2740 539.465
R16177 VGND VGND.t665 539.465
R16178 VGND.t2505 VGND.t846 539.465
R16179 VGND.t3185 VGND.t2308 539.465
R16180 VGND.t512 VGND.n7942 539.465
R16181 VGND VGND.t940 539.465
R16182 VGND.t2700 VGND.t3064 539.465
R16183 VGND VGND.t1470 539.465
R16184 VGND.t2857 VGND.t2714 539.465
R16185 VGND.t3169 VGND 539.465
R16186 VGND.t1327 VGND 539.465
R16187 VGND.t2008 VGND 539.465
R16188 VGND.t430 VGND 531.034
R16189 VGND.t238 VGND.t200 531.034
R16190 VGND.t279 VGND 531.034
R16191 VGND.t863 VGND 531.034
R16192 VGND.t1557 VGND 531.034
R16193 VGND VGND.t1627 531.034
R16194 VGND VGND.t1391 531.034
R16195 VGND.t1205 VGND 531.034
R16196 VGND.t1361 VGND 531.034
R16197 VGND.t1743 VGND 531.034
R16198 VGND.t467 VGND 531.034
R16199 VGND.t825 VGND.t2909 531.034
R16200 VGND VGND.t1421 531.034
R16201 VGND.t1231 VGND 531.034
R16202 VGND.t2504 VGND 531.034
R16203 VGND.t2988 VGND.t1775 531.034
R16204 VGND.t585 VGND 531.034
R16205 VGND VGND.t1814 531.034
R16206 VGND VGND.t1388 531.034
R16207 VGND VGND.t1504 531.034
R16208 VGND VGND.t1797 531.034
R16209 VGND.t1840 VGND 531.034
R16210 VGND VGND.t2637 531.034
R16211 VGND VGND.t1554 531.034
R16212 VGND VGND.t2207 531.034
R16213 VGND.t1285 VGND 531.034
R16214 VGND.t606 VGND 531.034
R16215 VGND.t1432 VGND 531.034
R16216 VGND.t1158 VGND 531.034
R16217 VGND.t2040 VGND.t3072 531.034
R16218 VGND.t1787 VGND.t376 530.187
R16219 VGND.t1844 VGND.t2724 530.187
R16220 VGND.t2478 VGND.t2861 522.606
R16221 VGND.t381 VGND 522.606
R16222 VGND.t2915 VGND 522.606
R16223 VGND.t2252 VGND.t3225 522.606
R16224 VGND.t2720 VGND 522.606
R16225 VGND.t33 VGND 522.606
R16226 VGND.t2817 VGND 522.606
R16227 VGND.t308 VGND.t2823 522.606
R16228 VGND.t2500 VGND.t835 522.606
R16229 VGND.t802 VGND 522.606
R16230 VGND.t693 VGND.t2268 522.606
R16231 VGND.t94 VGND 522.606
R16232 VGND.t722 VGND.t3143 522.606
R16233 VGND.t2752 VGND.t685 519.255
R16234 VGND.t714 VGND.t1697 519.255
R16235 VGND.t2952 VGND.t418 519.255
R16236 VGND.t2359 VGND.t3112 519.255
R16237 VGND.t37 VGND.t2010 519.255
R16238 VGND.t1725 VGND.t3027 519.255
R16239 VGND VGND.t413 514.177
R16240 VGND.t214 VGND 514.177
R16241 VGND VGND.t595 514.177
R16242 VGND VGND.t2280 514.177
R16243 VGND.t600 VGND 514.177
R16244 VGND.t3128 VGND 514.177
R16245 VGND.t2759 VGND 514.177
R16246 VGND.t2310 VGND 514.177
R16247 VGND.t3179 VGND 514.177
R16248 VGND.t774 VGND 514.177
R16249 VGND.t3202 VGND 514.177
R16250 VGND.t2570 VGND 514.177
R16251 VGND VGND.t1105 514.177
R16252 VGND.t20 VGND 514.177
R16253 VGND.t782 VGND 514.177
R16254 VGND VGND.t96 514.177
R16255 VGND VGND.t1825 514.177
R16256 VGND.t1827 VGND 514.177
R16257 VGND.t2457 VGND 514.177
R16258 VGND.t1856 VGND 514.177
R16259 VGND VGND.t2439 514.177
R16260 VGND.t1608 VGND.t1137 505.748
R16261 VGND VGND.t811 505.748
R16262 VGND.t2254 VGND.t2423 505.748
R16263 VGND.t516 VGND 505.748
R16264 VGND.t246 VGND.t262 505.748
R16265 VGND.t3069 VGND.t581 505.748
R16266 VGND.t2139 VGND.t277 505.748
R16267 VGND.t14 VGND 505.748
R16268 VGND.t2957 VGND 505.748
R16269 VGND.t2103 VGND.t2144 505.748
R16270 VGND VGND.t2991 505.748
R16271 VGND.t1640 VGND 505.748
R16272 VGND.t2300 VGND 505.748
R16273 VGND.t1774 VGND.t2758 505.748
R16274 VGND.t2689 VGND 497.318
R16275 VGND.t778 VGND 497.318
R16276 VGND.t2657 VGND 497.318
R16277 VGND.t2977 VGND.t1880 497.318
R16278 VGND.t1876 VGND.t256 497.318
R16279 VGND.t295 VGND.t2722 497.318
R16280 VGND.t1944 VGND 497.318
R16281 VGND.t492 VGND 497.318
R16282 VGND VGND.t62 497.318
R16283 VGND.t2867 VGND.t3119 497.318
R16284 VGND VGND.t2756 497.318
R16285 VGND.n7811 VGND.t1912 497.318
R16286 VGND.t2389 VGND 497.318
R16287 VGND.t3155 VGND 497.318
R16288 VGND VGND.t154 497.318
R16289 VGND.t765 VGND 497.318
R16290 VGND.t3248 VGND 497.318
R16291 VGND.t2018 VGND 497.318
R16292 VGND.t445 VGND 497.318
R16293 VGND.t1866 VGND 497.318
R16294 VGND.t2417 VGND.t2370 488.889
R16295 VGND.t1412 VGND.t2482 488.889
R16296 VGND.t473 VGND 488.889
R16297 VGND.t649 VGND 488.889
R16298 VGND.t2109 VGND.t2561 488.889
R16299 VGND VGND.t760 488.889
R16300 VGND VGND.t350 488.889
R16301 VGND VGND.t3017 488.889
R16302 VGND.t1680 VGND.t884 488.889
R16303 VGND.t2550 VGND.t3108 480.995
R16304 VGND.t3223 VGND.t2911 480.995
R16305 VGND.t2528 VGND 480.461
R16306 VGND VGND.t475 480.461
R16307 VGND.t3217 VGND 480.461
R16308 VGND VGND.t764 480.461
R16309 VGND.t2558 VGND 480.461
R16310 VGND.t2150 VGND 480.461
R16311 VGND.t2323 VGND 480.461
R16312 VGND.t1708 VGND 480.461
R16313 VGND.t2507 VGND.t2127 480.461
R16314 VGND VGND.t2125 480.461
R16315 VGND.t669 VGND.t2993 480.461
R16316 VGND.t2830 VGND 480.461
R16317 VGND.t2592 VGND.t484 480.461
R16318 VGND.t148 VGND 480.461
R16319 VGND.n3209 VGND.t2627 480.461
R16320 VGND.t591 VGND 480.461
R16321 VGND.t1589 VGND 480.461
R16322 VGND.t3001 VGND 480.461
R16323 VGND.t250 VGND 472.031
R16324 VGND.t3059 VGND.t516 472.031
R16325 VGND.t1609 VGND 472.031
R16326 VGND.t2372 VGND.t64 472.031
R16327 VGND.t2805 VGND 472.031
R16328 VGND.t3153 VGND 472.031
R16329 VGND.t1972 VGND.t184 472.031
R16330 VGND.t3145 VGND 472.031
R16331 VGND.t1952 VGND.t621 472.031
R16332 VGND.t716 VGND.t2693 472.031
R16333 VGND.t1781 VGND.t1783 470.062
R16334 VGND.t1783 VGND.t1785 470.062
R16335 VGND.t1785 VGND.t1787 470.062
R16336 VGND.t1846 VGND.t1848 470.062
R16337 VGND.t1848 VGND.t1842 470.062
R16338 VGND.t1842 VGND.t1844 470.062
R16339 VGND VGND.t3078 463.603
R16340 VGND.t2907 VGND 463.603
R16341 VGND.t747 VGND.t2403 463.603
R16342 VGND VGND.t2744 463.603
R16343 VGND.t2600 VGND.t18 463.603
R16344 VGND.t3019 VGND 463.603
R16345 VGND.t326 VGND.t2799 463.603
R16346 VGND.t793 VGND.t1633 463.603
R16347 VGND.t2318 VGND 463.603
R16348 VGND.t498 VGND.n3980 463.603
R16349 VGND.t769 VGND 463.603
R16350 VGND.t2531 VGND 463.603
R16351 VGND VGND.t2285 463.603
R16352 VGND VGND.t2217 463.603
R16353 VGND.t619 VGND.t1931 463.603
R16354 VGND.t685 VGND.t687 459.13
R16355 VGND.t1697 VGND.t1699 459.13
R16356 VGND.t88 VGND.t90 459.13
R16357 VGND.t2950 VGND.t2952 459.13
R16358 VGND.t2357 VGND.t2359 459.13
R16359 VGND.t39 VGND.t37 459.13
R16360 VGND.t3027 VGND.t3025 459.13
R16361 VGND VGND.t316 455.173
R16362 VGND VGND.t2925 455.173
R16363 VGND.t3215 VGND.t1338 455.173
R16364 VGND.t417 VGND.t1253 455.173
R16365 VGND.t1875 VGND.t66 455.173
R16366 VGND.t2961 VGND.t2793 455.173
R16367 VGND.t1199 VGND.t531 455.173
R16368 VGND.t366 VGND.t2644 455.173
R16369 VGND.t2791 VGND 455.173
R16370 VGND VGND.t1686 455.173
R16371 VGND VGND.t2807 455.173
R16372 VGND VGND.t2465 455.173
R16373 VGND.t1965 VGND.t2176 455.173
R16374 VGND.t2244 VGND.t2803 455.173
R16375 VGND.t2044 VGND.t1595 455.173
R16376 VGND.t127 VGND 446.743
R16377 VGND VGND.t252 446.743
R16378 VGND.t1921 VGND.t378 446.743
R16379 VGND.t739 VGND 446.743
R16380 VGND VGND.t234 446.743
R16381 VGND VGND.t583 446.743
R16382 VGND VGND.t2604 446.743
R16383 VGND.t840 VGND.t2502 446.743
R16384 VGND.t821 VGND.t2985 446.743
R16385 VGND.t2669 VGND 446.743
R16386 VGND.t3081 VGND 446.743
R16387 VGND.t1907 VGND 446.743
R16388 VGND.t2627 VGND 446.743
R16389 VGND.t607 VGND 446.743
R16390 VGND VGND.t3003 446.743
R16391 VGND VGND.t702 438.315
R16392 VGND VGND.t2276 438.315
R16393 VGND.t964 VGND.t2150 438.315
R16394 VGND.n7314 VGND.t70 438.315
R16395 VGND VGND.t3097 438.315
R16396 VGND.t2583 VGND 438.315
R16397 VGND VGND.t559 438.315
R16398 VGND.t2302 VGND 438.315
R16399 VGND.t447 VGND.t2592 438.315
R16400 VGND.t3017 VGND.n158 438.315
R16401 VGND.t2835 VGND 438.315
R16402 VGND VGND.t3110 438.315
R16403 VGND.n3209 VGND.t2532 438.315
R16404 VGND.t2026 VGND 438.315
R16405 VGND VGND.t2868 429.885
R16406 VGND VGND.t753 429.885
R16407 VGND.n5100 VGND.t757 429.885
R16408 VGND VGND.t2678 429.885
R16409 VGND.t823 VGND.t2984 429.885
R16410 VGND VGND.t2552 429.885
R16411 VGND.t1772 VGND.t372 429.885
R16412 VGND.t352 VGND.t1668 429.885
R16413 VGND.t1403 VGND.t2689 421.457
R16414 VGND.t811 VGND.n6338 421.457
R16415 VGND.t1265 VGND.t492 421.457
R16416 VGND.t2121 VGND.t2954 421.457
R16417 VGND.t982 VGND.t3248 421.457
R16418 VGND.t1510 VGND.t2018 421.457
R16419 VGND.n5814 VGND 420.87
R16420 VGND VGND.t1608 413.027
R16421 VGND VGND.t322 413.027
R16422 VGND VGND.t0 413.027
R16423 VGND.t3053 VGND.t1096 413.027
R16424 VGND.t2736 VGND 413.027
R16425 VGND.t1604 VGND.t562 413.027
R16426 VGND.t2982 VGND.t2121 413.027
R16427 VGND VGND.t2129 413.027
R16428 VGND.t1616 VGND.t827 413.027
R16429 VGND.t817 VGND.t2313 413.027
R16430 VGND.n8254 VGND.t20 413.027
R16431 VGND.t3231 VGND 413.027
R16432 VGND.t354 VGND.t1757 413.027
R16433 VGND.t1176 VGND 409.938
R16434 VGND.n5107 VGND 409.938
R16435 VGND VGND.n5813 409.938
R16436 VGND VGND.n5812 409.938
R16437 VGND VGND.n5811 409.938
R16438 VGND VGND.t2772 404.599
R16439 VGND VGND.t324 404.599
R16440 VGND.n1590 VGND.t121 404.599
R16441 VGND.t2306 VGND.t1291 404.599
R16442 VGND.t277 VGND.t2849 404.599
R16443 VGND.n5099 VGND.t2957 404.599
R16444 VGND VGND.t2901 404.599
R16445 VGND.t767 VGND.t2103 404.599
R16446 VGND.t2572 VGND 404.599
R16447 VGND VGND.t3087 404.599
R16448 VGND.t675 VGND 404.599
R16449 VGND.t3130 VGND.t137 404.599
R16450 VGND.t1619 VGND.t842 404.599
R16451 VGND.t1940 VGND.t167 404.599
R16452 VGND VGND.t1894 404.599
R16453 VGND.t301 VGND.t952 404.599
R16454 VGND.n8338 VGND.t2874 404.599
R16455 VGND.t1892 VGND 404.599
R16456 VGND VGND.t1888 404.599
R16457 VGND.t2801 VGND.t2462 404.599
R16458 VGND VGND.t2027 404.599
R16459 VGND.t2451 VGND 396.17
R16460 VGND VGND.t1601 396.17
R16461 VGND.t819 VGND.t2312 396.17
R16462 VGND VGND.t35 396.17
R16463 VGND.t2769 VGND 396.17
R16464 VGND VGND.t1704 396.17
R16465 VGND.t1194 VGND.t1373 387.74
R16466 VGND.t1519 VGND.n1624 387.74
R16467 VGND.t1490 VGND.n5337 387.74
R16468 VGND.t208 VGND.t444 387.74
R16469 VGND VGND.t2615 387.74
R16470 VGND.t1065 VGND 387.74
R16471 VGND.t1601 VGND 387.74
R16472 VGND.n7684 VGND.t1439 387.74
R16473 VGND.n7812 VGND.t1539 387.74
R16474 VGND.n306 VGND.t3114 387.74
R16475 VGND.t1504 VGND.t1155 387.74
R16476 VGND.t35 VGND 387.74
R16477 VGND VGND.t2769 387.74
R16478 VGND VGND.t2283 387.74
R16479 VGND.t1855 VGND.t2242 387.74
R16480 VGND VGND.t2742 379.31
R16481 VGND VGND.t2754 379.31
R16482 VGND.t452 VGND.t2567 379.31
R16483 VGND.t1789 VGND 379.31
R16484 VGND.t2901 VGND 379.31
R16485 VGND.t580 VGND.t1111 379.31
R16486 VGND VGND.t2304 379.31
R16487 VGND.t2974 VGND.t342 379.31
R16488 VGND.t372 VGND.t1666 379.31
R16489 VGND VGND.t2623 379.31
R16490 VGND.t2141 VGND.t2528 370.882
R16491 VGND.t281 VGND.t2923 370.882
R16492 VGND.n4661 VGND.t3219 370.882
R16493 VGND VGND.t2451 370.882
R16494 VGND.t3252 VGND.n4658 370.882
R16495 VGND.t4 VGND.t1660 370.882
R16496 VGND.t26 VGND.t1664 370.882
R16497 VGND.t2813 VGND.t893 370.882
R16498 VGND VGND.t2111 370.882
R16499 VGND.t2718 VGND.n7313 370.882
R16500 VGND.t3087 VGND 370.882
R16501 VGND.t2582 VGND 370.882
R16502 VGND.n7685 VGND.t3007 370.882
R16503 VGND.t2509 VGND.t1167 370.882
R16504 VGND.t1117 VGND.t482 370.882
R16505 VGND.n7943 VGND.t1712 370.882
R16506 VGND VGND.t88 366.212
R16507 VGND.t753 VGND 362.452
R16508 VGND.t1730 VGND 362.452
R16509 VGND.t186 VGND.t840 362.452
R16510 VGND VGND.t3231 362.452
R16511 VGND.t2072 VGND.t3015 362.452
R16512 VGND VGND.t260 362.452
R16513 VGND.t2462 VGND.t1965 362.452
R16514 VGND.t55 VGND 362.452
R16515 VGND.t376 VGND 360.745
R16516 VGND.t2724 VGND 360.745
R16517 VGND VGND.t2752 355.281
R16518 VGND VGND.t714 355.281
R16519 VGND.t3112 VGND 355.281
R16520 VGND.t2010 VGND 355.281
R16521 VGND.t1900 VGND.t1877 354.024
R16522 VGND.t303 VGND.t2573 354.024
R16523 VGND.t2105 VGND 354.024
R16524 VGND VGND.t3088 354.024
R16525 VGND.t2964 VGND.t3206 354.024
R16526 VGND VGND.t2596 354.024
R16527 VGND.t171 VGND.t793 354.024
R16528 VGND.t161 VGND.t2835 354.024
R16529 VGND.t720 VGND.t619 354.024
R16530 VGND.t496 VGND.t964 345.594
R16531 VGND.t829 VGND 345.594
R16532 VGND.t3084 VGND.t2908 345.594
R16533 VGND.t336 VGND.t2974 345.594
R16534 VGND.t1666 VGND.t366 345.594
R16535 VGND VGND.t1777 345.594
R16536 VGND VGND.t2550 344.349
R16537 VGND.t2911 VGND 344.349
R16538 VGND.t2276 VGND 337.166
R16539 VGND.t2923 VGND.t177 337.166
R16540 VGND.t2461 VGND.n4659 337.166
R16541 VGND.n4658 VGND.t3250 337.166
R16542 VGND VGND.t1729 337.166
R16543 VGND.t1660 VGND.t26 337.166
R16544 VGND.t1719 VGND.t640 337.166
R16545 VGND VGND.t1924 337.166
R16546 VGND.t3157 VGND.n306 337.166
R16547 VGND VGND.t1942 337.166
R16548 VGND.t2219 VGND.t1611 337.166
R16549 VGND VGND.t54 337.166
R16550 VGND.t2238 VGND.t1855 337.166
R16551 VGND.t3003 VGND 337.166
R16552 VGND.t2838 VGND 328.736
R16553 VGND VGND.t179 328.736
R16554 VGND VGND.t1874 328.736
R16555 VGND.t252 VGND 328.736
R16556 VGND VGND.t739 328.736
R16557 VGND VGND.t2250 328.736
R16558 VGND VGND.t2569 328.736
R16559 VGND.t559 VGND 328.736
R16560 VGND.t2312 VGND.t833 328.736
R16561 VGND VGND.t696 328.736
R16562 VGND VGND.t3081 328.736
R16563 VGND.t3227 VGND 328.736
R16564 VGND VGND.t85 328.736
R16565 VGND.t2465 VGND 328.736
R16566 VGND VGND.t607 328.736
R16567 VGND.t3086 VGND.t1495 320.307
R16568 VGND.t316 VGND 320.307
R16569 VGND.t240 VGND 320.307
R16570 VGND.t943 VGND.t1801 320.307
R16571 VGND.t2744 VGND 320.307
R16572 VGND.n4659 VGND.t3121 320.307
R16573 VGND.t764 VGND 320.307
R16574 VGND.t2113 VGND.t767 320.307
R16575 VGND VGND.t677 320.307
R16576 VGND.t2480 VGND 320.307
R16577 VGND.t3009 VGND 320.307
R16578 VGND.t846 VGND.t1619 320.307
R16579 VGND.t613 VGND 320.307
R16580 VGND VGND.t2706 320.307
R16581 VGND VGND.t2318 320.307
R16582 VGND VGND.t2669 320.307
R16583 VGND VGND.t2791 320.307
R16584 VGND.t2180 VGND.t1385 320.307
R16585 VGND.t2704 VGND 320.307
R16586 VGND.t615 VGND 320.307
R16587 VGND.t1288 VGND.t3125 320.307
R16588 VGND VGND.t625 320.307
R16589 VGND.t2127 VGND.t2982 311.877
R16590 VGND.t2125 VGND 311.877
R16591 VGND.t2313 VGND.t819 311.877
R16592 VGND.t1950 VGND.n7811 311.877
R16593 VGND.t1757 VGND.t346 311.877
R16594 VGND VGND.t148 311.877
R16595 VGND VGND.t769 311.877
R16596 VGND VGND.t748 311.877
R16597 VGND VGND.t3145 311.877
R16598 VGND.t2935 VGND 311.877
R16599 VGND.t1703 VGND 311.877
R16600 VGND VGND.t196 311.877
R16601 VGND.n9179 VGND.n20 306.625
R16602 VGND.n9181 VGND.n18 306.625
R16603 VGND.t2687 VGND.t1403 303.449
R16604 VGND VGND.t224 303.449
R16605 VGND.n6338 VGND.t809 303.449
R16606 VGND VGND.t1609 303.449
R16607 VGND VGND.t2166 303.449
R16608 VGND.t490 VGND.t1265 303.449
R16609 VGND.t2954 VGND.t2123 303.449
R16610 VGND VGND.t2575 303.449
R16611 VGND.t3089 VGND.t3130 303.449
R16612 VGND.t842 VGND.t1616 303.449
R16613 VGND VGND.t2928 303.449
R16614 VGND.t3244 VGND.t982 303.449
R16615 VGND.t1963 VGND 303.449
R16616 VGND VGND.t2847 303.449
R16617 VGND.t2022 VGND.t1510 303.449
R16618 VGND.t1860 VGND.t2801 303.449
R16619 VGND VGND.t104 303.449
R16620 VGND.t2879 VGND.t3123 295.019
R16621 VGND VGND.t533 295.019
R16622 VGND VGND.t2768 295.019
R16623 VGND VGND.t2461 295.019
R16624 VGND VGND.t2558 295.019
R16625 VGND VGND.t1638 295.019
R16626 VGND.t66 VGND.t1604 295.019
R16627 VGND.t3088 VGND.n7312 295.019
R16628 VGND.t760 VGND 295.019
R16629 VGND.t2984 VGND.t817 295.019
R16630 VGND VGND.t3205 295.019
R16631 VGND.n7942 VGND.t696 295.019
R16632 VGND.t330 VGND.t1772 295.019
R16633 VGND.t1668 VGND.t354 295.019
R16634 VGND VGND.t2889 295.019
R16635 VGND.t2939 VGND.t712 295.019
R16636 VGND.t157 VGND 295.019
R16637 VGND VGND.t1858 295.019
R16638 VGND VGND.t591 295.019
R16639 VGND.t1495 VGND.t226 286.591
R16640 VGND VGND.t3240 286.591
R16641 VGND.t236 VGND.t943 286.591
R16642 VGND VGND.t111 286.591
R16643 VGND.t8 VGND 286.591
R16644 VGND VGND.t2300 286.591
R16645 VGND.t1385 VGND.t2781 286.591
R16646 VGND VGND.t3171 286.591
R16647 VGND.t629 VGND.t1288 286.591
R16648 VGND.t568 VGND.t722 286.591
R16649 VGND.t413 VGND.t2074 278.161
R16650 VGND VGND.t3131 278.161
R16651 VGND VGND.t1864 278.161
R16652 VGND VGND.t1929 278.161
R16653 VGND VGND.t1921 278.161
R16654 VGND VGND.t2323 278.161
R16655 VGND VGND.t574 278.161
R16656 VGND.t2823 VGND.t2435 278.161
R16657 VGND.t2502 VGND.t844 278.161
R16658 VGND.t2985 VGND.t823 278.161
R16659 VGND.t2170 VGND 278.161
R16660 VGND.t2225 VGND 278.161
R16661 VGND VGND.t2620 278.161
R16662 VGND VGND.t2395 278.161
R16663 VGND VGND.t1589 278.161
R16664 VGND VGND.t2310 269.733
R16665 VGND VGND.t473 269.733
R16666 VGND.t893 VGND.t49 269.733
R16667 VGND.n7314 VGND.t60 269.733
R16668 VGND.t3119 VGND.t2785 269.733
R16669 VGND VGND.t334 269.733
R16670 VGND.t2991 VGND 269.733
R16671 VGND VGND.t27 269.733
R16672 VGND VGND.t2093 269.733
R16673 VGND.t1970 VGND.t1774 269.733
R16674 VGND VGND.t326 269.733
R16675 VGND.t2644 VGND.t344 269.733
R16676 VGND VGND.t2486 269.733
R16677 VGND.t2999 VGND 269.733
R16678 VGND.t3233 VGND 269.733
R16679 VGND.t621 VGND.t2219 269.733
R16680 VGND.t2803 VGND.t2238 269.733
R16681 VGND.t1595 VGND.t2038 269.733
R16682 VGND.t1931 VGND 269.733
R16683 VGND.t3074 VGND 269.733
R16684 VGND VGND.t1621 261.303
R16685 VGND VGND.t778 261.303
R16686 VGND VGND.t194 261.303
R16687 VGND.t1878 VGND 261.303
R16688 VGND.t2431 VGND.t747 261.303
R16689 VGND.t289 VGND 261.303
R16690 VGND.t780 VGND 261.303
R16691 VGND.t3219 VGND 261.303
R16692 VGND VGND.t3128 261.303
R16693 VGND VGND.t3252 261.303
R16694 VGND VGND.t3005 261.303
R16695 VGND VGND.t2032 261.303
R16696 VGND VGND.t1739 261.303
R16697 VGND.t2036 VGND 261.303
R16698 VGND.t165 VGND 261.303
R16699 VGND VGND.t3011 261.303
R16700 VGND VGND.t2185 261.303
R16701 VGND.t1896 VGND 261.303
R16702 VGND.t2511 VGND 261.303
R16703 VGND.t3095 VGND 261.303
R16704 VGND VGND.t1615 261.303
R16705 VGND VGND.t1831 261.303
R16706 VGND.t2758 VGND.t627 261.303
R16707 VGND VGND.t538 261.303
R16708 VGND.t1712 VGND 261.303
R16709 VGND.t2799 VGND.t336 261.303
R16710 VGND VGND.t1629 261.303
R16711 VGND VGND.t2014 261.303
R16712 VGND VGND.t2946 261.303
R16713 VGND.t3062 VGND 261.303
R16714 VGND VGND.t2131 261.303
R16715 VGND.t159 VGND 261.303
R16716 VGND.t3183 VGND 261.303
R16717 VGND VGND.t1769 261.303
R16718 VGND VGND.t92 261.303
R16719 VGND VGND.t3135 261.303
R16720 VGND VGND.t94 261.303
R16721 VGND VGND.t1866 261.303
R16722 VGND.t222 VGND.t1900 252.875
R16723 VGND.t2280 VGND 252.875
R16724 VGND VGND.t770 252.875
R16725 VGND.t1338 VGND.t3209 252.875
R16726 VGND VGND.t2209 252.875
R16727 VGND VGND.t2720 252.875
R16728 VGND VGND.t33 252.875
R16729 VGND VGND.t295 252.875
R16730 VGND VGND.t642 252.875
R16731 VGND.t64 VGND.t1875 252.875
R16732 VGND VGND.t2718 252.875
R16733 VGND VGND.t455 252.875
R16734 VGND.t2793 VGND.t2964 252.875
R16735 VGND VGND.t1723 252.875
R16736 VGND VGND.t453 252.875
R16737 VGND VGND.t3089 252.875
R16738 VGND VGND.t1640 252.875
R16739 VGND.t123 VGND.t1684 252.875
R16740 VGND.t3188 VGND 252.875
R16741 VGND VGND.t486 252.875
R16742 VGND.t3196 VGND 252.875
R16743 VGND.t2339 VGND 252.875
R16744 VGND VGND.t291 252.875
R16745 VGND.t146 VGND.t589 252.875
R16746 VGND VGND.t798 252.875
R16747 VGND.t2693 VGND.t720 252.875
R16748 VGND VGND.t1519 244.445
R16749 VGND.t1234 VGND 244.445
R16750 VGND VGND.t1490 244.445
R16751 VGND VGND.t1966 244.445
R16752 VGND.t2488 VGND 244.445
R16753 VGND.t1473 VGND 244.445
R16754 VGND.t1012 VGND 244.445
R16755 VGND.t1862 VGND 244.445
R16756 VGND.t426 VGND.t1851 244.445
R16757 VGND VGND.t1143 244.445
R16758 VGND.t700 VGND.t2205 244.445
R16759 VGND.t2827 VGND.t2433 244.445
R16760 VGND VGND.t994 244.445
R16761 VGND VGND.t1465 244.445
R16762 VGND.t2289 VGND.t2600 244.445
R16763 VGND.t18 VGND.t2288 244.445
R16764 VGND.t1638 VGND.t2355 244.445
R16765 VGND.t2115 VGND.t2507 244.445
R16766 VGND.t2123 VGND 244.445
R16767 VGND.t665 VGND 244.445
R16768 VGND VGND.t2936 244.445
R16769 VGND VGND.t1439 244.445
R16770 VGND.t1346 VGND 244.445
R16771 VGND.t1539 VGND 244.445
R16772 VGND VGND.t1303 244.445
R16773 VGND.t480 VGND 244.445
R16774 VGND.t3068 VGND.t2072 244.445
R16775 VGND.t478 VGND 244.445
R16776 VGND.t1370 VGND 244.445
R16777 VGND.t940 VGND 244.445
R16778 VGND.t911 VGND 244.445
R16779 VGND.t1470 VGND 244.445
R16780 VGND VGND.t1018 244.445
R16781 VGND.t2268 VGND.t2704 244.445
R16782 VGND VGND.t202 244.445
R16783 VGND VGND.t1546 244.445
R16784 VGND VGND.t1093 244.445
R16785 VGND VGND.t887 244.445
R16786 VGND VGND.t1432 244.445
R16787 VGND.t2370 VGND.t2415 236.016
R16788 VGND.t2837 VGND.t2498 236.016
R16789 VGND.t68 VGND.t2372 236.016
R16790 VGND.t2561 VGND.t2099 236.016
R16791 VGND.t2993 VGND.t681 236.016
R16792 VGND VGND.t3102 236.016
R16793 VGND.t2278 VGND.t1202 236.016
R16794 VGND VGND.t3239 236.016
R16795 VGND.t3198 VGND 236.016
R16796 VGND.t346 VGND 236.016
R16797 VGND.t1933 VGND.t2223 236.016
R16798 VGND.t86 VGND.t3029 236.016
R16799 VGND VGND.t1006 236.016
R16800 VGND.t1808 VGND.t1703 236.016
R16801 VGND VGND.t2691 227.587
R16802 VGND VGND.t287 227.587
R16803 VGND VGND.t130 227.587
R16804 VGND.t2076 VGND 227.587
R16805 VGND.t409 VGND 227.587
R16806 VGND.t471 VGND 227.587
R16807 VGND VGND.t2883 227.587
R16808 VGND VGND.t3211 227.587
R16809 VGND VGND.t273 227.587
R16810 VGND VGND.t708 227.587
R16811 VGND VGND.t2297 227.587
R16812 VGND VGND.t1980 227.587
R16813 VGND VGND.t1954 227.587
R16814 VGND VGND.t645 227.587
R16815 VGND.t644 VGND.t398 227.587
R16816 VGND.t1111 VGND.t1916 227.587
R16817 VGND.t2815 VGND.t305 227.587
R16818 VGND VGND.t494 227.587
R16819 VGND.t453 VGND.t669 227.587
R16820 VGND.t2211 VGND 227.587
R16821 VGND.t2308 VGND.t613 227.587
R16822 VGND VGND.t1761 227.587
R16823 VGND.t484 VGND.t391 227.587
R16824 VGND VGND.t2919 227.587
R16825 VGND VGND.t2893 227.587
R16826 VGND.t2387 VGND 227.587
R16827 VGND VGND.t3242 227.587
R16828 VGND VGND.t2020 227.587
R16829 VGND.t1282 VGND.t155 227.587
R16830 VGND VGND.t1804 227.587
R16831 VGND VGND.t1591 227.587
R16832 VGND VGND.t2776 227.587
R16833 VGND VGND.t2064 227.587
R16834 VGND.t2631 VGND.t405 219.157
R16835 VGND.t815 VGND 219.157
R16836 VGND.n6354 VGND.t2695 219.157
R16837 VGND.n6976 VGND.t0 219.157
R16838 VGND.t256 VGND.t208 219.157
R16839 VGND.t2144 VGND.t2109 219.157
R16840 VGND VGND.t3084 219.157
R16841 VGND.t299 VGND.t2584 219.157
R16842 VGND.t2555 VGND.t2553 219.157
R16843 VGND.t1888 VGND 219.157
R16844 VGND.t2263 VGND.t1182 219.157
R16845 VGND.t3039 VGND 219.157
R16846 VGND.t1070 VGND.t1937 219.157
R16847 VGND.t443 VGND 219.157
R16848 VGND VGND.t2921 219.157
R16849 VGND VGND.t2264 219.157
R16850 VGND.t955 VGND.t2966 219.157
R16851 VGND.n6019 VGND.t2880 215.036
R16852 VGND.n4892 VGND.t9 215.036
R16853 VGND.n4163 VGND.t1610 215.036
R16854 VGND.n4420 VGND.t1852 215.036
R16855 VGND.n2675 VGND.t2848 215.036
R16856 VGND.n8970 VGND.t1964 215.036
R16857 VGND.n8456 VGND.t3146 215.036
R16858 VGND.n7958 VGND.t2645 215.036
R16859 VGND.n357 VGND.t2929 215.036
R16860 VGND.n921 VGND.t1613 215.036
R16861 VGND.n811 VGND.t1639 215.036
R16862 VGND.n9130 VGND.t197 215.036
R16863 VGND.n1445 VGND.t2434 214.488
R16864 VGND.n1534 VGND.t3241 214.488
R16865 VGND.n2350 VGND.t2826 211.738
R16866 VGND.n2496 VGND.t2218 211.738
R16867 VGND.n5207 VGND.t395 211.738
R16868 VGND.n6647 VGND.t3148 211.738
R16869 VGND.n7024 VGND.t2400 211.738
R16870 VGND.n4080 VGND.t2082 211.738
R16871 VGND.n4235 VGND.t1905 211.738
R16872 VGND.n2923 VGND.t2161 211.738
R16873 VGND.n2750 VGND.t156 211.738
R16874 VGND.n3221 VGND.t2053 211.738
R16875 VGND.n3124 VGND.t1588 211.738
R16876 VGND.n9015 VGND.t170 211.738
R16877 VGND.n8746 VGND.t1600 211.738
R16878 VGND.n8609 VGND.t2877 211.738
R16879 VGND.n7900 VGND.t1707 211.738
R16880 VGND.n7659 VGND.t2230 211.738
R16881 VGND.n8156 VGND.t2057 211.738
R16882 VGND.n8303 VGND.t2335 211.738
R16883 VGND.n1156 VGND.t2436 211.738
R16884 VGND.n6300 VGND.t2438 211.738
R16885 VGND.n6405 VGND.t2697 211.738
R16886 VGND.n6388 VGND.t692 211.738
R16887 VGND.t1877 VGND 210.728
R16888 VGND.t1906 VGND 210.728
R16889 VGND.t2476 VGND.t1170 210.728
R16890 VGND.t2401 VGND.t2254 210.728
R16891 VGND.t2492 VGND.t1445 210.728
R16892 VGND.t106 VGND.t2977 210.728
R16893 VGND.t1513 VGND.t220 210.728
R16894 VGND.t2722 VGND.t115 210.728
R16895 VGND.t70 VGND 210.728
R16896 VGND.t2878 VGND.t2867 210.728
R16897 VGND.t3206 VGND 210.728
R16898 VGND.t1021 VGND.t1692 210.728
R16899 VGND VGND.t2282 210.728
R16900 VGND VGND.t2832 210.728
R16901 VGND.t1090 VGND.t2789 210.728
R16902 VGND.t125 VGND.t689 210.728
R16903 VGND VGND.t2656 210.728
R16904 VGND VGND.t133 210.728
R16905 VGND.t2441 VGND 210.728
R16906 VGND.t3225 VGND.t2246 202.299
R16907 VGND.t2336 VGND.t1730 202.299
R16908 VGND.t581 VGND.t2139 202.299
R16909 VGND VGND.t10 202.299
R16910 VGND.t1872 VGND.t293 202.299
R16911 VGND VGND.t1821 202.299
R16912 VGND.t1164 VGND.t2197 202.299
R16913 VGND.t27 VGND.t1612 202.299
R16914 VGND.t831 VGND.t2500 202.299
R16915 VGND.t3186 VGND.t3185 202.299
R16916 VGND.t1161 VGND.t269 202.299
R16917 VGND.t3143 VGND.t718 202.299
R16918 VGND.n3658 VGND.t3458 200.476
R16919 VGND.n3400 VGND.t3438 200.149
R16920 VGND.n8727 VGND.t3388 200.114
R16921 VGND.n7162 VGND.t588 197.79
R16922 VGND.n7181 VGND.t537 197.79
R16923 VGND.n7218 VGND.t1718 197.79
R16924 VGND.n4510 VGND.t2025 197.79
R16925 VGND.n7884 VGND.t2739 197.79
R16926 VGND.n7594 VGND.t100 197.79
R16927 VGND VGND.t2349 193.87
R16928 VGND VGND.t3126 193.87
R16929 VGND VGND.t3200 193.87
R16930 VGND VGND.t2580 193.87
R16931 VGND.t2909 VGND.t829 193.87
R16932 VGND VGND.t22 193.87
R16933 VGND.t1125 VGND.t432 193.87
R16934 VGND VGND.t1617 193.87
R16935 VGND VGND.t53 193.87
R16936 VGND.t82 VGND 193.87
R16937 VGND.t1611 VGND 193.87
R16938 VGND VGND.t3076 193.87
R16939 VGND VGND.t590 193.87
R16940 VGND.t2191 VGND.t55 193.87
R16941 VGND.t3072 VGND.t2042 193.87
R16942 VGND.n2646 VGND.t3498 193.488
R16943 VGND.n100 VGND.t3418 193.488
R16944 VGND.n3638 VGND.t3290 193.44
R16945 VGND.n1343 VGND.t2896 192.944
R16946 VGND.n1106 VGND.t2287 190.681
R16947 VGND.n1343 VGND.t2096 190.316
R16948 VGND.n4220 VGND.t427 190.316
R16949 VGND.n4631 VGND.t705 190.065
R16950 VGND.n479 VGND.t388 190.065
R16951 VGND.n1030 VGND.t565 190.065
R16952 VGND.n1581 VGND.t3060 190.065
R16953 VGND.n6829 VGND.t1960 190.065
R16954 VGND.n6688 VGND.t3440 189.316
R16955 VGND.n3456 VGND.t3397 189.316
R16956 VGND.n8699 VGND.t3257 189.316
R16957 VGND.n7675 VGND.t3381 189.316
R16958 VGND.n3033 VGND.t3376 189.308
R16959 VGND.n9184 VGND.t3357 189.298
R16960 VGND.n3428 VGND.t3273 189.298
R16961 VGND.n1292 VGND.t3336 189.298
R16962 VGND.n178 VGND.t3431 189.095
R16963 VGND.n2864 VGND.t3077 188.75
R16964 VGND.n2790 VGND.t1859 188.75
R16965 VGND.n3043 VGND.t158 188.75
R16966 VGND.n8348 VGND.t1632 188.75
R16967 VGND.n917 VGND.t3100 188.75
R16968 VGND.n5027 VGND.t2143 188.175
R16969 VGND.n152 VGND.t766 188.01
R16970 VGND.n3485 VGND.t3500 186.784
R16971 VGND.n3487 VGND.t3259 186.784
R16972 VGND.n7 VGND.t3472 186.784
R16973 VGND.n5234 VGND.t3327 186.784
R16974 VGND.n5236 VGND.t3346 186.784
R16975 VGND.n1711 VGND.t3281 186.784
R16976 VGND.n1713 VGND.t3306 186.784
R16977 VGND.n7012 VGND.t3478 186.784
R16978 VGND.n7014 VGND.t3295 186.784
R16979 VGND.n4767 VGND.t3429 186.784
R16980 VGND.n4768 VGND.t3503 186.784
R16981 VGND.n1409 VGND.t3480 186.784
R16982 VGND.n1411 VGND.t3490 186.784
R16983 VGND.n4099 VGND.t3437 186.784
R16984 VGND.n4100 VGND.t3446 186.784
R16985 VGND.n2908 VGND.t3493 186.784
R16986 VGND.n2909 VGND.t3501 186.784
R16987 VGND.n2048 VGND.t3423 186.784
R16988 VGND.n2050 VGND.t3430 186.784
R16989 VGND.n2681 VGND.t3415 186.784
R16990 VGND.n2682 VGND.t3324 186.784
R16991 VGND.n3670 VGND.t3355 186.784
R16992 VGND.n3672 VGND.t3280 186.784
R16993 VGND.n8915 VGND.t3298 186.784
R16994 VGND.n8462 VGND.t3320 186.784
R16995 VGND.n8464 VGND.t3329 186.784
R16996 VGND.n3779 VGND.t3278 186.784
R16997 VGND.n3780 VGND.t3283 186.784
R16998 VGND.n8353 VGND.t3502 186.784
R16999 VGND.n8355 VGND.t3508 186.784
R17000 VGND.n1884 VGND.t3463 186.784
R17001 VGND.n1885 VGND.t3466 186.784
R17002 VGND.n349 VGND.t3424 186.784
R17003 VGND.n350 VGND.t3436 186.784
R17004 VGND.n692 VGND.t3383 186.784
R17005 VGND.n693 VGND.t3394 186.784
R17006 VGND.n929 VGND.t3300 186.784
R17007 VGND.n930 VGND.t3363 186.784
R17008 VGND.n7459 VGND.t3505 186.784
R17009 VGND.n7461 VGND.t3322 186.784
R17010 VGND.n1490 VGND.t3405 186.784
R17011 VGND.n1492 VGND.t3413 186.784
R17012 VGND.n1588 VGND.t3468 186.784
R17013 VGND.n6117 VGND.t3364 186.784
R17014 VGND.n6119 VGND.t3372 186.784
R17015 VGND.n9119 VGND.t3313 186.784
R17016 VGND.n9120 VGND.t3331 186.784
R17017 VGND.n2424 VGND.t3407 186.719
R17018 VGND.n2295 VGND.t3356 186.719
R17019 VGND.n2601 VGND.t3482 186.719
R17020 VGND.n2606 VGND.t3469 186.719
R17021 VGND.n2230 VGND.t3325 186.719
R17022 VGND.n2218 VGND.t3294 186.719
R17023 VGND.n2206 VGND.t3433 186.719
R17024 VGND.n9189 VGND.t3302 186.719
R17025 VGND.n5171 VGND.t3416 186.719
R17026 VGND.n5718 VGND.t3442 186.719
R17027 VGND.n5518 VGND.t3481 186.719
R17028 VGND.n5909 VGND.t3304 186.719
R17029 VGND.n5949 VGND.t3311 186.719
R17030 VGND.n5247 VGND.t3487 186.719
R17031 VGND.n5269 VGND.t3368 186.719
R17032 VGND.n5269 VGND.t3391 186.719
R17033 VGND.n5443 VGND.t3305 186.719
R17034 VGND.n5435 VGND.t3467 186.719
R17035 VGND.n5389 VGND.t3398 186.719
R17036 VGND.n5361 VGND.t3262 186.719
R17037 VGND.n6717 VGND.t3315 186.719
R17038 VGND.n1643 VGND.t3296 186.719
R17039 VGND.n6601 VGND.t3287 186.719
R17040 VGND.n7027 VGND.t3384 186.719
R17041 VGND.n7053 VGND.t3261 186.719
R17042 VGND.n4938 VGND.t3361 186.719
R17043 VGND.n4267 VGND.t3285 186.719
R17044 VGND.n4539 VGND.t3293 186.719
R17045 VGND.n3433 VGND.t3479 186.719
R17046 VGND.n3405 VGND.t3350 186.719
R17047 VGND.n3383 VGND.t3495 186.719
R17048 VGND.n3307 VGND.t3264 186.719
R17049 VGND.n2655 VGND.t3255 186.719
R17050 VGND.n3123 VGND.t3370 186.719
R17051 VGND.n3094 VGND.t3486 186.719
R17052 VGND.n3647 VGND.t3404 186.719
R17053 VGND.n91 VGND.t3380 186.719
R17054 VGND.n8861 VGND.t3402 186.719
R17055 VGND.n9001 VGND.t3310 186.719
R17056 VGND.n3864 VGND.t3484 186.719
R17057 VGND.n7771 VGND.t3299 186.719
R17058 VGND.n7822 VGND.t3386 186.719
R17059 VGND.n335 VGND.t3387 186.719
R17060 VGND.n7574 VGND.t3291 186.719
R17061 VGND.n7656 VGND.t3403 186.719
R17062 VGND.n8170 VGND.t3497 186.719
R17063 VGND.n8300 VGND.t3362 186.719
R17064 VGND.n1127 VGND.t3378 186.719
R17065 VGND.n7361 VGND.t3421 186.719
R17066 VGND.n7394 VGND.t3333 186.719
R17067 VGND.n1508 VGND.t3288 186.719
R17068 VGND.n1501 VGND.t3326 186.719
R17069 VGND.n6883 VGND.t3337 186.719
R17070 VGND.n6848 VGND.t3473 186.719
R17071 VGND.n1593 VGND.t3374 186.719
R17072 VGND.n6312 VGND.t3352 186.719
R17073 VGND.n2900 VGND.t2858 185.452
R17074 VGND.n8452 VGND.t3065 185.452
R17075 VGND.n7831 VGND.t1618 185.452
R17076 VGND.n1022 VGND.t2373 185.452
R17077 VGND.t532 VGND.t192 185.441
R17078 VGND.t2742 VGND.t1816 185.441
R17079 VGND.t47 VGND.t2496 185.441
R17080 VGND.t2863 VGND.t2478 185.441
R17081 VGND.t383 VGND.t599 185.441
R17082 VGND VGND.t1982 185.441
R17083 VGND.t2032 VGND.t1917 185.441
R17084 VGND VGND.t2821 185.441
R17085 VGND VGND.t744 185.441
R17086 VGND.t1723 VGND.t308 185.441
R17087 VGND.t673 VGND 185.441
R17088 VGND.t835 VGND.t2505 185.441
R17089 VGND VGND.t805 185.441
R17090 VGND.t2588 VGND 185.441
R17091 VGND.t1676 VGND.t2999 185.441
R17092 VGND.t2532 VGND 185.441
R17093 VGND.t2266 VGND.t693 185.441
R17094 VGND.n1979 VGND.t2554 185.225
R17095 VGND.n3959 VGND.t2684 184.713
R17096 VGND.n5018 VGND.t1661 184.661
R17097 VGND.n4171 VGND.t1734 184.424
R17098 VGND.n8171 VGND.t390 184.424
R17099 VGND.n2400 VGND.t3258 183.082
R17100 VGND.n2475 VGND.t3443 183.082
R17101 VGND.n5135 VGND.t3494 183.082
R17102 VGND.n5738 VGND.t3289 183.082
R17103 VGND.n5593 VGND.t3297 183.082
R17104 VGND.n1856 VGND.t3349 183.082
R17105 VGND.n1803 VGND.t3369 183.082
R17106 VGND.n1628 VGND.t3339 183.082
R17107 VGND.n1709 VGND.t3373 183.082
R17108 VGND.n1345 VGND.t3492 183.082
R17109 VGND.n4035 VGND.t3282 183.082
R17110 VGND.n5048 VGND.t3312 183.082
R17111 VGND.n4238 VGND.t3451 183.082
R17112 VGND.n4452 VGND.t3417 183.082
R17113 VGND.n4653 VGND.t3432 183.082
R17114 VGND.n2903 VGND.t3396 183.082
R17115 VGND.n2046 VGND.t3254 183.082
R17116 VGND.n3668 VGND.t3441 183.082
R17117 VGND.n8889 VGND.t3371 183.082
R17118 VGND.n3796 VGND.t3344 183.082
R17119 VGND.n224 VGND.t3274 183.082
R17120 VGND.n1900 VGND.t3360 183.082
R17121 VGND.n495 VGND.t3316 183.082
R17122 VGND.n7741 VGND.t3338 183.082
R17123 VGND.n7842 VGND.t3332 183.082
R17124 VGND.n903 VGND.t3428 183.082
R17125 VGND.n7336 VGND.t3471 183.082
R17126 VGND.n7457 VGND.t3345 183.082
R17127 VGND.n6260 VGND.t3411 183.082
R17128 VGND.n6352 VGND.t3271 183.082
R17129 VGND.n6358 VGND.t3348 183.082
R17130 VGND.n1931 VGND.t46 182.812
R17131 VGND.n3797 VGND.t3082 182.792
R17132 VGND.n504 VGND.t3232 182.792
R17133 VGND.n6623 VGND.t3454 182.177
R17134 VGND.n7405 VGND.t2384 182.117
R17135 VGND.n7416 VGND.t2677 182.117
R17136 VGND.n8533 VGND.t3158 178.84
R17137 VGND.n1337 VGND.t2820 178.619
R17138 VGND.n517 VGND.t97 177.47
R17139 VGND.n2657 VGND.t3366 177.029
R17140 VGND.n233 VGND.t3256 177.029
R17141 VGND.t198 VGND.t238 177.012
R17142 VGND.t2411 VGND.t2330 177.012
R17143 VGND VGND.t1667 177.012
R17144 VGND.t1633 VGND.t2988 177.012
R17145 VGND.t2807 VGND.n78 177.012
R17146 VGND.t602 VGND.t2040 177.012
R17147 VGND.n7205 VGND.t2294 170.963
R17148 VGND.n4009 VGND.t741 170.963
R17149 VGND.t418 VGND 169.441
R17150 VGND VGND.t1725 169.441
R17151 VGND.t2277 VGND.t878 168.583
R17152 VGND.t2231 VGND.t1208 168.583
R17153 VGND VGND.t3013 168.583
R17154 VGND.t212 VGND.t3229 168.583
R17155 VGND.t1481 VGND.t1974 168.583
R17156 VGND.t697 VGND.t1364 168.583
R17157 VGND.t1766 VGND.t362 168.583
R17158 VGND VGND.t498 168.583
R17159 VGND.t2726 VGND.t1358 168.583
R17160 VGND.t1335 VGND.t2836 168.583
R17161 VGND.t2708 VGND.t109 168.583
R17162 VGND.t3111 VGND.t1330 168.583
R17163 VGND.t925 VGND.t2628 168.583
R17164 VGND.t2285 VGND.n9180 168.583
R17165 VGND.n4034 VGND.t2721 167.011
R17166 VGND.n8901 VGND.t3308 163.852
R17167 VGND.n1331 VGND.t2723 160.512
R17168 VGND VGND.t3192 160.154
R17169 VGND.t3147 VGND.t441 160.154
R17170 VGND.t2073 VGND 160.154
R17171 VGND.t691 VGND.t991 160.154
R17172 VGND VGND.t3177 160.154
R17173 VGND VGND.t2673 160.154
R17174 VGND.t2119 VGND.t1620 160.154
R17175 VGND VGND.t1714 160.154
R17176 VGND.t499 VGND.t1487 160.154
R17177 VGND.t3181 VGND 160.154
R17178 VGND.t2607 VGND 160.154
R17179 VGND.n7100 VGND.t1722 157.835
R17180 VGND.n4037 VGND.t19 154.006
R17181 VGND.n4765 VGND.t1871 154.006
R17182 VGND.n4386 VGND.t1881 154.006
R17183 VGND.n3268 VGND.t1861 154.006
R17184 VGND.n8952 VGND.t162 154.006
R17185 VGND.n8341 VGND.t1776 154.006
R17186 VGND.n1920 VGND.t2173 154.006
R17187 VGND.n7605 VGND.t3230 154.006
R17188 VGND.n1158 VGND.t2904 154.006
R17189 VGND.n6108 VGND.t129 154.006
R17190 VGND.n6108 VGND.t2841 154.006
R17191 VGND VGND.t1042 151.725
R17192 VGND.t2429 VGND.t401 151.725
R17193 VGND.n4660 VGND.t2865 151.725
R17194 VGND.t420 VGND.t2643 151.725
R17195 VGND.t2201 VGND.t536 151.725
R17196 VGND.t2184 VGND.t2564 151.725
R17197 VGND.t808 VGND.t2511 151.725
R17198 VGND.t190 VGND.t2174 151.725
R17199 VGND.t3033 VGND.t439 151.725
R17200 VGND.t1741 VGND.t2134 151.725
R17201 VGND.t2671 VGND.t2761 151.725
R17202 VGND.t2969 VGND.t2833 151.725
R17203 VGND.t291 VGND.t1701 151.725
R17204 VGND.n3489 VGND.t2346 150.786
R17205 VGND.n3489 VGND.t2155 150.786
R17206 VGND.n2472 VGND.t2045 150.786
R17207 VGND.n2560 VGND.t2241 150.786
R17208 VGND.n5663 VGND.t1847 150.786
R17209 VGND.n5572 VGND.t1782 150.786
R17210 VGND.n4784 VGND.t2249 150.786
R17211 VGND.n3778 VGND.t2670 150.786
R17212 VGND.n928 VGND.t2522 150.786
R17213 VGND.n6121 VGND.t1995 150.786
R17214 VGND.n6121 VGND.t3138 150.786
R17215 VGND.n1670 VGND.t810 150.786
R17216 VGND.n9111 VGND.t723 150.786
R17217 VGND.n9118 VGND.t2446 150.786
R17218 VGND.n7984 VGND.t375 149.567
R17219 VGND.n663 VGND.t841 149.567
R17220 VGND.n6445 VGND.t2422 149.567
R17221 VGND.n2401 VGND.t2856 149.471
R17222 VGND.n2342 VGND.t3073 149.471
R17223 VGND.n1649 VGND.t2075 149.471
R17224 VGND.n4554 VGND.t701 149.471
R17225 VGND.n2666 VGND.t3067 149.471
R17226 VGND.n242 VGND.t3160 149.471
R17227 VGND.n689 VGND.t2190 149.471
R17228 VGND.n982 VGND.t2992 149.471
R17229 VGND.n7806 VGND.t2365 148.808
R17230 VGND.n451 VGND.t3085 148.448
R17231 VGND.n6350 VGND.t323 148.448
R17232 VGND.n1619 VGND.t3425 148.102
R17233 VGND.n4439 VGND.t2577 148.075
R17234 VGND.n3785 VGND.t2015 148.075
R17235 VGND.n5451 VGND.t3303 147.107
R17236 VGND.n1715 VGND.t2688 146.9
R17237 VGND.n1407 VGND.t2165 146.9
R17238 VGND.n2052 VGND.t2023 146.9
R17239 VGND.n3674 VGND.t3245 146.9
R17240 VGND.n220 VGND.t3030 146.9
R17241 VGND.n8352 VGND.t2317 146.9
R17242 VGND.n8344 VGND.t521 146.9
R17243 VGND.n7463 VGND.t491 146.9
R17244 VGND.n6871 VGND.t3058 146.48
R17245 VGND.n167 VGND.t790 146.356
R17246 VGND.n3978 VGND.t461 146.272
R17247 VGND.n4436 VGND.t3129 146.058
R17248 VGND.n1639 VGND.t3265 145.972
R17249 VGND.n1921 VGND.t3385 145.958
R17250 VGND.n9165 VGND.t3483 145.958
R17251 VGND.n1194 VGND.t662 145.94
R17252 VGND.n1031 VGND.t2106 145.94
R17253 VGND.n613 VGND.t2910 145.811
R17254 VGND.n4904 VGND.t3176 145.583
R17255 VGND.n788 VGND.t1887 145.036
R17256 VGND.n448 VGND.t3426 144.952
R17257 VGND.n7951 VGND.t327 144.881
R17258 VGND.n1253 VGND.t335 144.881
R17259 VGND.n4170 VGND.t3253 143.998
R17260 VGND.n7479 VGND.t3191 143.498
R17261 VGND.t324 VGND.t283 143.296
R17262 VGND.t3055 VGND 143.296
R17263 VGND.t2979 VGND.t1834 143.296
R17264 VGND.t1096 VGND 143.296
R17265 VGND.t2849 VGND 143.296
R17266 VGND.n5101 VGND 143.296
R17267 VGND.t2963 VGND.t2870 143.296
R17268 VGND.t2261 VGND.t1717 143.296
R17269 VGND.t1276 VGND 143.296
R17270 VGND.t3099 VGND.t2583 143.296
R17271 VGND.t2734 VGND 143.296
R17272 VGND.t2659 VGND 143.296
R17273 VGND.t1315 VGND 143.296
R17274 VGND.n3980 VGND.t460 143.296
R17275 VGND.t1670 VGND 143.296
R17276 VGND.t1819 VGND.t1623 143.296
R17277 VGND VGND.t979 143.296
R17278 VGND.t2634 VGND.t204 143.296
R17279 VGND VGND.t1188 143.296
R17280 VGND.n3207 VGND 143.296
R17281 VGND.n1882 VGND.t2612 143.107
R17282 VGND.n3929 VGND.t153 142.871
R17283 VGND.n2509 VGND.t3427 142.308
R17284 VGND.n2345 VGND.t3263 142.308
R17285 VGND.n2307 VGND.t3399 142.308
R17286 VGND.n2178 VGND.t3400 142.308
R17287 VGND.n5496 VGND.t3354 142.308
R17288 VGND.n1799 VGND.t3317 142.308
R17289 VGND.n1736 VGND.t3395 142.308
R17290 VGND.n7111 VGND.t3455 142.308
R17291 VGND.n4085 VGND.t3268 142.308
R17292 VGND.n4865 VGND.t3367 142.308
R17293 VGND.n1415 VGND.t3390 142.308
R17294 VGND.n4149 VGND.t3409 142.308
R17295 VGND.n4688 VGND.t3314 142.308
R17296 VGND.n4667 VGND.t3393 142.308
R17297 VGND.n4302 VGND.t3452 142.308
R17298 VGND.n4509 VGND.t3461 142.308
R17299 VGND.n2749 VGND.t3340 142.308
R17300 VGND.n2833 VGND.t3464 142.308
R17301 VGND.n2785 VGND.t3334 142.308
R17302 VGND.n3064 VGND.t3379 142.308
R17303 VGND.n8471 VGND.t3489 142.308
R17304 VGND.n8487 VGND.t3392 142.308
R17305 VGND.n8759 VGND.t3491 142.308
R17306 VGND.n187 VGND.t3422 142.308
R17307 VGND.n1880 VGND.t3347 142.308
R17308 VGND.n7946 VGND.t3485 142.308
R17309 VGND.n7851 VGND.t3414 142.308
R17310 VGND.n8087 VGND.t3476 142.308
R17311 VGND.n396 VGND.t3266 142.308
R17312 VGND.n7616 VGND.t3260 142.308
R17313 VGND.n1006 VGND.t3353 142.308
R17314 VGND.n6857 VGND.t122 141.946
R17315 VGND.n6053 VGND.t42 141.739
R17316 VGND.n6583 VGND.t1969 141.739
R17317 VGND.n4870 VGND.t773 141.739
R17318 VGND.n4472 VGND.t384 141.739
R17319 VGND.n2716 VGND.t110 141.739
R17320 VGND.n1692 VGND.t2658 141.739
R17321 VGND.n165 VGND.t1650 141.232
R17322 VGND.n2942 VGND.t3044 140.959
R17323 VGND.n2857 VGND.t3038 140.959
R17324 VGND.n8502 VGND.t3050 140.959
R17325 VGND.n8346 VGND.t3048 140.959
R17326 VGND.n8573 VGND.t3052 140.631
R17327 VGND.n4432 VGND.t3343 139.754
R17328 VGND.n1924 VGND.t3496 139.754
R17329 VGND.n2796 VGND.t3046 139.725
R17330 VGND.n1053 VGND.t2216 138.477
R17331 VGND.n3806 VGND.t73 137.988
R17332 VGND.n3035 VGND.t3040 137.734
R17333 VGND.n7825 VGND.t182 137.333
R17334 VGND.n916 VGND.t3042 137.333
R17335 VGND.n1016 VGND.t1605 137.333
R17336 VGND.t258 VGND.t780 134.867
R17337 VGND.t1653 VGND.t139 134.867
R17338 VGND.t737 VGND.t742 134.867
R17339 VGND.t740 VGND.t2291 134.867
R17340 VGND.t667 VGND.t3237 134.867
R17341 VGND.n8253 VGND.t2756 134.867
R17342 VGND VGND.t1912 134.867
R17343 VGND.t2508 VGND.t1972 134.867
R17344 VGND.t364 VGND.t795 134.867
R17345 VGND.t3228 VGND.t2225 134.867
R17346 VGND.n2648 VGND.t1485 134.756
R17347 VGND.n1089 VGND.t339 134.397
R17348 VGND.n4910 VGND.t3180 134.382
R17349 VGND.n4111 VGND.t1628 134.382
R17350 VGND.n4384 VGND.t2978 134.382
R17351 VGND.n4613 VGND.t2916 134.382
R17352 VGND.n2661 VGND.t3184 134.382
R17353 VGND.n8972 VGND.t2514 134.382
R17354 VGND.n7872 VGND.t1832 134.382
R17355 VGND.n454 VGND.t1941 134.382
R17356 VGND.n1284 VGND.t3012 134.382
R17357 VGND.n1582 VGND.t517 134.382
R17358 VGND.n8267 VGND.t783 131.998
R17359 VGND.n166 VGND.t1648 131.714
R17360 VGND.n7382 VGND.t166 131.291
R17361 VGND.n2453 VGND.t799 131.248
R17362 VGND.n8896 VGND.t1505 130.938
R17363 VGND.n2301 VGND.t610 130.815
R17364 VGND.n5377 VGND.t2649 130.815
R17365 VGND.n1735 VGND.t3195 130.815
R17366 VGND.n1650 VGND.t414 130.815
R17367 VGND.n7005 VGND.t2931 130.815
R17368 VGND.n4791 VGND.t545 130.815
R17369 VGND.n4167 VGND.t3220 130.815
R17370 VGND.n2898 VGND.t2086 130.815
R17371 VGND.n2818 VGND.t2458 130.815
R17372 VGND.n2721 VGND.t2810 130.815
R17373 VGND.n3087 VGND.t2747 130.815
R17374 VGND.n8932 VGND.t2764 130.815
R17375 VGND.n8520 VGND.t1979 130.815
R17376 VGND.n213 VGND.t438 130.815
R17377 VGND.n8041 VGND.t1713 130.815
R17378 VGND.n334 VGND.t2733 130.815
R17379 VGND.n7686 VGND.t3008 130.815
R17380 VGND.n6796 VGND.t553 130.815
R17381 VGND.n6249 VGND.t215 130.815
R17382 VGND.n6449 VGND.t404 130.815
R17383 VGND.n1629 VGND.t1374 129.293
R17384 VGND.n6618 VGND.t950 127.472
R17385 VGND.n2576 VGND.t1329 127.406
R17386 VGND.t746 VGND.t2425 126.438
R17387 VGND.t2413 VGND.t2331 126.438
R17388 VGND.t396 VGND.t400 126.438
R17389 VGND.t2377 VGND.t387 126.438
R17390 VGND VGND.t370 126.438
R17391 VGND VGND.t710 126.438
R17392 VGND.t261 VGND.t3031 126.438
R17393 VGND.t3110 VGND.t469 126.438
R17394 VGND.t973 VGND.t2855 126.438
R17395 VGND.n5418 VGND.t935 125.927
R17396 VGND.n2596 VGND.t1089 125.478
R17397 VGND.n6675 VGND.t1195 125.478
R17398 VGND.n5341 VGND.t960 125.478
R17399 VGND.n5450 VGND.t865 125.454
R17400 VGND.n1922 VGND.t1380 125.433
R17401 VGND.n9166 VGND.t938 125.433
R17402 VGND.n2289 VGND.t1328 125.391
R17403 VGND.n5375 VGND.t1171 125.391
R17404 VGND.n6705 VGND.t1455 125.391
R17405 VGND.n182 VGND.t1174 125.391
R17406 VGND.n2109 VGND.t1530 125.368
R17407 VGND.n3283 VGND.t1556 125.368
R17408 VGND.n8881 VGND.t1506 125.368
R17409 VGND.n177 VGND.t1218 125.031
R17410 VGND.n8 VGND.t1547 124.46
R17411 VGND.n4949 VGND.t1449 124.46
R17412 VGND.n2798 VGND.t1016 124.46
R17413 VGND.n1515 VGND.t923 124.132
R17414 VGND.n81 VGND.t1038 124.124
R17415 VGND.n1620 VGND.t1235 124.088
R17416 VGND.n5452 VGND.t1491 124.088
R17417 VGND.n1640 VGND.t1517 124.079
R17418 VGND.n83 VGND.t999 124.07
R17419 VGND.n6852 VGND.t969 124.07
R17420 VGND.n9198 VGND.t870 123.546
R17421 VGND.n3442 VGND.t858 123.546
R17422 VGND.n7601 VGND.t1350 123.507
R17423 VGND.n3420 VGND.t1215 123.492
R17424 VGND.n93 VGND.t1192 123.492
R17425 VGND.n1691 VGND.t1582 123.492
R17426 VGND.n1628 VGND.t1375 123.406
R17427 VGND.n9164 VGND.t1274 122.907
R17428 VGND.n1399 VGND.t1466 122.907
R17429 VGND.n246 VGND.t912 122.907
R17430 VGND.n1482 VGND.t1013 122.907
R17431 VGND.n8900 VGND.t1389 122.892
R17432 VGND.n8265 VGND.t1323 122.63
R17433 VGND.n1619 VGND.t1236 121.987
R17434 VGND.n3487 VGND.t1571 121.956
R17435 VGND.n3487 VGND.t1572 121.956
R17436 VGND.n3485 VGND.t1032 121.956
R17437 VGND.n3485 VGND.t1031 121.956
R17438 VGND.n9101 VGND.t1275 121.956
R17439 VGND.n9165 VGND.t939 121.956
R17440 VGND.n2184 VGND.t1320 121.956
R17441 VGND.n2180 VGND.t1094 121.956
R17442 VGND.n2179 VGND.t1311 121.956
R17443 VGND.n2194 VGND.t1310 121.956
R17444 VGND.n2175 VGND.t1095 121.956
R17445 VGND.n2201 VGND.t888 121.956
R17446 VGND.n2213 VGND.t1433 121.956
R17447 VGND.n2171 VGND.t889 121.956
R17448 VGND.n2274 VGND.t1434 121.956
R17449 VGND.n2618 VGND.t1001 121.956
R17450 VGND.n2288 VGND.t1002 121.956
R17451 VGND.n2287 VGND.t1088 121.956
R17452 VGND.n2296 VGND.t1159 121.956
R17453 VGND.n2304 VGND.t1160 121.956
R17454 VGND.n2308 VGND.t1314 121.956
R17455 VGND.n2568 VGND.t1313 121.956
R17456 VGND.n2335 VGND.t1230 121.956
R17457 VGND.n2311 VGND.t1229 121.956
R17458 VGND.n2474 VGND.t1187 121.956
R17459 VGND.n2339 VGND.t1186 121.956
R17460 VGND.n2346 VGND.t957 121.956
R17461 VGND.n2343 VGND.t956 121.956
R17462 VGND.n2351 VGND.t1290 121.956
R17463 VGND.n2348 VGND.t1289 121.956
R17464 VGND.n2387 VGND.t975 121.956
R17465 VGND.n2406 VGND.t974 121.956
R17466 VGND.n9199 VGND.t1319 121.956
R17467 VGND.n15 VGND.t871 121.956
R17468 VGND.n10 VGND.t1548 121.956
R17469 VGND.n7 VGND.t1116 121.956
R17470 VGND.n7 VGND.t1115 121.956
R17471 VGND.n5136 VGND.t1568 121.956
R17472 VGND.n5134 VGND.t1567 121.956
R17473 VGND.n5498 VGND.t853 121.956
R17474 VGND.n5504 VGND.t852 121.956
R17475 VGND.n5540 VGND.t1034 121.956
R17476 VGND.n5560 VGND.t1035 121.956
R17477 VGND.n5497 VGND.t1242 121.956
R17478 VGND.n5564 VGND.t1241 121.956
R17479 VGND.n5594 VGND.t1420 121.956
R17480 VGND.n5586 VGND.t1419 121.956
R17481 VGND.n5635 VGND.t1537 121.956
R17482 VGND.n5470 VGND.t1538 121.956
R17483 VGND.n5679 VGND.t1579 121.956
R17484 VGND.n5698 VGND.t1580 121.956
R17485 VGND.n5469 VGND.t972 121.956
R17486 VGND.n5701 VGND.t971 121.956
R17487 VGND.n5755 VGND.t1444 121.956
R17488 VGND.n5735 VGND.t1443 121.956
R17489 VGND.n5127 VGND.t1047 121.956
R17490 VGND.n5799 VGND.t1046 121.956
R17491 VGND.n5154 VGND.t947 121.956
R17492 VGND.n5146 VGND.t948 121.956
R17493 VGND.n1857 VGND.t1248 121.956
R17494 VGND.n5970 VGND.t1247 121.956
R17495 VGND.n1860 VGND.t1384 121.956
R17496 VGND.n1859 VGND.t1383 121.956
R17497 VGND.n5111 VGND.t1408 121.956
R17498 VGND.n5926 VGND.t1407 121.956
R17499 VGND.n1800 VGND.t1357 121.956
R17500 VGND.n1808 VGND.t1356 121.956
R17501 VGND.n1801 VGND.t1178 121.956
R17502 VGND.n1804 VGND.t1177 121.956
R17503 VGND.n5223 VGND.t1221 121.956
R17504 VGND.n5225 VGND.t1222 121.956
R17505 VGND.n5225 VGND.t1438 121.956
R17506 VGND.n5223 VGND.t1437 121.956
R17507 VGND.n5228 VGND.t1077 121.956
R17508 VGND.n5231 VGND.t873 121.956
R17509 VGND.n5233 VGND.t874 121.956
R17510 VGND.n5233 VGND.t1078 121.956
R17511 VGND.n5236 VGND.t1353 121.956
R17512 VGND.n5236 VGND.t1354 121.956
R17513 VGND.n5234 VGND.t1543 121.956
R17514 VGND.n5234 VGND.t1542 121.956
R17515 VGND.n6668 VGND.t1213 121.956
R17516 VGND.n6656 VGND.t1212 121.956
R17517 VGND.n6656 VGND.t1532 121.956
R17518 VGND.n1631 VGND.t1533 121.956
R17519 VGND.n1627 VGND.t1196 121.956
R17520 VGND.n6689 VGND.t1520 121.956
R17521 VGND.n1621 VGND.t1521 121.956
R17522 VGND.n5363 VGND.t1456 121.956
R17523 VGND.n6706 VGND.t959 121.956
R17524 VGND.n5398 VGND.t1172 121.956
R17525 VGND.n5407 VGND.t1260 121.956
R17526 VGND.n5204 VGND.t1261 121.956
R17527 VGND.n5203 VGND.t936 121.956
R17528 VGND.n5419 VGND.t1004 121.956
R17529 VGND.n5200 VGND.t1005 121.956
R17530 VGND.n5428 VGND.t864 121.956
R17531 VGND.n5451 VGND.t1492 121.956
R17532 VGND.n1648 VGND.t883 121.956
R17533 VGND.n1644 VGND.t1518 121.956
R17534 VGND.n6612 VGND.t882 121.956
R17535 VGND.n1639 VGND.t951 121.956
R17536 VGND.n6619 VGND.t1044 121.956
R17537 VGND.n1638 VGND.t1043 121.956
R17538 VGND.n1739 VGND.t1345 121.956
R17539 VGND.n1732 VGND.t1344 121.956
R17540 VGND.n1710 VGND.t1405 121.956
R17541 VGND.n1716 VGND.t1404 121.956
R17542 VGND.n1713 VGND.t1479 121.956
R17543 VGND.n1713 VGND.t1480 121.956
R17544 VGND.n1711 VGND.t910 121.956
R17545 VGND.n1711 VGND.t909 121.956
R17546 VGND.n5047 VGND.t1426 121.956
R17547 VGND.n5045 VGND.t1425 121.956
R17548 VGND.n5062 VGND.t965 121.956
R17549 VGND.n4036 VGND.t966 121.956
R17550 VGND.n7150 VGND.t1112 121.956
R17551 VGND.n1346 VGND.t1113 121.956
R17552 VGND.n7105 VGND.t987 121.956
R17553 VGND.n1352 VGND.t986 121.956
R17554 VGND.n5088 VGND.t1410 121.956
R17555 VGND.n7003 VGND.t1411 121.956
R17556 VGND.n7067 VGND.t1526 121.956
R17557 VGND.n7006 VGND.t1527 121.956
R17558 VGND.n7011 VGND.t1166 121.956
R17559 VGND.n7010 VGND.t1165 121.956
R17560 VGND.n7014 VGND.t920 121.956
R17561 VGND.n7014 VGND.t921 121.956
R17562 VGND.n7012 VGND.t898 121.956
R17563 VGND.n7012 VGND.t897 121.956
R17564 VGND.n4851 VGND.t1463 121.956
R17565 VGND.n4089 VGND.t1464 121.956
R17566 VGND.n4087 VGND.t1515 121.956
R17567 VGND.n4911 VGND.t1514 121.956
R17568 VGND.n4082 VGND.t1255 121.956
R17569 VGND.n4919 VGND.t1254 121.956
R17570 VGND.n4982 VGND.t1450 121.956
R17571 VGND.n4950 VGND.t1074 121.956
R17572 VGND.n4984 VGND.t1075 121.956
R17573 VGND.n4768 VGND.t1068 121.956
R17574 VGND.n4768 VGND.t1069 121.956
R17575 VGND.n4767 VGND.t1041 121.956
R17576 VGND.n4767 VGND.t1040 121.956
R17577 VGND.n1408 VGND.t1399 121.956
R17578 VGND.n1422 VGND.t1398 121.956
R17579 VGND.n1411 VGND.t906 121.956
R17580 VGND.n1411 VGND.t907 121.956
R17581 VGND.n1409 VGND.t1124 121.956
R17582 VGND.n1409 VGND.t1123 121.956
R17583 VGND.n4589 VGND.t1181 121.956
R17584 VGND.n4568 VGND.t1180 121.956
R17585 VGND.n4565 VGND.t1340 121.956
R17586 VGND.n4630 VGND.t1339 121.956
R17587 VGND.n4552 VGND.t1097 121.956
R17588 VGND.n4652 VGND.t1098 121.956
R17589 VGND.n4173 VGND.t1502 121.956
R17590 VGND.n4547 VGND.t1503 121.956
R17591 VGND.n4477 VGND.t1028 121.956
R17592 VGND.n4515 VGND.t1029 121.956
R17593 VGND.n4451 VGND.t1293 121.956
R17594 VGND.n4450 VGND.t1292 121.956
R17595 VGND.n4434 VGND.t1363 121.956
R17596 VGND.n4433 VGND.t1362 121.956
R17597 VGND.n4218 VGND.t1145 121.956
R17598 VGND.n4424 VGND.t1144 121.956
R17599 VGND.n4307 VGND.t1207 121.956
R17600 VGND.n4294 VGND.t1206 121.956
R17601 VGND.n4236 VGND.t945 121.956
R17602 VGND.n4248 VGND.t944 121.956
R17603 VGND.n4239 VGND.t1210 121.956
R17604 VGND.n4240 VGND.t1209 121.956
R17605 VGND.n4666 VGND.t1393 121.956
R17606 VGND.n4166 VGND.t1392 121.956
R17607 VGND.n4162 VGND.t880 121.956
R17608 VGND.n4161 VGND.t879 121.956
R17609 VGND.n4150 VGND.t1326 121.956
R17610 VGND.n4117 VGND.t1325 121.956
R17611 VGND.n4100 VGND.t1057 121.956
R17612 VGND.n4100 VGND.t1058 121.956
R17613 VGND.n4099 VGND.t1252 121.956
R17614 VGND.n4099 VGND.t1251 121.956
R17615 VGND.n1393 VGND.t995 121.956
R17616 VGND.n1395 VGND.t996 121.956
R17617 VGND.n1398 VGND.t1467 121.956
R17618 VGND.n2963 VGND.t1071 121.956
R17619 VGND.n2899 VGND.t1072 121.956
R17620 VGND.n2904 VGND.t1122 121.956
R17621 VGND.n2924 VGND.t1121 121.956
R17622 VGND.n2909 VGND.t855 121.956
R17623 VGND.n2909 VGND.t856 121.956
R17624 VGND.n2908 VGND.t1570 121.956
R17625 VGND.n2908 VGND.t1569 121.956
R17626 VGND.n2758 VGND.t1296 121.956
R17627 VGND.n2772 VGND.t1295 121.956
R17628 VGND.n2808 VGND.t1017 121.956
R17629 VGND.n2801 VGND.t1286 121.956
R17630 VGND.n2817 VGND.t1287 121.956
R17631 VGND.n2836 VGND.t904 121.956
R17632 VGND.n2829 VGND.t903 121.956
R17633 VGND.n2751 VGND.t1284 121.956
R17634 VGND.n2849 VGND.t1283 121.956
R17635 VGND.n2866 VGND.t962 121.956
R17636 VGND.n2877 VGND.t963 121.956
R17637 VGND.n3222 VGND.t927 121.956
R17638 VGND.n3213 VGND.t926 121.956
R17639 VGND.n2658 VGND.t1190 121.956
R17640 VGND.n2656 VGND.t1189 121.956
R17641 VGND.n3310 VGND.t1555 121.956
R17642 VGND.n2652 VGND.t1486 121.956
R17643 VGND.n3305 VGND.t1053 121.956
R17644 VGND.n3322 VGND.t1052 121.956
R17645 VGND.n3320 VGND.t1565 121.956
R17646 VGND.n2123 VGND.t877 121.956
R17647 VGND.n2122 VGND.t1564 121.956
R17648 VGND.n2118 VGND.t876 121.956
R17649 VGND.n2121 VGND.t990 121.956
R17650 VGND.n2117 VGND.t1299 121.956
R17651 VGND.n2114 VGND.t989 121.956
R17652 VGND.n3421 VGND.t1298 121.956
R17653 VGND.n2113 VGND.t1216 121.956
R17654 VGND.n3443 VGND.t1529 121.956
R17655 VGND.n2106 VGND.t859 121.956
R17656 VGND.n2101 VGND.t1020 121.956
R17657 VGND.n3574 VGND.t1019 121.956
R17658 VGND.n3447 VGND.t1110 121.956
R17659 VGND.n2060 VGND.t1109 121.956
R17660 VGND.n2047 VGND.t1512 121.956
R17661 VGND.n2053 VGND.t1511 121.956
R17662 VGND.n2050 VGND.t1054 121.956
R17663 VGND.n2050 VGND.t1055 121.956
R17664 VGND.n2048 VGND.t1026 121.956
R17665 VGND.n2048 VGND.t1025 121.956
R17666 VGND.n2682 VGND.t1079 121.956
R17667 VGND.n2682 VGND.t1080 121.956
R17668 VGND.n2681 VGND.t1050 121.956
R17669 VGND.n2681 VGND.t1049 121.956
R17670 VGND.n9016 VGND.t1387 121.956
R17671 VGND.n8982 VGND.t1386 121.956
R17672 VGND.n3050 VGND.t1153 121.956
R17673 VGND.n3057 VGND.t1223 121.956
R17674 VGND.n3065 VGND.t1224 121.956
R17675 VGND.n3031 VGND.t1154 121.956
R17676 VGND.n3027 VGND.t1586 121.956
R17677 VGND.n3077 VGND.t1585 121.956
R17678 VGND.n3168 VGND.t1163 121.956
R17679 VGND.n3104 VGND.t1162 121.956
R17680 VGND.n3189 VGND.t1471 121.956
R17681 VGND.n2718 VGND.t1472 121.956
R17682 VGND.n2694 VGND.t1331 121.956
R17683 VGND.n2672 VGND.t1332 121.956
R17684 VGND.n8967 VGND.t1337 121.956
R17685 VGND.n8959 VGND.t1336 121.956
R17686 VGND.n79 VGND.t1008 121.956
R17687 VGND.n8919 VGND.t1007 121.956
R17688 VGND.n8915 VGND.t1063 121.956
R17689 VGND.n8915 VGND.t1064 121.956
R17690 VGND.n98 VGND.t1104 121.956
R17691 VGND.n97 VGND.t1037 121.956
R17692 VGND.n8876 VGND.t1103 121.956
R17693 VGND.n96 VGND.t1193 121.956
R17694 VGND.n8888 VGND.t1157 121.956
R17695 VGND.n8891 VGND.t1156 121.956
R17696 VGND.n8902 VGND.t1390 121.956
R17697 VGND.n3636 VGND.t998 121.956
R17698 VGND.n3637 VGND.t1086 121.956
R17699 VGND.n3633 VGND.t1227 121.956
R17700 VGND.n3661 VGND.t1085 121.956
R17701 VGND.n3630 VGND.t1308 121.956
R17702 VGND.n3690 VGND.t1226 121.956
R17703 VGND.n3690 VGND.t1307 121.956
R17704 VGND.n3669 VGND.t984 121.956
R17705 VGND.n3675 VGND.t983 121.956
R17706 VGND.n3672 VGND.t1268 121.956
R17707 VGND.n3672 VGND.t1269 121.956
R17708 VGND.n3670 VGND.t1239 121.956
R17709 VGND.n3670 VGND.t1238 121.956
R17710 VGND.n239 VGND.t941 121.956
R17711 VGND.n244 VGND.t942 121.956
R17712 VGND.n254 VGND.t913 121.956
R17713 VGND.n8536 VGND.t1183 121.956
R17714 VGND.n8451 VGND.t1184 121.956
R17715 VGND.n8455 VGND.t1360 121.956
R17716 VGND.n8454 VGND.t1359 121.956
R17717 VGND.n8460 VGND.t891 121.956
R17718 VGND.n8461 VGND.t892 121.956
R17719 VGND.n8464 VGND.t1368 121.956
R17720 VGND.n8464 VGND.t1369 121.956
R17721 VGND.n8462 VGND.t1553 121.956
R17722 VGND.n8462 VGND.t1552 121.956
R17723 VGND.n192 VGND.t1175 121.956
R17724 VGND.n189 VGND.t977 121.956
R17725 VGND.n188 VGND.t1250 121.956
R17726 VGND.n183 VGND.t1249 121.956
R17727 VGND.n178 VGND.t1219 121.956
R17728 VGND.n8749 VGND.t1458 121.956
R17729 VGND.n8740 VGND.t1459 121.956
R17730 VGND.n171 VGND.t885 121.956
R17731 VGND.n8756 VGND.t886 121.956
R17732 VGND.n163 VGND.t1130 121.956
R17733 VGND.n162 VGND.t1129 121.956
R17734 VGND.n3956 VGND.t1489 121.956
R17735 VGND.n3881 VGND.t1488 121.956
R17736 VGND.n1863 VGND.t1083 121.956
R17737 VGND.n3848 VGND.t1082 121.956
R17738 VGND.n3795 VGND.t1316 121.956
R17739 VGND.n3773 VGND.t1317 121.956
R17740 VGND.n3780 VGND.t1493 121.956
R17741 VGND.n3780 VGND.t1494 121.956
R17742 VGND.n3779 VGND.t933 121.956
R17743 VGND.n3779 VGND.t932 121.956
R17744 VGND.n8702 VGND.t1371 121.956
R17745 VGND.n206 VGND.t978 121.956
R17746 VGND.n215 VGND.t1372 121.956
R17747 VGND.n8619 VGND.t1523 121.956
R17748 VGND.n225 VGND.t1524 121.956
R17749 VGND.n226 VGND.t918 121.956
R17750 VGND.n8597 VGND.t919 121.956
R17751 VGND.n235 VGND.t980 121.956
R17752 VGND.n234 VGND.t981 121.956
R17753 VGND.n8355 VGND.t1010 121.956
R17754 VGND.n8355 VGND.t1011 121.956
R17755 VGND.n8353 VGND.t1198 121.956
R17756 VGND.n8353 VGND.t1197 121.956
R17757 VGND.n8381 VGND.t915 121.956
R17758 VGND.n8383 VGND.t916 121.956
R17759 VGND.n1898 VGND.t1452 121.956
R17760 VGND.n1901 VGND.t1453 121.956
R17761 VGND.n1881 VGND.t901 121.956
R17762 VGND.n1889 VGND.t900 121.956
R17763 VGND.n1885 VGND.t1141 121.956
R17764 VGND.n1885 VGND.t1142 121.956
R17765 VGND.n1884 VGND.t1342 121.956
R17766 VGND.n1884 VGND.t1341 121.956
R17767 VGND.n7906 VGND.t1118 121.956
R17768 VGND.n8068 VGND.t1119 121.956
R17769 VGND.n492 VGND.t1576 121.956
R17770 VGND.n496 VGND.t1577 121.956
R17771 VGND.n8036 VGND.t1091 121.956
R17772 VGND.n7948 VGND.t1092 121.956
R17773 VGND.n7901 VGND.t1366 121.956
R17774 VGND.n7893 VGND.t1365 121.956
R17775 VGND.n501 VGND.t1305 121.956
R17776 VGND.n7854 VGND.t1280 121.956
R17777 VGND.n502 VGND.t1281 121.956
R17778 VGND.n7854 VGND.t1304 121.956
R17779 VGND.n503 VGND.t954 121.956
R17780 VGND.n7845 VGND.t953 121.956
R17781 VGND.n505 VGND.t1541 121.956
R17782 VGND.n535 VGND.t1508 121.956
R17783 VGND.n537 VGND.t1509 121.956
R17784 VGND.n529 VGND.t1540 121.956
R17785 VGND.n523 VGND.t861 121.956
R17786 VGND.n528 VGND.t862 121.956
R17787 VGND.n528 VGND.t1061 121.956
R17788 VGND.n519 VGND.t1060 121.956
R17789 VGND.n516 VGND.t1127 121.956
R17790 VGND.n509 VGND.t1126 121.956
R17791 VGND.n1926 VGND.t1233 121.956
R17792 VGND.n1921 VGND.t1381 121.956
R17793 VGND.n1925 VGND.t1232 121.956
R17794 VGND.n433 VGND.t1422 121.956
R17795 VGND.n332 VGND.t1133 121.956
R17796 VGND.n401 VGND.t1132 121.956
R17797 VGND.n336 VGND.t1423 121.956
R17798 VGND.n342 VGND.t1200 121.956
R17799 VGND.n343 VGND.t1201 121.956
R17800 VGND.n350 VGND.t1263 121.956
R17801 VGND.n350 VGND.t1264 121.956
R17802 VGND.n349 VGND.t1436 121.956
R17803 VGND.n349 VGND.t1435 121.956
R17804 VGND.n8281 VGND.t1482 121.956
R17805 VGND.n441 VGND.t1483 121.956
R17806 VGND.n446 VGND.t1322 121.956
R17807 VGND.n8157 VGND.t1106 121.956
R17808 VGND.n8159 VGND.t1107 121.956
R17809 VGND.n8220 VGND.t1258 121.956
R17810 VGND.n455 VGND.t1257 121.956
R17811 VGND.n607 VGND.t1169 121.956
R17812 VGND.n673 VGND.t1168 121.956
R17813 VGND.n7608 VGND.t1022 121.956
R17814 VGND.n600 VGND.t1023 121.956
R17815 VGND.n7604 VGND.t1351 121.956
R17816 VGND.n7598 VGND.t1348 121.956
R17817 VGND.n7670 VGND.t1441 121.956
R17818 VGND.n7678 VGND.t1347 121.956
R17819 VGND.n7586 VGND.t1440 121.956
R17820 VGND.n686 VGND.t930 121.956
R17821 VGND.n7534 VGND.t929 121.956
R17822 VGND.n704 VGND.t1203 121.956
R17823 VGND.n690 VGND.t1204 121.956
R17824 VGND.n693 VGND.t1395 121.956
R17825 VGND.n693 VGND.t1396 121.956
R17826 VGND.n692 VGND.t1545 121.956
R17827 VGND.n692 VGND.t1544 121.956
R17828 VGND.n448 VGND.t1428 121.956
R17829 VGND.n448 VGND.t1427 121.956
R17830 VGND.n1191 VGND.t1478 121.956
R17831 VGND.n1215 VGND.t1477 121.956
R17832 VGND.n888 VGND.t1277 121.956
R17833 VGND.n904 VGND.t1278 121.956
R17834 VGND.n908 VGND.t867 121.956
R17835 VGND.n914 VGND.t868 121.956
R17836 VGND.n930 VGND.t1468 121.956
R17837 VGND.n930 VGND.t1469 121.956
R17838 VGND.n929 VGND.t1417 121.956
R17839 VGND.n929 VGND.t1416 121.956
R17840 VGND.n7435 VGND.t1100 121.956
R17841 VGND.n804 VGND.t1101 121.956
R17842 VGND.n805 VGND.t1561 121.956
R17843 VGND.n7387 VGND.t1562 121.956
R17844 VGND.n7383 VGND.t1301 121.956
R17845 VGND.n809 VGND.t1302 121.956
R17846 VGND.n7338 VGND.t895 121.956
R17847 VGND.n816 VGND.t894 121.956
R17848 VGND.n1075 VGND.t1066 121.956
R17849 VGND.n1097 VGND.t1067 121.956
R17850 VGND.n1007 VGND.t1245 121.956
R17851 VGND.n1103 VGND.t1244 121.956
R17852 VGND.n1112 VGND.t1150 121.956
R17853 VGND.n1119 VGND.t1550 121.956
R17854 VGND.n1146 VGND.t1151 121.956
R17855 VGND.n1149 VGND.t1551 121.956
R17856 VGND.n7458 VGND.t1267 121.956
R17857 VGND.n7464 VGND.t1266 121.956
R17858 VGND.n7461 VGND.t849 121.956
R17859 VGND.n7461 VGND.t850 121.956
R17860 VGND.n7459 VGND.t1535 121.956
R17861 VGND.n7459 VGND.t1534 121.956
R17862 VGND.n6863 VGND.t1377 121.956
R17863 VGND.n1586 VGND.t1378 121.956
R17864 VGND.n6934 VGND.t1414 121.956
R17865 VGND.n6910 VGND.t1413 121.956
R17866 VGND.n1478 VGND.t1474 121.956
R17867 VGND.n1480 VGND.t1475 121.956
R17868 VGND.n1484 VGND.t1014 121.956
R17869 VGND.n1486 VGND.t924 121.956
R17870 VGND.n1518 VGND.t1430 121.956
R17871 VGND.n1489 VGND.t1431 121.956
R17872 VGND.n1492 VGND.t1135 121.956
R17873 VGND.n1492 VGND.t1136 121.956
R17874 VGND.n1490 VGND.t1334 121.956
R17875 VGND.n1490 VGND.t1333 121.956
R17876 VGND.n6820 VGND.t1447 121.956
R17877 VGND.n6360 VGND.t1446 121.956
R17878 VGND.n6828 VGND.t968 121.956
R17879 VGND.n1588 VGND.t1148 121.956
R17880 VGND.n1588 VGND.t1147 121.956
R17881 VGND.n6359 VGND.t1500 121.956
R17882 VGND.n6356 VGND.t1499 121.956
R17883 VGND.n6353 VGND.t993 121.956
R17884 VGND.n6389 VGND.t992 121.956
R17885 VGND.n6258 VGND.t1138 121.956
R17886 VGND.n6261 VGND.t1139 121.956
R17887 VGND.n6301 VGND.t1497 121.956
R17888 VGND.n6257 VGND.t1496 121.956
R17889 VGND.n6250 VGND.t1583 121.956
R17890 VGND.n6235 VGND.t1559 121.956
R17891 VGND.n6226 VGND.t1558 121.956
R17892 VGND.n6119 VGND.t1271 121.956
R17893 VGND.n6119 VGND.t1272 121.956
R17894 VGND.n6117 VGND.t1461 121.956
R17895 VGND.n6117 VGND.t1460 121.956
R17896 VGND.n9120 VGND.t1401 121.956
R17897 VGND.n9120 VGND.t1402 121.956
R17898 VGND.n9119 VGND.t1573 121.956
R17899 VGND.n9119 VGND.t1574 121.956
R17900 VGND.n910 VGND.t2844 121.698
R17901 VGND.n23 VGND.t2606 121.698
R17902 VGND.n2405 VGND.n2404 121.002
R17903 VGND.n1337 VGND.n1336 119.064
R17904 VGND.n7158 VGND.n7157 118.763
R17905 VGND.n4781 VGND.n4780 118.1
R17906 VGND.n4381 VGND.n4380 118.1
R17907 VGND.n4643 VGND.n4642 118.1
R17908 VGND.n3274 VGND.n3273 118.1
R17909 VGND.n8947 VGND.n8946 118.1
R17910 VGND.n8396 VGND.n8395 118.1
R17911 VGND.n1978 VGND.n1977 118.1
R17912 VGND.n1232 VGND.n1231 118.1
R17913 VGND.n6143 VGND.n6142 118.1
R17914 VGND.n6143 VGND.n6141 118.1
R17915 VGND.t967 VGND.t2542 118.008
R17916 VGND VGND.t312 118.008
R17917 VGND.t671 VGND.t2903 118.008
R17918 VGND.t2391 VGND.t356 118.008
R17919 VGND.t2667 VGND.t1765 118.008
R17920 VGND.t1635 VGND.t1820 118.008
R17921 VGND.t2464 VGND.t794 118.008
R17922 VGND.t3144 VGND.t528 118.008
R17923 VGND.n2445 VGND.n2347 117.49
R17924 VGND.n4247 VGND.n4246 117.49
R17925 VGND.n8981 VGND.n8980 117.49
R17926 VGND.n6331 VGND.n6330 117.49
R17927 VGND.n6579 VGND.n6578 116.754
R17928 VGND.n2710 VGND.n2709 116.754
R17929 VGND.n8943 VGND.n8942 116.754
R17930 VGND.n8773 VGND.n8772 116.754
R17931 VGND.n384 VGND.n383 116.754
R17932 VGND.n8276 VGND.n8275 116.754
R17933 VGND.n1153 VGND.n1152 116.754
R17934 VGND.n9150 VGND.n9102 116.754
R17935 VGND.n7644 VGND.n7643 116.338
R17936 VGND.n4627 VGND.n4626 116.219
R17937 VGND.n482 VGND.n481 116.219
R17938 VGND.n1015 VGND.n1014 116.219
R17939 VGND.n1585 VGND.n1583 116.219
R17940 VGND.n6831 VGND.n6830 116.219
R17941 VGND.n5903 VGND.t91 116.115
R17942 VGND.n1760 VGND.t199 116.115
R17943 VGND.n2820 VGND.t2267 116.115
R17944 VGND.n3247 VGND.t2194 116.115
R17945 VGND.n3682 VGND.t79 116.115
R17946 VGND.n4097 VGND.t472 116.115
R17947 VGND.n2896 VGND.t2398 116.115
R17948 VGND.n173 VGND.t2224 116.115
R17949 VGND.n3268 VGND.n3267 115.561
R17950 VGND.n2827 VGND.n2826 115.525
R17951 VGND.n1351 VGND.n1350 115.466
R17952 VGND.n7200 VGND.n7199 115.466
R17953 VGND.n4019 VGND.n3996 115.466
R17954 VGND.n5034 VGND.n5033 115.466
R17955 VGND.n5038 VGND.n5037 115.466
R17956 VGND.n5030 VGND.n5029 115.466
R17957 VGND.n5026 VGND.n4041 115.466
R17958 VGND.n4528 VGND.n4526 115.466
R17959 VGND.n8165 VGND.n8164 115.466
R17960 VGND.n3509 VGND.t1592 115.118
R17961 VGND.n4034 VGND.t2298 115.118
R17962 VGND.n7172 VGND.n1334 114.713
R17963 VGND.n4014 VGND.n4013 114.713
R17964 VGND VGND.n5075 114.713
R17965 VGND.n4215 VGND.n4214 114.713
R17966 VGND.n7875 VGND.n7874 114.713
R17967 VGND.n647 VGND.n646 114.713
R17968 VGND.n7955 VGND.n7954 114.409
R17969 VGND.n7953 VGND.n7952 114.409
R17970 VGND.n615 VGND.n614 114.409
R17971 VGND.n617 VGND.n616 114.409
R17972 VGND.n1242 VGND.n1241 114.409
R17973 VGND.n6347 VGND.n6346 114.409
R17974 VGND.n5080 VGND.t2324 113.677
R17975 VGND.n3505 VGND.t1590 113.677
R17976 VGND.n5112 VGND.t89 113.677
R17977 VGND.n2825 VGND.t2269 113.677
R17978 VGND.n3234 VGND.t2196 113.677
R17979 VGND.n3665 VGND.t77 113.677
R17980 VGND.n172 VGND.t2226 113.677
R17981 VGND.n1154 VGND.t2965 113.677
R17982 VGND.n7483 VGND.t577 113.654
R17983 VGND.n8000 VGND.n7999 113.398
R17984 VGND.n612 VGND.n611 113.398
R17985 VGND.n637 VGND.n636 113.398
R17986 VGND.n1160 VGND.n1159 113.398
R17987 VGND.n1224 VGND.n1223 113.398
R17988 VGND.n1058 VGND.n1057 113.398
R17989 VGND.n6345 VGND.n6344 113.398
R17990 VGND.n6417 VGND.n6416 113.398
R17991 VGND.n1946 VGND.n1943 113.207
R17992 VGND.n7584 VGND.n685 113.207
R17993 VGND.n2464 VGND.n2463 113.04
R17994 VGND.n1647 VGND.n1645 113.04
R17995 VGND.n4039 VGND.n4038 113.04
R17996 VGND.n2734 VGND.n2733 113.04
R17997 VGND.n8590 VGND.n8589 113.04
R17998 VGND.n710 VGND.n709 113.04
R17999 VGND.n907 VGND.n905 113.04
R18000 VGND.n7966 VGND.n7965 112.981
R18001 VGND.n7964 VGND.n7963 112.981
R18002 VGND.n651 VGND.n608 112.981
R18003 VGND.n610 VGND.n609 112.981
R18004 VGND.n1163 VGND.n1162 112.981
R18005 VGND.n1048 VGND.n1047 112.981
R18006 VGND.n6343 VGND.n6342 112.981
R18007 VGND.n7479 VGND.t575 112.975
R18008 VGND.n2664 VGND.t2396 112.698
R18009 VGND.n3495 VGND.n3494 112.579
R18010 VGND.n3495 VGND.n3493 112.579
R18011 VGND.n5668 VGND.n5667 112.579
R18012 VGND.n5577 VGND.n5576 112.579
R18013 VGND.n4778 VGND.n4777 112.579
R18014 VGND.n3787 VGND.n3786 112.579
R18015 VGND.n219 VGND.n218 112.579
R18016 VGND.n925 VGND.n924 112.579
R18017 VGND.n6127 VGND.n6126 112.579
R18018 VGND.n6127 VGND.n6125 112.579
R18019 VGND.n6454 VGND.n6339 112.579
R18020 VGND.n9110 VGND.n9109 112.579
R18021 VGND.n9117 VGND.n9116 112.579
R18022 VGND.n6861 VGND.n1587 112.406
R18023 VGND.n1053 VGND.n1052 112.254
R18024 VGND.n4106 VGND.t476 112.243
R18025 VGND.n7957 VGND.n7956 112.192
R18026 VGND.n8011 VGND.n8010 112.192
R18027 VGND.n633 VGND.n632 112.192
R18028 VGND.n627 VGND.n626 112.192
R18029 VGND.n1228 VGND.n1227 112.192
R18030 VGND.n1236 VGND.n1235 112.192
R18031 VGND.n1012 VGND.n1011 112.192
R18032 VGND.n1036 VGND.n1013 112.192
R18033 VGND.n6413 VGND.n6412 112.192
R18034 VGND.n6028 VGND.n6027 111.957
R18035 VGND.n7844 VGND.n7841 111.701
R18036 VGND.n1903 VGND.n1902 111.606
R18037 VGND.n3501 VGND.n3500 111.118
R18038 VGND.n3501 VGND.n3499 111.118
R18039 VGND.n2310 VGND.n2309 111.118
R18040 VGND.n5673 VGND.n5672 111.118
R18041 VGND.n5582 VGND.n5581 111.118
R18042 VGND.n4774 VGND.n4773 111.118
R18043 VGND.n1406 VGND.n1405 111.118
R18044 VGND.n4441 VGND.n4440 111.118
R18045 VGND.n3685 VGND.n3684 111.118
R18046 VGND.n3775 VGND.n3774 111.118
R18047 VGND.n8774 VGND.n8771 111.118
R18048 VGND.n8370 VGND.n8351 111.118
R18049 VGND.n923 VGND.n922 111.118
R18050 VGND.n6133 VGND.n6132 111.118
R18051 VGND.n6133 VGND.n6131 111.118
R18052 VGND.n9129 VGND.n9113 111.118
R18053 VGND.n2565 VGND.n2564 111.026
R18054 VGND.n5388 VGND.n5387 111.026
R18055 VGND.n1769 VGND.n1768 111.026
R18056 VGND.n7048 VGND.n7047 111.026
R18057 VGND.n4086 VGND.n4083 111.026
R18058 VGND.n4861 VGND.n4860 111.026
R18059 VGND.n4121 VGND.n4120 111.026
R18060 VGND.n4392 VGND.n4222 111.026
R18061 VGND.n4604 VGND.n4603 111.026
R18062 VGND.n2946 VGND.n2945 111.026
R18063 VGND.n3098 VGND.n3097 111.026
R18064 VGND.n8506 VGND.n8505 111.026
R18065 VGND.n217 VGND.n216 111.026
R18066 VGND.n7947 VGND.n7944 111.026
R18067 VGND.n7883 VGND.n7882 111.026
R18068 VGND.n7607 VGND.n7606 111.026
R18069 VGND.n8239 VGND.n8238 111.026
R18070 VGND.n957 VGND.n915 111.026
R18071 VGND.n7373 VGND.n7372 111.026
R18072 VGND.n6904 VGND.n6903 111.026
R18073 VGND.n6366 VGND.n6365 111.026
R18074 VGND.n6437 VGND.n6436 111.026
R18075 VGND.n8897 VGND.t2779 110.934
R18076 VGND.n5256 VGND.t1928 110.934
R18077 VGND.n5197 VGND.t1869 110.934
R18078 VGND.n1630 VGND.t3134 110.934
R18079 VGND.n2041 VGND.t2619 110.934
R18080 VGND.n1268 VGND.t2962 110.934
R18081 VGND.n3991 VGND.n3990 110.719
R18082 VGND.n3992 VGND.t34 110.588
R18083 VGND.n2901 VGND.t292 110.588
R18084 VGND.n8484 VGND.t3197 110.588
R18085 VGND.n1222 VGND.t454 110.588
R18086 VGND.n810 VGND.t2356 110.588
R18087 VGND.n2354 VGND.t2009 110.588
R18088 VGND.n1260 VGND.t1724 110.588
R18089 VGND.n1727 VGND.n1726 110.46
R18090 VGND.n7475 VGND.n7474 110.46
R18091 VGND.n7968 VGND.n7967 110.4
R18092 VGND.n1246 VGND.n1245 110.224
R18093 VGND.n1081 VGND.n1080 110.224
R18094 VGND.n1074 VGND.n1073 110.224
R18095 VGND.n6399 VGND.n6398 110.224
R18096 VGND.n8370 VGND.t2920 110.01
R18097 VGND.n1151 VGND.n1150 109.849
R18098 VGND.n8346 VGND.t487 109.681
R18099 VGND.n7142 VGND.n7141 109.653
R18100 VGND.t647 VGND.t2956 109.579
R18101 VGND.t210 VGND.t2248 109.579
R18102 VGND.t772 VGND.t2257 109.579
R18103 VGND VGND.t2201 109.579
R18104 VGND.t1821 VGND.t2819 109.579
R18105 VGND VGND.t2101 109.579
R18106 VGND.t2845 VGND.t3041 109.579
R18107 VGND.t2379 VGND.t2948 109.579
R18108 VGND.t2002 VGND.t1773 109.579
R18109 VGND.t3083 VGND.t2945 109.579
R18110 VGND.t548 VGND.t1081 109.579
R18111 VGND VGND.t540 109.579
R18112 VGND.n5076 VGND.n5074 109.567
R18113 VGND.n3952 VGND.n3884 109.567
R18114 VGND.n1329 VGND.t3094 109.523
R18115 VGND.n2338 VGND.t446 109.35
R18116 VGND.n8053 VGND.n486 109.3
R18117 VGND.n7960 VGND.n7959 108.957
R18118 VGND.n5226 VGND.t1930 108.945
R18119 VGND.n5444 VGND.t1865 108.945
R18120 VGND.n6677 VGND.t3132 108.945
R18121 VGND.n1770 VGND.t201 108.945
R18122 VGND.n2067 VGND.t2621 108.945
R18123 VGND.n86 VGND.t2775 108.945
R18124 VGND.n1043 VGND.n1040 108.629
R18125 VGND.n1213 VGND.n1212 108.629
R18126 VGND.n6426 VGND.n6425 108.629
R18127 VGND.n1332 VGND.t2202 108.505
R18128 VGND.n2466 VGND.n2465 108.312
R18129 VGND.n2552 VGND.n2551 108.312
R18130 VGND.n1722 VGND.n1707 108.312
R18131 VGND.n1421 VGND.n1419 108.312
R18132 VGND.n2059 VGND.n2044 108.312
R18133 VGND.n3681 VGND.n3666 108.312
R18134 VGND.n8363 VGND.n8362 108.312
R18135 VGND.n8344 VGND.n8343 108.312
R18136 VGND.n7470 VGND.n7455 108.312
R18137 VGND.n3509 VGND.t735 108.153
R18138 VGND.n5726 VGND.t40 108.153
R18139 VGND.n5529 VGND.t2358 108.153
R18140 VGND.n1861 VGND.t1700 108.153
R18141 VGND.n1824 VGND.t688 108.153
R18142 VGND.n6898 VGND.t2864 108.153
R18143 VGND.n2357 VGND.t103 108.151
R18144 VGND.n5130 VGND.t3026 108.151
R18145 VGND.n5115 VGND.t2951 108.151
R18146 VGND.n2907 VGND.t3170 108.151
R18147 VGND.n2680 VGND.t2653 108.151
R18148 VGND.n9105 VGND.t529 108.151
R18149 VGND.n348 VGND.t2729 108.151
R18150 VGND.n1339 VGND.n1338 108.016
R18151 VGND.n4458 VGND.n4457 108.016
R18152 VGND.n485 VGND.n484 108.016
R18153 VGND.n656 VGND.n655 108.008
R18154 VGND.n1207 VGND.n1206 108.008
R18155 VGND.n1062 VGND.n1061 108.008
R18156 VGND.n6439 VGND.n6438 108.008
R18157 VGND.n6407 VGND.n6406 108.008
R18158 VGND.n2418 VGND.t136 107.82
R18159 VGND.n2902 VGND.t147 107.82
R18160 VGND.n8457 VGND.t145 107.82
R18161 VGND.n8349 VGND.t149 107.82
R18162 VGND.n8347 VGND.t151 107.82
R18163 VGND.n920 VGND.t138 107.82
R18164 VGND.n1161 VGND.t2994 107.82
R18165 VGND.n1155 VGND.t2824 107.82
R18166 VGND.n7355 VGND.t2565 107.82
R18167 VGND.n3995 VGND.t2571 107.784
R18168 VGND.n3777 VGND.n3776 107.731
R18169 VGND.n8255 VGND.t21 107.719
R18170 VGND.n7837 VGND.n7836 107.627
R18171 VGND.n6646 VGND.n6645 107.605
R18172 VGND.n4897 VGND.n4896 107.605
R18173 VGND.n4680 VGND.n4679 107.605
R18174 VGND.n453 VGND.n452 107.605
R18175 VGND.n1042 VGND.n1041 107.605
R18176 VGND.n7483 VGND.n7453 107.54
R18177 VGND.n6378 VGND.n6377 107.38
R18178 VGND.n3523 VGND.n3522 107.24
R18179 VGND.n2412 VGND.n2356 107.24
R18180 VGND.n2353 VGND.n2352 107.24
R18181 VGND.n2338 VGND.n2337 107.24
R18182 VGND.n5132 VGND.n5131 107.24
R18183 VGND.n5129 VGND.n5128 107.24
R18184 VGND.n5731 VGND.n5730 107.24
R18185 VGND.n5534 VGND.n5533 107.24
R18186 VGND.n5896 VGND.n5113 107.24
R18187 VGND.n5109 VGND.n5108 107.24
R18188 VGND.n1839 VGND.n1838 107.24
R18189 VGND.n1819 VGND.n1818 107.24
R18190 VGND.n6653 VGND.n1632 107.24
R18191 VGND.n6637 VGND.n1633 107.24
R18192 VGND.n1727 VGND.n1725 107.24
R18193 VGND.n6023 VGND.n6022 107.24
R18194 VGND.n7158 VGND.n1342 107.24
R18195 VGND.n3995 VGND.n3994 107.24
R18196 VGND.n3989 VGND.n3988 107.24
R18197 VGND.n4947 VGND.n4076 107.24
R18198 VGND.n4946 VGND.n4079 107.24
R18199 VGND.n4909 VGND.n4908 107.24
R18200 VGND.n4873 VGND.n4872 107.24
R18201 VGND.n1404 VGND.n1403 107.24
R18202 VGND.n4106 VGND.n4105 107.24
R18203 VGND.n4113 VGND.n4112 107.24
R18204 VGND.n4403 VGND.n4402 107.24
R18205 VGND.n4409 VGND.n4408 107.24
R18206 VGND.n4414 VGND.n4413 107.24
R18207 VGND.n1391 VGND.n1390 107.24
R18208 VGND.n2906 VGND.n2905 107.24
R18209 VGND.n2918 VGND.n2917 107.24
R18210 VGND.n2860 VGND.n2859 107.24
R18211 VGND.n3224 VGND.n3223 107.24
R18212 VGND.n2677 VGND.n2676 107.24
R18213 VGND.n2679 VGND.n2678 107.24
R18214 VGND.n8975 VGND.n8974 107.24
R18215 VGND.n8459 VGND.n8458 107.24
R18216 VGND.n3883 VGND.n3882 107.24
R18217 VGND.n3922 VGND.n3921 107.24
R18218 VGND.n8783 VGND.n159 107.24
R18219 VGND.n7950 VGND.n7949 107.24
R18220 VGND.n483 VGND.n480 107.24
R18221 VGND.n345 VGND.n344 107.24
R18222 VGND.n347 VGND.n346 107.24
R18223 VGND.n338 VGND.n337 107.24
R18224 VGND.n699 VGND.n698 107.24
R18225 VGND.n7644 VGND.n7642 107.24
R18226 VGND.n8143 VGND.n8142 107.24
R18227 VGND.n8271 VGND.n8270 107.24
R18228 VGND.n927 VGND.n926 107.24
R18229 VGND.n815 VGND.n814 107.24
R18230 VGND.n7475 VGND.n7473 107.24
R18231 VGND.n6213 VGND.n6212 107.24
R18232 VGND.n6264 VGND.n6263 107.24
R18233 VGND.n6349 VGND.n6348 107.24
R18234 VGND.n9104 VGND.n9103 107.24
R18235 VGND.n9115 VGND.n9114 107.24
R18236 VGND.n2459 VGND.n2341 107.162
R18237 VGND.n4656 VGND.n4551 107.162
R18238 VGND.n2043 VGND.n2042 107.162
R18239 VGND.n8633 VGND.n8632 107.162
R18240 VGND.n8386 VGND.n8382 107.162
R18241 VGND.n1891 VGND.n1890 107.162
R18242 VGND.n6450 VGND.n6448 107.162
R18243 VGND.n9108 VGND.n9107 107.162
R18244 VGND.n2671 VGND.n2670 107.028
R18245 VGND.n8958 VGND.n8957 107.028
R18246 VGND.n4288 VGND.n4287 106.465
R18247 VGND.n8573 VGND.n255 106.465
R18248 VGND.n8419 VGND.n8418 106.465
R18249 VGND.n7962 VGND.n7961 106.465
R18250 VGND.n813 VGND.n812 106.465
R18251 VGND.n1672 VGND.n1671 106.465
R18252 VGND.n1291 VGND.t456 106.055
R18253 VGND.n1330 VGND.t296 106.053
R18254 VGND.n4546 VGND.t2204 106.053
R18255 VGND.n3051 VGND.t2340 106.053
R18256 VGND.n946 VGND.t3090 106.053
R18257 VGND.n1341 VGND.n1340 105.975
R18258 VGND.n3859 VGND.n3858 105.749
R18259 VGND.n1945 VGND.n1944 105.749
R18260 VGND.n8258 VGND.n8257 104.96
R18261 VGND.n5210 VGND.n5205 104.743
R18262 VGND.n5060 VGND.n5059 104.719
R18263 VGND.n4620 VGND.n4619 104.719
R18264 VGND.n4563 VGND.n4557 104.719
R18265 VGND.n490 VGND.n489 104.719
R18266 VGND.n488 VGND.n487 104.719
R18267 VGND.n1066 VGND.n1065 104.719
R18268 VGND.n1023 VGND.n1017 104.719
R18269 VGND.n7318 VGND.n7317 104.719
R18270 VGND.n6880 VGND.n6879 104.719
R18271 VGND.n6887 VGND.n6886 104.719
R18272 VGND.n6839 VGND.n6838 104.719
R18273 VGND.n6845 VGND.n6844 104.719
R18274 VGND.n4040 VGND.t2228 104.609
R18275 VGND.n699 VGND.t3020 104.454
R18276 VGND.n3805 VGND.n3804 104.331
R18277 VGND.n1401 VGND.n1397 104.067
R18278 VGND.n17 VGND.t2031 103.968
R18279 VGND.n2586 VGND.t3168 103.966
R18280 VGND.n2242 VGND.t2275 103.966
R18281 VGND.n4026 VGND.t3203 103.966
R18282 VGND.n8466 VGND.t2448 103.966
R18283 VGND.n8357 VGND.t3162 103.966
R18284 VGND.n2434 VGND.n2433 103.942
R18285 VGND.n2556 VGND.n2555 103.942
R18286 VGND.n2292 VGND.n2290 103.942
R18287 VGND.n2227 VGND.n2226 103.942
R18288 VGND.n2183 VGND.n2181 103.942
R18289 VGND.n6546 VGND.n6545 103.942
R18290 VGND.n6044 VGND.n6043 103.942
R18291 VGND.n4792 VGND.n4790 103.942
R18292 VGND.n7019 VGND.n7018 103.942
R18293 VGND.n7008 VGND.n7007 103.942
R18294 VGND.n7127 VGND.n7126 103.942
R18295 VGND.n4927 VGND.n4926 103.942
R18296 VGND.n4898 VGND.n4895 103.942
R18297 VGND.n4715 VGND.n4712 103.942
R18298 VGND.n4165 VGND.n4164 103.942
R18299 VGND.n4714 VGND.n4713 103.942
R18300 VGND.n4676 VGND.n4675 103.942
R18301 VGND.n4258 VGND.n4257 103.942
R18302 VGND.n4280 VGND.n4279 103.942
R18303 VGND.n4393 VGND.n4221 103.942
R18304 VGND.n4422 VGND.n4421 103.942
R18305 VGND.n1439 VGND.n1438 103.942
R18306 VGND.n2844 VGND.n2843 103.942
R18307 VGND.n2936 VGND.n2935 103.942
R18308 VGND.n2654 VGND.n2653 103.942
R18309 VGND.n2840 VGND.n2839 103.942
R18310 VGND.n3212 VGND.n3211 103.942
R18311 VGND.n8918 VGND.n8917 103.942
R18312 VGND.n92 VGND.n90 103.942
R18313 VGND.n3130 VGND.n3129 103.942
R18314 VGND.n3108 VGND.n3107 103.942
R18315 VGND.n9041 VGND.n9040 103.942
R18316 VGND.n8992 VGND.n8991 103.942
R18317 VGND.n8473 VGND.n8470 103.942
R18318 VGND.n8496 VGND.n8495 103.942
R18319 VGND.n194 VGND.n193 103.942
R18320 VGND.n3847 VGND.n3846 103.942
R18321 VGND.n3931 VGND.n3930 103.942
R18322 VGND.n169 VGND.n168 103.942
R18323 VGND.n176 VGND.n174 103.942
R18324 VGND.n8624 VGND.n221 103.942
R18325 VGND.n8365 VGND.n8364 103.942
R18326 VGND.n7905 VGND.n7902 103.942
R18327 VGND.n8004 VGND.n8003 103.942
R18328 VGND.n8021 VGND.n8020 103.942
R18329 VGND.n522 VGND.n520 103.942
R18330 VGND.n7892 VGND.n7891 103.942
R18331 VGND.n7904 VGND.n7903 103.942
R18332 VGND.n340 VGND.n339 103.942
R18333 VGND.n7666 VGND.n7602 103.942
R18334 VGND.n657 VGND.n654 103.942
R18335 VGND.n8225 VGND.n8224 103.942
R18336 VGND.n8180 VGND.n8179 103.942
R18337 VGND.n8287 VGND.n8286 103.942
R18338 VGND.n947 VGND.n918 103.942
R18339 VGND.n1248 VGND.n1247 103.942
R18340 VGND.n1267 VGND.n1266 103.942
R18341 VGND.n7363 VGND.n7362 103.942
R18342 VGND.n1488 VGND.n1487 103.942
R18343 VGND.n1528 VGND.n1527 103.942
R18344 VGND.n6916 VGND.n6915 103.942
R18345 VGND.n6905 VGND.n6902 103.942
R18346 VGND.n6241 VGND.n1690 103.942
R18347 VGND.n6320 VGND.n6319 103.942
R18348 VGND.n6297 VGND.n6296 103.942
R18349 VGND.n6428 VGND.n6427 103.942
R18350 VGND.n6400 VGND.n6397 103.942
R18351 VGND.n9141 VGND.n9106 103.942
R18352 VGND.n4541 VGND.t1711 103.79
R18353 VGND.n4025 VGND.t2822 103.79
R18354 VGND.n1148 VGND.t634 103.79
R18355 VGND.n2479 VGND.t134 103.79
R18356 VGND.n7187 VGND.t116 103.79
R18357 VGND.n3056 VGND.t141 103.79
R18358 VGND.n4574 VGND.n4573 103.784
R18359 VGND.n5340 VGND.n5339 103.698
R18360 VGND.n4614 VGND.t3212 103.507
R18361 VGND.n866 VGND.t63 103.507
R18362 VGND.n5019 VGND.n5017 103.168
R18363 VGND.n4278 VGND.n4277 103.168
R18364 VGND.n4637 VGND.n4555 103.168
R18365 VGND.n2784 VGND.n2783 103.168
R18366 VGND.n3030 VGND.n3028 103.168
R18367 VGND.n9039 VGND.n9038 103.168
R18368 VGND.n6295 VGND.n6294 103.168
R18369 VGND.n4473 VGND.t1883 102.766
R18370 VGND.n7841 VGND.t185 101.43
R18371 VGND.n5054 VGND.t2601 101.156
R18372 VGND.n531 VGND.t2147 101.156
R18373 VGND.n498 VGND.t2976 101.156
R18374 VGND.n7579 VGND.t2188 101.156
R18375 VGND.t2842 VGND.t2773 101.15
R18376 VGND.n6630 VGND.t228 101.15
R18377 VGND.n5338 VGND.t2470 101.15
R18378 VGND.t1988 VGND.t2073 101.15
R18379 VGND.t2423 VGND.t248 101.15
R18380 VGND.t2405 VGND.t2696 101.15
R18381 VGND.t593 VGND.t1603 101.15
R18382 VGND.t131 VGND.t127 101.15
R18383 VGND.n6979 VGND.t2472 101.15
R18384 VGND.t2959 VGND.t1695 101.15
R18385 VGND.t2604 VGND.t1884 101.15
R18386 VGND.t3141 VGND.t2734 101.15
R18387 VGND.t2590 VGND.t3188 101.15
R18388 VGND.t2594 VGND.t728 101.15
R18389 VGND.t2586 VGND.t726 101.15
R18390 VGND.t2783 VGND.n222 101.15
R18391 VGND.t3246 VGND.t78 101.15
R18392 VGND.t2853 VGND.t2607 101.15
R18393 VGND.n3879 VGND.n3878 101.085
R18394 VGND.n7799 VGND.n7798 101.085
R18395 VGND.n7125 VGND.n7124 100.882
R18396 VGND.n4525 VGND.t112 100.653
R18397 VGND.n449 VGND.t3236 100.653
R18398 VGND.n5044 VGND.t11 100.653
R18399 VGND.n493 VGND.t725 100.21
R18400 VGND.n491 VGND.t2587 100.21
R18401 VGND.n6874 VGND.t507 100.21
R18402 VGND.n6851 VGND.t2539 100.21
R18403 VGND.n3868 VGND.n3867 100.162
R18404 VGND.n3945 VGND.n3944 100.162
R18405 VGND.n2347 VGND.t616 100.001
R18406 VGND.n2564 VGND.t2798 100.001
R18407 VGND.n5387 VGND.t2477 100.001
R18408 VGND.n1768 VGND.t239 100.001
R18409 VGND.n6578 VGND.t251 100.001
R18410 VGND.n7047 VGND.t2469 100.001
R18411 VGND.n4083 VGND.t221 100.001
R18412 VGND.n4860 VGND.t235 100.001
R18413 VGND.n4120 VGND.t243 100.001
R18414 VGND.n4246 VGND.t241 100.001
R18415 VGND.n4222 VGND.t253 100.001
R18416 VGND.n4603 VGND.t2491 100.001
R18417 VGND.n2945 VGND.t618 100.001
R18418 VGND.n2826 VGND.t2705 100.001
R18419 VGND.n3267 VGND.t2802 100.001
R18420 VGND.n2709 VGND.t2709 100.001
R18421 VGND.n3097 VGND.t632 100.001
R18422 VGND.n8942 VGND.t1687 100.001
R18423 VGND.n8980 VGND.t2808 100.001
R18424 VGND.n8505 VGND.t2711 100.001
R18425 VGND.n8772 VGND.t1677 100.001
R18426 VGND.n216 VGND.t2792 100.001
R18427 VGND.n7944 VGND.t2790 100.001
R18428 VGND.n7882 VGND.t628 100.001
R18429 VGND.n383 VGND.t2707 100.001
R18430 VGND.n7606 VGND.t1693 100.001
R18431 VGND.n8238 VGND.t2806 100.001
R18432 VGND.n8275 VGND.t614 100.001
R18433 VGND.n915 VGND.t2481 100.001
R18434 VGND.n1152 VGND.t2786 100.001
R18435 VGND.n7372 VGND.t255 100.001
R18436 VGND.n6903 VGND.t2479 100.001
R18437 VGND.n6365 VGND.t2493 100.001
R18438 VGND.n6330 VGND.t225 100.001
R18439 VGND.n6436 VGND.t245 100.001
R18440 VGND.n9102 VGND.t626 100.001
R18441 VGND.n1427 VGND.t1986 98.875
R18442 VGND.n4293 VGND.t132 98.875
R18443 VGND.n2796 VGND.t2467 98.875
R18444 VGND.n3046 VGND.t2639 98.875
R18445 VGND.n8340 VGND.t2989 98.875
R18446 VGND.n7968 VGND.t1780 98.875
R18447 VGND.n4553 VGND.t3006 98.0152
R18448 VGND.n4446 VGND.n4445 97.9005
R18449 VGND.n2879 VGND.t605 97.3829
R18450 VGND.n2489 VGND.n2488 96.9805
R18451 VGND.n230 VGND.n229 96.9805
R18452 VGND.n443 VGND.n442 96.9805
R18453 VGND.n2868 VGND.n2867 96.5538
R18454 VGND.n4301 VGND.t2840 96.4837
R18455 VGND.n3071 VGND.t2132 96.4837
R18456 VGND.n8580 VGND.t3116 96.4837
R18457 VGND.n7337 VGND.t2814 96.4837
R18458 VGND.n6286 VGND.t2077 96.4837
R18459 VGND.n6262 VGND.t1879 96.4837
R18460 VGND.n1865 VGND.t561 94.7488
R18461 VGND.n1347 VGND.t2037 93.2783
R18462 VGND.n3942 VGND.t1803 93.2783
R18463 VGND.n668 VGND.t2852 93.2783
R18464 VGND.n8085 VGND.t539 93.2779
R18465 VGND.t535 VGND.t41 92.7208
R18466 VGND.t807 VGND.t1256 92.7208
R18467 VGND.t2941 VGND.t72 92.7208
R18468 VGND.t526 VGND.t569 92.7208
R18469 VGND.n6045 VGND.n6042 92.5005
R18470 VGND.n6039 VGND.n6038 92.5005
R18471 VGND.n6564 VGND.n6563 92.5005
R18472 VGND.n1652 VGND.n1651 92.5005
R18473 VGND.n4883 VGND.n4882 92.5005
R18474 VGND.n4879 VGND.n4878 92.5005
R18475 VGND.n4460 VGND.n4459 92.5005
R18476 VGND.n4464 VGND.n4463 92.5005
R18477 VGND.n2706 VGND.n2705 92.5005
R18478 VGND.n2702 VGND.n2701 92.5005
R18479 VGND.n3887 VGND.n3886 92.5005
R18480 VGND.n1936 VGND.n1935 92.5005
R18481 VGND.n7565 VGND.n7564 92.5005
R18482 VGND.n7569 VGND.n7568 92.5005
R18483 VGND.n7141 VGND.t1657 87.1434
R18484 VGND.n1587 VGND.t703 86.3738
R18485 VGND.t2685 VGND.t2046 84.2917
R18486 VGND.t403 VGND.t813 84.2917
R18487 VGND.t1324 VGND.t1625 84.2917
R18488 VGND.t736 VGND.t457 84.2917
R18489 VGND.t2917 VGND.t1179 84.2917
R18490 VGND.t542 VGND.t1462 84.2917
R18491 VGND.t640 VGND 84.2917
R18492 VGND.t488 VGND.t638 84.2917
R18493 VGND.t2519 VGND.t556 84.2917
R18494 VGND.t2048 VGND 84.2917
R18495 VGND VGND.t447 84.2917
R18496 VGND.t152 VGND.t2943 84.2917
R18497 VGND.t2006 VGND 84.2917
R18498 VGND.t1649 VGND.t1128 84.2917
R18499 VGND.t611 VGND.t1312 84.2917
R18500 VGND.n5146 VGND.t3453 83.8949
R18501 VGND.n4218 VGND.t3474 83.8949
R18502 VGND.n2877 VGND.t3445 83.8949
R18503 VGND.n2672 VGND.t3323 83.8949
R18504 VGND.n8383 VGND.t3341 83.8949
R18505 VGND.n1398 VGND.t3309 83.8949
R18506 VGND.n8967 VGND.t3319 83.8949
R18507 VGND.n163 VGND.t3401 83.8949
R18508 VGND.n3990 VGND.t1873 83.8933
R18509 VGND.n6234 VGND.t3272 82.587
R18510 VGND.n1483 VGND.t3465 82.1249
R18511 VGND.n3886 VGND.t126 81.4291
R18512 VGND.n3878 VGND.t3071 81.4291
R18513 VGND.n7798 VGND.t433 81.4291
R18514 VGND.n6666 VGND.t3434 78.7329
R18515 VGND.n5202 VGND.t3277 78.7329
R18516 VGND.n2112 VGND.t3358 78.7329
R18517 VGND.n95 VGND.t3365 78.7329
R18518 VGND.n666 VGND.t3507 78.7329
R18519 VGND.n1204 VGND.t3269 78.7329
R18520 VGND.n6921 VGND.t3382 78.7329
R18521 VGND.n7063 VGND.t3389 78.7329
R18522 VGND.n4960 VGND.t3375 78.7329
R18523 VGND.n2806 VGND.t3449 78.7329
R18524 VGND.n8741 VGND.t3301 78.7329
R18525 VGND.n688 VGND.t3459 78.7329
R18526 VGND.n3630 VGND.t3330 76.4092
R18527 VGND.n7598 VGND.t3456 76.4092
R18528 VGND.n10 VGND.t3279 76.4077
R18529 VGND.n2101 VGND.t3448 76.4077
R18530 VGND.n5206 VGND.t3377 76.1558
R18531 VGND.n2300 VGND.n2299 76.0005
R18532 VGND.n5692 VGND.n5691 76.0005
R18533 VGND.n5655 VGND.n5654 76.0005
R18534 VGND.n5557 VGND.n5556 76.0005
R18535 VGND.n4561 VGND.n4560 76.0005
R18536 VGND.n4597 VGND.n4596 76.0005
R18537 VGND.n2952 VGND.n2951 76.0005
R18538 VGND.n2755 VGND.n2754 76.0005
R18539 VGND.n3302 VGND.n3301 76.0005
R18540 VGND.n3218 VGND.n3217 76.0005
R18541 VGND.n2724 VGND.n2723 76.0005
R18542 VGND.n8930 VGND.n8929 76.0005
R18543 VGND.n8512 VGND.n8511 76.0005
R18544 VGND.n251 VGND.n250 76.0005
R18545 VGND.n3965 VGND.n3964 76.0005
R18546 VGND.n8603 VGND.n8602 76.0005
R18547 VGND.n211 VGND.n210 76.0005
R18548 VGND.n513 VGND.n512 76.0005
R18549 VGND.n7863 VGND.n7862 76.0005
R18550 VGND.n7897 VGND.n7896 76.0005
R18551 VGND.n365 VGND.n364 76.0005
R18552 VGND.n8228 VGND.n8227 76.0005
R18553 VGND.n965 VGND.n964 76.0005
R18554 VGND.n1010 VGND.n1009 76.0005
R18555 VGND.n7420 VGND.n7419 76.0005
R18556 VGND.n6248 VGND.n6247 76.0005
R18557 VGND.n9158 VGND.n9157 76.0005
R18558 VGND.t2078 VGND.t415 75.8626
R18559 VGND.t642 VGND.t2897 75.8626
R18560 VGND VGND.t2322 75.8626
R18561 VGND.t2117 VGND.t2215 75.8626
R18562 VGND.t314 VGND.t310 75.8626
R18563 VGND.t45 VGND.t3153 75.8626
R18564 VGND.t2314 VGND.t3163 75.8626
R18565 VGND.t1678 VGND.t1802 75.8626
R18566 VGND.n1394 VGND.t3267 75.1361
R18567 VGND.n243 VGND.t3276 75.1361
R18568 VGND.n1479 VGND.t3359 75.1361
R18569 VGND.n1912 VGND.n1911 74.8382
R18570 VGND.n7400 VGND.n7399 74.8382
R18571 VGND.n792 VGND.n789 74.8382
R18572 VGND.n4956 VGND.t3420 74.3808
R18573 VGND.n7126 VGND.t306 74.2862
R18574 VGND.n3930 VGND.t2944 74.2862
R18575 VGND.n480 VGND.t485 74.2862
R18576 VGND.n654 VGND.t2503 74.2862
R18577 VGND.n8265 VGND.t3410 73.7549
R18578 VGND.n5240 VGND.t3506 73.7268
R18579 VGND.n526 VGND.t3307 73.7268
R18580 VGND.n2433 VGND.t630 72.8576
R18581 VGND.n2555 VGND.t2804 72.8576
R18582 VGND.n5339 VGND.t2471 72.8576
R18583 VGND.n6645 VGND.t2051 72.8576
R18584 VGND.n6545 VGND.t229 72.8576
R18585 VGND.n6043 VGND.t223 72.8576
R18586 VGND.n6027 VGND.t3124 72.8576
R18587 VGND.n7007 VGND.t2475 72.8576
R18588 VGND.n4926 VGND.t233 72.8576
R18589 VGND.n4896 VGND.t2140 72.8576
R18590 VGND.n4872 VGND.t257 72.8576
R18591 VGND.n4713 VGND.t247 72.8576
R18592 VGND.n4679 VGND.t1728 72.8576
R18593 VGND.n4257 VGND.t237 72.8576
R18594 VGND.n4402 VGND.t219 72.8576
R18595 VGND.n4573 VGND.t2473 72.8576
R18596 VGND.n2935 VGND.t2715 72.8576
R18597 VGND.n2839 VGND.t622 72.8576
R18598 VGND.n3211 VGND.t2788 72.8576
R18599 VGND.n2670 VGND.t2699 72.8576
R18600 VGND.n3107 VGND.t2713 72.8576
R18601 VGND.n8957 VGND.t1691 72.8576
R18602 VGND.n8991 VGND.t2782 72.8576
R18603 VGND.n8495 VGND.t2701 72.8576
R18604 VGND.n168 VGND.t1681 72.8576
R18605 VGND.n221 VGND.t2784 72.8576
R18606 VGND.n1902 VGND.t2171 72.8576
R18607 VGND.n8020 VGND.t2800 72.8576
R18608 VGND.n7891 VGND.t2717 72.8576
R18609 VGND.n339 VGND.t2703 72.8576
R18610 VGND.n7642 VGND.t1685 72.8576
R18611 VGND.n452 VGND.t2757 72.8576
R18612 VGND.n8224 VGND.t2796 72.8576
R18613 VGND.n8286 VGND.t624 72.8576
R18614 VGND.n918 VGND.t2485 72.8576
R18615 VGND.n1266 VGND.t2794 72.8576
R18616 VGND.n1041 VGND.t2145 72.8576
R18617 VGND.n7362 VGND.t231 72.8576
R18618 VGND.n6915 VGND.t2483 72.8576
R18619 VGND.n6319 VGND.t227 72.8576
R18620 VGND.n6427 VGND.t249 72.8576
R18621 VGND.n6377 VGND.t2489 72.8576
R18622 VGND.n9106 VGND.t620 72.8576
R18623 VGND.n8085 VGND.t483 70.4212
R18624 VGND.n1347 VGND.t304 70.4207
R18625 VGND.n3942 VGND.t2940 70.4207
R18626 VGND.n668 VGND.t2510 70.4207
R18627 VGND.n2347 VGND.t801 70.0005
R18628 VGND.n2564 VGND.t612 70.0005
R18629 VGND.n5387 VGND.t2651 70.0005
R18630 VGND.n1768 VGND.t3193 70.0005
R18631 VGND.n6578 VGND.t416 70.0005
R18632 VGND.n7047 VGND.t2933 70.0005
R18633 VGND.n4083 VGND.t3178 70.0005
R18634 VGND.n4860 VGND.t543 70.0005
R18635 VGND.n4120 VGND.t1626 70.0005
R18636 VGND.n4246 VGND.t3222 70.0005
R18637 VGND.n4222 VGND.t2980 70.0005
R18638 VGND.n4603 VGND.t2918 70.0005
R18639 VGND.n2945 VGND.t2084 70.0005
R18640 VGND.n2826 VGND.t2460 70.0005
R18641 VGND.n3267 VGND.t3182 70.0005
R18642 VGND.n2709 VGND.t2812 70.0005
R18643 VGND.n3097 VGND.t2749 70.0005
R18644 VGND.n8942 VGND.t2762 70.0005
R18645 VGND.n8980 VGND.t2516 70.0005
R18646 VGND.n8505 VGND.t1977 70.0005
R18647 VGND.n8772 VGND.t1652 70.0005
R18648 VGND.n216 VGND.t440 70.0005
R18649 VGND.n7944 VGND.t1715 70.0005
R18650 VGND.n7882 VGND.t1830 70.0005
R18651 VGND.n383 VGND.t2735 70.0005
R18652 VGND.n7606 VGND.t3010 70.0005
R18653 VGND.n8238 VGND.t1939 70.0005
R18654 VGND.n8275 VGND.t785 70.0005
R18655 VGND.n915 VGND.t2846 70.0005
R18656 VGND.n1152 VGND.t3014 70.0005
R18657 VGND.n7372 VGND.t164 70.0005
R18658 VGND.n6903 VGND.t515 70.0005
R18659 VGND.n6365 VGND.t551 70.0005
R18660 VGND.n6330 VGND.t217 70.0005
R18661 VGND.n6436 VGND.t402 70.0005
R18662 VGND.n9102 VGND.t2608 70.0005
R18663 VGND.n1622 VGND.t3286 68.7721
R18664 VGND.n4457 VGND.t379 68.3082
R18665 VGND.n1333 VGND.n1332 67.973
R18666 VGND.t2419 VGND.t2333 67.4335
R18667 VGND.t1498 VGND.t3154 67.4335
R18668 VGND.t514 VGND.t2997 67.4335
R18669 VGND.t776 VGND.t1716 67.4335
R18670 VGND.t3126 VGND.t2576 67.4335
R18671 VGND.t651 VGND.t3175 67.4335
R18672 VGND.t2142 VGND.t1658 67.4335
R18673 VGND.t2148 VGND.t16 67.4335
R18674 VGND.t2212 VGND.t12 67.4335
R18675 VGND.t2227 VGND.t14 67.4335
R18676 VGND.t1655 VGND.t1708 67.4335
R18677 VGND.t655 VGND.t1476 67.4335
R18678 VGND.t2521 VGND.t1747 67.4335
R18679 VGND.t3102 VGND.t3019 67.4335
R18680 VGND.t2908 VGND 67.4335
R18681 VGND.t2381 VGND.t1451 67.4335
R18682 VGND.t184 VGND 67.4335
R18683 VGND.t1829 VGND.t2738 67.4335
R18684 VGND.t1667 VGND.t2674 67.4335
R18685 VGND.t789 VGND.t1651 67.4335
R18686 VGND.t3035 VGND.t1908 67.4335
R18687 VGND.t2727 VGND.t3049 67.4335
R18688 VGND.t792 VGND.t157 67.4335
R18689 VGND.t3043 VGND.t1702 67.4335
R18690 VGND.t2240 VGND.t2681 67.4335
R18691 VGND.n7544 VGND.t3022 67.3107
R18692 VGND.n3867 VGND.t1689 67.1434
R18693 VGND.n3944 VGND.t1679 67.1434
R18694 VGND.n1935 VGND.t1683 67.1434
R18695 VGND.n7545 VGND.n7544 66.3713
R18696 VGND.n3838 VGND.t2013 65.3335
R18697 VGND.n3838 VGND.t3174 65.3335
R18698 VGND.n6223 VGND.t176 65.3335
R18699 VGND.n6223 VGND.t2662 65.3335
R18700 VGND.n6669 VGND.t3284 64.3579
R18701 VGND.n1102 VGND.n1101 62.9691
R18702 VGND.n1101 VGND.t2719 61.2134
R18703 VGND.n2433 VGND.t466 60.5809
R18704 VGND.n2555 VGND.t2682 60.5809
R18705 VGND.n5339 VGND.t2755 60.5809
R18706 VGND.n6545 VGND.t2743 60.5809
R18707 VGND.n6043 VGND.t406 60.5809
R18708 VGND.n7007 VGND.t2906 60.5809
R18709 VGND.n4926 VGND.t2882 60.5809
R18710 VGND.n4872 VGND.t2258 60.5809
R18711 VGND.n4713 VGND.t259 60.5809
R18712 VGND.n4257 VGND.t2055 60.5809
R18713 VGND.n4402 VGND.t2610 60.5809
R18714 VGND.n4573 VGND.t1790 60.5809
R18715 VGND.n2935 VGND.t2834 60.5809
R18716 VGND.n2839 VGND.t1705 60.5809
R18717 VGND.n3211 VGND.t2284 60.5809
R18718 VGND.n2670 VGND.t2770 60.5809
R18719 VGND.n3107 VGND.t2914 60.5809
R18720 VGND.n8957 VGND.t36 60.5809
R18721 VGND.n8991 VGND.t2362 60.5809
R18722 VGND.n8495 VGND.t1742 60.5809
R18723 VGND.n168 VGND.t1800 60.5809
R18724 VGND.n221 VGND.t87 60.5809
R18725 VGND.n8020 VGND.t3199 60.5809
R18726 VGND.n7891 VGND.t513 60.5809
R18727 VGND.n339 VGND.t2329 60.5809
R18728 VGND.n7642 VGND.t25 60.5809
R18729 VGND.n8224 VGND.t2342 60.5809
R18730 VGND.n8286 VGND.t756 60.5809
R18731 VGND.n918 VGND.t1602 60.5809
R18732 VGND.n1266 VGND.t2741 60.5809
R18733 VGND.n7362 VGND.t2626 60.5809
R18734 VGND.n6915 VGND.t695 60.5809
R18735 VGND.n6319 VGND.t189 60.5809
R18736 VGND.n6427 VGND.t2371 60.5809
R18737 VGND.n6377 VGND.t3105 60.5809
R18738 VGND.n9106 VGND.t2624 60.5809
R18739 VGND VGND.t2289 59.0043
R18740 VGND.t3093 VGND 59.0043
R18741 VGND.t587 VGND.t649 59.0043
R18742 VGND VGND.t68 59.0043
R18743 VGND.t318 VGND.t1753 59.0043
R18744 VGND VGND.t659 59.0043
R18745 VGND.t3149 VGND.t2068 59.0043
R18746 VGND.t2316 VGND.t3161 59.0043
R18747 VGND.n7133 VGND.n7132 58.7892
R18748 VGND.n4445 VGND.t3122 58.5719
R18749 VGND.n3776 VGND.t75 58.5719
R18750 VGND.n1150 VGND.t2579 58.5719
R18751 VGND.n7453 VGND.t2617 58.5719
R18752 VGND.n2341 VGND.t2043 55.7148
R18753 VGND.n3500 VGND.t2157 55.7148
R18754 VGND.n3499 VGND.t2347 55.7148
R18755 VGND.n2404 VGND.t2972 55.7148
R18756 VGND.n2463 VGND.t603 55.7148
R18757 VGND.n2309 VGND.t2243 55.7148
R18758 VGND.n5672 VGND.t1845 55.7148
R18759 VGND.n5581 VGND.t1788 55.7148
R18760 VGND.n1726 VGND.t2686 55.7148
R18761 VGND.n1645 VGND.t59 55.7148
R18762 VGND.n4038 VGND.t2290 55.7148
R18763 VGND.n4773 VGND.t2251 55.7148
R18764 VGND.n4780 VGND.t211 55.7148
R18765 VGND.n1405 VGND.t2167 55.7148
R18766 VGND.n4380 VGND.t107 55.7148
R18767 VGND.n4642 VGND.t648 55.7148
R18768 VGND.n2042 VGND.t2017 55.7148
R18769 VGND.n3273 VGND.t2463 55.7148
R18770 VGND.n2733 VGND.t2136 55.7148
R18771 VGND.n3684 VGND.t3247 55.7148
R18772 VGND.n8946 VGND.t2635 55.7148
R18773 VGND.n8589 VGND.t3118 55.7148
R18774 VGND.n3774 VGND.t2668 55.7148
R18775 VGND.n8632 VGND.t3034 55.7148
R18776 VGND.n8351 VGND.t2319 55.7148
R18777 VGND.n8382 VGND.t523 55.7148
R18778 VGND.n8395 VGND.t1634 55.7148
R18779 VGND.n1977 VGND.t2380 55.7148
R18780 VGND.n709 VGND.t2386 55.7148
R18781 VGND.n7643 VGND.t2563 55.7148
R18782 VGND.n905 VGND.t3098 55.7148
R18783 VGND.n922 VGND.t2524 55.7148
R18784 VGND.n1231 VGND.t3238 55.7148
R18785 VGND.n7474 VGND.t489 55.7148
R18786 VGND.n6448 VGND.t814 55.7148
R18787 VGND.n6132 VGND.t3137 55.7148
R18788 VGND.n6131 VGND.t1993 55.7148
R18789 VGND.n6142 VGND.t2633 55.7148
R18790 VGND.n6141 VGND.t174 55.7148
R18791 VGND.n9107 VGND.t721 55.7148
R18792 VGND.n9113 VGND.t2444 55.7148
R18793 VGND.n3867 VGND.t547 55.3018
R18794 VGND.n3944 VGND.t713 55.3018
R18795 VGND.n1935 VGND.t3152 55.3018
R18796 VGND.n3858 VGND.t549 54.2862
R18797 VGND.n3884 VGND.t711 54.2862
R18798 VGND.n1944 VGND.t3150 54.2862
R18799 VGND.n4551 VGND.t3251 52.8576
R18800 VGND.n4440 VGND.t3127 52.8576
R18801 VGND.n8771 VGND.t788 52.8576
R18802 VGND.n1890 VGND.t2614 52.8576
R18803 VGND.n3522 VGND.t203 51.4291
R18804 VGND.n2356 VGND.t1867 51.4291
R18805 VGND.n2290 VGND.t3136 51.4291
R18806 VGND.n2226 VGND.t93 51.4291
R18807 VGND.n2181 VGND.t2777 51.4291
R18808 VGND.n5128 VGND.t1726 51.4291
R18809 VGND.n5730 VGND.t2011 51.4291
R18810 VGND.n5533 VGND.t3113 51.4291
R18811 VGND.n5113 VGND.t419 51.4291
R18812 VGND.n5108 VGND.t715 51.4291
R18813 VGND.n1838 VGND.t2753 51.4291
R18814 VGND.n3994 VGND.t1955 51.4291
R18815 VGND.n2905 VGND.t1857 51.4291
R18816 VGND.n2678 VGND.t160 51.4291
R18817 VGND.n8470 VGND.t3063 51.4291
R18818 VGND.n8364 VGND.t1630 51.4291
R18819 VGND.n346 VGND.t3096 51.4291
R18820 VGND.n8257 VGND.t2495 51.4291
R18821 VGND.n6902 VGND.t2998 51.4291
R18822 VGND.n9103 VGND.t2854 51.4291
R18823 VGND.t58 VGND 50.5752
R18824 VGND.t475 VGND.t409 50.5752
R18825 VGND.t424 VGND.t2872 50.5752
R18826 VGND.t1300 VGND.t2181 50.5752
R18827 VGND.t558 VGND.t2990 50.5752
R18828 VGND.t2484 VGND 50.5752
R18829 VGND.t1349 VGND.t762 50.5752
R18830 VGND.t899 VGND.t2613 50.5752
R18831 VGND.t368 VGND.t1779 50.5752
R18832 VGND.t150 VGND.t1778 50.5752
R18833 VGND VGND.t125 50.5752
R18834 VGND.t1935 VGND.t1457 50.5752
R18835 VGND.t1909 VGND.t917 50.5752
R18836 VGND.t1643 VGND.t902 50.5752
R18837 VGND.n1340 VGND.t650 43.3851
R18838 VGND.t244 VGND.t2421 42.1461
R18839 VGND.t2369 VGND 42.1461
R18840 VGND.t663 VGND.t2750 42.1461
R18841 VGND.t24 VGND.t2562 42.1461
R18842 VGND.t2919 VGND.t3155 42.1461
R18843 VGND.t74 VGND.t6 42.1461
R18844 VGND.t3051 VGND.t2887 42.1461
R18845 VGND VGND.t2700 42.1461
R18846 VGND.t2449 VGND.t890 42.1461
R18847 VGND.t2714 VGND 42.1461
R18848 VGND.n7544 VGND.t2680 42.0669
R18849 VGND.n1342 VGND.t2098 41.6488
R18850 VGND.n1651 VGND.t57 41.539
R18851 VGND.n6563 VGND.t1817 41.539
R18852 VGND.n6042 VGND.t2632 41.539
R18853 VGND.n6038 VGND.t1901 41.539
R18854 VGND.n4878 VGND.t209 41.539
R18855 VGND.n4882 VGND.t2337 41.539
R18856 VGND.n4459 VGND.t1922 41.539
R18857 VGND.n4463 VGND.t2568 41.539
R18858 VGND.n2705 VGND.t143 41.539
R18859 VGND.n2701 VGND.t470 41.539
R18860 VGND.n7568 VGND.t429 41.539
R18861 VGND.n7564 VGND.t2938 40.6159
R18862 VGND.n2341 VGND.t2265 40.0005
R18863 VGND.n3494 VGND.t2159 40.0005
R18864 VGND.n3494 VGND.t2153 40.0005
R18865 VGND.n3493 VGND.t2348 40.0005
R18866 VGND.n3493 VGND.t2345 40.0005
R18867 VGND.n3500 VGND.t1987 40.0005
R18868 VGND.n3499 VGND.t3 40.0005
R18869 VGND.n2465 VGND.t2039 40.0005
R18870 VGND.n2465 VGND.t2041 40.0005
R18871 VGND.n2309 VGND.t2192 40.0005
R18872 VGND.n2551 VGND.t2245 40.0005
R18873 VGND.n2551 VGND.t2239 40.0005
R18874 VGND.n5672 VGND.t2725 40.0005
R18875 VGND.n5667 VGND.t1849 40.0005
R18876 VGND.n5667 VGND.t1843 40.0005
R18877 VGND.n5581 VGND.t377 40.0005
R18878 VGND.n5576 VGND.t1784 40.0005
R18879 VGND.n5576 VGND.t1786 40.0005
R18880 VGND.n1707 VGND.t2690 40.0005
R18881 VGND.n1707 VGND.t2692 40.0005
R18882 VGND.n1726 VGND.t1594 40.0005
R18883 VGND.n4773 VGND.t474 40.0005
R18884 VGND.n4777 VGND.t2253 40.0005
R18885 VGND.n4777 VGND.t2247 40.0005
R18886 VGND.n1419 VGND.t2169 40.0005
R18887 VGND.n1419 VGND.t2163 40.0005
R18888 VGND.n1405 VGND.t2311 40.0005
R18889 VGND.n4551 VGND.t3054 40.0005
R18890 VGND.n4440 VGND.t2886 40.0005
R18891 VGND.n2042 VGND.t2260 40.0005
R18892 VGND.n2044 VGND.t2019 40.0005
R18893 VGND.n2044 VGND.t2021 40.0005
R18894 VGND.n3666 VGND.t3249 40.0005
R18895 VGND.n3666 VGND.t3243 40.0005
R18896 VGND.n3684 VGND.t2344 40.0005
R18897 VGND.n3786 VGND.t2664 40.0005
R18898 VGND.n3786 VGND.t2666 40.0005
R18899 VGND.n3774 VGND.t7 40.0005
R18900 VGND.n8771 VGND.t3000 40.0005
R18901 VGND.n218 VGND.t3036 40.0005
R18902 VGND.n218 VGND.t3032 40.0005
R18903 VGND.n8632 VGND.t3234 40.0005
R18904 VGND.n8362 VGND.t2320 40.0005
R18905 VGND.n8362 VGND.t2315 40.0005
R18906 VGND.n8351 VGND.t3156 40.0005
R18907 VGND.n8343 VGND.t525 40.0005
R18908 VGND.n8343 VGND.t519 40.0005
R18909 VGND.n8382 VGND.t2487 40.0005
R18910 VGND.n7967 VGND.t369 40.0005
R18911 VGND.n7967 VGND.t371 40.0005
R18912 VGND.n7965 VGND.t361 40.0005
R18913 VGND.n7965 VGND.t365 40.0005
R18914 VGND.n7963 VGND.t357 40.0005
R18915 VGND.n7963 VGND.t359 40.0005
R18916 VGND.n7999 VGND.t351 40.0005
R18917 VGND.n1890 VGND.t2094 40.0005
R18918 VGND.n7959 VGND.t355 40.0005
R18919 VGND.n7959 VGND.t347 40.0005
R18920 VGND.n7956 VGND.t349 40.0005
R18921 VGND.n7956 VGND.t353 40.0005
R18922 VGND.n8010 VGND.t367 40.0005
R18923 VGND.n8010 VGND.t345 40.0005
R18924 VGND.n7954 VGND.t331 40.0005
R18925 VGND.n7954 VGND.t373 40.0005
R18926 VGND.n7952 VGND.t337 40.0005
R18927 VGND.n7952 VGND.t343 40.0005
R18928 VGND.n655 VGND.t845 40.0005
R18929 VGND.n655 VGND.t837 40.0005
R18930 VGND.n608 VGND.t839 40.0005
R18931 VGND.n608 VGND.t832 40.0005
R18932 VGND.n609 VGND.t836 40.0005
R18933 VGND.n609 VGND.t847 40.0005
R18934 VGND.n611 VGND.t828 40.0005
R18935 VGND.n636 VGND.t822 40.0005
R18936 VGND.n636 VGND.t824 40.0005
R18937 VGND.n632 VGND.t818 40.0005
R18938 VGND.n632 VGND.t820 40.0005
R18939 VGND.n626 VGND.t834 40.0005
R18940 VGND.n626 VGND.t826 40.0005
R18941 VGND.n614 VGND.t830 40.0005
R18942 VGND.n614 VGND.t2305 40.0005
R18943 VGND.n616 VGND.t2303 40.0005
R18944 VGND.n616 VGND.t2301 40.0005
R18945 VGND.n1040 VGND.t2104 40.0005
R18946 VGND.n1040 VGND.t2110 40.0005
R18947 VGND.n1212 VGND.t680 40.0005
R18948 VGND.n1212 VGND.t684 40.0005
R18949 VGND.n924 VGND.t2526 40.0005
R18950 VGND.n924 VGND.t2520 40.0005
R18951 VGND.n922 VGND.t28 40.0005
R18952 VGND.n1159 VGND.t670 40.0005
R18953 VGND.n1162 VGND.t676 40.0005
R18954 VGND.n1162 VGND.t678 40.0005
R18955 VGND.n1206 VGND.t656 40.0005
R18956 VGND.n1206 VGND.t658 40.0005
R18957 VGND.n1223 VGND.t674 40.0005
R18958 VGND.n1223 VGND.t666 40.0005
R18959 VGND.n1227 VGND.t668 40.0005
R18960 VGND.n1227 VGND.t672 40.0005
R18961 VGND.n1235 VGND.t654 40.0005
R18962 VGND.n1235 VGND.t664 40.0005
R18963 VGND.n1241 VGND.t313 40.0005
R18964 VGND.n1241 VGND.t660 40.0005
R18965 VGND.n1245 VGND.t315 40.0005
R18966 VGND.n1245 VGND.t319 40.0005
R18967 VGND.n1080 VGND.t329 40.0005
R18968 VGND.n1080 VGND.t333 40.0005
R18969 VGND.n1073 VGND.t2130 40.0005
R18970 VGND.n1073 VGND.t341 40.0005
R18971 VGND.n1011 VGND.t2124 40.0005
R18972 VGND.n1011 VGND.t2126 40.0005
R18973 VGND.n1061 VGND.t2128 40.0005
R18974 VGND.n1061 VGND.t2122 40.0005
R18975 VGND.n1057 VGND.t2120 40.0005
R18976 VGND.n1057 VGND.t2116 40.0005
R18977 VGND.n1052 VGND.t2118 40.0005
R18978 VGND.n1047 VGND.t2100 40.0005
R18979 VGND.n1047 VGND.t2102 40.0005
R18980 VGND.n1013 VGND.t2112 40.0005
R18981 VGND.n1013 VGND.t2114 40.0005
R18982 VGND.n7455 VGND.t493 40.0005
R18983 VGND.n7455 VGND.t495 40.0005
R18984 VGND.n7474 VGND.t573 40.0005
R18985 VGND.n6448 VGND.t2996 40.0005
R18986 VGND.n6126 VGND.t3139 40.0005
R18987 VGND.n6126 VGND.t3140 40.0005
R18988 VGND.n6125 VGND.t1997 40.0005
R18989 VGND.n6125 VGND.t1999 40.0005
R18990 VGND.n6132 VGND.t2622 40.0005
R18991 VGND.n6131 VGND.t81 40.0005
R18992 VGND.n6339 VGND.t812 40.0005
R18993 VGND.n6339 VGND.t816 40.0005
R18994 VGND.n6438 VGND.t2428 40.0005
R18995 VGND.n6438 VGND.t2430 40.0005
R18996 VGND.n6342 VGND.t2420 40.0005
R18997 VGND.n6342 VGND.t2426 40.0005
R18998 VGND.n6425 VGND.t2416 40.0005
R18999 VGND.n6425 VGND.t2418 40.0005
R19000 VGND.n6344 VGND.t2402 40.0005
R19001 VGND.n6416 VGND.t2404 40.0005
R19002 VGND.n6416 VGND.t2432 40.0005
R19003 VGND.n6412 VGND.t2412 40.0005
R19004 VGND.n6412 VGND.t2406 40.0005
R19005 VGND.n6406 VGND.t2408 40.0005
R19006 VGND.n6406 VGND.t2410 40.0005
R19007 VGND.n6398 VGND.t2414 40.0005
R19008 VGND.n6398 VGND.t325 40.0005
R19009 VGND.n6346 VGND.t317 40.0005
R19010 VGND.n6346 VGND.t321 40.0005
R19011 VGND.n9107 VGND.t1932 40.0005
R19012 VGND.n9109 VGND.t717 40.0005
R19013 VGND.n9109 VGND.t719 40.0005
R19014 VGND.n9113 VGND.t3075 40.0005
R19015 VGND.n9116 VGND.t2440 40.0005
R19016 VGND.n9116 VGND.t2442 40.0005
R19017 VGND.n1348 VGND.n1347 39.6134
R19018 VGND.n3943 VGND.n3942 39.6134
R19019 VGND.n669 VGND.n668 39.6134
R19020 VGND.n8086 VGND.n8085 39.6134
R19021 VGND.n1332 VGND.t1945 38.7697
R19022 VGND.n1065 VGND.t2955 38.7697
R19023 VGND.n2488 VGND.t3002 38.5719
R19024 VGND.n2488 VGND.t2065 38.5719
R19025 VGND.n2352 VGND.t434 38.5719
R19026 VGND.n2352 VGND.t2060 38.5719
R19027 VGND.n5205 VGND.t1949 38.5719
R19028 VGND.n5205 VGND.t1746 38.5719
R19029 VGND.n1632 VGND.t2529 38.5719
R19030 VGND.n1632 VGND.t288 38.5719
R19031 VGND.n6022 VGND.t534 38.5719
R19032 VGND.n6022 VGND.t280 38.5719
R19033 VGND.n7018 VGND.t2199 38.5719
R19034 VGND.n7018 VGND.t1760 38.5719
R19035 VGND.n7141 VGND.t2574 38.5719
R19036 VGND.n1342 VGND.t643 38.5719
R19037 VGND.n4079 VGND.t2559 38.5719
R19038 VGND.n4079 VGND.t274 38.5719
R19039 VGND.n4895 VGND.t582 38.5719
R19040 VGND.n4895 VGND.t278 38.5719
R19041 VGND.n4675 VGND.t178 38.5719
R19042 VGND.n4675 VGND.t282 38.5719
R19043 VGND.n4279 VGND.t2235 38.5719
R19044 VGND.n4279 VGND.t276 38.5719
R19045 VGND.n4421 VGND.t2641 38.5719
R19046 VGND.n4421 VGND.t286 38.5719
R19047 VGND.n1438 VGND.t1919 38.5719
R19048 VGND.n1438 VGND.t1756 38.5719
R19049 VGND.n2917 VGND.t592 38.5719
R19050 VGND.n2917 VGND.t1805 38.5719
R19051 VGND.n2859 VGND.t1645 38.5719
R19052 VGND.n2859 VGND.t1811 38.5719
R19053 VGND.n3223 VGND.t2534 38.5719
R19054 VGND.n3223 VGND.t1807 38.5719
R19055 VGND.n2676 VGND.t2088 38.5719
R19056 VGND.n2676 VGND.t2063 38.5719
R19057 VGND.n3129 VGND.t268 38.5719
R19058 VGND.n3129 VGND.t2080 38.5719
R19059 VGND.n9040 VGND.t2454 38.5719
R19060 VGND.n9040 VGND.t2059 38.5719
R19061 VGND.n8974 VGND.t206 38.5719
R19062 VGND.n8974 VGND.t1809 38.5719
R19063 VGND.n8458 VGND.t84 38.5719
R19064 VGND.n8458 VGND.t1815 38.5719
R19065 VGND.n3886 VGND.t1671 38.5719
R19066 VGND.n3878 VGND.t1675 38.5719
R19067 VGND.n3882 VGND.t2890 38.5719
R19068 VGND.n3882 VGND.t1893 38.5719
R19069 VGND.n159 VGND.t3018 38.5719
R19070 VGND.n159 VGND.t1889 38.5719
R19071 VGND.n174 VGND.t1936 38.5719
R19072 VGND.n174 VGND.t1891 38.5719
R19073 VGND.n229 VGND.t1910 38.5719
R19074 VGND.n229 VGND.t2067 38.5719
R19075 VGND.n7999 VGND.t363 38.5719
R19076 VGND.n8003 VGND.t1669 38.5719
R19077 VGND.n8003 VGND.t1758 38.5719
R19078 VGND.n7798 VGND.t1673 38.5719
R19079 VGND.n520 VGND.t1914 38.5719
R19080 VGND.n520 VGND.t1895 38.5719
R19081 VGND.n7903 VGND.t52 38.5719
R19082 VGND.n7903 VGND.t2061 38.5719
R19083 VGND.n344 VGND.t1794 38.5719
R19084 VGND.n344 VGND.t1750 38.5719
R19085 VGND.n442 VGND.t2831 38.5719
R19086 VGND.n442 VGND.t1762 38.5719
R19087 VGND.n7602 VGND.t1897 38.5719
R19088 VGND.n7602 VGND.t763 38.5719
R19089 VGND.n611 VGND.t843 38.5719
R19090 VGND.n8179 VGND.t298 38.5719
R19091 VGND.n8179 VGND.t1764 38.5719
R19092 VGND.n926 VGND.t557 38.5719
R19093 VGND.n926 VGND.t1748 38.5719
R19094 VGND.n1159 VGND.t682 38.5719
R19095 VGND.n1247 VGND.t311 38.5719
R19096 VGND.n1247 VGND.t1754 38.5719
R19097 VGND.n1052 VGND.t2108 38.5719
R19098 VGND.n814 VGND.t2183 38.5719
R19099 VGND.n814 VGND.t1885 38.5719
R19100 VGND.n1527 VGND.t2351 38.5719
R19101 VGND.n1527 VGND.t1752 38.5719
R19102 VGND.n6296 VGND.t1736 38.5719
R19103 VGND.n6296 VGND.t272 38.5719
R19104 VGND.n6344 VGND.t2424 38.5719
R19105 VGND.n6397 VGND.t2332 38.5719
R19106 VGND.n6397 VGND.t284 38.5719
R19107 VGND.n6348 VGND.t290 38.5719
R19108 VGND.n6348 VGND.t2367 38.5719
R19109 VGND.n9114 VGND.t567 38.5719
R19110 VGND.n9114 VGND.t1813 38.5719
R19111 VGND.n3839 VGND.n3838 37.2945
R19112 VGND.n6224 VGND.n6223 37.2945
R19113 VGND.n4221 VGND.t1835 36.9236
R19114 VGND.n7132 VGND.t2092 36.0005
R19115 VGND.n7132 VGND.t397 36.0005
R19116 VGND.n5074 VGND.t2960 36.0005
R19117 VGND.n5017 VGND.t2210 36.0005
R19118 VGND.n1101 VGND.t2296 35.03
R19119 VGND.n7139 VGND.n7138 34.6358
R19120 VGND.n7925 VGND.n7905 34.6358
R19121 VGND.n2459 VGND.n2458 34.6358
R19122 VGND.n2546 VGND.n2545 34.6358
R19123 VGND.n5933 VGND.n5932 34.6358
R19124 VGND.n1823 VGND.n1797 34.6358
R19125 VGND.n5403 VGND.n5402 34.6358
R19126 VGND.n6641 VGND.n6640 34.6358
R19127 VGND.n6036 VGND.n6035 34.6358
R19128 VGND.n6035 VGND.n6018 34.6358
R19129 VGND.n6588 VGND.n6587 34.6358
R19130 VGND.n7122 VGND.n7121 34.6358
R19131 VGND.n7138 VGND.n1349 34.6358
R19132 VGND.n7187 VGND.n7186 34.6358
R19133 VGND.n7191 VGND.n7190 34.6358
R19134 VGND.n4025 VGND.n3993 34.6358
R19135 VGND.n5020 VGND.n5016 34.6358
R19136 VGND.n4888 VGND.n4887 34.6358
R19137 VGND.n4788 VGND.n4787 34.6358
R19138 VGND.n4285 VGND.n4284 34.6358
R19139 VGND.n4387 VGND.n4223 34.6358
R19140 VGND.n4391 VGND.n4223 34.6358
R19141 VGND.n1451 VGND.n1450 34.6358
R19142 VGND.n2933 VGND.n2932 34.6358
R19143 VGND.n2848 VGND.n2752 34.6358
R19144 VGND.n2699 VGND.n2698 34.6358
R19145 VGND.n3845 VGND.n1865 34.6358
R19146 VGND.n8392 VGND.n8391 34.6358
R19147 VGND.n8403 VGND.n8402 34.6358
R19148 VGND.n1908 VGND.n1877 34.6358
R19149 VGND.n8001 VGND.n8000 34.6358
R19150 VGND.n8026 VGND.n8025 34.6358
R19151 VGND.n7887 VGND.n497 34.6358
R19152 VGND.n7638 VGND.n7637 34.6358
R19153 VGND.n940 VGND.n939 34.6358
R19154 VGND.n945 VGND.n919 34.6358
R19155 VGND.n1276 VGND.n1275 34.6358
R19156 VGND.n1032 VGND.n1029 34.6358
R19157 VGND.n6137 VGND.n6136 34.6358
R19158 VGND.n6280 VGND.n6279 34.6358
R19159 VGND.n9156 VGND.t3412 34.2973
R19160 VGND.n2298 VGND.t3450 34.2973
R19161 VGND.n5555 VGND.t3419 34.2973
R19162 VGND.n5653 VGND.t3504 34.2973
R19163 VGND.n5690 VGND.t3488 34.2973
R19164 VGND.n4595 VGND.t3462 34.2973
R19165 VGND.n4559 VGND.t3351 34.2973
R19166 VGND.n2950 VGND.t3406 34.2973
R19167 VGND.n2753 VGND.t3335 34.2973
R19168 VGND.n3216 VGND.t3457 34.2973
R19169 VGND.n3300 VGND.t3435 34.2973
R19170 VGND.n2722 VGND.t3275 34.2973
R19171 VGND.n8928 VGND.t3292 34.2973
R19172 VGND.n249 VGND.t3477 34.2973
R19173 VGND.n8510 VGND.t3444 34.2973
R19174 VGND.n3963 VGND.t3342 34.2973
R19175 VGND.n209 VGND.t3328 34.2973
R19176 VGND.n8601 VGND.t3475 34.2973
R19177 VGND.n7895 VGND.t3447 34.2973
R19178 VGND.n7861 VGND.t3470 34.2973
R19179 VGND.n511 VGND.t3270 34.2973
R19180 VGND.n363 VGND.t3460 34.2973
R19181 VGND.n8226 VGND.t3439 34.2973
R19182 VGND.n963 VGND.t3318 34.2973
R19183 VGND.n7418 VGND.t3499 34.2973
R19184 VGND.n1008 VGND.t3408 34.2973
R19185 VGND.n6246 VGND.t3321 34.2973
R19186 VGND.n8363 VGND.n8350 34.2593
R19187 VGND.n7121 VGND.n1351 33.8829
R19188 VGND.n7182 VGND.n7181 33.8829
R19189 VGND.n7172 VGND.n7171 33.8829
R19190 VGND.n4027 VGND.n4026 33.8829
R19191 VGND.n5055 VGND.n5054 33.8829
R19192 VGND.n4637 VGND.n4636 33.8829
R19193 VGND.n1253 VGND.n1252 33.8829
R19194 VGND.t2661 VGND.t1557 33.717
R19195 VGND.t1735 VGND.t1898 33.717
R19196 VGND.t595 VGND.t271 33.717
R19197 VGND.t411 VGND.t2234 33.717
R19198 VGND.t275 VGND.t600 33.717
R19199 VGND.t2162 VGND.t1397 33.717
R19200 VGND.t758 VGND.t3179 33.717
R19201 VGND.t273 VGND.t774 33.717
R19202 VGND.t1954 VGND.t2570 33.717
R19203 VGND.t2214 VGND.t2325 33.717
R19204 VGND.t2182 VGND.t2374 33.717
R19205 VGND.t1791 VGND.t1795 33.717
R19206 VGND.t1615 VGND.t3023 33.717
R19207 VGND.t51 VGND.t480 33.717
R19208 VGND.t2453 VGND.t1961 33.717
R19209 VGND.t1825 VGND.t2058 33.717
R19210 VGND.t1804 VGND.t1856 33.717
R19211 VGND.t2921 VGND.t445 33.717
R19212 VGND.t2439 VGND.t1812 33.717
R19213 VGND.n7195 VGND.n7194 33.5064
R19214 VGND.n3042 VGND.n3037 33.5064
R19215 VGND.n2337 VGND.t95 33.462
R19216 VGND.n2337 VGND.t2922 33.462
R19217 VGND.n5131 VGND.t3224 33.462
R19218 VGND.n5131 VGND.t2912 33.462
R19219 VGND.n1818 VGND.t3109 33.462
R19220 VGND.n1818 VGND.t2551 33.462
R19221 VGND.n1633 VGND.t1622 33.462
R19222 VGND.n1633 VGND.t48 33.462
R19223 VGND.n1725 VGND.t2047 33.462
R19224 VGND.n1725 VGND.t431 33.462
R19225 VGND.n4790 VGND.t571 33.462
R19226 VGND.n4790 VGND.t1744 33.462
R19227 VGND.n3988 VGND.t2871 33.462
R19228 VGND.n3988 VGND.t294 33.462
R19229 VGND.n4076 VGND.t775 33.462
R19230 VGND.n4076 VGND.t709 33.462
R19231 VGND.n4908 VGND.t652 33.462
R19232 VGND.n4908 VGND.t759 33.462
R19233 VGND.n4712 VGND.t781 33.462
R19234 VGND.n4712 VGND.t263 33.462
R19235 VGND.n1403 VGND.t1740 33.462
R19236 VGND.n1403 VGND.t1654 33.462
R19237 VGND.n4164 VGND.t2647 33.462
R19238 VGND.n4164 VGND.t2860 33.462
R19239 VGND.n4105 VGND.t2281 33.462
R19240 VGND.n4105 VGND.t410 33.462
R19241 VGND.n4112 VGND.t1863 33.462
R19242 VGND.n4112 VGND.t2499 33.462
R19243 VGND.n1390 VGND.t2033 33.462
R19244 VGND.n1390 VGND.t2828 33.462
R19245 VGND.n2843 VGND.t1953 33.462
R19246 VGND.n2843 VGND.t2220 33.462
R19247 VGND.n2653 VGND.t2927 33.462
R19248 VGND.n2653 VGND.t2208 33.462
R19249 VGND.n8917 VGND.t555 33.462
R19250 VGND.n8917 VGND.t1841 33.462
R19251 VGND.n90 VGND.t2630 33.462
R19252 VGND.n90 VGND.t1798 33.462
R19253 VGND.n193 VGND.t479 33.462
R19254 VGND.n193 VGND.t579 33.462
R19255 VGND.n3846 VGND.t3080 33.462
R19256 VGND.n3846 VGND.t586 33.462
R19257 VGND.n3921 VGND.t690 33.462
R19258 VGND.n3921 VGND.t1624 33.462
R19259 VGND.n7902 VGND.t481 33.462
R19260 VGND.n7902 VGND.t1926 33.462
R19261 VGND.n7949 VGND.t2675 33.462
R19262 VGND.n7949 VGND.t2003 33.462
R19263 VGND.n337 VGND.t3142 33.462
R19264 VGND.n337 VGND.t1792 33.462
R19265 VGND.n698 VGND.t1641 33.462
R19266 VGND.n698 VGND.t3103 33.462
R19267 VGND.n8142 VGND.t2512 33.462
R19268 VGND.n8142 VGND.t2585 33.462
R19269 VGND.n8270 VGND.t3187 33.462
R19270 VGND.n8270 VGND.t2309 33.462
R19271 VGND.n7473 VGND.t639 33.462
R19272 VGND.n7473 VGND.t468 33.462
R19273 VGND.n1487 VGND.t2001 33.462
R19274 VGND.n1487 VGND.t3107 33.462
R19275 VGND.n1690 VGND.t195 33.462
R19276 VGND.n1690 VGND.t2035 33.462
R19277 VGND.n6212 VGND.t779 33.462
R19278 VGND.n6212 VGND.t1967 33.462
R19279 VGND.n6263 VGND.t1989 33.462
R19280 VGND.n6263 VGND.t1850 33.462
R19281 VGND.n5059 VGND.t497 33.2313
R19282 VGND.n3952 VGND.n3951 32.377
R19283 VGND.n4277 VGND.t601 32.3082
R19284 VGND.n4287 VGND.t594 32.3082
R19285 VGND.n4555 VGND.t2206 32.3082
R19286 VGND.n1397 VGND.t2760 32.3082
R19287 VGND.n2867 VGND.t2394 32.3082
R19288 VGND.n2783 VGND.t1828 32.3082
R19289 VGND.n3028 VGND.t1824 32.3082
R19290 VGND.n9038 VGND.t1826 32.3082
R19291 VGND.n255 VGND.t2388 32.3082
R19292 VGND.n8418 VGND.t2390 32.3082
R19293 VGND.n7961 VGND.t2392 32.3082
R19294 VGND.n812 VGND.t2375 32.3082
R19295 VGND.n6294 VGND.t596 32.3082
R19296 VGND.n1671 VGND.t598 32.3082
R19297 VGND.n1909 VGND.n1908 32.0005
R19298 VGND.n1242 VGND.n1157 31.624
R19299 VGND.n8054 VGND.n8053 31.2476
R19300 VGND.n4020 VGND.n4019 30.8711
R19301 VGND.n6446 VGND.n6445 30.4946
R19302 VGND.n7124 VGND.t2816 30.462
R19303 VGND.n7124 VGND.t1720 30.462
R19304 VGND.n4893 VGND.n4892 29.7417
R19305 VGND.n680 VGND.n679 28.9887
R19306 VGND.n6636 VGND.n1634 28.9887
R19307 VGND.n1036 VGND.n1035 28.9887
R19308 VGND.n1021 VGND.n1018 28.9887
R19309 VGND.n3522 VGND.t733 28.7917
R19310 VGND.n2356 VGND.t105 28.7917
R19311 VGND.n2290 VGND.t3166 28.7917
R19312 VGND.n2226 VGND.t2273 28.7917
R19313 VGND.n2181 VGND.t2029 28.7917
R19314 VGND.n5128 VGND.t3028 28.7917
R19315 VGND.n5730 VGND.t38 28.7917
R19316 VGND.n5533 VGND.t2360 28.7917
R19317 VGND.n5113 VGND.t2953 28.7917
R19318 VGND.n5108 VGND.t1698 28.7917
R19319 VGND.n1838 VGND.t686 28.7917
R19320 VGND.n3994 VGND.t3201 28.7917
R19321 VGND.n2905 VGND.t3172 28.7917
R19322 VGND.n2678 VGND.t2655 28.7917
R19323 VGND.n8470 VGND.t2450 28.7917
R19324 VGND.n8364 VGND.t3164 28.7917
R19325 VGND.n346 VGND.t2731 28.7917
R19326 VGND.n8257 VGND.t23 28.7917
R19327 VGND.n6902 VGND.t2862 28.7917
R19328 VGND.n9103 VGND.t527 28.7917
R19329 VGND.n3927 VGND.n3926 28.6616
R19330 VGND.n9131 VGND.n9111 28.2358
R19331 VGND.n7835 VGND.n504 27.8593
R19332 VGND.n6282 VGND.n6262 27.8593
R19333 VGND.n2404 VGND.t2222 26.8576
R19334 VGND.n2463 VGND.t1596 26.8576
R19335 VGND.n1645 VGND.t2549 26.8576
R19336 VGND.n4038 VGND.t752 26.8576
R19337 VGND.n4780 VGND.t3226 26.8576
R19338 VGND.n4380 VGND.t2866 26.8576
R19339 VGND.n4642 VGND.t464 26.8576
R19340 VGND.n3273 VGND.t2177 26.8576
R19341 VGND.n2733 VGND.t2518 26.8576
R19342 VGND.n8946 VGND.t2672 26.8576
R19343 VGND.n8589 VGND.t2233 26.8576
R19344 VGND.n8395 VGND.t172 26.8576
R19345 VGND.n1977 VGND.t2556 26.8576
R19346 VGND.n709 VGND.t2279 26.8576
R19347 VGND.n7643 VGND.t124 26.8576
R19348 VGND.n905 VGND.t459 26.8576
R19349 VGND.n1231 VGND.t2751 26.8576
R19350 VGND.n6142 VGND.t1771 26.8576
R19351 VGND.n6141 VGND.t118 26.8576
R19352 VGND.n1340 VGND.t2902 26.7697
R19353 VGND.n4457 VGND.t2452 26.7697
R19354 VGND.n3505 VGND.n3504 26.7299
R19355 VGND.n5897 VGND.n5112 26.7299
R19356 VGND.n5080 VGND.n5079 26.7299
R19357 VGND.n3689 VGND.n3665 26.7299
R19358 VGND.n1261 VGND.n1154 26.7299
R19359 VGND.n5505 VGND.n5502 26.6009
R19360 VGND.n3849 VGND.n3845 26.6009
R19361 VGND.n8282 VGND.n8280 26.6009
R19362 VGND.n5163 VGND.n5162 26.314
R19363 VGND.n6592 VGND.n6591 26.314
R19364 VGND.n4275 VGND.n4274 26.314
R19365 VGND.n7651 VGND.n7650 26.314
R19366 VGND.n6893 VGND.n6892 26.314
R19367 VGND.n6303 VGND.n6302 26.314
R19368 VGND.n4027 VGND.n3992 25.977
R19369 VGND.n5086 VGND.n4034 25.977
R19370 VGND.n2928 VGND.n2901 25.977
R19371 VGND.n1222 VGND.n1160 25.977
R19372 VGND.n3858 VGND.t750 25.9346
R19373 VGND.n3884 VGND.t541 25.9346
R19374 VGND.n1944 VGND.t191 25.9346
R19375 VGND.n7841 VGND.t302 25.9346
R19376 VGND.n8047 VGND.n8046 25.7355
R19377 VGND.n2480 VGND.n2479 25.7355
R19378 VGND.n5141 VGND.n5140 25.7355
R19379 VGND.n5736 VGND.n5734 25.7355
R19380 VGND.n5587 VGND.n5585 25.7355
R19381 VGND.n6628 VGND.n1637 25.7355
R19382 VGND.n7147 VGND.n7146 25.7355
R19383 VGND.n5068 VGND.n5067 25.7355
R19384 VGND.n5063 VGND.n5058 25.7355
R19385 VGND.n7846 VGND.n7840 25.7355
R19386 VGND.n7346 VGND.n7345 25.7355
R19387 VGND.n6292 VGND.n6291 25.7355
R19388 VGND.n5541 VGND.n5539 25.6926
R19389 VGND.n1816 VGND.n1815 25.6926
R19390 VGND.n1731 VGND.n1706 25.6926
R19391 VGND.n7118 VGND.n7117 25.6926
R19392 VGND.n4118 VGND.n4116 25.6926
R19393 VGND.n4694 VGND.n4693 25.6926
R19394 VGND.n4686 VGND.n4685 25.6926
R19395 VGND.n4673 VGND.n4672 25.6926
R19396 VGND.n4636 VGND.n4556 25.6926
R19397 VGND.n2850 VGND.n2848 25.6926
R19398 VGND.n3263 VGND.n3214 25.6926
R19399 VGND.n8478 VGND.n8477 25.6926
R19400 VGND.n8493 VGND.n8492 25.6926
R19401 VGND.n8765 VGND.n8764 25.6926
R19402 VGND.n8391 VGND.n8342 25.6926
R19403 VGND.n8031 VGND.n8030 25.6926
R19404 VGND.n378 VGND.n377 25.6926
R19405 VGND.n703 VGND.n691 25.6926
R19406 VGND.n7637 VGND.n7609 25.6926
R19407 VGND.n679 VGND.n606 25.6926
R19408 VGND.n8244 VGND.n8243 25.6926
R19409 VGND.n1076 VGND.n1072 25.6926
R19410 VGND.n6911 VGND.n6909 25.6926
R19411 VGND.n6227 VGND.n6222 25.6926
R19412 VGND.n3043 VGND.n3042 25.6005
R19413 VGND.n1932 VGND.n1931 25.6005
R19414 VGND.n948 VGND.n917 25.6005
R19415 VGND.n9124 VGND.n9117 25.6005
R19416 VGND.n1723 VGND.n1722 25.5964
R19417 VGND.n7471 VGND.n7470 25.5964
R19418 VGND.n8064 VGND.n8063 25.4884
R19419 VGND.n8188 VGND.n8187 25.4715
R19420 VGND.n7126 VGND.t641 25.4291
R19421 VGND.n4445 VGND.t2307 25.4291
R19422 VGND.n3776 VGND.t2894 25.4291
R19423 VGND.n3930 VGND.t2007 25.4291
R19424 VGND.n480 VGND.t448 25.4291
R19425 VGND.n654 VGND.t2049 25.4291
R19426 VGND.n2545 VGND.n2313 25.4203
R19427 VGND.n4479 VGND.n4476 25.4203
R19428 VGND.n7921 VGND.n7920 25.4203
R19429 VGND.t322 VGND.t2366 25.2879
R19430 VGND.t2376 VGND.t2609 25.2879
R19431 VGND.t338 VGND.t1065 25.2879
R19432 VGND.t3151 VGND.t2949 25.2879
R19433 VGND.t3037 VGND.t1644 25.2879
R19434 VGND.n3505 VGND.n3484 25.224
R19435 VGND.n2413 VGND.n2354 25.224
R19436 VGND.n6054 VGND.n6053 25.224
R19437 VGND.n6584 VGND.n6583 25.224
R19438 VGND.n4107 VGND.n4097 25.224
R19439 VGND.n2932 VGND.n2901 25.224
R19440 VGND.n8753 VGND.n172 25.224
R19441 VGND.n652 VGND.n651 25.224
R19442 VGND.n1261 VGND.n1260 25.224
R19443 VGND.n7480 VGND.n7479 25.224
R19444 VGND.n8940 VGND.n8939 24.9894
R19445 VGND.n8638 VGND.n8637 24.9894
R19446 VGND.n7926 VGND.n7925 24.9894
R19447 VGND.n1098 VGND.n886 24.9894
R19448 VGND.n7453 VGND.t3190 24.9236
R19449 VGND.n1350 VGND.t2818 24.9236
R19450 VGND.n1350 VGND.t745 24.9236
R19451 VGND.n7157 VGND.t2898 24.9236
R19452 VGND.n7157 VGND.t2900 24.9236
R19453 VGND.n1338 VGND.t399 24.9236
R19454 VGND.n1338 VGND.t451 24.9236
R19455 VGND.n1336 VGND.t2958 24.9236
R19456 VGND.n1336 VGND.t1822 24.9236
R19457 VGND.n1334 VGND.t1709 24.9236
R19458 VGND.n1334 VGND.t646 24.9236
R19459 VGND.n7199 VGND.t2262 24.9236
R19460 VGND.n7199 VGND.t3092 24.9236
R19461 VGND.n3996 VGND.t2581 24.9236
R19462 VGND.n3996 VGND.t738 24.9236
R19463 VGND.n4013 VGND.t743 24.9236
R19464 VGND.n4013 VGND.t2292 24.9236
R19465 VGND.n5074 VGND.t32 24.9236
R19466 VGND.n5075 VGND.t1696 24.9236
R19467 VGND.n5075 VGND.t1694 24.9236
R19468 VGND.n5059 VGND.t2151 24.9236
R19469 VGND.n5033 VGND.t2149 24.9236
R19470 VGND.n5033 VGND.t2213 24.9236
R19471 VGND.n5037 VGND.t13 24.9236
R19472 VGND.n5037 VGND.t15 24.9236
R19473 VGND.n5029 VGND.t1659 24.9236
R19474 VGND.n5029 VGND.t17 24.9236
R19475 VGND.n4041 VGND.t1665 24.9236
R19476 VGND.n4041 VGND.t1663 24.9236
R19477 VGND.n5017 VGND.t5 24.9236
R19478 VGND.n4277 VGND.t412 24.9236
R19479 VGND.n4287 VGND.t1903 24.9236
R19480 VGND.n4221 VGND.t771 24.9236
R19481 VGND.n4408 VGND.t777 24.9236
R19482 VGND.n4408 VGND.t423 24.9236
R19483 VGND.n4413 VGND.t425 24.9236
R19484 VGND.n4413 VGND.t421 24.9236
R19485 VGND.n4214 VGND.t382 24.9236
R19486 VGND.n4214 VGND.t1983 24.9236
R19487 VGND.n4526 VGND.t114 24.9236
R19488 VGND.n4526 VGND.t1732 24.9236
R19489 VGND.n4555 VGND.t2884 24.9236
R19490 VGND.n4626 VGND.t699 24.9236
R19491 VGND.n4626 VGND.t3216 24.9236
R19492 VGND.n4619 VGND.t3210 24.9236
R19493 VGND.n4619 VGND.t3208 24.9236
R19494 VGND.n4557 VGND.t3214 24.9236
R19495 VGND.n4557 VGND.t3218 24.9236
R19496 VGND.n1397 VGND.t2005 24.9236
R19497 VGND.n2867 VGND.t1770 24.9236
R19498 VGND.n2783 VGND.t44 24.9236
R19499 VGND.n3028 VGND.t2179 24.9236
R19500 VGND.n9038 VGND.t1962 24.9236
R19501 VGND.n255 VGND.t2888 24.9236
R19502 VGND.n3804 VGND.t2947 24.9236
R19503 VGND.n3804 VGND.t2942 24.9236
R19504 VGND.n8418 VGND.t2875 24.9236
R19505 VGND.n7961 VGND.t1767 24.9236
R19506 VGND.n1911 VGND.t803 24.9236
R19507 VGND.n1911 VGND.t806 24.9236
R19508 VGND.n489 VGND.t727 24.9236
R19509 VGND.n489 VGND.t731 24.9236
R19510 VGND.n486 VGND.t3189 24.9236
R19511 VGND.n486 VGND.t729 24.9236
R19512 VGND.n487 VGND.t2591 24.9236
R19513 VGND.n487 VGND.t2595 24.9236
R19514 VGND.n484 VGND.t2589 24.9236
R19515 VGND.n484 VGND.t2597 24.9236
R19516 VGND.n481 VGND.t392 24.9236
R19517 VGND.n481 VGND.t2593 24.9236
R19518 VGND.n1943 VGND.t2175 24.9236
R19519 VGND.n1943 VGND.t2069 24.9236
R19520 VGND.n7836 VGND.t3024 24.9236
R19521 VGND.n7836 VGND.t1973 24.9236
R19522 VGND.n7874 VGND.t2987 24.9236
R19523 VGND.n7874 VGND.t1971 24.9236
R19524 VGND.n685 VGND.t2186 24.9236
R19525 VGND.n685 VGND.t2071 24.9236
R19526 VGND.n646 VGND.t2501 24.9236
R19527 VGND.n646 VGND.t2506 24.9236
R19528 VGND.n8164 VGND.t386 24.9236
R19529 VGND.n8164 VGND.t2354 24.9236
R19530 VGND.n1065 VGND.t2983 24.9236
R19531 VGND.n1014 VGND.t67 24.9236
R19532 VGND.n1014 VGND.t563 24.9236
R19533 VGND.n1017 VGND.t69 24.9236
R19534 VGND.n1017 VGND.t65 24.9236
R19535 VGND.n7317 VGND.t71 24.9236
R19536 VGND.n7317 VGND.t61 24.9236
R19537 VGND.n812 VGND.t707 24.9236
R19538 VGND.n7399 VGND.t2599 24.9236
R19539 VGND.n7399 VGND.t2603 24.9236
R19540 VGND.n789 VGND.t1839 24.9236
R19541 VGND.n789 VGND.t1837 24.9236
R19542 VGND.n6879 VGND.t505 24.9236
R19543 VGND.n6879 VGND.t511 24.9236
R19544 VGND.n6886 VGND.t503 24.9236
R19545 VGND.n6886 VGND.t509 24.9236
R19546 VGND.n1583 VGND.t501 24.9236
R19547 VGND.n1583 VGND.t3056 24.9236
R19548 VGND.n6830 VGND.t1957 24.9236
R19549 VGND.n6830 VGND.t2545 24.9236
R19550 VGND.n6838 VGND.t2541 24.9236
R19551 VGND.n6838 VGND.t2537 24.9236
R19552 VGND.n6844 VGND.t2543 24.9236
R19553 VGND.n6844 VGND.t2547 24.9236
R19554 VGND.n6294 VGND.t1899 24.9236
R19555 VGND.n1671 VGND.t2327 24.9236
R19556 VGND.n2413 VGND.n2412 24.8476
R19557 VGND.n5162 VGND.n5129 24.8476
R19558 VGND.n5897 VGND.n5896 24.8476
R19559 VGND.n4020 VGND.n3995 24.8476
R19560 VGND.n4392 VGND.n4391 24.8476
R19561 VGND.n8637 VGND.n217 24.8476
R19562 VGND.n8246 VGND.n454 24.8476
R19563 VGND.n6897 VGND.n1582 24.8476
R19564 VGND.n9149 VGND.n9104 24.8476
R19565 VGND.n4774 VGND.n4766 24.4711
R19566 VGND.n4442 VGND.n4441 24.4711
R19567 VGND.n8775 VGND.n8774 24.4711
R19568 VGND.n8371 VGND.n8349 24.4711
R19569 VGND.n8371 VGND.n8370 24.4711
R19570 VGND.n940 VGND.n920 24.4711
R19571 VGND.n939 VGND.n923 24.4711
R19572 VGND.n6454 VGND.n6453 24.4711
R19573 VGND.n6670 VGND.n6669 24.2743
R19574 VGND.n8042 VGND.n8041 24.2297
R19575 VGND.n4665 VGND.n4167 24.1867
R19576 VGND.n3509 VGND.n3484 24.0946
R19577 VGND.n1824 VGND.n1823 24.0946
R19578 VGND.n4775 VGND.n4774 24.0946
R19579 VGND.n8765 VGND.n167 24.0946
R19580 VGND.n8370 VGND.n8350 24.0946
R19581 VGND.n7988 VGND.n7968 24.0946
R19582 VGND.n6898 VGND.n6897 24.0946
R19583 VGND.n9142 VGND.n9105 24.0946
R19584 VGND.n1150 VGND.t3120 24.0005
R19585 VGND.n8252 VGND.n451 23.7181
R19586 VGND.n2454 VGND.n20 23.7181
R19587 VGND.n5148 VGND.n5145 23.7181
R19588 VGND.n5675 VGND.n5125 23.7181
R19589 VGND.n5815 VGND.n5123 23.7181
R19590 VGND.n7171 VGND.n1335 23.7181
R19591 VGND.n5087 VGND.n3987 23.7181
R19592 VGND.n5087 VGND.n5086 23.7181
R19593 VGND.n5082 VGND.n4034 23.7181
R19594 VGND.n5016 VGND.n3986 23.7181
R19595 VGND.n4769 VGND.n4766 23.7181
R19596 VGND.n1402 VGND.n1401 23.7181
R19597 VGND.n4101 VGND.n4098 23.7181
R19598 VGND.n4442 VGND.n4169 23.7181
R19599 VGND.n4473 VGND.n4215 23.7181
R19600 VGND.n3265 VGND.n3264 23.7181
R19601 VGND.n3264 VGND.n3263 23.7181
R19602 VGND.n8979 VGND.n77 23.7181
R19603 VGND.n8775 VGND.n166 23.7181
R19604 VGND.n1955 VGND.n1954 23.7181
R19605 VGND.n1949 VGND.n1928 23.7181
R19606 VGND.n7810 VGND.n508 23.7181
R19607 VGND.n7941 VGND.n497 23.7181
R19608 VGND.n697 VGND.n694 23.7181
R19609 VGND.n8259 VGND.n8255 23.7181
R19610 VGND.n8268 VGND.n8267 23.7181
R19611 VGND.n1269 VGND.n887 23.7181
R19612 VGND.n1272 VGND.n887 23.7181
R19613 VGND.n7479 VGND.n7454 23.7181
R19614 VGND.n6858 VGND.n6857 23.7181
R19615 VGND.n6336 VGND.n6335 23.7181
R19616 VGND.n2454 VGND.n2453 23.2027
R19617 VGND.n3802 VGND.n3801 23.1002
R19618 VGND.n8357 VGND.n8356 22.9652
R19619 VGND.n3510 VGND.n3509 22.9652
R19620 VGND.n6024 VGND.n6023 22.9652
R19621 VGND.n7837 VGND.n7835 22.9652
R19622 VGND.n7831 VGND.n7830 22.9257
R19623 VGND.n8903 VGND.n8902 22.9058
R19624 VGND.n2485 VGND.n2484 22.5887
R19625 VGND.n619 VGND.n451 22.5887
R19626 VGND.n6645 VGND.t442 22.3257
R19627 VGND.n6027 VGND.t193 22.3257
R19628 VGND.n4896 VGND.t2850 22.3257
R19629 VGND.n4679 VGND.t2924 22.3257
R19630 VGND.n1902 VGND.t2660 22.3257
R19631 VGND.n452 VGND.t168 22.3257
R19632 VGND.n1041 VGND.t768 22.3257
R19633 VGND.n1104 VGND.n1102 22.3044
R19634 VGND.n2480 VGND.n2338 22.2123
R19635 VGND.n2484 VGND.n2338 22.2123
R19636 VGND.n6637 VGND.n6636 22.2123
R19637 VGND.n1404 VGND.n1402 22.2123
R19638 VGND.n4106 VGND.n4098 22.2123
R19639 VGND.n4107 VGND.n4106 22.2123
R19640 VGND.n1450 VGND.n1391 22.2123
R19641 VGND.n3923 VGND.n3922 22.2123
R19642 VGND.n8376 VGND.n8346 22.2123
R19643 VGND.n8030 VGND.n7950 22.2123
R19644 VGND.n382 VGND.n338 22.2123
R19645 VGND.n699 VGND.n697 22.2123
R19646 VGND.n699 VGND.n691 22.2123
R19647 VGND.n6222 VGND.n1692 22.2123
R19648 VGND.n6279 VGND.n6264 22.2123
R19649 VGND.n1587 VGND.t120 22.1912
R19650 VGND.n3990 VGND.t1981 22.0959
R19651 VGND.n8063 VGND.n479 21.8358
R19652 VGND.n664 VGND.n663 21.5514
R19653 VGND.n6654 VGND.n6653 21.4593
R19654 VGND.n7159 VGND.n7158 21.4593
R19655 VGND.n7182 VGND.n1333 21.4593
R19656 VGND.n7190 VGND.n1331 21.4593
R19657 VGND.n7194 VGND.n1329 21.4593
R19658 VGND.n1023 VGND.n1022 21.4593
R19659 VGND.n8259 VGND.n8258 21.2097
R19660 VGND.n5417 VGND.n5204 20.966
R19661 VGND.n4425 VGND.n4420 20.7985
R19662 VGND.n8001 VGND.n7960 20.7064
R19663 VGND.n3978 VGND.n3977 20.422
R19664 VGND.n8624 VGND.n8623 20.3299
R19665 VGND.n8022 VGND.n8021 20.3299
R19666 VGND.n9141 VGND.n9140 20.3299
R19667 VGND.n6671 VGND.n6670 20.103
R19668 VGND.n2679 VGND.n2675 19.9534
R19669 VGND.n357 VGND.n347 19.9534
R19670 VGND.n947 VGND.n946 19.9534
R19671 VGND.n5904 VGND.n5903 19.914
R19672 VGND.n2412 VGND.n2355 19.577
R19673 VGND.n3995 VGND.n3993 19.577
R19674 VGND.n2913 VGND.n2906 19.577
R19675 VGND.n1163 VGND.n1161 19.577
R19676 VGND.n9130 VGND.n9129 19.577
R19677 VGND.n2473 VGND.n2472 19.3355
R19678 VGND.n6287 VGND.n6286 19.3355
R19679 VGND.n2561 VGND.n2560 19.2926
R19680 VGND.n5572 VGND.n5571 19.2926
R19681 VGND.n2964 VGND.n2896 19.2926
R19682 VGND.n8750 VGND.n173 19.2926
R19683 VGND.n3682 VGND.n3681 19.1964
R19684 VGND.n2864 VGND.n2863 18.824
R19685 VGND.n2791 VGND.n2790 18.824
R19686 VGND.n3044 VGND.n3043 18.824
R19687 VGND.n8249 VGND.n453 18.824
R19688 VGND.n5663 VGND.n5662 18.5894
R19689 VGND.n2820 VGND.n2819 18.5894
R19690 VGND.n3248 VGND.n3247 18.5894
R19691 VGND.n4458 VGND.n4216 18.5826
R19692 VGND.n5402 VGND.n5340 18.4613
R19693 VGND.n6332 VGND.n6331 18.3084
R19694 VGND.n2190 VGND.n2189 18.2791
R19695 VGND.n7043 VGND.n7042 18.2791
R19696 VGND.n3105 VGND.n3103 18.2791
R19697 VGND.n3078 VGND.n3076 18.2791
R19698 VGND.n7584 VGND.n7583 18.1
R19699 VGND.n622 VGND.n615 18.0711
R19700 VGND.n1243 VGND.n1242 18.0711
R19701 VGND.n6827 VGND.n1591 18.0105
R19702 VGND.n5965 VGND.n5964 17.7007
R19703 VGND.n8276 VGND.n8274 17.6946
R19704 VGND.n4920 VGND.n4918 17.6577
R19705 VGND.n1113 VGND.n1111 17.6577
R19706 VGND.n6864 VGND.n6861 17.5656
R19707 VGND.n2061 VGND.n2059 17.5615
R19708 VGND.n4522 VGND.n4521 17.4535
R19709 VGND.n3489 VGND.n3488 17.3181
R19710 VGND.n3781 VGND.n3778 17.3181
R19711 VGND.n931 VGND.n928 17.3181
R19712 VGND.n7484 VGND.n7483 17.3181
R19713 VGND.n6121 VGND.n6120 17.3181
R19714 VGND.n9121 VGND.n9118 17.3181
R19715 VGND.n2658 VGND.n2657 17.2527
R19716 VGND.n234 VGND.n233 17.2527
R19717 VGND.n5261 VGND.n5260 17.1563
R19718 VGND.n716 VGND.n715 17.0312
R19719 VGND.n5418 VGND.n5417 16.9936
R19720 VGND.n6621 VGND.n6618 16.9936
R19721 VGND.n7413 VGND.n7412 16.9545
R19722 VGND.n1156 VGND.n1155 16.9417
R19723 VGND.n7767 VGND.n7766 16.9331
R19724 VGND.n7807 VGND.n7806 16.886
R19725 VGND.t1343 VGND.t3194 16.8587
R19726 VGND.t2527 VGND.t56 16.8587
R19727 VGND.t2034 VGND.t1581 16.8587
R19728 VGND.t1376 VGND.t506 16.8587
R19729 VGND.t1391 VGND.t2859 16.8587
R19730 VGND.t2839 VGND.t1205 16.8587
R19731 VGND.t2873 VGND.t108 16.8587
R19732 VGND VGND.t3091 16.8587
R19733 VGND.t2899 VGND.t2097 16.8587
R19734 VGND.t2895 VGND.t2095 16.8587
R19735 VGND.t2321 VGND.t2091 16.8587
R19736 VGND.t1099 VGND.t1838 16.8587
R19737 VGND.t2602 VGND.t1560 16.8587
R19738 VGND.t866 VGND.t2843 16.8587
R19739 VGND.t1775 VGND 16.8587
R19740 VGND.t914 VGND.t524 16.8587
R19741 VGND.t2014 VGND.t2663 16.8587
R19742 VGND.t976 VGND.t578 16.8587
R19743 VGND.t3115 VGND.t911 16.8587
R19744 VGND.t2637 VGND.t2638 16.8587
R19745 VGND.t142 VGND.t2811 16.8587
R19746 VGND.t2193 VGND.t2533 16.8587
R19747 VGND.t2195 VGND.t1806 16.8587
R19748 VGND.t1294 VGND.t43 16.8587
R19749 VGND.t1810 VGND.t606 16.8587
R19750 VGND.t2605 VGND.t1273 16.8587
R19751 VGND.t2443 VGND.t566 16.8587
R19752 VGND.n1809 VGND.n1807 16.7924
R19753 VGND.n8616 VGND.n8615 16.7924
R19754 VGND.n1897 VGND.n1883 16.7924
R19755 VGND.n976 VGND.n975 16.7924
R19756 VGND.n2790 VGND.n2789 16.6573
R19757 VGND.n4904 VGND.n3985 16.5652
R19758 VGND.n6621 VGND.n6620 16.5522
R19759 VGND.n4870 VGND.n4869 16.2808
R19760 VGND.n8485 VGND.n8484 16.2808
R19761 VGND.n2419 VGND.n2418 16.1492
R19762 VGND.n7356 VGND.n7355 16.1492
R19763 VGND.n7151 VGND.n1343 15.9473
R19764 VGND.n4912 VGND.n4910 15.9044
R19765 VGND.n4613 VGND.n4612 15.9044
R19766 VGND.n7855 VGND.n7850 15.9033
R19767 VGND.n1435 VGND.n1434 15.8505
R19768 VGND.n8585 VGND.n8584 15.8505
R19769 VGND.n1524 VGND.n1523 15.8505
R19770 VGND.n4681 VGND.n4680 15.8123
R19771 VGND.n8252 VGND.n453 15.8123
R19772 VGND.n1063 VGND.n1062 15.8123
R19773 VGND.n1043 VGND.n1042 15.8123
R19774 VGND.n5726 VGND.n5725 15.7728
R19775 VGND.n5529 VGND.n5528 15.7728
R19776 VGND.n2619 VGND.n18 15.6833
R19777 VGND.n1446 VGND.n1445 15.6771
R19778 VGND.n1535 VGND.n1534 15.6771
R19779 VGND.n2717 VGND.n2716 15.5776
R19780 VGND.n2925 VGND.n2902 15.5708
R19781 VGND.n5046 VGND.n4039 15.5708
R19782 VGND.n2857 VGND.n2856 15.5279
R19783 VGND.n7128 VGND.n7125 15.4358
R19784 VGND.n1337 VGND.n1335 15.4358
R19785 VGND.n3953 VGND.n3952 15.4358
R19786 VGND.n8349 VGND.n8348 15.4358
R19787 VGND.n5941 VGND.n5940 15.3963
R19788 VGND.n7016 VGND.n7015 15.3963
R19789 VGND.n3979 VGND.n1864 15.3963
R19790 VGND.n1494 VGND.n1493 15.3963
R19791 VGND.n8255 VGND.n449 15.3068
R19792 VGND.n958 VGND.n957 15.2011
R19793 VGND.n5043 VGND.n4040 15.1944
R19794 VGND.n5155 VGND.n5130 15.1514
R19795 VGND.n1423 VGND.n1406 15.1514
R19796 VGND.n4295 VGND.n4293 15.1514
R19797 VGND.n4433 VGND.n4432 15.1259
R19798 VGND.n1925 VGND.n1924 15.1259
R19799 VGND.n4898 VGND.n4897 15.0593
R19800 VGND.n4111 VGND.n4097 15.0593
R19801 VGND.n3840 VGND.n3839 15.0593
R19802 VGND.n1920 VGND.n1919 15.0593
R19803 VGND.n6624 VGND.n6623 15.0266
R19804 VGND.n7788 VGND.n7787 14.9303
R19805 VGND.n2943 VGND.n2942 14.8247
R19806 VGND.n8503 VGND.n8502 14.8247
R19807 VGND.n1717 VGND.n1714 14.8179
R19808 VGND.n4657 VGND.n4656 14.8179
R19809 VGND.n2054 VGND.n2051 14.8179
R19810 VGND.n3676 VGND.n3673 14.8179
R19811 VGND.n7465 VGND.n7462 14.8179
R19812 VGND.n6390 VGND.n6350 14.8179
R19813 VGND.n6385 VGND.n6384 14.8179
R19814 VGND.n6384 VGND.n6383 14.8179
R19815 VGND.n2569 VGND.n19 14.775
R19816 VGND.n5680 VGND.n5125 14.775
R19817 VGND.n5565 VGND.n5124 14.775
R19818 VGND.n1413 VGND.n1412 14.775
R19819 VGND.n8920 VGND.n8916 14.775
R19820 VGND.n240 VGND.n237 14.775
R19821 VGND.n1888 VGND.n1886 14.775
R19822 VGND.n7941 VGND.n7940 14.775
R19823 VGND.n4892 VGND.n4891 14.6829
R19824 VGND.n4685 VGND.n4163 14.6829
R19825 VGND.n1016 VGND.n1015 14.6829
R19826 VGND.n6455 VGND.n6454 14.6829
R19827 VGND.n9131 VGND.n9130 14.6829
R19828 VGND.n4946 VGND.n4945 14.6434
R19829 VGND.n8466 VGND.n8465 14.6388
R19830 VGND.n2557 VGND.n2556 14.3064
R19831 VGND.n7159 VGND.n1341 14.3064
R19832 VGND.n5026 VGND.n5025 14.3064
R19833 VGND.n4715 VGND.n4714 14.3064
R19834 VGND.n8625 VGND.n8624 14.3064
R19835 VGND.n6429 VGND.n6428 14.3064
R19836 VGND.n2937 VGND.n2936 14.3064
R19837 VGND.n2841 VGND.n2840 14.3064
R19838 VGND.n8497 VGND.n8496 14.3064
R19839 VGND.n948 VGND.n947 14.3064
R19840 VGND.n9142 VGND.n9141 14.3064
R19841 VGND.n5561 VGND.n5124 14.0717
R19842 VGND.n6336 VGND.n1688 14.0717
R19843 VGND.n2919 VGND.n2918 14.065
R19844 VGND.n5238 VGND.n5237 14.0503
R19845 VGND.n3046 VGND.n3035 13.9824
R19846 VGND.n1427 VGND.n1406 13.9299
R19847 VGND.n3923 VGND.n3887 13.8312
R19848 VGND.n8346 VGND.n8345 13.5534
R19849 VGND.n8021 VGND.n7951 13.5534
R19850 VGND.n1072 VGND.n1012 13.5534
R19851 VGND.n8901 VGND.n8900 13.48
R19852 VGND.n8574 VGND.n8573 13.3188
R19853 VGND.n5940 VGND.n1861 13.177
R19854 VGND.n6547 VGND.n6546 13.177
R19855 VGND.n5027 VGND.n5026 13.177
R19856 VGND.n2910 VGND.n2907 13.177
R19857 VGND.n2797 VGND.n2796 13.177
R19858 VGND.n2683 VGND.n2680 13.177
R19859 VGND.n351 VGND.n348 13.177
R19860 VGND.n1285 VGND.n1284 13.1375
R19861 VGND.n4461 VGND.n4458 13.0724
R19862 VGND.n1330 VGND.n1329 12.8005
R19863 VGND.n8459 VGND.n8457 12.8005
R19864 VGND.n8060 VGND.n479 12.8005
R19865 VGND.n1268 VGND.n1267 12.8005
R19866 VGND.n6857 VGND.n1589 12.8005
R19867 VGND.n6213 VGND.n1692 12.8005
R19868 VGND.n3794 VGND.n3777 12.5591
R19869 VGND.n8783 VGND.n8782 12.5161
R19870 VGND.n5019 VGND.n5018 12.424
R19871 VGND.n4113 VGND.n4111 12.424
R19872 VGND.n2865 VGND.n2864 12.424
R19873 VGND.n8054 VGND.n485 12.424
R19874 VGND.n1090 VGND.n1089 12.0894
R19875 VGND.n8310 VGND.n8309 12.0818
R19876 VGND.n3992 VGND.n3991 12.0476
R19877 VGND.n8784 VGND.n8783 12.0476
R19878 VGND.n7872 VGND.n7871 11.8129
R19879 VGND.n1216 VGND.n1163 11.7632
R19880 VGND.n2918 VGND.n2906 11.6711
R19881 VGND.n911 VGND.n910 11.5456
R19882 VGND.n25 VGND.n23 11.5456
R19883 VGND.n4948 VGND.n4947 11.2946
R19884 VGND.n4614 VGND.n4613 11.2946
R19885 VGND.n6408 VGND.n6407 11.2946
R19886 VGND.n4657 VGND.n4170 11.2016
R19887 VGND.n1428 VGND.n1427 10.9181
R19888 VGND.n3787 VGND.n3785 10.9181
R19889 VGND.n3319 VGND.n3318 10.9091
R19890 VGND.n4949 VGND.n4948 10.7135
R19891 VGND.n4436 VGND.n4435 10.7135
R19892 VGND.n2798 VGND.n2797 10.7135
R19893 VGND.n1954 VGND.n1922 10.7135
R19894 VGND.n1928 VGND.n1927 10.7135
R19895 VGND.n2459 VGND.n2342 10.5417
R19896 VGND.n4473 VGND.n4472 10.5417
R19897 VGND.n4638 VGND.n4554 10.5417
R19898 VGND.n2661 VGND.n2660 10.5417
R19899 VGND.n2660 VGND.n2659 10.4353
R19900 VGND.n4615 VGND.n4614 10.307
R19901 VGND.n2827 VGND.n2825 10.2756
R19902 VGND.n2467 VGND.n2464 10.1652
R19903 VGND.n5053 VGND.n4039 10.1652
R19904 VGND.n4449 VGND.n4446 10.0005
R19905 VGND.n8634 VGND.n217 9.78874
R19906 VGND.n7885 VGND.n7883 9.78874
R19907 VGND.n957 VGND.n956 9.78874
R19908 VGND.n1024 VGND.n1023 9.78874
R19909 VGND.n6440 VGND.n6437 9.78874
R19910 VGND.n1903 VGND.n1877 9.53804
R19911 VGND.n8534 VGND.n8533 9.41937
R19912 VGND.n4441 VGND.n4439 9.41227
R19913 VGND.n3785 VGND.n3778 9.41227
R19914 VGND.n6349 VGND.n6347 9.41227
R19915 VGND.n4247 VGND.n4245 9.40819
R19916 VGND.n385 VGND.n384 9.37278
R19917 VGND.n2446 VGND.n2445 9.36527
R19918 VGND.n8739 VGND.n177 9.32922
R19919 VGND.n7104 VGND.n7103 9.3005
R19920 VGND.n7107 VGND.n7106 9.3005
R19921 VGND.n7196 VGND.n7195 9.3005
R19922 VGND.n7198 VGND.n7197 9.3005
R19923 VGND.n7207 VGND.n7206 9.3005
R19924 VGND.n7209 VGND.n7208 9.3005
R19925 VGND.n4008 VGND.n4007 9.3005
R19926 VGND.n4006 VGND.n4005 9.3005
R19927 VGND.n4980 VGND.n4979 9.3005
R19928 VGND.n4850 VGND.n4849 9.3005
R19929 VGND.n4853 VGND.n4852 9.3005
R19930 VGND.n4797 VGND.n4796 9.3005
R19931 VGND.n4795 VGND.n4794 9.3005
R19932 VGND.n4521 VGND.n4520 9.3005
R19933 VGND.n4322 VGND.n4321 9.3005
R19934 VGND.n4500 VGND.n4499 9.3005
R19935 VGND.n4498 VGND.n4497 9.3005
R19936 VGND.n4212 VGND.n4211 9.3005
R19937 VGND.n4519 VGND.n4518 9.3005
R19938 VGND.n4334 VGND.n4333 9.3005
R19939 VGND.n4332 VGND.n4331 9.3005
R19940 VGND.n4320 VGND.n4319 9.3005
R19941 VGND.n4726 VGND.n4725 9.3005
R19942 VGND.n4724 VGND.n4723 9.3005
R19943 VGND.n4127 VGND.n4126 9.3005
R19944 VGND.n4125 VGND.n4124 9.3005
R19945 VGND.n3370 VGND.n3369 9.3005
R19946 VGND.n3360 VGND.n3359 9.3005
R19947 VGND.n3368 VGND.n3367 9.3005
R19948 VGND.n3228 VGND.n3227 9.3005
R19949 VGND.n2782 VGND.n2781 9.3005
R19950 VGND.n3226 VGND.n3225 9.3005
R19951 VGND.n2780 VGND.n2779 9.3005
R19952 VGND.n2076 VGND.n2075 9.3005
R19953 VGND.n2074 VGND.n2073 9.3005
R19954 VGND.n8848 VGND.n8847 9.3005
R19955 VGND.n8846 VGND.n8845 9.3005
R19956 VGND.n8838 VGND.n8837 9.3005
R19957 VGND.n9027 VGND.n9026 9.3005
R19958 VGND.n3040 VGND.n3037 9.3005
R19959 VGND.n9029 VGND.n9028 9.3005
R19960 VGND.n3039 VGND.n3038 9.3005
R19961 VGND.n3167 VGND.n3166 9.3005
R19962 VGND.n3170 VGND.n3169 9.3005
R19963 VGND.n9022 VGND.n9021 9.3005
R19964 VGND.n9020 VGND.n9019 9.3005
R19965 VGND.n3905 VGND.n3904 9.3005
R19966 VGND.n8660 VGND.n8659 9.3005
R19967 VGND.n8662 VGND.n8661 9.3005
R19968 VGND.n8566 VGND.n8565 9.3005
R19969 VGND.n8568 VGND.n8567 9.3005
R19970 VGND.n8655 VGND.n8654 9.3005
R19971 VGND.n8653 VGND.n8652 9.3005
R19972 VGND.n3907 VGND.n3906 9.3005
R19973 VGND.n3829 VGND.n3828 9.3005
R19974 VGND.n3831 VGND.n3830 9.3005
R19975 VGND.n3808 VGND.n3807 9.3005
R19976 VGND.n3803 VGND.n3802 9.3005
R19977 VGND.n7818 VGND.n506 9.3005
R19978 VGND.n7743 VGND.n7742 9.3005
R19979 VGND.n8076 VGND.n8075 9.3005
R19980 VGND.n8067 VGND.n8066 9.3005
R19981 VGND.n8074 VGND.n8073 9.3005
R19982 VGND.n7917 VGND.n7916 9.3005
R19983 VGND.n8065 VGND.n8064 9.3005
R19984 VGND.n1914 VGND.n1913 9.3005
R19985 VGND.n1910 VGND.n1909 9.3005
R19986 VGND.n8189 VGND.n8188 9.3005
R19987 VGND.n681 VGND.n680 9.3005
R19988 VGND.n7550 VGND.n7549 9.3005
R19989 VGND.n7622 VGND.n7621 9.3005
R19990 VGND.n7688 VGND.n7687 9.3005
R19991 VGND.n8136 VGND.n8135 9.3005
R19992 VGND.n439 VGND.n438 9.3005
R19993 VGND.n437 VGND.n436 9.3005
R19994 VGND.n8191 VGND.n8190 9.3005
R19995 VGND.n7620 VGND.n7619 9.3005
R19996 VGND.n7611 VGND.n7610 9.3005
R19997 VGND.n7552 VGND.n7551 9.3005
R19998 VGND.n8131 VGND.n8130 9.3005
R19999 VGND.n8205 VGND.n8204 9.3005
R20000 VGND.n719 VGND.n718 9.3005
R20001 VGND.n717 VGND.n716 9.3005
R20002 VGND.n7316 VGND.n7315 9.3005
R20003 VGND.n1129 VGND.n1128 9.3005
R20004 VGND.n1193 VGND.n1192 9.3005
R20005 VGND.n1190 VGND.n1189 9.3005
R20006 VGND.n1301 VGND.n1300 9.3005
R20007 VGND.n1019 VGND.n1018 9.3005
R20008 VGND.n876 VGND.n875 9.3005
R20009 VGND.n874 VGND.n873 9.3005
R20010 VGND.n7439 VGND.n7438 9.3005
R20011 VGND.n7437 VGND.n7436 9.3005
R20012 VGND.n7487 VGND.n7486 9.3005
R20013 VGND.n7485 VGND.n7484 9.3005
R20014 VGND.n6798 VGND.n6797 9.3005
R20015 VGND.n6800 VGND.n6799 9.3005
R20016 VGND.n6805 VGND.n6804 9.3005
R20017 VGND.n6936 VGND.n6935 9.3005
R20018 VGND.n6938 VGND.n6937 9.3005
R20019 VGND.n6825 VGND.n1591 9.3005
R20020 VGND.n6824 VGND.n6823 9.3005
R20021 VGND.n6807 VGND.n6806 9.3005
R20022 VGND.n6180 VGND.n6179 9.3005
R20023 VGND.n6182 VGND.n6181 9.3005
R20024 VGND.n6149 VGND.n6148 9.3005
R20025 VGND.n6147 VGND.n6146 9.3005
R20026 VGND.n6632 VGND.n6631 9.3005
R20027 VGND.n5350 VGND.n5349 9.3005
R20028 VGND.n5372 VGND.n5371 9.3005
R20029 VGND.n6722 VGND.n6721 9.3005
R20030 VGND.n6634 VGND.n1634 9.3005
R20031 VGND.n6550 VGND.n6549 9.3005
R20032 VGND.n6552 VGND.n6551 9.3005
R20033 VGND.n6560 VGND.n6559 9.3005
R20034 VGND.n6562 VGND.n6561 9.3005
R20035 VGND.n6065 VGND.n6064 9.3005
R20036 VGND.n6063 VGND.n6062 9.3005
R20037 VGND.n1743 VGND.n1742 9.3005
R20038 VGND.n1741 VGND.n1740 9.3005
R20039 VGND.n5879 VGND.n5878 9.3005
R20040 VGND.n5596 VGND.n5595 9.3005
R20041 VGND.n5757 VGND.n5756 9.3005
R20042 VGND.n5759 VGND.n5758 9.3005
R20043 VGND.n5645 VGND.n5644 9.3005
R20044 VGND.n5643 VGND.n5642 9.3005
R20045 VGND.n5592 VGND.n5591 9.3005
R20046 VGND.n5601 VGND.n5600 9.3005
R20047 VGND.n5881 VGND.n5880 9.3005
R20048 VGND.n5869 VGND.n5868 9.3005
R20049 VGND.n5871 VGND.n5870 9.3005
R20050 VGND.n5994 VGND.n5993 9.3005
R20051 VGND.n5992 VGND.n5991 9.3005
R20052 VGND.n1829 VGND.n1828 9.3005
R20053 VGND.n1827 VGND.n1826 9.3005
R20054 VGND.n2487 VGND.n2486 9.3005
R20055 VGND.n2255 VGND.n2254 9.3005
R20056 VGND.n2265 VGND.n2264 9.3005
R20057 VGND.n2257 VGND.n2256 9.3005
R20058 VGND.n2498 VGND.n2497 9.3005
R20059 VGND.n2492 VGND.n2491 9.3005
R20060 VGND.n2389 VGND.n2388 9.3005
R20061 VGND.n2386 VGND.n2385 9.3005
R20062 VGND.n2500 VGND.n2499 9.3005
R20063 VGND.n2316 VGND.n2315 9.3005
R20064 VGND.n3513 VGND.n3512 9.3005
R20065 VGND.n3511 VGND.n3510 9.3005
R20066 VGND.n1770 VGND.n1769 9.03579
R20067 VGND.n1650 VGND.n1649 9.03579
R20068 VGND.n4947 VGND.n4946 9.03579
R20069 VGND.n4910 VGND.n4909 9.03579
R20070 VGND.n4393 VGND.n4392 9.03579
R20071 VGND.n7071 VGND.n7070 9.02922
R20072 VGND.n8526 VGND.n8525 9.02922
R20073 VGND.n405 VGND.n404 9.02922
R20074 VGND.n5286 VGND.n5285 9.02922
R20075 VGND.n4800 VGND.n4799 9.0005
R20076 VGND.n4847 VGND.n4846 9.0005
R20077 VGND.n4855 VGND.n4854 9.0005
R20078 VGND.n4011 VGND.n4010 9.0005
R20079 VGND.n7109 VGND.n7108 9.0005
R20080 VGND.n7102 VGND.n7101 9.0005
R20081 VGND.n7202 VGND.n7201 9.0005
R20082 VGND.n7211 VGND.n7210 9.0005
R20083 VGND.n4991 VGND.n4986 9.0005
R20084 VGND.n4517 VGND.n4516 9.0005
R20085 VGND.n4480 VGND.n4479 9.0005
R20086 VGND.n4130 VGND.n4129 9.0005
R20087 VGND.n4159 VGND.n4146 9.0005
R20088 VGND.n4729 VGND.n4728 9.0005
R20089 VGND.n4722 VGND.n4721 9.0005
R20090 VGND.n4502 VGND.n4501 9.0005
R20091 VGND.n1463 VGND.n1462 9.0005
R20092 VGND.n4576 VGND.n4575 9.0005
R20093 VGND.n4358 VGND.n4357 9.0005
R20094 VGND.n4340 VGND.n4335 9.0005
R20095 VGND.n4308 VGND.n4307 9.0005
R20096 VGND.n4324 VGND 9.0005
R20097 VGND VGND.n4323 9.0005
R20098 VGND.n2079 VGND.n2078 9.0005
R20099 VGND.n52 VGND.n51 9.0005
R20100 VGND.n2778 VGND.n2777 9.0005
R20101 VGND.n2990 VGND.n2989 9.0005
R20102 VGND.n2980 VGND.n2979 9.0005
R20103 VGND.n3233 VGND.n3232 9.0005
R20104 VGND.n3366 VGND.n3365 9.0005
R20105 VGND.n3372 VGND.n3371 9.0005
R20106 VGND.n3357 VGND.n2125 9.0005
R20107 VGND.n9018 VGND.n9017 9.0005
R20108 VGND.n9031 VGND.n9030 9.0005
R20109 VGND.n76 VGND.n75 9.0005
R20110 VGND.n3172 VGND.n3171 9.0005
R20111 VGND.n3165 VGND.n3164 9.0005
R20112 VGND.n8850 VGND.n8849 9.0005
R20113 VGND.n8844 VGND.n8843 9.0005
R20114 VGND.n8835 VGND.n101 9.0005
R20115 VGND.n196 VGND.n195 9.0005
R20116 VGND.n3811 VGND.n3810 9.0005
R20117 VGND.n3826 VGND.n3825 9.0005
R20118 VGND.n3833 VGND.n3832 9.0005
R20119 VGND.n8664 VGND.n8663 9.0005
R20120 VGND.n8570 VGND.n8569 9.0005
R20121 VGND.n8564 VGND.n8563 9.0005
R20122 VGND.n3909 VGND.n3908 9.0005
R20123 VGND.n3903 VGND.n3902 9.0005
R20124 VGND.n7920 VGND.n7919 9.0005
R20125 VGND.n1917 VGND.n1916 9.0005
R20126 VGND.n8078 VGND.n8077 9.0005
R20127 VGND.n8070 VGND.n8069 9.0005
R20128 VGND.n7815 VGND.n7814 9.0005
R20129 VGND.n7749 VGND.n7748 9.0005
R20130 VGND.n7739 VGND.n539 9.0005
R20131 VGND.n8311 VGND.n8310 9.0005
R20132 VGND.n8192 VGND.n8154 9.0005
R20133 VGND.n8133 VGND.n8132 9.0005
R20134 VGND.n435 VGND.n434 9.0005
R20135 VGND.n7547 VGND.n7546 9.0005
R20136 VGND.n7554 VGND.n7553 9.0005
R20137 VGND.n8203 VGND.n8202 9.0005
R20138 VGND.n7690 VGND.n7689 9.0005
R20139 VGND.n7624 VGND.n7623 9.0005
R20140 VGND.n7618 VGND.n7617 9.0005
R20141 VGND.n7705 VGND.n602 9.0005
R20142 VGND.n7490 VGND.n7489 9.0005
R20143 VGND.n7442 VGND.n7441 9.0005
R20144 VGND.n7434 VGND.n7433 9.0005
R20145 VGND.n1196 VGND.n1195 9.0005
R20146 VGND.n1133 VGND.n1132 9.0005
R20147 VGND.n1188 VGND.n1187 9.0005
R20148 VGND.n7333 VGND.n7332 9.0005
R20149 VGND.n879 VGND.n877 9.0005
R20150 VGND.n7320 VGND.n7319 9.0005
R20151 VGND.n6795 VGND.n6794 9.0005
R20152 VGND.n6152 VGND.n6151 9.0005
R20153 VGND.n6114 VGND.n6100 9.0005
R20154 VGND.n6177 VGND.n6176 9.0005
R20155 VGND.n6184 VGND.n6183 9.0005
R20156 VGND.n6822 VGND.n6821 9.0005
R20157 VGND.n6933 VGND.n6932 9.0005
R20158 VGND.n6963 VGND.n6962 9.0005
R20159 VGND.n6940 VGND.n6939 9.0005
R20160 VGND.n6809 VGND.n6808 9.0005
R20161 VGND.n1745 VGND.n1744 9.0005
R20162 VGND.n6068 VGND.n6067 9.0005
R20163 VGND.n6061 VGND.n6060 9.0005
R20164 VGND.n6548 VGND.n6547 9.0005
R20165 VGND.n6726 VGND.n6725 9.0005
R20166 VGND.n1636 VGND.n1635 9.0005
R20167 VGND.n6566 VGND.n6565 9.0005
R20168 VGND.n6558 VGND.n6557 9.0005
R20169 VGND.n1832 VGND.n1831 9.0005
R20170 VGND.n5997 VGND.n5996 9.0005
R20171 VGND.n5990 VGND.n5989 9.0005
R20172 VGND.n5605 VGND.n5604 9.0005
R20173 VGND.n5641 VGND.n5640 9.0005
R20174 VGND.n5754 VGND.n5753 9.0005
R20175 VGND.n5761 VGND.n5760 9.0005
R20176 VGND.n5590 VGND.n5589 9.0005
R20177 VGND.n5883 VGND.n5882 9.0005
R20178 VGND.n5877 VGND.n5876 9.0005
R20179 VGND.n5867 VGND.n5866 9.0005
R20180 VGND.n2391 VGND.n2390 9.0005
R20181 VGND.n2493 VGND.n2336 9.0005
R20182 VGND.n2318 VGND.n2313 9.0005
R20183 VGND.n3516 VGND.n3515 9.0005
R20184 VGND.n2259 VGND.n2258 9.0005
R20185 VGND.n2253 VGND.n2252 9.0005
R20186 VGND.n2277 VGND.n2276 9.0005
R20187 VGND.n2502 VGND.n2501 9.0005
R20188 VGND.n2384 VGND.n2383 9.0005
R20189 VGND.n4784 VGND.n4765 8.65932
R20190 VGND.n8348 VGND.n8347 8.65932
R20191 VGND.n1582 VGND.n1581 8.65932
R20192 VGND.t1593 VGND.t430 8.42962
R20193 VGND.t320 VGND.t289 8.42962
R20194 VGND VGND.t751 8.42962
R20195 VGND.t572 VGND.t467 8.42962
R20196 VGND.t1793 VGND.t2730 8.42962
R20197 VGND.t1749 VGND.t2728 8.42962
R20198 VGND VGND.t2364 8.42962
R20199 VGND.t486 VGND.t3047 8.42962
R20200 VGND.t76 VGND.t2343 8.42962
R20201 VGND.t2087 VGND.t2654 8.42962
R20202 VGND.t2062 VGND.t2652 8.42962
R20203 VGND.t3045 VGND.t2466 8.42962
R20204 VGND.n6647 VGND.n6646 8.28285
R20205 VGND.n5031 VGND.n5030 8.28285
R20206 VGND.n3946 VGND.n3945 8.28285
R20207 VGND.n2592 VGND.n2591 8.23546
R20208 VGND.n2228 VGND.n2225 8.23546
R20209 VGND.n5255 VGND.n5254 8.23546
R20210 VGND.n6683 VGND.n6682 8.23546
R20211 VGND.n6687 VGND.n1629 8.23546
R20212 VGND.n4529 VGND.n4525 8.23546
R20213 VGND.n4537 VGND.n4172 8.23546
R20214 VGND.n4538 VGND.n4537 8.23546
R20215 VGND.n4541 VGND.n4540 8.23546
R20216 VGND.n2065 VGND.n2043 8.23546
R20217 VGND.n2068 VGND.n2065 8.23546
R20218 VGND.n3427 VGND.n2108 8.23546
R20219 VGND.n3085 VGND.n3084 8.23546
R20220 VGND.n3072 VGND.n3069 8.23546
R20221 VGND.n3056 VGND.n3034 8.23546
R20222 VGND.n8882 VGND.n92 8.23546
R20223 VGND.n3855 VGND.n3853 8.23546
R20224 VGND.n3855 VGND.n3854 8.23546
R20225 VGND.n8735 VGND.n8734 8.23546
R20226 VGND.n8720 VGND.n194 8.23546
R20227 VGND.n7783 VGND.n7782 8.23546
R20228 VGND.n7826 VGND.n7823 8.23546
R20229 VGND.n7576 VGND.n7575 8.23546
R20230 VGND.n7683 VGND.n683 8.23546
R20231 VGND.n7683 VGND.n684 8.23546
R20232 VGND.n8177 VGND.n8176 8.23546
R20233 VGND.n8176 VGND.n8158 8.23546
R20234 VGND.n8172 VGND.n8158 8.23546
R20235 VGND.n1290 VGND.n1147 8.23546
R20236 VGND.n1148 VGND.n1147 8.23546
R20237 VGND.n1004 VGND.n1003 8.23546
R20238 VGND.n1118 VGND.n1004 8.23546
R20239 VGND.n7409 VGND.n7408 8.23546
R20240 VGND.n7393 VGND.n807 8.23546
R20241 VGND.n7386 VGND.n807 8.23546
R20242 VGND.n1498 VGND.n1488 8.23546
R20243 VGND.n6833 VGND.n6832 8.23546
R20244 VGND.n6674 VGND.n1631 8.16157
R20245 VGND.n2490 VGND.n2489 8.10717
R20246 VGND.n231 VGND.n230 8.10717
R20247 VGND.n444 VGND.n443 8.10717
R20248 VGND.n6236 VGND.n6235 8.10717
R20249 VGND.n2586 VGND.n2585 8.05644
R20250 VGND.n9183 VGND.n17 8.05644
R20251 VGND.n6677 VGND.n6676 8.05644
R20252 VGND.n2067 VGND.n2066 8.05644
R20253 VGND.n3084 VGND.n3030 8.05644
R20254 VGND.n86 VGND.n85 8.05644
R20255 VGND.n7783 VGND.n522 8.05644
R20256 VGND.n531 VGND.n530 8.05644
R20257 VGND.n7667 VGND.n7666 8.05644
R20258 VGND.n9151 VGND.n9150 8.0482
R20259 VGND.n7825 VGND.n7824 7.96693
R20260 VGND.n2679 VGND.n2677 7.90638
R20261 VGND.n3777 VGND.n3775 7.90638
R20262 VGND.n347 VGND.n345 7.90638
R20263 VGND.n5257 VGND.n5256 7.87742
R20264 VGND.n5442 VGND.n5197 7.87742
R20265 VGND.n5378 VGND.n5377 7.87742
R20266 VGND.n6676 VGND.n1630 7.87742
R20267 VGND.n7060 VGND.n7005 7.87742
R20268 VGND.n2066 VGND.n2041 7.87742
R20269 VGND.n2618 VGND.n2617 7.6984
R20270 VGND.n2193 VGND.n2180 7.6984
R20271 VGND.n5469 VGND.n5468 7.6984
R20272 VGND.n5504 VGND.n5503 7.6984
R20273 VGND.n5111 VGND.n5110 7.6984
R20274 VGND.n1859 VGND.n1858 7.6984
R20275 VGND.n5257 VGND.n5228 7.6984
R20276 VGND.n7010 VGND.n7009 7.6984
R20277 VGND.n4082 VGND.n4081 7.6984
R20278 VGND.n4525 VGND.n4173 7.6984
R20279 VGND.n4529 VGND.n4528 7.6984
R20280 VGND.n3027 VGND.n3026 7.6984
R20281 VGND.n3070 VGND.n3031 7.6984
R20282 VGND.n3848 VGND.n3847 7.6984
R20283 VGND.n7580 VGND.n686 7.6984
R20284 VGND.n7586 VGND.n7585 7.6984
R20285 VGND.n7604 VGND.n7603 7.6984
R20286 VGND.n441 VGND.n440 7.6984
R20287 VGND.n1149 VGND.n1148 7.6984
R20288 VGND.n809 VGND.n808 7.6984
R20289 VGND.n7409 VGND.n805 7.6984
R20290 VGND.n7387 VGND.n7386 7.6984
R20291 VGND.n6863 VGND.n6862 7.6984
R20292 VGND.n6257 VGND.n6256 7.6984
R20293 VGND.n2869 VGND.n2868 7.6805
R20294 VGND.n2292 VGND.n2291 7.60889
R20295 VGND.n2183 VGND.n2182 7.60889
R20296 VGND.n4547 VGND.n4546 7.60889
R20297 VGND.n2073 VGND.n2072 7.60889
R20298 VGND.n3051 VGND.n3050 7.60889
R20299 VGND.n518 VGND.n517 7.6005
R20300 VGND.n1435 VGND.n1394 7.56414
R20301 VGND.n8585 VGND.n243 7.56414
R20302 VGND.n1524 VGND.n1479 7.56414
R20303 VGND.n6648 VGND.n6647 7.52991
R20304 VGND.n1946 VGND.n1945 7.52991
R20305 VGND.n1254 VGND.n1156 7.52991
R20306 VGND.n6408 VGND.n6405 7.52991
R20307 VGND.n5206 VGND.n5204 7.50395
R20308 VGND.n8981 VGND.n8979 7.3908
R20309 VGND.n7536 VGND.n7535 7.34036
R20310 VGND.n6234 VGND.n6233 7.23528
R20311 VGND.n4447 VGND.n4169 7.15344
R20312 VGND.n8774 VGND.n8773 7.15344
R20313 VGND.n483 VGND.n482 7.15344
R20314 VGND.n1032 VGND.n1031 7.15344
R20315 VGND.n6905 VGND.n6904 7.15344
R20316 VGND.n2617 VGND.n2616 7.15139
R20317 VGND.n1120 VGND.n1118 7.15139
R20318 VGND.n2225 VGND.n2172 7.11268
R20319 VGND.n5445 VGND.n5441 7.11268
R20320 VGND.n6597 VGND.n6596 7.11268
R20321 VGND.n3289 VGND.n3288 7.11268
R20322 VGND.n8721 VGND.n8720 7.11268
R20323 VGND.n1499 VGND.n1498 7.11268
R20324 VGND.n8893 VGND.n8892 6.90655
R20325 VGND.n8887 VGND.n87 6.90655
R20326 VGND.n7762 VGND.n7761 6.90655
R20327 VGND.n7821 VGND.n506 6.89281
R20328 VGND.n2585 VGND.n2297 6.88949
R20329 VGND.n2195 VGND.n2193 6.88949
R20330 VGND.n5254 VGND.n5232 6.88949
R20331 VGND.n7061 VGND.n7060 6.88949
R20332 VGND.n3058 VGND.n3056 6.88949
R20333 VGND.n8734 VGND.n184 6.88949
R20334 VGND.n7782 VGND.n524 6.88949
R20335 VGND.n394 VGND.n393 6.88949
R20336 VGND.n3932 VGND.n3929 6.77697
R20337 VGND.n7832 VGND.n504 6.77697
R20338 VGND.n6285 VGND.n6262 6.77697
R20339 VGND.n3071 VGND.n3070 6.62428
R20340 VGND.n6704 VGND.n1620 6.61527
R20341 VGND.n5453 VGND.n5452 6.57117
R20342 VGND.n6701 VGND.n1620 6.57117
R20343 VGND.n6701 VGND.n6700 6.57117
R20344 VGND.n3420 VGND.n2110 6.57117
R20345 VGND.n8880 VGND.n93 6.57117
R20346 VGND.n6236 VGND.n1691 6.57117
R20347 VGND.n2350 VGND.n2349 6.44526
R20348 VGND.n4235 VGND.n4234 6.44526
R20349 VGND.n180 VGND.n179 6.44345
R20350 VGND.n6029 VGND.n6028 6.4005
R20351 VGND.n3282 VGND.n2659 6.4005
R20352 VGND.n8598 VGND.n236 6.4005
R20353 VGND.n6286 VGND.n6285 6.4005
R20354 VGND.n8925 VGND.n80 6.26433
R20355 VGND.n8779 VGND.n8778 6.26433
R20356 VGND.n675 VGND.n674 6.26433
R20357 VGND.n971 VGND.n970 6.26433
R20358 VGND.n7427 VGND.n7426 6.26433
R20359 VGND.n7426 VGND.n793 6.26433
R20360 VGND.n6241 VGND.n6239 6.26433
R20361 VGND.n8386 VGND.n8385 6.19624
R20362 VGND.n5399 VGND.n5340 6.15761
R20363 VGND.n2405 VGND.n2357 6.14752
R20364 VGND.n8741 VGND.n176 6.12816
R20365 VGND.n8902 VGND.n8901 6.06366
R20366 VGND.n3394 VGND.n3393 6.02861
R20367 VGND.n3654 VGND.n3653 6.02861
R20368 VGND.n2214 VGND.n2212 6.0286
R20369 VGND.n8484 VGND.n8456 6.02403
R20370 VGND.n648 VGND.n647 6.02403
R20371 VGND.n634 VGND.n633 6.02403
R20372 VGND.n1161 VGND.n1160 6.02403
R20373 VGND.n1229 VGND.n1228 6.02403
R20374 VGND.n6414 VGND.n6413 6.02403
R20375 VGND.n6400 VGND.n6399 6.02403
R20376 VGND.n2962 VGND.n2898 5.99199
R20377 VGND.n2476 VGND.n2339 5.98311
R20378 VGND.n5134 VGND.n5133 5.98311
R20379 VGND.n1802 VGND.n1801 5.98311
R20380 VGND.n6625 VGND.n1638 5.98311
R20381 VGND.n5062 VGND.n5061 5.98311
R20382 VGND.n5049 VGND.n5045 5.98311
R20383 VGND.n4453 VGND.n4450 5.98311
R20384 VGND.n4654 VGND.n4552 5.98311
R20385 VGND.n3798 VGND.n3795 5.98311
R20386 VGND.n1899 VGND.n1898 5.98311
R20387 VGND.n8157 VGND.n8156 5.90819
R20388 VGND.n1629 VGND.n1628 5.8885
R20389 VGND.n5154 VGND.n5153 5.85582
R20390 VGND.n5679 VGND.n5678 5.85582
R20391 VGND.n1733 VGND.n1732 5.85582
R20392 VGND.n4161 VGND.n4160 5.85582
R20393 VGND.n4166 VGND.n4165 5.85582
R20394 VGND.n4424 VGND.n4423 5.85582
R20395 VGND.n1393 VGND.n1392 5.85582
R20396 VGND.n2963 VGND.n2962 5.85582
R20397 VGND.n2829 VGND.n2828 5.85582
R20398 VGND.n2694 VGND.n2693 5.85582
R20399 VGND.n8919 VGND.n8918 5.85582
R20400 VGND.n8474 VGND.n8460 5.85582
R20401 VGND.n8454 VGND.n8453 5.85582
R20402 VGND.n3881 VGND.n3880 5.85582
R20403 VGND.n8779 VGND.n162 5.85582
R20404 VGND.n171 VGND.n170 5.85582
R20405 VGND.n8741 VGND.n8740 5.85582
R20406 VGND.n8387 VGND.n8381 5.85582
R20407 VGND.n1892 VGND.n1889 5.85582
R20408 VGND.n342 VGND.n341 5.85582
R20409 VGND.n705 VGND.n704 5.85582
R20410 VGND.n675 VGND.n673 5.85582
R20411 VGND.n447 VGND.n446 5.85582
R20412 VGND.n1478 VGND.n1477 5.85582
R20413 VGND.n6226 VGND.n6225 5.85582
R20414 VGND.n1647 VGND.n1646 5.81868
R20415 VGND.n2202 VGND.n2200 5.80542
R20416 VGND.n5429 VGND.n5427 5.80542
R20417 VGND.n3416 VGND.n3415 5.80542
R20418 VGND.n8872 VGND.n8871 5.80542
R20419 VGND.n1422 VGND.n1421 5.78773
R20420 VGND.n8473 VGND.n8472 5.78773
R20421 VGND.n7844 VGND.n7843 5.70485
R20422 VGND.n2729 VGND.n2728 5.65809
R20423 VGND.n8934 VGND.n8925 5.65809
R20424 VGND.n6241 VGND.n6240 5.65809
R20425 VGND.n1031 VGND.n1030 5.64756
R20426 VGND.n2592 VGND.n2289 5.63966
R20427 VGND.n5450 VGND.n5449 5.63966
R20428 VGND.n5378 VGND.n5375 5.63966
R20429 VGND.n6678 VGND.n6675 5.63966
R20430 VGND.n2109 VGND.n2108 5.63966
R20431 VGND.n3284 VGND.n3283 5.63966
R20432 VGND.n8898 VGND.n8896 5.63966
R20433 VGND.n8882 VGND.n8881 5.63966
R20434 VGND.n8735 VGND.n182 5.63966
R20435 VGND.n7667 VGND.n7601 5.63966
R20436 VGND.n6853 VGND.n6852 5.63966
R20437 VGND.n8907 VGND.n83 5.5878
R20438 VGND.n793 VGND.n792 5.57042
R20439 VGND.n6696 VGND.n6695 5.53969
R20440 VGND.n3311 VGND.n3306 5.48128
R20441 VGND.n8267 VGND.n8266 5.35702
R20442 VGND.n7139 VGND.n1348 5.27109
R20443 VGND.n4381 VGND.n4168 5.27109
R20444 VGND.n3946 VGND.n3943 5.27109
R20445 VGND.n1067 VGND.n1066 5.27109
R20446 VGND.n811 VGND.n810 5.27109
R20447 VGND.n1623 VGND.n1622 5.13241
R20448 VGND.n3488 VGND.n3485 5.13108
R20449 VGND.n3488 VGND.n3487 5.13108
R20450 VGND.n9 VGND.n7 5.13108
R20451 VGND.n5237 VGND.n5234 5.13108
R20452 VGND.n5237 VGND.n5236 5.13108
R20453 VGND.n1714 VGND.n1711 5.13108
R20454 VGND.n1714 VGND.n1713 5.13108
R20455 VGND.n7015 VGND.n7012 5.13108
R20456 VGND.n7015 VGND.n7014 5.13108
R20457 VGND.n4769 VGND.n4767 5.13108
R20458 VGND.n4769 VGND.n4768 5.13108
R20459 VGND.n1412 VGND.n1409 5.13108
R20460 VGND.n1412 VGND.n1411 5.13108
R20461 VGND.n4101 VGND.n4099 5.13108
R20462 VGND.n4101 VGND.n4100 5.13108
R20463 VGND.n2910 VGND.n2908 5.13108
R20464 VGND.n2910 VGND.n2909 5.13108
R20465 VGND.n2051 VGND.n2048 5.13108
R20466 VGND.n2051 VGND.n2050 5.13108
R20467 VGND.n2683 VGND.n2681 5.13108
R20468 VGND.n2683 VGND.n2682 5.13108
R20469 VGND.n3673 VGND.n3670 5.13108
R20470 VGND.n3673 VGND.n3672 5.13108
R20471 VGND.n8916 VGND.n8915 5.13108
R20472 VGND.n8465 VGND.n8462 5.13108
R20473 VGND.n8465 VGND.n8464 5.13108
R20474 VGND.n3781 VGND.n3779 5.13108
R20475 VGND.n3781 VGND.n3780 5.13108
R20476 VGND.n8356 VGND.n8353 5.13108
R20477 VGND.n8356 VGND.n8355 5.13108
R20478 VGND.n1886 VGND.n1884 5.13108
R20479 VGND.n1886 VGND.n1885 5.13108
R20480 VGND.n351 VGND.n349 5.13108
R20481 VGND.n351 VGND.n350 5.13108
R20482 VGND.n694 VGND.n692 5.13108
R20483 VGND.n694 VGND.n693 5.13108
R20484 VGND.n931 VGND.n929 5.13108
R20485 VGND.n931 VGND.n930 5.13108
R20486 VGND.n7462 VGND.n7459 5.13108
R20487 VGND.n7462 VGND.n7461 5.13108
R20488 VGND.n1493 VGND.n1490 5.13108
R20489 VGND.n1493 VGND.n1492 5.13108
R20490 VGND.n1589 VGND.n1588 5.13108
R20491 VGND.n6120 VGND.n6117 5.13108
R20492 VGND.n6120 VGND.n6119 5.13108
R20493 VGND.n9121 VGND.n9119 5.13108
R20494 VGND.n9121 VGND.n9120 5.13108
R20495 VGND VGND.n1804 5.09003
R20496 VGND.n5137 VGND.n5136 5.06789
R20497 VGND.n1485 VGND.n1484 5.04614
R20498 VGND.n358 VGND.n357 5.03644
R20499 VGND.n1396 VGND.n1395 5.02529
R20500 VGND.n245 VGND.n244 5.02529
R20501 VGND.n1481 VGND.n1480 5.02529
R20502 VGND.n8644 VGND.n8643 4.93346
R20503 VGND.n3979 VGND.n3978 4.89462
R20504 VGND.n9157 VGND.n9156 4.85762
R20505 VGND.n2299 VGND.n2298 4.85762
R20506 VGND.n5556 VGND.n5555 4.85762
R20507 VGND.n5654 VGND.n5653 4.85762
R20508 VGND.n5691 VGND.n5690 4.85762
R20509 VGND.n4596 VGND.n4595 4.85762
R20510 VGND.n4560 VGND.n4559 4.85762
R20511 VGND.n2951 VGND.n2950 4.85762
R20512 VGND.n2754 VGND.n2753 4.85762
R20513 VGND.n3217 VGND.n3216 4.85762
R20514 VGND.n3301 VGND.n3300 4.85762
R20515 VGND.n2723 VGND.n2722 4.85762
R20516 VGND.n8929 VGND.n8928 4.85762
R20517 VGND.n250 VGND.n249 4.85762
R20518 VGND.n8511 VGND.n8510 4.85762
R20519 VGND.n3964 VGND.n3963 4.85762
R20520 VGND.n210 VGND.n209 4.85762
R20521 VGND.n8602 VGND.n8601 4.85762
R20522 VGND.n7896 VGND.n7895 4.85762
R20523 VGND.n7862 VGND.n7861 4.85762
R20524 VGND.n512 VGND.n511 4.85762
R20525 VGND.n364 VGND.n363 4.85762
R20526 VGND.n8227 VGND.n8226 4.85762
R20527 VGND.n964 VGND.n963 4.85762
R20528 VGND.n7419 VGND.n7418 4.85762
R20529 VGND.n1009 VGND.n1008 4.85762
R20530 VGND.n6247 VGND.n6246 4.85762
R20531 VGND.n6620 VGND.n6619 4.85567
R20532 VGND.n2476 VGND.n2475 4.8005
R20533 VGND.n5739 VGND.n5738 4.8005
R20534 VGND.n1803 VGND.n1802 4.8005
R20535 VGND.n1709 VGND.n1708 4.8005
R20536 VGND.n1345 VGND.n1344 4.8005
R20537 VGND.n5049 VGND.n5048 4.8005
R20538 VGND.n4238 VGND.n4237 4.8005
R20539 VGND.n4453 VGND.n4452 4.8005
R20540 VGND.n4654 VGND.n4653 4.8005
R20541 VGND.n2046 VGND.n2045 4.8005
R20542 VGND.n3668 VGND.n3667 4.8005
R20543 VGND.n224 VGND.n223 4.8005
R20544 VGND.n1900 VGND.n1899 4.8005
R20545 VGND.n495 VGND.n494 4.8005
R20546 VGND.n7843 VGND.n7842 4.8005
R20547 VGND.n7457 VGND.n7456 4.8005
R20548 VGND.n6260 VGND.n6259 4.8005
R20549 VGND.n6352 VGND.n6351 4.8005
R20550 VGND.n6358 VGND.n6357 4.8005
R20551 VGND.n4575 VGND.n4574 4.79833
R20552 VGND.n7866 VGND.n7860 4.76901
R20553 VGND.n2595 VGND.n2289 4.72533
R20554 VGND.n5375 VGND.n5374 4.72533
R20555 VGND.n6705 VGND.n6704 4.72533
R20556 VGND.n182 VGND.n180 4.72533
R20557 VGND.n2110 VGND.n2109 4.69383
R20558 VGND.n3283 VGND.n3282 4.69383
R20559 VGND.n8881 VGND.n8880 4.69383
R20560 VGND.n2286 VGND.n2285 4.67352
R20561 VGND.n2170 VGND.n2169 4.67352
R20562 VGND.n2174 VGND.n2173 4.67352
R20563 VGND.n14 VGND.n13 4.67352
R20564 VGND.n5199 VGND.n5198 4.67352
R20565 VGND.n1642 VGND.n1641 4.67352
R20566 VGND.n2105 VGND.n2104 4.67352
R20567 VGND.n2116 VGND.n2115 4.67352
R20568 VGND.n2120 VGND.n2119 4.67352
R20569 VGND.n3309 VGND.n3308 4.67352
R20570 VGND.n3660 VGND.n3659 4.67352
R20571 VGND.n3635 VGND.n3634 4.67352
R20572 VGND.n191 VGND.n190 4.67352
R20573 VGND.n1517 VGND.n1516 4.67352
R20574 VGND.n2578 VGND.n2577 4.65776
R20575 VGND.n6829 VGND.n6828 4.65505
R20576 VGND.n4867 VGND.n4866 4.6505
R20577 VGND.n4871 VGND.n4870 4.6505
R20578 VGND.n4892 VGND.n4088 4.6505
R20579 VGND.n4903 VGND.n3985 4.6505
R20580 VGND.n4905 VGND.n4904 4.6505
R20581 VGND.n4910 VGND.n4907 4.6505
R20582 VGND.n4946 VGND.n4078 4.6505
R20583 VGND.n4947 VGND.n4077 4.6505
R20584 VGND.n4948 VGND.n4075 4.6505
R20585 VGND.n4774 VGND.n4772 4.6505
R20586 VGND.n4779 VGND.n4778 4.6505
R20587 VGND.n4785 VGND.n4784 4.6505
R20588 VGND.n4869 VGND.n4868 4.6505
R20589 VGND.n4881 VGND.n4880 4.6505
R20590 VGND.n4952 VGND.n4951 4.6505
R20591 VGND.n4954 VGND.n4953 4.6505
R20592 VGND.n5021 VGND.n5020 4.6505
R20593 VGND.n5028 VGND.n5027 4.6505
R20594 VGND.n5041 VGND.n4040 4.6505
R20595 VGND.n5077 VGND.n5076 4.6505
R20596 VGND.n5081 VGND.n5080 4.6505
R20597 VGND.n5084 VGND.n4034 4.6505
R20598 VGND.n5087 VGND.n4033 4.6505
R20599 VGND.n4031 VGND.n3989 4.6505
R20600 VGND.n4030 VGND.n3991 4.6505
R20601 VGND.n4029 VGND.n3992 4.6505
R20602 VGND.n4022 VGND.n3995 4.6505
R20603 VGND.n7184 VGND.n1333 4.6505
R20604 VGND.n7169 VGND.n1335 4.6505
R20605 VGND.n7168 VGND.n1337 4.6505
R20606 VGND.n7165 VGND.n1339 4.6505
R20607 VGND.n7161 VGND.n1341 4.6505
R20608 VGND.n7158 VGND.n7156 4.6505
R20609 VGND.n7153 VGND.n1343 4.6505
R20610 VGND.n7057 VGND.n7056 4.6505
R20611 VGND.n7055 VGND.n7054 4.6505
R20612 VGND.n7052 VGND.n7051 4.6505
R20613 VGND.n7050 VGND.n7049 4.6505
R20614 VGND.n7046 VGND.n7045 4.6505
R20615 VGND.n7044 VGND.n7043 4.6505
R20616 VGND.n7042 VGND.n7041 4.6505
R20617 VGND.n7039 VGND.n7038 4.6505
R20618 VGND.n7037 VGND.n7036 4.6505
R20619 VGND.n7035 VGND.n7034 4.6505
R20620 VGND.n7033 VGND.n7032 4.6505
R20621 VGND.n7031 VGND.n7030 4.6505
R20622 VGND.n7029 VGND.n7028 4.6505
R20623 VGND.n7026 VGND.n7025 4.6505
R20624 VGND.n7023 VGND.n7022 4.6505
R20625 VGND.n7021 VGND.n7020 4.6505
R20626 VGND.n7017 VGND.n7016 4.6505
R20627 VGND.n7079 VGND.n7078 4.6505
R20628 VGND.n7069 VGND.n7068 4.6505
R20629 VGND.n7066 VGND.n7065 4.6505
R20630 VGND.n7064 VGND.n7063 4.6505
R20631 VGND.n7062 VGND.n7061 4.6505
R20632 VGND.n7060 VGND.n7059 4.6505
R20633 VGND.n7194 VGND.n7193 4.6505
R20634 VGND.n7192 VGND.n7191 4.6505
R20635 VGND.n7190 VGND.n7189 4.6505
R20636 VGND.n7188 VGND.n7187 4.6505
R20637 VGND.n7186 VGND.n7185 4.6505
R20638 VGND.n7183 VGND.n7182 4.6505
R20639 VGND.n7180 VGND.n7179 4.6505
R20640 VGND.n7178 VGND.n7177 4.6505
R20641 VGND.n7176 VGND.n7175 4.6505
R20642 VGND.n7174 VGND.n7173 4.6505
R20643 VGND.n7171 VGND.n7170 4.6505
R20644 VGND.n7167 VGND.n7166 4.6505
R20645 VGND.n7164 VGND.n7163 4.6505
R20646 VGND.n7160 VGND.n7159 4.6505
R20647 VGND.n7155 VGND.n7154 4.6505
R20648 VGND.n7152 VGND.n7151 4.6505
R20649 VGND.n7148 VGND.n7147 4.6505
R20650 VGND.n7146 VGND.n7145 4.6505
R20651 VGND.n7144 VGND.n7143 4.6505
R20652 VGND.n7140 VGND.n7139 4.6505
R20653 VGND.n7138 VGND.n7137 4.6505
R20654 VGND.n7136 VGND.n1349 4.6505
R20655 VGND.n7135 VGND.n7134 4.6505
R20656 VGND.n7131 VGND.n7130 4.6505
R20657 VGND.n7129 VGND.n7128 4.6505
R20658 VGND.n7123 VGND.n7122 4.6505
R20659 VGND.n7121 VGND.n7120 4.6505
R20660 VGND.n7119 VGND.n7118 4.6505
R20661 VGND.n7117 VGND.n7116 4.6505
R20662 VGND.n7115 VGND.n7114 4.6505
R20663 VGND.n7113 VGND.n7112 4.6505
R20664 VGND.n5023 VGND.n5022 4.6505
R20665 VGND.n5025 VGND.n5024 4.6505
R20666 VGND.n5032 VGND.n5031 4.6505
R20667 VGND.n5036 VGND.n5035 4.6505
R20668 VGND.n5040 VGND.n5039 4.6505
R20669 VGND.n5043 VGND.n5042 4.6505
R20670 VGND.n5050 VGND.n5049 4.6505
R20671 VGND.n5053 VGND.n5052 4.6505
R20672 VGND.n5056 VGND.n5055 4.6505
R20673 VGND.n5058 VGND.n5057 4.6505
R20674 VGND.n5064 VGND.n5063 4.6505
R20675 VGND.n5067 VGND.n5066 4.6505
R20676 VGND.n5069 VGND.n5068 4.6505
R20677 VGND.n5071 VGND.n5070 4.6505
R20678 VGND.n5073 VGND.n5072 4.6505
R20679 VGND.n5079 VGND.n5078 4.6505
R20680 VGND.n5083 VGND.n5082 4.6505
R20681 VGND.n5086 VGND.n5085 4.6505
R20682 VGND.n4032 VGND.n3987 4.6505
R20683 VGND.n4028 VGND.n4027 4.6505
R20684 VGND.n4025 VGND.n4024 4.6505
R20685 VGND.n4023 VGND.n3993 4.6505
R20686 VGND.n4021 VGND.n4020 4.6505
R20687 VGND.n4018 VGND.n4017 4.6505
R20688 VGND.n4016 VGND.n4015 4.6505
R20689 VGND.n5016 VGND.n5015 4.6505
R20690 VGND.n4945 VGND.n4944 4.6505
R20691 VGND.n4942 VGND.n4941 4.6505
R20692 VGND.n4940 VGND.n4939 4.6505
R20693 VGND.n4937 VGND.n4936 4.6505
R20694 VGND.n4935 VGND.n4934 4.6505
R20695 VGND.n4933 VGND.n4932 4.6505
R20696 VGND.n4931 VGND.n4930 4.6505
R20697 VGND.n4929 VGND.n4928 4.6505
R20698 VGND.n4925 VGND.n4924 4.6505
R20699 VGND.n4923 VGND.n4922 4.6505
R20700 VGND.n4921 VGND.n4920 4.6505
R20701 VGND.n4918 VGND.n4917 4.6505
R20702 VGND.n4915 VGND.n4914 4.6505
R20703 VGND.n4913 VGND.n4912 4.6505
R20704 VGND.n4902 VGND.n4901 4.6505
R20705 VGND.n4900 VGND.n4899 4.6505
R20706 VGND.n4894 VGND.n4893 4.6505
R20707 VGND.n4891 VGND.n4890 4.6505
R20708 VGND.n4889 VGND.n4888 4.6505
R20709 VGND.n4887 VGND.n4886 4.6505
R20710 VGND.n4885 VGND.n4884 4.6505
R20711 VGND.n4877 VGND.n4876 4.6505
R20712 VGND.n4875 VGND.n4874 4.6505
R20713 VGND.n4771 VGND.n4766 4.6505
R20714 VGND.n4776 VGND.n4775 4.6505
R20715 VGND.n4783 VGND.n4782 4.6505
R20716 VGND.n4787 VGND.n4786 4.6505
R20717 VGND.n4789 VGND.n4788 4.6505
R20718 VGND.n4793 VGND.n4792 4.6505
R20719 VGND.n4657 VGND.n4550 4.6505
R20720 VGND.n4614 VGND.n4566 4.6505
R20721 VGND.n4613 VGND.n4567 4.6505
R20722 VGND.n4385 VGND.n4384 4.6505
R20723 VGND.n4410 VGND.n4409 4.6505
R20724 VGND.n4415 VGND.n4414 4.6505
R20725 VGND.n4418 VGND.n4220 4.6505
R20726 VGND.n4420 VGND.n4419 4.6505
R20727 VGND.n4439 VGND.n4438 4.6505
R20728 VGND.n4441 VGND.n4217 4.6505
R20729 VGND.n4443 VGND.n4169 4.6505
R20730 VGND.n4458 VGND.n4456 4.6505
R20731 VGND.n4472 VGND.n4471 4.6505
R20732 VGND.n4474 VGND.n4473 4.6505
R20733 VGND.n4683 VGND.n4163 4.6505
R20734 VGND.n4289 VGND.n4288 4.6505
R20735 VGND.n4293 VGND.n4292 4.6505
R20736 VGND.n4106 VGND.n4104 4.6505
R20737 VGND.n4109 VGND.n4097 4.6505
R20738 VGND.n4111 VGND.n4110 4.6505
R20739 VGND.n4114 VGND.n4113 4.6505
R20740 VGND.n4678 VGND.n4677 4.6505
R20741 VGND.n4663 VGND.n4662 4.6505
R20742 VGND.n4282 VGND.n4281 4.6505
R20743 VGND.n4437 VGND.n4436 4.6505
R20744 VGND.n4523 VGND.n4522 4.6505
R20745 VGND.n4525 VGND.n4524 4.6505
R20746 VGND.n4530 VGND.n4529 4.6505
R20747 VGND.n4533 VGND.n4532 4.6505
R20748 VGND.n4534 VGND.n4172 4.6505
R20749 VGND.n4537 VGND.n4536 4.6505
R20750 VGND.n4542 VGND.n4541 4.6505
R20751 VGND.n4545 VGND.n4544 4.6505
R20752 VGND.n4549 VGND.n4548 4.6505
R20753 VGND.n4656 VGND.n4655 4.6505
R20754 VGND VGND.n4654 4.6505
R20755 VGND.n4651 VGND.n4650 4.6505
R20756 VGND.n4634 VGND.n4556 4.6505
R20757 VGND.n4633 VGND.n4632 4.6505
R20758 VGND.n4629 VGND.n4628 4.6505
R20759 VGND.n4625 VGND.n4624 4.6505
R20760 VGND.n4623 VGND.n4622 4.6505
R20761 VGND.n4616 VGND.n4615 4.6505
R20762 VGND.n1448 VGND.n1391 4.6505
R20763 VGND.n1431 VGND.n1402 4.6505
R20764 VGND.n1430 VGND.n1404 4.6505
R20765 VGND.n1427 VGND.n1426 4.6505
R20766 VGND.n1425 VGND.n1406 4.6505
R20767 VGND.n1466 VGND.n1465 4.6505
R20768 VGND.n1452 VGND.n1451 4.6505
R20769 VGND.n1450 VGND.n1449 4.6505
R20770 VGND.n1447 VGND.n1446 4.6505
R20771 VGND.n1444 VGND.n1443 4.6505
R20772 VGND.n1441 VGND.n1440 4.6505
R20773 VGND.n1437 VGND.n1436 4.6505
R20774 VGND.n1429 VGND.n1428 4.6505
R20775 VGND.n1424 VGND.n1423 4.6505
R20776 VGND.n1417 VGND.n1416 4.6505
R20777 VGND.n1414 VGND.n1413 4.6505
R20778 VGND.n4594 VGND.n4593 4.6505
R20779 VGND.n4599 VGND.n4598 4.6505
R20780 VGND.n4602 VGND.n4601 4.6505
R20781 VGND.n4606 VGND.n4605 4.6505
R20782 VGND.n4608 VGND.n4607 4.6505
R20783 VGND.n4610 VGND.n4609 4.6505
R20784 VGND.n4612 VGND.n4611 4.6505
R20785 VGND.n4636 VGND.n4635 4.6505
R20786 VGND.n4639 VGND.n4638 4.6505
R20787 VGND.n4641 VGND.n4640 4.6505
R20788 VGND.n4645 VGND.n4644 4.6505
R20789 VGND.n4647 VGND.n4646 4.6505
R20790 VGND.n4649 VGND.n4648 4.6505
R20791 VGND.n4476 VGND.n4475 4.6505
R20792 VGND.n4470 VGND.n4469 4.6505
R20793 VGND.n4468 VGND.n4467 4.6505
R20794 VGND.n4466 VGND.n4465 4.6505
R20795 VGND.n4462 VGND.n4461 4.6505
R20796 VGND.n4455 VGND.n4216 4.6505
R20797 VGND.n4454 VGND.n4453 4.6505
R20798 VGND VGND.n4442 4.6505
R20799 VGND.n4429 VGND.n4428 4.6505
R20800 VGND.n4426 VGND.n4425 4.6505
R20801 VGND.n4417 VGND.n4416 4.6505
R20802 VGND.n4412 VGND.n4411 4.6505
R20803 VGND.n4407 VGND.n4406 4.6505
R20804 VGND.n4405 VGND.n4404 4.6505
R20805 VGND.n4401 VGND.n4400 4.6505
R20806 VGND.n4399 VGND.n4398 4.6505
R20807 VGND.n4397 VGND.n4396 4.6505
R20808 VGND.n4395 VGND.n4394 4.6505
R20809 VGND.n4391 VGND.n4390 4.6505
R20810 VGND.n4389 VGND.n4223 4.6505
R20811 VGND.n4388 VGND.n4387 4.6505
R20812 VGND.n4383 VGND.n4382 4.6505
R20813 VGND.n4298 VGND.n4297 4.6505
R20814 VGND.n4296 VGND.n4295 4.6505
R20815 VGND.n4291 VGND.n4290 4.6505
R20816 VGND.n4286 VGND.n4285 4.6505
R20817 VGND.n4284 VGND.n4283 4.6505
R20818 VGND.n4276 VGND.n4275 4.6505
R20819 VGND.n4274 VGND.n4273 4.6505
R20820 VGND.n4271 VGND.n4270 4.6505
R20821 VGND.n4269 VGND.n4268 4.6505
R20822 VGND.n4266 VGND.n4265 4.6505
R20823 VGND.n4264 VGND.n4263 4.6505
R20824 VGND.n4262 VGND.n4261 4.6505
R20825 VGND.n4260 VGND.n4259 4.6505
R20826 VGND.n4256 VGND.n4255 4.6505
R20827 VGND.n4254 VGND.n4253 4.6505
R20828 VGND.n4252 VGND.n4251 4.6505
R20829 VGND.n4250 VGND.n4249 4.6505
R20830 VGND.n4245 VGND.n4244 4.6505
R20831 VGND.n4242 VGND.n4241 4.6505
R20832 VGND.n4665 VGND.n4664 4.6505
R20833 VGND.n4669 VGND.n4668 4.6505
R20834 VGND.n4672 VGND.n4671 4.6505
R20835 VGND.n4674 VGND.n4673 4.6505
R20836 VGND.n4682 VGND.n4681 4.6505
R20837 VGND.n4685 VGND.n4684 4.6505
R20838 VGND.n4687 VGND.n4686 4.6505
R20839 VGND.n4690 VGND.n4689 4.6505
R20840 VGND.n4693 VGND.n4692 4.6505
R20841 VGND.n4695 VGND.n4694 4.6505
R20842 VGND.n4103 VGND.n4098 4.6505
R20843 VGND.n4108 VGND.n4107 4.6505
R20844 VGND.n4116 VGND.n4115 4.6505
R20845 VGND.n4119 VGND.n4118 4.6505
R20846 VGND.n4123 VGND.n4122 4.6505
R20847 VGND.n3280 VGND.n2660 4.6505
R20848 VGND.n3279 VGND.n2661 4.6505
R20849 VGND.n3264 VGND.n3210 4.6505
R20850 VGND.n3247 VGND.n3246 4.6505
R20851 VGND.n3245 VGND.n3224 4.6505
R20852 VGND.n3451 VGND.n3450 4.6505
R20853 VGND.n3449 VGND.n3448 4.6505
R20854 VGND.n3445 VGND.n3444 4.6505
R20855 VGND.n3441 VGND.n3440 4.6505
R20856 VGND.n3439 VGND.n3438 4.6505
R20857 VGND.n3437 VGND.n3436 4.6505
R20858 VGND.n3435 VGND.n3434 4.6505
R20859 VGND.n3430 VGND.n3429 4.6505
R20860 VGND.n3427 VGND.n3426 4.6505
R20861 VGND.n3425 VGND.n2108 4.6505
R20862 VGND.n3423 VGND.n3422 4.6505
R20863 VGND.n3417 VGND.n3416 4.6505
R20864 VGND.n3415 VGND.n3414 4.6505
R20865 VGND.n3413 VGND.n3412 4.6505
R20866 VGND.n3411 VGND.n3410 4.6505
R20867 VGND.n3409 VGND.n3408 4.6505
R20868 VGND.n3407 VGND.n3406 4.6505
R20869 VGND.n3402 VGND.n3401 4.6505
R20870 VGND.n3399 VGND.n3398 4.6505
R20871 VGND.n3395 VGND.n3394 4.6505
R20872 VGND.n3393 VGND.n3392 4.6505
R20873 VGND.n3391 VGND.n3390 4.6505
R20874 VGND.n3389 VGND.n3388 4.6505
R20875 VGND.n3387 VGND.n3386 4.6505
R20876 VGND.n3385 VGND.n3384 4.6505
R20877 VGND.n3324 VGND.n3323 4.6505
R20878 VGND.n3317 VGND.n3316 4.6505
R20879 VGND.n3312 VGND.n3311 4.6505
R20880 VGND.n3296 VGND.n3295 4.6505
R20881 VGND.n3294 VGND.n3293 4.6505
R20882 VGND.n3292 VGND.n3291 4.6505
R20883 VGND.n3290 VGND.n3289 4.6505
R20884 VGND.n3288 VGND.n3287 4.6505
R20885 VGND.n3285 VGND.n3284 4.6505
R20886 VGND.n2790 VGND.n2757 4.6505
R20887 VGND.n2796 VGND.n2795 4.6505
R20888 VGND.n2797 VGND.n2756 4.6505
R20889 VGND.n2821 VGND.n2820 4.6505
R20890 VGND.n2825 VGND.n2824 4.6505
R20891 VGND.n2858 VGND.n2857 4.6505
R20892 VGND.n2861 VGND.n2860 4.6505
R20893 VGND.n2864 VGND.n2747 4.6505
R20894 VGND.n2966 VGND.n2896 4.6505
R20895 VGND.n2942 VGND.n2941 4.6505
R20896 VGND.n2930 VGND.n2901 4.6505
R20897 VGND.n2927 VGND.n2902 4.6505
R20898 VGND.n2918 VGND.n2916 4.6505
R20899 VGND.n2915 VGND.n2906 4.6505
R20900 VGND.n2912 VGND.n2907 4.6505
R20901 VGND.n2965 VGND.n2964 4.6505
R20902 VGND.n2962 VGND.n2961 4.6505
R20903 VGND.n2959 VGND.n2958 4.6505
R20904 VGND.n2957 VGND.n2956 4.6505
R20905 VGND.n2954 VGND.n2953 4.6505
R20906 VGND.n2949 VGND.n2948 4.6505
R20907 VGND.n2944 VGND.n2943 4.6505
R20908 VGND.n2940 VGND.n2939 4.6505
R20909 VGND.n2938 VGND.n2937 4.6505
R20910 VGND.n2934 VGND.n2933 4.6505
R20911 VGND.n2932 VGND.n2931 4.6505
R20912 VGND.n2929 VGND.n2928 4.6505
R20913 VGND.n2926 VGND.n2925 4.6505
R20914 VGND.n2920 VGND.n2919 4.6505
R20915 VGND.n2914 VGND.n2913 4.6505
R20916 VGND.n2983 VGND.n2982 4.6505
R20917 VGND.n2787 VGND.n2786 4.6505
R20918 VGND.n2789 VGND.n2788 4.6505
R20919 VGND.n2792 VGND.n2791 4.6505
R20920 VGND.n2794 VGND.n2793 4.6505
R20921 VGND.n2803 VGND.n2802 4.6505
R20922 VGND.n2807 VGND.n2806 4.6505
R20923 VGND.n2811 VGND.n2810 4.6505
R20924 VGND.n2812 VGND.n2663 4.6505
R20925 VGND.n2815 VGND.n2814 4.6505
R20926 VGND.n2823 VGND.n2822 4.6505
R20927 VGND.n2831 VGND.n2830 4.6505
R20928 VGND.n2835 VGND.n2834 4.6505
R20929 VGND.n2838 VGND.n2837 4.6505
R20930 VGND.n2842 VGND.n2841 4.6505
R20931 VGND.n2845 VGND.n2844 4.6505
R20932 VGND.n2846 VGND.n2752 4.6505
R20933 VGND.n2848 VGND.n2847 4.6505
R20934 VGND.n2851 VGND.n2850 4.6505
R20935 VGND.n2853 VGND.n2852 4.6505
R20936 VGND.n2856 VGND.n2855 4.6505
R20937 VGND.n2863 VGND.n2862 4.6505
R20938 VGND.n2871 VGND.n2870 4.6505
R20939 VGND.n2873 VGND.n2872 4.6505
R20940 VGND.n2875 VGND.n2874 4.6505
R20941 VGND.n3249 VGND.n3248 4.6505
R20942 VGND.n3254 VGND.n3253 4.6505
R20943 VGND.n3256 VGND.n3255 4.6505
R20944 VGND.n3258 VGND.n3257 4.6505
R20945 VGND.n3260 VGND.n3259 4.6505
R20946 VGND.n3261 VGND.n3214 4.6505
R20947 VGND.n3263 VGND.n3262 4.6505
R20948 VGND.n3266 VGND.n3265 4.6505
R20949 VGND.n3270 VGND.n3269 4.6505
R20950 VGND.n3272 VGND.n3271 4.6505
R20951 VGND.n3276 VGND.n3275 4.6505
R20952 VGND.n3278 VGND.n3277 4.6505
R20953 VGND.n2055 VGND.n2054 4.6505
R20954 VGND.n2058 VGND.n2057 4.6505
R20955 VGND.n2062 VGND.n2061 4.6505
R20956 VGND.n2065 VGND.n2064 4.6505
R20957 VGND.n2069 VGND.n2068 4.6505
R20958 VGND.n2072 VGND.n2071 4.6505
R20959 VGND.n8971 VGND.n8970 4.6505
R20960 VGND.n8973 VGND.n8972 4.6505
R20961 VGND.n8976 VGND.n8975 4.6505
R20962 VGND.n8979 VGND.n8978 4.6505
R20963 VGND.n3683 VGND.n3682 4.6505
R20964 VGND.n3686 VGND.n3685 4.6505
R20965 VGND.n3687 VGND.n3665 4.6505
R20966 VGND.n3663 VGND.n3662 4.6505
R20967 VGND.n3655 VGND.n3654 4.6505
R20968 VGND.n3653 VGND.n3652 4.6505
R20969 VGND.n3649 VGND.n3648 4.6505
R20970 VGND.n3646 VGND.n3645 4.6505
R20971 VGND.n3644 VGND.n3643 4.6505
R20972 VGND.n3642 VGND.n3641 4.6505
R20973 VGND.n3640 VGND.n3639 4.6505
R20974 VGND.n8907 VGND.n8906 4.6505
R20975 VGND.n8904 VGND.n8903 4.6505
R20976 VGND.n8899 VGND.n8898 4.6505
R20977 VGND.n8894 VGND.n8893 4.6505
R20978 VGND.n8887 VGND.n8886 4.6505
R20979 VGND.n8885 VGND.n87 4.6505
R20980 VGND.n8883 VGND.n8882 4.6505
R20981 VGND.n8878 VGND.n8877 4.6505
R20982 VGND.n8873 VGND.n8872 4.6505
R20983 VGND.n8871 VGND.n8870 4.6505
R20984 VGND.n8869 VGND.n8868 4.6505
R20985 VGND.n8867 VGND.n8866 4.6505
R20986 VGND.n8865 VGND.n8864 4.6505
R20987 VGND.n8863 VGND.n8862 4.6505
R20988 VGND.n8921 VGND.n8920 4.6505
R20989 VGND.n8923 VGND.n80 4.6505
R20990 VGND.n8925 VGND.n8924 4.6505
R20991 VGND.n8935 VGND.n8934 4.6505
R20992 VGND.n8939 VGND.n8938 4.6505
R20993 VGND.n8961 VGND.n8960 4.6505
R20994 VGND.n8963 VGND.n8962 4.6505
R20995 VGND.n8965 VGND.n8964 4.6505
R20996 VGND.n3043 VGND.n3036 4.6505
R20997 VGND.n3047 VGND.n3046 4.6505
R20998 VGND.n3049 VGND.n3048 4.6505
R20999 VGND.n2716 VGND.n2715 4.6505
R21000 VGND.n2688 VGND.n2675 4.6505
R21001 VGND.n2687 VGND.n2679 4.6505
R21002 VGND.n2685 VGND.n2680 4.6505
R21003 VGND.n2736 VGND.n2735 4.6505
R21004 VGND.n2732 VGND.n2731 4.6505
R21005 VGND.n2730 VGND.n2729 4.6505
R21006 VGND.n2728 VGND.n2727 4.6505
R21007 VGND.n2726 VGND.n2725 4.6505
R21008 VGND.n2714 VGND.n2713 4.6505
R21009 VGND.n2712 VGND.n2711 4.6505
R21010 VGND.n2708 VGND.n2707 4.6505
R21011 VGND.n2704 VGND.n2703 4.6505
R21012 VGND.n2700 VGND.n2699 4.6505
R21013 VGND.n2698 VGND.n2697 4.6505
R21014 VGND.n2696 VGND.n2695 4.6505
R21015 VGND.n2691 VGND.n2690 4.6505
R21016 VGND.n3191 VGND.n3190 4.6505
R21017 VGND.n3042 VGND.n3041 4.6505
R21018 VGND.n3045 VGND.n3044 4.6505
R21019 VGND.n3053 VGND.n3052 4.6505
R21020 VGND.n3056 VGND.n3055 4.6505
R21021 VGND.n3059 VGND.n3058 4.6505
R21022 VGND.n3067 VGND.n3066 4.6505
R21023 VGND.n3069 VGND.n3068 4.6505
R21024 VGND.n3073 VGND.n3072 4.6505
R21025 VGND.n3076 VGND.n3075 4.6505
R21026 VGND.n3079 VGND.n3078 4.6505
R21027 VGND.n3081 VGND.n3080 4.6505
R21028 VGND.n3084 VGND.n3083 4.6505
R21029 VGND.n3086 VGND.n3085 4.6505
R21030 VGND.n3089 VGND.n3088 4.6505
R21031 VGND.n3091 VGND.n3090 4.6505
R21032 VGND.n3093 VGND.n3092 4.6505
R21033 VGND.n3096 VGND.n3095 4.6505
R21034 VGND.n3100 VGND.n3099 4.6505
R21035 VGND.n3103 VGND.n3102 4.6505
R21036 VGND.n3106 VGND.n3105 4.6505
R21037 VGND.n3110 VGND.n3109 4.6505
R21038 VGND.n3112 VGND.n3111 4.6505
R21039 VGND.n3114 VGND.n3113 4.6505
R21040 VGND.n3116 VGND.n3115 4.6505
R21041 VGND.n3118 VGND.n3117 4.6505
R21042 VGND.n3120 VGND.n3119 4.6505
R21043 VGND.n3122 VGND.n3121 4.6505
R21044 VGND.n3126 VGND.n3125 4.6505
R21045 VGND.n3128 VGND.n3127 4.6505
R21046 VGND.n3132 VGND.n3131 4.6505
R21047 VGND.n9007 VGND.n9006 4.6505
R21048 VGND.n9005 VGND.n9004 4.6505
R21049 VGND.n9003 VGND.n9002 4.6505
R21050 VGND.n9000 VGND.n8999 4.6505
R21051 VGND.n8998 VGND.n8997 4.6505
R21052 VGND.n8996 VGND.n8995 4.6505
R21053 VGND.n8994 VGND.n8993 4.6505
R21054 VGND.n8990 VGND.n8989 4.6505
R21055 VGND.n8988 VGND.n8987 4.6505
R21056 VGND.n8986 VGND.n8985 4.6505
R21057 VGND.n8984 VGND.n8983 4.6505
R21058 VGND.n8977 VGND.n77 4.6505
R21059 VGND.n8956 VGND.n8955 4.6505
R21060 VGND.n8954 VGND.n8953 4.6505
R21061 VGND.n8951 VGND.n8950 4.6505
R21062 VGND.n8949 VGND.n8948 4.6505
R21063 VGND.n8945 VGND.n8944 4.6505
R21064 VGND.n8941 VGND.n8940 4.6505
R21065 VGND.n3677 VGND.n3676 4.6505
R21066 VGND.n3680 VGND.n3679 4.6505
R21067 VGND.n3689 VGND.n3688 4.6505
R21068 VGND.n3692 VGND.n3691 4.6505
R21069 VGND.n3695 VGND.n3694 4.6505
R21070 VGND.n8783 VGND.n161 4.6505
R21071 VGND.n8774 VGND.n8770 4.6505
R21072 VGND.n8767 VGND.n167 4.6505
R21073 VGND.n8755 VGND.n172 4.6505
R21074 VGND.n8752 VGND.n173 4.6505
R21075 VGND.n3979 VGND.n3876 4.6505
R21076 VGND.n3978 VGND.n3877 4.6505
R21077 VGND.n3955 VGND.n3883 4.6505
R21078 VGND.n3952 VGND.n3885 4.6505
R21079 VGND.n3922 VGND.n3920 4.6505
R21080 VGND.n3783 VGND.n3778 4.6505
R21081 VGND.n3785 VGND.n3784 4.6505
R21082 VGND.n3788 VGND.n3787 4.6505
R21083 VGND.n3792 VGND.n3777 4.6505
R21084 VGND.n3870 VGND.n3869 4.6505
R21085 VGND.n3962 VGND.n3961 4.6505
R21086 VGND.n3947 VGND.n3946 4.6505
R21087 VGND.n3933 VGND.n3932 4.6505
R21088 VGND.n8782 VGND.n8781 4.6505
R21089 VGND.n8780 VGND.n8779 4.6505
R21090 VGND.n8778 VGND.n8777 4.6505
R21091 VGND.n8764 VGND.n8763 4.6505
R21092 VGND.n8761 VGND.n8760 4.6505
R21093 VGND.n8758 VGND.n8757 4.6505
R21094 VGND.n8751 VGND.n8750 4.6505
R21095 VGND.n8748 VGND.n8747 4.6505
R21096 VGND.n8745 VGND.n8744 4.6505
R21097 VGND.n8742 VGND.n8741 4.6505
R21098 VGND.n8739 VGND.n8738 4.6505
R21099 VGND.n8736 VGND.n8735 4.6505
R21100 VGND.n8734 VGND.n8733 4.6505
R21101 VGND.n8732 VGND.n184 4.6505
R21102 VGND.n8729 VGND.n8728 4.6505
R21103 VGND.n8726 VGND.n8725 4.6505
R21104 VGND.n8722 VGND.n8721 4.6505
R21105 VGND.n8718 VGND.n194 4.6505
R21106 VGND.n8629 VGND.n219 4.6505
R21107 VGND.n8593 VGND.n240 4.6505
R21108 VGND.n8573 VGND.n8572 4.6505
R21109 VGND.n8502 VGND.n8501 4.6505
R21110 VGND.n8484 VGND.n8483 4.6505
R21111 VGND.n8482 VGND.n8456 4.6505
R21112 VGND.n8481 VGND.n8457 4.6505
R21113 VGND.n8480 VGND.n8459 4.6505
R21114 VGND.n8524 VGND.n8523 4.6505
R21115 VGND.n8522 VGND.n8521 4.6505
R21116 VGND.n8519 VGND.n8518 4.6505
R21117 VGND.n8517 VGND.n8516 4.6505
R21118 VGND.n8514 VGND.n8513 4.6505
R21119 VGND.n8509 VGND.n8508 4.6505
R21120 VGND.n8504 VGND.n8503 4.6505
R21121 VGND.n8500 VGND.n8499 4.6505
R21122 VGND.n8498 VGND.n8497 4.6505
R21123 VGND.n8494 VGND.n8493 4.6505
R21124 VGND.n8492 VGND.n8491 4.6505
R21125 VGND.n8489 VGND.n8488 4.6505
R21126 VGND.n8486 VGND.n8485 4.6505
R21127 VGND.n8479 VGND.n8478 4.6505
R21128 VGND.n8477 VGND.n8476 4.6505
R21129 VGND.n8475 VGND.n8474 4.6505
R21130 VGND.n8468 VGND.n8467 4.6505
R21131 VGND.n8538 VGND.n8537 4.6505
R21132 VGND.n8648 VGND.n8647 4.6505
R21133 VGND.n8645 VGND.n8644 4.6505
R21134 VGND.n8643 VGND.n8642 4.6505
R21135 VGND.n8639 VGND.n8638 4.6505
R21136 VGND.n8637 VGND.n8636 4.6505
R21137 VGND.n8635 VGND.n8634 4.6505
R21138 VGND.n8631 VGND.n8630 4.6505
R21139 VGND.n8628 VGND.n8627 4.6505
R21140 VGND.n8626 VGND.n8625 4.6505
R21141 VGND.n8623 VGND.n8622 4.6505
R21142 VGND.n8621 VGND.n8620 4.6505
R21143 VGND.n8617 VGND.n8616 4.6505
R21144 VGND.n8615 VGND.n8614 4.6505
R21145 VGND.n8613 VGND.n8612 4.6505
R21146 VGND.n8611 VGND.n8610 4.6505
R21147 VGND.n8608 VGND.n8607 4.6505
R21148 VGND.n8605 VGND.n8604 4.6505
R21149 VGND.n8596 VGND.n8595 4.6505
R21150 VGND.n8594 VGND.n237 4.6505
R21151 VGND.n8592 VGND.n8591 4.6505
R21152 VGND.n8587 VGND.n8586 4.6505
R21153 VGND.n8582 VGND.n8581 4.6505
R21154 VGND.n8579 VGND.n8578 4.6505
R21155 VGND.n8575 VGND.n8574 4.6505
R21156 VGND.n8720 VGND.n8719 4.6505
R21157 VGND.n8754 VGND.n8753 4.6505
R21158 VGND.n8766 VGND.n8765 4.6505
R21159 VGND.n8769 VGND.n8768 4.6505
R21160 VGND VGND.n8775 4.6505
R21161 VGND.n3924 VGND.n3923 4.6505
R21162 VGND.n3926 VGND.n3925 4.6505
R21163 VGND.n3928 VGND.n3927 4.6505
R21164 VGND.n3935 VGND.n3934 4.6505
R21165 VGND.n3937 VGND.n3936 4.6505
R21166 VGND.n3939 VGND.n3938 4.6505
R21167 VGND.n3941 VGND.n3940 4.6505
R21168 VGND.n3949 VGND.n3948 4.6505
R21169 VGND.n3951 VGND.n3950 4.6505
R21170 VGND.n3954 VGND.n3953 4.6505
R21171 VGND.n3958 VGND.n3957 4.6505
R21172 VGND.n3967 VGND.n3966 4.6505
R21173 VGND.n3970 VGND.n3969 4.6505
R21174 VGND.n3972 VGND.n3971 4.6505
R21175 VGND.n3974 VGND.n3973 4.6505
R21176 VGND.n3977 VGND.n3976 4.6505
R21177 VGND.n3875 VGND.n1864 4.6505
R21178 VGND.n3874 VGND.n3873 4.6505
R21179 VGND.n3872 VGND.n3871 4.6505
R21180 VGND.n3866 VGND.n3865 4.6505
R21181 VGND.n3863 VGND.n3862 4.6505
R21182 VGND.n3861 VGND.n3860 4.6505
R21183 VGND.n3856 VGND.n3855 4.6505
R21184 VGND.n3853 VGND.n3852 4.6505
R21185 VGND.n3850 VGND.n3849 4.6505
R21186 VGND.n3845 VGND.n3844 4.6505
R21187 VGND.n3843 VGND.n1865 4.6505
R21188 VGND.n3790 VGND.n3789 4.6505
R21189 VGND.n3794 VGND.n3793 4.6505
R21190 VGND.n3799 VGND.n3798 4.6505
R21191 VGND.n3801 VGND.n3800 4.6505
R21192 VGND.n7838 VGND.n7837 4.6505
R21193 VGND.n7873 VGND.n7872 4.6505
R21194 VGND.n7941 VGND.n7890 4.6505
R21195 VGND.n1957 VGND.n1919 4.6505
R21196 VGND.n1951 VGND.n1928 4.6505
R21197 VGND.n7810 VGND.n7809 4.6505
R21198 VGND.n1954 VGND.n1953 4.6505
R21199 VGND.n1938 VGND.n1937 4.6505
R21200 VGND.n7801 VGND.n7800 4.6505
R21201 VGND.n7790 VGND.n7789 4.6505
R21202 VGND.n7780 VGND.n524 4.6505
R21203 VGND.n7779 VGND.n7778 4.6505
R21204 VGND.n7777 VGND.n7776 4.6505
R21205 VGND.n7775 VGND.n7774 4.6505
R21206 VGND.n7773 VGND.n7772 4.6505
R21207 VGND.n7768 VGND.n7767 4.6505
R21208 VGND.n7763 VGND.n7762 4.6505
R21209 VGND.n7827 VGND.n7826 4.6505
R21210 VGND.n7833 VGND.n7832 4.6505
R21211 VGND.n7856 VGND.n7855 4.6505
R21212 VGND.n7860 VGND.n7859 4.6505
R21213 VGND.n7923 VGND.n7905 4.6505
R21214 VGND.n8057 VGND.n483 4.6505
R21215 VGND.n8056 VGND.n485 4.6505
R21216 VGND.n8028 VGND.n7950 4.6505
R21217 VGND.n8019 VGND.n7953 4.6505
R21218 VGND.n8016 VGND.n7955 4.6505
R21219 VGND.n8009 VGND.n7958 4.6505
R21220 VGND.n8000 VGND.n7998 4.6505
R21221 VGND.n7997 VGND.n7962 4.6505
R21222 VGND.n7996 VGND.n7964 4.6505
R21223 VGND.n7993 VGND.n7966 4.6505
R21224 VGND.n7990 VGND.n7968 4.6505
R21225 VGND.n8394 VGND.n8340 4.6505
R21226 VGND.n8378 VGND.n8346 4.6505
R21227 VGND.n8375 VGND.n8347 4.6505
R21228 VGND.n8374 VGND.n8348 4.6505
R21229 VGND.n8373 VGND.n8349 4.6505
R21230 VGND.n8370 VGND.n8369 4.6505
R21231 VGND.n8404 VGND.n8403 4.6505
R21232 VGND.n8402 VGND.n8401 4.6505
R21233 VGND.n8400 VGND.n8399 4.6505
R21234 VGND.n8398 VGND.n8397 4.6505
R21235 VGND.n8393 VGND.n8392 4.6505
R21236 VGND.n8391 VGND.n8390 4.6505
R21237 VGND.n8389 VGND.n8342 4.6505
R21238 VGND.n8388 VGND.n8387 4.6505
R21239 VGND.n8377 VGND.n8376 4.6505
R21240 VGND.n8372 VGND.n8371 4.6505
R21241 VGND.n8368 VGND.n8350 4.6505
R21242 VGND.n8367 VGND.n8366 4.6505
R21243 VGND.n8361 VGND.n8360 4.6505
R21244 VGND.n8359 VGND.n8358 4.6505
R21245 VGND.n8061 VGND.n8060 4.6505
R21246 VGND.n8059 VGND.n8058 4.6505
R21247 VGND.n8055 VGND.n8054 4.6505
R21248 VGND.n8052 VGND.n8051 4.6505
R21249 VGND.n8050 VGND.n8049 4.6505
R21250 VGND.n8048 VGND.n8047 4.6505
R21251 VGND.n8046 VGND.n8045 4.6505
R21252 VGND.n8043 VGND.n8042 4.6505
R21253 VGND.n8040 VGND.n8039 4.6505
R21254 VGND.n8038 VGND.n8037 4.6505
R21255 VGND.n8035 VGND.n8034 4.6505
R21256 VGND.n8032 VGND.n8031 4.6505
R21257 VGND.n8030 VGND.n8029 4.6505
R21258 VGND.n8027 VGND.n8026 4.6505
R21259 VGND.n8025 VGND.n8024 4.6505
R21260 VGND.n8023 VGND.n8022 4.6505
R21261 VGND.n8018 VGND.n8017 4.6505
R21262 VGND.n8015 VGND.n8014 4.6505
R21263 VGND.n8013 VGND.n8012 4.6505
R21264 VGND.n8008 VGND.n8007 4.6505
R21265 VGND.n8006 VGND.n8005 4.6505
R21266 VGND.n8002 VGND.n8001 4.6505
R21267 VGND.n7995 VGND.n7994 4.6505
R21268 VGND.n7992 VGND.n7991 4.6505
R21269 VGND.n7989 VGND.n7988 4.6505
R21270 VGND.n8063 VGND.n8062 4.6505
R21271 VGND.n7922 VGND.n7921 4.6505
R21272 VGND.n7925 VGND.n7924 4.6505
R21273 VGND.n7927 VGND.n7926 4.6505
R21274 VGND.n7932 VGND.n7931 4.6505
R21275 VGND.n7934 VGND.n7933 4.6505
R21276 VGND.n7936 VGND.n7935 4.6505
R21277 VGND.n7938 VGND.n7937 4.6505
R21278 VGND.n7940 VGND.n7939 4.6505
R21279 VGND.n7889 VGND.n497 4.6505
R21280 VGND.n7888 VGND.n7887 4.6505
R21281 VGND.n7886 VGND.n7885 4.6505
R21282 VGND.n7881 VGND.n7880 4.6505
R21283 VGND.n7879 VGND.n7878 4.6505
R21284 VGND.n7877 VGND.n7876 4.6505
R21285 VGND.n7871 VGND.n7870 4.6505
R21286 VGND.n7867 VGND.n7866 4.6505
R21287 VGND.n7850 VGND.n7849 4.6505
R21288 VGND.n7847 VGND.n7846 4.6505
R21289 VGND.n7840 VGND.n7839 4.6505
R21290 VGND.n7835 VGND.n7834 4.6505
R21291 VGND.n7830 VGND.n7829 4.6505
R21292 VGND.n7821 VGND.n7820 4.6505
R21293 VGND.n7766 VGND.n7765 4.6505
R21294 VGND.n7782 VGND.n7781 4.6505
R21295 VGND.n7784 VGND.n7783 4.6505
R21296 VGND.n7787 VGND.n7786 4.6505
R21297 VGND.n7795 VGND.n7794 4.6505
R21298 VGND.n7797 VGND.n7796 4.6505
R21299 VGND.n7803 VGND.n7802 4.6505
R21300 VGND.n7805 VGND.n7804 4.6505
R21301 VGND.n7808 VGND.n7807 4.6505
R21302 VGND.n1929 VGND.n508 4.6505
R21303 VGND.n1934 VGND.n1933 4.6505
R21304 VGND.n1940 VGND.n1939 4.6505
R21305 VGND.n1942 VGND.n1941 4.6505
R21306 VGND.n1948 VGND.n1947 4.6505
R21307 VGND.n1950 VGND.n1949 4.6505
R21308 VGND.n1956 VGND.n1955 4.6505
R21309 VGND.n1888 VGND 4.6505
R21310 VGND.n1893 VGND.n1892 4.6505
R21311 VGND.n1895 VGND.n1883 4.6505
R21312 VGND.n1897 VGND.n1896 4.6505
R21313 VGND.n1905 VGND.n1904 4.6505
R21314 VGND.n1906 VGND.n1877 4.6505
R21315 VGND.n1908 VGND.n1907 4.6505
R21316 VGND.n8255 VGND.n450 4.6505
R21317 VGND.n8272 VGND.n8271 4.6505
R21318 VGND.n663 VGND.n662 4.6505
R21319 VGND.n651 VGND.n650 4.6505
R21320 VGND.n645 VGND.n610 4.6505
R21321 VGND.n642 VGND.n612 4.6505
R21322 VGND.n625 VGND.n613 4.6505
R21323 VGND.n624 VGND.n615 4.6505
R21324 VGND.n621 VGND.n617 4.6505
R21325 VGND.n618 VGND.n451 4.6505
R21326 VGND.n8248 VGND.n454 4.6505
R21327 VGND.n700 VGND.n699 4.6505
R21328 VGND.n7563 VGND.n7562 4.6505
R21329 VGND.n7567 VGND.n7566 4.6505
R21330 VGND.n7571 VGND.n7570 4.6505
R21331 VGND.n7573 VGND.n7572 4.6505
R21332 VGND.n7577 VGND.n7576 4.6505
R21333 VGND.n7581 VGND.n7580 4.6505
R21334 VGND.n7583 VGND.n7582 4.6505
R21335 VGND.n7588 VGND.n7587 4.6505
R21336 VGND.n7591 VGND.n7590 4.6505
R21337 VGND.n7593 VGND.n7592 4.6505
R21338 VGND.n7596 VGND.n7595 4.6505
R21339 VGND.n7597 VGND.n683 4.6505
R21340 VGND.n7683 VGND.n7682 4.6505
R21341 VGND.n7681 VGND.n684 4.6505
R21342 VGND.n7680 VGND.n7679 4.6505
R21343 VGND.n7672 VGND.n7671 4.6505
R21344 VGND.n7668 VGND.n7667 4.6505
R21345 VGND.n7665 VGND.n7664 4.6505
R21346 VGND.n7663 VGND.n7662 4.6505
R21347 VGND.n7661 VGND.n7660 4.6505
R21348 VGND.n7658 VGND.n7657 4.6505
R21349 VGND.n7655 VGND.n7654 4.6505
R21350 VGND.n7652 VGND.n7651 4.6505
R21351 VGND.n7635 VGND.n7609 4.6505
R21352 VGND.n671 VGND.n670 4.6505
R21353 VGND.n659 VGND.n658 4.6505
R21354 VGND.n8243 VGND.n8242 4.6505
R21355 VGND.n8241 VGND.n8240 4.6505
R21356 VGND.n8237 VGND.n8236 4.6505
R21357 VGND.n8235 VGND.n8234 4.6505
R21358 VGND.n8233 VGND.n8232 4.6505
R21359 VGND.n8230 VGND.n8229 4.6505
R21360 VGND.n8223 VGND.n8222 4.6505
R21361 VGND.n8187 VGND.n8186 4.6505
R21362 VGND.n8184 VGND.n8183 4.6505
R21363 VGND.n8182 VGND.n8181 4.6505
R21364 VGND.n8178 VGND.n8177 4.6505
R21365 VGND.n8176 VGND.n8175 4.6505
R21366 VGND.n8173 VGND.n8172 4.6505
R21367 VGND.n8167 VGND.n8166 4.6505
R21368 VGND.n8163 VGND.n8162 4.6505
R21369 VGND.n8161 VGND.n8160 4.6505
R21370 VGND.n8262 VGND.n447 4.6505
R21371 VGND.n8283 VGND.n8282 4.6505
R21372 VGND.n8285 VGND.n8284 4.6505
R21373 VGND.n8289 VGND.n8288 4.6505
R21374 VGND.n8291 VGND.n8290 4.6505
R21375 VGND.n8293 VGND.n8292 4.6505
R21376 VGND.n8295 VGND.n8294 4.6505
R21377 VGND.n8297 VGND.n8296 4.6505
R21378 VGND.n8299 VGND.n8298 4.6505
R21379 VGND.n8302 VGND.n8301 4.6505
R21380 VGND.n8305 VGND.n8304 4.6505
R21381 VGND.n8308 VGND.n8307 4.6505
R21382 VGND.n380 VGND.n338 4.6505
R21383 VGND.n357 VGND.n356 4.6505
R21384 VGND.n355 VGND.n347 4.6505
R21385 VGND.n353 VGND.n348 4.6505
R21386 VGND.n379 VGND.n378 4.6505
R21387 VGND.n377 VGND.n376 4.6505
R21388 VGND.n374 VGND.n373 4.6505
R21389 VGND.n372 VGND.n371 4.6505
R21390 VGND.n370 VGND.n369 4.6505
R21391 VGND.n367 VGND.n366 4.6505
R21392 VGND.n362 VGND.n361 4.6505
R21393 VGND.n359 VGND.n358 4.6505
R21394 VGND.n330 VGND.n329 4.6505
R21395 VGND.n403 VGND.n402 4.6505
R21396 VGND.n400 VGND.n399 4.6505
R21397 VGND.n398 VGND.n397 4.6505
R21398 VGND.n395 VGND.n394 4.6505
R21399 VGND.n393 VGND.n392 4.6505
R21400 VGND.n390 VGND.n389 4.6505
R21401 VGND.n388 VGND.n387 4.6505
R21402 VGND.n386 VGND.n385 4.6505
R21403 VGND.n382 VGND.n381 4.6505
R21404 VGND.n8280 VGND.n8279 4.6505
R21405 VGND.n8278 VGND.n8277 4.6505
R21406 VGND.n8274 VGND.n8273 4.6505
R21407 VGND.n8269 VGND.n8268 4.6505
R21408 VGND.n8260 VGND.n8259 4.6505
R21409 VGND.n8245 VGND.n8244 4.6505
R21410 VGND.n8247 VGND.n8246 4.6505
R21411 VGND.n8250 VGND.n8249 4.6505
R21412 VGND.n8252 VGND.n8251 4.6505
R21413 VGND.n620 VGND.n619 4.6505
R21414 VGND.n623 VGND.n622 4.6505
R21415 VGND.n629 VGND.n628 4.6505
R21416 VGND.n631 VGND.n630 4.6505
R21417 VGND.n635 VGND.n634 4.6505
R21418 VGND.n639 VGND.n638 4.6505
R21419 VGND.n641 VGND.n640 4.6505
R21420 VGND.n644 VGND.n643 4.6505
R21421 VGND.n649 VGND.n648 4.6505
R21422 VGND.n653 VGND.n652 4.6505
R21423 VGND.n661 VGND.n660 4.6505
R21424 VGND.n665 VGND.n664 4.6505
R21425 VGND.n667 VGND.n666 4.6505
R21426 VGND.n676 VGND.n675 4.6505
R21427 VGND.n677 VGND.n606 4.6505
R21428 VGND.n679 VGND.n678 4.6505
R21429 VGND.n7637 VGND.n7636 4.6505
R21430 VGND.n7639 VGND.n7638 4.6505
R21431 VGND.n7641 VGND.n7640 4.6505
R21432 VGND.n7646 VGND.n7645 4.6505
R21433 VGND.n7648 VGND.n7647 4.6505
R21434 VGND.n7650 VGND.n7649 4.6505
R21435 VGND.n697 VGND.n696 4.6505
R21436 VGND.n701 VGND.n691 4.6505
R21437 VGND.n703 VGND.n702 4.6505
R21438 VGND.n706 VGND.n705 4.6505
R21439 VGND.n708 VGND.n707 4.6505
R21440 VGND.n712 VGND.n711 4.6505
R21441 VGND.n715 VGND.n714 4.6505
R21442 VGND.n7426 VGND.n7425 4.6505
R21443 VGND.n7355 VGND.n7354 4.6505
R21444 VGND.n7351 VGND.n810 4.6505
R21445 VGND.n7350 VGND.n811 4.6505
R21446 VGND.n7349 VGND.n813 4.6505
R21447 VGND.n7348 VGND.n815 4.6505
R21448 VGND.n7476 VGND.n7475 4.6505
R21449 VGND.n7479 VGND.n7478 4.6505
R21450 VGND.n7483 VGND.n7482 4.6505
R21451 VGND.n7424 VGND.n793 4.6505
R21452 VGND.n7422 VGND.n7421 4.6505
R21453 VGND.n7417 VGND.n7416 4.6505
R21454 VGND.n7414 VGND.n7413 4.6505
R21455 VGND.n7412 VGND.n7411 4.6505
R21456 VGND.n7410 VGND.n7409 4.6505
R21457 VGND.n7406 VGND.n7405 4.6505
R21458 VGND.n7404 VGND.n7403 4.6505
R21459 VGND.n7402 VGND.n7401 4.6505
R21460 VGND.n7398 VGND.n7397 4.6505
R21461 VGND.n7396 VGND.n7395 4.6505
R21462 VGND.n7393 VGND.n7392 4.6505
R21463 VGND.n7391 VGND.n807 4.6505
R21464 VGND.n7389 VGND.n7388 4.6505
R21465 VGND.n7385 VGND.n7384 4.6505
R21466 VGND.n7381 VGND.n7380 4.6505
R21467 VGND.n7379 VGND.n7378 4.6505
R21468 VGND.n7377 VGND.n7376 4.6505
R21469 VGND.n7375 VGND.n7374 4.6505
R21470 VGND.n7371 VGND.n7370 4.6505
R21471 VGND.n7369 VGND.n7368 4.6505
R21472 VGND.n7367 VGND.n7366 4.6505
R21473 VGND.n7365 VGND.n7364 4.6505
R21474 VGND.n7360 VGND.n7359 4.6505
R21475 VGND.n7357 VGND.n7356 4.6505
R21476 VGND.n1284 VGND.n1283 4.6505
R21477 VGND.n1278 VGND.n1151 4.6505
R21478 VGND.n1271 VGND.n887 4.6505
R21479 VGND.n1263 VGND.n1154 4.6505
R21480 VGND.n1260 VGND.n1259 4.6505
R21481 VGND.n1256 VGND.n1155 4.6505
R21482 VGND.n1242 VGND.n1240 4.6505
R21483 VGND.n1222 VGND.n1221 4.6505
R21484 VGND.n1219 VGND.n1161 4.6505
R21485 VGND.n1218 VGND.n1163 4.6505
R21486 VGND.n1294 VGND.n1293 4.6505
R21487 VGND.n1290 VGND.n1289 4.6505
R21488 VGND.n1288 VGND.n1147 4.6505
R21489 VGND.n1286 VGND.n1285 4.6505
R21490 VGND.n1255 VGND.n1254 4.6505
R21491 VGND.n1250 VGND.n1249 4.6505
R21492 VGND.n1214 VGND.n1213 4.6505
R21493 VGND.n985 VGND.n984 4.6505
R21494 VGND.n950 VGND.n917 4.6505
R21495 VGND.n937 VGND.n923 4.6505
R21496 VGND.n933 VGND.n928 4.6505
R21497 VGND.n934 VGND.n927 4.6505
R21498 VGND.n935 VGND.n925 4.6505
R21499 VGND.n939 VGND.n938 4.6505
R21500 VGND.n941 VGND.n940 4.6505
R21501 VGND.n942 VGND.n920 4.6505
R21502 VGND.n943 VGND.n919 4.6505
R21503 VGND.n945 VGND.n944 4.6505
R21504 VGND.n949 VGND.n948 4.6505
R21505 VGND.n952 VGND.n951 4.6505
R21506 VGND.n977 VGND.n976 4.6505
R21507 VGND.n975 VGND.n974 4.6505
R21508 VGND.n972 VGND.n971 4.6505
R21509 VGND.n970 VGND.n969 4.6505
R21510 VGND.n967 VGND.n966 4.6505
R21511 VGND.n962 VGND.n961 4.6505
R21512 VGND.n959 VGND.n958 4.6505
R21513 VGND.n956 VGND.n955 4.6505
R21514 VGND.n954 VGND.n953 4.6505
R21515 VGND.n1205 VGND.n1204 4.6505
R21516 VGND.n1209 VGND.n1208 4.6505
R21517 VGND.n1211 VGND.n1210 4.6505
R21518 VGND.n1217 VGND.n1216 4.6505
R21519 VGND.n1226 VGND.n1225 4.6505
R21520 VGND.n1230 VGND.n1229 4.6505
R21521 VGND.n1234 VGND.n1233 4.6505
R21522 VGND.n1238 VGND.n1237 4.6505
R21523 VGND.n1239 VGND.n1157 4.6505
R21524 VGND.n1244 VGND.n1243 4.6505
R21525 VGND.n1252 VGND.n1251 4.6505
R21526 VGND.n1258 VGND.n1257 4.6505
R21527 VGND.n1262 VGND.n1261 4.6505
R21528 VGND.n1265 VGND.n1264 4.6505
R21529 VGND.n1270 VGND.n1269 4.6505
R21530 VGND.n1273 VGND.n1272 4.6505
R21531 VGND.n1275 VGND.n1274 4.6505
R21532 VGND.n1277 VGND.n1276 4.6505
R21533 VGND.n1280 VGND.n1279 4.6505
R21534 VGND.n1282 VGND.n1281 4.6505
R21535 VGND.n1027 VGND.n1026 4.6505
R21536 VGND.n1029 VGND.n1028 4.6505
R21537 VGND.n1033 VGND.n1032 4.6505
R21538 VGND.n1035 VGND.n1034 4.6505
R21539 VGND.n1037 VGND.n1036 4.6505
R21540 VGND.n1039 VGND.n1038 4.6505
R21541 VGND.n1044 VGND.n1043 4.6505
R21542 VGND.n1046 VGND.n1045 4.6505
R21543 VGND.n1049 VGND.n1048 4.6505
R21544 VGND.n1051 VGND.n1050 4.6505
R21545 VGND.n1054 VGND.n1053 4.6505
R21546 VGND.n1056 VGND.n1055 4.6505
R21547 VGND.n1060 VGND.n1059 4.6505
R21548 VGND.n1064 VGND.n1063 4.6505
R21549 VGND.n1068 VGND.n1067 4.6505
R21550 VGND.n1070 VGND.n1069 4.6505
R21551 VGND.n1072 VGND.n1071 4.6505
R21552 VGND.n1077 VGND.n1076 4.6505
R21553 VGND.n1079 VGND.n1078 4.6505
R21554 VGND.n1083 VGND.n1082 4.6505
R21555 VGND.n1092 VGND.n1091 4.6505
R21556 VGND.n1095 VGND.n1094 4.6505
R21557 VGND.n1099 VGND.n1098 4.6505
R21558 VGND.n1100 VGND.n886 4.6505
R21559 VGND.n1105 VGND.n1104 4.6505
R21560 VGND.n1108 VGND.n1107 4.6505
R21561 VGND.n1111 VGND.n1110 4.6505
R21562 VGND.n1114 VGND.n1113 4.6505
R21563 VGND.n1116 VGND.n1004 4.6505
R21564 VGND.n1118 VGND.n1117 4.6505
R21565 VGND.n1121 VGND.n1120 4.6505
R21566 VGND.n1123 VGND.n1122 4.6505
R21567 VGND.n1125 VGND.n1124 4.6505
R21568 VGND.n1021 VGND.n1020 4.6505
R21569 VGND.n1025 VGND.n1024 4.6505
R21570 VGND.n7343 VGND.n7342 4.6505
R21571 VGND.n7345 VGND.n7344 4.6505
R21572 VGND.n7347 VGND.n7346 4.6505
R21573 VGND.n7353 VGND.n7352 4.6505
R21574 VGND.n7466 VGND.n7465 4.6505
R21575 VGND.n7469 VGND.n7468 4.6505
R21576 VGND.n7472 VGND.n7471 4.6505
R21577 VGND.n7477 VGND.n7454 4.6505
R21578 VGND.n7481 VGND.n7480 4.6505
R21579 VGND.n6454 VGND.n6341 4.6505
R21580 VGND.n6445 VGND.n6444 4.6505
R21581 VGND.n6433 VGND.n6343 4.6505
R21582 VGND.n6422 VGND.n6345 4.6505
R21583 VGND.n6394 VGND.n6347 4.6505
R21584 VGND.n6393 VGND.n6349 4.6505
R21585 VGND.n6392 VGND.n6350 4.6505
R21586 VGND.n6384 VGND.n6355 4.6505
R21587 VGND.n6220 VGND.n1692 4.6505
R21588 VGND.n6336 VGND.n6255 4.6505
R21589 VGND.n6122 VGND.n6121 4.6505
R21590 VGND.n6128 VGND.n6127 4.6505
R21591 VGND.n6134 VGND.n6133 4.6505
R21592 VGND.n6228 VGND.n6227 4.6505
R21593 VGND.n6232 VGND.n6231 4.6505
R21594 VGND.n6242 VGND.n6241 4.6505
R21595 VGND.n6299 VGND.n6298 4.6505
R21596 VGND.n6291 VGND.n6290 4.6505
R21597 VGND.n6288 VGND.n6287 4.6505
R21598 VGND.n6285 VGND.n6284 4.6505
R21599 VGND.n6451 VGND.n6450 4.6505
R21600 VGND.n6402 VGND.n6401 4.6505
R21601 VGND.n6857 VGND.n6856 4.6505
R21602 VGND.n1536 VGND.n1535 4.6505
R21603 VGND.n1533 VGND.n1532 4.6505
R21604 VGND.n1530 VGND.n1529 4.6505
R21605 VGND.n1526 VGND.n1525 4.6505
R21606 VGND.n1520 VGND.n1519 4.6505
R21607 VGND.n1512 VGND.n1511 4.6505
R21608 VGND.n1510 VGND.n1509 4.6505
R21609 VGND.n1507 VGND.n1506 4.6505
R21610 VGND.n1505 VGND.n1504 4.6505
R21611 VGND.n1503 VGND.n1502 4.6505
R21612 VGND.n1500 VGND.n1499 4.6505
R21613 VGND.n1498 VGND.n1497 4.6505
R21614 VGND.n1495 VGND.n1494 4.6505
R21615 VGND.n6966 VGND.n6965 4.6505
R21616 VGND.n6922 VGND.n6921 4.6505
R21617 VGND.n6920 VGND.n6919 4.6505
R21618 VGND.n6918 VGND.n6917 4.6505
R21619 VGND.n6914 VGND.n6913 4.6505
R21620 VGND.n6912 VGND.n6911 4.6505
R21621 VGND.n6909 VGND.n6908 4.6505
R21622 VGND.n6907 VGND.n6906 4.6505
R21623 VGND.n6901 VGND.n6900 4.6505
R21624 VGND.n6899 VGND.n6898 4.6505
R21625 VGND.n6897 VGND.n6896 4.6505
R21626 VGND.n6895 VGND.n1582 4.6505
R21627 VGND.n6865 VGND.n6864 4.6505
R21628 VGND.n6868 VGND.n6867 4.6505
R21629 VGND.n6870 VGND.n6869 4.6505
R21630 VGND.n6873 VGND.n6872 4.6505
R21631 VGND.n6876 VGND.n6875 4.6505
R21632 VGND.n6878 VGND.n6877 4.6505
R21633 VGND.n6882 VGND.n6881 4.6505
R21634 VGND.n6885 VGND.n6884 4.6505
R21635 VGND.n6889 VGND.n6888 4.6505
R21636 VGND.n6892 VGND.n6891 4.6505
R21637 VGND.n6894 VGND.n6893 4.6505
R21638 VGND.n6861 VGND.n6860 4.6505
R21639 VGND.n6834 VGND.n6833 4.6505
R21640 VGND.n6837 VGND.n6836 4.6505
R21641 VGND.n6841 VGND.n6840 4.6505
R21642 VGND.n6843 VGND.n6842 4.6505
R21643 VGND.n6847 VGND.n6846 4.6505
R21644 VGND.n6850 VGND.n6849 4.6505
R21645 VGND.n6854 VGND.n6853 4.6505
R21646 VGND.n6859 VGND.n6858 4.6505
R21647 VGND.n6827 VGND.n6826 4.6505
R21648 VGND.n1595 VGND.n1594 4.6505
R21649 VGND.n6362 VGND.n6361 4.6505
R21650 VGND.n6364 VGND.n6363 4.6505
R21651 VGND.n6368 VGND.n6367 4.6505
R21652 VGND.n6370 VGND.n6369 4.6505
R21653 VGND.n6372 VGND.n6371 4.6505
R21654 VGND.n6374 VGND.n6373 4.6505
R21655 VGND.n6376 VGND.n6375 4.6505
R21656 VGND.n6380 VGND.n6379 4.6505
R21657 VGND.n6383 VGND.n6382 4.6505
R21658 VGND.n6386 VGND.n6385 4.6505
R21659 VGND.n6391 VGND.n6390 4.6505
R21660 VGND.n6396 VGND.n6395 4.6505
R21661 VGND.n6404 VGND.n6403 4.6505
R21662 VGND.n6409 VGND.n6408 4.6505
R21663 VGND.n6411 VGND.n6410 4.6505
R21664 VGND.n6415 VGND.n6414 4.6505
R21665 VGND.n6419 VGND.n6418 4.6505
R21666 VGND.n6421 VGND.n6420 4.6505
R21667 VGND.n6424 VGND.n6423 4.6505
R21668 VGND.n6430 VGND.n6429 4.6505
R21669 VGND.n6432 VGND.n6431 4.6505
R21670 VGND.n6435 VGND.n6434 4.6505
R21671 VGND.n6441 VGND.n6440 4.6505
R21672 VGND.n6443 VGND.n6442 4.6505
R21673 VGND.n6447 VGND.n6446 4.6505
R21674 VGND.n6453 VGND.n6452 4.6505
R21675 VGND.n6279 VGND.n6278 4.6505
R21676 VGND.n6281 VGND.n6280 4.6505
R21677 VGND.n6283 VGND.n6282 4.6505
R21678 VGND.n6293 VGND.n6292 4.6505
R21679 VGND.n6304 VGND.n6303 4.6505
R21680 VGND.n6307 VGND.n6306 4.6505
R21681 VGND.n6309 VGND.n6308 4.6505
R21682 VGND.n6311 VGND.n6310 4.6505
R21683 VGND.n6314 VGND.n6313 4.6505
R21684 VGND.n6316 VGND.n6315 4.6505
R21685 VGND.n6318 VGND.n6317 4.6505
R21686 VGND.n6322 VGND.n6321 4.6505
R21687 VGND.n6324 VGND.n6323 4.6505
R21688 VGND.n6326 VGND.n6325 4.6505
R21689 VGND.n6329 VGND.n6328 4.6505
R21690 VGND.n6333 VGND.n6332 4.6505
R21691 VGND.n6335 VGND.n6334 4.6505
R21692 VGND.n6253 VGND.n6252 4.6505
R21693 VGND.n6245 VGND.n6244 4.6505
R21694 VGND.n6239 VGND.n6238 4.6505
R21695 VGND.n6222 VGND.n6221 4.6505
R21696 VGND.n6124 VGND.n6123 4.6505
R21697 VGND.n6130 VGND.n6129 4.6505
R21698 VGND.n6136 VGND.n6135 4.6505
R21699 VGND.n6138 VGND.n6137 4.6505
R21700 VGND.n6140 VGND.n6139 4.6505
R21701 VGND.n6145 VGND.n6144 4.6505
R21702 VGND.n6053 VGND.n6052 4.6505
R21703 VGND.n6026 VGND.n6019 4.6505
R21704 VGND.n6023 VGND.n6021 4.6505
R21705 VGND.n6583 VGND.n6582 4.6505
R21706 VGND.n1728 VGND.n1727 4.6505
R21707 VGND.n6628 VGND.n6627 4.6505
R21708 VGND.n6626 VGND.n6625 4.6505
R21709 VGND.n6622 VGND.n6621 4.6505
R21710 VGND.n6614 VGND.n6613 4.6505
R21711 VGND.n6611 VGND.n6610 4.6505
R21712 VGND.n6609 VGND.n6608 4.6505
R21713 VGND.n6607 VGND.n6606 4.6505
R21714 VGND.n6605 VGND.n6604 4.6505
R21715 VGND.n6603 VGND.n6602 4.6505
R21716 VGND.n6598 VGND.n6597 4.6505
R21717 VGND.n6638 VGND.n6637 4.6505
R21718 VGND.n6653 VGND.n6652 4.6505
R21719 VGND.n5284 VGND.n5224 4.6505
R21720 VGND.n5254 VGND.n5253 4.6505
R21721 VGND.n5252 VGND.n5232 4.6505
R21722 VGND.n5249 VGND.n5248 4.6505
R21723 VGND.n5246 VGND.n5245 4.6505
R21724 VGND.n5244 VGND.n5243 4.6505
R21725 VGND.n5242 VGND.n5241 4.6505
R21726 VGND.n5239 VGND.n5238 4.6505
R21727 VGND.n5283 VGND.n5282 4.6505
R21728 VGND.n5281 VGND.n5280 4.6505
R21729 VGND.n5279 VGND.n5278 4.6505
R21730 VGND.n5277 VGND.n5276 4.6505
R21731 VGND.n5275 VGND.n5274 4.6505
R21732 VGND.n5273 VGND.n5272 4.6505
R21733 VGND.n5271 VGND.n5270 4.6505
R21734 VGND.n5268 VGND.n5267 4.6505
R21735 VGND.n5266 VGND.n5265 4.6505
R21736 VGND.n5264 VGND.n5263 4.6505
R21737 VGND.n5262 VGND.n5261 4.6505
R21738 VGND.n5260 VGND.n5259 4.6505
R21739 VGND.n5258 VGND.n5257 4.6505
R21740 VGND.n5406 VGND.n5405 4.6505
R21741 VGND.n5409 VGND.n5408 4.6505
R21742 VGND.n5411 VGND.n5410 4.6505
R21743 VGND.n5413 VGND.n5412 4.6505
R21744 VGND.n5417 VGND.n5416 4.6505
R21745 VGND.n5421 VGND.n5420 4.6505
R21746 VGND.n5423 VGND.n5422 4.6505
R21747 VGND.n5427 VGND.n5426 4.6505
R21748 VGND.n5430 VGND.n5429 4.6505
R21749 VGND.n5432 VGND.n5431 4.6505
R21750 VGND.n5434 VGND.n5433 4.6505
R21751 VGND.n5437 VGND.n5436 4.6505
R21752 VGND.n5441 VGND.n5440 4.6505
R21753 VGND.n5446 VGND.n5445 4.6505
R21754 VGND.n5449 VGND.n5448 4.6505
R21755 VGND.n5379 VGND.n5378 4.6505
R21756 VGND.n5382 VGND.n5381 4.6505
R21757 VGND.n5384 VGND.n5383 4.6505
R21758 VGND.n5386 VGND.n5385 4.6505
R21759 VGND.n5391 VGND.n5390 4.6505
R21760 VGND.n5393 VGND.n5392 4.6505
R21761 VGND.n5395 VGND.n5394 4.6505
R21762 VGND.n5397 VGND.n5396 4.6505
R21763 VGND.n5400 VGND.n5399 4.6505
R21764 VGND.n5402 VGND.n5401 4.6505
R21765 VGND.n5404 VGND.n5403 4.6505
R21766 VGND.n6640 VGND.n6639 4.6505
R21767 VGND.n6642 VGND.n6641 4.6505
R21768 VGND.n6644 VGND.n6643 4.6505
R21769 VGND.n6649 VGND.n6648 4.6505
R21770 VGND.n6651 VGND.n6650 4.6505
R21771 VGND.n6655 VGND.n6654 4.6505
R21772 VGND.n6658 VGND.n6657 4.6505
R21773 VGND.n6660 VGND.n6659 4.6505
R21774 VGND.n6662 VGND.n6661 4.6505
R21775 VGND.n6672 VGND.n6671 4.6505
R21776 VGND.n6679 VGND.n6678 4.6505
R21777 VGND.n6682 VGND.n6681 4.6505
R21778 VGND.n6684 VGND.n6683 4.6505
R21779 VGND.n6687 VGND.n6686 4.6505
R21780 VGND.n6691 VGND.n6690 4.6505
R21781 VGND.n6695 VGND.n6694 4.6505
R21782 VGND.n6697 VGND.n6696 4.6505
R21783 VGND.n6699 VGND.n6698 4.6505
R21784 VGND.n6708 VGND.n6707 4.6505
R21785 VGND.n6710 VGND.n6709 4.6505
R21786 VGND.n6712 VGND.n6711 4.6505
R21787 VGND.n6714 VGND.n6713 4.6505
R21788 VGND.n6716 VGND.n6715 4.6505
R21789 VGND.n6719 VGND.n6718 4.6505
R21790 VGND.n6636 VGND.n6635 4.6505
R21791 VGND.n6577 VGND.n6576 4.6505
R21792 VGND.n6581 VGND.n6580 4.6505
R21793 VGND.n6585 VGND.n6584 4.6505
R21794 VGND.n6587 VGND.n6586 4.6505
R21795 VGND.n6589 VGND.n6588 4.6505
R21796 VGND.n6591 VGND.n6590 4.6505
R21797 VGND.n6593 VGND.n6592 4.6505
R21798 VGND.n6596 VGND.n6595 4.6505
R21799 VGND.n6020 VGND.n1637 4.6505
R21800 VGND.n6025 VGND.n6024 4.6505
R21801 VGND.n6030 VGND.n6029 4.6505
R21802 VGND.n6032 VGND.n6031 4.6505
R21803 VGND.n6033 VGND.n6018 4.6505
R21804 VGND.n6035 VGND.n6034 4.6505
R21805 VGND.n6037 VGND.n6036 4.6505
R21806 VGND.n6041 VGND.n6040 4.6505
R21807 VGND.n6047 VGND.n6046 4.6505
R21808 VGND.n6049 VGND.n6048 4.6505
R21809 VGND.n6051 VGND.n6050 4.6505
R21810 VGND.n1718 VGND.n1717 4.6505
R21811 VGND.n1721 VGND.n1720 4.6505
R21812 VGND.n1724 VGND.n1723 4.6505
R21813 VGND.n1729 VGND.n1706 4.6505
R21814 VGND.n1731 VGND.n1730 4.6505
R21815 VGND.n1734 VGND.n1733 4.6505
R21816 VGND.n1738 VGND.n1737 4.6505
R21817 VGND.n1820 VGND.n1819 4.6505
R21818 VGND.n1825 VGND.n1824 4.6505
R21819 VGND.n5940 VGND.n5939 4.6505
R21820 VGND.n5938 VGND.n1861 4.6505
R21821 VGND.n5935 VGND.n5109 4.6505
R21822 VGND.n5903 VGND.n5902 4.6505
R21823 VGND.n5899 VGND.n5112 4.6505
R21824 VGND.n5896 VGND.n5895 4.6505
R21825 VGND.n5500 VGND.n5123 4.6505
R21826 VGND.n5530 VGND.n5529 4.6505
R21827 VGND.n5535 VGND.n5534 4.6505
R21828 VGND.n5563 VGND.n5124 4.6505
R21829 VGND.n5573 VGND.n5572 4.6505
R21830 VGND.n5578 VGND.n5577 4.6505
R21831 VGND.n5583 VGND.n5582 4.6505
R21832 VGND.n5140 VGND.n5139 4.6505
R21833 VGND.n5142 VGND.n5141 4.6505
R21834 VGND.n5143 VGND.n5132 4.6505
R21835 VGND.n5145 VGND.n5144 4.6505
R21836 VGND.n5151 VGND.n5150 4.6505
R21837 VGND.n5156 VGND.n5155 4.6505
R21838 VGND.n5157 VGND.n5130 4.6505
R21839 VGND.n5159 VGND.n5158 4.6505
R21840 VGND.n5160 VGND.n5129 4.6505
R21841 VGND.n5162 VGND.n5161 4.6505
R21842 VGND.n5164 VGND.n5163 4.6505
R21843 VGND.n5166 VGND.n5165 4.6505
R21844 VGND.n5168 VGND.n5167 4.6505
R21845 VGND.n5170 VGND.n5169 4.6505
R21846 VGND.n5173 VGND.n5172 4.6505
R21847 VGND.n5175 VGND.n5174 4.6505
R21848 VGND.n5177 VGND.n5176 4.6505
R21849 VGND.n5179 VGND.n5178 4.6505
R21850 VGND.n5181 VGND.n5180 4.6505
R21851 VGND.n5183 VGND.n5182 4.6505
R21852 VGND.n5185 VGND.n5184 4.6505
R21853 VGND.n5801 VGND.n5800 4.6505
R21854 VGND.n5740 VGND.n5739 4.6505
R21855 VGND.n5737 VGND.n5736 4.6505
R21856 VGND.n5734 VGND.n5733 4.6505
R21857 VGND.n5732 VGND.n5731 4.6505
R21858 VGND.n5729 VGND.n5728 4.6505
R21859 VGND.n5727 VGND.n5726 4.6505
R21860 VGND.n5725 VGND.n5724 4.6505
R21861 VGND.n5722 VGND.n5721 4.6505
R21862 VGND.n5720 VGND.n5719 4.6505
R21863 VGND.n5717 VGND.n5716 4.6505
R21864 VGND.n5715 VGND.n5714 4.6505
R21865 VGND.n5713 VGND.n5712 4.6505
R21866 VGND.n5711 VGND.n5710 4.6505
R21867 VGND.n5709 VGND.n5708 4.6505
R21868 VGND.n5707 VGND.n5706 4.6505
R21869 VGND.n5705 VGND.n5704 4.6505
R21870 VGND.n5703 VGND.n5702 4.6505
R21871 VGND.n5700 VGND.n5699 4.6505
R21872 VGND.n5697 VGND.n5696 4.6505
R21873 VGND.n5694 VGND.n5693 4.6505
R21874 VGND.n5689 VGND.n5688 4.6505
R21875 VGND.n5686 VGND.n5685 4.6505
R21876 VGND.n5684 VGND.n5683 4.6505
R21877 VGND.n5681 VGND.n5680 4.6505
R21878 VGND.n5677 VGND.n5125 4.6505
R21879 VGND.n5676 VGND.n5675 4.6505
R21880 VGND.n5674 VGND.n5673 4.6505
R21881 VGND.n5671 VGND.n5670 4.6505
R21882 VGND.n5669 VGND.n5668 4.6505
R21883 VGND.n5666 VGND.n5665 4.6505
R21884 VGND.n5664 VGND.n5663 4.6505
R21885 VGND.n5662 VGND.n5661 4.6505
R21886 VGND.n5660 VGND.n5659 4.6505
R21887 VGND.n5657 VGND.n5656 4.6505
R21888 VGND.n5652 VGND.n5651 4.6505
R21889 VGND.n5649 VGND.n5648 4.6505
R21890 VGND.n5647 VGND.n5646 4.6505
R21891 VGND.n5502 VGND.n5501 4.6505
R21892 VGND.n5506 VGND.n5505 4.6505
R21893 VGND.n5509 VGND.n5508 4.6505
R21894 VGND.n5511 VGND.n5510 4.6505
R21895 VGND.n5513 VGND.n5512 4.6505
R21896 VGND.n5515 VGND.n5514 4.6505
R21897 VGND.n5517 VGND.n5516 4.6505
R21898 VGND.n5520 VGND.n5519 4.6505
R21899 VGND.n5522 VGND.n5521 4.6505
R21900 VGND.n5524 VGND.n5523 4.6505
R21901 VGND.n5526 VGND.n5525 4.6505
R21902 VGND.n5528 VGND.n5527 4.6505
R21903 VGND.n5532 VGND.n5531 4.6505
R21904 VGND.n5537 VGND.n5536 4.6505
R21905 VGND.n5539 VGND.n5538 4.6505
R21906 VGND.n5542 VGND.n5541 4.6505
R21907 VGND.n5544 VGND.n5543 4.6505
R21908 VGND.n5546 VGND.n5545 4.6505
R21909 VGND.n5548 VGND.n5547 4.6505
R21910 VGND.n5551 VGND.n5550 4.6505
R21911 VGND.n5562 VGND.n5561 4.6505
R21912 VGND.n5566 VGND.n5565 4.6505
R21913 VGND.n5568 VGND.n5567 4.6505
R21914 VGND.n5571 VGND.n5570 4.6505
R21915 VGND.n5575 VGND.n5574 4.6505
R21916 VGND.n5580 VGND.n5579 4.6505
R21917 VGND.n5585 VGND.n5584 4.6505
R21918 VGND.n5588 VGND.n5587 4.6505
R21919 VGND.n5968 VGND.n5967 4.6505
R21920 VGND.n5966 VGND.n5965 4.6505
R21921 VGND.n5964 VGND.n5963 4.6505
R21922 VGND.n5961 VGND.n5960 4.6505
R21923 VGND.n5959 VGND.n5958 4.6505
R21924 VGND.n5957 VGND.n5956 4.6505
R21925 VGND.n5955 VGND.n5954 4.6505
R21926 VGND.n5953 VGND.n5952 4.6505
R21927 VGND.n5951 VGND.n5950 4.6505
R21928 VGND.n5948 VGND.n5947 4.6505
R21929 VGND.n5946 VGND.n5945 4.6505
R21930 VGND.n5944 VGND.n5943 4.6505
R21931 VGND.n5942 VGND.n5941 4.6505
R21932 VGND.n5937 VGND.n5936 4.6505
R21933 VGND.n5934 VGND.n5933 4.6505
R21934 VGND.n5932 VGND.n5931 4.6505
R21935 VGND.n5930 VGND.n5929 4.6505
R21936 VGND.n5928 VGND.n5927 4.6505
R21937 VGND.n5925 VGND.n5924 4.6505
R21938 VGND.n5923 VGND.n5922 4.6505
R21939 VGND.n5921 VGND.n5920 4.6505
R21940 VGND.n5919 VGND.n5918 4.6505
R21941 VGND.n5917 VGND.n5916 4.6505
R21942 VGND.n5915 VGND.n5914 4.6505
R21943 VGND.n5913 VGND.n5912 4.6505
R21944 VGND.n5911 VGND.n5910 4.6505
R21945 VGND.n5908 VGND.n5907 4.6505
R21946 VGND.n5905 VGND.n5904 4.6505
R21947 VGND.n5901 VGND.n5900 4.6505
R21948 VGND.n5898 VGND.n5897 4.6505
R21949 VGND.n5894 VGND.n5893 4.6505
R21950 VGND.n1807 VGND.n1806 4.6505
R21951 VGND.n1810 VGND.n1809 4.6505
R21952 VGND.n1812 VGND.n1811 4.6505
R21953 VGND.n1815 VGND.n1814 4.6505
R21954 VGND.n1817 VGND.n1816 4.6505
R21955 VGND.n1821 VGND.n1797 4.6505
R21956 VGND.n1823 VGND.n1822 4.6505
R21957 VGND.n2482 VGND.n2338 4.6505
R21958 VGND.n2472 VGND.n2471 4.6505
R21959 VGND.n2456 VGND.n20 4.6505
R21960 VGND.n2418 VGND.n2417 4.6505
R21961 VGND.n2416 VGND.n2353 4.6505
R21962 VGND.n2415 VGND.n2354 4.6505
R21963 VGND.n2412 VGND.n2411 4.6505
R21964 VGND.n2409 VGND.n2357 4.6505
R21965 VGND.n2571 VGND.n19 4.6505
R21966 VGND.n2560 VGND.n2559 4.6505
R21967 VGND.n2548 VGND.n2310 4.6505
R21968 VGND.n9183 VGND.n16 4.6505
R21969 VGND.n3490 VGND.n3489 4.6505
R21970 VGND.n3496 VGND.n3495 4.6505
R21971 VGND.n3502 VGND.n3501 4.6505
R21972 VGND.n3506 VGND.n3505 4.6505
R21973 VGND.n3509 VGND.n3508 4.6505
R21974 VGND.n9201 VGND.n9200 4.6505
R21975 VGND.n9197 VGND.n9196 4.6505
R21976 VGND.n9195 VGND.n9194 4.6505
R21977 VGND.n9193 VGND.n9192 4.6505
R21978 VGND.n9191 VGND.n9190 4.6505
R21979 VGND.n9186 VGND.n9185 4.6505
R21980 VGND.n2186 VGND.n2185 4.6505
R21981 VGND.n2189 VGND.n2188 4.6505
R21982 VGND.n2191 VGND.n2190 4.6505
R21983 VGND.n2193 VGND.n2192 4.6505
R21984 VGND.n2196 VGND.n2195 4.6505
R21985 VGND.n2200 VGND.n2199 4.6505
R21986 VGND.n2203 VGND.n2202 4.6505
R21987 VGND.n2205 VGND.n2204 4.6505
R21988 VGND.n2208 VGND.n2207 4.6505
R21989 VGND.n2212 VGND.n2211 4.6505
R21990 VGND.n2215 VGND.n2214 4.6505
R21991 VGND.n2217 VGND.n2216 4.6505
R21992 VGND.n2220 VGND.n2219 4.6505
R21993 VGND.n2223 VGND.n2172 4.6505
R21994 VGND.n2225 VGND.n2224 4.6505
R21995 VGND.n2229 VGND.n2228 4.6505
R21996 VGND.n2232 VGND.n2231 4.6505
R21997 VGND.n2620 VGND.n2619 4.6505
R21998 VGND.n2616 VGND.n2615 4.6505
R21999 VGND.n2612 VGND.n2611 4.6505
R22000 VGND.n2610 VGND.n2609 4.6505
R22001 VGND.n2608 VGND.n2607 4.6505
R22002 VGND.n2605 VGND.n2604 4.6505
R22003 VGND.n2603 VGND.n2602 4.6505
R22004 VGND.n2600 VGND.n2599 4.6505
R22005 VGND.n2598 VGND.n2597 4.6505
R22006 VGND.n2593 VGND.n2592 4.6505
R22007 VGND.n2591 VGND.n2590 4.6505
R22008 VGND.n2588 VGND.n2587 4.6505
R22009 VGND.n2585 VGND.n2584 4.6505
R22010 VGND.n2583 VGND.n2297 4.6505
R22011 VGND.n2580 VGND.n2579 4.6505
R22012 VGND.n2479 VGND.n2478 4.6505
R22013 VGND.n2452 VGND.n2451 4.6505
R22014 VGND.n2403 VGND.n2402 4.6505
R22015 VGND.n2408 VGND.n2407 4.6505
R22016 VGND.n2410 VGND.n2355 4.6505
R22017 VGND.n2414 VGND.n2413 4.6505
R22018 VGND.n2420 VGND.n2419 4.6505
R22019 VGND.n2423 VGND.n2422 4.6505
R22020 VGND.n2426 VGND.n2425 4.6505
R22021 VGND.n2428 VGND.n2427 4.6505
R22022 VGND.n2430 VGND.n2429 4.6505
R22023 VGND.n2432 VGND.n2431 4.6505
R22024 VGND.n2436 VGND.n2435 4.6505
R22025 VGND.n2438 VGND.n2437 4.6505
R22026 VGND.n2440 VGND.n2439 4.6505
R22027 VGND.n2442 VGND.n2441 4.6505
R22028 VGND.n2444 VGND.n2443 4.6505
R22029 VGND.n2447 VGND.n2446 4.6505
R22030 VGND.n2450 VGND.n2449 4.6505
R22031 VGND.n2455 VGND.n2454 4.6505
R22032 VGND.n2458 VGND.n2457 4.6505
R22033 VGND.n2460 VGND.n2459 4.6505
R22034 VGND.n2462 VGND.n2461 4.6505
R22035 VGND.n2468 VGND.n2467 4.6505
R22036 VGND.n2470 VGND.n2469 4.6505
R22037 VGND.n2477 VGND.n2476 4.6505
R22038 VGND.n2481 VGND.n2480 4.6505
R22039 VGND.n2484 VGND.n2483 4.6505
R22040 VGND.n2545 VGND.n2544 4.6505
R22041 VGND.n2547 VGND.n2546 4.6505
R22042 VGND.n2550 VGND.n2549 4.6505
R22043 VGND.n2554 VGND.n2553 4.6505
R22044 VGND.n2558 VGND.n2557 4.6505
R22045 VGND.n2562 VGND.n2561 4.6505
R22046 VGND.n2567 VGND.n2566 4.6505
R22047 VGND.n2570 VGND.n2569 4.6505
R22048 VGND VGND.n2305 4.6505
R22049 VGND.n2574 VGND.n2573 4.6505
R22050 VGND.n3492 VGND.n3491 4.6505
R22051 VGND.n3498 VGND.n3497 4.6505
R22052 VGND.n3504 VGND.n3503 4.6505
R22053 VGND.n3507 VGND.n3484 4.6505
R22054 VGND.n9163 VGND.n9162 4.6505
R22055 VGND.n9160 VGND.n9159 4.6505
R22056 VGND.n9155 VGND.n9154 4.6505
R22057 VGND.n9152 VGND.n9151 4.6505
R22058 VGND.n9149 VGND.n9148 4.6505
R22059 VGND.n9147 VGND.n9104 4.6505
R22060 VGND.n9146 VGND.n9145 4.6505
R22061 VGND.n9144 VGND.n9105 4.6505
R22062 VGND.n9143 VGND.n9142 4.6505
R22063 VGND.n9140 VGND.n9139 4.6505
R22064 VGND.n9138 VGND.n9137 4.6505
R22065 VGND.n9136 VGND.n9110 4.6505
R22066 VGND.n9135 VGND.n9134 4.6505
R22067 VGND.n9133 VGND.n9111 4.6505
R22068 VGND.n9132 VGND.n9131 4.6505
R22069 VGND.n9130 VGND.n9112 4.6505
R22070 VGND.n9129 VGND.n9128 4.6505
R22071 VGND.n9127 VGND.n9115 4.6505
R22072 VGND.n9126 VGND.n9117 4.6505
R22073 VGND.n9125 VGND.n9124 4.6505
R22074 VGND.n9123 VGND.n9118 4.6505
R22075 VGND.n2596 VGND.n2595 4.63943
R22076 VGND.n5374 VGND.n5341 4.63943
R22077 VGND.n6675 VGND.n6674 4.63943
R22078 VGND.n5453 VGND.n5450 4.6085
R22079 VGND.n2597 VGND.n2596 4.60638
R22080 VGND.n2924 VGND.n2923 4.5918
R22081 VGND.n4863 VGND.n4862 4.57427
R22082 VGND.n5097 VGND.n5096 4.57427
R22083 VGND.n7220 VGND.n7219 4.57427
R22084 VGND.n4810 VGND.n4809 4.57427
R22085 VGND.n4963 VGND.n4962 4.57427
R22086 VGND.n4512 VGND.n4511 4.57427
R22087 VGND.n6981 VGND.n6980 4.57427
R22088 VGND.n4716 VGND.n4715 4.57427
R22089 VGND.n4152 VGND.n4151 4.57427
R22090 VGND.n4304 VGND.n4303 4.57427
R22091 VGND.n3577 VGND.n3576 4.57427
R22092 VGND.n2894 VGND.n2664 4.57427
R22093 VGND.n2774 VGND.n2773 4.57427
R22094 VGND.n3458 VGND.n3457 4.57427
R22095 VGND.n3381 VGND.n3380 4.57427
R22096 VGND.n3708 VGND.n3707 4.57427
R22097 VGND.n3200 VGND.n3199 4.57427
R22098 VGND.n9043 VGND.n9042 4.57427
R22099 VGND.n8859 VGND.n8858 4.57427
R22100 VGND.n3841 VGND.n3840 4.57427
R22101 VGND.n305 VGND.n304 4.57427
R22102 VGND.n8704 VGND.n8703 4.57427
R22103 VGND.n3818 VGND.n3817 4.57427
R22104 VGND.n3918 VGND.n3917 4.57427
R22105 VGND.n8428 VGND.n8339 4.57427
R22106 VGND.n8089 VGND.n8088 4.57427
R22107 VGND.n1971 VGND.n1970 4.57427
R22108 VGND.n1990 VGND.n1989 4.57427
R22109 VGND.n7761 VGND.n7760 4.57427
R22110 VGND.n7560 VGND.n7559 4.57427
R22111 VGND.n8334 VGND.n8333 4.57427
R22112 VGND.n8195 VGND.n8143 4.57427
R22113 VGND.n7537 VGND.n7536 4.57427
R22114 VGND.n7633 VGND.n7632 4.57427
R22115 VGND.n7428 VGND.n7427 4.57427
R22116 VGND.n1315 VGND.n1314 4.57427
R22117 VGND.n7310 VGND.n7309 4.57427
R22118 VGND.n778 VGND.n777 4.57427
R22119 VGND.n7340 VGND.n7339 4.57427
R22120 VGND.n6214 VGND.n6213 4.57427
R22121 VGND.n6975 VGND.n6974 4.57427
R22122 VGND.n6817 VGND.n6816 4.57427
R22123 VGND.n6276 VGND.n6264 4.57427
R22124 VGND.n6110 VGND.n6109 4.57427
R22125 VGND.n6574 VGND.n1653 4.57427
R22126 VGND.n5366 VGND.n5365 4.57427
R22127 VGND.n6055 VGND.n6054 4.57427
R22128 VGND.n1761 VGND.n1760 4.57427
R22129 VGND.n5810 VGND.n5809 4.57427
R22130 VGND.n5637 VGND.n5636 4.57427
R22131 VGND.n5891 VGND.n5115 4.57427
R22132 VGND.n5972 VGND.n5971 4.57427
R22133 VGND.n1840 VGND.n1839 4.57427
R22134 VGND.n2244 VGND.n2243 4.57427
R22135 VGND.n9177 VGND.n9176 4.57427
R22136 VGND.n2511 VGND.n2510 4.57427
R22137 VGND.n3524 VGND.n3523 4.57427
R22138 VGND.n4377 VGND.n4168 4.57412
R22139 VGND.n8785 VGND.n8784 4.57412
R22140 VGND.n6456 VGND.n6455 4.57412
R22141 VGND.n2623 VGND.n18 4.57412
R22142 VGND.n5012 VGND.n3986 4.57412
R22143 VGND.n3327 VGND.n2644 4.57412
R22144 VGND.n8911 VGND.n8910 4.57412
R22145 VGND.n5816 VGND.n5815 4.57412
R22146 VGND.n5209 VGND.n5208 4.5622
R22147 VGND.n1436 VGND.n1435 4.5622
R22148 VGND.n8586 VGND.n8585 4.5622
R22149 VGND.n1525 VGND.n1524 4.5622
R22150 VGND.n9200 VGND.n9198 4.55559
R22151 VGND.n6707 VGND.n6705 4.55559
R22152 VGND.n6613 VGND.n1640 4.55559
R22153 VGND.n3444 VGND.n3442 4.55559
R22154 VGND.n1519 VGND.n1515 4.55559
R22155 VGND.n1747 VGND.n1746 4.53348
R22156 VGND.n4798 VGND.n4764 4.53348
R22157 VGND.n1915 VGND.n1876 4.53348
R22158 VGND.n7527 VGND.n7526 4.53348
R22159 VGND.n6017 VGND.n6016 4.5303
R22160 VGND.n803 VGND.n802 4.5303
R22161 VGND.n6219 VGND.n6218 4.5303
R22162 VGND.n4420 VGND.n4220 4.51815
R22163 VGND.n8341 VGND.n8340 4.51815
R22164 VGND.n491 VGND.n490 4.51815
R22165 VGND.n638 VGND.n637 4.51815
R22166 VGND.n1225 VGND.n1224 4.51815
R22167 VGND.n1059 VGND.n1058 4.51815
R22168 VGND.n6429 VGND.n6426 4.51815
R22169 VGND.n6418 VGND.n6417 4.51815
R22170 VGND.n3926 VGND.n3887 4.51198
R22171 VGND.n4989 VGND.n4988 4.5005
R22172 VGND.n4338 VGND.n4337 4.5005
R22173 VGND.n8799 VGND.n8798 4.5005
R22174 VGND.n565 VGND.n564 4.5005
R22175 VGND.n7703 VGND.n7702 4.5005
R22176 VGND.n883 VGND.n882 4.5005
R22177 VGND.n6515 VGND.n6514 4.5005
R22178 VGND.n5863 VGND.n5862 4.5005
R22179 VGND.n2282 VGND.n2281 4.5005
R22180 VGND.n1585 VGND.n1584 4.47602
R22181 VGND.n5371 VGND.n5341 4.454
R22182 VGND.n2402 VGND.n2401 4.45267
R22183 VGND.n8900 VGND.n84 4.43378
R22184 VGND.n8580 VGND.n8579 4.43256
R22185 VGND.n6696 VGND.n1623 4.42603
R22186 VGND.n1314 VGND.n1311 4.41955
R22187 VGND.n2287 VGND.n2286 4.36875
R22188 VGND.n2171 VGND.n2170 4.36875
R22189 VGND.n2175 VGND.n2174 4.36875
R22190 VGND.n15 VGND.n14 4.36875
R22191 VGND.n5200 VGND.n5199 4.36875
R22192 VGND.n2106 VGND.n2105 4.36875
R22193 VGND.n2117 VGND.n2116 4.36875
R22194 VGND.n2121 VGND.n2120 4.36875
R22195 VGND.n3310 VGND.n3309 4.36875
R22196 VGND.n3661 VGND.n3660 4.36875
R22197 VGND.n3636 VGND.n3635 4.36875
R22198 VGND.n192 VGND.n191 4.36875
R22199 VGND.n1518 VGND.n1517 4.36875
R22200 VGND.n242 VGND.n241 4.35795
R22201 VGND.n689 VGND.n688 4.35795
R22202 VGND.n907 VGND.n906 4.35795
R22203 VGND.n1086 VGND.n1085 4.35795
R22204 VGND.n6700 VGND.n6699 4.28986
R22205 VGND.n4428 VGND.n4219 4.28986
R22206 VGND.n8581 VGND.n246 4.28986
R22207 VGND.n8385 VGND.n8384 4.28986
R22208 VGND.n8266 VGND.n447 4.28986
R22209 VGND.n6233 VGND.n6232 4.28986
R22210 VGND.n6239 VGND.n1691 4.28986
R22211 VGND.n9164 VGND.n9163 4.28986
R22212 VGND.n970 VGND.n913 4.22178
R22213 VGND.n9163 VGND.n27 4.22178
R22214 VGND.n1146 VGND.n1145 4.21637
R22215 VGND.n4957 VGND.n4956 4.18553
R22216 VGND.n1465 VGND.n1464 4.14168
R22217 VGND.n2982 VGND.n2981 4.14168
R22218 VGND.n8625 VGND.n220 4.14168
R22219 VGND.n8358 VGND.n8352 4.14168
R22220 VGND.n7958 VGND.n7957 4.14168
R22221 VGND.n923 VGND.n921 4.14168
R22222 VGND.n6965 VGND.n6964 4.14168
R22223 VGND.n6440 VGND.n6439 4.14168
R22224 VGND.n2425 VGND.n2424 4.11798
R22225 VGND.n2231 VGND.n2230 4.11798
R22226 VGND.n5172 VGND.n5171 4.11798
R22227 VGND.n5719 VGND.n5718 4.11798
R22228 VGND.n5519 VGND.n5518 4.11798
R22229 VGND.n5910 VGND.n5909 4.11798
R22230 VGND.n5950 VGND.n5949 4.11798
R22231 VGND.n5443 VGND.n5442 4.11798
R22232 VGND.n5390 VGND.n5389 4.11798
R22233 VGND.n7028 VGND.n7027 4.11798
R22234 VGND.n7054 VGND.n7053 4.11798
R22235 VGND.n4939 VGND.n4938 4.11798
R22236 VGND.n4268 VGND.n4267 4.11798
R22237 VGND.n4539 VGND.n4538 4.11798
R22238 VGND.n4541 VGND.n4539 4.11798
R22239 VGND.n3288 VGND.n2655 4.11798
R22240 VGND.n2655 VGND.n2654 4.11798
R22241 VGND.n3095 VGND.n3094 4.11798
R22242 VGND.n92 VGND.n91 4.11798
R22243 VGND.n9002 VGND.n9001 4.11798
R22244 VGND.n3865 VGND.n3864 4.11798
R22245 VGND.n7822 VGND.n7821 4.11798
R22246 VGND.n7823 VGND.n7822 4.11798
R22247 VGND.n393 VGND.n335 4.11798
R22248 VGND.n7574 VGND.n7573 4.11798
R22249 VGND.n7576 VGND.n7574 4.11798
R22250 VGND.n7657 VGND.n7656 4.11798
R22251 VGND.n8170 VGND.n8169 4.11798
R22252 VGND.n8301 VGND.n8300 4.11798
R22253 VGND.n7364 VGND.n7361 4.11798
R22254 VGND.n7395 VGND.n7394 4.11798
R22255 VGND.n7394 VGND.n7393 4.11798
R22256 VGND.n6884 VGND.n6883 4.11798
R22257 VGND.n6849 VGND.n6848 4.11798
R22258 VGND.n6313 VGND.n6312 4.11798
R22259 VGND.n1594 VGND.n1593 4.11798
R22260 VGND.n6617 VGND.n6616 4.09013
R22261 VGND.n9 VGND.n8 4.07323
R22262 VGND.n5148 VGND.n5147 4.07323
R22263 VGND.n4431 VGND.n4219 4.07323
R22264 VGND.n4435 VGND.n4431 4.07323
R22265 VGND.n1401 VGND.n1400 4.07323
R22266 VGND.n1399 VGND.n1396 4.07323
R22267 VGND.n2879 VGND.n2878 4.07323
R22268 VGND.n2674 VGND.n2673 4.07323
R22269 VGND.n8969 VGND.n8968 4.07323
R22270 VGND.n246 VGND.n245 4.07323
R22271 VGND.n1927 VGND.n1923 4.07323
R22272 VGND.n1923 VGND.n1922 4.07323
R22273 VGND.n1482 VGND.n1481 4.07323
R22274 VGND.n9167 VGND.n9164 4.07323
R22275 VGND.n9167 VGND.n9166 4.07323
R22276 VGND.n6688 VGND.n6687 4.03876
R22277 VGND.n3457 VGND.n3456 4.03876
R22278 VGND.n7675 VGND.n684 4.03876
R22279 VGND.n9184 VGND.n9183 3.97459
R22280 VGND.n3428 VGND.n3427 3.97459
R22281 VGND.n2294 VGND.n2293 3.96548
R22282 VGND.n2177 VGND.n2176 3.96548
R22283 VGND.n5230 VGND.n5229 3.96548
R22284 VGND.n5202 VGND.n5201 3.96548
R22285 VGND.n1626 VGND.n1625 3.96548
R22286 VGND.n2112 VGND.n2111 3.96548
R22287 VGND.n3063 VGND.n3062 3.96548
R22288 VGND.n95 VGND.n94 3.96548
R22289 VGND.n186 VGND.n185 3.96548
R22290 VGND.n7677 VGND.n7676 3.96548
R22291 VGND.n5365 VGND.n5364 3.9624
R22292 VGND.n1314 VGND.n1313 3.9624
R22293 VGND.n3069 VGND.n3033 3.96015
R22294 VGND.n5444 VGND.n5443 3.93896
R22295 VGND.n8264 VGND.n448 3.90948
R22296 VGND.n1292 VGND.n1291 3.88508
R22297 VGND.n165 VGND.n164 3.88135
R22298 VGND.n8647 VGND.n8646 3.83619
R22299 VGND.n3797 VGND.n3796 3.82659
R22300 VGND.n6045 VGND.n6044 3.79309
R22301 VGND.n7143 VGND.n7142 3.76521
R22302 VGND.n4019 VGND.n4018 3.76521
R22303 VGND.n5020 VGND.n5019 3.76521
R22304 VGND.n2675 VGND.n2674 3.76521
R22305 VGND.n8970 VGND.n8969 3.76521
R22306 VGND.n8052 VGND.n488 3.76521
R22307 VGND.n335 VGND.n334 3.75994
R22308 VGND.n6832 VGND.n6831 3.75994
R22309 VGND.n8891 VGND.n8890 3.7575
R22310 VGND.n5231 VGND.n5230 3.7069
R22311 VGND.n5203 VGND.n5202 3.7069
R22312 VGND.n1627 VGND.n1626 3.7069
R22313 VGND.n2113 VGND.n2112 3.7069
R22314 VGND.n3322 VGND.n3321 3.7069
R22315 VGND.n3321 VGND.n3320 3.7069
R22316 VGND.n96 VGND.n95 3.7069
R22317 VGND.n528 VGND.n527 3.7069
R22318 VGND.n7678 VGND.n7677 3.7069
R22319 VGND.n3694 VGND.n3693 3.6638
R22320 VGND.n5210 VGND.n5209 3.62403
R22321 VGND.n493 VGND.n492 3.61789
R22322 VGND.n5420 VGND.n5418 3.59021
R22323 VGND.n3422 VGND.n3420 3.59021
R22324 VGND.n8877 VGND.n93 3.59021
R22325 VGND.n4631 VGND.n4630 3.54093
R22326 VGND.n3707 VGND.n3706 3.53451
R22327 VGND.n2575 VGND.n2574 3.50735
R22328 VGND.n2725 VGND.n2667 3.50735
R22329 VGND.n8604 VGND.n232 3.50735
R22330 VGND.n7865 VGND.n7864 3.50735
R22331 VGND.n1088 VGND.n1087 3.50735
R22332 VGND.n6245 VGND.n1689 3.50735
R22333 VGND.n179 VGND.n177 3.50486
R22334 VGND.n535 VGND.n534 3.49538
R22335 VGND.n4435 VGND.n4434 3.47876
R22336 VGND.n1927 VGND.n1926 3.47876
R22337 VGND.n6666 VGND.n6665 3.44377
R22338 VGND.n2800 VGND.n2799 3.44377
R22339 VGND.n7853 VGND.n7852 3.44377
R22340 VGND.n4815 VGND.n4814 3.4105
R22341 VGND VGND.n4843 3.4105
R22342 VGND.n7074 VGND.n7073 3.4105
R22343 VGND.n7085 VGND.n7084 3.4105
R22344 VGND.n7096 VGND.n7095 3.4105
R22345 VGND.n4807 VGND.n4806 3.4105
R22346 VGND.n5009 VGND.n5008 3.4105
R22347 VGND.n4569 VGND.n1388 3.4105
R22348 VGND.n4135 VGND.n4134 3.4105
R22349 VGND.n4733 VGND 3.4105
R22350 VGND.n4158 VGND.n4157 3.4105
R22351 VGND.n4353 VGND.n4352 3.4105
R22352 VGND.n4374 VGND.n4373 3.4105
R22353 VGND.n2084 VGND.n2083 3.4105
R22354 VGND VGND.n3559 3.4105
R22355 VGND.n9075 VGND.n9074 3.4105
R22356 VGND.n3005 VGND.n3004 3.4105
R22357 VGND.n2770 VGND.n2769 3.4105
R22358 VGND.n3462 VGND.n3461 3.4105
R22359 VGND.n3331 VGND.n3330 3.4105
R22360 VGND.n3160 VGND.n3159 3.4105
R22361 VGND.n131 VGND.n130 3.4105
R22362 VGND.n8695 VGND.n8694 3.4105
R22363 VGND.n8529 VGND.n8528 3.4105
R22364 VGND.n8544 VGND.n8543 3.4105
R22365 VGND.n8789 VGND.n8788 3.4105
R22366 VGND.n1995 VGND.n1994 3.4105
R22367 VGND.n7979 VGND.n299 3.4105
R22368 VGND.n568 VGND.n567 3.4105
R22369 VGND.n429 VGND.n428 3.4105
R22370 VGND.n8330 VGND.n8329 3.4105
R22371 VGND.n409 VGND.n408 3.4105
R22372 VGND.n8138 VGND.n8137 3.4105
R22373 VGND.n8206 VGND.n8205 3.4105
R22374 VGND.n7693 VGND.n7692 3.4105
R22375 VGND.n7494 VGND.n7493 3.4105
R22376 VGND.n7446 VGND 3.4105
R22377 VGND.n7306 VGND.n7305 3.4105
R22378 VGND.n1183 VGND.n1182 3.4105
R22379 VGND.n785 VGND.n784 3.4105
R22380 VGND.n7323 VGND.n7322 3.4105
R22381 VGND.n6156 VGND.n6155 3.4105
R22382 VGND VGND.n6170 3.4105
R22383 VGND.n6189 VGND.n6188 3.4105
R22384 VGND.n6944 VGND.n1578 3.4105
R22385 VGND.n6113 VGND.n6112 3.4105
R22386 VGND.n6217 VGND.n6216 3.4105
R22387 VGND.n6467 VGND.n6466 3.4105
R22388 VGND.n1756 VGND.n1755 3.4105
R22389 VGND.n6519 VGND.n6518 3.4105
R22390 VGND.n5289 VGND.n5288 3.4105
R22391 VGND.n5330 VGND.n5329 3.4105
R22392 VGND.n5988 VGND.n5987 3.4105
R22393 VGND.n5765 VGND.n5467 3.4105
R22394 VGND.n5860 VGND.n5859 3.4105
R22395 VGND.n9216 VGND.n9215 3.4105
R22396 VGND.n2379 VGND.n2378 3.4105
R22397 VGND.n3528 VGND.n3527 3.4105
R22398 VGND.n2627 VGND.n2626 3.4105
R22399 VGND.n2435 VGND.n2434 3.4019
R22400 VGND.n7009 VGND.n7008 3.4019
R22401 VGND.n4928 VGND.n4927 3.4019
R22402 VGND.n4259 VGND.n4258 3.4019
R22403 VGND.n3109 VGND.n3108 3.4019
R22404 VGND.n8993 VGND.n8992 3.4019
R22405 VGND.n8288 VGND.n8287 3.4019
R22406 VGND.n7364 VGND.n7363 3.4019
R22407 VGND.n6321 VGND.n6320 3.4019
R22408 VGND.n7201 VGND.n7200 3.38874
R22409 VGND.n2933 VGND.n2900 3.38874
R22410 VGND.n8493 VGND.n8452 3.38874
R22411 VGND.n8053 VGND.n8052 3.38874
R22412 VGND.n7832 VGND.n7831 3.38874
R22413 VGND.n657 VGND.n656 3.38874
R22414 VGND.n1102 VGND.n886 3.38874
R22415 VGND.n1022 VGND.n1021 3.38874
R22416 VGND.n3576 VGND.n3575 3.36212
R22417 VGND.n8933 VGND.n8932 3.33201
R22418 VGND.n214 VGND.n213 3.33201
R22419 VGND.n5076 VGND 3.29747
R22420 VGND.n8171 VGND.n8170 3.22288
R22421 VGND.n1586 VGND.n1585 3.22288
R22422 VGND.n4962 VGND.n4961 3.21921
R22423 VGND.n2801 VGND.n2800 3.21921
R22424 VGND.n7854 VGND.n7853 3.21921
R22425 VGND.n5558 VGND.n5557 3.2005
R22426 VGND.n4562 VGND.n4561 3.2005
R22427 VGND.n2815 VGND.n2755 3.2005
R22428 VGND.n3219 VGND.n3218 3.2005
R22429 VGND.n8930 VGND.n8927 3.2005
R22430 VGND.n252 VGND.n251 3.2005
R22431 VGND.n8603 VGND.n8600 3.2005
R22432 VGND.n211 VGND.n208 3.2005
R22433 VGND.n514 VGND.n513 3.2005
R22434 VGND.n7898 VGND.n7897 3.2005
R22435 VGND.n1095 VGND.n1010 3.2005
R22436 VGND.n6252 VGND.n6248 3.2005
R22437 VGND.n2345 VGND.n2344 3.13241
R22438 VGND.n2510 VGND.n2509 3.13241
R22439 VGND.n2307 VGND.n2306 3.13241
R22440 VGND.n5496 VGND.n5495 3.13241
R22441 VGND.n1799 VGND.n1798 3.13241
R22442 VGND.n1737 VGND.n1736 3.13241
R22443 VGND.n7112 VGND.n7111 3.13241
R22444 VGND.n4085 VGND.n4084 3.13241
R22445 VGND.n4866 VGND.n4865 3.13241
R22446 VGND.n1416 VGND.n1415 3.13241
R22447 VGND.n4689 VGND.n4688 3.13241
R22448 VGND.n4668 VGND.n4667 3.13241
R22449 VGND.n4303 VGND.n4302 3.13241
R22450 VGND.n2749 VGND.n2748 3.13241
R22451 VGND.n2834 VGND.n2833 3.13241
R22452 VGND.n2786 VGND.n2785 3.13241
R22453 VGND.n8472 VGND.n8471 3.13241
R22454 VGND.n8488 VGND.n8487 3.13241
R22455 VGND.n8760 VGND.n8759 3.13241
R22456 VGND.n1880 VGND.n1879 3.13241
R22457 VGND.n7946 VGND.n7945 3.13241
R22458 VGND.n8088 VGND.n8087 3.13241
R22459 VGND.n1006 VGND.n1005 3.13241
R22460 VGND.n8702 VGND.n8701 3.10353
R22461 VGND.n3318 VGND.n2648 3.09945
R22462 VGND.n5 VGND.n3 3.06298
R22463 VGND.n1980 VGND.n1979 3.06297
R22464 VGND.n153 VGND.n152 3.06215
R22465 VGND.n1686 VGND.n1670 3.06215
R22466 VGND.n3235 VGND.n3234 3.06214
R22467 VGND.n2659 VGND.n2658 3.06137
R22468 VGND.n9185 VGND.n9184 3.05276
R22469 VGND.n3429 VGND.n3428 3.05276
R22470 VGND.n1293 VGND.n1292 3.05276
R22471 VGND.n6833 VGND.n6829 3.04386
R22472 VGND.n2301 VGND.n2300 3.02516
R22473 VGND.n2724 VGND.n2721 3.02516
R22474 VGND.n4300 VGND.n4299 3.01896
R22475 VGND.n3919 VGND.n3897 3.01896
R22476 VGND.n7341 VGND.n817 3.01896
R22477 VGND.n6277 VGND.n6271 3.01896
R22478 VGND.n2241 VGND.n2240 3.01896
R22479 VGND.n5892 VGND.n5114 3.01896
R22480 VGND.n8890 VGND.n8889 3.01483
R22481 VGND.n1979 VGND.n1978 3.01226
R22482 VGND.n1933 VGND.n1932 3.01226
R22483 VGND.n7319 VGND.n7318 3.01226
R22484 VGND.n4731 VGND.n4730 3.0005
R22485 VGND.n4328 VGND.n4327 3.0005
R22486 VGND.n9078 VGND.n9077 3.0005
R22487 VGND.n8679 VGND.n8678 3.0005
R22488 VGND.n7444 VGND.n7443 3.0005
R22489 VGND.n6175 VGND.n6174 3.0005
R22490 VGND.n1683 VGND.n1682 3.0005
R22491 VGND.n6070 VGND.n6069 3.0005
R22492 VGND.n5629 VGND.n5628 3.0005
R22493 VGND.n5999 VGND.n5998 3.0005
R22494 VGND.n9231 VGND.n9230 3.0005
R22495 VGND.n4510 VGND.n4509 2.99624
R22496 VGND.n8266 VGND.n8264 2.9514
R22497 VGND.n6616 VGND.n1640 2.92166
R22498 VGND.n6670 VGND.n1631 2.92131
R22499 VGND.n84 VGND.n83 2.90959
R22500 VGND.n6852 VGND.n1589 2.90959
R22501 VGND.n6235 VGND.n6234 2.90183
R22502 VGND.n2486 VGND.n2485 2.90012
R22503 VGND.n1515 VGND.n1485 2.86855
R22504 VGND.n4628 VGND.n4627 2.86007
R22505 VGND.n8916 VGND.n81 2.8567
R22506 VGND.n3066 VGND.n3033 2.84782
R22507 VGND.n3631 VGND.n3630 2.83202
R22508 VGND.n7599 VGND.n7598 2.83202
R22509 VGND.n11 VGND.n10 2.79323
R22510 VGND.n2102 VGND.n2101 2.79323
R22511 VGND.n6625 VGND.n6624 2.78311
R22512 VGND.n6690 VGND.n6688 2.77203
R22513 VGND.n8703 VGND.n8699 2.77203
R22514 VGND.n7679 VGND.n7675 2.77203
R22515 VGND.n2809 VGND.n2663 2.76214
R22516 VGND.n2346 VGND.n2345 2.7239
R22517 VGND.n2308 VGND.n2307 2.7239
R22518 VGND.n5497 VGND.n5496 2.7239
R22519 VGND.n1800 VGND.n1799 2.7239
R22520 VGND.n4150 VGND.n4149 2.7239
R22521 VGND.n4667 VGND.n4666 2.7239
R22522 VGND.n1881 VGND.n1880 2.7239
R22523 VGND.n1007 VGND.n1006 2.7239
R22524 VGND.n6225 VGND.n6224 2.7239
R22525 VGND.n6580 VGND.n6579 2.63579
R22526 VGND.n2711 VGND.n2710 2.63579
R22527 VGND.n8944 VGND.n8943 2.63579
R22528 VGND.n8366 VGND.n8365 2.63579
R22529 VGND.n384 VGND.n382 2.63579
R22530 VGND.n8277 VGND.n8276 2.63579
R22531 VGND.n1276 VGND.n1153 2.63579
R22532 VGND.n6906 VGND.n6905 2.63579
R22533 VGND.n9150 VGND.n9149 2.63579
R22534 VGND.n2304 VGND.n2303 2.63064
R22535 VGND.n5560 VGND.n5559 2.63064
R22536 VGND.n4565 VGND.n4564 2.63064
R22537 VGND.n2817 VGND.n2816 2.63064
R22538 VGND.n2719 VGND.n2718 2.63064
R22539 VGND.n254 VGND.n253 2.63064
R22540 VGND.n516 VGND.n515 2.63064
R22541 VGND.n501 VGND.n500 2.63064
R22542 VGND.n8221 VGND.n8220 2.63064
R22543 VGND.n1097 VGND.n1096 2.63064
R22544 VGND.n6251 VGND.n6250 2.63064
R22545 VGND.n8309 VGND.n8308 2.5963
R22546 VGND.n170 VGND.n169 2.58773
R22547 VGND.n341 VGND.n340 2.58773
R22548 VGND.n6917 VGND.n6916 2.58773
R22549 VGND.n3299 VGND.n2649 2.55412
R22550 VGND.n4985 VGND.n4984 2.50485
R22551 VGND.n5092 VGND.n5091 2.47351
R22552 VGND.n4992 VGND.n4991 2.47351
R22553 VGND.n6984 VGND.n6983 2.47351
R22554 VGND.n4341 VGND.n4340 2.47351
R22555 VGND.n2892 VGND.n2891 2.47351
R22556 VGND.n3357 VGND.n3356 2.47351
R22557 VGND.n3140 VGND.n3139 2.47351
R22558 VGND.n8835 VGND.n8834 2.47351
R22559 VGND.n8558 VGND.n8557 2.47351
R22560 VGND.n8802 VGND.n8801 2.47351
R22561 VGND.n8431 VGND.n8430 2.47351
R22562 VGND.n7739 VGND.n7738 2.47351
R22563 VGND.n419 VGND.n418 2.47351
R22564 VGND.n7706 VGND.n7705 2.47351
R22565 VGND.n1171 VGND.n1170 2.47351
R22566 VGND.n880 VGND.n879 2.47351
R22567 VGND.n6946 VGND.n6945 2.47351
R22568 VGND.n6472 VGND.n6471 2.47351
R22569 VGND.n6548 VGND.n6544 2.47351
R22570 VGND.n5316 VGND.n5315 2.47351
R22571 VGND.n5767 VGND.n5766 2.47351
R22572 VGND.n5867 VGND.n5865 2.47351
R22573 VGND.n2277 VGND.n2273 2.47351
R22574 VGND.n2365 VGND.n2364 2.47351
R22575 VGND.n5209 VGND.n5206 2.44756
R22576 VGND.n6379 VGND.n6378 2.40286
R22577 VGND.n6618 VGND.n6617 2.38348
R22578 VGND.n494 VGND.n493 2.36572
R22579 VGND.n2607 VGND.n2606 2.33701
R22580 VGND.n2602 VGND.n2601 2.33701
R22581 VGND.n2219 VGND.n2218 2.33701
R22582 VGND.n2207 VGND.n2206 2.33701
R22583 VGND.n9190 VGND.n9189 2.33701
R22584 VGND.n5270 VGND.n5269 2.33701
R22585 VGND.n5436 VGND.n5435 2.33701
R22586 VGND.n6718 VGND.n6717 2.33701
R22587 VGND.n5365 VGND.n5361 2.33701
R22588 VGND.n6602 VGND.n6601 2.33701
R22589 VGND.n1643 VGND.n1642 2.33701
R22590 VGND.n3434 VGND.n3433 2.33701
R22591 VGND.n3406 VGND.n3405 2.33701
R22592 VGND.n3384 VGND.n3383 2.33701
R22593 VGND.n3308 VGND.n3307 2.33701
R22594 VGND.n3648 VGND.n3647 2.33701
R22595 VGND.n8862 VGND.n8861 2.33701
R22596 VGND.n1509 VGND.n1508 2.33701
R22597 VGND.n1502 VGND.n1501 2.33701
R22598 VGND.n3303 VGND.n3302 2.33067
R22599 VGND.n5390 VGND.n5388 2.32777
R22600 VGND.n7049 VGND.n7048 2.32777
R22601 VGND.n3124 VGND.n3123 2.32777
R22602 VGND.n3099 VGND.n3098 2.32777
R22603 VGND.n7374 VGND.n7373 2.32777
R22604 VGND.n6888 VGND.n6887 2.32777
R22605 VGND.n6840 VGND.n6839 2.32777
R22606 VGND.n6367 VGND.n6366 2.32777
R22607 VGND.n4632 VGND.n4631 2.31539
R22608 VGND.n1400 VGND.n1399 2.31539
R22609 VGND.n3424 VGND.n2110 2.29662
R22610 VGND.n3282 VGND.n3281 2.29662
R22611 VGND.n3664 VGND.n3632 2.29662
R22612 VGND.n8880 VGND.n8879 2.29662
R22613 VGND.n8737 VGND.n180 2.29662
R22614 VGND.n6237 VGND.n6236 2.29662
R22615 VGND.n5374 VGND.n5373 2.29662
R22616 VGND.n6674 VGND.n6673 2.29662
R22617 VGND.n6702 VGND.n6701 2.29662
R22618 VGND.n6704 VGND.n6703 2.29662
R22619 VGND.n9203 VGND.n9 2.29662
R22620 VGND.n2595 VGND.n2594 2.29662
R22621 VGND.n8267 VGND.n445 2.29643
R22622 VGND.n8420 VGND.n8419 2.2824
R22623 VGND.n5336 VGND.n5335 2.2824
R22624 VGND.n9168 VGND.n9167 2.28222
R22625 VGND.n7985 VGND.n7984 2.28171
R22626 VGND.n5454 VGND.n5453 2.28171
R22627 VGND.n3010 VGND.n2879 2.28159
R22628 VGND.n867 VGND.n866 2.28144
R22629 VGND.n1677 VGND.n1672 2.28144
R22630 VGND.n3658 VGND.n3632 2.26126
R22631 VGND.n5035 VGND.n5034 2.25932
R22632 VGND.n5039 VGND.n5038 2.25932
R22633 VGND.n4782 VGND.n4781 2.25932
R22634 VGND.n4382 VGND.n4381 2.25932
R22635 VGND.n4644 VGND.n4643 2.25932
R22636 VGND.n3275 VGND.n3274 2.25932
R22637 VGND.n8948 VGND.n8947 2.25932
R22638 VGND.n8397 VGND.n8396 2.25932
R22639 VGND.n8047 VGND.n491 2.25932
R22640 VGND.n1224 VGND.n1222 2.25932
R22641 VGND.n1233 VGND.n1232 2.25932
R22642 VGND.n1249 VGND.n1246 2.25932
R22643 VGND.n6144 VGND.n6143 2.25932
R22644 VGND.n4592 VGND.n4591 2.23612
R22645 VGND.n4010 VGND.n4009 2.2005
R22646 VGND.n3213 VGND.n3212 2.17922
R22647 VGND.n7893 VGND.n7892 2.17922
R22648 VGND.n6040 VGND.n6039 2.13383
R22649 VGND.n4884 VGND.n4883 2.13383
R22650 VGND.n4461 VGND.n4460 2.13383
R22651 VGND.n2703 VGND.n2702 2.13383
R22652 VGND.n7601 VGND.n7600 2.13383
R22653 VGND.n1620 VGND.n1619 2.11085
R22654 VGND.n9198 VGND.n12 2.09505
R22655 VGND.n3442 VGND.n2103 2.09505
R22656 VGND.n6378 VGND.n6376 2.09362
R22657 VGND.n5361 VGND.n5360 2.08304
R22658 VGND.n526 VGND.n525 2.06919
R22659 VGND.n1644 VGND.n1643 2.03225
R22660 VGND.n4448 VGND.n4447 2.01789
R22661 VGND.n3221 VGND.n3220 2.01694
R22662 VGND.n7900 VGND.n7899 2.01694
R22663 VGND.n1933 VGND.n1930 1.99869
R22664 VGND.n2295 VGND.n2294 1.98299
R22665 VGND.n2178 VGND.n2177 1.98299
R22666 VGND.n5248 VGND.n5247 1.98299
R22667 VGND.n3064 VGND.n3063 1.98299
R22668 VGND.n187 VGND.n186 1.98299
R22669 VGND.n7772 VGND.n7771 1.98299
R22670 VGND.n397 VGND.n396 1.98299
R22671 VGND.n2870 VGND.n2865 1.97497
R22672 VGND.n7617 VGND.n7616 1.97497
R22673 VGND.n3860 VGND.n3859 1.96973
R22674 VGND.n3869 VGND.n3868 1.96973
R22675 VGND.n2695 VGND.n2671 1.93149
R22676 VGND.n8960 VGND.n8958 1.93149
R22677 VGND.n2698 VGND.n2671 1.92649
R22678 VGND.n8958 VGND.n8956 1.92649
R22679 VGND.n3305 VGND.n3304 1.91571
R22680 VGND.n2729 VGND.n2666 1.90688
R22681 VGND.n8586 VGND.n242 1.90688
R22682 VGND.n5241 VGND.n5240 1.8968
R22683 VGND.n527 VGND.n526 1.8968
R22684 VGND.n1904 VGND.n1903 1.89065
R22685 VGND.n179 VGND.n178 1.89043
R22686 VGND.n4874 VGND.n4873 1.88285
R22687 VGND.n4404 VGND.n4403 1.88285
R22688 VGND.n7645 VGND.n7644 1.88285
R22689 VGND.n7687 VGND.n7686 1.88285
R22690 VGND.n2445 VGND.n2444 1.88081
R22691 VGND.n4249 VGND.n4247 1.88081
R22692 VGND.n8983 VGND.n8981 1.88081
R22693 VGND.n6331 VGND.n6329 1.88081
R22694 VGND.n1648 VGND.n1647 1.88022
R22695 VGND.n2659 VGND.n2656 1.87783
R22696 VGND.n6699 VGND.n1623 1.8388
R22697 VGND.n2735 VGND.n2734 1.8388
R22698 VGND.n8591 VGND.n8590 1.8388
R22699 VGND.n711 VGND.n710 1.8388
R22700 VGND.n1484 VGND.n1483 1.80631
R22701 VGND.n1395 VGND.n1394 1.79885
R22702 VGND.n244 VGND.n243 1.79885
R22703 VGND.n1480 VGND.n1479 1.79885
R22704 VGND.n6667 VGND.n6666 1.79699
R22705 VGND.n7025 VGND.n7024 1.79071
R22706 VGND.n4081 VGND.n4080 1.79071
R22707 VGND.n3125 VGND.n3124 1.79071
R22708 VGND.n7660 VGND.n7659 1.79071
R22709 VGND.n8156 VGND.n8155 1.79071
R22710 VGND.n8304 VGND.n8303 1.79071
R22711 VGND.n2566 VGND.n2565 1.77071
R22712 VGND.n4862 VGND.n4861 1.77071
R22713 VGND.n4122 VGND.n4121 1.77071
R22714 VGND.n4605 VGND.n4604 1.77071
R22715 VGND.n2750 VGND.n2749 1.77071
R22716 VGND.n8240 VGND.n8239 1.77071
R22717 VGND.n8598 VGND.n8597 1.75392
R22718 VGND.n5452 VGND.n5451 1.73963
R22719 VGND.n2296 VGND.n2295 1.72441
R22720 VGND.n2179 VGND.n2178 1.72441
R22721 VGND.n3065 VGND.n3064 1.72441
R22722 VGND.n188 VGND.n187 1.72441
R22723 VGND.n7852 VGND.n7851 1.72214
R22724 VGND.n1128 VGND.n1127 1.67669
R22725 VGND.n3072 VGND.n3071 1.61169
R22726 VGND.n6700 VGND.n1621 1.5365
R22727 VGND.n2407 VGND.n2405 1.50935
R22728 VGND.n4770 VGND.n4769 1.50646
R22729 VGND.n4102 VGND.n4101 1.50646
R22730 VGND.n2051 VGND.n2049 1.50646
R22731 VGND.n3673 VGND.n3671 1.50646
R22732 VGND.n3782 VGND.n3781 1.50646
R22733 VGND.n1887 VGND.n1886 1.50646
R22734 VGND.n695 VGND.n694 1.50646
R22735 VGND.n7462 VGND.n7460 1.50646
R22736 VGND.n6120 VGND.n6118 1.50646
R22737 VGND.n1714 VGND.n1712 1.50646
R22738 VGND.n3488 VGND.n3486 1.50646
R22739 VGND.n6588 VGND.n1650 1.50638
R22740 VGND.n5058 VGND.n4037 1.50638
R22741 VGND.n4787 VGND.n4765 1.50638
R22742 VGND.n4792 VGND.n4791 1.50638
R22743 VGND.n4662 VGND.n4167 1.50638
R22744 VGND.n4387 VGND.n4386 1.50638
R22745 VGND.n3269 VGND.n3268 1.50638
R22746 VGND.n8953 VGND.n8952 1.50638
R22747 VGND.n3807 VGND.n3806 1.50638
R22748 VGND.n8392 VGND.n8341 1.50638
R22749 VGND.n1955 VGND.n1920 1.50638
R22750 VGND.n8012 VGND.n8011 1.50638
R22751 VGND.n8041 VGND.n8040 1.50638
R22752 VGND.n7638 VGND.n7605 1.50638
R22753 VGND.n628 VGND.n627 1.50638
R22754 VGND.n1225 VGND.n1158 1.50638
R22755 VGND.n1237 VGND.n1236 1.50638
R22756 VGND.n1269 VGND.n1268 1.50638
R22757 VGND.n1069 VGND.n1012 1.50638
R22758 VGND.n6109 VGND.n6108 1.50638
R22759 VGND.n6450 VGND.n6449 1.50638
R22760 VGND.n4431 VGND.n4430 1.49961
R22761 VGND.n1433 VGND.n1396 1.49961
R22762 VGND.n1432 VGND.n1401 1.49961
R22763 VGND.n8905 VGND.n84 1.49961
R22764 VGND.n2689 VGND.n2674 1.49961
R22765 VGND.n8583 VGND.n245 1.49961
R22766 VGND.n1952 VGND.n1923 1.49961
R22767 VGND.n8379 VGND.n8345 1.49961
R22768 VGND.n1522 VGND.n1481 1.49961
R22769 VGND.n1521 VGND.n1485 1.49961
R22770 VGND.n6855 VGND.n1589 1.49961
R22771 VGND.n6616 VGND.n6615 1.49961
R22772 VGND.n5415 VGND.n5210 1.49961
R22773 VGND.n5149 VGND.n5148 1.49933
R22774 VGND.n7015 VGND.n7013 1.49932
R22775 VGND.n1412 VGND.n1410 1.49932
R22776 VGND.n2911 VGND.n2910 1.49932
R22777 VGND.n8916 VGND.n8914 1.49932
R22778 VGND.n8969 VGND.n8966 1.49932
R22779 VGND.n2684 VGND.n2683 1.49932
R22780 VGND.n8776 VGND.n166 1.49932
R22781 VGND.n8465 VGND.n8463 1.49932
R22782 VGND.n8356 VGND.n8354 1.49932
R22783 VGND.n352 VGND.n351 1.49932
R22784 VGND.n932 VGND.n931 1.49932
R22785 VGND.n1493 VGND.n1491 1.49932
R22786 VGND.n5237 VGND.n5235 1.49932
R22787 VGND.n9122 VGND.n9121 1.49932
R22788 VGND.n690 VGND.n689 1.49837
R22789 VGND.n908 VGND.n907 1.49837
R22790 VGND.n2830 VGND.n2827 1.48166
R22791 VGND.n3401 VGND.n3400 1.46398
R22792 VGND.n913 VGND.n912 1.43682
R22793 VGND.n27 VGND.n26 1.43682
R22794 VGND.n3400 VGND.n3399 1.42915
R22795 VGND.n6668 VGND.n6667 1.42272
R22796 VGND.n6565 VGND.n6564 1.42272
R22797 VGND.n8727 VGND.n8726 1.40924
R22798 VGND.n2923 VGND.n2922 1.3918
R22799 VGND.n5208 VGND.n5207 1.3622
R22800 VGND.n4086 VGND.n4085 1.3622
R22801 VGND.n4087 VGND.n4086 1.3622
R22802 VGND.n8747 VGND.n8746 1.3622
R22803 VGND.n8610 VGND.n8609 1.3622
R22804 VGND.n7947 VGND.n7946 1.3622
R22805 VGND.n7948 VGND.n7947 1.3622
R22806 VGND.n7608 VGND.n7607 1.3622
R22807 VGND.n5969 VGND.n1855 1.35467
R22808 VGND.n4864 VGND.n4090 1.35465
R22809 VGND.n4711 VGND.n4710 1.35465
R22810 VGND.n3579 VGND.n3578 1.35465
R22811 VGND.n3725 VGND.n3724 1.35465
R22812 VGND.n3842 VGND.n3772 1.35465
R22813 VGND.n1969 VGND.n1968 1.35465
R22814 VGND.n7561 VGND.n687 1.35465
R22815 VGND.n9210 VGND.n9209 1.35465
R22816 VGND.n4012 VGND.n4003 1.35464
R22817 VGND.n6728 VGND.n6727 1.35464
R22818 VGND.n5607 VGND.n5606 1.35464
R22819 VGND.n4482 VGND.n4481 1.35464
R22820 VGND.n3244 VGND.n3243 1.35464
R22821 VGND.n9014 VGND.n9013 1.35464
R22822 VGND.n8717 VGND.n8716 1.35464
R22823 VGND.n7914 VGND.n7913 1.35464
R22824 VGND.n8217 VGND.n8216 1.35464
R22825 VGND.n1135 VGND.n1134 1.35464
R22826 VGND.n6793 VGND.n6792 1.35464
R22827 VGND.n2543 VGND.n2542 1.35464
R22828 VGND.n988 VGND.n987 1.35459
R22829 VGND.n5795 VGND.n5794 1.35459
R22830 VGND.n9099 VGND.n9098 1.35459
R22831 VGND.n1461 VGND.n1460 1.35457
R22832 VGND.n2978 VGND.n2977 1.35457
R22833 VGND.n3185 VGND.n3184 1.35457
R22834 VGND.n8416 VGND.n8415 1.35457
R22835 VGND.n6961 VGND.n6960 1.35457
R22836 VGND.n4587 VGND.n4586 1.35455
R22837 VGND.n8313 VGND.n8312 1.35455
R22838 VGND.n1203 VGND.n1202 1.35455
R22839 VGND.n6931 VGND.n6930 1.35455
R22840 VGND.n5752 VGND.n5751 1.35455
R22841 VGND.n2399 VGND.n2398 1.35455
R22842 VGND.n7110 VGND.n1353 1.35455
R22843 VGND.n3013 VGND.n3012 1.35455
R22844 VGND.n3174 VGND.n3173 1.35455
R22845 VGND.n8571 VGND.n256 1.35455
R22846 VGND.n7987 VGND.n7978 1.35455
R22847 VGND.n5457 VGND.n5456 1.35455
R22848 VGND.n3639 VGND.n3638 1.3469
R22849 VGND.n6617 VGND.n1639 1.3283
R22850 VGND.n4435 VGND.n4433 1.32281
R22851 VGND.n1927 VGND.n1925 1.32281
R22852 VGND.n1922 VGND.n1921 1.32281
R22853 VGND.n9166 VGND.n9165 1.32281
R22854 VGND.n228 VGND.n227 1.30065
R22855 VGND.n1091 VGND.n1086 1.30065
R22856 VGND.n3662 VGND.n3658 1.29559
R22857 VGND.n3880 VGND.n3879 1.29412
R22858 VGND.n7800 VGND.n7799 1.29412
R22859 VGND.n8596 VGND.n237 1.27173
R22860 VGND.n7789 VGND.n7788 1.27173
R22861 VGND.n8728 VGND.n8727 1.26145
R22862 VGND.n2351 VGND.n2350 1.25365
R22863 VGND.n4236 VGND.n4235 1.25365
R22864 VGND.n9016 VGND.n9015 1.25365
R22865 VGND.n6301 VGND.n6300 1.25365
R22866 VGND.n3323 VGND.n2647 1.25033
R22867 VGND.n8532 VGND.n8531 1.22603
R22868 VGND.n8581 VGND.n8580 1.22603
R22869 VGND.n2646 VGND.n2125 1.1942
R22870 VGND.n101 VGND.n100 1.1942
R22871 VGND.n2475 VGND.n2474 1.18311
R22872 VGND.n5136 VGND.n5135 1.18311
R22873 VGND.n1857 VGND.n1856 1.18311
R22874 VGND.n1804 VGND.n1803 1.18311
R22875 VGND.n1710 VGND.n1709 1.18311
R22876 VGND.n1346 VGND.n1345 1.18311
R22877 VGND.n4036 VGND.n4035 1.18311
R22878 VGND.n5048 VGND.n5047 1.18311
R22879 VGND.n4239 VGND.n4238 1.18311
R22880 VGND.n4452 VGND.n4451 1.18311
R22881 VGND.n4653 VGND.n4652 1.18311
R22882 VGND.n2904 VGND.n2903 1.18311
R22883 VGND.n2047 VGND.n2046 1.18311
R22884 VGND.n3669 VGND.n3668 1.18311
R22885 VGND.n3796 VGND.n3773 1.18311
R22886 VGND.n225 VGND.n224 1.18311
R22887 VGND.n1901 VGND.n1900 1.18311
R22888 VGND.n496 VGND.n495 1.18311
R22889 VGND.n7842 VGND.n503 1.18311
R22890 VGND.n904 VGND.n903 1.18311
R22891 VGND.n7458 VGND.n7457 1.18311
R22892 VGND.n6261 VGND.n6260 1.18311
R22893 VGND.n6353 VGND.n6352 1.18311
R22894 VGND.n6359 VGND.n6358 1.18311
R22895 VGND.n7223 VGND.n7222 1.17646
R22896 VGND.n2776 VGND.n2764 1.17646
R22897 VGND.n9046 VGND.n9045 1.17646
R22898 VGND.n8707 VGND.n8706 1.17646
R22899 VGND.n8092 VGND.n8091 1.17646
R22900 VGND.n6819 VGND.n1592 1.17646
R22901 VGND.n5368 VGND.n5346 1.17646
R22902 VGND.n5639 VGND.n5471 1.17646
R22903 VGND.n4514 VGND.n4494 1.17642
R22904 VGND.n8193 VGND.n8153 1.17642
R22905 VGND.n1318 VGND.n1317 1.17642
R22906 VGND.n2514 VGND.n2513 1.17642
R22907 VGND.n4303 VGND.n4301 1.15795
R22908 VGND.n2303 VGND.n2302 1.14023
R22909 VGND.n5696 VGND.n5695 1.14023
R22910 VGND.n5659 VGND.n5658 1.14023
R22911 VGND.n5559 VGND.n5558 1.14023
R22912 VGND.n4593 VGND.n4592 1.14023
R22913 VGND.n2948 VGND.n2946 1.14023
R22914 VGND.n2948 VGND.n2947 1.14023
R22915 VGND.n2816 VGND.n2815 1.14023
R22916 VGND.n3220 VGND.n3219 1.14023
R22917 VGND.n2720 VGND.n2719 1.14023
R22918 VGND.n8927 VGND.n8926 1.14023
R22919 VGND.n8508 VGND.n8506 1.14023
R22920 VGND.n8508 VGND.n8507 1.14023
R22921 VGND.n253 VGND.n252 1.14023
R22922 VGND.n3961 VGND.n3960 1.14023
R22923 VGND.n8600 VGND.n8599 1.14023
R22924 VGND.n208 VGND.n207 1.14023
R22925 VGND.n515 VGND.n514 1.14023
R22926 VGND.n500 VGND.n499 1.14023
R22927 VGND.n7899 VGND.n7898 1.14023
R22928 VGND.n361 VGND.n360 1.14023
R22929 VGND.n8222 VGND.n8221 1.14023
R22930 VGND.n961 VGND.n960 1.14023
R22931 VGND.n1096 VGND.n1095 1.14023
R22932 VGND.n7416 VGND.n7415 1.14023
R22933 VGND.n6252 VGND.n6251 1.14023
R22934 VGND.n9154 VGND.n9153 1.14023
R22935 VGND.n6736 VGND.n1613 1.13896
R22936 VGND.n5003 VGND.n5002 1.13896
R22937 VGND.n1457 VGND.n1378 1.13896
R22938 VGND.n2761 VGND.n47 1.13896
R22939 VGND.n3345 VGND.n3334 1.13896
R22940 VGND.n9050 VGND.n9049 1.13896
R22941 VGND.n8823 VGND.n134 1.13896
R22942 VGND.n8711 VGND.n8710 1.13896
R22943 VGND.n8793 VGND.n135 1.13896
R22944 VGND.n8096 VGND.n8095 1.13896
R22945 VGND.n7727 VGND.n571 1.13896
R22946 VGND.n8320 VGND.n412 1.13896
R22947 VGND.n7697 VGND.n582 1.13896
R22948 VGND.n4363 VGND.n4362 1.13896
R22949 VGND.n8320 VGND.n8319 1.13896
R22950 VGND.n4582 VGND.n1378 1.13896
R22951 VGND.n8096 VGND.n461 1.13896
R22952 VGND.n8712 VGND.n8711 1.13896
R22953 VGND.n9050 VGND.n57 1.13896
R22954 VGND.n3239 VGND.n47 1.13896
R22955 VGND.n8212 VGND.n8211 1.13896
R22956 VGND.n4489 VGND.n4488 1.13896
R22957 VGND.n2003 VGND.n2002 1.13896
R22958 VGND.n3767 VGND.n3766 1.13896
R22959 VGND.n3621 VGND.n3620 1.13896
R22960 VGND.n2092 VGND.n2091 1.13896
R22961 VGND.n7520 VGND.n7519 1.13896
R22962 VGND.n4823 VGND.n4822 1.13896
R22963 VGND.n1750 VGND.n1697 1.13896
R22964 VGND.n4143 VGND.n4142 1.13896
R22965 VGND.n6999 VGND.n6998 1.13885
R22966 VGND.n7227 VGND.n7226 1.13885
R22967 VGND.n2974 VGND.n2744 1.13885
R22968 VGND.n3181 VGND.n3180 1.13885
R22969 VGND.n8447 VGND.n8446 1.13885
R22970 VGND.n8412 VGND.n279 1.13885
R22971 VGND.n2235 VGND.n2163 1.13885
R22972 VGND.n6523 VGND.n6522 1.13885
R22973 VGND.n5219 VGND.n5192 1.13885
R22974 VGND.n5791 VGND.n5790 1.13885
R22975 VGND.n2394 VGND.n43 1.13885
R22976 VGND.n5619 VGND.n5618 1.13885
R22977 VGND.n2538 VGND.n2537 1.13885
R22978 VGND.n6007 VGND.n1789 1.13885
R22979 VGND.n5854 VGND.n5853 1.13885
R22980 VGND.n6734 VGND.n6733 1.13717
R22981 VGND.n6014 VGND.n6013 1.13717
R22982 VGND.n6996 VGND.n6995 1.13717
R22983 VGND.n4002 VGND.n4001 1.13717
R22984 VGND.n4762 VGND.n4761 1.13717
R22985 VGND.n4054 VGND.n4053 1.13717
R22986 VGND.n4709 VGND.n4708 1.13717
R22987 VGND.n4493 VGND.n4492 1.13717
R22988 VGND.n4370 VGND.n4369 1.13717
R22989 VGND.n3017 VGND.n3016 1.13717
R22990 VGND.n3581 VGND.n3580 1.13717
R22991 VGND.n3333 VGND.n3332 1.13717
R22992 VGND.n3343 VGND.n3342 1.13717
R22993 VGND.n3178 VGND.n3177 1.13717
R22994 VGND.n3727 VGND.n3726 1.13717
R22995 VGND.n133 VGND.n132 1.13717
R22996 VGND.n8821 VGND.n8820 1.13717
R22997 VGND.n8444 VGND.n8443 1.13717
R22998 VGND.n3771 VGND.n3770 1.13717
R22999 VGND.n8795 VGND.n8794 1.13717
R23000 VGND.n3895 VGND.n3894 1.13717
R23001 VGND.n7977 VGND.n7976 1.13717
R23002 VGND.n1967 VGND.n1966 1.13717
R23003 VGND.n570 VGND.n569 1.13717
R23004 VGND.n7725 VGND.n7724 1.13717
R23005 VGND.n7517 VGND.n7516 1.13717
R23006 VGND.n8152 VGND.n8151 1.13717
R23007 VGND.n7699 VGND.n7698 1.13717
R23008 VGND.n580 VGND.n579 1.13717
R23009 VGND.n1320 VGND.n1319 1.13717
R23010 VGND.n800 VGND.n799 1.13717
R23011 VGND.n6929 VGND.n6928 1.13717
R23012 VGND.n6211 VGND.n6210 1.13717
R23013 VGND.n6463 VGND.n6462 1.13717
R23014 VGND.n2629 VGND.n2628 1.13717
R23015 VGND.n2272 VGND.n2271 1.13717
R23016 VGND.n2161 VGND.n2160 1.13717
R23017 VGND.n6475 VGND.n6473 1.13717
R23018 VGND.n6491 VGND.n6490 1.13717
R23019 VGND.n7330 VGND.n7329 1.13717
R23020 VGND.n7736 VGND.n7735 1.13717
R23021 VGND.n7729 VGND.n555 1.13717
R23022 VGND.n8804 VGND.n8803 1.13717
R23023 VGND.n8810 VGND.n148 1.13717
R23024 VGND.n8832 VGND.n8831 1.13717
R23025 VGND.n8825 VGND.n117 1.13717
R23026 VGND.n3354 VGND.n3353 1.13717
R23027 VGND.n3347 VGND.n2141 1.13717
R23028 VGND.n7708 VGND.n7707 1.13717
R23029 VGND.n7714 VGND.n595 1.13717
R23030 VGND.n5005 VGND.n5004 1.13717
R23031 VGND.n4994 VGND.n4993 1.13717
R23032 VGND.n5000 VGND.n4071 1.13717
R23033 VGND.n4343 VGND.n4342 1.13717
R23034 VGND.n4350 VGND.n4349 1.13717
R23035 VGND.n4361 VGND.n4359 1.13717
R23036 VGND.n7325 VGND.n7324 1.13717
R23037 VGND.n860 VGND.n859 1.13717
R23038 VGND.n841 VGND.n840 1.13717
R23039 VGND.n6269 VGND.n6268 1.13717
R23040 VGND.n2238 VGND.n2237 1.13717
R23041 VGND.n6504 VGND.n6501 1.13717
R23042 VGND.n6521 VGND.n6520 1.13717
R23043 VGND.n6543 VGND.n6542 1.13717
R23044 VGND.n6536 VGND.n6535 1.13717
R23045 VGND.n5461 VGND.n5460 1.13717
R23046 VGND.n5750 VGND.n5749 1.13717
R23047 VGND.n9097 VGND.n9096 1.13717
R23048 VGND.n39 VGND.n38 1.13717
R23049 VGND.n2377 VGND.n2376 1.13717
R23050 VGND.n6953 VGND.n6948 1.13717
R23051 VGND.n1553 VGND.n1551 1.13717
R23052 VGND.n6959 VGND.n6958 1.13717
R23053 VGND.n8318 VGND.n8316 1.13717
R23054 VGND.n8434 VGND.n8433 1.13717
R23055 VGND.n289 VGND.n288 1.13717
R23056 VGND.n8414 VGND.n8413 1.13717
R23057 VGND.n8553 VGND.n8552 1.13717
R23058 VGND.n8546 VGND.n8545 1.13717
R23059 VGND.n8449 VGND.n8448 1.13717
R23060 VGND.n3158 VGND.n3157 1.13717
R23061 VGND.n3151 VGND.n3150 1.13717
R23062 VGND.n3183 VGND.n3182 1.13717
R23063 VGND.n3003 VGND.n3002 1.13717
R23064 VGND.n2996 VGND.n2995 1.13717
R23065 VGND.n2976 VGND.n2975 1.13717
R23066 VGND.n8325 VGND.n8324 1.13717
R23067 VGND.n411 VGND.n410 1.13717
R23068 VGND.n427 VGND.n426 1.13717
R23069 VGND.n990 VGND.n989 1.13717
R23070 VGND.n7301 VGND.n7300 1.13717
R23071 VGND.n1181 VGND.n1180 1.13717
R23072 VGND.n1201 VGND.n1200 1.13717
R23073 VGND.n4585 VGND.n4584 1.13717
R23074 VGND.n7094 VGND.n7093 1.13717
R23075 VGND.n7087 VGND.n7086 1.13717
R23076 VGND.n7001 VGND.n7000 1.13717
R23077 VGND.n5319 VGND.n5318 1.13717
R23078 VGND.n5326 VGND.n5325 1.13717
R23079 VGND.n5221 VGND.n5220 1.13717
R23080 VGND.n1459 VGND.n1458 1.13717
R23081 VGND.n1567 VGND.n1566 1.13717
R23082 VGND.n6987 VGND.n6986 1.13717
R23083 VGND.n5793 VGND.n5792 1.13717
R23084 VGND.n5788 VGND.n5785 1.13717
R23085 VGND.n5770 VGND.n5769 1.13717
R23086 VGND.n2397 VGND.n2396 1.13717
R23087 VGND.n5612 VGND.n5611 1.13717
R23088 VGND.n2516 VGND.n2515 1.13717
R23089 VGND.n2326 VGND.n2325 1.13717
R23090 VGND.n2535 VGND.n2534 1.13717
R23091 VGND.n5617 VGND.n5616 1.13717
R23092 VGND.n5624 VGND.n5623 1.13717
R23093 VGND.n6791 VGND.n6790 1.13717
R23094 VGND.n7290 VGND.n7288 1.13717
R23095 VGND.n8094 VGND.n8093 1.13717
R23096 VGND.n8110 VGND.n8107 1.13717
R23097 VGND.n475 VGND.n471 1.13717
R23098 VGND.n7912 VGND.n7911 1.13717
R23099 VGND.n8709 VGND.n8708 1.13717
R23100 VGND.n8692 VGND.n8691 1.13717
R23101 VGND.n8674 VGND.n8673 1.13717
R23102 VGND.n8715 VGND.n8714 1.13717
R23103 VGND.n9048 VGND.n9047 1.13717
R23104 VGND.n71 VGND.n68 1.13717
R23105 VGND.n9064 VGND.n9060 1.13717
R23106 VGND.n9012 VGND.n9011 1.13717
R23107 VGND.n2763 VGND.n2762 1.13717
R23108 VGND.n9072 VGND.n9071 1.13717
R23109 VGND.n9086 VGND.n9082 1.13717
R23110 VGND.n3242 VGND.n3241 1.13717
R23111 VGND.n8122 VGND.n8121 1.13717
R23112 VGND.n8209 VGND.n8208 1.13717
R23113 VGND.n8215 VGND.n8214 1.13717
R23114 VGND.n1139 VGND.n1138 1.13717
R23115 VGND.n7271 VGND.n7270 1.13717
R23116 VGND.n4202 VGND.n4201 1.13717
R23117 VGND.n4208 VGND.n4195 1.13717
R23118 VGND.n7251 VGND.n7250 1.13717
R23119 VGND.n7236 VGND.n7235 1.13717
R23120 VGND.n7225 VGND.n7224 1.13717
R23121 VGND.n6741 VGND.n6740 1.13717
R23122 VGND.n6760 VGND.n6757 1.13717
R23123 VGND.n5345 VGND.n5344 1.13717
R23124 VGND.n4487 VGND.n4485 1.13717
R23125 VGND.n6784 VGND.n6783 1.13717
R23126 VGND.n6779 VGND.n6778 1.13717
R23127 VGND.n1611 VGND.n1610 1.13717
R23128 VGND.n5483 VGND.n5482 1.13717
R23129 VGND.n2541 VGND.n2540 1.13717
R23130 VGND.n6194 VGND.n6191 1.13717
R23131 VGND.n6167 VGND.n6166 1.13717
R23132 VGND.n764 VGND.n762 1.13717
R23133 VGND.n7449 VGND.n7448 1.13717
R23134 VGND.n2023 VGND.n2022 1.13717
R23135 VGND.n2029 VGND.n2015 1.13717
R23136 VGND.n2001 VGND.n1999 1.13717
R23137 VGND.n3750 VGND.n3749 1.13717
R23138 VGND.n3756 VGND.n3742 1.13717
R23139 VGND.n3765 VGND.n3763 1.13717
R23140 VGND.n3604 VGND.n3603 1.13717
R23141 VGND.n3610 VGND.n3596 1.13717
R23142 VGND.n3619 VGND.n3617 1.13717
R23143 VGND.n3548 VGND.n3547 1.13717
R23144 VGND.n3555 VGND.n3554 1.13717
R23145 VGND.n2090 VGND.n2088 1.13717
R23146 VGND.n741 VGND.n740 1.13717
R23147 VGND.n747 VGND.n733 1.13717
R23148 VGND.n7523 VGND.n7522 1.13717
R23149 VGND.n4832 VGND.n4831 1.13717
R23150 VGND.n4839 VGND.n4838 1.13717
R23151 VGND.n4821 VGND.n4819 1.13717
R23152 VGND.n6082 VGND.n6081 1.13717
R23153 VGND.n6088 VGND.n6074 1.13717
R23154 VGND.n1753 VGND.n1752 1.13717
R23155 VGND.n4743 VGND.n4742 1.13717
R23156 VGND.n4749 VGND.n4735 1.13717
R23157 VGND.n4141 VGND.n4139 1.13717
R23158 VGND.n7498 VGND.n7497 1.13717
R23159 VGND.n6159 VGND.n6158 1.13717
R23160 VGND.n9226 VGND.n9225 1.13717
R23161 VGND.n3533 VGND.n3532 1.13717
R23162 VGND.n1788 VGND.n1785 1.13717
R23163 VGND.n1854 VGND.n1853 1.13717
R23164 VGND.n5984 VGND.n5983 1.13717
R23165 VGND.n6004 VGND.n6003 1.13717
R23166 VGND.n5833 VGND.n5829 1.13717
R23167 VGND.n5851 VGND.n5121 1.13717
R23168 VGND.n5856 VGND.n5855 1.13717
R23169 VGND.n5843 VGND.n5842 1.13717
R23170 VGND.n5852 VGND.n5851 1.1368
R23171 VGND.n7729 VGND.n7728 1.1368
R23172 VGND.n8811 VGND.n8810 1.1368
R23173 VGND.n8825 VGND.n8824 1.1368
R23174 VGND.n3347 VGND.n3346 1.1368
R23175 VGND.n7715 VGND.n7714 1.1368
R23176 VGND.n5001 VGND.n5000 1.1368
R23177 VGND.n4349 VGND.n4231 1.1368
R23178 VGND.n2162 VGND.n2161 1.1368
R23179 VGND.n5789 VGND.n5788 1.1368
R23180 VGND.n2376 VGND.n2370 1.1368
R23181 VGND.n5623 VGND.n5620 1.1368
R23182 VGND.n476 VGND.n475 1.1368
R23183 VGND.n8673 VGND.n203 1.1368
R23184 VGND.n9065 VGND.n9064 1.1368
R23185 VGND.n9087 VGND.n9086 1.1368
R23186 VGND.n8210 VGND.n8209 1.1368
R23187 VGND.n4209 VGND.n4208 1.1368
R23188 VGND.n2536 VGND.n2535 1.1368
R23189 VGND.n2030 VGND.n2029 1.1368
R23190 VGND.n3757 VGND.n3756 1.1368
R23191 VGND.n3611 VGND.n3610 1.1368
R23192 VGND.n3554 VGND.n3540 1.1368
R23193 VGND.n748 VGND.n747 1.1368
R23194 VGND.n4838 VGND.n4824 1.1368
R23195 VGND.n6089 VGND.n6088 1.1368
R23196 VGND.n4750 VGND.n4749 1.1368
R23197 VGND.n3534 VGND.n3533 1.1368
R23198 VGND.n7726 VGND.n7725 1.13669
R23199 VGND.n3894 VGND.n3892 1.13669
R23200 VGND.n8822 VGND.n8821 1.13669
R23201 VGND.n3344 VGND.n3343 1.13669
R23202 VGND.n581 VGND.n580 1.13669
R23203 VGND.n4055 VGND.n4054 1.13669
R23204 VGND.n4369 VGND.n4367 1.13669
R23205 VGND.n5834 VGND.n5833 1.13669
R23206 VGND.n2630 VGND.n2629 1.13669
R23207 VGND.n6505 VGND.n6504 1.13669
R23208 VGND.n6536 VGND.n6524 1.13669
R23209 VGND.n7976 VGND.n7974 1.13669
R23210 VGND.n8435 VGND.n8434 1.13669
R23211 VGND.n8445 VGND.n8444 1.13669
R23212 VGND.n8552 VGND.n265 1.13669
R23213 VGND.n3179 VGND.n3178 1.13669
R23214 VGND.n3157 VGND.n3021 1.13669
R23215 VGND.n3018 VGND.n3017 1.13669
R23216 VGND.n3002 VGND.n2887 1.13669
R23217 VGND.n8324 VGND.n8321 1.13669
R23218 VGND.n426 VGND.n318 1.13669
R23219 VGND.n6997 VGND.n6996 1.13669
R23220 VGND.n7093 VGND.n1364 1.13669
R23221 VGND.n5462 VGND.n5461 1.13669
R23222 VGND.n5319 VGND.n5299 1.13669
R23223 VGND.n1568 VGND.n1567 1.13669
R23224 VGND.n6988 VGND.n6987 1.13669
R23225 VGND.n5749 VGND.n5191 1.13669
R23226 VGND.n9096 VGND.n9094 1.13669
R23227 VGND.n8111 VGND.n8110 1.13669
R23228 VGND.n8691 VGND.n200 1.13669
R23229 VGND.n72 VGND.n71 1.13669
R23230 VGND.n9071 VGND.n9068 1.13669
R23231 VGND.n8151 VGND.n460 1.13669
R23232 VGND.n4492 VGND.n4490 1.13669
R23233 VGND.n4001 VGND.n1322 1.13669
R23234 VGND.n7252 VGND.n7251 1.13669
R23235 VGND.n6761 VGND.n6760 1.13669
R23236 VGND.n6735 VGND.n6734 1.13669
R23237 VGND.n5613 VGND.n5612 1.13669
R23238 VGND.n2517 VGND.n2516 1.13669
R23239 VGND.n1966 VGND.n1875 1.13669
R23240 VGND.n3770 VGND.n3768 1.13669
R23241 VGND.n3728 VGND.n3727 1.13669
R23242 VGND.n3582 VGND.n3581 1.13669
R23243 VGND.n7518 VGND.n7517 1.13669
R23244 VGND.n4763 VGND.n4762 1.13669
R23245 VGND.n6013 VGND.n6011 1.13669
R23246 VGND.n4708 VGND.n4706 1.13669
R23247 VGND.n6008 VGND.n1788 1.13669
R23248 VGND.n6006 VGND.n6004 1.13669
R23249 VGND.n956 VGND.n916 1.12991
R23250 VGND.n1029 VGND.n1016 1.12991
R23251 VGND.n983 VGND.n982 1.11354
R23252 VGND.n3446 VGND.n2103 1.09272
R23253 VGND.n7669 VGND.n7600 1.09272
R23254 VGND.n8264 VGND.n8263 1.09272
R23255 VGND.n9202 VGND.n12 1.09272
R23256 VGND.n4951 VGND.n4949 1.08588
R23257 VGND.n4958 VGND.n4957 1.08588
R23258 VGND.n2802 VGND.n2798 1.08588
R23259 VGND.n329 VGND.n328 1.07463
R23260 VGND.n1107 VGND.n1106 1.02178
R23261 VGND.n2810 VGND.n2809 1.00931
R23262 VGND.n2577 VGND.n2576 1.00568
R23263 VGND.n5800 VGND.n5797 0.985115
R23264 VGND.n329 VGND.n327 0.985115
R23265 VGND.n3798 VGND.n3797 0.974413
R23266 VGND.n6389 VGND.n6388 0.974413
R23267 VGND.n4986 VGND.n4985 0.973599
R23268 VGND.n2751 VGND.n2750 0.953691
R23269 VGND.n8088 VGND.n8086 0.953691
R23270 VGND.n670 VGND.n669 0.953691
R23271 VGND.n5147 VGND.n5146 0.952566
R23272 VGND.n4219 VGND.n4218 0.952566
R23273 VGND.n1400 VGND.n1398 0.952566
R23274 VGND.n2878 VGND.n2877 0.952566
R23275 VGND.n2673 VGND.n2672 0.952566
R23276 VGND.n8968 VGND.n8967 0.952566
R23277 VGND.n164 VGND.n163 0.952566
R23278 VGND.n8384 VGND.n8383 0.952566
R23279 VGND.n7570 VGND.n7569 0.944279
R23280 VGND.n1445 VGND.n1444 0.931411
R23281 VGND.n1534 VGND.n1533 0.931411
R23282 VGND.n8345 VGND.n8344 0.899674
R23283 VGND.n4172 VGND.n4171 0.895605
R23284 VGND.n8172 VGND.n8171 0.895605
R23285 VGND.n6881 VGND.n6880 0.895605
R23286 VGND.n6846 VGND.n6845 0.895605
R23287 VGND.n12 VGND.n11 0.892621
R23288 VGND.n2103 VGND.n2102 0.892621
R23289 VGND.n8599 VGND.n8598 0.877212
R23290 VGND.n7806 VGND.n7805 0.860318
R23291 VGND.n3632 VGND.n3631 0.853833
R23292 VGND.n7600 VGND.n7599 0.853833
R23293 VGND.n984 VGND.n983 0.835283
R23294 VGND.n2574 VGND.n2300 0.833377
R23295 VGND.n5693 VGND.n5692 0.833377
R23296 VGND.n5656 VGND.n5655 0.833377
R23297 VGND.n5557 VGND.n5554 0.833377
R23298 VGND.n4561 VGND.n4558 0.833377
R23299 VGND.n4598 VGND.n4597 0.833377
R23300 VGND.n2953 VGND.n2952 0.833377
R23301 VGND.n2755 VGND.n2663 0.833377
R23302 VGND.n3218 VGND.n3215 0.833377
R23303 VGND.n2725 VGND.n2724 0.833377
R23304 VGND.n8931 VGND.n8930 0.833377
R23305 VGND.n8513 VGND.n8512 0.833377
R23306 VGND.n251 VGND.n248 0.833377
R23307 VGND.n3966 VGND.n3965 0.833377
R23308 VGND.n8604 VGND.n8603 0.833377
R23309 VGND.n212 VGND.n211 0.833377
R23310 VGND.n513 VGND.n510 0.833377
R23311 VGND.n7864 VGND.n7863 0.833377
R23312 VGND.n7897 VGND.n7894 0.833377
R23313 VGND.n366 VGND.n365 0.833377
R23314 VGND.n8229 VGND.n8228 0.833377
R23315 VGND.n8228 VGND.n8225 0.833377
R23316 VGND.n966 VGND.n965 0.833377
R23317 VGND.n1087 VGND.n1010 0.833377
R23318 VGND.n7421 VGND.n7420 0.833377
R23319 VGND.n6248 VGND.n6245 0.833377
R23320 VGND.n9159 VGND.n9158 0.833377
R23321 VGND.n3304 VGND.n3303 0.830425
R23322 VGND.n7078 VGND.n7077 0.817521
R23323 VGND.n1075 VGND.n1074 0.817521
R23324 VGND.n3318 VGND.n3317 0.798505
R23325 VGND.n5595 VGND.n5593 0.765717
R23326 VGND.n984 VGND.n981 0.765717
R23327 VGND.n7338 VGND.n7337 0.765717
R23328 VGND.n2467 VGND.n2466 0.753441
R23329 VGND.n2553 VGND.n2552 0.753441
R23330 VGND.n6054 VGND.n1770 0.753441
R23331 VGND.n7118 VGND.n1351 0.753441
R23332 VGND.n7128 VGND.n7127 0.753441
R23333 VGND.n7163 VGND.n7162 0.753441
R23334 VGND.n7181 VGND.n7180 0.753441
R23335 VGND.n7173 VGND.n7172 0.753441
R23336 VGND.n7219 VGND.n7218 0.753441
R23337 VGND.n4015 VGND.n4014 0.753441
R23338 VGND.n4026 VGND.n4025 0.753441
R23339 VGND.n5054 VGND.n5053 0.753441
R23340 VGND.n4899 VGND.n4898 0.753441
R23341 VGND.n4677 VGND.n4676 0.753441
R23342 VGND.n4281 VGND.n4278 0.753441
R23343 VGND.n4281 VGND.n4280 0.753441
R23344 VGND.n4394 VGND.n4393 0.753441
R23345 VGND.n4476 VGND.n4215 0.753441
R23346 VGND.n4638 VGND.n4637 0.753441
R23347 VGND.n9042 VGND.n9039 0.753441
R23348 VGND.n9042 VGND.n9041 0.753441
R23349 VGND.n3807 VGND.n3805 0.753441
R23350 VGND.n3932 VGND.n3931 0.753441
R23351 VGND.n8358 VGND.n8357 0.753441
R23352 VGND.n1913 VGND.n1912 0.753441
R23353 VGND.n8005 VGND.n8004 0.753441
R23354 VGND.n8025 VGND.n7951 0.753441
R23355 VGND.n1947 VGND.n1946 0.753441
R23356 VGND.n7876 VGND.n7875 0.753441
R23357 VGND.n7885 VGND.n7884 0.753441
R23358 VGND.n7905 VGND.n7904 0.753441
R23359 VGND.n658 VGND.n657 0.753441
R23360 VGND.n1249 VGND.n1248 0.753441
R23361 VGND.n1254 VGND.n1253 0.753441
R23362 VGND.n6298 VGND.n6295 0.753441
R23363 VGND.n6298 VGND.n6297 0.753441
R23364 VGND.n6401 VGND.n6400 0.753441
R23365 VGND.n7078 VGND.n7076 0.749436
R23366 VGND.n3190 VGND.n3187 0.749436
R23367 VGND.n1208 VGND.n1207 0.749436
R23368 VGND.n8889 VGND.n8888 0.743162
R23369 VGND.n6821 VGND.n6820 0.716584
R23370 VGND.n6046 VGND.n6045 0.711611
R23371 VGND.n1653 VGND.n1652 0.711611
R23372 VGND.n4880 VGND.n4879 0.711611
R23373 VGND.n4465 VGND.n4464 0.711611
R23374 VGND.n2707 VGND.n2706 0.711611
R23375 VGND.n1313 VGND.n1312 0.711611
R23376 VGND.n4564 VGND.n4563 0.70187
R23377 VGND.n5061 VGND.n5060 0.696152
R23378 VGND.n236 VGND.n234 0.696152
R23379 VGND.n1937 VGND.n1936 0.689731
R23380 VGND.n4651 VGND.n4553 0.629895
R23381 VGND.n2591 VGND.n2292 0.627073
R23382 VGND.n2228 VGND.n2227 0.627073
R23383 VGND.n7546 VGND.n7545 0.627073
R23384 VGND.n4621 VGND.n4620 0.614199
R23385 VGND.n3222 VGND.n3221 0.614199
R23386 VGND.n7901 VGND.n7900 0.614199
R23387 VGND.n8534 VGND.n8532 0.613266
R23388 VGND.n3302 VGND.n3299 0.606984
R23389 VGND.n8701 VGND.n8700 0.603867
R23390 VGND.n2038 VGND.n2037 0.546928
R23391 VGND.n3538 VGND.n45 0.546928
R23392 VGND.n2497 VGND.n2496 0.545181
R23393 VGND.n2336 VGND.n2335 0.545181
R23394 VGND.n4516 VGND.n4515 0.545181
R23395 VGND.n8069 VGND.n8068 0.545181
R23396 VGND.n2444 VGND.n2348 0.537563
R23397 VGND.n2419 VGND.n2351 0.537563
R23398 VGND.n2619 VGND.n2618 0.537563
R23399 VGND.n2275 VGND.n2274 0.537563
R23400 VGND.n2190 VGND.n2180 0.537563
R23401 VGND.n2189 VGND.n2184 0.537563
R23402 VGND.n5800 VGND.n5799 0.537563
R23403 VGND.n5799 VGND.n5798 0.537563
R23404 VGND.n5163 VGND.n5127 0.537563
R23405 VGND.n5702 VGND.n5701 0.537563
R23406 VGND.n5725 VGND.n5469 0.537563
R23407 VGND.n5505 VGND.n5504 0.537563
R23408 VGND.n5528 VGND.n5498 0.537563
R23409 VGND.n5927 VGND.n5926 0.537563
R23410 VGND.n5904 VGND.n5111 0.537563
R23411 VGND.n5964 VGND.n1859 0.537563
R23412 VGND.n5941 VGND.n1860 0.537563
R23413 VGND.n5399 VGND.n5398 0.537563
R23414 VGND.n6592 VGND.n1648 0.537563
R23415 VGND.n7042 VGND.n7010 0.537563
R23416 VGND.n7016 VGND.n7011 0.537563
R23417 VGND.n7043 VGND.n7006 0.537563
R23418 VGND.n4920 VGND.n4919 0.537563
R23419 VGND.n4945 VGND.n4082 0.537563
R23420 VGND.n4249 VGND.n4248 0.537563
R23421 VGND.n4274 VGND.n4236 0.537563
R23422 VGND.n4522 VGND.n4173 0.537563
R23423 VGND.n4528 VGND.n4527 0.537563
R23424 VGND.n4548 VGND.n4547 0.537563
R23425 VGND.n2061 VGND.n2060 0.537563
R23426 VGND.n3105 VGND.n3104 0.537563
R23427 VGND.n3078 VGND.n3077 0.537563
R23428 VGND.n3103 VGND.n3027 0.537563
R23429 VGND.n3076 VGND.n3031 0.537563
R23430 VGND.n3050 VGND.n3049 0.537563
R23431 VGND.n8983 VGND.n8982 0.537563
R23432 VGND.n3849 VGND.n3848 0.537563
R23433 VGND.n1864 VGND.n1863 0.537563
R23434 VGND.n7787 VGND.n519 0.537563
R23435 VGND.n7766 VGND.n529 0.537563
R23436 VGND.n7830 VGND.n505 0.537563
R23437 VGND.n385 VGND.n336 0.537563
R23438 VGND.n7583 VGND.n686 0.537563
R23439 VGND.n7587 VGND.n7586 0.537563
R23440 VGND.n7651 VGND.n7604 0.537563
R23441 VGND.n8187 VGND.n8157 0.537563
R23442 VGND.n8166 VGND.n8165 0.537563
R23443 VGND.n8160 VGND.n8159 0.537563
R23444 VGND.n8282 VGND.n8281 0.537563
R23445 VGND.n1285 VGND.n1149 0.537563
R23446 VGND.n1113 VGND.n1112 0.537563
R23447 VGND.n7384 VGND.n7383 0.537563
R23448 VGND.n7356 VGND.n809 0.537563
R23449 VGND.n7412 VGND.n805 0.537563
R23450 VGND.n7388 VGND.n7387 0.537563
R23451 VGND.n1494 VGND.n1489 0.537563
R23452 VGND.n6864 VGND.n6863 0.537563
R23453 VGND.n6875 VGND.n6874 0.537563
R23454 VGND.n6892 VGND.n1586 0.537563
R23455 VGND.n6828 VGND.n6827 0.537563
R23456 VGND.n6853 VGND.n6851 0.537563
R23457 VGND.n6329 VGND.n6257 0.537563
R23458 VGND.n6302 VGND.n6301 0.537563
R23459 VGND.n6376 VGND.n6360 0.537563
R23460 VGND.n5688 VGND.n5687 0.526527
R23461 VGND.n5651 VGND.n5650 0.526527
R23462 VGND.n5550 VGND.n5549 0.526527
R23463 VGND.n4622 VGND.n4621 0.526527
R23464 VGND.n4601 VGND.n4600 0.526527
R23465 VGND.n2956 VGND.n2955 0.526527
R23466 VGND.n3253 VGND.n3252 0.526527
R23467 VGND.n2728 VGND.n2667 0.526527
R23468 VGND.n8934 VGND.n8933 0.526527
R23469 VGND.n8516 VGND.n8515 0.526527
R23470 VGND.n8579 VGND.n247 0.526527
R23471 VGND.n3969 VGND.n3968 0.526527
R23472 VGND.n8643 VGND.n214 0.526527
R23473 VGND.n7794 VGND.n7793 0.526527
R23474 VGND.n7866 VGND.n7865 0.526527
R23475 VGND.n7931 VGND.n7930 0.526527
R23476 VGND.n369 VGND.n368 0.526527
R23477 VGND.n8232 VGND.n8231 0.526527
R23478 VGND.n791 VGND.n790 0.526527
R23479 VGND.n6240 VGND.n1689 0.526527
R23480 VGND.n2577 VGND.n2575 0.519731
R23481 VGND.n8266 VGND.n8265 0.507715
R23482 VGND.n7206 VGND.n7205 0.5005
R23483 VGND.n911 VGND.n909 0.482692
R23484 VGND.n25 VGND.n24 0.482692
R23485 VGND.n4323 VGND.n4322 0.477096
R23486 VGND.n8474 VGND.n8473 0.477096
R23487 VGND.n444 VGND.n441 0.448052
R23488 VGND.n6797 VGND.n6796 0.448052
R23489 VGND.n4563 VGND.n4562 0.438856
R23490 VGND.n1090 VGND.n1088 0.438856
R23491 VGND.n533 VGND.n532 0.43736
R23492 VGND.n3706 VGND.n3705 0.431476
R23493 VGND.n236 VGND.n235 0.427167
R23494 VGND.n2407 VGND.n2406 0.417891
R23495 VGND.n2479 VGND.n2339 0.417891
R23496 VGND.n2474 VGND.n2473 0.417891
R23497 VGND.n5140 VGND.n5134 0.417891
R23498 VGND.n5736 VGND.n5735 0.417891
R23499 VGND.n5587 VGND.n5586 0.417891
R23500 VGND.n5595 VGND.n5594 0.417891
R23501 VGND.n5971 VGND.n5970 0.417891
R23502 VGND.n5965 VGND.n1857 0.417891
R23503 VGND.n1807 VGND.n1801 0.417891
R23504 VGND.n1717 VGND.n1716 0.417891
R23505 VGND.n1721 VGND.n1710 0.417891
R23506 VGND.n6628 VGND.n1638 0.417891
R23507 VGND.n7151 VGND.n7150 0.417891
R23508 VGND.n7147 VGND.n1346 0.417891
R23509 VGND.n5063 VGND.n5062 0.417891
R23510 VGND.n5067 VGND.n4036 0.417891
R23511 VGND.n5047 VGND.n5046 0.417891
R23512 VGND.n4241 VGND.n4240 0.417891
R23513 VGND.n4245 VGND.n4239 0.417891
R23514 VGND.n4451 VGND.n4216 0.417891
R23515 VGND.n4656 VGND.n4552 0.417891
R23516 VGND.n4652 VGND.n4651 0.417891
R23517 VGND.n2925 VGND.n2924 0.417891
R23518 VGND.n2919 VGND.n2904 0.417891
R23519 VGND.n2054 VGND.n2053 0.417891
R23520 VGND.n2058 VGND.n2047 0.417891
R23521 VGND.n3676 VGND.n3675 0.417891
R23522 VGND.n3680 VGND.n3669 0.417891
R23523 VGND.n3795 VGND.n3794 0.417891
R23524 VGND.n3801 VGND.n3773 0.417891
R23525 VGND.n8620 VGND.n8619 0.417891
R23526 VGND.n8616 VGND.n225 0.417891
R23527 VGND.n1898 VGND.n1897 0.417891
R23528 VGND.n1904 VGND.n1901 0.417891
R23529 VGND.n8046 VGND.n492 0.417891
R23530 VGND.n8042 VGND.n496 0.417891
R23531 VGND.n7846 VGND.n7845 0.417891
R23532 VGND.n7850 VGND.n503 0.417891
R23533 VGND.n7310 VGND.n888 0.417891
R23534 VGND.n976 VGND.n904 0.417891
R23535 VGND.n7345 VGND.n816 0.417891
R23536 VGND.n7337 VGND.n7336 0.417891
R23537 VGND.n7339 VGND.n7338 0.417891
R23538 VGND.n7465 VGND.n7464 0.417891
R23539 VGND.n7469 VGND.n7458 0.417891
R23540 VGND.n6291 VGND.n6258 0.417891
R23541 VGND.n6287 VGND.n6261 0.417891
R23542 VGND.n6390 VGND.n6389 0.417891
R23543 VGND.n6385 VGND.n6353 0.417891
R23544 VGND.n6383 VGND.n6356 0.417891
R23545 VGND.n6379 VGND.n6359 0.417891
R23546 VGND.n2452 VGND.n2343 0.409011
R23547 VGND.n2446 VGND.n2346 0.409011
R23548 VGND.n2312 VGND.n2311 0.409011
R23549 VGND.n2569 VGND.n2568 0.409011
R23550 VGND.n2561 VGND.n2308 0.409011
R23551 VGND.n5155 VGND.n5154 0.409011
R23552 VGND.n5680 VGND.n5679 0.409011
R23553 VGND.n5636 VGND.n5635 0.409011
R23554 VGND.n5565 VGND.n5564 0.409011
R23555 VGND.n5571 VGND.n5497 0.409011
R23556 VGND.n5541 VGND.n5540 0.409011
R23557 VGND.n1809 VGND.n1808 0.409011
R23558 VGND.n1815 VGND.n1800 0.409011
R23559 VGND.n5408 VGND.n5407 0.409011
R23560 VGND.n1732 VGND.n1731 0.409011
R23561 VGND.n5097 VGND.n5088 0.409011
R23562 VGND.n7117 VGND.n1352 0.409011
R23563 VGND.n7101 VGND.n7100 0.409011
R23564 VGND.n4912 VGND.n4911 0.409011
R23565 VGND.n4918 VGND.n4087 0.409011
R23566 VGND.n4869 VGND.n4089 0.409011
R23567 VGND.n1423 VGND.n1422 0.409011
R23568 VGND.n1413 VGND.n1408 0.409011
R23569 VGND.n4118 VGND.n4117 0.409011
R23570 VGND.n4151 VGND.n4150 0.409011
R23571 VGND.n4693 VGND.n4161 0.409011
R23572 VGND.n4686 VGND.n4162 0.409011
R23573 VGND.n4672 VGND.n4166 0.409011
R23574 VGND.n4666 VGND.n4665 0.409011
R23575 VGND.n4295 VGND.n4294 0.409011
R23576 VGND.n4425 VGND.n4424 0.409011
R23577 VGND.n4478 VGND.n4477 0.409011
R23578 VGND.n4630 VGND.n4556 0.409011
R23579 VGND.n4612 VGND.n4568 0.409011
R23580 VGND.n1444 VGND.n1393 0.409011
R23581 VGND.n2964 VGND.n2963 0.409011
R23582 VGND.n2850 VGND.n2849 0.409011
R23583 VGND.n2856 VGND.n2751 0.409011
R23584 VGND.n2830 VGND.n2829 0.409011
R23585 VGND.n2837 VGND.n2836 0.409011
R23586 VGND.n2773 VGND.n2772 0.409011
R23587 VGND.n2789 VGND.n2758 0.409011
R23588 VGND.n3214 VGND.n3213 0.409011
R23589 VGND.n2695 VGND.n2694 0.409011
R23590 VGND.n3190 VGND.n3189 0.409011
R23591 VGND.n3189 VGND.n3188 0.409011
R23592 VGND.n8920 VGND.n8919 0.409011
R23593 VGND.n8960 VGND.n8959 0.409011
R23594 VGND.n8477 VGND.n8460 0.409011
R23595 VGND.n8467 VGND.n8461 0.409011
R23596 VGND.n8492 VGND.n8454 0.409011
R23597 VGND.n8485 VGND.n8455 0.409011
R23598 VGND.n8537 VGND.n8536 0.409011
R23599 VGND.n8536 VGND.n8535 0.409011
R23600 VGND.n240 VGND.n239 0.409011
R23601 VGND.n3977 VGND.n3881 0.409011
R23602 VGND.n8782 VGND.n162 0.409011
R23603 VGND.n8778 VGND.n165 0.409011
R23604 VGND.n8764 VGND.n171 0.409011
R23605 VGND.n8757 VGND.n8756 0.409011
R23606 VGND.n8750 VGND.n8749 0.409011
R23607 VGND.n8740 VGND.n8739 0.409011
R23608 VGND.n8615 VGND.n226 0.409011
R23609 VGND.n8381 VGND.n8342 0.409011
R23610 VGND.n1889 VGND.n1888 0.409011
R23611 VGND.n8037 VGND.n8036 0.409011
R23612 VGND.n8031 VGND.n7948 0.409011
R23613 VGND.n7805 VGND.n509 0.409011
R23614 VGND.n7940 VGND.n7893 0.409011
R23615 VGND.n7907 VGND.n7906 0.409011
R23616 VGND.n377 VGND.n342 0.409011
R23617 VGND.n704 VGND.n703 0.409011
R23618 VGND.n715 VGND.n690 0.409011
R23619 VGND.n7609 VGND.n7608 0.409011
R23620 VGND.n601 VGND.n600 0.409011
R23621 VGND.n673 VGND.n606 0.409011
R23622 VGND.n664 VGND.n607 0.409011
R23623 VGND.n8243 VGND.n455 0.409011
R23624 VGND.n975 VGND.n908 0.409011
R23625 VGND.n1216 VGND.n1215 0.409011
R23626 VGND.n1104 VGND.n1103 0.409011
R23627 VGND.n1111 VGND.n1007 0.409011
R23628 VGND.n1076 VGND.n1075 0.409011
R23629 VGND.n1082 VGND.n1081 0.409011
R23630 VGND.n7427 VGND.n788 0.409011
R23631 VGND.n1533 VGND.n1478 0.409011
R23632 VGND.n6911 VGND.n6910 0.409011
R23633 VGND.n6227 VGND.n6226 0.409011
R23634 VGND.n5364 VGND.n5363 0.406849
R23635 VGND.n7742 VGND.n7741 0.393674
R23636 VGND.n3572 VGND.n3571 0.388379
R23637 VGND.n3317 VGND.n2649 0.383542
R23638 VGND.n7328 VGND.n7327 0.3805
R23639 VGND.n7327 VGND.n841 0.3805
R23640 VGND.n7327 VGND.n7326 0.3805
R23641 VGND.n7298 VGND.n991 0.3805
R23642 VGND.n7298 VGND.n998 0.3805
R23643 VGND.n7300 VGND.n7298 0.3805
R23644 VGND.n6476 VGND.n1660 0.3805
R23645 VGND.n7291 VGND.n1321 0.3805
R23646 VGND.n7291 VGND.n1140 0.3805
R23647 VGND.n7291 VGND.n7290 0.3805
R23648 VGND.n7500 VGND.n7499 0.3805
R23649 VGND.n7500 VGND.n764 0.3805
R23650 VGND.n7500 VGND.n751 0.3805
R23651 VGND.n7134 VGND.n7133 0.376971
R23652 VGND.n7191 VGND.n1330 0.376971
R23653 VGND.n8634 VGND.n8633 0.376971
R23654 VGND.n8366 VGND.n8363 0.376971
R23655 VGND.n946 VGND.n945 0.376971
R23656 VGND.n9140 VGND.n9108 0.376971
R23657 VGND.n4960 VGND.n4959 0.374769
R23658 VGND.n5228 VGND.n5226 0.358542
R23659 VGND.n5256 VGND.n5255 0.358542
R23660 VGND.n5449 VGND.n5197 0.358542
R23661 VGND.n5377 VGND.n5376 0.358542
R23662 VGND.n6682 VGND.n1630 0.358542
R23663 VGND.n7005 VGND.n7004 0.358542
R23664 VGND.n2072 VGND.n2041 0.358542
R23665 VGND.n3088 VGND.n3087 0.358542
R23666 VGND.n8898 VGND.n8897 0.358542
R23667 VGND.n334 VGND.n333 0.358542
R23668 VGND.n7535 VGND.n7534 0.358542
R23669 VGND.n4548 VGND.n4170 0.357094
R23670 VGND.n2037 VGND.n2035 0.356928
R23671 VGND.n2035 VGND.n2032 0.356928
R23672 VGND.n9090 VGND.n45 0.356928
R23673 VGND.n9091 VGND.n9090 0.356928
R23674 VGND.n7566 VGND.n7565 0.354417
R23675 VGND.n829 VGND.n752 0.352216
R23676 VGND.n6206 VGND.n6204 0.352216
R23677 VGND.n2401 VGND.n2400 0.348326
R23678 VGND.n1716 VGND.n1715 0.348326
R23679 VGND.n5045 VGND.n5044 0.348326
R23680 VGND.n2053 VGND.n2052 0.348326
R23681 VGND.n3675 VGND.n3674 0.348326
R23682 VGND.n7464 VGND.n7463 0.348326
R23683 VGND.n7297 VGND.n7296 0.348099
R23684 VGND.n6202 VGND.n6201 0.347759
R23685 VGND.n7294 VGND.n7293 0.347759
R23686 VGND.n3575 VGND.n3574 0.345281
R23687 VGND.n6199 VGND.n6198 0.34507
R23688 VGND.n859 VGND.n842 0.342516
R23689 VGND.n1180 VGND.n895 0.342516
R23690 VGND.n7272 VGND.n7271 0.342516
R23691 VGND.n7450 VGND.n7449 0.342516
R23692 VGND.n6492 VGND.n6491 0.342503
R23693 VGND.n6955 VGND.n1553 0.3424
R23694 VGND.n6476 VGND.n6475 0.3424
R23695 VGND.n6476 VGND.n1663 0.341811
R23696 VGND.n6956 VGND.n6955 0.341811
R23697 VGND.n6789 VGND.n6787 0.341811
R23698 VGND.n6787 VGND.n6786 0.341811
R23699 VGND.n6208 VGND.n6207 0.341811
R23700 VGND.n1408 VGND.n1407 0.340926
R23701 VGND.n2869 VGND.n2866 0.340926
R23702 VGND.n1883 VGND.n1882 0.340926
R23703 VGND.n6166 VGND.n1696 0.31175
R23704 VGND.n6780 VGND.n6779 0.311379
R23705 VGND.n1612 VGND.n1611 0.311379
R23706 VGND.n6954 VGND.n6953 0.311321
R23707 VGND.n6195 VGND.n6194 0.311321
R23708 VGND.n4591 VGND.n4590 0.307349
R23709 VGND.n232 VGND.n231 0.307349
R23710 VGND.n2616 VGND.n2287 0.305262
R23711 VGND.n2597 VGND.n2288 0.305262
R23712 VGND.n2214 VGND.n2213 0.305262
R23713 VGND.n2172 VGND.n2171 0.305262
R23714 VGND.n2202 VGND.n2201 0.305262
R23715 VGND.n2212 VGND.n2175 0.305262
R23716 VGND.n9200 VGND.n9199 0.305262
R23717 VGND.n9185 VGND.n15 0.305262
R23718 VGND.n5224 VGND.n5223 0.305262
R23719 VGND.n5261 VGND.n5225 0.305262
R23720 VGND.n5429 VGND.n5428 0.305262
R23721 VGND.n5441 VGND.n5200 0.305262
R23722 VGND.n6707 VGND.n6706 0.305262
R23723 VGND.n5363 VGND.n5362 0.305262
R23724 VGND.n6613 VGND.n6612 0.305262
R23725 VGND.n6597 VGND.n1644 0.305262
R23726 VGND.n3444 VGND.n3443 0.305262
R23727 VGND.n3429 VGND.n2106 0.305262
R23728 VGND.n3415 VGND.n2114 0.305262
R23729 VGND.n3401 VGND.n2117 0.305262
R23730 VGND.n3399 VGND.n2118 0.305262
R23731 VGND.n3394 VGND.n2121 0.305262
R23732 VGND.n3393 VGND.n2122 0.305262
R23733 VGND.n2124 VGND.n2123 0.305262
R23734 VGND.n3311 VGND.n3310 0.305262
R23735 VGND.n3289 VGND.n2652 0.305262
R23736 VGND.n3662 VGND.n3661 0.305262
R23737 VGND.n3654 VGND.n3633 0.305262
R23738 VGND.n3653 VGND.n3636 0.305262
R23739 VGND.n3639 VGND.n3637 0.305262
R23740 VGND.n8871 VGND.n97 0.305262
R23741 VGND.n99 VGND.n98 0.305262
R23742 VGND.n8726 VGND.n189 0.305262
R23743 VGND.n8721 VGND.n192 0.305262
R23744 VGND.n1120 VGND.n1119 0.305262
R23745 VGND.n1293 VGND.n1146 0.305262
R23746 VGND.n1519 VGND.n1518 0.305262
R23747 VGND.n1499 VGND.n1486 0.305262
R23748 VGND.n7384 VGND.n7382 0.295551
R23749 VGND.n8258 VGND.n8256 0.294628
R23750 VGND.n5604 VGND.n5603 0.278761
R23751 VGND.n7845 VGND.n7844 0.278761
R23752 VGND VGND.n3446 0.274365
R23753 VGND VGND.n7669 0.274365
R23754 VGND.n2313 VGND.n2312 0.27284
R23755 VGND.n1737 VGND.n1735 0.27284
R23756 VGND.n4479 VGND.n4478 0.27284
R23757 VGND.n2898 VGND.n2897 0.27284
R23758 VGND.n8521 VGND.n8520 0.27284
R23759 VGND.n7920 VGND.n7907 0.27284
R23760 VGND.n1195 VGND.n1194 0.27284
R23761 VGND.n2276 VGND.n2275 0.269031
R23762 VGND.n7826 VGND.n7825 0.269031
R23763 VGND.n2305 VGND.n2304 0.263514
R23764 VGND.n5699 VGND.n5698 0.263514
R23765 VGND.n5662 VGND.n5470 0.263514
R23766 VGND.n5561 VGND.n5560 0.263514
R23767 VGND.n4615 VGND.n4565 0.263514
R23768 VGND.n4589 VGND.n4588 0.263514
R23769 VGND.n2943 VGND.n2899 0.263514
R23770 VGND.n3248 VGND.n3222 0.263514
R23771 VGND.n2718 VGND.n2717 0.263514
R23772 VGND.n8939 VGND.n79 0.263514
R23773 VGND.n8503 VGND.n8451 0.263514
R23774 VGND.n8574 VGND.n254 0.263514
R23775 VGND.n3957 VGND.n3956 0.263514
R23776 VGND.n8597 VGND.n8596 0.263514
R23777 VGND.n8638 VGND.n215 0.263514
R23778 VGND.n7871 VGND.n501 0.263514
R23779 VGND.n7926 VGND.n7901 0.263514
R23780 VGND.n358 VGND.n343 0.263514
R23781 VGND.n958 VGND.n914 0.263514
R23782 VGND.n1098 VGND.n1097 0.263514
R23783 VGND.n7413 VGND.n804 0.263514
R23784 VGND.n9151 VGND.n9101 0.263514
R23785 VGND.n8892 VGND.n8891 0.262616
R23786 VGND.n8888 VGND.n8887 0.262616
R23787 VGND.n7761 VGND.n535 0.262616
R23788 VGND.n534 VGND.n533 0.262616
R23789 VGND.n538 VGND.n537 0.262616
R23790 VGND.n4959 VGND.n4958 0.262488
R23791 VGND.n2297 VGND.n2296 0.259086
R23792 VGND.n2195 VGND.n2194 0.259086
R23793 VGND.n2200 VGND.n2179 0.259086
R23794 VGND.n5232 VGND.n5231 0.259086
R23795 VGND.n5238 VGND.n5233 0.259086
R23796 VGND.n5420 VGND.n5419 0.259086
R23797 VGND.n5427 VGND.n5203 0.259086
R23798 VGND.n6690 VGND.n6689 0.259086
R23799 VGND.n6695 VGND.n1627 0.259086
R23800 VGND.n7068 VGND.n7067 0.259086
R23801 VGND.n7061 VGND.n7003 0.259086
R23802 VGND.n3448 VGND.n3447 0.259086
R23803 VGND.n3422 VGND.n3421 0.259086
R23804 VGND.n3416 VGND.n2113 0.259086
R23805 VGND.n3323 VGND.n3322 0.259086
R23806 VGND.n3320 VGND.n3319 0.259086
R23807 VGND.n3058 VGND.n3057 0.259086
R23808 VGND.n3066 VGND.n3065 0.259086
R23809 VGND.n3691 VGND.n3690 0.259086
R23810 VGND.n8877 VGND.n8876 0.259086
R23811 VGND.n8872 VGND.n96 0.259086
R23812 VGND.n184 VGND.n183 0.259086
R23813 VGND.n8728 VGND.n188 0.259086
R23814 VGND.n8703 VGND.n8702 0.259086
R23815 VGND.n8644 VGND.n206 0.259086
R23816 VGND.n524 VGND.n523 0.259086
R23817 VGND.n7767 VGND.n528 0.259086
R23818 VGND.n402 VGND.n401 0.259086
R23819 VGND.n394 VGND.n332 0.259086
R23820 VGND.n7679 VGND.n7678 0.259086
R23821 VGND.n7671 VGND.n7670 0.259086
R23822 VGND.n5360 VGND.n5359 0.254468
R23823 VGND.n1311 VGND.n1310 0.254468
R23824 VGND.n2032 VGND 0.242831
R23825 VGND.n9091 VGND 0.242831
R23826 VGND.n2691 VGND.n2689 0.239569
R23827 VGND.n8380 VGND.n8379 0.239569
R23828 VGND.n5415 VGND.n5414 0.239569
R23829 VGND.n6196 VGND 0.239202
R23830 VGND.n5151 VGND.n5149 0.238116
R23831 VGND.n8966 VGND.n8965 0.237885
R23832 VGND.n8777 VGND.n8776 0.237885
R23833 VGND.n999 VGND 0.237242
R23834 VGND.n8263 VGND 0.236604
R23835 VGND VGND.n9202 0.236604
R23836 VGND.n6657 VGND.n6656 0.225061
R23837 VGND.n6671 VGND.n6668 0.225061
R23838 VGND.n4951 VGND.n4950 0.225061
R23839 VGND.n4961 VGND.n4960 0.225061
R23840 VGND.n4983 VGND.n4982 0.225061
R23841 VGND.n2802 VGND.n2801 0.225061
R23842 VGND.n2810 VGND.n2808 0.225061
R23843 VGND.n7855 VGND.n7854 0.225061
R23844 VGND.n7860 VGND.n502 0.225061
R23845 VGND.n231 VGND.n228 0.219678
R23846 VGND.n3573 VGND.n3572 0.215988
R23847 VGND.n4449 VGND.n4448 0.209196
R23848 VGND.n4450 VGND.n4449 0.209196
R23849 VGND.n2453 VGND.n2452 0.207909
R23850 VGND.n602 VGND.n601 0.204755
R23851 VGND.n6725 VGND.n6724 0.203675
R23852 VGND.n1132 VGND.n1131 0.203675
R23853 VGND.n3446 VGND 0.196835
R23854 VGND.n8263 VGND 0.196835
R23855 VGND.n7669 VGND 0.196835
R23856 VGND.n9202 VGND 0.196835
R23857 VGND.n3306 VGND.n3305 0.192021
R23858 VGND.n2037 VGND.n2036 0.1905
R23859 VGND.n2035 VGND.n2034 0.1905
R23860 VGND.n9090 VGND.n9089 0.1905
R23861 VGND.n9092 VGND.n9091 0.1905
R23862 VGND.n2632 VGND.n45 0.1905
R23863 VGND.n2876 VGND.n2875 0.180551
R23864 VGND.n4430 VGND 0.179673
R23865 VGND VGND.n1433 0.179673
R23866 VGND VGND.n1432 0.179673
R23867 VGND VGND.n8905 0.179673
R23868 VGND VGND.n8583 0.179673
R23869 VGND VGND.n1952 0.179673
R23870 VGND.n6855 VGND 0.179673
R23871 VGND VGND.n1522 0.179673
R23872 VGND VGND.n1521 0.179673
R23873 VGND.n6615 VGND 0.179673
R23874 VGND.n2587 VGND.n2586 0.179521
R23875 VGND.n2243 VGND.n2242 0.179521
R23876 VGND.n2185 VGND.n17 0.179521
R23877 VGND.n5260 VGND.n5226 0.179521
R23878 VGND.n5445 VGND.n5444 0.179521
R23879 VGND.n6678 VGND.n6677 0.179521
R23880 VGND.n7020 VGND.n7019 0.179521
R23881 VGND.n2068 VGND.n2067 0.179521
R23882 VGND.n3131 VGND.n3130 0.179521
R23883 VGND.n3169 VGND.n3168 0.179521
R23884 VGND.n3030 VGND.n3029 0.179521
R23885 VGND.n8893 VGND.n86 0.179521
R23886 VGND.n9017 VGND.n9016 0.179521
R23887 VGND.n522 VGND.n521 0.179521
R23888 VGND.n7762 VGND.n531 0.179521
R23889 VGND.n7814 VGND.n7813 0.179521
R23890 VGND.n7580 VGND.n7579 0.179521
R23891 VGND.n7587 VGND.n7584 0.179521
R23892 VGND.n7595 VGND.n7594 0.179521
R23893 VGND.n7666 VGND.n7665 0.179521
R23894 VGND.n8181 VGND.n8180 0.179521
R23895 VGND.n434 VGND.n433 0.179521
R23896 VGND.n7401 VGND.n7400 0.179521
R23897 VGND.n6872 VGND.n6871 0.179521
R23898 VGND VGND.n9122 0.178345
R23899 VGND.n7013 VGND 0.177989
R23900 VGND.n1410 VGND 0.177989
R23901 VGND VGND.n2911 0.177989
R23902 VGND.n8914 VGND 0.177989
R23903 VGND VGND.n2684 0.177989
R23904 VGND.n8463 VGND 0.177989
R23905 VGND.n8354 VGND 0.177989
R23906 VGND VGND.n352 0.177989
R23907 VGND VGND.n932 0.177989
R23908 VGND.n1491 VGND 0.177989
R23909 VGND.n5235 VGND 0.177989
R23910 VGND.n2302 VGND.n2301 0.175842
R23911 VGND.n2819 VGND.n2818 0.175842
R23912 VGND.n2721 VGND.n2720 0.175842
R23913 VGND.n8932 VGND.n8931 0.175842
R23914 VGND.n213 VGND.n212 0.175842
R23915 VGND.n8219 VGND.n8218 0.175842
R23916 VGND.n6249 VGND.n1688 0.175842
R23917 VGND.n3049 VGND.n3035 0.17139
R23918 VGND VGND.n4770 0.171212
R23919 VGND VGND.n4102 0.171212
R23920 VGND.n2049 VGND 0.171212
R23921 VGND.n3671 VGND 0.171212
R23922 VGND VGND.n3782 0.171212
R23923 VGND VGND.n1887 0.171212
R23924 VGND VGND.n695 0.171212
R23925 VGND.n7460 VGND 0.171212
R23926 VGND.n6118 VGND 0.171212
R23927 VGND.n1712 VGND 0.171212
R23928 VGND.n3486 VGND 0.171212
R23929 VGND.n3724 VGND.n3664 0.165322
R23930 VGND.n9210 VGND.n9203 0.165322
R23931 VGND.n5373 VGND 0.158415
R23932 VGND.n2594 VGND 0.158415
R23933 VGND.n2125 VGND.n2124 0.152881
R23934 VGND.n101 VGND.n99 0.152881
R23935 VGND.n3335 VGND.n118 0.151488
R23936 VGND.n8813 VGND.n8812 0.151488
R23937 VGND.n7717 VGND.n7716 0.151488
R23938 VGND.n4230 VGND.n4229 0.151488
R23939 VGND.n5835 VGND.n1658 0.151488
R23940 VGND.n3020 VGND.n3019 0.151488
R23941 VGND.n3023 VGND.n3022 0.151488
R23942 VGND.n7973 VGND.n7972 0.151488
R23943 VGND.n6990 VGND.n6989 0.151488
R23944 VGND.n5464 VGND.n5463 0.151488
R23945 VGND.n9067 VGND.n9066 0.151488
R23946 VGND.n202 VGND.n201 0.151488
R23947 VGND.n8113 VGND.n8112 0.151488
R23948 VGND.n4184 VGND.n4183 0.151488
R23949 VGND.n5489 VGND.n1614 0.151488
R23950 VGND.n3584 VGND.n3583 0.151488
R23951 VGND.n3730 VGND.n3729 0.151488
R23952 VGND.n1874 VGND.n1873 0.151488
R23953 VGND.n4752 VGND.n4751 0.151488
R23954 VGND.n6010 VGND.n6009 0.151488
R23955 VGND.n7507 VGND.n7506 0.151341
R23956 VGND.n6495 VGND.n6494 0.148403
R23957 VGND.n5298 VGND.n5297 0.148403
R23958 VGND.n6763 VGND.n6762 0.148403
R23959 VGND.n6091 VGND.n6090 0.148403
R23960 VGND.n4366 VGND.n4365 0.145562
R23961 VGND.n1570 VGND.n1569 0.145562
R23962 VGND.n4182 VGND.n4181 0.145562
R23963 VGND.n4705 VGND.n4704 0.145562
R23964 VGND.n5149 VGND 0.141328
R23965 VGND.n4058 VGND.n4057 0.141179
R23966 VGND.n1363 VGND.n1362 0.141179
R23967 VGND.n7254 VGND.n7253 0.141179
R23968 VGND.n4095 VGND.n4094 0.141179
R23969 VGND.n4430 VGND 0.140863
R23970 VGND.n1433 VGND 0.140863
R23971 VGND.n1432 VGND 0.140863
R23972 VGND.n8905 VGND 0.140863
R23973 VGND.n2689 VGND 0.140863
R23974 VGND.n8583 VGND 0.140863
R23975 VGND.n1952 VGND 0.140863
R23976 VGND.n8379 VGND 0.140863
R23977 VGND VGND.n6855 0.140863
R23978 VGND.n1522 VGND 0.140863
R23979 VGND.n1521 VGND 0.140863
R23980 VGND.n6615 VGND 0.140863
R23981 VGND VGND.n5415 0.140863
R23982 VGND.n7013 VGND 0.140584
R23983 VGND.n1410 VGND 0.140584
R23984 VGND.n2911 VGND 0.140584
R23985 VGND.n8914 VGND 0.140584
R23986 VGND.n8966 VGND 0.140584
R23987 VGND.n2684 VGND 0.140584
R23988 VGND.n8776 VGND 0.140584
R23989 VGND.n8463 VGND 0.140584
R23990 VGND.n8354 VGND 0.140584
R23991 VGND.n352 VGND 0.140584
R23992 VGND.n932 VGND 0.140584
R23993 VGND.n1491 VGND 0.140584
R23994 VGND.n5235 VGND 0.140584
R23995 VGND.n9122 VGND 0.140228
R23996 VGND.n2388 VGND.n2387 0.13963
R23997 VGND.n5756 VGND.n5755 0.13963
R23998 VGND.n1722 VGND.n1721 0.13963
R23999 VGND.n2059 VGND.n2058 0.13963
R24000 VGND.n3681 VGND.n3680 0.13963
R24001 VGND.n7470 VGND.n7469 0.13963
R24002 VGND.n9100 VGND.n9099 0.136751
R24003 VGND.n7106 VGND.n7105 0.13667
R24004 VGND.n4423 VGND.n4422 0.13667
R24005 VGND.n4511 VGND.n4510 0.13667
R24006 VGND.n1440 VGND.n1439 0.13667
R24007 VGND.n2786 VGND.n2784 0.13667
R24008 VGND.n8467 VGND.n8466 0.13667
R24009 VGND.n8537 VGND.n8534 0.13667
R24010 VGND.n176 VGND.n175 0.13667
R24011 VGND.n1192 VGND.n1191 0.13667
R24012 VGND.n1529 VGND.n1528 0.13667
R24013 VGND.n6935 VGND.n6934 0.13667
R24014 VGND.n518 VGND.n516 0.132007
R24015 VGND.n7789 VGND.n518 0.132007
R24016 VGND.n539 VGND.n538 0.131558
R24017 VGND.n3012 VGND.n2876 0.127051
R24018 VGND.n2647 VGND.n2646 0.126617
R24019 VGND.n100 VGND.n81 0.126617
R24020 VGND.n3638 VGND.n83 0.126304
R24021 VGND.n2036 VGND.n556 0.122994
R24022 VGND.n8437 VGND.n8436 0.122994
R24023 VGND.n2034 VGND.n2033 0.122994
R24024 VGND.n2038 VGND.n2031 0.122994
R24025 VGND VGND.n3424 0.120655
R24026 VGND.n3281 VGND 0.120655
R24027 VGND.n8879 VGND 0.120655
R24028 VGND VGND.n8737 0.120655
R24029 VGND.n6237 VGND 0.120655
R24030 VGND.n6673 VGND 0.120655
R24031 VGND.n6702 VGND 0.120655
R24032 VGND.n6703 VGND 0.120655
R24033 VGND.n4779 VGND.n4776 0.120292
R24034 VGND.n4783 VGND.n4779 0.120292
R24035 VGND.n4785 VGND.n4783 0.120292
R24036 VGND.n4793 VGND.n4789 0.120292
R24037 VGND.n4868 VGND.n4867 0.120292
R24038 VGND.n4875 VGND.n4871 0.120292
R24039 VGND.n4877 VGND.n4875 0.120292
R24040 VGND.n4881 VGND.n4877 0.120292
R24041 VGND.n4885 VGND.n4881 0.120292
R24042 VGND.n4886 VGND.n4885 0.120292
R24043 VGND.n4890 VGND.n4889 0.120292
R24044 VGND.n4900 VGND.n4894 0.120292
R24045 VGND.n4902 VGND.n4900 0.120292
R24046 VGND.n4906 VGND.n4905 0.120292
R24047 VGND.n4907 VGND.n4906 0.120292
R24048 VGND.n4915 VGND.n4913 0.120292
R24049 VGND.n4916 VGND.n4915 0.120292
R24050 VGND.n4917 VGND.n4916 0.120292
R24051 VGND.n4923 VGND.n4921 0.120292
R24052 VGND.n4925 VGND.n4923 0.120292
R24053 VGND.n4929 VGND.n4925 0.120292
R24054 VGND.n4931 VGND.n4929 0.120292
R24055 VGND.n4933 VGND.n4931 0.120292
R24056 VGND.n4935 VGND.n4933 0.120292
R24057 VGND.n4937 VGND.n4935 0.120292
R24058 VGND.n4940 VGND.n4937 0.120292
R24059 VGND.n4942 VGND.n4940 0.120292
R24060 VGND.n4943 VGND.n4942 0.120292
R24061 VGND.n4944 VGND.n4943 0.120292
R24062 VGND.n4954 VGND.n4952 0.120292
R24063 VGND.n5023 VGND.n5021 0.120292
R24064 VGND.n5024 VGND.n5023 0.120292
R24065 VGND.n5032 VGND.n5028 0.120292
R24066 VGND.n5036 VGND.n5032 0.120292
R24067 VGND.n5040 VGND.n5036 0.120292
R24068 VGND.n5041 VGND.n5040 0.120292
R24069 VGND.n5051 VGND.n5050 0.120292
R24070 VGND.n5057 VGND.n5056 0.120292
R24071 VGND.n5065 VGND.n5064 0.120292
R24072 VGND.n5066 VGND.n5065 0.120292
R24073 VGND.n5071 VGND.n5069 0.120292
R24074 VGND.n5073 VGND.n5071 0.120292
R24075 VGND.n5077 VGND.n5073 0.120292
R24076 VGND.n5078 VGND.n5077 0.120292
R24077 VGND.n4032 VGND.n4031 0.120292
R24078 VGND.n4031 VGND.n4030 0.120292
R24079 VGND.n4017 VGND.n4016 0.120292
R24080 VGND.n7189 VGND.n7188 0.120292
R24081 VGND.n7185 VGND.n7184 0.120292
R24082 VGND.n7179 VGND.n7178 0.120292
R24083 VGND.n7178 VGND.n7176 0.120292
R24084 VGND.n7176 VGND.n7174 0.120292
R24085 VGND.n7167 VGND.n7165 0.120292
R24086 VGND.n7165 VGND.n7164 0.120292
R24087 VGND.n7164 VGND.n7161 0.120292
R24088 VGND.n7156 VGND.n7155 0.120292
R24089 VGND.n7155 VGND.n7153 0.120292
R24090 VGND.n7152 VGND.n7149 0.120292
R24091 VGND.n7149 VGND.n7148 0.120292
R24092 VGND.n7145 VGND.n7144 0.120292
R24093 VGND.n7144 VGND.n7140 0.120292
R24094 VGND.n7136 VGND.n7135 0.120292
R24095 VGND.n7135 VGND.n7131 0.120292
R24096 VGND.n7131 VGND.n7129 0.120292
R24097 VGND.n7129 VGND.n7123 0.120292
R24098 VGND.n7116 VGND.n7115 0.120292
R24099 VGND.n7115 VGND.n7113 0.120292
R24100 VGND.n7069 VGND.n7066 0.120292
R24101 VGND.n7066 VGND.n7064 0.120292
R24102 VGND.n7064 VGND.n7062 0.120292
R24103 VGND.n7059 VGND.n7058 0.120292
R24104 VGND.n7058 VGND.n7057 0.120292
R24105 VGND.n7057 VGND.n7055 0.120292
R24106 VGND.n7055 VGND.n7052 0.120292
R24107 VGND.n7052 VGND.n7050 0.120292
R24108 VGND.n7050 VGND.n7046 0.120292
R24109 VGND.n7046 VGND.n7044 0.120292
R24110 VGND.n7041 VGND.n7040 0.120292
R24111 VGND.n7040 VGND.n7039 0.120292
R24112 VGND.n7039 VGND.n7037 0.120292
R24113 VGND.n7037 VGND.n7035 0.120292
R24114 VGND.n7035 VGND.n7033 0.120292
R24115 VGND.n7033 VGND.n7031 0.120292
R24116 VGND.n7031 VGND.n7029 0.120292
R24117 VGND.n7029 VGND.n7026 0.120292
R24118 VGND.n7026 VGND.n7023 0.120292
R24119 VGND.n7023 VGND.n7021 0.120292
R24120 VGND.n7021 VGND.n7017 0.120292
R24121 VGND.n4115 VGND.n4114 0.120292
R24122 VGND.n4123 VGND.n4119 0.120292
R24123 VGND.n4692 VGND.n4691 0.120292
R24124 VGND.n4691 VGND.n4690 0.120292
R24125 VGND.n4690 VGND.n4687 0.120292
R24126 VGND.n4683 VGND.n4682 0.120292
R24127 VGND.n4682 VGND.n4678 0.120292
R24128 VGND.n4678 VGND.n4674 0.120292
R24129 VGND.n4671 VGND.n4670 0.120292
R24130 VGND.n4670 VGND.n4669 0.120292
R24131 VGND.n4243 VGND.n4242 0.120292
R24132 VGND.n4244 VGND.n4243 0.120292
R24133 VGND.n4252 VGND.n4250 0.120292
R24134 VGND.n4254 VGND.n4252 0.120292
R24135 VGND.n4256 VGND.n4254 0.120292
R24136 VGND.n4260 VGND.n4256 0.120292
R24137 VGND.n4262 VGND.n4260 0.120292
R24138 VGND.n4264 VGND.n4262 0.120292
R24139 VGND.n4266 VGND.n4264 0.120292
R24140 VGND.n4269 VGND.n4266 0.120292
R24141 VGND.n4271 VGND.n4269 0.120292
R24142 VGND.n4272 VGND.n4271 0.120292
R24143 VGND.n4273 VGND.n4272 0.120292
R24144 VGND.n4282 VGND.n4276 0.120292
R24145 VGND.n4283 VGND.n4282 0.120292
R24146 VGND.n4289 VGND.n4286 0.120292
R24147 VGND.n4291 VGND.n4289 0.120292
R24148 VGND.n4292 VGND.n4291 0.120292
R24149 VGND.n4298 VGND.n4296 0.120292
R24150 VGND.n4385 VGND.n4383 0.120292
R24151 VGND.n4388 VGND.n4385 0.120292
R24152 VGND.n4397 VGND.n4395 0.120292
R24153 VGND.n4399 VGND.n4397 0.120292
R24154 VGND.n4401 VGND.n4399 0.120292
R24155 VGND.n4405 VGND.n4401 0.120292
R24156 VGND.n4407 VGND.n4405 0.120292
R24157 VGND.n4410 VGND.n4407 0.120292
R24158 VGND.n4412 VGND.n4410 0.120292
R24159 VGND.n4415 VGND.n4412 0.120292
R24160 VGND.n4417 VGND.n4415 0.120292
R24161 VGND.n4418 VGND.n4417 0.120292
R24162 VGND.n4427 VGND.n4426 0.120292
R24163 VGND.n4429 VGND.n4427 0.120292
R24164 VGND VGND.n4217 0.120292
R24165 VGND.n4454 VGND.n4444 0.120292
R24166 VGND.n4466 VGND.n4462 0.120292
R24167 VGND.n4468 VGND.n4466 0.120292
R24168 VGND.n4470 VGND.n4468 0.120292
R24169 VGND.n4471 VGND.n4470 0.120292
R24170 VGND.n4531 VGND.n4530 0.120292
R24171 VGND.n4533 VGND.n4531 0.120292
R24172 VGND.n4534 VGND.n4533 0.120292
R24173 VGND.n4536 VGND.n4535 0.120292
R24174 VGND.n4543 VGND.n4542 0.120292
R24175 VGND.n4544 VGND.n4543 0.120292
R24176 VGND.n4655 VGND 0.120292
R24177 VGND.n4649 VGND.n4647 0.120292
R24178 VGND.n4647 VGND.n4645 0.120292
R24179 VGND.n4645 VGND.n4641 0.120292
R24180 VGND.n4641 VGND.n4639 0.120292
R24181 VGND.n4633 VGND.n4629 0.120292
R24182 VGND.n4629 VGND.n4625 0.120292
R24183 VGND.n4625 VGND.n4623 0.120292
R24184 VGND.n4623 VGND.n4618 0.120292
R24185 VGND.n4618 VGND.n4617 0.120292
R24186 VGND.n4617 VGND.n4616 0.120292
R24187 VGND.n4611 VGND.n4610 0.120292
R24188 VGND.n4610 VGND.n4608 0.120292
R24189 VGND.n4608 VGND.n4606 0.120292
R24190 VGND.n4606 VGND.n4602 0.120292
R24191 VGND.n4602 VGND.n4599 0.120292
R24192 VGND.n4599 VGND.n4594 0.120292
R24193 VGND.n1448 VGND.n1447 0.120292
R24194 VGND.n1443 VGND.n1442 0.120292
R24195 VGND.n1442 VGND.n1441 0.120292
R24196 VGND.n1441 VGND.n1437 0.120292
R24197 VGND.n1430 VGND.n1429 0.120292
R24198 VGND.n1424 VGND.n1418 0.120292
R24199 VGND.n1418 VGND.n1417 0.120292
R24200 VGND.n1417 VGND.n1414 0.120292
R24201 VGND.n2056 VGND.n2055 0.120292
R24202 VGND.n2057 VGND.n2056 0.120292
R24203 VGND.n2063 VGND.n2062 0.120292
R24204 VGND.n2064 VGND.n2063 0.120292
R24205 VGND.n2071 VGND.n2070 0.120292
R24206 VGND.n3451 VGND.n3449 0.120292
R24207 VGND.n3445 VGND.n3441 0.120292
R24208 VGND.n3441 VGND.n3439 0.120292
R24209 VGND.n3439 VGND.n3437 0.120292
R24210 VGND.n3437 VGND.n3435 0.120292
R24211 VGND.n3435 VGND.n3432 0.120292
R24212 VGND.n3432 VGND.n3431 0.120292
R24213 VGND.n3431 VGND.n3430 0.120292
R24214 VGND.n3423 VGND.n3419 0.120292
R24215 VGND.n3419 VGND.n3418 0.120292
R24216 VGND.n3418 VGND.n3417 0.120292
R24217 VGND.n3414 VGND.n3413 0.120292
R24218 VGND.n3413 VGND.n3411 0.120292
R24219 VGND.n3411 VGND.n3409 0.120292
R24220 VGND.n3409 VGND.n3407 0.120292
R24221 VGND.n3407 VGND.n3404 0.120292
R24222 VGND.n3404 VGND.n3403 0.120292
R24223 VGND.n3403 VGND.n3402 0.120292
R24224 VGND.n3398 VGND.n3397 0.120292
R24225 VGND.n3397 VGND.n3396 0.120292
R24226 VGND.n3396 VGND.n3395 0.120292
R24227 VGND.n3392 VGND.n3391 0.120292
R24228 VGND.n3391 VGND.n3389 0.120292
R24229 VGND.n3389 VGND.n3387 0.120292
R24230 VGND.n3387 VGND.n3385 0.120292
R24231 VGND.n3324 VGND.n2645 0.120292
R24232 VGND.n2650 VGND.n2645 0.120292
R24233 VGND.n3316 VGND.n2651 0.120292
R24234 VGND.n3316 VGND.n3315 0.120292
R24235 VGND.n3315 VGND.n3314 0.120292
R24236 VGND.n3314 VGND.n3313 0.120292
R24237 VGND.n3312 VGND.n3298 0.120292
R24238 VGND.n3298 VGND.n3297 0.120292
R24239 VGND.n3297 VGND.n3296 0.120292
R24240 VGND.n3296 VGND.n3294 0.120292
R24241 VGND.n3294 VGND.n3292 0.120292
R24242 VGND.n3292 VGND.n3290 0.120292
R24243 VGND.n3287 VGND.n3286 0.120292
R24244 VGND.n3286 VGND.n3285 0.120292
R24245 VGND.n3279 VGND.n3278 0.120292
R24246 VGND.n3278 VGND.n3276 0.120292
R24247 VGND.n3276 VGND.n3272 0.120292
R24248 VGND.n3272 VGND.n3270 0.120292
R24249 VGND.n3261 VGND.n3260 0.120292
R24250 VGND.n3260 VGND.n3258 0.120292
R24251 VGND.n3258 VGND.n3256 0.120292
R24252 VGND.n3256 VGND.n3254 0.120292
R24253 VGND.n3254 VGND.n3251 0.120292
R24254 VGND.n3251 VGND.n3250 0.120292
R24255 VGND.n3250 VGND.n3249 0.120292
R24256 VGND.n3246 VGND.n3245 0.120292
R24257 VGND.n2788 VGND.n2787 0.120292
R24258 VGND.n2794 VGND.n2792 0.120292
R24259 VGND.n2795 VGND.n2794 0.120292
R24260 VGND.n2804 VGND.n2803 0.120292
R24261 VGND.n2805 VGND.n2804 0.120292
R24262 VGND.n2807 VGND.n2805 0.120292
R24263 VGND.n2811 VGND.n2807 0.120292
R24264 VGND.n2814 VGND.n2813 0.120292
R24265 VGND.n2823 VGND.n2821 0.120292
R24266 VGND.n2824 VGND.n2823 0.120292
R24267 VGND.n2832 VGND.n2831 0.120292
R24268 VGND.n2835 VGND.n2832 0.120292
R24269 VGND.n2838 VGND.n2835 0.120292
R24270 VGND.n2845 VGND.n2842 0.120292
R24271 VGND.n2846 VGND.n2845 0.120292
R24272 VGND.n2853 VGND.n2851 0.120292
R24273 VGND.n2854 VGND.n2853 0.120292
R24274 VGND.n2855 VGND.n2854 0.120292
R24275 VGND.n2861 VGND.n2858 0.120292
R24276 VGND.n2862 VGND.n2861 0.120292
R24277 VGND.n2873 VGND.n2871 0.120292
R24278 VGND.n2875 VGND.n2873 0.120292
R24279 VGND.n2961 VGND.n2960 0.120292
R24280 VGND.n2960 VGND.n2959 0.120292
R24281 VGND.n2959 VGND.n2957 0.120292
R24282 VGND.n2957 VGND.n2954 0.120292
R24283 VGND.n2954 VGND.n2949 0.120292
R24284 VGND.n2949 VGND.n2944 0.120292
R24285 VGND.n2941 VGND.n2940 0.120292
R24286 VGND.n2940 VGND.n2938 0.120292
R24287 VGND.n2938 VGND.n2934 0.120292
R24288 VGND.n2929 VGND.n2927 0.120292
R24289 VGND.n2926 VGND.n2921 0.120292
R24290 VGND.n2921 VGND.n2920 0.120292
R24291 VGND.n2914 VGND.n2912 0.120292
R24292 VGND.n3678 VGND.n3677 0.120292
R24293 VGND.n3679 VGND.n3678 0.120292
R24294 VGND.n3686 VGND.n3683 0.120292
R24295 VGND.n3687 VGND.n3686 0.120292
R24296 VGND.n3695 VGND.n3692 0.120292
R24297 VGND.n3663 VGND.n3657 0.120292
R24298 VGND.n3657 VGND.n3656 0.120292
R24299 VGND.n3656 VGND.n3655 0.120292
R24300 VGND.n3652 VGND.n3651 0.120292
R24301 VGND.n3651 VGND.n3650 0.120292
R24302 VGND.n3650 VGND.n3649 0.120292
R24303 VGND.n3649 VGND.n3646 0.120292
R24304 VGND.n3646 VGND.n3644 0.120292
R24305 VGND.n3644 VGND.n3642 0.120292
R24306 VGND.n3642 VGND.n3640 0.120292
R24307 VGND.n8899 VGND.n8895 0.120292
R24308 VGND.n8895 VGND.n8894 0.120292
R24309 VGND.n89 VGND.n88 0.120292
R24310 VGND.n8886 VGND.n89 0.120292
R24311 VGND.n8885 VGND.n8884 0.120292
R24312 VGND.n8884 VGND.n8883 0.120292
R24313 VGND.n8878 VGND.n8875 0.120292
R24314 VGND.n8875 VGND.n8874 0.120292
R24315 VGND.n8874 VGND.n8873 0.120292
R24316 VGND.n8870 VGND.n8869 0.120292
R24317 VGND.n8869 VGND.n8867 0.120292
R24318 VGND.n8867 VGND.n8865 0.120292
R24319 VGND.n8865 VGND.n8863 0.120292
R24320 VGND.n8922 VGND.n8921 0.120292
R24321 VGND.n8923 VGND.n8922 0.120292
R24322 VGND.n8936 VGND.n8935 0.120292
R24323 VGND.n8937 VGND.n8936 0.120292
R24324 VGND.n8938 VGND.n8937 0.120292
R24325 VGND.n8945 VGND.n8941 0.120292
R24326 VGND.n8949 VGND.n8945 0.120292
R24327 VGND.n8951 VGND.n8949 0.120292
R24328 VGND.n8954 VGND.n8951 0.120292
R24329 VGND.n8963 VGND.n8961 0.120292
R24330 VGND.n8965 VGND.n8963 0.120292
R24331 VGND.n8973 VGND.n8971 0.120292
R24332 VGND.n8976 VGND.n8973 0.120292
R24333 VGND.n8977 VGND.n8976 0.120292
R24334 VGND.n8986 VGND.n8984 0.120292
R24335 VGND.n8988 VGND.n8986 0.120292
R24336 VGND.n8990 VGND.n8988 0.120292
R24337 VGND.n8994 VGND.n8990 0.120292
R24338 VGND.n8996 VGND.n8994 0.120292
R24339 VGND.n8998 VGND.n8996 0.120292
R24340 VGND.n9000 VGND.n8998 0.120292
R24341 VGND.n9003 VGND.n9000 0.120292
R24342 VGND.n9005 VGND.n9003 0.120292
R24343 VGND.n9007 VGND.n9005 0.120292
R24344 VGND.n3047 VGND.n3045 0.120292
R24345 VGND.n3055 VGND.n3054 0.120292
R24346 VGND.n3060 VGND.n3059 0.120292
R24347 VGND.n3061 VGND.n3060 0.120292
R24348 VGND.n3067 VGND.n3061 0.120292
R24349 VGND.n3075 VGND.n3074 0.120292
R24350 VGND.n3081 VGND.n3079 0.120292
R24351 VGND.n3082 VGND.n3081 0.120292
R24352 VGND.n3083 VGND.n3082 0.120292
R24353 VGND.n3089 VGND.n3086 0.120292
R24354 VGND.n3091 VGND.n3089 0.120292
R24355 VGND.n3093 VGND.n3091 0.120292
R24356 VGND.n3096 VGND.n3093 0.120292
R24357 VGND.n3100 VGND.n3096 0.120292
R24358 VGND.n3101 VGND.n3100 0.120292
R24359 VGND.n3102 VGND.n3101 0.120292
R24360 VGND.n3110 VGND.n3106 0.120292
R24361 VGND.n3112 VGND.n3110 0.120292
R24362 VGND.n3114 VGND.n3112 0.120292
R24363 VGND.n3116 VGND.n3114 0.120292
R24364 VGND.n3118 VGND.n3116 0.120292
R24365 VGND.n3120 VGND.n3118 0.120292
R24366 VGND.n3122 VGND.n3120 0.120292
R24367 VGND.n3126 VGND.n3122 0.120292
R24368 VGND.n3128 VGND.n3126 0.120292
R24369 VGND.n3132 VGND.n3128 0.120292
R24370 VGND.n2736 VGND.n2732 0.120292
R24371 VGND.n2732 VGND.n2730 0.120292
R24372 VGND.n2726 VGND.n2668 0.120292
R24373 VGND.n2669 VGND.n2668 0.120292
R24374 VGND.n2715 VGND.n2714 0.120292
R24375 VGND.n2714 VGND.n2712 0.120292
R24376 VGND.n2712 VGND.n2708 0.120292
R24377 VGND.n2708 VGND.n2704 0.120292
R24378 VGND.n2704 VGND.n2700 0.120292
R24379 VGND.n2696 VGND.n2692 0.120292
R24380 VGND.n2692 VGND.n2691 0.120292
R24381 VGND.n2687 VGND.n2686 0.120292
R24382 VGND.n2686 VGND.n2685 0.120292
R24383 VGND.n3790 VGND.n3788 0.120292
R24384 VGND.n3791 VGND.n3790 0.120292
R24385 VGND.n3792 VGND.n3791 0.120292
R24386 VGND.n3851 VGND.n3850 0.120292
R24387 VGND.n3852 VGND.n3851 0.120292
R24388 VGND.n3857 VGND.n3856 0.120292
R24389 VGND.n3861 VGND.n3857 0.120292
R24390 VGND.n3863 VGND.n3861 0.120292
R24391 VGND.n3866 VGND.n3863 0.120292
R24392 VGND.n3870 VGND.n3866 0.120292
R24393 VGND.n3872 VGND.n3870 0.120292
R24394 VGND.n3874 VGND.n3872 0.120292
R24395 VGND.n3875 VGND.n3874 0.120292
R24396 VGND.n3976 VGND.n3975 0.120292
R24397 VGND.n3975 VGND.n3974 0.120292
R24398 VGND.n3974 VGND.n3972 0.120292
R24399 VGND.n3972 VGND.n3970 0.120292
R24400 VGND.n3970 VGND.n3967 0.120292
R24401 VGND.n3967 VGND.n3962 0.120292
R24402 VGND.n3962 VGND.n3958 0.120292
R24403 VGND.n3955 VGND.n3954 0.120292
R24404 VGND.n3950 VGND.n3949 0.120292
R24405 VGND.n3949 VGND.n3947 0.120292
R24406 VGND.n3947 VGND.n3941 0.120292
R24407 VGND.n3941 VGND.n3939 0.120292
R24408 VGND.n3939 VGND.n3937 0.120292
R24409 VGND.n3937 VGND.n3935 0.120292
R24410 VGND.n3935 VGND.n3933 0.120292
R24411 VGND.n3933 VGND.n3928 0.120292
R24412 VGND.n8770 VGND.n8769 0.120292
R24413 VGND.n8769 VGND.n8767 0.120292
R24414 VGND.n8763 VGND.n8762 0.120292
R24415 VGND.n8762 VGND.n8761 0.120292
R24416 VGND.n8761 VGND.n8758 0.120292
R24417 VGND.n8754 VGND.n8752 0.120292
R24418 VGND.n8751 VGND.n8748 0.120292
R24419 VGND.n8748 VGND.n8745 0.120292
R24420 VGND.n8745 VGND.n8743 0.120292
R24421 VGND.n8743 VGND.n8742 0.120292
R24422 VGND.n8732 VGND.n8731 0.120292
R24423 VGND.n8731 VGND.n8730 0.120292
R24424 VGND.n8730 VGND.n8729 0.120292
R24425 VGND.n8725 VGND.n8724 0.120292
R24426 VGND.n8724 VGND.n8723 0.120292
R24427 VGND.n8723 VGND.n8722 0.120292
R24428 VGND.n8648 VGND.n8645 0.120292
R24429 VGND.n8642 VGND.n8641 0.120292
R24430 VGND.n8641 VGND.n8640 0.120292
R24431 VGND.n8640 VGND.n8639 0.120292
R24432 VGND.n8635 VGND.n8631 0.120292
R24433 VGND.n8631 VGND.n8629 0.120292
R24434 VGND.n8629 VGND.n8628 0.120292
R24435 VGND.n8628 VGND.n8626 0.120292
R24436 VGND.n8621 VGND.n8618 0.120292
R24437 VGND.n8618 VGND.n8617 0.120292
R24438 VGND.n8614 VGND.n8613 0.120292
R24439 VGND.n8613 VGND.n8611 0.120292
R24440 VGND.n8611 VGND.n8608 0.120292
R24441 VGND.n8608 VGND.n8606 0.120292
R24442 VGND.n8606 VGND.n8605 0.120292
R24443 VGND.n8595 VGND.n238 0.120292
R24444 VGND.n8593 VGND.n8592 0.120292
R24445 VGND.n8592 VGND.n8588 0.120292
R24446 VGND.n8588 VGND.n8587 0.120292
R24447 VGND.n8578 VGND.n8577 0.120292
R24448 VGND.n8577 VGND.n8576 0.120292
R24449 VGND.n8576 VGND.n8575 0.120292
R24450 VGND.n8524 VGND.n8522 0.120292
R24451 VGND.n8522 VGND.n8519 0.120292
R24452 VGND.n8519 VGND.n8517 0.120292
R24453 VGND.n8517 VGND.n8514 0.120292
R24454 VGND.n8514 VGND.n8509 0.120292
R24455 VGND.n8509 VGND.n8504 0.120292
R24456 VGND.n8501 VGND.n8500 0.120292
R24457 VGND.n8500 VGND.n8498 0.120292
R24458 VGND.n8498 VGND.n8494 0.120292
R24459 VGND.n8491 VGND.n8490 0.120292
R24460 VGND.n8490 VGND.n8489 0.120292
R24461 VGND.n8489 VGND.n8486 0.120292
R24462 VGND.n8482 VGND.n8481 0.120292
R24463 VGND.n8480 VGND.n8479 0.120292
R24464 VGND.n8475 VGND.n8469 0.120292
R24465 VGND.n8469 VGND.n8468 0.120292
R24466 VGND.n1894 VGND.n1893 0.120292
R24467 VGND.n1895 VGND.n1894 0.120292
R24468 VGND.n1905 VGND.n1878 0.120292
R24469 VGND.n1950 VGND.n1948 0.120292
R24470 VGND.n1948 VGND.n1942 0.120292
R24471 VGND.n1942 VGND.n1940 0.120292
R24472 VGND.n1940 VGND.n1938 0.120292
R24473 VGND.n1938 VGND.n1934 0.120292
R24474 VGND.n1934 VGND.n1929 0.120292
R24475 VGND.n7804 VGND.n7803 0.120292
R24476 VGND.n7803 VGND.n7801 0.120292
R24477 VGND.n7801 VGND.n7797 0.120292
R24478 VGND.n7797 VGND.n7795 0.120292
R24479 VGND.n7795 VGND.n7792 0.120292
R24480 VGND.n7792 VGND.n7791 0.120292
R24481 VGND.n7791 VGND.n7790 0.120292
R24482 VGND.n7786 VGND.n7785 0.120292
R24483 VGND.n7785 VGND.n7784 0.120292
R24484 VGND.n7780 VGND.n7779 0.120292
R24485 VGND.n7779 VGND.n7777 0.120292
R24486 VGND.n7777 VGND.n7775 0.120292
R24487 VGND.n7775 VGND.n7773 0.120292
R24488 VGND.n7773 VGND.n7770 0.120292
R24489 VGND.n7770 VGND.n7769 0.120292
R24490 VGND.n7769 VGND.n7768 0.120292
R24491 VGND.n7765 VGND.n7764 0.120292
R24492 VGND.n7764 VGND.n7763 0.120292
R24493 VGND.n7820 VGND.n7819 0.120292
R24494 VGND.n7828 VGND.n7827 0.120292
R24495 VGND.n7829 VGND.n7828 0.120292
R24496 VGND.n7839 VGND.n7838 0.120292
R24497 VGND.n7848 VGND.n7847 0.120292
R24498 VGND.n7857 VGND.n7856 0.120292
R24499 VGND.n7858 VGND.n7857 0.120292
R24500 VGND.n7859 VGND.n7858 0.120292
R24501 VGND.n7868 VGND.n7867 0.120292
R24502 VGND.n7869 VGND.n7868 0.120292
R24503 VGND.n7877 VGND.n7873 0.120292
R24504 VGND.n7879 VGND.n7877 0.120292
R24505 VGND.n7881 VGND.n7879 0.120292
R24506 VGND.n7886 VGND.n7881 0.120292
R24507 VGND.n7888 VGND.n7886 0.120292
R24508 VGND.n7939 VGND.n7938 0.120292
R24509 VGND.n7938 VGND.n7936 0.120292
R24510 VGND.n7936 VGND.n7934 0.120292
R24511 VGND.n7934 VGND.n7932 0.120292
R24512 VGND.n7932 VGND.n7929 0.120292
R24513 VGND.n7929 VGND.n7928 0.120292
R24514 VGND.n7928 VGND.n7927 0.120292
R24515 VGND.n7923 VGND.n7922 0.120292
R24516 VGND.n8061 VGND.n8059 0.120292
R24517 VGND.n8059 VGND.n8057 0.120292
R24518 VGND.n8057 VGND.n8056 0.120292
R24519 VGND.n8051 VGND.n8050 0.120292
R24520 VGND.n8050 VGND.n8048 0.120292
R24521 VGND.n8045 VGND.n8044 0.120292
R24522 VGND.n8038 VGND.n8035 0.120292
R24523 VGND.n8035 VGND.n8033 0.120292
R24524 VGND.n8033 VGND.n8032 0.120292
R24525 VGND.n8028 VGND.n8027 0.120292
R24526 VGND.n8023 VGND.n8019 0.120292
R24527 VGND.n8019 VGND.n8018 0.120292
R24528 VGND.n8018 VGND.n8016 0.120292
R24529 VGND.n8016 VGND.n8015 0.120292
R24530 VGND.n8015 VGND.n8013 0.120292
R24531 VGND.n8013 VGND.n8009 0.120292
R24532 VGND.n8009 VGND.n8008 0.120292
R24533 VGND.n8008 VGND.n8006 0.120292
R24534 VGND.n8006 VGND.n8002 0.120292
R24535 VGND.n7998 VGND.n7997 0.120292
R24536 VGND.n7997 VGND.n7996 0.120292
R24537 VGND.n7996 VGND.n7995 0.120292
R24538 VGND.n7995 VGND.n7993 0.120292
R24539 VGND.n7993 VGND.n7992 0.120292
R24540 VGND.n7992 VGND.n7990 0.120292
R24541 VGND.n8401 VGND.n8400 0.120292
R24542 VGND.n8400 VGND.n8398 0.120292
R24543 VGND.n8398 VGND.n8394 0.120292
R24544 VGND.n8388 VGND.n8380 0.120292
R24545 VGND.n8377 VGND.n8375 0.120292
R24546 VGND.n8367 VGND.n8361 0.120292
R24547 VGND.n8361 VGND.n8359 0.120292
R24548 VGND.n708 VGND.n706 0.120292
R24549 VGND.n712 VGND.n708 0.120292
R24550 VGND.n713 VGND.n712 0.120292
R24551 VGND.n714 VGND.n713 0.120292
R24552 VGND.n7567 VGND.n7563 0.120292
R24553 VGND.n7571 VGND.n7567 0.120292
R24554 VGND.n7572 VGND.n7571 0.120292
R24555 VGND.n7578 VGND.n7577 0.120292
R24556 VGND.n7581 VGND.n7578 0.120292
R24557 VGND.n7589 VGND.n7588 0.120292
R24558 VGND.n7591 VGND.n7589 0.120292
R24559 VGND.n7593 VGND.n7591 0.120292
R24560 VGND.n7596 VGND.n7593 0.120292
R24561 VGND.n7597 VGND.n7596 0.120292
R24562 VGND.n7680 VGND.n7674 0.120292
R24563 VGND.n7674 VGND.n7673 0.120292
R24564 VGND.n7673 VGND.n7672 0.120292
R24565 VGND.n7664 VGND.n7663 0.120292
R24566 VGND.n7663 VGND.n7661 0.120292
R24567 VGND.n7661 VGND.n7658 0.120292
R24568 VGND.n7658 VGND.n7655 0.120292
R24569 VGND.n7655 VGND.n7653 0.120292
R24570 VGND.n7653 VGND.n7652 0.120292
R24571 VGND.n7649 VGND.n7648 0.120292
R24572 VGND.n7648 VGND.n7646 0.120292
R24573 VGND.n7646 VGND.n7641 0.120292
R24574 VGND.n7641 VGND.n7639 0.120292
R24575 VGND.n676 VGND.n672 0.120292
R24576 VGND.n672 VGND.n671 0.120292
R24577 VGND.n671 VGND.n667 0.120292
R24578 VGND.n667 VGND.n665 0.120292
R24579 VGND.n662 VGND.n661 0.120292
R24580 VGND.n661 VGND.n659 0.120292
R24581 VGND.n659 VGND.n653 0.120292
R24582 VGND.n650 VGND.n649 0.120292
R24583 VGND.n649 VGND.n645 0.120292
R24584 VGND.n645 VGND.n644 0.120292
R24585 VGND.n644 VGND.n642 0.120292
R24586 VGND.n642 VGND.n641 0.120292
R24587 VGND.n641 VGND.n639 0.120292
R24588 VGND.n639 VGND.n635 0.120292
R24589 VGND.n635 VGND.n631 0.120292
R24590 VGND.n631 VGND.n629 0.120292
R24591 VGND.n629 VGND.n625 0.120292
R24592 VGND.n625 VGND.n624 0.120292
R24593 VGND.n623 VGND.n621 0.120292
R24594 VGND.n8250 VGND.n8248 0.120292
R24595 VGND.n8247 VGND.n8245 0.120292
R24596 VGND.n8242 VGND.n8241 0.120292
R24597 VGND.n8241 VGND.n8237 0.120292
R24598 VGND.n8237 VGND.n8235 0.120292
R24599 VGND.n8235 VGND.n8233 0.120292
R24600 VGND.n8233 VGND.n8230 0.120292
R24601 VGND.n8230 VGND.n8223 0.120292
R24602 VGND.n8186 VGND.n8185 0.120292
R24603 VGND.n8185 VGND.n8184 0.120292
R24604 VGND.n8184 VGND.n8182 0.120292
R24605 VGND.n8182 VGND.n8178 0.120292
R24606 VGND.n8175 VGND.n8174 0.120292
R24607 VGND.n8173 VGND.n8168 0.120292
R24608 VGND.n8168 VGND.n8167 0.120292
R24609 VGND.n8167 VGND.n8163 0.120292
R24610 VGND.n8163 VGND.n8161 0.120292
R24611 VGND.n8262 VGND.n8261 0.120292
R24612 VGND.n8272 VGND.n8269 0.120292
R24613 VGND.n8273 VGND.n8272 0.120292
R24614 VGND.n8279 VGND.n8278 0.120292
R24615 VGND.n8285 VGND.n8283 0.120292
R24616 VGND.n8289 VGND.n8285 0.120292
R24617 VGND.n8291 VGND.n8289 0.120292
R24618 VGND.n8293 VGND.n8291 0.120292
R24619 VGND.n8295 VGND.n8293 0.120292
R24620 VGND.n8297 VGND.n8295 0.120292
R24621 VGND.n8299 VGND.n8297 0.120292
R24622 VGND.n8302 VGND.n8299 0.120292
R24623 VGND.n8305 VGND.n8302 0.120292
R24624 VGND.n8306 VGND.n8305 0.120292
R24625 VGND.n8307 VGND.n8306 0.120292
R24626 VGND.n403 VGND.n400 0.120292
R24627 VGND.n400 VGND.n398 0.120292
R24628 VGND.n398 VGND.n395 0.120292
R24629 VGND.n392 VGND.n391 0.120292
R24630 VGND.n391 VGND.n390 0.120292
R24631 VGND.n390 VGND.n388 0.120292
R24632 VGND.n388 VGND.n386 0.120292
R24633 VGND.n380 VGND.n379 0.120292
R24634 VGND.n376 VGND.n375 0.120292
R24635 VGND.n375 VGND.n374 0.120292
R24636 VGND.n374 VGND.n372 0.120292
R24637 VGND.n372 VGND.n370 0.120292
R24638 VGND.n370 VGND.n367 0.120292
R24639 VGND.n367 VGND.n362 0.120292
R24640 VGND.n362 VGND.n359 0.120292
R24641 VGND.n355 VGND.n354 0.120292
R24642 VGND.n354 VGND.n353 0.120292
R24643 VGND.n7467 VGND.n7466 0.120292
R24644 VGND.n7468 VGND.n7467 0.120292
R24645 VGND.n7476 VGND.n7472 0.120292
R24646 VGND.n7477 VGND.n7476 0.120292
R24647 VGND.n7482 VGND.n7481 0.120292
R24648 VGND.n7424 VGND.n7423 0.120292
R24649 VGND.n7423 VGND.n7422 0.120292
R24650 VGND.n7422 VGND.n7417 0.120292
R24651 VGND.n7417 VGND.n7414 0.120292
R24652 VGND.n7410 VGND.n7407 0.120292
R24653 VGND.n7407 VGND.n7406 0.120292
R24654 VGND.n7406 VGND.n7404 0.120292
R24655 VGND.n7404 VGND.n7402 0.120292
R24656 VGND.n7402 VGND.n7398 0.120292
R24657 VGND.n7398 VGND.n7396 0.120292
R24658 VGND.n7391 VGND.n7390 0.120292
R24659 VGND.n7385 VGND.n7381 0.120292
R24660 VGND.n7381 VGND.n7379 0.120292
R24661 VGND.n7379 VGND.n7377 0.120292
R24662 VGND.n7377 VGND.n7375 0.120292
R24663 VGND.n7375 VGND.n7371 0.120292
R24664 VGND.n7371 VGND.n7369 0.120292
R24665 VGND.n7369 VGND.n7367 0.120292
R24666 VGND.n7367 VGND.n7365 0.120292
R24667 VGND.n7365 VGND.n7360 0.120292
R24668 VGND.n7360 VGND.n7358 0.120292
R24669 VGND.n7358 VGND.n7357 0.120292
R24670 VGND.n7354 VGND.n7353 0.120292
R24671 VGND.n7353 VGND.n7351 0.120292
R24672 VGND.n7350 VGND.n7349 0.120292
R24673 VGND.n7349 VGND.n7348 0.120292
R24674 VGND.n7348 VGND.n7347 0.120292
R24675 VGND.n7344 VGND.n7343 0.120292
R24676 VGND.n1027 VGND.n1025 0.120292
R24677 VGND.n1028 VGND.n1027 0.120292
R24678 VGND.n1034 VGND.n1033 0.120292
R24679 VGND.n1039 VGND.n1037 0.120292
R24680 VGND.n1044 VGND.n1039 0.120292
R24681 VGND.n1046 VGND.n1044 0.120292
R24682 VGND.n1049 VGND.n1046 0.120292
R24683 VGND.n1054 VGND.n1051 0.120292
R24684 VGND.n1056 VGND.n1054 0.120292
R24685 VGND.n1060 VGND.n1056 0.120292
R24686 VGND.n1064 VGND.n1060 0.120292
R24687 VGND.n1068 VGND.n1064 0.120292
R24688 VGND.n1070 VGND.n1068 0.120292
R24689 VGND.n1079 VGND.n1077 0.120292
R24690 VGND.n1083 VGND.n1079 0.120292
R24691 VGND.n1084 VGND.n1083 0.120292
R24692 VGND.n1092 VGND.n1084 0.120292
R24693 VGND.n1094 VGND.n1093 0.120292
R24694 VGND.n1108 VGND.n1105 0.120292
R24695 VGND.n1109 VGND.n1108 0.120292
R24696 VGND.n1110 VGND.n1109 0.120292
R24697 VGND.n1115 VGND.n1114 0.120292
R24698 VGND.n1116 VGND.n1115 0.120292
R24699 VGND.n1123 VGND.n1121 0.120292
R24700 VGND.n1125 VGND.n1123 0.120292
R24701 VGND.n1288 VGND.n1287 0.120292
R24702 VGND.n1283 VGND.n1282 0.120292
R24703 VGND.n1282 VGND.n1280 0.120292
R24704 VGND.n1280 VGND.n1278 0.120292
R24705 VGND.n1278 VGND.n1277 0.120292
R24706 VGND.n1274 VGND.n1273 0.120292
R24707 VGND.n1270 VGND.n1265 0.120292
R24708 VGND.n1265 VGND.n1263 0.120292
R24709 VGND.n1258 VGND.n1256 0.120292
R24710 VGND.n1251 VGND.n1250 0.120292
R24711 VGND.n1250 VGND.n1244 0.120292
R24712 VGND.n1239 VGND.n1238 0.120292
R24713 VGND.n1238 VGND.n1234 0.120292
R24714 VGND.n1234 VGND.n1230 0.120292
R24715 VGND.n1230 VGND.n1226 0.120292
R24716 VGND.n1220 VGND.n1219 0.120292
R24717 VGND.n1217 VGND.n1214 0.120292
R24718 VGND.n1214 VGND.n1211 0.120292
R24719 VGND.n1211 VGND.n1209 0.120292
R24720 VGND.n1209 VGND.n1205 0.120292
R24721 VGND.n974 VGND.n973 0.120292
R24722 VGND.n973 VGND.n972 0.120292
R24723 VGND.n969 VGND.n968 0.120292
R24724 VGND.n968 VGND.n967 0.120292
R24725 VGND.n967 VGND.n962 0.120292
R24726 VGND.n962 VGND.n959 0.120292
R24727 VGND.n955 VGND.n954 0.120292
R24728 VGND.n954 VGND.n952 0.120292
R24729 VGND.n952 VGND.n950 0.120292
R24730 VGND.n943 VGND.n942 0.120292
R24731 VGND.n937 VGND.n936 0.120292
R24732 VGND.n936 VGND.n935 0.120292
R24733 VGND.n935 VGND.n934 0.120292
R24734 VGND.n934 VGND.n933 0.120292
R24735 VGND.n6124 VGND.n6122 0.120292
R24736 VGND.n6128 VGND.n6124 0.120292
R24737 VGND.n6130 VGND.n6128 0.120292
R24738 VGND.n6134 VGND.n6130 0.120292
R24739 VGND.n6135 VGND.n6134 0.120292
R24740 VGND.n6140 VGND.n6138 0.120292
R24741 VGND.n6145 VGND.n6140 0.120292
R24742 VGND.n6229 VGND.n6228 0.120292
R24743 VGND.n6231 VGND.n6229 0.120292
R24744 VGND.n6231 VGND.n6230 0.120292
R24745 VGND.n6243 VGND.n6242 0.120292
R24746 VGND.n6254 VGND.n6253 0.120292
R24747 VGND.n6334 VGND.n6333 0.120292
R24748 VGND.n6328 VGND.n6327 0.120292
R24749 VGND.n6327 VGND.n6326 0.120292
R24750 VGND.n6326 VGND.n6324 0.120292
R24751 VGND.n6324 VGND.n6322 0.120292
R24752 VGND.n6322 VGND.n6318 0.120292
R24753 VGND.n6318 VGND.n6316 0.120292
R24754 VGND.n6316 VGND.n6314 0.120292
R24755 VGND.n6314 VGND.n6311 0.120292
R24756 VGND.n6311 VGND.n6309 0.120292
R24757 VGND.n6309 VGND.n6307 0.120292
R24758 VGND.n6307 VGND.n6305 0.120292
R24759 VGND.n6304 VGND.n6299 0.120292
R24760 VGND.n6299 VGND.n6293 0.120292
R24761 VGND.n6290 VGND.n6289 0.120292
R24762 VGND.n6289 VGND.n6288 0.120292
R24763 VGND.n6283 VGND.n6281 0.120292
R24764 VGND.n6452 VGND.n6451 0.120292
R24765 VGND.n6451 VGND.n6447 0.120292
R24766 VGND.n6444 VGND.n6443 0.120292
R24767 VGND.n6443 VGND.n6441 0.120292
R24768 VGND.n6441 VGND.n6435 0.120292
R24769 VGND.n6435 VGND.n6433 0.120292
R24770 VGND.n6433 VGND.n6432 0.120292
R24771 VGND.n6432 VGND.n6430 0.120292
R24772 VGND.n6430 VGND.n6424 0.120292
R24773 VGND.n6424 VGND.n6422 0.120292
R24774 VGND.n6422 VGND.n6421 0.120292
R24775 VGND.n6421 VGND.n6419 0.120292
R24776 VGND.n6419 VGND.n6415 0.120292
R24777 VGND.n6415 VGND.n6411 0.120292
R24778 VGND.n6411 VGND.n6409 0.120292
R24779 VGND.n6409 VGND.n6404 0.120292
R24780 VGND.n6404 VGND.n6402 0.120292
R24781 VGND.n6402 VGND.n6396 0.120292
R24782 VGND.n6393 VGND.n6392 0.120292
R24783 VGND.n6391 VGND.n6387 0.120292
R24784 VGND.n6387 VGND.n6386 0.120292
R24785 VGND.n6382 VGND.n6381 0.120292
R24786 VGND.n6381 VGND.n6380 0.120292
R24787 VGND.n6375 VGND.n6374 0.120292
R24788 VGND.n6374 VGND.n6372 0.120292
R24789 VGND.n6372 VGND.n6370 0.120292
R24790 VGND.n6370 VGND.n6368 0.120292
R24791 VGND.n6368 VGND.n6364 0.120292
R24792 VGND.n6364 VGND.n6362 0.120292
R24793 VGND.n6362 VGND.n1595 0.120292
R24794 VGND.n6835 VGND.n6834 0.120292
R24795 VGND.n6837 VGND.n6835 0.120292
R24796 VGND.n6841 VGND.n6837 0.120292
R24797 VGND.n6843 VGND.n6841 0.120292
R24798 VGND.n6847 VGND.n6843 0.120292
R24799 VGND.n6850 VGND.n6847 0.120292
R24800 VGND.n6854 VGND.n6850 0.120292
R24801 VGND.n6860 VGND.n6859 0.120292
R24802 VGND.n6866 VGND.n6865 0.120292
R24803 VGND.n6868 VGND.n6866 0.120292
R24804 VGND.n6870 VGND.n6868 0.120292
R24805 VGND.n6873 VGND.n6870 0.120292
R24806 VGND.n6878 VGND.n6876 0.120292
R24807 VGND.n6882 VGND.n6878 0.120292
R24808 VGND.n6885 VGND.n6882 0.120292
R24809 VGND.n6889 VGND.n6885 0.120292
R24810 VGND.n6890 VGND.n6889 0.120292
R24811 VGND.n6891 VGND.n6890 0.120292
R24812 VGND.n6895 VGND.n6894 0.120292
R24813 VGND.n6901 VGND.n6899 0.120292
R24814 VGND.n6907 VGND.n6901 0.120292
R24815 VGND.n6908 VGND.n6907 0.120292
R24816 VGND.n6914 VGND.n6912 0.120292
R24817 VGND.n6918 VGND.n6914 0.120292
R24818 VGND.n6920 VGND.n6918 0.120292
R24819 VGND.n6922 VGND.n6920 0.120292
R24820 VGND.n1532 VGND.n1531 0.120292
R24821 VGND.n1531 VGND.n1530 0.120292
R24822 VGND.n1530 VGND.n1526 0.120292
R24823 VGND.n1520 VGND.n1514 0.120292
R24824 VGND.n1514 VGND.n1513 0.120292
R24825 VGND.n1513 VGND.n1512 0.120292
R24826 VGND.n1512 VGND.n1510 0.120292
R24827 VGND.n1510 VGND.n1507 0.120292
R24828 VGND.n1507 VGND.n1505 0.120292
R24829 VGND.n1505 VGND.n1503 0.120292
R24830 VGND.n1503 VGND.n1500 0.120292
R24831 VGND.n1497 VGND.n1496 0.120292
R24832 VGND.n1496 VGND.n1495 0.120292
R24833 VGND.n1719 VGND.n1718 0.120292
R24834 VGND.n1720 VGND.n1719 0.120292
R24835 VGND.n1728 VGND.n1724 0.120292
R24836 VGND.n1729 VGND.n1728 0.120292
R24837 VGND.n1738 VGND.n1734 0.120292
R24838 VGND.n6052 VGND.n6051 0.120292
R24839 VGND.n6051 VGND.n6049 0.120292
R24840 VGND.n6049 VGND.n6047 0.120292
R24841 VGND.n6047 VGND.n6041 0.120292
R24842 VGND.n6041 VGND.n6037 0.120292
R24843 VGND.n6033 VGND.n6032 0.120292
R24844 VGND.n6032 VGND.n6030 0.120292
R24845 VGND.n6030 VGND.n6026 0.120292
R24846 VGND.n6026 VGND.n6025 0.120292
R24847 VGND.n6021 VGND.n6020 0.120292
R24848 VGND.n6614 VGND.n6611 0.120292
R24849 VGND.n6611 VGND.n6609 0.120292
R24850 VGND.n6609 VGND.n6607 0.120292
R24851 VGND.n6607 VGND.n6605 0.120292
R24852 VGND.n6605 VGND.n6603 0.120292
R24853 VGND.n6603 VGND.n6600 0.120292
R24854 VGND.n6600 VGND.n6599 0.120292
R24855 VGND.n6599 VGND.n6598 0.120292
R24856 VGND.n6595 VGND.n6594 0.120292
R24857 VGND.n6594 VGND.n6593 0.120292
R24858 VGND.n6590 VGND.n6589 0.120292
R24859 VGND.n6586 VGND.n6585 0.120292
R24860 VGND.n6582 VGND.n6581 0.120292
R24861 VGND.n6581 VGND.n6577 0.120292
R24862 VGND.n6639 VGND.n6638 0.120292
R24863 VGND.n6644 VGND.n6642 0.120292
R24864 VGND.n6649 VGND.n6644 0.120292
R24865 VGND.n6651 VGND.n6649 0.120292
R24866 VGND.n6652 VGND.n6651 0.120292
R24867 VGND.n6660 VGND.n6658 0.120292
R24868 VGND.n6662 VGND.n6660 0.120292
R24869 VGND.n6663 VGND.n6662 0.120292
R24870 VGND.n6664 VGND.n6663 0.120292
R24871 VGND.n6672 VGND.n6664 0.120292
R24872 VGND.n6681 VGND.n6680 0.120292
R24873 VGND.n6685 VGND.n6684 0.120292
R24874 VGND.n6686 VGND.n6685 0.120292
R24875 VGND.n6692 VGND.n6691 0.120292
R24876 VGND.n6693 VGND.n6692 0.120292
R24877 VGND.n6694 VGND.n6693 0.120292
R24878 VGND.n6710 VGND.n6708 0.120292
R24879 VGND.n6712 VGND.n6710 0.120292
R24880 VGND.n6714 VGND.n6712 0.120292
R24881 VGND.n6716 VGND.n6714 0.120292
R24882 VGND.n6719 VGND.n6716 0.120292
R24883 VGND.n5380 VGND.n5379 0.120292
R24884 VGND.n5382 VGND.n5380 0.120292
R24885 VGND.n5384 VGND.n5382 0.120292
R24886 VGND.n5386 VGND.n5384 0.120292
R24887 VGND.n5391 VGND.n5386 0.120292
R24888 VGND.n5393 VGND.n5391 0.120292
R24889 VGND.n5395 VGND.n5393 0.120292
R24890 VGND.n5397 VGND.n5395 0.120292
R24891 VGND.n5400 VGND.n5397 0.120292
R24892 VGND.n5406 VGND.n5404 0.120292
R24893 VGND.n5411 VGND.n5409 0.120292
R24894 VGND.n5413 VGND.n5411 0.120292
R24895 VGND.n5414 VGND.n5413 0.120292
R24896 VGND.n5423 VGND.n5421 0.120292
R24897 VGND.n5424 VGND.n5423 0.120292
R24898 VGND.n5425 VGND.n5424 0.120292
R24899 VGND.n5426 VGND.n5425 0.120292
R24900 VGND.n5432 VGND.n5430 0.120292
R24901 VGND.n5434 VGND.n5432 0.120292
R24902 VGND.n5437 VGND.n5434 0.120292
R24903 VGND.n5438 VGND.n5437 0.120292
R24904 VGND.n5439 VGND.n5438 0.120292
R24905 VGND.n5440 VGND.n5439 0.120292
R24906 VGND.n5448 VGND.n5447 0.120292
R24907 VGND.n5284 VGND.n5283 0.120292
R24908 VGND.n5283 VGND.n5281 0.120292
R24909 VGND.n5281 VGND.n5279 0.120292
R24910 VGND.n5279 VGND.n5277 0.120292
R24911 VGND.n5277 VGND.n5275 0.120292
R24912 VGND.n5275 VGND.n5273 0.120292
R24913 VGND.n5273 VGND.n5271 0.120292
R24914 VGND.n5271 VGND.n5268 0.120292
R24915 VGND.n5268 VGND.n5266 0.120292
R24916 VGND.n5266 VGND.n5264 0.120292
R24917 VGND.n5264 VGND.n5262 0.120292
R24918 VGND.n5258 VGND.n5227 0.120292
R24919 VGND.n5252 VGND.n5251 0.120292
R24920 VGND.n5251 VGND.n5250 0.120292
R24921 VGND.n5250 VGND.n5249 0.120292
R24922 VGND.n5249 VGND.n5246 0.120292
R24923 VGND.n5246 VGND.n5244 0.120292
R24924 VGND.n5244 VGND.n5242 0.120292
R24925 VGND.n5242 VGND.n5239 0.120292
R24926 VGND.n1806 VGND.n1805 0.120292
R24927 VGND.n1812 VGND.n1810 0.120292
R24928 VGND.n1813 VGND.n1812 0.120292
R24929 VGND.n1814 VGND.n1813 0.120292
R24930 VGND.n1820 VGND.n1817 0.120292
R24931 VGND.n1821 VGND.n1820 0.120292
R24932 VGND.n5968 VGND.n5966 0.120292
R24933 VGND.n5963 VGND.n5962 0.120292
R24934 VGND.n5962 VGND.n5961 0.120292
R24935 VGND.n5961 VGND.n5959 0.120292
R24936 VGND.n5959 VGND.n5957 0.120292
R24937 VGND.n5957 VGND.n5955 0.120292
R24938 VGND.n5955 VGND.n5953 0.120292
R24939 VGND.n5953 VGND.n5951 0.120292
R24940 VGND.n5951 VGND.n5948 0.120292
R24941 VGND.n5948 VGND.n5946 0.120292
R24942 VGND.n5946 VGND.n5944 0.120292
R24943 VGND.n5944 VGND.n5942 0.120292
R24944 VGND.n5938 VGND.n5937 0.120292
R24945 VGND.n5937 VGND.n5935 0.120292
R24946 VGND.n5935 VGND.n5934 0.120292
R24947 VGND.n5931 VGND.n5930 0.120292
R24948 VGND.n5928 VGND.n5925 0.120292
R24949 VGND.n5925 VGND.n5923 0.120292
R24950 VGND.n5923 VGND.n5921 0.120292
R24951 VGND.n5921 VGND.n5919 0.120292
R24952 VGND.n5919 VGND.n5917 0.120292
R24953 VGND.n5917 VGND.n5915 0.120292
R24954 VGND.n5915 VGND.n5913 0.120292
R24955 VGND.n5913 VGND.n5911 0.120292
R24956 VGND.n5911 VGND.n5908 0.120292
R24957 VGND.n5908 VGND.n5906 0.120292
R24958 VGND.n5906 VGND.n5905 0.120292
R24959 VGND.n5902 VGND.n5901 0.120292
R24960 VGND.n5901 VGND.n5899 0.120292
R24961 VGND.n5895 VGND.n5894 0.120292
R24962 VGND.n5501 VGND.n5500 0.120292
R24963 VGND.n5507 VGND.n5506 0.120292
R24964 VGND.n5509 VGND.n5507 0.120292
R24965 VGND.n5511 VGND.n5509 0.120292
R24966 VGND.n5513 VGND.n5511 0.120292
R24967 VGND.n5515 VGND.n5513 0.120292
R24968 VGND.n5517 VGND.n5515 0.120292
R24969 VGND.n5520 VGND.n5517 0.120292
R24970 VGND.n5522 VGND.n5520 0.120292
R24971 VGND.n5524 VGND.n5522 0.120292
R24972 VGND.n5526 VGND.n5524 0.120292
R24973 VGND.n5527 VGND.n5526 0.120292
R24974 VGND.n5532 VGND.n5530 0.120292
R24975 VGND.n5535 VGND.n5532 0.120292
R24976 VGND.n5537 VGND.n5535 0.120292
R24977 VGND.n5544 VGND.n5542 0.120292
R24978 VGND.n5546 VGND.n5544 0.120292
R24979 VGND.n5548 VGND.n5546 0.120292
R24980 VGND.n5551 VGND.n5548 0.120292
R24981 VGND.n5552 VGND.n5551 0.120292
R24982 VGND.n5553 VGND.n5552 0.120292
R24983 VGND.n5562 VGND.n5553 0.120292
R24984 VGND.n5568 VGND.n5566 0.120292
R24985 VGND.n5569 VGND.n5568 0.120292
R24986 VGND.n5570 VGND.n5569 0.120292
R24987 VGND.n5575 VGND.n5573 0.120292
R24988 VGND.n5578 VGND.n5575 0.120292
R24989 VGND.n5580 VGND.n5578 0.120292
R24990 VGND.n5583 VGND.n5580 0.120292
R24991 VGND.n5584 VGND.n5583 0.120292
R24992 VGND.n5649 VGND.n5647 0.120292
R24993 VGND.n5652 VGND.n5649 0.120292
R24994 VGND.n5657 VGND.n5652 0.120292
R24995 VGND.n5660 VGND.n5657 0.120292
R24996 VGND.n5661 VGND.n5660 0.120292
R24997 VGND.n5666 VGND.n5664 0.120292
R24998 VGND.n5669 VGND.n5666 0.120292
R24999 VGND.n5671 VGND.n5669 0.120292
R25000 VGND.n5674 VGND.n5671 0.120292
R25001 VGND.n5676 VGND.n5674 0.120292
R25002 VGND.n5682 VGND.n5681 0.120292
R25003 VGND.n5684 VGND.n5682 0.120292
R25004 VGND.n5686 VGND.n5684 0.120292
R25005 VGND.n5689 VGND.n5686 0.120292
R25006 VGND.n5694 VGND.n5689 0.120292
R25007 VGND.n5697 VGND.n5694 0.120292
R25008 VGND.n5700 VGND.n5697 0.120292
R25009 VGND.n5705 VGND.n5703 0.120292
R25010 VGND.n5707 VGND.n5705 0.120292
R25011 VGND.n5709 VGND.n5707 0.120292
R25012 VGND.n5711 VGND.n5709 0.120292
R25013 VGND.n5713 VGND.n5711 0.120292
R25014 VGND.n5715 VGND.n5713 0.120292
R25015 VGND.n5717 VGND.n5715 0.120292
R25016 VGND.n5720 VGND.n5717 0.120292
R25017 VGND.n5722 VGND.n5720 0.120292
R25018 VGND.n5723 VGND.n5722 0.120292
R25019 VGND.n5724 VGND.n5723 0.120292
R25020 VGND.n5729 VGND.n5727 0.120292
R25021 VGND.n5732 VGND.n5729 0.120292
R25022 VGND.n5733 VGND.n5732 0.120292
R25023 VGND.n5740 VGND.n5737 0.120292
R25024 VGND.n5185 VGND.n5183 0.120292
R25025 VGND.n5183 VGND.n5181 0.120292
R25026 VGND.n5181 VGND.n5179 0.120292
R25027 VGND.n5179 VGND.n5177 0.120292
R25028 VGND.n5177 VGND.n5175 0.120292
R25029 VGND.n5175 VGND.n5173 0.120292
R25030 VGND.n5173 VGND.n5170 0.120292
R25031 VGND.n5170 VGND.n5168 0.120292
R25032 VGND.n5168 VGND.n5166 0.120292
R25033 VGND.n5166 VGND.n5164 0.120292
R25034 VGND.n5160 VGND.n5159 0.120292
R25035 VGND.n5159 VGND.n5157 0.120292
R25036 VGND.n5156 VGND.n5152 0.120292
R25037 VGND.n5152 VGND.n5151 0.120292
R25038 VGND.n5144 VGND.n5143 0.120292
R25039 VGND.n5143 VGND.n5142 0.120292
R25040 VGND.n5139 VGND.n5138 0.120292
R25041 VGND.n5138 VGND.n5137 0.120292
R25042 VGND.n3492 VGND.n3490 0.120292
R25043 VGND.n3496 VGND.n3492 0.120292
R25044 VGND.n3498 VGND.n3496 0.120292
R25045 VGND.n3502 VGND.n3498 0.120292
R25046 VGND.n3503 VGND.n3502 0.120292
R25047 VGND.n9201 VGND.n9197 0.120292
R25048 VGND.n9197 VGND.n9195 0.120292
R25049 VGND.n9195 VGND.n9193 0.120292
R25050 VGND.n9193 VGND.n9191 0.120292
R25051 VGND.n9191 VGND.n9188 0.120292
R25052 VGND.n9188 VGND.n9187 0.120292
R25053 VGND.n9187 VGND.n9186 0.120292
R25054 VGND.n2187 VGND.n2186 0.120292
R25055 VGND.n2188 VGND.n2187 0.120292
R25056 VGND.n2197 VGND.n2196 0.120292
R25057 VGND.n2198 VGND.n2197 0.120292
R25058 VGND.n2199 VGND.n2198 0.120292
R25059 VGND.n2205 VGND.n2203 0.120292
R25060 VGND.n2208 VGND.n2205 0.120292
R25061 VGND.n2209 VGND.n2208 0.120292
R25062 VGND.n2210 VGND.n2209 0.120292
R25063 VGND.n2211 VGND.n2210 0.120292
R25064 VGND.n2217 VGND.n2215 0.120292
R25065 VGND.n2220 VGND.n2217 0.120292
R25066 VGND.n2221 VGND.n2220 0.120292
R25067 VGND.n2222 VGND.n2221 0.120292
R25068 VGND.n2223 VGND.n2222 0.120292
R25069 VGND.n2232 VGND.n2229 0.120292
R25070 VGND.n2620 VGND.n2284 0.120292
R25071 VGND.n2615 VGND.n2614 0.120292
R25072 VGND.n2614 VGND.n2613 0.120292
R25073 VGND.n2613 VGND.n2612 0.120292
R25074 VGND.n2612 VGND.n2610 0.120292
R25075 VGND.n2610 VGND.n2608 0.120292
R25076 VGND.n2608 VGND.n2605 0.120292
R25077 VGND.n2605 VGND.n2603 0.120292
R25078 VGND.n2603 VGND.n2600 0.120292
R25079 VGND.n2600 VGND.n2598 0.120292
R25080 VGND.n2590 VGND.n2589 0.120292
R25081 VGND.n2589 VGND.n2588 0.120292
R25082 VGND.n2583 VGND.n2582 0.120292
R25083 VGND.n2582 VGND.n2581 0.120292
R25084 VGND.n2581 VGND.n2580 0.120292
R25085 VGND.n2580 VGND.n2578 0.120292
R25086 VGND.n2573 VGND.n2572 0.120292
R25087 VGND.n2572 VGND 0.120292
R25088 VGND.n2570 VGND.n2567 0.120292
R25089 VGND.n2567 VGND.n2563 0.120292
R25090 VGND.n2563 VGND.n2562 0.120292
R25091 VGND.n2559 VGND.n2558 0.120292
R25092 VGND.n2558 VGND.n2554 0.120292
R25093 VGND.n2554 VGND.n2550 0.120292
R25094 VGND.n2550 VGND.n2548 0.120292
R25095 VGND.n2548 VGND.n2547 0.120292
R25096 VGND.n2477 VGND.n2340 0.120292
R25097 VGND.n2471 VGND.n2470 0.120292
R25098 VGND.n2470 VGND.n2468 0.120292
R25099 VGND.n2468 VGND.n2462 0.120292
R25100 VGND.n2462 VGND.n2460 0.120292
R25101 VGND.n2451 VGND.n2450 0.120292
R25102 VGND.n2450 VGND.n2448 0.120292
R25103 VGND.n2448 VGND.n2447 0.120292
R25104 VGND.n2443 VGND.n2442 0.120292
R25105 VGND.n2442 VGND.n2440 0.120292
R25106 VGND.n2440 VGND.n2438 0.120292
R25107 VGND.n2438 VGND.n2436 0.120292
R25108 VGND.n2436 VGND.n2432 0.120292
R25109 VGND.n2432 VGND.n2430 0.120292
R25110 VGND.n2430 VGND.n2428 0.120292
R25111 VGND.n2428 VGND.n2426 0.120292
R25112 VGND.n2426 VGND.n2423 0.120292
R25113 VGND.n2423 VGND.n2421 0.120292
R25114 VGND.n2421 VGND.n2420 0.120292
R25115 VGND.n2417 VGND.n2416 0.120292
R25116 VGND.n2416 VGND.n2415 0.120292
R25117 VGND.n2410 VGND.n2409 0.120292
R25118 VGND.n2408 VGND.n2403 0.120292
R25119 VGND.n9162 VGND.n9161 0.120292
R25120 VGND.n9161 VGND.n9160 0.120292
R25121 VGND.n9160 VGND.n9155 0.120292
R25122 VGND.n9155 VGND.n9152 0.120292
R25123 VGND.n9147 VGND.n9146 0.120292
R25124 VGND.n9146 VGND.n9144 0.120292
R25125 VGND.n9139 VGND.n9138 0.120292
R25126 VGND.n9138 VGND.n9136 0.120292
R25127 VGND.n9136 VGND.n9135 0.120292
R25128 VGND.n9135 VGND.n9133 0.120292
R25129 VGND.n9128 VGND.n9127 0.120292
R25130 VGND.n9127 VGND.n9126 0.120292
R25131 VGND.n9125 VGND.n9123 0.120292
R25132 VGND VGND.n445 0.12003
R25133 VGND.n2787 VGND.n2782 0.116385
R25134 VGND.n8649 VGND.n8648 0.116385
R25135 VGND.n1295 VGND.n1294 0.116385
R25136 VGND.n5647 VGND.n5645 0.116385
R25137 VGND.n4986 VGND.n4983 0.112781
R25138 VGND.n4795 VGND.n4793 0.111177
R25139 VGND.n4125 VGND.n4123 0.111177
R25140 VGND.n3696 VGND.n3695 0.111177
R25141 VGND.n6147 VGND.n6145 0.111177
R25142 VGND.n1741 VGND.n1738 0.111177
R25143 VGND.n1827 VGND.n1825 0.111177
R25144 VGND.n6577 VGND.n6575 0.106288
R25145 VGND.n4955 VGND.n4954 0.106288
R25146 VGND.n4300 VGND.n4298 0.106288
R25147 VGND.n3385 VGND.n3382 0.106288
R25148 VGND.n8863 VGND.n8860 0.106288
R25149 VGND.n3920 VGND.n3919 0.106288
R25150 VGND.n7635 VGND.n7634 0.106288
R25151 VGND.n7343 VGND.n7341 0.106288
R25152 VGND.n2241 VGND.n2232 0.106288
R25153 VGND.n5894 VGND.n5892 0.106288
R25154 VGND.n4867 VGND.n4864 0.105063
R25155 VGND.n4711 VGND.n4695 0.105063
R25156 VGND.n3578 VGND.n3451 0.105063
R25157 VGND.n3843 VGND.n3842 0.105063
R25158 VGND.n1969 VGND.n1957 0.105063
R25159 VGND.n7563 VGND.n7561 0.105063
R25160 VGND.n5969 VGND.n5968 0.104289
R25161 VGND.n4770 VGND 0.104136
R25162 VGND.n4102 VGND 0.104136
R25163 VGND.n2049 VGND 0.104136
R25164 VGND.n3671 VGND 0.104136
R25165 VGND.n3782 VGND 0.104136
R25166 VGND.n1887 VGND 0.104136
R25167 VGND.n695 VGND 0.104136
R25168 VGND.n7460 VGND 0.104136
R25169 VGND.n6118 VGND 0.104136
R25170 VGND.n1712 VGND 0.104136
R25171 VGND.n3486 VGND 0.104136
R25172 VGND.n2633 VGND.n2632 0.103019
R25173 VGND.n9092 VGND.n44 0.103019
R25174 VGND.n9089 VGND.n9088 0.103019
R25175 VGND.n3539 VGND.n3538 0.103019
R25176 VGND.n5056 VGND 0.0994583
R25177 VGND VGND.n7167 0.0994583
R25178 VGND.n701 VGND 0.0994583
R25179 VGND.n4772 VGND 0.0981562
R25180 VGND.n4894 VGND 0.0981562
R25181 VGND VGND.n4078 0.0981562
R25182 VGND VGND.n4077 0.0981562
R25183 VGND.n5083 VGND 0.0981562
R25184 VGND VGND.n4021 0.0981562
R25185 VGND.n7179 VGND 0.0981562
R25186 VGND VGND.n7136 0.0981562
R25187 VGND.n7041 VGND 0.0981562
R25188 VGND.n4108 VGND 0.0981562
R25189 VGND VGND.n4683 0.0981562
R25190 VGND.n4276 VGND 0.0981562
R25191 VGND VGND.n4217 0.0981562
R25192 VGND.n4462 VGND 0.0981562
R25193 VGND.n4550 VGND 0.0981562
R25194 VGND VGND.n1448 0.0981562
R25195 VGND VGND.n1430 0.0981562
R25196 VGND.n2070 VGND 0.0981562
R25197 VGND.n3426 VGND 0.0981562
R25198 VGND VGND.n3423 0.0981562
R25199 VGND.n3398 VGND 0.0981562
R25200 VGND.n3392 VGND 0.0981562
R25201 VGND.n2651 VGND 0.0981562
R25202 VGND.n3287 VGND 0.0981562
R25203 VGND VGND.n3280 0.0981562
R25204 VGND.n2792 VGND 0.0981562
R25205 VGND VGND.n2915 0.0981562
R25206 VGND.n3652 VGND 0.0981562
R25207 VGND.n8906 VGND 0.0981562
R25208 VGND VGND.n8904 0.0981562
R25209 VGND VGND.n8878 0.0981562
R25210 VGND.n3045 VGND 0.0981562
R25211 VGND.n3074 VGND 0.0981562
R25212 VGND.n3079 VGND 0.0981562
R25213 VGND.n3106 VGND 0.0981562
R25214 VGND VGND.n2687 0.0981562
R25215 VGND.n3788 VGND 0.0981562
R25216 VGND.n3800 VGND 0.0981562
R25217 VGND.n3876 VGND 0.0981562
R25218 VGND.n3920 VGND 0.0981562
R25219 VGND.n8770 VGND 0.0981562
R25220 VGND VGND.n8754 0.0981562
R25221 VGND.n8719 VGND 0.0981562
R25222 VGND.n8642 VGND 0.0981562
R25223 VGND VGND.n8635 0.0981562
R25224 VGND.n8578 VGND 0.0981562
R25225 VGND VGND.n8475 0.0981562
R25226 VGND.n1893 VGND 0.0981562
R25227 VGND VGND.n1878 0.0981562
R25228 VGND.n1907 VGND 0.0981562
R25229 VGND.n7833 VGND 0.0981562
R25230 VGND.n7838 VGND 0.0981562
R25231 VGND VGND.n8023 0.0981562
R25232 VGND VGND.n8388 0.0981562
R25233 VGND.n8369 VGND 0.0981562
R25234 VGND VGND.n8367 0.0981562
R25235 VGND.n7588 VGND 0.0981562
R25236 VGND.n7664 VGND 0.0981562
R25237 VGND.n7649 VGND 0.0981562
R25238 VGND VGND.n618 0.0981562
R25239 VGND.n381 VGND 0.0981562
R25240 VGND VGND.n355 0.0981562
R25241 VGND.n7481 VGND 0.0981562
R25242 VGND VGND.n7424 0.0981562
R25243 VGND VGND.n7385 0.0981562
R25244 VGND.n7354 VGND 0.0981562
R25245 VGND.n1025 VGND 0.0981562
R25246 VGND.n1289 VGND 0.0981562
R25247 VGND.n1283 VGND 0.0981562
R25248 VGND.n1251 VGND 0.0981562
R25249 VGND VGND.n937 0.0981562
R25250 VGND.n6242 VGND 0.0981562
R25251 VGND VGND.n6304 0.0981562
R25252 VGND VGND.n6393 0.0981562
R25253 VGND.n6894 VGND 0.0981562
R25254 VGND.n1497 VGND 0.0981562
R25255 VGND.n6595 VGND 0.0981562
R25256 VGND.n6590 VGND 0.0981562
R25257 VGND.n6638 VGND 0.0981562
R25258 VGND.n6680 VGND 0.0981562
R25259 VGND.n6697 VGND 0.0981562
R25260 VGND.n5379 VGND 0.0981562
R25261 VGND.n5401 VGND 0.0981562
R25262 VGND.n5446 VGND 0.0981562
R25263 VGND.n5447 VGND 0.0981562
R25264 VGND.n5259 VGND 0.0981562
R25265 VGND VGND.n5258 0.0981562
R25266 VGND.n1805 VGND 0.0981562
R25267 VGND.n5939 VGND 0.0981562
R25268 VGND.n5902 VGND 0.0981562
R25269 VGND.n5895 VGND 0.0981562
R25270 VGND.n5530 VGND 0.0981562
R25271 VGND.n5727 VGND 0.0981562
R25272 VGND.n5161 VGND 0.0981562
R25273 VGND VGND.n5160 0.0981562
R25274 VGND.n3507 VGND 0.0981562
R25275 VGND.n16 VGND 0.0981562
R25276 VGND.n2191 VGND 0.0981562
R25277 VGND.n2215 VGND 0.0981562
R25278 VGND.n2224 VGND 0.0981562
R25279 VGND.n2229 VGND 0.0981562
R25280 VGND VGND.n2593 0.0981562
R25281 VGND.n2590 VGND 0.0981562
R25282 VGND.n2573 VGND 0.0981562
R25283 VGND.n2417 VGND 0.0981562
R25284 VGND.n2411 VGND 0.0981562
R25285 VGND VGND.n9147 0.0981562
R25286 VGND.n9139 VGND 0.0981562
R25287 VGND.n9128 VGND 0.0981562
R25288 VGND.n7189 VGND 0.0968542
R25289 VGND.n7156 VGND 0.0968542
R25290 VGND.n4395 VGND 0.0968542
R25291 VGND.n4530 VGND 0.0968542
R25292 VGND VGND.n4633 0.0968542
R25293 VGND VGND.n2929 0.0968542
R25294 VGND.n3054 VGND 0.0968542
R25295 VGND VGND.n8482 0.0968542
R25296 VGND VGND.n8061 0.0968542
R25297 VGND.n8051 VGND 0.0968542
R25298 VGND VGND.n8377 0.0968542
R25299 VGND VGND.n1288 0.0968542
R25300 VGND VGND.n1258 0.0968542
R25301 VGND VGND.n1220 0.0968542
R25302 VGND VGND.n943 0.0968542
R25303 VGND.n6834 VGND 0.0968542
R25304 VGND VGND.n2481 0.0968542
R25305 VGND.n4114 VGND 0.0955521
R25306 VGND VGND.n8718 0.0955521
R25307 VGND VGND.n7923 0.0955521
R25308 VGND VGND.n8028 0.0955521
R25309 VGND VGND.n380 0.0955521
R25310 VGND.n4016 VGND.n4012 0.0946561
R25311 VGND.n6727 VGND.n6719 0.0946561
R25312 VGND.n5606 VGND.n5588 0.0946561
R25313 VGND.n3245 VGND.n3244 0.0946561
R25314 VGND.n9014 VGND.n9007 0.0946561
R25315 VGND.n8718 VGND.n8717 0.0946561
R25316 VGND.n8223 VGND.n8217 0.0946561
R25317 VGND.n1134 VGND.n1125 0.0946561
R25318 VGND.n6793 VGND.n1595 0.0946561
R25319 VGND.n7327 VGND.n829 0.0942472
R25320 VGND.n7298 VGND.n7297 0.0942472
R25321 VGND.n7294 VGND.n7291 0.0942472
R25322 VGND.n2184 VGND.n2183 0.0900105
R25323 VGND.n4546 VGND.n4545 0.0900105
R25324 VGND.n3052 VGND.n3051 0.0900105
R25325 VGND.n8160 VGND.n449 0.0900105
R25326 VGND.n8308 VGND.n444 0.0900105
R25327 VGND.n1291 VGND.n1290 0.0900105
R25328 VGND.n4590 VGND.n4589 0.0881712
R25329 VGND.n2818 VGND.n2817 0.0881712
R25330 VGND.n3961 VGND.n3959 0.0881712
R25331 VGND.n499 VGND.n498 0.0881712
R25332 VGND.n8220 VGND.n8219 0.0881712
R25333 VGND.n1091 VGND.n1090 0.0881712
R25334 VGND.n792 VGND.n791 0.0881712
R25335 VGND.n6250 VGND.n6249 0.0881712
R25336 VGND VGND.n6277 0.0841522
R25337 VGND.n3281 VGND 0.0826382
R25338 VGND.n3424 VGND 0.0826382
R25339 VGND.n3664 VGND 0.0826382
R25340 VGND.n8879 VGND 0.0826382
R25341 VGND.n8737 VGND 0.0826382
R25342 VGND VGND.n6237 0.0826382
R25343 VGND.n6673 VGND 0.0826382
R25344 VGND VGND.n6702 0.0826382
R25345 VGND.n6703 VGND 0.0826382
R25346 VGND.n5373 VGND 0.0826382
R25347 VGND.n2594 VGND 0.0826382
R25348 VGND.n9203 VGND 0.0826382
R25349 VGND VGND.n9100 0.0826382
R25350 VGND.n445 VGND 0.0822696
R25351 VGND.n1461 VGND.n1452 0.0772651
R25352 VGND.n2978 VGND.n2966 0.0772651
R25353 VGND.n3185 VGND.n2736 0.0772651
R25354 VGND.n8416 VGND.n8404 0.0772651
R25355 VGND.n6961 VGND.n1536 0.0772651
R25356 VGND.n987 VGND.n977 0.0764916
R25357 VGND.n5795 VGND.n5185 0.0764916
R25358 VGND.n4514 VGND.n4513 0.0711194
R25359 VGND.n8194 VGND.n8193 0.0711194
R25360 VGND.n1317 VGND.n1316 0.0711194
R25361 VGND.n2513 VGND.n2512 0.0711194
R25362 VGND.n7222 VGND.n7221 0.0709266
R25363 VGND.n9045 VGND.n9044 0.0709266
R25364 VGND.n8706 VGND.n8705 0.0709266
R25365 VGND.n8091 VGND.n8090 0.0709266
R25366 VGND.n6819 VGND.n6818 0.0709266
R25367 VGND.n5368 VGND.n5367 0.0709266
R25368 VGND.n5639 VGND.n5638 0.0709266
R25369 VGND.n5044 VGND.n5043 0.0700652
R25370 VGND.n2491 VGND.n2490 0.0685851
R25371 VGND.n1740 VGND.n1739 0.0685851
R25372 VGND.n4852 VGND.n4851 0.0685851
R25373 VGND.n1421 VGND.n1420 0.0685851
R25374 VGND.n2870 VGND.n2869 0.0685851
R25375 VGND.n8387 VGND.n8386 0.0685851
R25376 VGND.n1892 VGND.n1891 0.0685851
R25377 VGND.n1882 VGND.n1881 0.0685851
R25378 VGND.n7436 VGND.n7435 0.0685851
R25379 VGND.n7113 VGND.n7110 0.0670478
R25380 VGND.n4594 VGND.n4587 0.0670478
R25381 VGND.n3173 VGND.n3132 0.0670478
R25382 VGND.n8572 VGND.n8571 0.0670478
R25383 VGND.n7989 VGND.n7987 0.0670478
R25384 VGND.n1205 VGND.n1203 0.0670478
R25385 VGND.n6931 VGND.n6922 0.0670478
R25386 VGND.n5456 VGND.n5195 0.0670478
R25387 VGND.n5752 VGND.n5740 0.0670478
R25388 VGND.n2403 VGND.n2399 0.0670478
R25389 VGND.n4771 VGND 0.0603958
R25390 VGND.n4776 VGND 0.0603958
R25391 VGND VGND.n4785 0.0603958
R25392 VGND.n4786 VGND 0.0603958
R25393 VGND.n4789 VGND 0.0603958
R25394 VGND.n4871 VGND 0.0603958
R25395 VGND.n4889 VGND 0.0603958
R25396 VGND VGND.n4088 0.0603958
R25397 VGND.n4903 VGND 0.0603958
R25398 VGND.n4905 VGND 0.0603958
R25399 VGND.n4913 VGND 0.0603958
R25400 VGND.n4921 VGND 0.0603958
R25401 VGND VGND.n4075 0.0603958
R25402 VGND.n4075 VGND 0.0603958
R25403 VGND.n4952 VGND 0.0603958
R25404 VGND.n5015 VGND 0.0603958
R25405 VGND.n5021 VGND 0.0603958
R25406 VGND.n5024 VGND 0.0603958
R25407 VGND.n5028 VGND 0.0603958
R25408 VGND.n5042 VGND 0.0603958
R25409 VGND.n5050 VGND 0.0603958
R25410 VGND.n5052 VGND 0.0603958
R25411 VGND.n5064 VGND 0.0603958
R25412 VGND.n5069 VGND 0.0603958
R25413 VGND.n5081 VGND 0.0603958
R25414 VGND.n5084 VGND 0.0603958
R25415 VGND.n5085 VGND 0.0603958
R25416 VGND VGND.n4033 0.0603958
R25417 VGND VGND.n4032 0.0603958
R25418 VGND VGND.n4029 0.0603958
R25419 VGND VGND.n4028 0.0603958
R25420 VGND.n4024 VGND 0.0603958
R25421 VGND.n4024 VGND 0.0603958
R25422 VGND VGND.n4023 0.0603958
R25423 VGND VGND.n4022 0.0603958
R25424 VGND.n4017 VGND 0.0603958
R25425 VGND.n7193 VGND 0.0603958
R25426 VGND VGND.n7192 0.0603958
R25427 VGND.n7188 VGND 0.0603958
R25428 VGND.n7185 VGND 0.0603958
R25429 VGND VGND.n7183 0.0603958
R25430 VGND.n7170 VGND 0.0603958
R25431 VGND VGND.n7169 0.0603958
R25432 VGND VGND.n7168 0.0603958
R25433 VGND VGND.n7160 0.0603958
R25434 VGND.n7153 VGND 0.0603958
R25435 VGND VGND.n7152 0.0603958
R25436 VGND.n7145 VGND 0.0603958
R25437 VGND.n7140 VGND 0.0603958
R25438 VGND.n7137 VGND 0.0603958
R25439 VGND.n7120 VGND 0.0603958
R25440 VGND.n7120 VGND 0.0603958
R25441 VGND VGND.n7119 0.0603958
R25442 VGND.n7116 VGND 0.0603958
R25443 VGND.n7059 VGND 0.0603958
R25444 VGND.n4103 VGND 0.0603958
R25445 VGND.n4104 VGND 0.0603958
R25446 VGND.n4109 VGND 0.0603958
R25447 VGND VGND.n4109 0.0603958
R25448 VGND.n4110 VGND 0.0603958
R25449 VGND.n4115 VGND 0.0603958
R25450 VGND.n4119 VGND 0.0603958
R25451 VGND.n4695 VGND 0.0603958
R25452 VGND.n4692 VGND 0.0603958
R25453 VGND.n4684 VGND 0.0603958
R25454 VGND.n4671 VGND 0.0603958
R25455 VGND.n4664 VGND 0.0603958
R25456 VGND VGND.n4663 0.0603958
R25457 VGND.n4242 VGND 0.0603958
R25458 VGND.n4250 VGND 0.0603958
R25459 VGND.n4286 VGND 0.0603958
R25460 VGND.n4296 VGND 0.0603958
R25461 VGND.n4383 VGND 0.0603958
R25462 VGND.n4389 VGND 0.0603958
R25463 VGND.n4390 VGND 0.0603958
R25464 VGND VGND.n4418 0.0603958
R25465 VGND.n4419 VGND 0.0603958
R25466 VGND.n4426 VGND 0.0603958
R25467 VGND.n4437 VGND 0.0603958
R25468 VGND.n4438 VGND 0.0603958
R25469 VGND.n4443 VGND 0.0603958
R25470 VGND.n4444 VGND 0.0603958
R25471 VGND VGND.n4454 0.0603958
R25472 VGND.n4455 VGND 0.0603958
R25473 VGND.n4456 VGND 0.0603958
R25474 VGND.n4471 VGND 0.0603958
R25475 VGND.n4474 VGND 0.0603958
R25476 VGND VGND.n4474 0.0603958
R25477 VGND.n4475 VGND 0.0603958
R25478 VGND.n4523 VGND 0.0603958
R25479 VGND.n4524 VGND 0.0603958
R25480 VGND VGND.n4534 0.0603958
R25481 VGND.n4536 VGND 0.0603958
R25482 VGND.n4542 VGND 0.0603958
R25483 VGND.n4549 VGND 0.0603958
R25484 VGND.n4655 VGND 0.0603958
R25485 VGND.n4650 VGND 0.0603958
R25486 VGND VGND.n4649 0.0603958
R25487 VGND.n4635 VGND 0.0603958
R25488 VGND VGND.n4634 0.0603958
R25489 VGND.n4566 VGND 0.0603958
R25490 VGND VGND.n4566 0.0603958
R25491 VGND.n4567 VGND 0.0603958
R25492 VGND.n4611 VGND 0.0603958
R25493 VGND.n1449 VGND 0.0603958
R25494 VGND.n1447 VGND 0.0603958
R25495 VGND.n1443 VGND 0.0603958
R25496 VGND.n1434 VGND 0.0603958
R25497 VGND VGND.n1431 0.0603958
R25498 VGND.n1429 VGND 0.0603958
R25499 VGND.n1426 VGND 0.0603958
R25500 VGND VGND.n1425 0.0603958
R25501 VGND VGND.n1424 0.0603958
R25502 VGND.n2055 VGND 0.0603958
R25503 VGND.n2062 VGND 0.0603958
R25504 VGND.n2069 VGND 0.0603958
R25505 VGND.n2071 VGND 0.0603958
R25506 VGND VGND.n3445 0.0603958
R25507 VGND VGND.n3425 0.0603958
R25508 VGND.n3414 VGND 0.0603958
R25509 VGND VGND.n3324 0.0603958
R25510 VGND VGND.n3312 0.0603958
R25511 VGND VGND.n3279 0.0603958
R25512 VGND VGND.n3266 0.0603958
R25513 VGND.n3210 VGND 0.0603958
R25514 VGND.n3262 VGND 0.0603958
R25515 VGND VGND.n3261 0.0603958
R25516 VGND.n3246 VGND 0.0603958
R25517 VGND VGND.n2757 0.0603958
R25518 VGND VGND.n2756 0.0603958
R25519 VGND.n2803 VGND 0.0603958
R25520 VGND.n2812 VGND 0.0603958
R25521 VGND.n2814 VGND 0.0603958
R25522 VGND.n2821 VGND 0.0603958
R25523 VGND.n2831 VGND 0.0603958
R25524 VGND.n2842 VGND 0.0603958
R25525 VGND.n2847 VGND 0.0603958
R25526 VGND.n2851 VGND 0.0603958
R25527 VGND.n2858 VGND 0.0603958
R25528 VGND VGND.n2747 0.0603958
R25529 VGND.n2871 VGND 0.0603958
R25530 VGND VGND.n2965 0.0603958
R25531 VGND.n2961 VGND 0.0603958
R25532 VGND.n2941 VGND 0.0603958
R25533 VGND.n2931 VGND 0.0603958
R25534 VGND VGND.n2930 0.0603958
R25535 VGND.n2927 VGND 0.0603958
R25536 VGND VGND.n2926 0.0603958
R25537 VGND.n2916 VGND 0.0603958
R25538 VGND VGND.n2914 0.0603958
R25539 VGND.n3677 VGND 0.0603958
R25540 VGND.n3683 VGND 0.0603958
R25541 VGND.n3688 VGND 0.0603958
R25542 VGND.n3692 VGND 0.0603958
R25543 VGND VGND.n3663 0.0603958
R25544 VGND VGND.n8899 0.0603958
R25545 VGND.n88 VGND 0.0603958
R25546 VGND VGND.n8885 0.0603958
R25547 VGND.n8870 VGND 0.0603958
R25548 VGND.n8921 VGND 0.0603958
R25549 VGND.n8924 VGND 0.0603958
R25550 VGND.n8935 VGND 0.0603958
R25551 VGND.n8941 VGND 0.0603958
R25552 VGND.n8955 VGND 0.0603958
R25553 VGND.n8961 VGND 0.0603958
R25554 VGND.n8971 VGND 0.0603958
R25555 VGND.n8978 VGND 0.0603958
R25556 VGND.n8984 VGND 0.0603958
R25557 VGND.n3041 VGND 0.0603958
R25558 VGND VGND.n3036 0.0603958
R25559 VGND.n3048 VGND 0.0603958
R25560 VGND.n3048 VGND 0.0603958
R25561 VGND.n3053 VGND 0.0603958
R25562 VGND.n3055 VGND 0.0603958
R25563 VGND.n3059 VGND 0.0603958
R25564 VGND.n3068 VGND 0.0603958
R25565 VGND.n3073 VGND 0.0603958
R25566 VGND.n3083 VGND 0.0603958
R25567 VGND.n3086 VGND 0.0603958
R25568 VGND.n2727 VGND 0.0603958
R25569 VGND VGND.n2726 0.0603958
R25570 VGND.n2715 VGND 0.0603958
R25571 VGND.n2697 VGND 0.0603958
R25572 VGND VGND.n2696 0.0603958
R25573 VGND VGND.n2688 0.0603958
R25574 VGND.n3783 VGND 0.0603958
R25575 VGND.n3784 VGND 0.0603958
R25576 VGND.n3793 VGND 0.0603958
R25577 VGND.n3793 VGND 0.0603958
R25578 VGND.n3799 VGND 0.0603958
R25579 VGND VGND.n3843 0.0603958
R25580 VGND.n3844 VGND 0.0603958
R25581 VGND.n3850 VGND 0.0603958
R25582 VGND.n3856 VGND 0.0603958
R25583 VGND.n3877 VGND 0.0603958
R25584 VGND.n3976 VGND 0.0603958
R25585 VGND VGND.n3955 0.0603958
R25586 VGND.n3885 VGND 0.0603958
R25587 VGND.n3950 VGND 0.0603958
R25588 VGND.n3925 VGND 0.0603958
R25589 VGND VGND.n3924 0.0603958
R25590 VGND.n161 VGND 0.0603958
R25591 VGND.n8781 VGND 0.0603958
R25592 VGND VGND.n8780 0.0603958
R25593 VGND.n8777 VGND 0.0603958
R25594 VGND.n8767 VGND 0.0603958
R25595 VGND VGND.n8766 0.0603958
R25596 VGND.n8763 VGND 0.0603958
R25597 VGND VGND.n8755 0.0603958
R25598 VGND.n8752 VGND 0.0603958
R25599 VGND VGND.n8751 0.0603958
R25600 VGND.n8738 VGND 0.0603958
R25601 VGND VGND.n8736 0.0603958
R25602 VGND.n8733 VGND 0.0603958
R25603 VGND VGND.n8732 0.0603958
R25604 VGND.n8725 VGND 0.0603958
R25605 VGND.n8636 VGND 0.0603958
R25606 VGND.n8626 VGND 0.0603958
R25607 VGND.n8622 VGND 0.0603958
R25608 VGND VGND.n8621 0.0603958
R25609 VGND.n8614 VGND 0.0603958
R25610 VGND.n238 VGND 0.0603958
R25611 VGND VGND.n8594 0.0603958
R25612 VGND VGND.n8593 0.0603958
R25613 VGND.n8584 VGND 0.0603958
R25614 VGND VGND.n8582 0.0603958
R25615 VGND.n8572 VGND 0.0603958
R25616 VGND.n8501 VGND 0.0603958
R25617 VGND.n8491 VGND 0.0603958
R25618 VGND.n8483 VGND 0.0603958
R25619 VGND.n8481 VGND 0.0603958
R25620 VGND VGND.n8480 0.0603958
R25621 VGND.n8476 VGND 0.0603958
R25622 VGND.n1896 VGND 0.0603958
R25623 VGND.n1906 VGND 0.0603958
R25624 VGND.n1907 VGND 0.0603958
R25625 VGND.n1957 VGND 0.0603958
R25626 VGND VGND.n1956 0.0603958
R25627 VGND.n1953 VGND 0.0603958
R25628 VGND VGND.n1951 0.0603958
R25629 VGND VGND.n1950 0.0603958
R25630 VGND.n7809 VGND 0.0603958
R25631 VGND VGND.n7808 0.0603958
R25632 VGND.n7804 VGND 0.0603958
R25633 VGND.n7786 VGND 0.0603958
R25634 VGND.n7781 VGND 0.0603958
R25635 VGND VGND.n7780 0.0603958
R25636 VGND.n7765 VGND 0.0603958
R25637 VGND.n7820 VGND 0.0603958
R25638 VGND.n7827 VGND 0.0603958
R25639 VGND.n7834 VGND 0.0603958
R25640 VGND.n7847 VGND 0.0603958
R25641 VGND VGND.n7848 0.0603958
R25642 VGND.n7849 VGND 0.0603958
R25643 VGND.n7856 VGND 0.0603958
R25644 VGND.n7867 VGND 0.0603958
R25645 VGND.n7870 VGND 0.0603958
R25646 VGND.n7873 VGND 0.0603958
R25647 VGND.n7889 VGND 0.0603958
R25648 VGND.n7890 VGND 0.0603958
R25649 VGND.n7939 VGND 0.0603958
R25650 VGND.n7924 VGND 0.0603958
R25651 VGND.n8062 VGND 0.0603958
R25652 VGND VGND.n8055 0.0603958
R25653 VGND.n8048 VGND 0.0603958
R25654 VGND.n8045 VGND 0.0603958
R25655 VGND.n8044 VGND 0.0603958
R25656 VGND VGND.n8043 0.0603958
R25657 VGND.n8039 VGND 0.0603958
R25658 VGND VGND.n8038 0.0603958
R25659 VGND.n8029 VGND 0.0603958
R25660 VGND.n8027 VGND 0.0603958
R25661 VGND.n8024 VGND 0.0603958
R25662 VGND.n7998 VGND 0.0603958
R25663 VGND VGND.n7989 0.0603958
R25664 VGND.n8401 VGND 0.0603958
R25665 VGND VGND.n8393 0.0603958
R25666 VGND.n8390 VGND 0.0603958
R25667 VGND VGND.n8389 0.0603958
R25668 VGND VGND.n8378 0.0603958
R25669 VGND.n8375 VGND 0.0603958
R25670 VGND VGND.n8374 0.0603958
R25671 VGND VGND.n8373 0.0603958
R25672 VGND VGND.n8372 0.0603958
R25673 VGND VGND.n8368 0.0603958
R25674 VGND.n8359 VGND 0.0603958
R25675 VGND.n696 VGND 0.0603958
R25676 VGND.n700 VGND 0.0603958
R25677 VGND.n702 VGND 0.0603958
R25678 VGND.n702 VGND 0.0603958
R25679 VGND.n706 VGND 0.0603958
R25680 VGND.n7572 VGND 0.0603958
R25681 VGND.n7577 VGND 0.0603958
R25682 VGND.n7582 VGND 0.0603958
R25683 VGND.n7682 VGND 0.0603958
R25684 VGND VGND.n7681 0.0603958
R25685 VGND VGND.n7680 0.0603958
R25686 VGND VGND.n7668 0.0603958
R25687 VGND.n7636 VGND 0.0603958
R25688 VGND VGND.n7635 0.0603958
R25689 VGND.n678 VGND 0.0603958
R25690 VGND.n678 VGND 0.0603958
R25691 VGND VGND.n677 0.0603958
R25692 VGND VGND.n676 0.0603958
R25693 VGND.n662 VGND 0.0603958
R25694 VGND.n650 VGND 0.0603958
R25695 VGND VGND.n623 0.0603958
R25696 VGND VGND.n620 0.0603958
R25697 VGND.n8251 VGND 0.0603958
R25698 VGND VGND.n8250 0.0603958
R25699 VGND.n8248 VGND 0.0603958
R25700 VGND VGND.n8247 0.0603958
R25701 VGND.n8242 VGND 0.0603958
R25702 VGND.n8186 VGND 0.0603958
R25703 VGND.n8175 VGND 0.0603958
R25704 VGND VGND.n8173 0.0603958
R25705 VGND VGND.n450 0.0603958
R25706 VGND.n8260 VGND 0.0603958
R25707 VGND.n8261 VGND 0.0603958
R25708 VGND.n8269 VGND 0.0603958
R25709 VGND.n8278 VGND 0.0603958
R25710 VGND.n8283 VGND 0.0603958
R25711 VGND.n392 VGND 0.0603958
R25712 VGND.n379 VGND 0.0603958
R25713 VGND.n376 VGND 0.0603958
R25714 VGND.n356 VGND 0.0603958
R25715 VGND.n7466 VGND 0.0603958
R25716 VGND.n7472 VGND 0.0603958
R25717 VGND.n7478 VGND 0.0603958
R25718 VGND.n7482 VGND 0.0603958
R25719 VGND.n7425 VGND 0.0603958
R25720 VGND.n7411 VGND 0.0603958
R25721 VGND.n7411 VGND 0.0603958
R25722 VGND VGND.n7410 0.0603958
R25723 VGND.n7392 VGND 0.0603958
R25724 VGND VGND.n7391 0.0603958
R25725 VGND VGND.n7389 0.0603958
R25726 VGND VGND.n7350 0.0603958
R25727 VGND.n7344 VGND 0.0603958
R25728 VGND.n1020 VGND 0.0603958
R25729 VGND.n1028 VGND 0.0603958
R25730 VGND.n1033 VGND 0.0603958
R25731 VGND.n1037 VGND 0.0603958
R25732 VGND.n1051 VGND 0.0603958
R25733 VGND.n1071 VGND 0.0603958
R25734 VGND.n1077 VGND 0.0603958
R25735 VGND.n1093 VGND 0.0603958
R25736 VGND.n1099 VGND 0.0603958
R25737 VGND.n1100 VGND 0.0603958
R25738 VGND.n1105 VGND 0.0603958
R25739 VGND.n1114 VGND 0.0603958
R25740 VGND VGND.n1116 0.0603958
R25741 VGND.n1117 VGND 0.0603958
R25742 VGND.n1121 VGND 0.0603958
R25743 VGND.n1287 VGND 0.0603958
R25744 VGND VGND.n1286 0.0603958
R25745 VGND.n1274 VGND 0.0603958
R25746 VGND VGND.n1271 0.0603958
R25747 VGND VGND.n1270 0.0603958
R25748 VGND VGND.n1262 0.0603958
R25749 VGND.n1259 VGND 0.0603958
R25750 VGND.n1256 VGND 0.0603958
R25751 VGND VGND.n1255 0.0603958
R25752 VGND.n1240 VGND 0.0603958
R25753 VGND VGND.n1239 0.0603958
R25754 VGND.n1221 VGND 0.0603958
R25755 VGND.n1219 VGND 0.0603958
R25756 VGND VGND.n1218 0.0603958
R25757 VGND VGND.n1217 0.0603958
R25758 VGND.n974 VGND 0.0603958
R25759 VGND.n972 VGND 0.0603958
R25760 VGND.n969 VGND 0.0603958
R25761 VGND.n955 VGND 0.0603958
R25762 VGND VGND.n949 0.0603958
R25763 VGND.n944 VGND 0.0603958
R25764 VGND.n942 VGND 0.0603958
R25765 VGND VGND.n941 0.0603958
R25766 VGND.n938 VGND 0.0603958
R25767 VGND.n6122 VGND 0.0603958
R25768 VGND.n6138 VGND 0.0603958
R25769 VGND.n6220 VGND 0.0603958
R25770 VGND VGND.n6220 0.0603958
R25771 VGND.n6221 VGND 0.0603958
R25772 VGND.n6228 VGND 0.0603958
R25773 VGND.n6238 VGND 0.0603958
R25774 VGND VGND.n6243 0.0603958
R25775 VGND.n6244 VGND 0.0603958
R25776 VGND.n6253 VGND 0.0603958
R25777 VGND.n6255 VGND 0.0603958
R25778 VGND.n6334 VGND 0.0603958
R25779 VGND.n6328 VGND 0.0603958
R25780 VGND.n6290 VGND 0.0603958
R25781 VGND.n6284 VGND 0.0603958
R25782 VGND VGND.n6283 0.0603958
R25783 VGND.n6278 VGND 0.0603958
R25784 VGND.n6341 VGND 0.0603958
R25785 VGND.n6452 VGND 0.0603958
R25786 VGND.n6444 VGND 0.0603958
R25787 VGND VGND.n6394 0.0603958
R25788 VGND VGND.n6391 0.0603958
R25789 VGND.n6355 VGND 0.0603958
R25790 VGND.n6382 VGND 0.0603958
R25791 VGND.n6375 VGND 0.0603958
R25792 VGND.n6826 VGND 0.0603958
R25793 VGND VGND.n6854 0.0603958
R25794 VGND.n6856 VGND 0.0603958
R25795 VGND.n6859 VGND 0.0603958
R25796 VGND.n6865 VGND 0.0603958
R25797 VGND.n6876 VGND 0.0603958
R25798 VGND.n6896 VGND 0.0603958
R25799 VGND.n6899 VGND 0.0603958
R25800 VGND.n6912 VGND 0.0603958
R25801 VGND.n1532 VGND 0.0603958
R25802 VGND.n1523 VGND 0.0603958
R25803 VGND VGND.n1520 0.0603958
R25804 VGND.n1718 VGND 0.0603958
R25805 VGND.n1724 VGND 0.0603958
R25806 VGND.n1730 VGND 0.0603958
R25807 VGND.n1734 VGND 0.0603958
R25808 VGND.n6052 VGND 0.0603958
R25809 VGND.n6034 VGND 0.0603958
R25810 VGND VGND.n6033 0.0603958
R25811 VGND.n6021 VGND 0.0603958
R25812 VGND.n6627 VGND 0.0603958
R25813 VGND VGND.n6626 0.0603958
R25814 VGND VGND.n6622 0.0603958
R25815 VGND VGND.n6614 0.0603958
R25816 VGND.n6586 VGND 0.0603958
R25817 VGND.n6582 VGND 0.0603958
R25818 VGND.n6635 VGND 0.0603958
R25819 VGND.n6639 VGND 0.0603958
R25820 VGND.n6642 VGND 0.0603958
R25821 VGND.n6655 VGND 0.0603958
R25822 VGND.n6658 VGND 0.0603958
R25823 VGND.n6679 VGND 0.0603958
R25824 VGND.n6681 VGND 0.0603958
R25825 VGND.n6684 VGND 0.0603958
R25826 VGND.n6691 VGND 0.0603958
R25827 VGND.n6698 VGND 0.0603958
R25828 VGND.n6708 VGND 0.0603958
R25829 VGND.n5404 VGND 0.0603958
R25830 VGND.n5409 VGND 0.0603958
R25831 VGND.n5416 VGND 0.0603958
R25832 VGND.n5421 VGND 0.0603958
R25833 VGND.n5430 VGND 0.0603958
R25834 VGND.n5448 VGND 0.0603958
R25835 VGND VGND.n5195 0.0603958
R25836 VGND VGND.n5227 0.0603958
R25837 VGND.n5253 VGND 0.0603958
R25838 VGND VGND.n5252 0.0603958
R25839 VGND.n1806 VGND 0.0603958
R25840 VGND.n1810 VGND 0.0603958
R25841 VGND.n1817 VGND 0.0603958
R25842 VGND.n1822 VGND 0.0603958
R25843 VGND.n1825 VGND 0.0603958
R25844 VGND.n5963 VGND 0.0603958
R25845 VGND VGND.n5938 0.0603958
R25846 VGND.n5931 VGND 0.0603958
R25847 VGND VGND.n5928 0.0603958
R25848 VGND VGND.n5898 0.0603958
R25849 VGND.n5500 VGND 0.0603958
R25850 VGND.n5506 VGND 0.0603958
R25851 VGND.n5538 VGND 0.0603958
R25852 VGND.n5542 VGND 0.0603958
R25853 VGND.n5563 VGND 0.0603958
R25854 VGND.n5566 VGND 0.0603958
R25855 VGND.n5573 VGND 0.0603958
R25856 VGND.n5588 VGND 0.0603958
R25857 VGND.n5664 VGND 0.0603958
R25858 VGND.n5677 VGND 0.0603958
R25859 VGND.n5681 VGND 0.0603958
R25860 VGND.n5703 VGND 0.0603958
R25861 VGND.n5737 VGND 0.0603958
R25862 VGND.n5157 VGND 0.0603958
R25863 VGND VGND.n5156 0.0603958
R25864 VGND.n5144 VGND 0.0603958
R25865 VGND.n5139 VGND 0.0603958
R25866 VGND.n3490 VGND 0.0603958
R25867 VGND.n3506 VGND 0.0603958
R25868 VGND.n3508 VGND 0.0603958
R25869 VGND.n3508 VGND 0.0603958
R25870 VGND VGND.n9201 0.0603958
R25871 VGND.n2186 VGND 0.0603958
R25872 VGND.n2192 VGND 0.0603958
R25873 VGND.n2196 VGND 0.0603958
R25874 VGND.n2203 VGND 0.0603958
R25875 VGND VGND.n2620 0.0603958
R25876 VGND.n2615 VGND 0.0603958
R25877 VGND.n2588 VGND 0.0603958
R25878 VGND.n2584 VGND 0.0603958
R25879 VGND VGND.n2583 0.0603958
R25880 VGND VGND.n2571 0.0603958
R25881 VGND VGND.n2570 0.0603958
R25882 VGND.n2559 VGND 0.0603958
R25883 VGND.n2544 VGND 0.0603958
R25884 VGND.n2483 VGND 0.0603958
R25885 VGND VGND.n2482 0.0603958
R25886 VGND.n2478 VGND 0.0603958
R25887 VGND.n2478 VGND 0.0603958
R25888 VGND VGND.n2477 0.0603958
R25889 VGND.n2471 VGND 0.0603958
R25890 VGND.n2457 VGND 0.0603958
R25891 VGND VGND.n2456 0.0603958
R25892 VGND VGND.n2455 0.0603958
R25893 VGND.n2451 VGND 0.0603958
R25894 VGND.n2443 VGND 0.0603958
R25895 VGND VGND.n2414 0.0603958
R25896 VGND VGND.n2410 0.0603958
R25897 VGND.n2409 VGND 0.0603958
R25898 VGND VGND.n2408 0.0603958
R25899 VGND.n9162 VGND 0.0603958
R25900 VGND.n9148 VGND 0.0603958
R25901 VGND.n9144 VGND 0.0603958
R25902 VGND VGND.n9143 0.0603958
R25903 VGND.n9133 VGND 0.0603958
R25904 VGND VGND.n9132 0.0603958
R25905 VGND.n9112 VGND 0.0603958
R25906 VGND VGND.n9125 0.0603958
R25907 VGND.n8189 VGND 0.0564896
R25908 VGND.n7500 VGND.n752 0.0548679
R25909 VGND.n6207 VGND.n6206 0.0548679
R25910 VGND.n4863 VGND.n4859 0.0525833
R25911 VGND.n4717 VGND.n4716 0.0525833
R25912 VGND.n3577 VGND.n3570 0.0525833
R25913 VGND.n3723 VGND.n3722 0.0525833
R25914 VGND.n3841 VGND.n3837 0.0525833
R25915 VGND.n1972 VGND.n1971 0.0525833
R25916 VGND.n7560 VGND.n7558 0.0525833
R25917 VGND.n7429 VGND.n7428 0.0525833
R25918 VGND.n6056 VGND.n6055 0.0525833
R25919 VGND.n5973 VGND.n5972 0.0525833
R25920 VGND.n9212 VGND.n9211 0.0525833
R25921 VGND.n2074 VGND 0.0512812
R25922 VGND.n3803 VGND 0.0512812
R25923 VGND.n1910 VGND 0.0512812
R25924 VGND.n717 VGND 0.0512812
R25925 VGND.n7485 VGND 0.0512812
R25926 VGND.n3511 VGND 0.0512812
R25927 VGND.n2632 VGND.n2631 0.0489687
R25928 VGND.n9093 VGND.n9092 0.0489687
R25929 VGND.n9089 VGND.n46 0.0489687
R25930 VGND.n3538 VGND.n3537 0.0489687
R25931 VGND.n7070 VGND.n7069 0.0486771
R25932 VGND.n8525 VGND.n8524 0.0486771
R25933 VGND.n405 VGND.n403 0.0486771
R25934 VGND.n5285 VGND.n5284 0.0486771
R25935 VGND.n536 VGND 0.0463917
R25936 VGND.n4133 VGND.n4132 0.0460729
R25937 VGND.n2082 VGND.n2081 0.0460729
R25938 VGND.n2643 VGND.n2642 0.0460729
R25939 VGND.n3703 VGND.n3702 0.0460729
R25940 VGND.n128 VGND.n127 0.0460729
R25941 VGND.n3815 VGND.n3814 0.0460729
R25942 VGND.n7532 VGND.n7531 0.0460729
R25943 VGND.n1836 VGND.n1835 0.0460729
R25944 VGND.n3520 VGND.n3519 0.0460729
R25945 VGND.n8312 VGND 0.0449123
R25946 VGND.n5315 VGND.n5310 0.0447708
R25947 VGND.n912 VGND.n911 0.0443356
R25948 VGND.n26 VGND.n25 0.0443356
R25949 VGND.n3574 VGND.n3573 0.0435976
R25950 VGND.n4967 VGND.n4966 0.0395625
R25951 VGND.n3377 VGND.n3376 0.0395625
R25952 VGND.n8855 VGND.n8854 0.0395625
R25953 VGND.n7757 VGND.n7756 0.0395625
R25954 VGND.n7629 VGND.n7628 0.0395625
R25955 VGND.n6273 VGND.n6272 0.0395625
R25956 VGND.n6571 VGND.n6570 0.0395625
R25957 VGND.n1785 VGND.n1784 0.0393514
R25958 VGND.n5345 VGND.n5342 0.0393514
R25959 VGND.n1753 VGND.n1749 0.0393514
R25960 VGND.n7224 VGND.n1328 0.0393514
R25961 VGND.n4819 VGND.n4818 0.0393514
R25962 VGND.n4139 VGND.n4138 0.0393514
R25963 VGND.n4493 VGND.n4176 0.0393514
R25964 VGND.n2088 VGND.n2087 0.0393514
R25965 VGND.n2763 VGND.n2759 0.0393514
R25966 VGND.n3617 VGND.n3616 0.0393514
R25967 VGND.n9047 VGND.n74 0.0393514
R25968 VGND.n3763 VGND.n3762 0.0393514
R25969 VGND.n8708 VGND.n205 0.0393514
R25970 VGND.n1999 VGND.n1998 0.0393514
R25971 VGND.n8093 VGND.n478 0.0393514
R25972 VGND.n7523 VGND.n721 0.0393514
R25973 VGND.n8152 VGND.n8146 0.0393514
R25974 VGND.n1319 VGND.n1144 0.0393514
R25975 VGND.n7497 VGND.n7496 0.0393514
R25976 VGND.n6783 VGND.n6782 0.0393514
R25977 VGND.n5616 VGND.n5615 0.0393514
R25978 VGND.n2515 VGND.n2334 0.0393514
R25979 VGND.n3479 VGND.n3478 0.0393514
R25980 VGND.n1849 VGND.n1848 0.0376622
R25981 VGND.n1775 VGND.n1774 0.0376622
R25982 VGND.n4760 VGND.n4759 0.0376622
R25983 VGND.n4699 VGND.n4698 0.0376622
R25984 VGND.n2100 VGND.n2099 0.0376622
R25985 VGND.n3629 VGND.n3628 0.0376622
R25986 VGND.n1869 VGND.n1868 0.0376622
R25987 VGND.n1961 VGND.n1960 0.0376622
R25988 VGND.n7515 VGND.n7514 0.0376622
R25989 VGND.n796 VGND.n795 0.0376622
R25990 VGND.n1694 VGND.n1693 0.0376622
R25991 VGND.n9207 VGND.n9206 0.0376622
R25992 VGND.n7110 VGND.n7109 0.0371114
R25993 VGND.n4587 VGND.n4579 0.0371114
R25994 VGND.n3012 VGND.n3011 0.0371114
R25995 VGND.n3173 VGND.n3172 0.0371114
R25996 VGND.n8571 VGND.n8570 0.0371114
R25997 VGND.n7987 VGND.n7986 0.0371114
R25998 VGND.n8312 VGND.n8311 0.0371114
R25999 VGND.n1203 VGND.n1196 0.0371114
R26000 VGND.n6933 VGND.n6931 0.0371114
R26001 VGND.n5456 VGND.n5455 0.0371114
R26002 VGND.n5754 VGND.n5752 0.0371114
R26003 VGND.n2399 VGND.n2391 0.0371114
R26004 VGND.n3898 VGND.n153 0.0370003
R26005 VGND.n1686 VGND.n1685 0.0370003
R26006 VGND.n7215 VGND.n7214 0.0369583
R26007 VGND.n4506 VGND.n4505 0.0369583
R26008 VGND.n9035 VGND.n9034 0.0369583
R26009 VGND.n8082 VGND.n8081 0.0369583
R26010 VGND.n8199 VGND.n8198 0.0369583
R26011 VGND.n1307 VGND.n1306 0.0369583
R26012 VGND.n5356 VGND.n5355 0.0369583
R26013 VGND.n2506 VGND.n2505 0.0369583
R26014 VGND.n4481 VGND 0.0347603
R26015 VGND.n7914 VGND 0.0347603
R26016 VGND VGND.n2543 0.0347603
R26017 VGND.n4772 VGND 0.0343542
R26018 VGND.n4890 VGND 0.0343542
R26019 VGND VGND.n5083 0.0343542
R26020 VGND.n7184 VGND 0.0343542
R26021 VGND.n4535 VGND 0.0343542
R26022 VGND.n1452 VGND 0.0343542
R26023 VGND.n2966 VGND 0.0343542
R26024 VGND.n2912 VGND 0.0343542
R26025 VGND.n7819 VGND 0.0343542
R26026 VGND.n8404 VGND 0.0343542
R26027 VGND.n8373 VGND 0.0343542
R26028 VGND.n677 VGND 0.0343542
R26029 VGND.n621 VGND 0.0343542
R26030 VGND.n8245 VGND 0.0343542
R26031 VGND.n8174 VGND 0.0343542
R26032 VGND.n8279 VGND 0.0343542
R26033 VGND.n7390 VGND 0.0343542
R26034 VGND.n1094 VGND 0.0343542
R26035 VGND.n1273 VGND 0.0343542
R26036 VGND.n6333 VGND 0.0343542
R26037 VGND.n6281 VGND 0.0343542
R26038 VGND.n6860 VGND 0.0343542
R26039 VGND.n1536 VGND 0.0343542
R26040 VGND.n6585 VGND 0.0343542
R26041 VGND VGND.n5406 0.0343542
R26042 VGND.n5930 VGND 0.0343542
R26043 VGND.n5501 VGND 0.0343542
R26044 VGND VGND.n3507 0.0343542
R26045 VGND VGND.n2284 0.0343542
R26046 VGND.n2411 VGND 0.0343542
R26047 VGND.n9123 VGND 0.0343542
R26048 VGND VGND.n4812 0.0330521
R26049 VGND VGND.n4903 0.0330521
R26050 VGND.n4033 VGND 0.0330521
R26051 VGND.n7169 VGND 0.0330521
R26052 VGND.n4663 VGND 0.0330521
R26053 VGND VGND.n4443 0.0330521
R26054 VGND VGND.n4550 0.0330521
R26055 VGND.n3426 VGND 0.0330521
R26056 VGND VGND.n3210 0.0330521
R26057 VGND VGND.n2812 0.0330521
R26058 VGND.n8906 VGND 0.0330521
R26059 VGND.n8978 VGND 0.0330521
R26060 VGND.n3068 VGND 0.0330521
R26061 VGND VGND.n3876 0.0330521
R26062 VGND.n8736 VGND 0.0330521
R26063 VGND.n8622 VGND 0.0330521
R26064 VGND VGND.n1992 0.0330521
R26065 VGND.n7809 VGND 0.0330521
R26066 VGND VGND.n7890 0.0330521
R26067 VGND.n8039 VGND 0.0330521
R26068 VGND.n7682 VGND 0.0330521
R26069 VGND.n8251 VGND 0.0330521
R26070 VGND.n450 VGND 0.0330521
R26071 VGND.n7392 VGND 0.0330521
R26072 VGND VGND.n1100 0.0330521
R26073 VGND.n1271 VGND 0.0330521
R26074 VGND VGND.n6255 0.0330521
R26075 VGND VGND.n6355 0.0330521
R26076 VGND.n6856 VGND 0.0330521
R26077 VGND.n1758 VGND 0.0330521
R26078 VGND.n6627 VGND 0.0330521
R26079 VGND VGND.n6697 0.0330521
R26080 VGND.n5401 VGND 0.0330521
R26081 VGND.n5939 VGND 0.0330521
R26082 VGND VGND.n5563 0.0330521
R26083 VGND VGND.n5677 0.0330521
R26084 VGND VGND.n16 0.0330521
R26085 VGND.n2571 VGND 0.0330521
R26086 VGND.n2456 VGND 0.0330521
R26087 VGND.n6532 VGND.n6531 0.0325946
R26088 VGND.n5091 VGND.n5090 0.0325946
R26089 VGND.n4068 VGND.n4067 0.0325946
R26090 VGND.n6984 VGND.n1389 0.0325946
R26091 VGND.n4327 VGND.n4325 0.0325946
R26092 VGND.n2891 VGND.n2890 0.0325946
R26093 VGND.n2138 VGND.n2137 0.0325946
R26094 VGND.n3140 VGND.n3138 0.0325946
R26095 VGND.n114 VGND.n113 0.0325946
R26096 VGND.n8557 VGND.n8556 0.0325946
R26097 VGND.n145 VGND.n144 0.0325946
R26098 VGND.n8431 VGND.n301 0.0325946
R26099 VGND.n552 VGND.n551 0.0325946
R26100 VGND.n419 VGND.n417 0.0325946
R26101 VGND.n592 VGND.n591 0.0325946
R26102 VGND.n1171 VGND.n1169 0.0325946
R26103 VGND.n6946 VGND.n1580 0.0325946
R26104 VGND.n2157 VGND.n2156 0.0325946
R26105 VGND.n5316 VGND.n5306 0.0325946
R26106 VGND.n2365 VGND.n2363 0.0325946
R26107 VGND.n1463 VGND.n1461 0.0317953
R26108 VGND.n2980 VGND.n2978 0.0317953
R26109 VGND.n3186 VGND.n3185 0.0317953
R26110 VGND.n8417 VGND.n8416 0.0317953
R26111 VGND.n6963 VGND.n6961 0.0317953
R26112 VGND.n5085 VGND 0.03175
R26113 VGND.n4028 VGND 0.03175
R26114 VGND.n4023 VGND 0.03175
R26115 VGND.n7193 VGND 0.03175
R26116 VGND.n7170 VGND 0.03175
R26117 VGND.n7119 VGND 0.03175
R26118 VGND VGND.n4103 0.03175
R26119 VGND VGND.n4159 0.03175
R26120 VGND VGND.n4389 0.03175
R26121 VGND.n4419 VGND 0.03175
R26122 VGND.n4475 VGND 0.03175
R26123 VGND VGND.n4523 0.03175
R26124 VGND.n4635 VGND 0.03175
R26125 VGND VGND.n4567 0.03175
R26126 VGND.n1434 VGND 0.03175
R26127 VGND.n1425 VGND 0.03175
R26128 VGND.n3425 VGND 0.03175
R26129 VGND.n3266 VGND 0.03175
R26130 VGND.n3262 VGND 0.03175
R26131 VGND.n2756 VGND 0.03175
R26132 VGND.n2847 VGND 0.03175
R26133 VGND.n2965 VGND 0.03175
R26134 VGND.n2931 VGND 0.03175
R26135 VGND.n3688 VGND 0.03175
R26136 VGND.n3712 VGND.n3711 0.03175
R26137 VGND.n8924 VGND 0.03175
R26138 VGND.n8955 VGND 0.03175
R26139 VGND.n3041 VGND 0.03175
R26140 VGND.n2727 VGND 0.03175
R26141 VGND.n2697 VGND 0.03175
R26142 VGND VGND.n3783 0.03175
R26143 VGND.n3822 VGND.n3821 0.03175
R26144 VGND VGND.n3877 0.03175
R26145 VGND VGND.n3885 0.03175
R26146 VGND.n3925 VGND 0.03175
R26147 VGND VGND.n161 0.03175
R26148 VGND.n8780 VGND 0.03175
R26149 VGND.n8766 VGND 0.03175
R26150 VGND.n8733 VGND 0.03175
R26151 VGND.n8584 VGND 0.03175
R26152 VGND.n1986 VGND.n1985 0.03175
R26153 VGND.n1953 VGND 0.03175
R26154 VGND.n7808 VGND 0.03175
R26155 VGND.n7781 VGND 0.03175
R26156 VGND VGND.n7889 0.03175
R26157 VGND.n8390 VGND 0.03175
R26158 VGND.n696 VGND 0.03175
R26159 VGND.n7541 VGND.n7540 0.03175
R26160 VGND.n7681 VGND 0.03175
R26161 VGND.n7636 VGND 0.03175
R26162 VGND VGND.n8260 0.03175
R26163 VGND.n1071 VGND 0.03175
R26164 VGND.n1117 VGND 0.03175
R26165 VGND.n1262 VGND 0.03175
R26166 VGND.n1240 VGND 0.03175
R26167 VGND.n1218 VGND 0.03175
R26168 VGND.n949 VGND 0.03175
R26169 VGND.n941 VGND 0.03175
R26170 VGND VGND.n6100 0.03175
R26171 VGND.n6221 VGND 0.03175
R26172 VGND.n6244 VGND 0.03175
R26173 VGND VGND.n6341 0.03175
R26174 VGND.n6896 VGND 0.03175
R26175 VGND.n1523 VGND 0.03175
R26176 VGND.n1730 VGND 0.03175
R26177 VGND.n1765 VGND.n1764 0.03175
R26178 VGND.n6034 VGND 0.03175
R26179 VGND.n6626 VGND 0.03175
R26180 VGND.n6698 VGND 0.03175
R26181 VGND.n5253 VGND 0.03175
R26182 VGND.n1822 VGND 0.03175
R26183 VGND.n1844 VGND.n1843 0.03175
R26184 VGND.n5538 VGND 0.03175
R26185 VGND.n2192 VGND 0.03175
R26186 VGND.n2584 VGND 0.03175
R26187 VGND.n2544 VGND 0.03175
R26188 VGND.n2455 VGND 0.03175
R26189 VGND.n9132 VGND 0.03175
R26190 VGND.n5796 VGND.n5795 0.0315717
R26191 VGND.n9099 VGND.n22 0.0315717
R26192 VGND.n1848 VGND.n1847 0.0309054
R26193 VGND.n6732 VGND.n6731 0.0309054
R26194 VGND.n6731 VGND.n6730 0.0309054
R26195 VGND.n1774 VGND.n1773 0.0309054
R26196 VGND.n6514 VGND.n6513 0.0309054
R26197 VGND.n3998 VGND.n3997 0.0309054
R26198 VGND.n1328 VGND.n1327 0.0309054
R26199 VGND.n4759 VGND.n4758 0.0309054
R26200 VGND.n4988 VGND.n4987 0.0309054
R26201 VGND.n4698 VGND.n4697 0.0309054
R26202 VGND.n4484 VGND.n4483 0.0309054
R26203 VGND.n4176 VGND.n4175 0.0309054
R26204 VGND.n4337 VGND.n4336 0.0309054
R26205 VGND.n2099 VGND.n2098 0.0309054
R26206 VGND.n3238 VGND.n3237 0.0309054
R26207 VGND.n2638 VGND.n2637 0.0309054
R26208 VGND.n3628 VGND.n3627 0.0309054
R26209 VGND.n9009 VGND.n9008 0.0309054
R26210 VGND.n123 VGND.n122 0.0309054
R26211 VGND.n1868 VGND.n1867 0.0309054
R26212 VGND.n198 VGND.n197 0.0309054
R26213 VGND.n8798 VGND.n8797 0.0309054
R26214 VGND.n1960 VGND.n1959 0.0309054
R26215 VGND.n7909 VGND.n7908 0.0309054
R26216 VGND.n564 VGND.n563 0.0309054
R26217 VGND.n7514 VGND.n7513 0.0309054
R26218 VGND.n458 VGND.n457 0.0309054
R26219 VGND.n8146 VGND.n8145 0.0309054
R26220 VGND.n7702 VGND.n7701 0.0309054
R26221 VGND.n1137 VGND.n1136 0.0309054
R26222 VGND.n850 VGND.n849 0.0309054
R26223 VGND.n6174 VGND.n6173 0.0309054
R26224 VGND.n1597 VGND.n1596 0.0309054
R26225 VGND.n1681 VGND.n1680 0.0309054
R26226 VGND.n2281 VGND.n2280 0.0309054
R26227 VGND.n5610 VGND.n5609 0.0309054
R26228 VGND.n5609 VGND.n5608 0.0309054
R26229 VGND.n2320 VGND.n2319 0.0309054
R26230 VGND.n2334 VGND.n2333 0.0309054
R26231 VGND.n9230 VGND.n9229 0.0309054
R26232 VGND.n9206 VGND.n9205 0.0309054
R26233 VGND.n5827 VGND.n5826 0.0309054
R26234 VGND.n5119 VGND.n5118 0.0309054
R26235 VGND.n5092 VGND 0.0304479
R26236 VGND.n6983 VGND 0.0304479
R26237 VGND.n2892 VGND 0.0304479
R26238 VGND.n3139 VGND 0.0304479
R26239 VGND VGND.n8558 0.0304479
R26240 VGND.n8430 VGND 0.0304479
R26241 VGND.n418 VGND 0.0304479
R26242 VGND.n1170 VGND 0.0304479
R26243 VGND.n6945 VGND 0.0304479
R26244 VGND.n5766 VGND 0.0304479
R26245 VGND.n2364 VGND 0.0304479
R26246 VGND.n6513 VGND.n6509 0.0292162
R26247 VGND.n6995 VGND.n6994 0.0292162
R26248 VGND.n4987 VGND.n4043 0.0292162
R26249 VGND.n4585 VGND.n4581 0.0292162
R26250 VGND.n4336 VGND.n4225 0.0292162
R26251 VGND.n3016 VGND.n3015 0.0292162
R26252 VGND.n2639 VGND.n2638 0.0292162
R26253 VGND.n3177 VGND.n3176 0.0292162
R26254 VGND.n124 VGND.n123 0.0292162
R26255 VGND.n8443 VGND.n8442 0.0292162
R26256 VGND.n8797 VGND.n8796 0.0292162
R26257 VGND.n7977 VGND.n7970 0.0292162
R26258 VGND.n563 VGND.n560 0.0292162
R26259 VGND.n8316 VGND.n8315 0.0292162
R26260 VGND.n7701 VGND.n7700 0.0292162
R26261 VGND.n1201 VGND.n1198 0.0292162
R26262 VGND.n845 VGND.n844 0.0292162
R26263 VGND.n6929 VGND.n6923 0.0292162
R26264 VGND.n1574 VGND.n1573 0.0292162
R26265 VGND.n6460 VGND.n6459 0.0292162
R26266 VGND.n2280 VGND.n2166 0.0292162
R26267 VGND.n5460 VGND.n5459 0.0292162
R26268 VGND.n5750 VGND.n5744 0.0292162
R26269 VGND.n5743 VGND.n5742 0.0292162
R26270 VGND.n2397 VGND.n2393 0.0292162
R26271 VGND.n5820 VGND.n5819 0.0292162
R26272 VGND.n7207 VGND.n7204 0.0291458
R26273 VGND.n4498 VGND.n4496 0.0291458
R26274 VGND.n3229 VGND.n3228 0.0291458
R26275 VGND.n9027 VGND.n9025 0.0291458
R26276 VGND.n8660 VGND.n8658 0.0291458
R26277 VGND.n8074 VGND.n8072 0.0291458
R26278 VGND.n8137 VGND.n8136 0.0291458
R26279 VGND.n1301 VGND.n1299 0.0291458
R26280 VGND.n6805 VGND.n6803 0.0291458
R26281 VGND.n5350 VGND.n5348 0.0291458
R26282 VGND.n5597 VGND.n5596 0.0291458
R26283 VGND.n2498 VGND.n2495 0.0291458
R26284 VGND.n8438 VGND.n8437 0.0289937
R26285 VGND.n2039 VGND.n2038 0.0289937
R26286 VGND.n4357 VGND 0.0278438
R26287 VGND.n3914 VGND 0.0278438
R26288 VGND.n7333 VGND 0.0278438
R26289 VGND.n5888 VGND 0.0278438
R26290 VGND VGND.n2247 0.0278438
R26291 VGND.n2765 VGND 0.0265417
R26292 VGND VGND.n2775 0.0265417
R26293 VGND.n8696 VGND 0.0265417
R26294 VGND.n6813 VGND 0.0265417
R26295 VGND.n5632 VGND 0.0265417
R26296 VGND.n4517 VGND.n4514 0.0264488
R26297 VGND.n8193 VGND.n8192 0.0264488
R26298 VGND.n1317 VGND.n1297 0.0264488
R26299 VGND.n2513 VGND.n2493 0.0264488
R26300 VGND.n6730 VGND.n6729 0.0258378
R26301 VGND.n6514 VGND.n6512 0.0258378
R26302 VGND.n1356 VGND.n1355 0.0258378
R26303 VGND.n7243 VGND.n7242 0.0258378
R26304 VGND.n4188 VGND.n4187 0.0258378
R26305 VGND.n1386 VGND.n1385 0.0258378
R26306 VGND.n1559 VGND.n1558 0.0258378
R26307 VGND.n1563 VGND.n1562 0.0258378
R26308 VGND.n2882 VGND.n2881 0.0258378
R26309 VGND.n3232 VGND.n3231 0.0258378
R26310 VGND.n3135 VGND.n3134 0.0258378
R26311 VGND.n9054 VGND.n9053 0.0258378
R26312 VGND.n260 VGND.n259 0.0258378
R26313 VGND.n8666 VGND.n8665 0.0258378
R26314 VGND.n297 VGND.n296 0.0258378
R26315 VGND.n465 VGND.n464 0.0258378
R26316 VGND.n8132 VGND.n8128 0.0258378
R26317 VGND.n415 VGND.n414 0.0258378
R26318 VGND.n312 VGND.n311 0.0258378
R26319 VGND.n8327 VGND.n8326 0.0258378
R26320 VGND.n7264 VGND.n7263 0.0258378
R26321 VGND.n1166 VGND.n1165 0.0258378
R26322 VGND.n7303 VGND.n7302 0.0258378
R26323 VGND.n882 VGND.n881 0.0258378
R26324 VGND.n1576 VGND.n1575 0.0258378
R26325 VGND.n1548 VGND.n1547 0.0258378
R26326 VGND.n1605 VGND.n1604 0.0258378
R26327 VGND.n1669 VGND.n1668 0.0258378
R26328 VGND.n2281 VGND.n2279 0.0258378
R26329 VGND.n5302 VGND.n5301 0.0258378
R26330 VGND.n5778 VGND.n5777 0.0258378
R26331 VGND.n5782 VGND.n5781 0.0258378
R26332 VGND.n2360 VGND.n2359 0.0258378
R26333 VGND.n29 VGND.n28 0.0258378
R26334 VGND.n2527 VGND.n2526 0.0258378
R26335 VGND.n5864 VGND.n5863 0.0258378
R26336 VGND.n7222 VGND.n7202 0.0256464
R26337 VGND.n2778 VGND.n2776 0.0256464
R26338 VGND.n9045 VGND.n76 0.0256464
R26339 VGND.n8706 VGND.n8651 0.0256464
R26340 VGND.n8091 VGND.n8070 0.0256464
R26341 VGND.n6822 VGND.n6819 0.0256464
R26342 VGND.n5369 VGND.n5368 0.0256464
R26343 VGND.n5641 VGND.n5639 0.0256464
R26344 VGND.n4976 VGND.n4975 0.0252396
R26345 VGND.n4006 VGND.n4004 0.0252396
R26346 VGND.n5093 VGND.n5092 0.0252396
R26347 VGND.n4110 VGND 0.0252396
R26348 VGND.n4131 VGND.n4130 0.0252396
R26349 VGND.n4328 VGND.n4318 0.0252396
R26350 VGND.n4212 VGND.n4210 0.0252396
R26351 VGND.n6983 VGND.n6982 0.0252396
R26352 VGND.n2080 VGND.n2079 0.0252396
R26353 VGND.n3364 VGND.n3363 0.0252396
R26354 VGND.n2893 VGND.n2892 0.0252396
R26355 VGND.n3700 VGND.n3699 0.0252396
R26356 VGND.n8842 VGND.n8841 0.0252396
R26357 VGND.n3139 VGND.n2665 0.0252396
R26358 VGND.n3812 VGND.n3811 0.0252396
R26359 VGND.n3901 VGND.n3900 0.0252396
R26360 VGND.n8719 VGND 0.0252396
R26361 VGND.n8656 VGND.n8655 0.0252396
R26362 VGND.n8558 VGND.n257 0.0252396
R26363 VGND.n7747 VGND.n7746 0.0252396
R26364 VGND.n7924 VGND 0.0252396
R26365 VGND.n7917 VGND.n7915 0.0252396
R26366 VGND.n8029 VGND 0.0252396
R26367 VGND.n8430 VGND.n8429 0.0252396
R26368 VGND.n7615 VGND.n7614 0.0252396
R26369 VGND.n418 VGND.n309 0.0252396
R26370 VGND.n381 VGND 0.0252396
R26371 VGND.n7491 VGND.n7490 0.0252396
R26372 VGND.n870 VGND.n869 0.0252396
R26373 VGND.n1129 VGND.n1126 0.0252396
R26374 VGND.n1170 VGND.n889 0.0252396
R26375 VGND.n6153 VGND.n6152 0.0252396
R26376 VGND.n1683 VGND.n1679 0.0252396
R26377 VGND.n6801 VGND.n6800 0.0252396
R26378 VGND.n6945 VGND.n1476 0.0252396
R26379 VGND.n6556 VGND.n6555 0.0252396
R26380 VGND.n6722 VGND.n6720 0.0252396
R26381 VGND.n5315 VGND.n5314 0.0252396
R26382 VGND.n1833 VGND.n1832 0.0252396
R26383 VGND.n5875 VGND.n5874 0.0252396
R26384 VGND.n5601 VGND.n5599 0.0252396
R26385 VGND.n5766 VGND.n5126 0.0252396
R26386 VGND.n3517 VGND.n3516 0.0252396
R26387 VGND.n2261 VGND.n2260 0.0252396
R26388 VGND.n2316 VGND.n2314 0.0252396
R26389 VGND.n2364 VGND.n21 0.0252396
R26390 VGND.n987 VGND 0.0250613
R26391 VGND.n1793 VGND.n1792 0.0241486
R26392 VGND.n6748 VGND.n6747 0.0241486
R26393 VGND.n1701 VGND.n1700 0.0241486
R26394 VGND.n7247 VGND.n7246 0.0241486
R26395 VGND.n4804 VGND.n4803 0.0241486
R26396 VGND.n4155 VGND.n4154 0.0241486
R26397 VGND.n4192 VGND.n4191 0.0241486
R26398 VGND.n3453 VGND.n3452 0.0241486
R26399 VGND.n9079 VGND.n9078 0.0241486
R26400 VGND.n3588 VGND.n3587 0.0241486
R26401 VGND.n9057 VGND.n9056 0.0241486
R26402 VGND.n3734 VGND.n3733 0.0241486
R26403 VGND.n8678 VGND.n8677 0.0241486
R26404 VGND.n2007 VGND.n2006 0.0241486
R26405 VGND.n468 VGND.n467 0.0241486
R26406 VGND.n725 VGND.n724 0.0241486
R26407 VGND.n8141 VGND.n8140 0.0241486
R26408 VGND.n7267 VGND.n7266 0.0241486
R26409 VGND.n782 VGND.n781 0.0241486
R26410 VGND.n6104 VGND.n6103 0.0241486
R26411 VGND.n5628 VGND.n5472 0.0241486
R26412 VGND.n2531 VGND.n2530 0.0241486
R26413 VGND.n3482 VGND.n3481 0.0241486
R26414 VGND.n4847 VGND.n4845 0.0239375
R26415 VGND.n4978 VGND.n4977 0.0239375
R26416 VGND VGND.n4042 0.0239375
R26417 VGND.n5015 VGND 0.0239375
R26418 VGND VGND.n5084 0.0239375
R26419 VGND.n4029 VGND 0.0239375
R26420 VGND.n7192 VGND 0.0239375
R26421 VGND.n7160 VGND 0.0239375
R26422 VGND.n4731 VGND.n4729 0.0239375
R26423 VGND VGND.n4224 0.0239375
R26424 VGND.n4390 VGND 0.0239375
R26425 VGND.n4524 VGND 0.0239375
R26426 VGND.n4634 VGND 0.0239375
R26427 VGND.n3562 VGND.n3561 0.0239375
R26428 VGND.n3362 VGND.n3361 0.0239375
R26429 VGND.n2930 VGND 0.0239375
R26430 VGND.n3715 VGND.n3714 0.0239375
R26431 VGND.n8840 VGND.n8839 0.0239375
R26432 VGND VGND.n3053 0.0239375
R26433 VGND.n3826 VGND.n3824 0.0239375
R26434 VGND.n3899 VGND.n3898 0.0239375
R26435 VGND.n156 VGND 0.0239375
R26436 VGND.n8483 VGND 0.0239375
R26437 VGND.n1983 VGND.n1982 0.0239375
R26438 VGND.n7763 VGND 0.0239375
R26439 VGND.n7745 VGND.n7744 0.0239375
R26440 VGND.n566 VGND 0.0239375
R26441 VGND VGND.n7869 0.0239375
R26442 VGND.n8062 VGND 0.0239375
R26443 VGND.n8055 VGND 0.0239375
R26444 VGND.n8378 VGND 0.0239375
R26445 VGND.n7547 VGND.n7543 0.0239375
R26446 VGND VGND.n7581 0.0239375
R26447 VGND.n7613 VGND.n7612 0.0239375
R26448 VGND.n605 VGND 0.0239375
R26449 VGND.n7444 VGND.n7442 0.0239375
R26450 VGND.n872 VGND.n871 0.0239375
R26451 VGND.n884 VGND 0.0239375
R26452 VGND.n1289 VGND 0.0239375
R26453 VGND.n1259 VGND 0.0239375
R26454 VGND.n1221 VGND 0.0239375
R26455 VGND.n944 VGND 0.0239375
R26456 VGND.n6177 VGND.n6175 0.0239375
R26457 VGND VGND.n6468 0.0239375
R26458 VGND.n6826 VGND 0.0239375
R26459 VGND.n6069 VGND.n6068 0.0239375
R26460 VGND.n6554 VGND.n6553 0.0239375
R26461 VGND.n6516 VGND 0.0239375
R26462 VGND.n5998 VGND.n5997 0.0239375
R26463 VGND.n5873 VGND.n5872 0.0239375
R26464 VGND VGND.n5861 0.0239375
R26465 VGND.n9231 VGND.n0 0.0239375
R26466 VGND.n2263 VGND.n2262 0.0239375
R26467 VGND.n2283 VGND 0.0239375
R26468 VGND.n2482 VGND 0.0239375
R26469 VGND.n4012 VGND.n4011 0.0238078
R26470 VGND.n6727 VGND.n6726 0.0238078
R26471 VGND.n5606 VGND.n5605 0.0238078
R26472 VGND.n4481 VGND.n4480 0.0238078
R26473 VGND.n3244 VGND.n3236 0.0238078
R26474 VGND.n9018 VGND.n9014 0.0238078
R26475 VGND.n8717 VGND.n196 0.0238078
R26476 VGND.n7919 VGND.n7914 0.0238078
R26477 VGND.n8217 VGND.n456 0.0238078
R26478 VGND.n1134 VGND.n1133 0.0238078
R26479 VGND.n6795 VGND.n6793 0.0238078
R26480 VGND.n2543 VGND.n2318 0.0238078
R26481 VGND VGND.n803 0.0231359
R26482 VGND VGND.n6219 0.0231359
R26483 VGND VGND.n6017 0.0231359
R26484 VGND VGND.n4771 0.0226354
R26485 VGND.n4786 VGND 0.0226354
R26486 VGND.n4868 VGND 0.0226354
R26487 VGND.n4886 VGND 0.0226354
R26488 VGND.n4088 VGND 0.0226354
R26489 VGND VGND.n4902 0.0226354
R26490 VGND.n4907 VGND 0.0226354
R26491 VGND.n4917 VGND 0.0226354
R26492 VGND.n4944 VGND 0.0226354
R26493 VGND.n4078 VGND 0.0226354
R26494 VGND.n4077 VGND 0.0226354
R26495 VGND.n4980 VGND.n4978 0.0226354
R26496 VGND.n4989 VGND 0.0226354
R26497 VGND VGND.n5051 0.0226354
R26498 VGND.n5057 VGND 0.0226354
R26499 VGND.n5066 VGND 0.0226354
R26500 VGND VGND.n5081 0.0226354
R26501 VGND.n4030 VGND 0.0226354
R26502 VGND.n4022 VGND 0.0226354
R26503 VGND.n4021 VGND 0.0226354
R26504 VGND.n7183 VGND 0.0226354
R26505 VGND.n7174 VGND 0.0226354
R26506 VGND.n7161 VGND 0.0226354
R26507 VGND.n7148 VGND 0.0226354
R26508 VGND.n7137 VGND 0.0226354
R26509 VGND.n7062 VGND 0.0226354
R26510 VGND.n7044 VGND 0.0226354
R26511 VGND.n7017 VGND 0.0226354
R26512 VGND.n4104 VGND 0.0226354
R26513 VGND.n4687 VGND 0.0226354
R26514 VGND.n4684 VGND 0.0226354
R26515 VGND.n4674 VGND 0.0226354
R26516 VGND.n4669 VGND 0.0226354
R26517 VGND.n4664 VGND 0.0226354
R26518 VGND.n4244 VGND 0.0226354
R26519 VGND.n4273 VGND 0.0226354
R26520 VGND.n4283 VGND 0.0226354
R26521 VGND.n4292 VGND 0.0226354
R26522 VGND.n4332 VGND.n4330 0.0226354
R26523 VGND.n4338 VGND 0.0226354
R26524 VGND VGND.n4388 0.0226354
R26525 VGND VGND.n4429 0.0226354
R26526 VGND VGND.n4437 0.0226354
R26527 VGND.n4438 VGND 0.0226354
R26528 VGND VGND.n4455 0.0226354
R26529 VGND.n4456 VGND 0.0226354
R26530 VGND VGND.n4549 0.0226354
R26531 VGND.n4650 VGND 0.0226354
R26532 VGND.n4639 VGND 0.0226354
R26533 VGND.n4616 VGND 0.0226354
R26534 VGND.n1449 VGND 0.0226354
R26535 VGND.n1437 VGND 0.0226354
R26536 VGND.n1431 VGND 0.0226354
R26537 VGND.n1426 VGND 0.0226354
R26538 VGND.n1414 VGND 0.0226354
R26539 VGND.n2057 VGND 0.0226354
R26540 VGND.n2064 VGND 0.0226354
R26541 VGND VGND.n2069 0.0226354
R26542 VGND.n3449 VGND 0.0226354
R26543 VGND.n3430 VGND 0.0226354
R26544 VGND.n3417 VGND 0.0226354
R26545 VGND.n3402 VGND 0.0226354
R26546 VGND.n3395 VGND 0.0226354
R26547 VGND.n3361 VGND.n3360 0.0226354
R26548 VGND VGND.n2650 0.0226354
R26549 VGND.n3313 VGND 0.0226354
R26550 VGND.n3290 VGND 0.0226354
R26551 VGND.n3280 VGND 0.0226354
R26552 VGND.n3270 VGND 0.0226354
R26553 VGND.n3249 VGND 0.0226354
R26554 VGND.n2788 VGND 0.0226354
R26555 VGND.n2757 VGND 0.0226354
R26556 VGND.n2795 VGND 0.0226354
R26557 VGND VGND.n2811 0.0226354
R26558 VGND.n2813 VGND 0.0226354
R26559 VGND.n2824 VGND 0.0226354
R26560 VGND VGND.n2838 0.0226354
R26561 VGND.n2855 VGND 0.0226354
R26562 VGND.n2862 VGND 0.0226354
R26563 VGND.n2747 VGND 0.0226354
R26564 VGND.n2944 VGND 0.0226354
R26565 VGND.n2934 VGND 0.0226354
R26566 VGND.n2920 VGND 0.0226354
R26567 VGND.n2916 VGND 0.0226354
R26568 VGND.n2915 VGND 0.0226354
R26569 VGND.n3679 VGND 0.0226354
R26570 VGND VGND.n3687 0.0226354
R26571 VGND.n3655 VGND 0.0226354
R26572 VGND.n3640 VGND 0.0226354
R26573 VGND.n8904 VGND 0.0226354
R26574 VGND.n8894 VGND 0.0226354
R26575 VGND.n8886 VGND 0.0226354
R26576 VGND.n8873 VGND 0.0226354
R26577 VGND.n8839 VGND.n8838 0.0226354
R26578 VGND.n8938 VGND 0.0226354
R26579 VGND VGND.n8954 0.0226354
R26580 VGND VGND.n8977 0.0226354
R26581 VGND.n3036 VGND 0.0226354
R26582 VGND VGND.n3047 0.0226354
R26583 VGND VGND.n3067 0.0226354
R26584 VGND VGND.n3073 0.0226354
R26585 VGND.n3075 VGND 0.0226354
R26586 VGND.n3102 VGND 0.0226354
R26587 VGND.n2730 VGND 0.0226354
R26588 VGND VGND.n2669 0.0226354
R26589 VGND.n2700 VGND 0.0226354
R26590 VGND.n2688 VGND 0.0226354
R26591 VGND.n2685 VGND 0.0226354
R26592 VGND.n3784 VGND 0.0226354
R26593 VGND VGND.n3792 0.0226354
R26594 VGND VGND.n3799 0.0226354
R26595 VGND.n3800 VGND 0.0226354
R26596 VGND.n3844 VGND 0.0226354
R26597 VGND VGND.n3875 0.0226354
R26598 VGND.n3958 VGND 0.0226354
R26599 VGND.n3954 VGND 0.0226354
R26600 VGND.n3924 VGND 0.0226354
R26601 VGND.n8799 VGND 0.0226354
R26602 VGND.n8781 VGND 0.0226354
R26603 VGND.n8758 VGND 0.0226354
R26604 VGND.n8755 VGND 0.0226354
R26605 VGND.n8742 VGND 0.0226354
R26606 VGND.n8738 VGND 0.0226354
R26607 VGND.n8729 VGND 0.0226354
R26608 VGND.n8722 VGND 0.0226354
R26609 VGND.n8645 VGND 0.0226354
R26610 VGND.n8639 VGND 0.0226354
R26611 VGND.n8636 VGND 0.0226354
R26612 VGND.n8617 VGND 0.0226354
R26613 VGND.n8605 VGND 0.0226354
R26614 VGND.n8595 VGND 0.0226354
R26615 VGND.n8594 VGND 0.0226354
R26616 VGND.n8587 VGND 0.0226354
R26617 VGND.n8582 VGND 0.0226354
R26618 VGND.n8575 VGND 0.0226354
R26619 VGND.n8504 VGND 0.0226354
R26620 VGND.n8494 VGND 0.0226354
R26621 VGND.n8486 VGND 0.0226354
R26622 VGND.n8479 VGND 0.0226354
R26623 VGND.n8476 VGND 0.0226354
R26624 VGND.n8468 VGND 0.0226354
R26625 VGND VGND.n1895 0.0226354
R26626 VGND.n1896 VGND 0.0226354
R26627 VGND VGND.n1905 0.0226354
R26628 VGND VGND.n1906 0.0226354
R26629 VGND.n1956 VGND 0.0226354
R26630 VGND.n1951 VGND 0.0226354
R26631 VGND.n1929 VGND 0.0226354
R26632 VGND.n7790 VGND 0.0226354
R26633 VGND.n7784 VGND 0.0226354
R26634 VGND.n7768 VGND 0.0226354
R26635 VGND.n7744 VGND.n7743 0.0226354
R26636 VGND VGND.n565 0.0226354
R26637 VGND.n7829 VGND 0.0226354
R26638 VGND VGND.n7833 0.0226354
R26639 VGND.n7834 VGND 0.0226354
R26640 VGND.n7849 VGND 0.0226354
R26641 VGND.n7859 VGND 0.0226354
R26642 VGND.n7870 VGND 0.0226354
R26643 VGND VGND.n7888 0.0226354
R26644 VGND.n7927 VGND 0.0226354
R26645 VGND.n7922 VGND 0.0226354
R26646 VGND.n8043 VGND 0.0226354
R26647 VGND.n8032 VGND 0.0226354
R26648 VGND.n8024 VGND 0.0226354
R26649 VGND.n8002 VGND 0.0226354
R26650 VGND.n7990 VGND 0.0226354
R26651 VGND.n8394 VGND 0.0226354
R26652 VGND.n8393 VGND 0.0226354
R26653 VGND.n8389 VGND 0.0226354
R26654 VGND.n8374 VGND 0.0226354
R26655 VGND.n8372 VGND 0.0226354
R26656 VGND.n8368 VGND 0.0226354
R26657 VGND.n714 VGND 0.0226354
R26658 VGND.n7582 VGND 0.0226354
R26659 VGND VGND.n7597 0.0226354
R26660 VGND.n7672 VGND 0.0226354
R26661 VGND.n7668 VGND 0.0226354
R26662 VGND.n7652 VGND 0.0226354
R26663 VGND.n7639 VGND 0.0226354
R26664 VGND.n7612 VGND.n7611 0.0226354
R26665 VGND.n7703 VGND 0.0226354
R26666 VGND.n665 VGND 0.0226354
R26667 VGND.n620 VGND 0.0226354
R26668 VGND.n618 VGND 0.0226354
R26669 VGND.n8178 VGND 0.0226354
R26670 VGND VGND.n8262 0.0226354
R26671 VGND.n8273 VGND 0.0226354
R26672 VGND.n8307 VGND 0.0226354
R26673 VGND.n395 VGND 0.0226354
R26674 VGND.n386 VGND 0.0226354
R26675 VGND.n359 VGND 0.0226354
R26676 VGND.n356 VGND 0.0226354
R26677 VGND.n353 VGND 0.0226354
R26678 VGND.n7468 VGND 0.0226354
R26679 VGND.n7478 VGND 0.0226354
R26680 VGND.n7425 VGND 0.0226354
R26681 VGND.n7414 VGND 0.0226354
R26682 VGND.n7396 VGND 0.0226354
R26683 VGND.n7389 VGND 0.0226354
R26684 VGND.n7357 VGND 0.0226354
R26685 VGND.n7347 VGND 0.0226354
R26686 VGND.n874 VGND.n872 0.0226354
R26687 VGND VGND.n883 0.0226354
R26688 VGND.n1020 VGND 0.0226354
R26689 VGND VGND.n1049 0.0226354
R26690 VGND VGND.n1092 0.0226354
R26691 VGND VGND.n1099 0.0226354
R26692 VGND.n1110 VGND 0.0226354
R26693 VGND.n1294 VGND 0.0226354
R26694 VGND.n1286 VGND 0.0226354
R26695 VGND.n1263 VGND 0.0226354
R26696 VGND.n1255 VGND 0.0226354
R26697 VGND.n1244 VGND 0.0226354
R26698 VGND.n1226 VGND 0.0226354
R26699 VGND.n977 VGND 0.0226354
R26700 VGND.n959 VGND 0.0226354
R26701 VGND.n950 VGND 0.0226354
R26702 VGND.n938 VGND 0.0226354
R26703 VGND.n933 VGND 0.0226354
R26704 VGND.n6135 VGND 0.0226354
R26705 VGND.n6215 VGND 0.0226354
R26706 VGND.n6230 VGND 0.0226354
R26707 VGND.n6238 VGND 0.0226354
R26708 VGND VGND.n6254 0.0226354
R26709 VGND.n6305 VGND 0.0226354
R26710 VGND.n6293 VGND 0.0226354
R26711 VGND.n6288 VGND 0.0226354
R26712 VGND.n6284 VGND 0.0226354
R26713 VGND.n6278 VGND 0.0226354
R26714 VGND.n6469 VGND 0.0226354
R26715 VGND.n6447 VGND 0.0226354
R26716 VGND.n6396 VGND 0.0226354
R26717 VGND.n6394 VGND 0.0226354
R26718 VGND.n6392 VGND 0.0226354
R26719 VGND.n6386 VGND 0.0226354
R26720 VGND.n6380 VGND 0.0226354
R26721 VGND VGND.n6873 0.0226354
R26722 VGND.n6891 VGND 0.0226354
R26723 VGND.n6908 VGND 0.0226354
R26724 VGND.n1526 VGND 0.0226354
R26725 VGND.n1500 VGND 0.0226354
R26726 VGND.n1495 VGND 0.0226354
R26727 VGND.n1720 VGND 0.0226354
R26728 VGND.n6037 VGND 0.0226354
R26729 VGND.n6025 VGND 0.0226354
R26730 VGND.n6020 VGND 0.0226354
R26731 VGND.n6622 VGND 0.0226354
R26732 VGND.n6598 VGND 0.0226354
R26733 VGND.n6593 VGND 0.0226354
R26734 VGND.n6589 VGND 0.0226354
R26735 VGND.n6553 VGND.n6552 0.0226354
R26736 VGND VGND.n6515 0.0226354
R26737 VGND.n6635 VGND 0.0226354
R26738 VGND.n6652 VGND 0.0226354
R26739 VGND VGND.n6655 0.0226354
R26740 VGND VGND.n6672 0.0226354
R26741 VGND VGND.n6679 0.0226354
R26742 VGND.n6686 VGND 0.0226354
R26743 VGND.n6694 VGND 0.0226354
R26744 VGND VGND.n5400 0.0226354
R26745 VGND.n5416 VGND 0.0226354
R26746 VGND.n5426 VGND 0.0226354
R26747 VGND.n5440 VGND 0.0226354
R26748 VGND VGND.n5446 0.0226354
R26749 VGND.n5262 VGND 0.0226354
R26750 VGND.n5259 VGND 0.0226354
R26751 VGND.n5239 VGND 0.0226354
R26752 VGND.n1814 VGND 0.0226354
R26753 VGND.n5966 VGND 0.0226354
R26754 VGND.n5942 VGND 0.0226354
R26755 VGND.n5934 VGND 0.0226354
R26756 VGND.n5905 VGND 0.0226354
R26757 VGND.n5899 VGND 0.0226354
R26758 VGND.n5898 VGND 0.0226354
R26759 VGND.n5872 VGND.n5871 0.0226354
R26760 VGND.n5862 VGND 0.0226354
R26761 VGND.n5527 VGND 0.0226354
R26762 VGND VGND.n5537 0.0226354
R26763 VGND VGND.n5562 0.0226354
R26764 VGND.n5570 VGND 0.0226354
R26765 VGND.n5584 VGND 0.0226354
R26766 VGND.n5661 VGND 0.0226354
R26767 VGND VGND.n5676 0.0226354
R26768 VGND VGND.n5700 0.0226354
R26769 VGND.n5724 VGND 0.0226354
R26770 VGND.n5733 VGND 0.0226354
R26771 VGND.n5164 VGND 0.0226354
R26772 VGND.n5161 VGND 0.0226354
R26773 VGND.n5137 VGND 0.0226354
R26774 VGND.n3503 VGND 0.0226354
R26775 VGND VGND.n3506 0.0226354
R26776 VGND.n9186 VGND 0.0226354
R26777 VGND.n2188 VGND 0.0226354
R26778 VGND VGND.n2191 0.0226354
R26779 VGND.n2199 VGND 0.0226354
R26780 VGND.n2211 VGND 0.0226354
R26781 VGND VGND.n2223 0.0226354
R26782 VGND.n2224 VGND 0.0226354
R26783 VGND.n2265 VGND.n2263 0.0226354
R26784 VGND VGND.n2282 0.0226354
R26785 VGND.n2598 VGND 0.0226354
R26786 VGND.n2593 VGND 0.0226354
R26787 VGND.n2578 VGND 0.0226354
R26788 VGND.n2562 VGND 0.0226354
R26789 VGND.n2547 VGND 0.0226354
R26790 VGND.n2483 VGND 0.0226354
R26791 VGND VGND.n2340 0.0226354
R26792 VGND.n2460 VGND 0.0226354
R26793 VGND.n2457 VGND 0.0226354
R26794 VGND.n2447 VGND 0.0226354
R26795 VGND.n2420 VGND 0.0226354
R26796 VGND.n2414 VGND 0.0226354
R26797 VGND.n9152 VGND 0.0226354
R26798 VGND.n9148 VGND 0.0226354
R26799 VGND.n9143 VGND 0.0226354
R26800 VGND VGND.n9112 0.0226354
R26801 VGND.n9126 VGND 0.0226354
R26802 VGND.n6002 VGND.n6001 0.0224595
R26803 VGND.n5978 VGND.n5977 0.0224595
R26804 VGND.n6740 VGND.n6737 0.0224595
R26805 VGND.n6739 VGND.n6738 0.0224595
R26806 VGND.n6751 VGND.n6750 0.0224595
R26807 VGND.n6073 VGND.n6072 0.0224595
R26808 VGND.n6077 VGND.n6076 0.0224595
R26809 VGND.n1656 VGND.n1655 0.0224595
R26810 VGND.n6544 VGND.n6543 0.0224595
R26811 VGND.n7095 VGND.n7094 0.0224595
R26812 VGND.n5091 VGND.n1358 0.0224595
R26813 VGND.n7086 VGND.n7085 0.0224595
R26814 VGND.n7250 VGND.n7244 0.0224595
R26815 VGND.n7249 VGND.n7248 0.0224595
R26816 VGND.n7231 VGND.n7230 0.0224595
R26817 VGND.n4843 VGND.n4840 0.0224595
R26818 VGND.n4827 VGND.n4826 0.0224595
R26819 VGND.n4073 VGND.n4072 0.0224595
R26820 VGND.n4993 VGND.n4992 0.0224595
R26821 VGND.n4734 VGND.n4733 0.0224595
R26822 VGND.n4738 VGND.n4737 0.0224595
R26823 VGND.n4195 VGND.n4189 0.0224595
R26824 VGND.n4194 VGND.n4193 0.0224595
R26825 VGND.n4197 VGND.n4196 0.0224595
R26826 VGND.n6986 VGND.n1388 0.0224595
R26827 VGND.n6985 VGND.n6984 0.0224595
R26828 VGND.n1566 VGND.n1565 0.0224595
R26829 VGND.n4316 VGND.n4315 0.0224595
R26830 VGND.n4342 VGND.n4341 0.0224595
R26831 VGND.n3004 VGND.n3003 0.0224595
R26832 VGND.n2891 VGND.n2884 0.0224595
R26833 VGND.n2995 VGND.n2994 0.0224595
R26834 VGND.n3559 VGND.n3556 0.0224595
R26835 VGND.n3543 VGND.n3542 0.0224595
R26836 VGND.n9082 VGND.n50 0.0224595
R26837 VGND.n9081 VGND.n9080 0.0224595
R26838 VGND.n9074 VGND.n9073 0.0224595
R26839 VGND.n2128 VGND.n2127 0.0224595
R26840 VGND.n3356 VGND.n3354 0.0224595
R26841 VGND.n3159 VGND.n3158 0.0224595
R26842 VGND.n3141 VGND.n3140 0.0224595
R26843 VGND.n3150 VGND.n3149 0.0224595
R26844 VGND.n3595 VGND.n3594 0.0224595
R26845 VGND.n3599 VGND.n3598 0.0224595
R26846 VGND.n9060 VGND.n9055 0.0224595
R26847 VGND.n9059 VGND.n9058 0.0224595
R26848 VGND.n62 VGND.n61 0.0224595
R26849 VGND.n104 VGND.n103 0.0224595
R26850 VGND.n8834 VGND.n8832 0.0224595
R26851 VGND.n8553 VGND.n262 0.0224595
R26852 VGND.n8557 VGND.n8554 0.0224595
R26853 VGND.n8545 VGND.n8544 0.0224595
R26854 VGND.n3741 VGND.n3740 0.0224595
R26855 VGND.n3745 VGND.n3744 0.0224595
R26856 VGND.n8674 VGND.n8667 0.0224595
R26857 VGND.n8676 VGND.n8675 0.0224595
R26858 VGND.n8694 VGND.n8693 0.0224595
R26859 VGND.n150 VGND.n149 0.0224595
R26860 VGND.n8803 VGND.n8802 0.0224595
R26861 VGND.n8433 VGND.n299 0.0224595
R26862 VGND.n8432 VGND.n8431 0.0224595
R26863 VGND.n288 VGND.n287 0.0224595
R26864 VGND.n2014 VGND.n2013 0.0224595
R26865 VGND.n2018 VGND.n2017 0.0224595
R26866 VGND.n471 VGND.n466 0.0224595
R26867 VGND.n470 VGND.n469 0.0224595
R26868 VGND.n8101 VGND.n8100 0.0224595
R26869 VGND.n542 VGND.n541 0.0224595
R26870 VGND.n7738 VGND.n7736 0.0224595
R26871 VGND.n732 VGND.n731 0.0224595
R26872 VGND.n736 VGND.n735 0.0224595
R26873 VGND.n8208 VGND.n8138 0.0224595
R26874 VGND.n8207 VGND.n8206 0.0224595
R26875 VGND.n8117 VGND.n8116 0.0224595
R26876 VGND.n428 VGND.n427 0.0224595
R26877 VGND.n420 VGND.n419 0.0224595
R26878 VGND.n8329 VGND.n8325 0.0224595
R26879 VGND.n597 VGND.n596 0.0224595
R26880 VGND.n7707 VGND.n7706 0.0224595
R26881 VGND.n7270 VGND.n7265 0.0224595
R26882 VGND.n7269 VGND.n7268 0.0224595
R26883 VGND.n7282 VGND.n7281 0.0224595
R26884 VGND.n1182 VGND.n1181 0.0224595
R26885 VGND.n1172 VGND.n1171 0.0224595
R26886 VGND.n7305 VGND.n7301 0.0224595
R26887 VGND.n7447 VGND.n7446 0.0224595
R26888 VGND.n756 VGND.n755 0.0224595
R26889 VGND.n851 VGND.n850 0.0224595
R26890 VGND.n880 VGND.n860 0.0224595
R26891 VGND.n6948 VGND.n1578 0.0224595
R26892 VGND.n6947 VGND.n6946 0.0224595
R26893 VGND.n1551 VGND.n1550 0.0224595
R26894 VGND.n6170 VGND.n6168 0.0224595
R26895 VGND.n6172 VGND.n6096 0.0224595
R26896 VGND.n1610 VGND.n1606 0.0224595
R26897 VGND.n1609 VGND.n1608 0.0224595
R26898 VGND.n6772 VGND.n6771 0.0224595
R26899 VGND.n1680 VGND.n1667 0.0224595
R26900 VGND.n6473 VGND.n6472 0.0224595
R26901 VGND.n2268 VGND.n2267 0.0224595
R26902 VGND.n2273 VGND.n2272 0.0224595
R26903 VGND.n5318 VGND.n5304 0.0224595
R26904 VGND.n5317 VGND.n5316 0.0224595
R26905 VGND.n5329 VGND.n5326 0.0224595
R26906 VGND.n5769 VGND.n5467 0.0224595
R26907 VGND.n5768 VGND.n5767 0.0224595
R26908 VGND.n5785 VGND.n5784 0.0224595
R26909 VGND.n2378 VGND.n2377 0.0224595
R26910 VGND.n2366 VGND.n2365 0.0224595
R26911 VGND.n38 VGND.n37 0.0224595
R26912 VGND.n5482 VGND.n5479 0.0224595
R26913 VGND.n5481 VGND.n5480 0.0224595
R26914 VGND.n5626 VGND.n5625 0.0224595
R26915 VGND.n2534 VGND.n2528 0.0224595
R26916 VGND.n2533 VGND.n2532 0.0224595
R26917 VGND.n2322 VGND.n2321 0.0224595
R26918 VGND.n3531 VGND.n3530 0.0224595
R26919 VGND.n9228 VGND.n9227 0.0224595
R26920 VGND.n5120 VGND.n5119 0.0224595
R26921 VGND.n5865 VGND.n5121 0.0224595
R26922 VGND.n4966 VGND.n4965 0.0213333
R26923 VGND VGND.n5041 0.0213333
R26924 VGND.n5042 VGND 0.0213333
R26925 VGND.n5052 VGND 0.0213333
R26926 VGND.n5078 VGND 0.0213333
R26927 VGND.n7168 VGND 0.0213333
R26928 VGND.n7123 VGND 0.0213333
R26929 VGND.n4544 VGND 0.0213333
R26930 VGND.n3378 VGND.n3377 0.0213333
R26931 VGND.n8856 VGND.n8855 0.0213333
R26932 VGND.n3928 VGND 0.0213333
R26933 VGND.n3915 VGND.n3914 0.0213333
R26934 VGND.n7758 VGND.n7757 0.0213333
R26935 VGND.n7839 VGND 0.0213333
R26936 VGND.n8056 VGND 0.0213333
R26937 VGND.n8369 VGND 0.0213333
R26938 VGND VGND.n700 0.0213333
R26939 VGND.n7630 VGND.n7629 0.0213333
R26940 VGND.n653 VGND 0.0213333
R26941 VGND.n624 VGND 0.0213333
R26942 VGND.n8161 VGND 0.0213333
R26943 VGND.n7351 VGND 0.0213333
R26944 VGND.n1034 VGND 0.0213333
R26945 VGND VGND.n1070 0.0213333
R26946 VGND.n1277 VGND 0.0213333
R26947 VGND.n6274 VGND.n6273 0.0213333
R26948 VGND VGND.n6895 0.0213333
R26949 VGND.n6572 VGND.n6571 0.0213333
R26950 VGND.n5889 VGND.n5888 0.0213333
R26951 VGND.n2247 VGND.n2246 0.0213333
R26952 VGND.n2415 VGND 0.0213333
R26953 VGND.n5987 VGND.n5985 0.0207703
R26954 VGND.n1847 VGND.n1846 0.0207703
R26955 VGND.n6749 VGND.n6748 0.0207703
R26956 VGND.n6080 VGND.n6079 0.0207703
R26957 VGND.n1773 VGND.n1772 0.0207703
R26958 VGND.n6500 VGND.n6499 0.0207703
R26959 VGND.n6511 VGND.n6510 0.0207703
R26960 VGND.n1373 VGND.n1372 0.0207703
R26961 VGND.n7001 VGND.n1374 0.0207703
R26962 VGND.n7246 VGND.n7245 0.0207703
R26963 VGND.n4830 VGND.n4829 0.0207703
R26964 VGND.n4758 VGND.n4757 0.0207703
R26965 VGND.n4052 VGND.n4051 0.0207703
R26966 VGND.n5007 VGND.n5006 0.0207703
R26967 VGND.n4741 VGND.n4740 0.0207703
R26968 VGND.n4697 VGND.n4696 0.0207703
R26969 VGND.n4191 VGND.n4190 0.0207703
R26970 VGND.n1454 VGND.n1453 0.0207703
R26971 VGND.n1459 VGND.n1455 0.0207703
R26972 VGND.n4358 VGND.n4233 0.0207703
R26973 VGND.n4372 VGND.n4371 0.0207703
R26974 VGND.n2969 VGND.n2968 0.0207703
R26975 VGND.n2976 VGND.n2970 0.0207703
R26976 VGND.n3546 VGND.n3545 0.0207703
R26977 VGND.n2098 VGND.n2097 0.0207703
R26978 VGND.n3341 VGND.n3340 0.0207703
R26979 VGND.n2641 VGND.n2640 0.0207703
R26980 VGND.n2739 VGND.n2738 0.0207703
R26981 VGND.n3183 VGND.n2740 0.0207703
R26982 VGND.n3602 VGND.n3601 0.0207703
R26983 VGND.n3627 VGND.n3626 0.0207703
R26984 VGND.n8819 VGND.n8818 0.0207703
R26985 VGND.n126 VGND.n125 0.0207703
R26986 VGND.n274 VGND.n273 0.0207703
R26987 VGND.n8449 VGND.n275 0.0207703
R26988 VGND.n3748 VGND.n3747 0.0207703
R26989 VGND.n1867 VGND.n1866 0.0207703
R26990 VGND.n3889 VGND.n3888 0.0207703
R26991 VGND.n155 VGND.n154 0.0207703
R26992 VGND.n8407 VGND.n8406 0.0207703
R26993 VGND.n8414 VGND.n8408 0.0207703
R26994 VGND.n2021 VGND.n2020 0.0207703
R26995 VGND.n1959 VGND.n1958 0.0207703
R26996 VGND.n7723 VGND.n7722 0.0207703
R26997 VGND.n562 VGND.n561 0.0207703
R26998 VGND.n739 VGND.n738 0.0207703
R26999 VGND.n7513 VGND.n7512 0.0207703
R27000 VGND.n8140 VGND.n8139 0.0207703
R27001 VGND.n321 VGND.n320 0.0207703
R27002 VGND.n410 VGND.n322 0.0207703
R27003 VGND.n578 VGND.n577 0.0207703
R27004 VGND.n604 VGND.n603 0.0207703
R27005 VGND.n901 VGND.n900 0.0207703
R27006 VGND.n989 VGND.n902 0.0207703
R27007 VGND.n761 VGND.n760 0.0207703
R27008 VGND.n758 VGND.n757 0.0207703
R27009 VGND.n7332 VGND.n7331 0.0207703
R27010 VGND.n847 VGND.n846 0.0207703
R27011 VGND.n1538 VGND.n1537 0.0207703
R27012 VGND.n6959 VGND.n1539 0.0207703
R27013 VGND.n6190 VGND.n6189 0.0207703
R27014 VGND.n6098 VGND.n6097 0.0207703
R27015 VGND.n6770 VGND.n6769 0.0207703
R27016 VGND.n6266 VGND.n6265 0.0207703
R27017 VGND.n6465 VGND.n6464 0.0207703
R27018 VGND.n2234 VGND.n2233 0.0207703
R27019 VGND.n2168 VGND.n2167 0.0207703
R27020 VGND.n5214 VGND.n5213 0.0207703
R27021 VGND.n5221 VGND.n5215 0.0207703
R27022 VGND.n5187 VGND.n5186 0.0207703
R27023 VGND.n5793 VGND.n5188 0.0207703
R27024 VGND.n31 VGND.n30 0.0207703
R27025 VGND.n9097 VGND.n32 0.0207703
R27026 VGND.n5628 VGND.n5627 0.0207703
R27027 VGND.n2530 VGND.n2529 0.0207703
R27028 VGND.n9217 VGND.n9216 0.0207703
R27029 VGND.n9205 VGND.n9204 0.0207703
R27030 VGND.n5828 VGND.n5827 0.0207703
R27031 VGND.n5858 VGND.n5857 0.0207703
R27032 VGND.n3717 VGND.n3716 0.0204349
R27033 VGND.n1981 VGND.n1980 0.0204349
R27034 VGND.n1617 VGND.n1616 0.0202124
R27035 VGND.n6759 VGND.n6758 0.0202124
R27036 VGND.n1699 VGND.n1698 0.0202124
R27037 VGND.n1777 VGND.n1776 0.0202124
R27038 VGND.n1360 VGND.n1359 0.0202124
R27039 VGND.n1376 VGND.n1375 0.0202124
R27040 VGND.n7229 VGND.n7228 0.0202124
R27041 VGND.n1324 VGND.n1323 0.0202124
R27042 VGND.n4093 VGND.n4092 0.0202124
R27043 VGND.n4754 VGND.n4753 0.0202124
R27044 VGND.n4060 VGND.n4059 0.0202124
R27045 VGND.n4045 VGND.n4044 0.0202124
R27046 VGND.n4145 VGND.n4144 0.0202124
R27047 VGND.n4701 VGND.n4700 0.0202124
R27048 VGND.n4186 VGND.n4185 0.0202124
R27049 VGND.n4178 VGND.n4177 0.0202124
R27050 VGND.n1380 VGND.n1379 0.0202124
R27051 VGND.n1557 VGND.n1556 0.0202124
R27052 VGND.n4314 VGND.n4313 0.0202124
R27053 VGND.n4227 VGND.n4226 0.0202124
R27054 VGND.n2886 VGND.n2885 0.0202124
R27055 VGND.n2972 VGND.n2971 0.0202124
R27056 VGND.n3465 VGND.n3464 0.0202124
R27057 VGND.n2094 VGND.n2093 0.0202124
R27058 VGND.n49 VGND.n48 0.0202124
R27059 VGND.n9070 VGND.n9069 0.0202124
R27060 VGND.n2130 VGND.n2129 0.0202124
R27061 VGND.n2635 VGND.n2634 0.0202124
R27062 VGND.n3143 VGND.n3142 0.0202124
R27063 VGND.n2742 VGND.n2741 0.0202124
R27064 VGND.n3586 VGND.n3585 0.0202124
R27065 VGND.n3623 VGND.n3622 0.0202124
R27066 VGND.n9052 VGND.n9051 0.0202124
R27067 VGND.n70 VGND.n69 0.0202124
R27068 VGND.n106 VGND.n105 0.0202124
R27069 VGND.n120 VGND.n119 0.0202124
R27070 VGND.n264 VGND.n263 0.0202124
R27071 VGND.n277 VGND.n276 0.0202124
R27072 VGND.n3732 VGND.n3731 0.0202124
R27073 VGND.n1871 VGND.n1870 0.0202124
R27074 VGND.n8669 VGND.n8668 0.0202124
R27075 VGND.n8690 VGND.n8689 0.0202124
R27076 VGND.n137 VGND.n136 0.0202124
R27077 VGND.n8791 VGND.n8790 0.0202124
R27078 VGND.n281 VGND.n280 0.0202124
R27079 VGND.n8410 VGND.n8409 0.0202124
R27080 VGND.n2005 VGND.n2004 0.0202124
R27081 VGND.n1963 VGND.n1962 0.0202124
R27082 VGND.n463 VGND.n462 0.0202124
R27083 VGND.n8109 VGND.n8108 0.0202124
R27084 VGND.n544 VGND.n543 0.0202124
R27085 VGND.n558 VGND.n557 0.0202124
R27086 VGND.n723 VGND.n722 0.0202124
R27087 VGND.n7509 VGND.n7508 0.0202124
R27088 VGND.n8115 VGND.n8114 0.0202124
R27089 VGND.n8148 VGND.n8147 0.0202124
R27090 VGND.n422 VGND.n421 0.0202124
R27091 VGND.n8323 VGND.n8322 0.0202124
R27092 VGND.n584 VGND.n583 0.0202124
R27093 VGND.n7695 VGND.n7694 0.0202124
R27094 VGND.n7258 VGND.n7257 0.0202124
R27095 VGND.n1175 VGND.n1174 0.0202124
R27096 VGND.n768 VGND.n767 0.0202124
R27097 VGND.n858 VGND.n857 0.0202124
R27098 VGND.n6925 VGND.n1572 0.0202124
R27099 VGND.n6163 VGND.n6162 0.0202124
R27100 VGND.n6193 VGND.n6192 0.0202124
R27101 VGND.n1600 VGND.n1599 0.0202124
R27102 VGND.n6768 VGND.n6767 0.0202124
R27103 VGND.n6479 VGND.n6478 0.0202124
R27104 VGND.n5831 VGND.n5830 0.0202124
R27105 VGND.n5850 VGND.n5849 0.0202124
R27106 VGND.n2144 VGND.n2143 0.0202124
R27107 VGND.n2270 VGND.n2269 0.0202124
R27108 VGND.n6507 VGND.n6506 0.0202124
R27109 VGND.n5295 VGND.n5294 0.0202124
R27110 VGND.n5217 VGND.n5216 0.0202124
R27111 VGND.n5747 VGND.n5746 0.0202124
R27112 VGND.n5787 VGND.n5786 0.0202124
R27113 VGND.n2368 VGND.n2367 0.0202124
R27114 VGND.n41 VGND.n40 0.0202124
R27115 VGND.n5493 VGND.n5492 0.0202124
R27116 VGND.n5622 VGND.n5621 0.0202124
R27117 VGND.n2520 VGND.n2519 0.0202124
R27118 VGND.n2328 VGND.n2327 0.0202124
R27119 VGND.n3471 VGND.n3470 0.0202124
R27120 VGND.n9224 VGND.n9223 0.0202124
R27121 VGND.n1851 VGND.n1850 0.0202124
R27122 VGND.n5 VGND.n4 0.0200989
R27123 VGND.n5096 VGND.n5095 0.0200312
R27124 VGND.n7082 VGND.n7081 0.0200312
R27125 VGND VGND.n4108 0.0200312
R27126 VGND.n4330 VGND 0.0200312
R27127 VGND.n6981 VGND.n1473 0.0200312
R27128 VGND.n1469 VGND.n1468 0.0200312
R27129 VGND.n3285 VGND 0.0200312
R27130 VGND VGND.n3233 0.0200312
R27131 VGND VGND.n2846 0.0200312
R27132 VGND.n2895 VGND.n2894 0.0200312
R27133 VGND.n2986 VGND.n2985 0.0200312
R27134 VGND.n8883 VGND 0.0200312
R27135 VGND VGND.n8923 0.0200312
R27136 VGND.n9023 VGND 0.0200312
R27137 VGND.n9024 VGND.n9023 0.0200312
R27138 VGND.n3199 VGND.n3198 0.0200312
R27139 VGND.n3194 VGND.n3193 0.0200312
R27140 VGND.n3852 VGND 0.0200312
R27141 VGND.n8562 VGND.n8561 0.0200312
R27142 VGND.n304 VGND.n303 0.0200312
R27143 VGND.n8541 VGND.n8540 0.0200312
R27144 VGND.n7982 VGND.n7981 0.0200312
R27145 VGND.n8428 VGND.n8427 0.0200312
R27146 VGND.n8423 VGND.n8422 0.0200312
R27147 VGND VGND.n701 0.0200312
R27148 VGND.n8133 VGND 0.0200312
R27149 VGND.n8333 VGND.n8332 0.0200312
R27150 VGND.n325 VGND.n324 0.0200312
R27151 VGND VGND.n7477 0.0200312
R27152 VGND.n7309 VGND.n7308 0.0200312
R27153 VGND.n979 VGND.n978 0.0200312
R27154 VGND.n1685 VGND 0.0200312
R27155 VGND.n6470 VGND.n6469 0.0200312
R27156 VGND.n6802 VGND.n6801 0.0200312
R27157 VGND.n6974 VGND.n6973 0.0200312
R27158 VGND.n6969 VGND.n6968 0.0200312
R27159 VGND VGND.n1729 0.0200312
R27160 VGND.n5313 VGND.n5312 0.0200312
R27161 VGND.n5333 VGND.n5332 0.0200312
R27162 VGND VGND.n1821 0.0200312
R27163 VGND.n5599 VGND.n5598 0.0200312
R27164 VGND.n5809 VGND.n5808 0.0200312
R27165 VGND.n5804 VGND.n5803 0.0200312
R27166 VGND.n5142 VGND 0.0200312
R27167 VGND.n2481 VGND 0.0200312
R27168 VGND.n9176 VGND.n9175 0.0200312
R27169 VGND.n9171 VGND.n9170 0.0200312
R27170 VGND.n3235 VGND 0.0199818
R27171 VGND.n4864 VGND.n4863 0.0195896
R27172 VGND.n4716 VGND.n4711 0.0195896
R27173 VGND.n3578 VGND.n3577 0.0195896
R27174 VGND.n3724 VGND.n3723 0.0195896
R27175 VGND.n3842 VGND.n3841 0.0195896
R27176 VGND.n1971 VGND.n1969 0.0195896
R27177 VGND.n7561 VGND.n7560 0.0195896
R27178 VGND.n9211 VGND.n9210 0.0195896
R27179 VGND.n5972 VGND.n5969 0.0193669
R27180 VGND.n1784 VGND.n1783 0.0190811
R27181 VGND.n1795 VGND.n1794 0.0190811
R27182 VGND.n6001 VGND.n6000 0.0190811
R27183 VGND.n5987 VGND.n5986 0.0190811
R27184 VGND.n6755 VGND.n6754 0.0190811
R27185 VGND.n1749 VGND.n1748 0.0190811
R27186 VGND.n1703 VGND.n1702 0.0190811
R27187 VGND.n6072 VGND.n6071 0.0190811
R27188 VGND.n6079 VGND.n6078 0.0190811
R27189 VGND.n6501 VGND.n6500 0.0190811
R27190 VGND.n6528 VGND.n6527 0.0190811
R27191 VGND.n1374 VGND.n1373 0.0190811
R27192 VGND.n7244 VGND.n7243 0.0190811
R27193 VGND.n7233 VGND.n7232 0.0190811
R27194 VGND.n4818 VGND.n4817 0.0190811
R27195 VGND.n4806 VGND.n4805 0.0190811
R27196 VGND.n4843 VGND.n4842 0.0190811
R27197 VGND.n4829 VGND.n4828 0.0190811
R27198 VGND.n4053 VGND.n4052 0.0190811
R27199 VGND.n4064 VGND.n4063 0.0190811
R27200 VGND.n4992 VGND.n4074 0.0190811
R27201 VGND.n4138 VGND.n4137 0.0190811
R27202 VGND.n4157 VGND.n4156 0.0190811
R27203 VGND.n4733 VGND.n4147 0.0190811
R27204 VGND.n4740 VGND.n4739 0.0190811
R27205 VGND.n4189 VGND.n4188 0.0190811
R27206 VGND.n4199 VGND.n4198 0.0190811
R27207 VGND.n1455 VGND.n1454 0.0190811
R27208 VGND.n4359 VGND.n4358 0.0190811
R27209 VGND.n4352 VGND.n4311 0.0190811
R27210 VGND.n4341 VGND.n4317 0.0190811
R27211 VGND.n2970 VGND.n2969 0.0190811
R27212 VGND.n2087 VGND.n2086 0.0190811
R27213 VGND.n3462 VGND.n3454 0.0190811
R27214 VGND.n3559 VGND.n3558 0.0190811
R27215 VGND.n3545 VGND.n3544 0.0190811
R27216 VGND.n3231 VGND.n50 0.0190811
R27217 VGND.n2769 VGND.n2768 0.0190811
R27218 VGND.n3342 VGND.n3341 0.0190811
R27219 VGND.n2134 VGND.n2133 0.0190811
R27220 VGND.n3356 VGND.n3355 0.0190811
R27221 VGND.n2740 VGND.n2739 0.0190811
R27222 VGND.n3616 VGND.n3615 0.0190811
R27223 VGND.n3590 VGND.n3589 0.0190811
R27224 VGND.n3594 VGND.n3593 0.0190811
R27225 VGND.n3601 VGND.n3600 0.0190811
R27226 VGND.n9055 VGND.n9054 0.0190811
R27227 VGND.n66 VGND.n65 0.0190811
R27228 VGND.n8820 VGND.n8819 0.0190811
R27229 VGND.n110 VGND.n109 0.0190811
R27230 VGND.n8834 VGND.n8833 0.0190811
R27231 VGND.n275 VGND.n274 0.0190811
R27232 VGND.n3762 VGND.n3761 0.0190811
R27233 VGND.n3736 VGND.n3735 0.0190811
R27234 VGND.n3740 VGND.n3739 0.0190811
R27235 VGND.n3747 VGND.n3746 0.0190811
R27236 VGND.n8667 VGND.n8666 0.0190811
R27237 VGND.n8685 VGND.n8684 0.0190811
R27238 VGND.n3895 VGND.n3889 0.0190811
R27239 VGND.n141 VGND.n140 0.0190811
R27240 VGND.n8802 VGND.n151 0.0190811
R27241 VGND.n8408 VGND.n8407 0.0190811
R27242 VGND.n1998 VGND.n1997 0.0190811
R27243 VGND.n2009 VGND.n2008 0.0190811
R27244 VGND.n2013 VGND.n2012 0.0190811
R27245 VGND.n2020 VGND.n2019 0.0190811
R27246 VGND.n466 VGND.n465 0.0190811
R27247 VGND.n8105 VGND.n8104 0.0190811
R27248 VGND.n7724 VGND.n7723 0.0190811
R27249 VGND.n548 VGND.n547 0.0190811
R27250 VGND.n7738 VGND.n7737 0.0190811
R27251 VGND.n721 VGND.n720 0.0190811
R27252 VGND.n727 VGND.n726 0.0190811
R27253 VGND.n731 VGND.n730 0.0190811
R27254 VGND.n738 VGND.n737 0.0190811
R27255 VGND.n8138 VGND.n8128 0.0190811
R27256 VGND.n8119 VGND.n8118 0.0190811
R27257 VGND.n322 VGND.n321 0.0190811
R27258 VGND.n579 VGND.n578 0.0190811
R27259 VGND.n588 VGND.n587 0.0190811
R27260 VGND.n7706 VGND.n598 0.0190811
R27261 VGND.n7265 VGND.n7264 0.0190811
R27262 VGND.n7286 VGND.n7285 0.0190811
R27263 VGND.n902 VGND.n901 0.0190811
R27264 VGND.n784 VGND.n783 0.0190811
R27265 VGND.n7446 VGND.n774 0.0190811
R27266 VGND.n760 VGND.n759 0.0190811
R27267 VGND.n7332 VGND.n7330 0.0190811
R27268 VGND.n835 VGND.n834 0.0190811
R27269 VGND.n881 VGND.n880 0.0190811
R27270 VGND.n1539 VGND.n1538 0.0190811
R27271 VGND.n6102 VGND.n6101 0.0190811
R27272 VGND.n6113 VGND.n6105 0.0190811
R27273 VGND.n6170 VGND.n6169 0.0190811
R27274 VGND.n6189 VGND.n6099 0.0190811
R27275 VGND.n1606 VGND.n1605 0.0190811
R27276 VGND.n6776 VGND.n6775 0.0190811
R27277 VGND.n6269 VGND.n6266 0.0190811
R27278 VGND.n6485 VGND.n6484 0.0190811
R27279 VGND.n6472 VGND.n1669 0.0190811
R27280 VGND.n2238 VGND.n2234 0.0190811
R27281 VGND.n2153 VGND.n2152 0.0190811
R27282 VGND.n5215 VGND.n5214 0.0190811
R27283 VGND.n5188 VGND.n5187 0.0190811
R27284 VGND.n32 VGND.n31 0.0190811
R27285 VGND.n5479 VGND.n5478 0.0190811
R27286 VGND.n5476 VGND.n5475 0.0190811
R27287 VGND.n2528 VGND.n2527 0.0190811
R27288 VGND.n3480 VGND.n3479 0.0190811
R27289 VGND.n3528 VGND.n3483 0.0190811
R27290 VGND.n3530 VGND.n1 0.0190811
R27291 VGND.n9216 VGND.n2 0.0190811
R27292 VGND.n5829 VGND.n5828 0.0190811
R27293 VGND.n5837 VGND.n5836 0.0190811
R27294 VGND.n5865 VGND.n5864 0.0190811
R27295 VGND.n2776 VGND 0.0188432
R27296 VGND.n4801 VGND 0.0187292
R27297 VGND.n4811 VGND.n4810 0.0187292
R27298 VGND.n4981 VGND.n4980 0.0187292
R27299 VGND.n7212 VGND.n7211 0.0187292
R27300 VGND.n7202 VGND.n7198 0.0187292
R27301 VGND.n7196 VGND 0.0187292
R27302 VGND.n4152 VGND.n4148 0.0187292
R27303 VGND.n4334 VGND.n4332 0.0187292
R27304 VGND.n4503 VGND.n4502 0.0187292
R27305 VGND.n4519 VGND.n4517 0.0187292
R27306 VGND.n4520 VGND 0.0187292
R27307 VGND.n3458 VGND.n3455 0.0187292
R27308 VGND.n3360 VGND.n3358 0.0187292
R27309 VGND.n3233 VGND 0.0187292
R27310 VGND.n9077 VGND.n52 0.0187292
R27311 VGND.n2780 VGND.n2778 0.0187292
R27312 VGND.n3708 VGND.n3704 0.0187292
R27313 VGND.n8838 VGND.n8836 0.0187292
R27314 VGND.n9032 VGND.n9031 0.0187292
R27315 VGND.n3039 VGND.n76 0.0187292
R27316 VGND VGND.n3040 0.0187292
R27317 VGND.n3818 VGND.n3816 0.0187292
R27318 VGND VGND.n8656 0.0187292
R27319 VGND.n8679 VGND.n8664 0.0187292
R27320 VGND.n8651 VGND.n8650 0.0187292
R27321 VGND VGND.n1917 0.0187292
R27322 VGND.n1991 VGND.n1990 0.0187292
R27323 VGND.n7743 VGND.n7740 0.0187292
R27324 VGND.n8079 VGND.n8078 0.0187292
R27325 VGND.n8070 VGND.n8067 0.0187292
R27326 VGND.n8065 VGND 0.0187292
R27327 VGND.n7537 VGND.n7533 0.0187292
R27328 VGND.n7611 VGND.n599 0.0187292
R27329 VGND VGND.n8133 0.0187292
R27330 VGND.n8192 VGND.n8191 0.0187292
R27331 VGND.n778 VGND.n776 0.0187292
R27332 VGND.n876 VGND.n874 0.0187292
R27333 VGND.n1304 VGND.n1303 0.0187292
R27334 VGND.n1297 VGND.n1296 0.0187292
R27335 VGND.n6110 VGND.n6107 0.0187292
R27336 VGND.n6810 VGND.n6809 0.0187292
R27337 VGND.n6824 VGND.n6822 0.0187292
R27338 VGND VGND.n6825 0.0187292
R27339 VGND.n1761 VGND.n1759 0.0187292
R27340 VGND.n6552 VGND.n6550 0.0187292
R27341 VGND.n5353 VGND.n5352 0.0187292
R27342 VGND.n5370 VGND.n5369 0.0187292
R27343 VGND VGND.n5372 0.0187292
R27344 VGND.n1840 VGND.n1837 0.0187292
R27345 VGND.n5871 VGND.n5869 0.0187292
R27346 VGND.n5643 VGND.n5641 0.0187292
R27347 VGND.n3524 VGND.n3521 0.0187292
R27348 VGND.n2266 VGND.n2265 0.0187292
R27349 VGND.n2503 VGND.n2502 0.0187292
R27350 VGND.n2493 VGND.n2492 0.0187292
R27351 VGND.n2487 VGND 0.0187292
R27352 VGND.n803 VGND 0.0179232
R27353 VGND.n4008 VGND.n4006 0.0174271
R27354 VGND.n4213 VGND.n4212 0.0174271
R27355 VGND.n9022 VGND.n9020 0.0174271
R27356 VGND.n8655 VGND.n8653 0.0174271
R27357 VGND.n7918 VGND.n7917 0.0174271
R27358 VGND.n8131 VGND.n8129 0.0174271
R27359 VGND.n1130 VGND.n1129 0.0174271
R27360 VGND.n6800 VGND.n6798 0.0174271
R27361 VGND.n6723 VGND.n6722 0.0174271
R27362 VGND.n5602 VGND.n5601 0.0174271
R27363 VGND.n2317 VGND.n2316 0.0174271
R27364 VGND.n1796 VGND.n1795 0.0173919
R27365 VGND.n1704 VGND.n1703 0.0173919
R27366 VGND.n6527 VGND.n6526 0.0173919
R27367 VGND.n1357 VGND.n1356 0.0173919
R27368 VGND.n4806 VGND.n4091 0.0173919
R27369 VGND.n4063 VGND.n4062 0.0173919
R27370 VGND.n4157 VGND.n4146 0.0173919
R27371 VGND.n1387 VGND.n1386 0.0173919
R27372 VGND.n4311 VGND.n4310 0.0173919
R27373 VGND.n2883 VGND.n2882 0.0173919
R27374 VGND.n3463 VGND.n3462 0.0173919
R27375 VGND.n2133 VGND.n2132 0.0173919
R27376 VGND.n3136 VGND.n3135 0.0173919
R27377 VGND.n3591 VGND.n3590 0.0173919
R27378 VGND.n109 VGND.n108 0.0173919
R27379 VGND.n261 VGND.n260 0.0173919
R27380 VGND.n3737 VGND.n3736 0.0173919
R27381 VGND.n140 VGND.n139 0.0173919
R27382 VGND.n298 VGND.n297 0.0173919
R27383 VGND.n2010 VGND.n2009 0.0173919
R27384 VGND.n547 VGND.n546 0.0173919
R27385 VGND.n728 VGND.n727 0.0173919
R27386 VGND.n416 VGND.n415 0.0173919
R27387 VGND.n587 VGND.n586 0.0173919
R27388 VGND.n1167 VGND.n1166 0.0173919
R27389 VGND.n784 VGND.n773 0.0173919
R27390 VGND.n834 VGND.n833 0.0173919
R27391 VGND.n1577 VGND.n1576 0.0173919
R27392 VGND.n6114 VGND.n6113 0.0173919
R27393 VGND.n6484 VGND.n6483 0.0173919
R27394 VGND.n2152 VGND.n2151 0.0173919
R27395 VGND.n5303 VGND.n5302 0.0173919
R27396 VGND.n5466 VGND.n5465 0.0173919
R27397 VGND.n2361 VGND.n2360 0.0173919
R27398 VGND.n3529 VGND.n3528 0.0173919
R27399 VGND.n7985 VGND.n7983 0.017391
R27400 VGND.n5454 VGND.n5196 0.017391
R27401 VGND.n9168 VGND.n22 0.0172667
R27402 VGND.n3010 VGND.n3009 0.0172634
R27403 VGND.n868 VGND.n867 0.0172616
R27404 VGND.n1678 VGND.n1677 0.0172616
R27405 VGND.n6734 VGND.n1618 0.0168788
R27406 VGND.n5344 VGND.n5343 0.0168788
R27407 VGND.n1752 VGND.n1751 0.0168788
R27408 VGND.n6013 VGND.n1778 0.0168788
R27409 VGND.n6996 VGND.n6992 0.0168788
R27410 VGND.n7000 VGND.n1377 0.0168788
R27411 VGND.n4001 VGND.n4000 0.0168788
R27412 VGND.n7225 VGND.n1325 0.0168788
R27413 VGND.n4821 VGND.n4820 0.0168788
R27414 VGND.n4762 VGND.n4755 0.0168788
R27415 VGND.n4054 VGND.n4048 0.0168788
R27416 VGND.n5004 VGND.n4046 0.0168788
R27417 VGND.n4141 VGND.n4140 0.0168788
R27418 VGND.n4708 VGND.n4702 0.0168788
R27419 VGND.n4487 VGND.n4486 0.0168788
R27420 VGND.n4492 VGND.n4179 0.0168788
R27421 VGND.n4584 VGND.n4583 0.0168788
R27422 VGND.n1458 VGND.n1456 0.0168788
R27423 VGND.n4361 VGND.n4360 0.0168788
R27424 VGND.n4369 VGND.n4228 0.0168788
R27425 VGND.n3017 VGND.n2746 0.0168788
R27426 VGND.n2975 VGND.n2973 0.0168788
R27427 VGND.n2090 VGND.n2089 0.0168788
R27428 VGND.n3581 VGND.n2095 0.0168788
R27429 VGND.n3241 VGND.n3240 0.0168788
R27430 VGND.n2762 VGND.n2760 0.0168788
R27431 VGND.n3343 VGND.n3337 0.0168788
R27432 VGND.n3333 VGND.n2636 0.0168788
R27433 VGND.n3178 VGND.n3025 0.0168788
R27434 VGND.n3182 VGND.n2743 0.0168788
R27435 VGND.n3619 VGND.n3618 0.0168788
R27436 VGND.n3727 VGND.n3624 0.0168788
R27437 VGND.n9011 VGND.n9010 0.0168788
R27438 VGND.n9048 VGND.n73 0.0168788
R27439 VGND.n8821 VGND.n8815 0.0168788
R27440 VGND.n133 VGND.n121 0.0168788
R27441 VGND.n8444 VGND.n8440 0.0168788
R27442 VGND.n8448 VGND.n278 0.0168788
R27443 VGND.n3765 VGND.n3764 0.0168788
R27444 VGND.n3770 VGND.n1872 0.0168788
R27445 VGND.n8714 VGND.n8713 0.0168788
R27446 VGND.n8709 VGND.n204 0.0168788
R27447 VGND.n3894 VGND.n3893 0.0168788
R27448 VGND.n8794 VGND.n8792 0.0168788
R27449 VGND.n7976 VGND.n7975 0.0168788
R27450 VGND.n8413 VGND.n8411 0.0168788
R27451 VGND.n2001 VGND.n2000 0.0168788
R27452 VGND.n1966 VGND.n1964 0.0168788
R27453 VGND.n7911 VGND.n7910 0.0168788
R27454 VGND.n8094 VGND.n477 0.0168788
R27455 VGND.n7725 VGND.n7719 0.0168788
R27456 VGND.n570 VGND.n559 0.0168788
R27457 VGND.n7522 VGND.n7521 0.0168788
R27458 VGND.n7517 VGND.n7510 0.0168788
R27459 VGND.n8214 VGND.n8213 0.0168788
R27460 VGND.n8151 VGND.n8149 0.0168788
R27461 VGND.n8318 VGND.n8317 0.0168788
R27462 VGND.n411 VGND.n319 0.0168788
R27463 VGND.n580 VGND.n574 0.0168788
R27464 VGND.n7698 VGND.n7696 0.0168788
R27465 VGND.n5833 VGND.n5832 0.0168788
R27466 VGND.n5855 VGND.n5821 0.0168788
R27467 VGND.n2237 VGND.n2236 0.0168788
R27468 VGND.n2629 VGND.n2164 0.0168788
R27469 VGND.n6504 VGND.n6503 0.0168788
R27470 VGND.n6521 VGND.n6508 0.0168788
R27471 VGND.n5461 VGND.n5194 0.0168788
R27472 VGND.n5220 VGND.n5218 0.0168788
R27473 VGND.n5749 VGND.n5748 0.0168788
R27474 VGND.n5792 VGND.n5189 0.0168788
R27475 VGND.n2396 VGND.n2395 0.0168788
R27476 VGND.n9096 VGND.n42 0.0168788
R27477 VGND.n5612 VGND.n5494 0.0168788
R27478 VGND.n5617 VGND.n5614 0.0168788
R27479 VGND.n2540 VGND.n2539 0.0168788
R27480 VGND.n2516 VGND.n2329 0.0168788
R27481 VGND.n3469 VGND.n3468 0.0168788
R27482 VGND.n9222 VGND.n9221 0.0168788
R27483 VGND.n1788 VGND.n1787 0.0168788
R27484 VGND.n1853 VGND.n1852 0.0168788
R27485 VGND.n8420 VGND.n8417 0.0166396
R27486 VGND.n5335 VGND.n5290 0.0166396
R27487 VGND.n9169 VGND.n9168 0.016628
R27488 VGND.n3011 VGND.n3010 0.0166244
R27489 VGND.n867 VGND.n865 0.0166226
R27490 VGND.n1677 VGND.n1676 0.0166226
R27491 VGND.n6017 VGND 0.0166211
R27492 VGND.n7986 VGND.n7985 0.0164962
R27493 VGND.n5455 VGND.n5454 0.0164962
R27494 VGND.n4963 VGND.n4955 0.016464
R27495 VGND.n4304 VGND.n4300 0.016464
R27496 VGND.n3382 VGND.n3381 0.016464
R27497 VGND.n8860 VGND.n8859 0.016464
R27498 VGND.n3919 VGND.n3918 0.016464
R27499 VGND.n7760 VGND.n536 0.016464
R27500 VGND.n7634 VGND.n7633 0.016464
R27501 VGND.n7341 VGND.n7340 0.016464
R27502 VGND.n6277 VGND.n6276 0.016464
R27503 VGND.n6575 VGND.n6574 0.016464
R27504 VGND.n5892 VGND.n5891 0.016464
R27505 VGND.n2244 VGND.n2241 0.016464
R27506 VGND.n5335 VGND.n5334 0.0162568
R27507 VGND.n8421 VGND.n8420 0.0162568
R27508 VGND.n4856 VGND.n4855 0.016125
R27509 VGND.n4859 VGND.n4858 0.016125
R27510 VGND VGND.n4989 0.016125
R27511 VGND.n5011 VGND.n5010 0.016125
R27512 VGND.n7209 VGND.n7207 0.016125
R27513 VGND.n7213 VGND.n7212 0.016125
R27514 VGND.n7079 VGND.n7075 0.016125
R27515 VGND.n7075 VGND 0.016125
R27516 VGND.n4718 VGND.n4717 0.016125
R27517 VGND.n4339 VGND 0.016125
R27518 VGND.n4376 VGND.n4375 0.016125
R27519 VGND.n4500 VGND.n4498 0.016125
R27520 VGND.n4504 VGND.n4503 0.016125
R27521 VGND.n1466 VGND.n1463 0.016125
R27522 VGND.n3567 VGND.n3566 0.016125
R27523 VGND.n3570 VGND.n3569 0.016125
R27524 VGND.n2642 VGND 0.016125
R27525 VGND.n3329 VGND.n3328 0.016125
R27526 VGND.n3228 VGND.n3226 0.016125
R27527 VGND.n2983 VGND.n2980 0.016125
R27528 VGND.n3719 VGND.n3718 0.016125
R27529 VGND.n3722 VGND.n3721 0.016125
R27530 VGND.n127 VGND 0.016125
R27531 VGND.n129 VGND.n82 0.016125
R27532 VGND.n9029 VGND.n9027 0.016125
R27533 VGND.n9033 VGND.n9032 0.016125
R27534 VGND.n3191 VGND.n3186 0.016125
R27535 VGND.n3834 VGND.n3833 0.016125
R27536 VGND.n3837 VGND.n3836 0.016125
R27537 VGND.n8800 VGND 0.016125
R27538 VGND.n8787 VGND.n8786 0.016125
R27539 VGND.n8662 VGND.n8660 0.016125
R27540 VGND.n8538 VGND.n8530 0.016125
R27541 VGND VGND.n8529 0.016125
R27542 VGND.n1976 VGND.n1975 0.016125
R27543 VGND.n1973 VGND.n1972 0.016125
R27544 VGND.n565 VGND 0.016125
R27545 VGND.n7815 VGND.n507 0.016125
R27546 VGND.n8076 VGND.n8074 0.016125
R27547 VGND.n8080 VGND.n8079 0.016125
R27548 VGND.n7529 VGND 0.016125
R27549 VGND.n7555 VGND.n7554 0.016125
R27550 VGND.n7558 VGND.n7557 0.016125
R27551 VGND VGND.n7703 0.016125
R27552 VGND.n7691 VGND.n7690 0.016125
R27553 VGND.n8203 VGND 0.016125
R27554 VGND.n8201 VGND.n8200 0.016125
R27555 VGND.n331 VGND.n330 0.016125
R27556 VGND VGND.n331 0.016125
R27557 VGND.n7434 VGND.n7432 0.016125
R27558 VGND.n7430 VGND.n7429 0.016125
R27559 VGND.n878 VGND 0.016125
R27560 VGND.n7321 VGND.n7320 0.016125
R27561 VGND.n1302 VGND.n1301 0.016125
R27562 VGND.n1305 VGND.n1304 0.016125
R27563 VGND.n986 VGND.n985 0.016125
R27564 VGND.n6186 VGND.n6185 0.016125
R27565 VGND.n6458 VGND.n6457 0.016125
R27566 VGND.n6807 VGND.n6805 0.016125
R27567 VGND.n6811 VGND.n6810 0.016125
R27568 VGND.n6966 VGND.n6963 0.016125
R27569 VGND VGND.n1705 0.016125
R27570 VGND.n6061 VGND.n6059 0.016125
R27571 VGND.n6057 VGND.n6056 0.016125
R27572 VGND.n6515 VGND 0.016125
R27573 VGND.n6517 VGND.n1636 0.016125
R27574 VGND.n5351 VGND.n5350 0.016125
R27575 VGND.n5354 VGND.n5353 0.016125
R27576 VGND VGND.n5116 0.016125
R27577 VGND.n5818 VGND.n5817 0.016125
R27578 VGND.n5596 VGND.n5592 0.016125
R27579 VGND.n5590 VGND 0.016125
R27580 VGND.n5630 VGND.n5629 0.016125
R27581 VGND.n5801 VGND.n5796 0.016125
R27582 VGND.n2625 VGND.n2624 0.016125
R27583 VGND.n2500 VGND.n2498 0.016125
R27584 VGND.n2504 VGND.n2503 0.016125
R27585 VGND.n6754 VGND.n6753 0.0157027
R27586 VGND.n2768 VGND.n2767 0.0157027
R27587 VGND.n65 VGND.n64 0.0157027
R27588 VGND.n8684 VGND.n8683 0.0157027
R27589 VGND.n8104 VGND.n8103 0.0157027
R27590 VGND.n7285 VGND.n7284 0.0157027
R27591 VGND.n6775 VGND.n6774 0.0157027
R27592 VGND.n5475 VGND.n5474 0.0157027
R27593 VGND.n2332 VGND.n2331 0.0157027
R27594 VGND.n4808 VGND.n4807 0.0148229
R27595 VGND.n4844 VGND 0.0148229
R27596 VGND.n4857 VGND.n4856 0.0148229
R27597 VGND.n4970 VGND.n4969 0.0148229
R27598 VGND.n4991 VGND.n4990 0.0148229
R27599 VGND.n5009 VGND.n4042 0.0148229
R27600 VGND.n7204 VGND.n7203 0.0148229
R27601 VGND.n7217 VGND.n7216 0.0148229
R27602 VGND.n7096 VGND 0.0148229
R27603 VGND.n7080 VGND.n7079 0.0148229
R27604 VGND.n4158 VGND.n4153 0.0148229
R27605 VGND VGND.n4732 0.0148229
R27606 VGND.n4720 VGND.n4719 0.0148229
R27607 VGND.n4354 VGND.n4353 0.0148229
R27608 VGND.n4340 VGND.n4339 0.0148229
R27609 VGND.n4374 VGND.n4224 0.0148229
R27610 VGND.n4496 VGND.n4495 0.0148229
R27611 VGND.n4508 VGND.n4507 0.0148229
R27612 VGND.n4569 VGND 0.0148229
R27613 VGND.n1467 VGND.n1466 0.0148229
R27614 VGND.n3461 VGND.n3459 0.0148229
R27615 VGND.n3560 VGND 0.0148229
R27616 VGND.n3568 VGND.n3567 0.0148229
R27617 VGND.n3374 VGND.n3373 0.0148229
R27618 VGND.n3357 VGND.n2126 0.0148229
R27619 VGND.n3330 VGND.n2643 0.0148229
R27620 VGND.n3230 VGND.n3229 0.0148229
R27621 VGND.n2771 VGND.n2770 0.0148229
R27622 VGND.n3005 VGND 0.0148229
R27623 VGND.n2984 VGND.n2983 0.0148229
R27624 VGND.n3710 VGND.n3709 0.0148229
R27625 VGND.n3713 VGND.n3712 0.0148229
R27626 VGND.n3720 VGND.n3719 0.0148229
R27627 VGND.n8852 VGND.n8851 0.0148229
R27628 VGND.n8835 VGND.n102 0.0148229
R27629 VGND.n130 VGND.n128 0.0148229
R27630 VGND.n9025 VGND.n9024 0.0148229
R27631 VGND.n9037 VGND.n9036 0.0148229
R27632 VGND.n3160 VGND 0.0148229
R27633 VGND.n3192 VGND.n3191 0.0148229
R27634 VGND.n3820 VGND.n3819 0.0148229
R27635 VGND.n3823 VGND.n3822 0.0148229
R27636 VGND.n3835 VGND.n3834 0.0148229
R27637 VGND.n3911 VGND.n3910 0.0148229
R27638 VGND.n8801 VGND.n8800 0.0148229
R27639 VGND.n8788 VGND.n156 0.0148229
R27640 VGND.n8658 VGND.n8657 0.0148229
R27641 VGND.n8698 VGND.n8697 0.0148229
R27642 VGND.n8559 VGND 0.0148229
R27643 VGND.n8539 VGND.n8538 0.0148229
R27644 VGND.n1988 VGND.n1987 0.0148229
R27645 VGND.n1985 VGND.n1984 0.0148229
R27646 VGND.n1975 VGND.n1974 0.0148229
R27647 VGND.n7754 VGND.n7753 0.0148229
R27648 VGND.n7739 VGND.n540 0.0148229
R27649 VGND.n567 VGND.n566 0.0148229
R27650 VGND.n8072 VGND.n8071 0.0148229
R27651 VGND.n8084 VGND.n8083 0.0148229
R27652 VGND.n7979 VGND 0.0148229
R27653 VGND.n7539 VGND.n7538 0.0148229
R27654 VGND.n7542 VGND.n7541 0.0148229
R27655 VGND.n7556 VGND.n7555 0.0148229
R27656 VGND.n7626 VGND.n7625 0.0148229
R27657 VGND.n7705 VGND.n7704 0.0148229
R27658 VGND.n7692 VGND.n605 0.0148229
R27659 VGND.n8137 VGND.n8134 0.0148229
R27660 VGND.n8197 VGND.n8196 0.0148229
R27661 VGND.n429 VGND 0.0148229
R27662 VGND.n330 VGND.n326 0.0148229
R27663 VGND.n785 VGND.n779 0.0148229
R27664 VGND VGND.n7445 0.0148229
R27665 VGND.n7432 VGND.n7431 0.0148229
R27666 VGND.n864 VGND.n863 0.0148229
R27667 VGND.n879 VGND.n878 0.0148229
R27668 VGND.n7322 VGND.n884 0.0148229
R27669 VGND.n1299 VGND.n1298 0.0148229
R27670 VGND.n1309 VGND.n1308 0.0148229
R27671 VGND.n1183 VGND 0.0148229
R27672 VGND.n985 VGND.n980 0.0148229
R27673 VGND.n6112 VGND.n6111 0.0148229
R27674 VGND.n6171 VGND 0.0148229
R27675 VGND.n6188 VGND.n6187 0.0148229
R27676 VGND.n1675 VGND.n1674 0.0148229
R27677 VGND.n6471 VGND.n6470 0.0148229
R27678 VGND.n6468 VGND.n6467 0.0148229
R27679 VGND.n6803 VGND.n6802 0.0148229
R27680 VGND.n6815 VGND.n6814 0.0148229
R27681 VGND VGND.n6944 0.0148229
R27682 VGND.n6967 VGND.n6966 0.0148229
R27683 VGND.n1763 VGND.n1762 0.0148229
R27684 VGND.n1766 VGND.n1765 0.0148229
R27685 VGND.n6059 VGND.n6058 0.0148229
R27686 VGND.n6568 VGND.n6567 0.0148229
R27687 VGND.n6548 VGND.n1654 0.0148229
R27688 VGND.n6518 VGND.n6516 0.0148229
R27689 VGND.n5348 VGND.n5347 0.0148229
R27690 VGND.n5358 VGND.n5357 0.0148229
R27691 VGND.n1842 VGND.n1841 0.0148229
R27692 VGND.n1845 VGND.n1844 0.0148229
R27693 VGND.n5988 VGND.n5975 0.0148229
R27694 VGND.n5885 VGND.n5884 0.0148229
R27695 VGND.n5867 VGND.n5116 0.0148229
R27696 VGND.n5861 VGND.n5860 0.0148229
R27697 VGND.n5598 VGND.n5597 0.0148229
R27698 VGND.n5634 VGND.n5633 0.0148229
R27699 VGND VGND.n5765 0.0148229
R27700 VGND.n5802 VGND.n5801 0.0148229
R27701 VGND.n3527 VGND.n3525 0.0148229
R27702 VGND VGND.n9232 0.0148229
R27703 VGND.n9215 VGND.n9214 0.0148229
R27704 VGND.n2251 VGND.n2250 0.0148229
R27705 VGND.n2278 VGND.n2277 0.0148229
R27706 VGND.n2626 VGND.n2283 0.0148229
R27707 VGND.n2495 VGND.n2494 0.0148229
R27708 VGND.n2508 VGND.n2507 0.0148229
R27709 VGND.n2379 VGND 0.0148229
R27710 VGND.n6744 VGND.n6743 0.0145155
R27711 VGND.n6745 VGND.n6744 0.0145155
R27712 VGND.n6086 VGND.n6085 0.0145155
R27713 VGND.n6085 VGND.n6084 0.0145155
R27714 VGND.n7091 VGND.n7090 0.0145155
R27715 VGND.n7090 VGND.n7089 0.0145155
R27716 VGND.n7240 VGND.n7239 0.0145155
R27717 VGND.n7239 VGND.n7238 0.0145155
R27718 VGND.n4836 VGND.n4835 0.0145155
R27719 VGND.n4835 VGND.n4834 0.0145155
R27720 VGND.n4998 VGND.n4997 0.0145155
R27721 VGND.n4997 VGND.n4996 0.0145155
R27722 VGND.n4747 VGND.n4746 0.0145155
R27723 VGND.n4746 VGND.n4745 0.0145155
R27724 VGND.n4206 VGND.n4205 0.0145155
R27725 VGND.n4205 VGND.n4204 0.0145155
R27726 VGND.n1382 VGND.n1381 0.0145155
R27727 VGND.n4347 VGND.n4346 0.0145155
R27728 VGND.n4346 VGND.n4345 0.0145155
R27729 VGND.n3000 VGND.n2999 0.0145155
R27730 VGND.n2999 VGND.n2998 0.0145155
R27731 VGND.n3552 VGND.n3551 0.0145155
R27732 VGND.n3551 VGND.n3550 0.0145155
R27733 VGND.n9084 VGND.n9083 0.0145155
R27734 VGND.n3350 VGND.n3349 0.0145155
R27735 VGND.n3351 VGND.n3350 0.0145155
R27736 VGND.n3155 VGND.n3154 0.0145155
R27737 VGND.n3154 VGND.n3153 0.0145155
R27738 VGND.n3608 VGND.n3607 0.0145155
R27739 VGND.n3607 VGND.n3606 0.0145155
R27740 VGND.n9062 VGND.n9061 0.0145155
R27741 VGND.n8828 VGND.n8827 0.0145155
R27742 VGND.n8829 VGND.n8828 0.0145155
R27743 VGND.n8550 VGND.n8549 0.0145155
R27744 VGND.n8549 VGND.n8548 0.0145155
R27745 VGND.n3754 VGND.n3753 0.0145155
R27746 VGND.n3753 VGND.n3752 0.0145155
R27747 VGND.n8671 VGND.n8670 0.0145155
R27748 VGND.n8808 VGND.n8807 0.0145155
R27749 VGND.n8807 VGND.n8806 0.0145155
R27750 VGND.n293 VGND.n292 0.0145155
R27751 VGND.n292 VGND.n291 0.0145155
R27752 VGND.n2027 VGND.n2026 0.0145155
R27753 VGND.n2026 VGND.n2025 0.0145155
R27754 VGND.n473 VGND.n472 0.0145155
R27755 VGND.n7732 VGND.n7731 0.0145155
R27756 VGND.n7733 VGND.n7732 0.0145155
R27757 VGND.n745 VGND.n744 0.0145155
R27758 VGND.n744 VGND.n743 0.0145155
R27759 VGND.n8126 VGND.n8125 0.0145155
R27760 VGND.n8125 VGND.n8124 0.0145155
R27761 VGND.n424 VGND.n423 0.0145155
R27762 VGND.n7712 VGND.n7711 0.0145155
R27763 VGND.n7711 VGND.n7710 0.0145155
R27764 VGND.n7261 VGND.n7260 0.0145155
R27765 VGND.n7260 VGND.n7259 0.0145155
R27766 VGND.n1178 VGND.n1177 0.0145155
R27767 VGND.n1177 VGND.n1176 0.0145155
R27768 VGND.n771 VGND.n770 0.0145155
R27769 VGND.n770 VGND.n769 0.0145155
R27770 VGND.n853 VGND.n852 0.0145155
R27771 VGND.n854 VGND.n853 0.0145155
R27772 VGND.n6951 VGND.n6950 0.0145155
R27773 VGND.n6950 VGND.n6949 0.0145155
R27774 VGND.n6094 VGND.n6093 0.0145155
R27775 VGND.n1602 VGND.n1601 0.0145155
R27776 VGND.n1665 VGND.n1664 0.0145155
R27777 VGND.n5846 VGND.n5845 0.0145155
R27778 VGND.n5847 VGND.n5846 0.0145155
R27779 VGND.n2148 VGND.n2147 0.0145155
R27780 VGND.n2147 VGND.n2146 0.0145155
R27781 VGND.n6539 VGND.n6538 0.0145155
R27782 VGND.n6540 VGND.n6539 0.0145155
R27783 VGND.n5322 VGND.n5321 0.0145155
R27784 VGND.n5323 VGND.n5322 0.0145155
R27785 VGND.n5773 VGND.n5772 0.0145155
R27786 VGND.n5774 VGND.n5773 0.0145155
R27787 VGND.n2374 VGND.n2373 0.0145155
R27788 VGND.n2373 VGND.n2372 0.0145155
R27789 VGND.n5486 VGND.n5485 0.0145155
R27790 VGND.n5487 VGND.n5486 0.0145155
R27791 VGND.n2524 VGND.n2523 0.0145155
R27792 VGND.n2523 VGND.n2522 0.0145155
R27793 VGND.n3473 VGND.n3472 0.0145155
R27794 VGND.n5980 VGND.n5979 0.0145155
R27795 VGND.n5981 VGND.n5980 0.0145155
R27796 VGND.n5013 VGND.n5012 0.014042
R27797 VGND.n4378 VGND.n4377 0.014042
R27798 VGND.n3327 VGND.n3326 0.014042
R27799 VGND.n8912 VGND.n8911 0.014042
R27800 VGND.n8785 VGND.n157 0.014042
R27801 VGND.n6456 VGND.n1687 0.014042
R27802 VGND.n5816 VGND.n5122 0.014042
R27803 VGND.n2623 VGND.n2622 0.014042
R27804 VGND.n6003 VGND.n6002 0.0140135
R27805 VGND.n6000 VGND.n5999 0.0140135
R27806 VGND.n5984 VGND.n5978 0.0140135
R27807 VGND.n6740 VGND.n6739 0.0140135
R27808 VGND.n6757 VGND.n6751 0.0140135
R27809 VGND.n6074 VGND.n6073 0.0140135
R27810 VGND.n6071 VGND.n6070 0.0140135
R27811 VGND.n6081 VGND.n6077 0.0140135
R27812 VGND.n6535 VGND.n6529 0.0140135
R27813 VGND.n6535 VGND.n6534 0.0140135
R27814 VGND.n6543 VGND.n1656 0.0140135
R27815 VGND.n7094 VGND.n1358 0.0140135
R27816 VGND.n1367 VGND.n1366 0.0140135
R27817 VGND.n7086 VGND.n1367 0.0140135
R27818 VGND.n7250 VGND.n7249 0.0140135
R27819 VGND.n7235 VGND.n7231 0.0140135
R27820 VGND.n4840 VGND.n4839 0.0140135
R27821 VGND.n4842 VGND.n4841 0.0140135
R27822 VGND.n4831 VGND.n4827 0.0140135
R27823 VGND.n4071 VGND.n4065 0.0140135
R27824 VGND.n4071 VGND.n4070 0.0140135
R27825 VGND.n4993 VGND.n4073 0.0140135
R27826 VGND.n4735 VGND.n4734 0.0140135
R27827 VGND.n4730 VGND.n4147 0.0140135
R27828 VGND.n4742 VGND.n4738 0.0140135
R27829 VGND.n4195 VGND.n4194 0.0140135
R27830 VGND.n4201 VGND.n4197 0.0140135
R27831 VGND.n6986 VGND.n6985 0.0140135
R27832 VGND.n1561 VGND.n1560 0.0140135
R27833 VGND.n1566 VGND.n1561 0.0140135
R27834 VGND.n4351 VGND.n4350 0.0140135
R27835 VGND.n4350 VGND.n4312 0.0140135
R27836 VGND.n4342 VGND.n4316 0.0140135
R27837 VGND.n3003 VGND.n2884 0.0140135
R27838 VGND.n2991 VGND.n2990 0.0140135
R27839 VGND.n2995 VGND.n2991 0.0140135
R27840 VGND.n3556 VGND.n3555 0.0140135
R27841 VGND.n3558 VGND.n3557 0.0140135
R27842 VGND.n3547 VGND.n3543 0.0140135
R27843 VGND.n9082 VGND.n9081 0.0140135
R27844 VGND.n9073 VGND.n9072 0.0140135
R27845 VGND.n2141 VGND.n2135 0.0140135
R27846 VGND.n2141 VGND.n2140 0.0140135
R27847 VGND.n3354 VGND.n2128 0.0140135
R27848 VGND.n3158 VGND.n3141 0.0140135
R27849 VGND.n3146 VGND.n3145 0.0140135
R27850 VGND.n3150 VGND.n3146 0.0140135
R27851 VGND.n3596 VGND.n3595 0.0140135
R27852 VGND.n3593 VGND.n3592 0.0140135
R27853 VGND.n3603 VGND.n3599 0.0140135
R27854 VGND.n9060 VGND.n9059 0.0140135
R27855 VGND.n68 VGND.n62 0.0140135
R27856 VGND.n117 VGND.n111 0.0140135
R27857 VGND.n117 VGND.n116 0.0140135
R27858 VGND.n8832 VGND.n104 0.0140135
R27859 VGND.n8554 VGND.n8553 0.0140135
R27860 VGND.n268 VGND.n267 0.0140135
R27861 VGND.n8545 VGND.n268 0.0140135
R27862 VGND.n3742 VGND.n3741 0.0140135
R27863 VGND.n3739 VGND.n3738 0.0140135
R27864 VGND.n3749 VGND.n3745 0.0140135
R27865 VGND.n8675 VGND.n8674 0.0140135
R27866 VGND.n8693 VGND.n8692 0.0140135
R27867 VGND.n148 VGND.n142 0.0140135
R27868 VGND.n148 VGND.n147 0.0140135
R27869 VGND.n8803 VGND.n150 0.0140135
R27870 VGND.n8433 VGND.n8432 0.0140135
R27871 VGND.n284 VGND.n283 0.0140135
R27872 VGND.n288 VGND.n284 0.0140135
R27873 VGND.n2015 VGND.n2014 0.0140135
R27874 VGND.n2012 VGND.n2011 0.0140135
R27875 VGND.n2022 VGND.n2018 0.0140135
R27876 VGND.n471 VGND.n470 0.0140135
R27877 VGND.n8107 VGND.n8101 0.0140135
R27878 VGND.n555 VGND.n549 0.0140135
R27879 VGND.n555 VGND.n554 0.0140135
R27880 VGND.n7736 VGND.n542 0.0140135
R27881 VGND.n733 VGND.n732 0.0140135
R27882 VGND.n730 VGND.n729 0.0140135
R27883 VGND.n740 VGND.n736 0.0140135
R27884 VGND.n8208 VGND.n8207 0.0140135
R27885 VGND.n8121 VGND.n8117 0.0140135
R27886 VGND.n427 VGND.n420 0.0140135
R27887 VGND.n314 VGND.n313 0.0140135
R27888 VGND.n8325 VGND.n314 0.0140135
R27889 VGND.n595 VGND.n589 0.0140135
R27890 VGND.n595 VGND.n594 0.0140135
R27891 VGND.n7707 VGND.n597 0.0140135
R27892 VGND.n7270 VGND.n7269 0.0140135
R27893 VGND.n7288 VGND.n7282 0.0140135
R27894 VGND.n1181 VGND.n1172 0.0140135
R27895 VGND.n893 VGND.n892 0.0140135
R27896 VGND.n7301 VGND.n893 0.0140135
R27897 VGND.n7448 VGND.n7447 0.0140135
R27898 VGND.n7443 VGND.n774 0.0140135
R27899 VGND.n762 VGND.n756 0.0140135
R27900 VGND.n840 VGND.n836 0.0140135
R27901 VGND.n840 VGND.n839 0.0140135
R27902 VGND.n860 VGND.n851 0.0140135
R27903 VGND.n6948 VGND.n6947 0.0140135
R27904 VGND.n1546 VGND.n1545 0.0140135
R27905 VGND.n1551 VGND.n1546 0.0140135
R27906 VGND.n6168 VGND.n6167 0.0140135
R27907 VGND.n6191 VGND.n6096 0.0140135
R27908 VGND.n1610 VGND.n1609 0.0140135
R27909 VGND.n6778 VGND.n6772 0.0140135
R27910 VGND.n6490 VGND.n6486 0.0140135
R27911 VGND.n6490 VGND.n6489 0.0140135
R27912 VGND.n6473 VGND.n1667 0.0140135
R27913 VGND.n2160 VGND.n2154 0.0140135
R27914 VGND.n2160 VGND.n2159 0.0140135
R27915 VGND.n2272 VGND.n2268 0.0140135
R27916 VGND.n5318 VGND.n5317 0.0140135
R27917 VGND.n5293 VGND.n5292 0.0140135
R27918 VGND.n5326 VGND.n5293 0.0140135
R27919 VGND.n5769 VGND.n5768 0.0140135
R27920 VGND.n5780 VGND.n5779 0.0140135
R27921 VGND.n5785 VGND.n5780 0.0140135
R27922 VGND.n2377 VGND.n2366 0.0140135
R27923 VGND.n35 VGND.n34 0.0140135
R27924 VGND.n38 VGND.n35 0.0140135
R27925 VGND.n5482 VGND.n5481 0.0140135
R27926 VGND.n5625 VGND.n5624 0.0140135
R27927 VGND.n2534 VGND.n2533 0.0140135
R27928 VGND.n2325 VGND.n2322 0.0140135
R27929 VGND.n3532 VGND.n3531 0.0140135
R27930 VGND.n9230 VGND.n1 0.0140135
R27931 VGND.n9227 VGND.n9226 0.0140135
R27932 VGND.n5842 VGND.n5838 0.0140135
R27933 VGND.n5842 VGND.n5841 0.0140135
R27934 VGND.n5121 VGND.n5120 0.0140135
R27935 VGND.n4813 VGND 0.0135208
R27936 VGND.n4807 VGND.n4802 0.0135208
R27937 VGND.n4969 VGND.n4968 0.0135208
R27938 VGND.n4973 VGND.n4972 0.0135208
R27939 VGND.n7098 VGND.n7097 0.0135208
R27940 VGND.n4355 VGND.n4354 0.0135208
R27941 VGND.n4321 VGND.n4320 0.0135208
R27942 VGND VGND.n4379 0.0135208
R27943 VGND.n4571 VGND.n4570 0.0135208
R27944 VGND.n3461 VGND.n3460 0.0135208
R27945 VGND.n3375 VGND.n3374 0.0135208
R27946 VGND.n3370 VGND.n3368 0.0135208
R27947 VGND.n3325 VGND 0.0135208
R27948 VGND.n3007 VGND.n3006 0.0135208
R27949 VGND.n3711 VGND.n3710 0.0135208
R27950 VGND.n8853 VGND.n8852 0.0135208
R27951 VGND.n8848 VGND.n8846 0.0135208
R27952 VGND VGND.n8913 0.0135208
R27953 VGND.n3162 VGND.n3161 0.0135208
R27954 VGND.n3821 VGND.n3820 0.0135208
R27955 VGND.n3912 VGND.n3911 0.0135208
R27956 VGND.n3907 VGND.n3905 0.0135208
R27957 VGND VGND.n160 0.0135208
R27958 VGND.n8561 VGND.n8560 0.0135208
R27959 VGND.n1993 VGND 0.0135208
R27960 VGND.n1987 VGND.n1986 0.0135208
R27961 VGND.n7755 VGND.n7754 0.0135208
R27962 VGND.n7751 VGND.n7750 0.0135208
R27963 VGND VGND.n7818 0.0135208
R27964 VGND.n7540 VGND.n7539 0.0135208
R27965 VGND.n7627 VGND.n7626 0.0135208
R27966 VGND.n7622 VGND.n7620 0.0135208
R27967 VGND.n681 VGND 0.0135208
R27968 VGND.n431 VGND.n430 0.0135208
R27969 VGND.n786 VGND.n785 0.0135208
R27970 VGND.n863 VGND.n862 0.0135208
R27971 VGND VGND.n1019 0.0135208
R27972 VGND.n1185 VGND.n1184 0.0135208
R27973 VGND.n1674 VGND.n1673 0.0135208
R27974 VGND VGND.n6340 0.0135208
R27975 VGND.n6943 VGND.n6942 0.0135208
R27976 VGND VGND.n1757 0.0135208
R27977 VGND.n1764 VGND.n1763 0.0135208
R27978 VGND.n6569 VGND.n6568 0.0135208
R27979 VGND.n6562 VGND.n6560 0.0135208
R27980 VGND VGND.n6634 0.0135208
R27981 VGND.n5309 VGND.n5308 0.0135208
R27982 VGND.n1843 VGND.n1842 0.0135208
R27983 VGND.n5886 VGND.n5885 0.0135208
R27984 VGND.n5881 VGND.n5879 0.0135208
R27985 VGND VGND.n5499 0.0135208
R27986 VGND.n5764 VGND.n5763 0.0135208
R27987 VGND.n3527 VGND.n3526 0.0135208
R27988 VGND.n2250 VGND.n2249 0.0135208
R27989 VGND.n2257 VGND.n2255 0.0135208
R27990 VGND.n2621 VGND 0.0135208
R27991 VGND.n2381 VGND.n2380 0.0135208
R27992 VGND.n1618 VGND.n1617 0.0130912
R27993 VGND.n1778 VGND.n1777 0.0130912
R27994 VGND.n1377 VGND.n1376 0.0130912
R27995 VGND.n1325 VGND.n1324 0.0130912
R27996 VGND.n4755 VGND.n4754 0.0130912
R27997 VGND.n4046 VGND.n4045 0.0130912
R27998 VGND.n4702 VGND.n4701 0.0130912
R27999 VGND.n4179 VGND.n4178 0.0130912
R28000 VGND.n4228 VGND.n4227 0.0130912
R28001 VGND.n2973 VGND.n2972 0.0130912
R28002 VGND.n2095 VGND.n2094 0.0130912
R28003 VGND.n2636 VGND.n2635 0.0130912
R28004 VGND.n2743 VGND.n2742 0.0130912
R28005 VGND.n3624 VGND.n3623 0.0130912
R28006 VGND.n121 VGND.n120 0.0130912
R28007 VGND.n278 VGND.n277 0.0130912
R28008 VGND.n1872 VGND.n1871 0.0130912
R28009 VGND.n8792 VGND.n8791 0.0130912
R28010 VGND.n8411 VGND.n8410 0.0130912
R28011 VGND.n1964 VGND.n1963 0.0130912
R28012 VGND.n559 VGND.n558 0.0130912
R28013 VGND.n7510 VGND.n7509 0.0130912
R28014 VGND.n8149 VGND.n8148 0.0130912
R28015 VGND.n7696 VGND.n7695 0.0130912
R28016 VGND.n7257 VGND.n7256 0.0130912
R28017 VGND.n1142 VGND.n1141 0.0130912
R28018 VGND.n1174 VGND.n1173 0.0130912
R28019 VGND.n897 VGND.n896 0.0130912
R28020 VGND.n767 VGND.n766 0.0130912
R28021 VGND.n750 VGND.n749 0.0130912
R28022 VGND.n822 VGND.n821 0.0130912
R28023 VGND.n857 VGND.n856 0.0130912
R28024 VGND.n6926 VGND.n6925 0.0130912
R28025 VGND.n1541 VGND.n1540 0.0130912
R28026 VGND.n6162 VGND.n6161 0.0130912
R28027 VGND.n6478 VGND.n6477 0.0130912
R28028 VGND.n1662 VGND.n1661 0.0130912
R28029 VGND.n5832 VGND.n5831 0.0130912
R28030 VGND.n2269 VGND.n2164 0.0130912
R28031 VGND.n6503 VGND.n6502 0.0130912
R28032 VGND.n6508 VGND.n6507 0.0130912
R28033 VGND.n5218 VGND.n5217 0.0130912
R28034 VGND.n5748 VGND.n5747 0.0130912
R28035 VGND.n42 VGND.n41 0.0130912
R28036 VGND.n5494 VGND.n5493 0.0130912
R28037 VGND.n2329 VGND.n2328 0.0130912
R28038 VGND.n3470 VGND.n3469 0.0130912
R28039 VGND.n9223 VGND.n9222 0.0130912
R28040 VGND.n1787 VGND.n1786 0.0130912
R28041 VGND.n1852 VGND.n1851 0.0130912
R28042 VGND.n1140 VGND.n1139 0.0126061
R28043 VGND.n1321 VGND.n1320 0.0126061
R28044 VGND.n1200 VGND.n998 0.0126061
R28045 VGND.n991 VGND.n990 0.0126061
R28046 VGND.n7499 VGND.n7498 0.0126061
R28047 VGND.n799 VGND.n751 0.0126061
R28048 VGND.n7329 VGND.n7328 0.0126061
R28049 VGND.n7326 VGND.n7325 0.0126061
R28050 VGND.n6928 VGND.n6927 0.0126061
R28051 VGND.n6160 VGND.n6159 0.0126061
R28052 VGND.n6268 VGND.n1660 0.0126061
R28053 VGND.n6750 VGND.n6749 0.0123243
R28054 VGND.n6757 VGND.n6756 0.0123243
R28055 VGND.n6534 VGND.n6533 0.0123243
R28056 VGND.n7235 VGND.n7234 0.0123243
R28057 VGND.n4070 VGND.n4069 0.0123243
R28058 VGND.n4201 VGND.n4200 0.0123243
R28059 VGND.n4324 VGND.n4312 0.0123243
R28060 VGND.n9074 VGND.n53 0.0123243
R28061 VGND.n9072 VGND.n54 0.0123243
R28062 VGND.n2140 VGND.n2139 0.0123243
R28063 VGND.n61 VGND.n60 0.0123243
R28064 VGND.n68 VGND.n67 0.0123243
R28065 VGND.n116 VGND.n115 0.0123243
R28066 VGND.n8694 VGND.n8681 0.0123243
R28067 VGND.n8692 VGND.n8686 0.0123243
R28068 VGND.n147 VGND.n146 0.0123243
R28069 VGND.n8100 VGND.n8099 0.0123243
R28070 VGND.n8107 VGND.n8106 0.0123243
R28071 VGND.n554 VGND.n553 0.0123243
R28072 VGND.n8121 VGND.n8120 0.0123243
R28073 VGND.n594 VGND.n593 0.0123243
R28074 VGND.n7281 VGND.n7280 0.0123243
R28075 VGND.n7288 VGND.n7287 0.0123243
R28076 VGND.n781 VGND.n780 0.0123243
R28077 VGND.n839 VGND.n838 0.0123243
R28078 VGND.n6103 VGND.n6102 0.0123243
R28079 VGND.n6771 VGND.n6770 0.0123243
R28080 VGND.n6778 VGND.n6777 0.0123243
R28081 VGND.n6489 VGND.n6488 0.0123243
R28082 VGND.n2159 VGND.n2158 0.0123243
R28083 VGND.n5627 VGND.n5626 0.0123243
R28084 VGND.n5624 VGND.n5477 0.0123243
R28085 VGND.n2325 VGND.n2324 0.0123243
R28086 VGND.n3481 VGND.n3480 0.0123243
R28087 VGND.n5841 VGND.n5840 0.0123243
R28088 VGND.n4855 VGND.n4853 0.0122188
R28089 VGND.n7220 VGND.n7217 0.0122188
R28090 VGND.n7070 VGND 0.0122188
R28091 VGND.n4724 VGND.n4722 0.0122188
R28092 VGND VGND.n4720 0.0122188
R28093 VGND VGND.n4356 0.0122188
R28094 VGND.n4512 VGND.n4508 0.0122188
R28095 VGND.n3566 VGND.n3565 0.0122188
R28096 VGND.n2774 VGND.n2771 0.0122188
R28097 VGND.n9043 VGND.n9037 0.0122188
R28098 VGND.n3833 VGND.n3831 0.0122188
R28099 VGND VGND.n3913 0.0122188
R28100 VGND.n8704 VGND.n8698 0.0122188
R28101 VGND.n8525 VGND 0.0122188
R28102 VGND.n7817 VGND.n7816 0.0122188
R28103 VGND.n8089 VGND.n8084 0.0122188
R28104 VGND.n7554 VGND.n7552 0.0122188
R28105 VGND.n7688 VGND.n682 0.0122188
R28106 VGND.n8196 VGND.n8195 0.0122188
R28107 VGND VGND.n405 0.0122188
R28108 VGND.n7437 VGND.n7434 0.0122188
R28109 VGND.n861 VGND 0.0122188
R28110 VGND.n7316 VGND.n885 0.0122188
R28111 VGND.n1315 VGND.n1309 0.0122188
R28112 VGND.n6184 VGND.n6182 0.0122188
R28113 VGND.n6188 VGND 0.0122188
R28114 VGND.n6817 VGND.n6815 0.0122188
R28115 VGND.n6063 VGND.n6061 0.0122188
R28116 VGND.n6633 VGND.n6632 0.0122188
R28117 VGND.n5366 VGND.n5358 0.0122188
R28118 VGND.n5285 VGND 0.0122188
R28119 VGND.n5992 VGND.n5990 0.0122188
R28120 VGND VGND.n5988 0.0122188
R28121 VGND VGND.n5887 0.0122188
R28122 VGND.n5637 VGND.n5634 0.0122188
R28123 VGND.n9215 VGND 0.0122188
R28124 VGND.n2248 VGND 0.0122188
R28125 VGND.n2511 VGND.n2508 0.0122188
R28126 VGND.n6958 VGND.n6956 0.0118576
R28127 VGND.n6210 VGND.n6208 0.0118576
R28128 VGND.n6462 VGND.n1663 0.0118576
R28129 VGND.n6790 VGND.n6789 0.0118576
R28130 VGND.n6786 VGND.n6784 0.0118576
R28131 VGND.n4057 VGND.n4056 0.0117818
R28132 VGND.n1362 VGND.n1361 0.0117818
R28133 VGND.n7255 VGND.n7254 0.0117818
R28134 VGND.n4094 VGND.n765 0.0117818
R28135 VGND.n6 VGND.n5 0.0115273
R28136 VGND.n4798 VGND.n4797 0.0114169
R28137 VGND.n4128 VGND.n4127 0.0114169
R28138 VGND.n2077 VGND.n2076 0.0114169
R28139 VGND.n3698 VGND.n3697 0.0114169
R28140 VGND.n3809 VGND.n3808 0.0114169
R28141 VGND.n1915 VGND.n1914 0.0114169
R28142 VGND.n7527 VGND.n719 0.0114169
R28143 VGND.n7488 VGND.n7487 0.0114169
R28144 VGND.n6150 VGND.n6149 0.0114169
R28145 VGND.n1746 VGND.n1743 0.0114169
R28146 VGND.n1830 VGND.n1829 0.0114169
R28147 VGND.n3514 VGND.n3513 0.0114169
R28148 VGND.n3718 VGND.n3717 0.0111911
R28149 VGND.n1980 VGND.n1976 0.0111911
R28150 VGND.n4845 VGND.n4844 0.0109167
R28151 VGND.n4850 VGND.n4848 0.0109167
R28152 VGND.n7107 VGND.n7104 0.0109167
R28153 VGND.n7104 VGND.n7102 0.0109167
R28154 VGND.n7099 VGND 0.0109167
R28155 VGND VGND.n7002 0.0109167
R28156 VGND.n4732 VGND.n4731 0.0109167
R28157 VGND.n4727 VGND.n4726 0.0109167
R28158 VGND VGND.n4306 0.0109167
R28159 VGND.n4357 VGND 0.0109167
R28160 VGND.n4578 VGND.n4577 0.0109167
R28161 VGND.n4577 VGND.n4576 0.0109167
R28162 VGND.n4572 VGND 0.0109167
R28163 VGND.n3561 VGND.n3560 0.0109167
R28164 VGND.n3564 VGND.n3563 0.0109167
R28165 VGND.n9075 VGND 0.0109167
R28166 VGND.n3008 VGND 0.0109167
R28167 VGND.n3714 VGND.n3713 0.0109167
R28168 VGND.n3170 VGND.n3167 0.0109167
R28169 VGND.n3167 VGND.n3165 0.0109167
R28170 VGND.n3163 VGND 0.0109167
R28171 VGND.n3824 VGND.n3823 0.0109167
R28172 VGND.n3829 VGND.n3827 0.0109167
R28173 VGND VGND.n8695 0.0109167
R28174 VGND.n8568 VGND.n8566 0.0109167
R28175 VGND.n8566 VGND.n8564 0.0109167
R28176 VGND VGND.n8450 0.0109167
R28177 VGND.n1984 VGND.n1983 0.0109167
R28178 VGND VGND.n7980 0.0109167
R28179 VGND.n7543 VGND.n7542 0.0109167
R28180 VGND.n7550 VGND.n7548 0.0109167
R28181 VGND.n439 VGND.n437 0.0109167
R28182 VGND.n437 VGND.n435 0.0109167
R28183 VGND.n432 VGND 0.0109167
R28184 VGND.n406 VGND 0.0109167
R28185 VGND.n7445 VGND.n7444 0.0109167
R28186 VGND.n7440 VGND.n7439 0.0109167
R28187 VGND.n7334 VGND 0.0109167
R28188 VGND VGND.n7333 0.0109167
R28189 VGND.n1193 VGND.n1190 0.0109167
R28190 VGND.n1190 VGND.n1188 0.0109167
R28191 VGND.n1186 VGND 0.0109167
R28192 VGND.n6175 VGND.n6171 0.0109167
R28193 VGND.n6180 VGND.n6178 0.0109167
R28194 VGND VGND.n6812 0.0109167
R28195 VGND.n6938 VGND.n6936 0.0109167
R28196 VGND.n6940 VGND.n6938 0.0109167
R28197 VGND VGND.n6941 0.0109167
R28198 VGND.n6069 VGND.n1766 0.0109167
R28199 VGND.n6066 VGND.n6065 0.0109167
R28200 VGND VGND.n1771 0.0109167
R28201 VGND VGND.n5307 0.0109167
R28202 VGND VGND.n5222 0.0109167
R28203 VGND.n5998 VGND.n1845 0.0109167
R28204 VGND.n5995 VGND.n5994 0.0109167
R28205 VGND VGND.n5631 0.0109167
R28206 VGND.n5759 VGND.n5757 0.0109167
R28207 VGND.n5761 VGND.n5759 0.0109167
R28208 VGND VGND.n5762 0.0109167
R28209 VGND.n9232 VGND.n9231 0.0109167
R28210 VGND.n2389 VGND.n2386 0.0109167
R28211 VGND.n2386 VGND.n2384 0.0109167
R28212 VGND.n2382 VGND 0.0109167
R28213 VGND.n6756 VGND.n6755 0.0106351
R28214 VGND.n6753 VGND.n6752 0.0106351
R28215 VGND.n6533 VGND.n6532 0.0106351
R28216 VGND.n6520 VGND.n6509 0.0106351
R28217 VGND.n6994 VGND.n6993 0.0106351
R28218 VGND.n7085 VGND.n1369 0.0106351
R28219 VGND.n1372 VGND.n1371 0.0106351
R28220 VGND.n7072 VGND.n7071 0.0106351
R28221 VGND.n7234 VGND.n7233 0.0106351
R28222 VGND.n1327 VGND.n1326 0.0106351
R28223 VGND.n4069 VGND.n4068 0.0106351
R28224 VGND.n5005 VGND.n4043 0.0106351
R28225 VGND.n4200 VGND.n4199 0.0106351
R28226 VGND.n4175 VGND.n4174 0.0106351
R28227 VGND.n4581 VGND.n4580 0.0106351
R28228 VGND.n1565 VGND.n1564 0.0106351
R28229 VGND.n4325 VGND.n4324 0.0106351
R28230 VGND.n4370 VGND.n4225 0.0106351
R28231 VGND.n3015 VGND.n3014 0.0106351
R28232 VGND.n2994 VGND.n2993 0.0106351
R28233 VGND.n2968 VGND.n2967 0.0106351
R28234 VGND.n2769 VGND.n54 0.0106351
R28235 VGND.n2767 VGND.n2766 0.0106351
R28236 VGND.n2139 VGND.n2138 0.0106351
R28237 VGND.n3332 VGND.n2639 0.0106351
R28238 VGND.n3176 VGND.n3175 0.0106351
R28239 VGND.n3149 VGND.n3148 0.0106351
R28240 VGND.n2738 VGND.n2737 0.0106351
R28241 VGND.n67 VGND.n66 0.0106351
R28242 VGND.n64 VGND.n63 0.0106351
R28243 VGND.n115 VGND.n114 0.0106351
R28244 VGND.n132 VGND.n124 0.0106351
R28245 VGND.n8442 VGND.n8441 0.0106351
R28246 VGND.n8544 VGND.n270 0.0106351
R28247 VGND.n273 VGND.n272 0.0106351
R28248 VGND.n8527 VGND.n8526 0.0106351
R28249 VGND.n8686 VGND.n8685 0.0106351
R28250 VGND.n8683 VGND.n8682 0.0106351
R28251 VGND.n146 VGND.n145 0.0106351
R28252 VGND.n8796 VGND.n8795 0.0106351
R28253 VGND.n7970 VGND.n7969 0.0106351
R28254 VGND.n287 VGND.n286 0.0106351
R28255 VGND.n8406 VGND.n8405 0.0106351
R28256 VGND.n8106 VGND.n8105 0.0106351
R28257 VGND.n8103 VGND.n8102 0.0106351
R28258 VGND.n553 VGND.n552 0.0106351
R28259 VGND.n569 VGND.n560 0.0106351
R28260 VGND.n8120 VGND.n8119 0.0106351
R28261 VGND.n8145 VGND.n8144 0.0106351
R28262 VGND.n8315 VGND.n8314 0.0106351
R28263 VGND.n8329 VGND.n8328 0.0106351
R28264 VGND.n404 VGND.n323 0.0106351
R28265 VGND.n593 VGND.n592 0.0106351
R28266 VGND.n7700 VGND.n7699 0.0106351
R28267 VGND.n7287 VGND.n7286 0.0106351
R28268 VGND.n7284 VGND.n7283 0.0106351
R28269 VGND.n1198 VGND.n1197 0.0106351
R28270 VGND.n7305 VGND.n7304 0.0106351
R28271 VGND.n838 VGND.n837 0.0106351
R28272 VGND.n7324 VGND.n845 0.0106351
R28273 VGND.n1550 VGND.n1549 0.0106351
R28274 VGND.n6777 VGND.n6776 0.0106351
R28275 VGND.n6774 VGND.n6773 0.0106351
R28276 VGND.n6488 VGND.n6487 0.0106351
R28277 VGND.n6463 VGND.n6460 0.0106351
R28278 VGND.n2158 VGND.n2157 0.0106351
R28279 VGND.n2628 VGND.n2166 0.0106351
R28280 VGND.n5459 VGND.n5458 0.0106351
R28281 VGND.n5329 VGND.n5328 0.0106351
R28282 VGND.n5213 VGND.n5212 0.0106351
R28283 VGND.n5287 VGND.n5286 0.0106351
R28284 VGND.n5744 VGND.n5743 0.0106351
R28285 VGND.n5784 VGND.n5783 0.0106351
R28286 VGND.n2393 VGND.n2392 0.0106351
R28287 VGND.n37 VGND.n36 0.0106351
R28288 VGND.n30 VGND.n29 0.0106351
R28289 VGND.n5477 VGND.n5476 0.0106351
R28290 VGND.n5474 VGND.n5473 0.0106351
R28291 VGND.n2324 VGND.n2323 0.0106351
R28292 VGND.n2333 VGND.n2332 0.0106351
R28293 VGND.n5840 VGND.n5839 0.0106351
R28294 VGND.n5856 VGND.n5820 0.0106351
R28295 VGND.n3236 VGND.n3235 0.0103319
R28296 VGND.n8801 VGND.n153 0.0102388
R28297 VGND.n6471 VGND.n1686 0.0102388
R28298 VGND.n6743 VGND.n6742 0.00975758
R28299 VGND.n6746 VGND.n6745 0.00975758
R28300 VGND.n6760 VGND.n6759 0.00975758
R28301 VGND.n6088 VGND.n1699 0.00975758
R28302 VGND.n6087 VGND.n6086 0.00975758
R28303 VGND.n6084 VGND.n6083 0.00975758
R28304 VGND.n7093 VGND.n1360 0.00975758
R28305 VGND.n7092 VGND.n7091 0.00975758
R28306 VGND.n7089 VGND.n7088 0.00975758
R28307 VGND.n7251 VGND.n7229 0.00975758
R28308 VGND.n7241 VGND.n7240 0.00975758
R28309 VGND.n7238 VGND.n7237 0.00975758
R28310 VGND.n4838 VGND.n4093 0.00975758
R28311 VGND.n4837 VGND.n4836 0.00975758
R28312 VGND.n4834 VGND.n4833 0.00975758
R28313 VGND.n5000 VGND.n4060 0.00975758
R28314 VGND.n4999 VGND.n4998 0.00975758
R28315 VGND.n4996 VGND.n4995 0.00975758
R28316 VGND.n4749 VGND.n4145 0.00975758
R28317 VGND.n4748 VGND.n4747 0.00975758
R28318 VGND.n4745 VGND.n4744 0.00975758
R28319 VGND.n4208 VGND.n4186 0.00975758
R28320 VGND.n4207 VGND.n4206 0.00975758
R28321 VGND.n4204 VGND.n4203 0.00975758
R28322 VGND.n6987 VGND.n1380 0.00975758
R28323 VGND.n1383 VGND.n1382 0.00975758
R28324 VGND.n1555 VGND.n1554 0.00975758
R28325 VGND.n1567 VGND.n1557 0.00975758
R28326 VGND.n4349 VGND.n4314 0.00975758
R28327 VGND.n4348 VGND.n4347 0.00975758
R28328 VGND.n4345 VGND.n4344 0.00975758
R28329 VGND.n3002 VGND.n2886 0.00975758
R28330 VGND.n3001 VGND.n3000 0.00975758
R28331 VGND.n2998 VGND.n2997 0.00975758
R28332 VGND.n3554 VGND.n3465 0.00975758
R28333 VGND.n3553 VGND.n3552 0.00975758
R28334 VGND.n3550 VGND.n3549 0.00975758
R28335 VGND.n9086 VGND.n49 0.00975758
R28336 VGND.n9085 VGND.n9084 0.00975758
R28337 VGND.n56 VGND.n55 0.00975758
R28338 VGND.n9071 VGND.n9070 0.00975758
R28339 VGND.n3347 VGND.n2130 0.00975758
R28340 VGND.n3349 VGND.n3348 0.00975758
R28341 VGND.n3352 VGND.n3351 0.00975758
R28342 VGND.n3157 VGND.n3143 0.00975758
R28343 VGND.n3156 VGND.n3155 0.00975758
R28344 VGND.n3153 VGND.n3152 0.00975758
R28345 VGND.n3610 VGND.n3586 0.00975758
R28346 VGND.n3609 VGND.n3608 0.00975758
R28347 VGND.n3606 VGND.n3605 0.00975758
R28348 VGND.n9064 VGND.n9052 0.00975758
R28349 VGND.n9063 VGND.n9062 0.00975758
R28350 VGND.n59 VGND.n58 0.00975758
R28351 VGND.n71 VGND.n70 0.00975758
R28352 VGND.n8825 VGND.n106 0.00975758
R28353 VGND.n8827 VGND.n8826 0.00975758
R28354 VGND.n8830 VGND.n8829 0.00975758
R28355 VGND.n8552 VGND.n264 0.00975758
R28356 VGND.n8551 VGND.n8550 0.00975758
R28357 VGND.n8548 VGND.n8547 0.00975758
R28358 VGND.n3756 VGND.n3732 0.00975758
R28359 VGND.n3755 VGND.n3754 0.00975758
R28360 VGND.n3752 VGND.n3751 0.00975758
R28361 VGND.n8673 VGND.n8669 0.00975758
R28362 VGND.n8672 VGND.n8671 0.00975758
R28363 VGND.n8688 VGND.n8687 0.00975758
R28364 VGND.n8691 VGND.n8690 0.00975758
R28365 VGND.n8810 VGND.n137 0.00975758
R28366 VGND.n8809 VGND.n8808 0.00975758
R28367 VGND.n8806 VGND.n8805 0.00975758
R28368 VGND.n8434 VGND.n281 0.00975758
R28369 VGND.n294 VGND.n293 0.00975758
R28370 VGND.n291 VGND.n290 0.00975758
R28371 VGND.n2029 VGND.n2005 0.00975758
R28372 VGND.n2028 VGND.n2027 0.00975758
R28373 VGND.n2025 VGND.n2024 0.00975758
R28374 VGND.n475 VGND.n463 0.00975758
R28375 VGND.n474 VGND.n473 0.00975758
R28376 VGND.n8098 VGND.n8097 0.00975758
R28377 VGND.n8110 VGND.n8109 0.00975758
R28378 VGND.n7729 VGND.n544 0.00975758
R28379 VGND.n7731 VGND.n7730 0.00975758
R28380 VGND.n7734 VGND.n7733 0.00975758
R28381 VGND.n747 VGND.n723 0.00975758
R28382 VGND.n746 VGND.n745 0.00975758
R28383 VGND.n743 VGND.n742 0.00975758
R28384 VGND.n8209 VGND.n8115 0.00975758
R28385 VGND.n8127 VGND.n8126 0.00975758
R28386 VGND.n8124 VGND.n8123 0.00975758
R28387 VGND.n426 VGND.n422 0.00975758
R28388 VGND.n425 VGND.n424 0.00975758
R28389 VGND.n316 VGND.n315 0.00975758
R28390 VGND.n8324 VGND.n8323 0.00975758
R28391 VGND.n7714 VGND.n584 0.00975758
R28392 VGND.n7713 VGND.n7712 0.00975758
R28393 VGND.n7710 VGND.n7709 0.00975758
R28394 VGND.n7271 VGND.n7258 0.00975758
R28395 VGND.n7262 VGND.n7261 0.00975758
R28396 VGND.n7290 VGND.n7289 0.00975758
R28397 VGND.n1180 VGND.n1175 0.00975758
R28398 VGND.n1179 VGND.n1178 0.00975758
R28399 VGND.n7300 VGND.n7299 0.00975758
R28400 VGND.n7449 VGND.n768 0.00975758
R28401 VGND.n772 VGND.n771 0.00975758
R28402 VGND.n764 VGND.n763 0.00975758
R28403 VGND.n841 VGND.n830 0.00975758
R28404 VGND.n855 VGND.n854 0.00975758
R28405 VGND.n859 VGND.n858 0.00975758
R28406 VGND.n6953 VGND.n1572 0.00975758
R28407 VGND.n6952 VGND.n6951 0.00975758
R28408 VGND.n1553 VGND.n1552 0.00975758
R28409 VGND.n6166 VGND.n6163 0.00975758
R28410 VGND.n6165 VGND.n6164 0.00975758
R28411 VGND.n6095 VGND.n6094 0.00975758
R28412 VGND.n6194 VGND.n6193 0.00975758
R28413 VGND.n1611 VGND.n1600 0.00975758
R28414 VGND.n1603 VGND.n1602 0.00975758
R28415 VGND.n6766 VGND.n6765 0.00975758
R28416 VGND.n6779 VGND.n6768 0.00975758
R28417 VGND.n6491 VGND.n6479 0.00975758
R28418 VGND.n6481 VGND.n6480 0.00975758
R28419 VGND.n1666 VGND.n1665 0.00975758
R28420 VGND.n6475 VGND.n6474 0.00975758
R28421 VGND.n5845 VGND.n5844 0.00975758
R28422 VGND.n5848 VGND.n5847 0.00975758
R28423 VGND.n5851 VGND.n5850 0.00975758
R28424 VGND.n2161 VGND.n2144 0.00975758
R28425 VGND.n2149 VGND.n2148 0.00975758
R28426 VGND.n2146 VGND.n2145 0.00975758
R28427 VGND.n2271 VGND.n2270 0.00975758
R28428 VGND.n6536 VGND.n1657 0.00975758
R28429 VGND.n6538 VGND.n6537 0.00975758
R28430 VGND.n6541 VGND.n6540 0.00975758
R28431 VGND.n5319 VGND.n5295 0.00975758
R28432 VGND.n5321 VGND.n5320 0.00975758
R28433 VGND.n5324 VGND.n5323 0.00975758
R28434 VGND.n5772 VGND.n5771 0.00975758
R28435 VGND.n5775 VGND.n5774 0.00975758
R28436 VGND.n5788 VGND.n5787 0.00975758
R28437 VGND.n2376 VGND.n2368 0.00975758
R28438 VGND.n2375 VGND.n2374 0.00975758
R28439 VGND.n2372 VGND.n2371 0.00975758
R28440 VGND.n40 VGND.n39 0.00975758
R28441 VGND.n5485 VGND.n5484 0.00975758
R28442 VGND.n5488 VGND.n5487 0.00975758
R28443 VGND.n5623 VGND.n5622 0.00975758
R28444 VGND.n2535 VGND.n2520 0.00975758
R28445 VGND.n2525 VGND.n2524 0.00975758
R28446 VGND.n2522 VGND.n2521 0.00975758
R28447 VGND.n2327 VGND.n2326 0.00975758
R28448 VGND.n3533 VGND.n3471 0.00975758
R28449 VGND.n3474 VGND.n3473 0.00975758
R28450 VGND.n9219 VGND.n9218 0.00975758
R28451 VGND.n9225 VGND.n9224 0.00975758
R28452 VGND.n6004 VGND.n1790 0.00975758
R28453 VGND.n5979 VGND.n1791 0.00975758
R28454 VGND.n5982 VGND.n5981 0.00975758
R28455 VGND.n4797 VGND.n4795 0.00961458
R28456 VGND.n4812 VGND.n4811 0.00961458
R28457 VGND.n4974 VGND.n4973 0.00961458
R28458 VGND.n7214 VGND.n7213 0.00961458
R28459 VGND.n7109 VGND.n7107 0.00961458
R28460 VGND VGND.n7098 0.00961458
R28461 VGND.n4127 VGND.n4125 0.00961458
R28462 VGND VGND.n4321 0.00961458
R28463 VGND.n4505 VGND.n4504 0.00961458
R28464 VGND.n4579 VGND.n4578 0.00961458
R28465 VGND VGND.n4571 0.00961458
R28466 VGND.n2076 VGND.n2074 0.00961458
R28467 VGND.n3368 VGND.n3366 0.00961458
R28468 VGND VGND.n9076 0.00961458
R28469 VGND.n9076 VGND.n9075 0.00961458
R28470 VGND VGND.n3007 0.00961458
R28471 VGND.n3697 VGND.n3696 0.00961458
R28472 VGND.n3704 VGND.n3703 0.00961458
R28473 VGND.n8846 VGND.n8844 0.00961458
R28474 VGND.n9034 VGND.n9033 0.00961458
R28475 VGND.n3172 VGND.n3170 0.00961458
R28476 VGND VGND.n3162 0.00961458
R28477 VGND.n3808 VGND.n3803 0.00961458
R28478 VGND.n3816 VGND.n3815 0.00961458
R28479 VGND.n3905 VGND.n3903 0.00961458
R28480 VGND.n8680 VGND 0.00961458
R28481 VGND.n8695 VGND.n8680 0.00961458
R28482 VGND.n8570 VGND.n8568 0.00961458
R28483 VGND.n1914 VGND.n1910 0.00961458
R28484 VGND.n1992 VGND.n1991 0.00961458
R28485 VGND.n7750 VGND.n7749 0.00961458
R28486 VGND.n8081 VGND.n8080 0.00961458
R28487 VGND.n719 VGND.n717 0.00961458
R28488 VGND VGND.n7528 0.00961458
R28489 VGND.n7533 VGND.n7532 0.00961458
R28490 VGND.n7620 VGND.n7618 0.00961458
R28491 VGND.n8200 VGND.n8199 0.00961458
R28492 VGND.n8311 VGND.n439 0.00961458
R28493 VGND VGND.n431 0.00961458
R28494 VGND.n7487 VGND.n7485 0.00961458
R28495 VGND.n776 VGND.n775 0.00961458
R28496 VGND VGND.n794 0.00961458
R28497 VGND.n1306 VGND.n1305 0.00961458
R28498 VGND.n1196 VGND.n1193 0.00961458
R28499 VGND VGND.n1185 0.00961458
R28500 VGND.n6149 VGND.n6147 0.00961458
R28501 VGND.n6107 VGND.n6106 0.00961458
R28502 VGND.n6812 VGND.n6811 0.00961458
R28503 VGND.n6936 VGND.n6933 0.00961458
R28504 VGND.n6942 VGND 0.00961458
R28505 VGND.n1743 VGND.n1741 0.00961458
R28506 VGND.n1745 VGND 0.00961458
R28507 VGND.n1759 VGND.n1758 0.00961458
R28508 VGND.n6560 VGND.n6558 0.00961458
R28509 VGND.n5355 VGND.n5354 0.00961458
R28510 VGND.n5308 VGND 0.00961458
R28511 VGND.n1829 VGND.n1827 0.00961458
R28512 VGND.n1837 VGND.n1836 0.00961458
R28513 VGND.n5879 VGND.n5877 0.00961458
R28514 VGND.n5631 VGND.n5630 0.00961458
R28515 VGND.n5757 VGND.n5754 0.00961458
R28516 VGND.n5763 VGND 0.00961458
R28517 VGND.n3513 VGND.n3511 0.00961458
R28518 VGND.n3521 VGND.n3520 0.00961458
R28519 VGND.n2259 VGND.n2257 0.00961458
R28520 VGND.n2505 VGND.n2504 0.00961458
R28521 VGND.n2391 VGND.n2389 0.00961458
R28522 VGND VGND.n2381 0.00961458
R28523 VGND.n1855 VGND.n1854 0.00894595
R28524 VGND.n6733 VGND.n6728 0.00894595
R28525 VGND.n6733 VGND.n6732 0.00894595
R28526 VGND.n5346 VGND.n5345 0.00894595
R28527 VGND.n6015 VGND.n6014 0.00894595
R28528 VGND.n6501 VGND.n6498 0.00894595
R28529 VGND.n6526 VGND.n6525 0.00894595
R28530 VGND.n6529 VGND.n6528 0.00894595
R28531 VGND.n6520 VGND.n6519 0.00894595
R28532 VGND.n6995 VGND.n1353 0.00894595
R28533 VGND.n1366 VGND.n1365 0.00894595
R28534 VGND.n1369 VGND.n1368 0.00894595
R28535 VGND.n7073 VGND.n7001 0.00894595
R28536 VGND.n4003 VGND.n4002 0.00894595
R28537 VGND.n4002 VGND.n3998 0.00894595
R28538 VGND.n7248 VGND.n7247 0.00894595
R28539 VGND.n7224 VGND.n7223 0.00894595
R28540 VGND.n4761 VGND.n4090 0.00894595
R28541 VGND.n4053 VGND.n4050 0.00894595
R28542 VGND.n4062 VGND.n4061 0.00894595
R28543 VGND.n4065 VGND.n4064 0.00894595
R28544 VGND.n5008 VGND.n5005 0.00894595
R28545 VGND.n4710 VGND.n4709 0.00894595
R28546 VGND.n4485 VGND.n4482 0.00894595
R28547 VGND.n4485 VGND.n4484 0.00894595
R28548 VGND.n4193 VGND.n4192 0.00894595
R28549 VGND.n4494 VGND.n4493 0.00894595
R28550 VGND.n4586 VGND.n4585 0.00894595
R28551 VGND.n1560 VGND.n1559 0.00894595
R28552 VGND.n1564 VGND.n1563 0.00894595
R28553 VGND.n1460 VGND.n1459 0.00894595
R28554 VGND.n4359 VGND.n4232 0.00894595
R28555 VGND.n4310 VGND.n4309 0.00894595
R28556 VGND.n4352 VGND.n4351 0.00894595
R28557 VGND.n4373 VGND.n4370 0.00894595
R28558 VGND.n3016 VGND.n3013 0.00894595
R28559 VGND.n2990 VGND.n2888 0.00894595
R28560 VGND.n2993 VGND.n2992 0.00894595
R28561 VGND.n2977 VGND.n2976 0.00894595
R28562 VGND.n3580 VGND.n3579 0.00894595
R28563 VGND.n3243 VGND.n3242 0.00894595
R28564 VGND.n3242 VGND.n3238 0.00894595
R28565 VGND.n9080 VGND.n9079 0.00894595
R28566 VGND.n2764 VGND.n2763 0.00894595
R28567 VGND.n3342 VGND.n3339 0.00894595
R28568 VGND.n2132 VGND.n2131 0.00894595
R28569 VGND.n2135 VGND.n2134 0.00894595
R28570 VGND.n3332 VGND.n3331 0.00894595
R28571 VGND.n3177 VGND.n3174 0.00894595
R28572 VGND.n3145 VGND.n3144 0.00894595
R28573 VGND.n3148 VGND.n3147 0.00894595
R28574 VGND.n3184 VGND.n3183 0.00894595
R28575 VGND.n3726 VGND.n3725 0.00894595
R28576 VGND.n9013 VGND.n9012 0.00894595
R28577 VGND.n9012 VGND.n9009 0.00894595
R28578 VGND.n9058 VGND.n9057 0.00894595
R28579 VGND.n9047 VGND.n9046 0.00894595
R28580 VGND.n8820 VGND.n8817 0.00894595
R28581 VGND.n108 VGND.n107 0.00894595
R28582 VGND.n111 VGND.n110 0.00894595
R28583 VGND.n132 VGND.n131 0.00894595
R28584 VGND.n8443 VGND.n256 0.00894595
R28585 VGND.n267 VGND.n266 0.00894595
R28586 VGND.n270 VGND.n269 0.00894595
R28587 VGND.n8528 VGND.n8449 0.00894595
R28588 VGND.n3772 VGND.n3771 0.00894595
R28589 VGND.n8716 VGND.n8715 0.00894595
R28590 VGND.n8715 VGND.n198 0.00894595
R28591 VGND.n8677 VGND.n8676 0.00894595
R28592 VGND.n8708 VGND.n8707 0.00894595
R28593 VGND.n3896 VGND.n3895 0.00894595
R28594 VGND.n139 VGND.n138 0.00894595
R28595 VGND.n142 VGND.n141 0.00894595
R28596 VGND.n8795 VGND.n8789 0.00894595
R28597 VGND.n7978 VGND.n7977 0.00894595
R28598 VGND.n283 VGND.n282 0.00894595
R28599 VGND.n286 VGND.n285 0.00894595
R28600 VGND.n8415 VGND.n8414 0.00894595
R28601 VGND.n1968 VGND.n1967 0.00894595
R28602 VGND.n7913 VGND.n7912 0.00894595
R28603 VGND.n7912 VGND.n7909 0.00894595
R28604 VGND.n469 VGND.n468 0.00894595
R28605 VGND.n8093 VGND.n8092 0.00894595
R28606 VGND.n7724 VGND.n7721 0.00894595
R28607 VGND.n546 VGND.n545 0.00894595
R28608 VGND.n549 VGND.n548 0.00894595
R28609 VGND.n569 VGND.n568 0.00894595
R28610 VGND.n7516 VGND.n687 0.00894595
R28611 VGND.n8216 VGND.n8215 0.00894595
R28612 VGND.n8215 VGND.n458 0.00894595
R28613 VGND.n8206 VGND.n8141 0.00894595
R28614 VGND.n8153 VGND.n8152 0.00894595
R28615 VGND.n8316 VGND.n8313 0.00894595
R28616 VGND.n313 VGND.n312 0.00894595
R28617 VGND.n8328 VGND.n8327 0.00894595
R28618 VGND.n410 VGND.n409 0.00894595
R28619 VGND.n579 VGND.n576 0.00894595
R28620 VGND.n586 VGND.n585 0.00894595
R28621 VGND.n589 VGND.n588 0.00894595
R28622 VGND.n7699 VGND.n7693 0.00894595
R28623 VGND.n1138 VGND.n1135 0.00894595
R28624 VGND.n1138 VGND.n1137 0.00894595
R28625 VGND.n7268 VGND.n7267 0.00894595
R28626 VGND.n1319 VGND.n1318 0.00894595
R28627 VGND.n1202 VGND.n1201 0.00894595
R28628 VGND.n892 VGND.n891 0.00894595
R28629 VGND.n7304 VGND.n7303 0.00894595
R28630 VGND.n989 VGND.n988 0.00894595
R28631 VGND.n801 VGND.n800 0.00894595
R28632 VGND.n7330 VGND.n818 0.00894595
R28633 VGND.n833 VGND.n832 0.00894595
R28634 VGND.n836 VGND.n835 0.00894595
R28635 VGND.n7324 VGND.n7323 0.00894595
R28636 VGND.n6930 VGND.n6929 0.00894595
R28637 VGND.n1545 VGND.n1544 0.00894595
R28638 VGND.n1549 VGND.n1548 0.00894595
R28639 VGND.n6960 VGND.n6959 0.00894595
R28640 VGND.n6217 VGND.n6211 0.00894595
R28641 VGND.n6792 VGND.n6791 0.00894595
R28642 VGND.n6791 VGND.n1597 0.00894595
R28643 VGND.n1608 VGND.n1607 0.00894595
R28644 VGND.n6783 VGND.n1592 0.00894595
R28645 VGND.n6270 VGND.n6269 0.00894595
R28646 VGND.n6483 VGND.n6482 0.00894595
R28647 VGND.n6486 VGND.n6485 0.00894595
R28648 VGND.n6466 VGND.n6463 0.00894595
R28649 VGND.n2239 VGND.n2238 0.00894595
R28650 VGND.n2151 VGND.n2150 0.00894595
R28651 VGND.n2154 VGND.n2153 0.00894595
R28652 VGND.n2628 VGND.n2627 0.00894595
R28653 VGND.n5460 VGND.n5457 0.00894595
R28654 VGND.n5292 VGND.n5291 0.00894595
R28655 VGND.n5328 VGND.n5327 0.00894595
R28656 VGND.n5288 VGND.n5221 0.00894595
R28657 VGND.n5751 VGND.n5750 0.00894595
R28658 VGND.n5779 VGND.n5778 0.00894595
R28659 VGND.n5783 VGND.n5782 0.00894595
R28660 VGND.n5794 VGND.n5793 0.00894595
R28661 VGND.n2398 VGND.n2397 0.00894595
R28662 VGND.n34 VGND.n33 0.00894595
R28663 VGND.n9098 VGND.n9097 0.00894595
R28664 VGND.n5611 VGND.n5607 0.00894595
R28665 VGND.n5611 VGND.n5610 0.00894595
R28666 VGND.n5616 VGND.n5471 0.00894595
R28667 VGND.n2542 VGND.n2541 0.00894595
R28668 VGND.n2541 VGND.n2320 0.00894595
R28669 VGND.n2532 VGND.n2531 0.00894595
R28670 VGND.n2515 VGND.n2514 0.00894595
R28671 VGND.n9209 VGND.n9208 0.00894595
R28672 VGND.n5829 VGND.n5824 0.00894595
R28673 VGND.n5826 VGND.n5825 0.00894595
R28674 VGND.n5838 VGND.n5837 0.00894595
R28675 VGND.n5859 VGND.n5856 0.00894595
R28676 VGND.n7293 VGND.n7292 0.00837842
R28677 VGND.n6198 VGND.n6197 0.00837842
R28678 VGND.n6203 VGND.n6202 0.00837842
R28679 VGND.n6200 VGND.n6199 0.00837842
R28680 VGND.n4964 VGND.n4963 0.0083125
R28681 VGND.n4972 VGND.n4971 0.0083125
R28682 VGND.n4975 VGND.n4974 0.0083125
R28683 VGND.n5014 VGND.n5013 0.0083125
R28684 VGND.n7216 VGND.n7215 0.0083125
R28685 VGND.n7221 VGND.n7220 0.0083125
R28686 VGND.n7084 VGND.n7083 0.0083125
R28687 VGND.n7081 VGND.n7080 0.0083125
R28688 VGND.n7002 VGND.n1370 0.0083125
R28689 VGND.n4305 VGND.n4304 0.0083125
R28690 VGND.n4320 VGND.n4308 0.0083125
R28691 VGND VGND.n4318 0.0083125
R28692 VGND.n4379 VGND.n4378 0.0083125
R28693 VGND.n4507 VGND.n4506 0.0083125
R28694 VGND.n4513 VGND.n4512 0.0083125
R28695 VGND.n1471 VGND.n1470 0.0083125
R28696 VGND.n1468 VGND.n1467 0.0083125
R28697 VGND.n3381 VGND.n3379 0.0083125
R28698 VGND.n3372 VGND.n3370 0.0083125
R28699 VGND.n3366 VGND.n3364 0.0083125
R28700 VGND.n3326 VGND.n3325 0.0083125
R28701 VGND.n2770 VGND.n2765 0.0083125
R28702 VGND.n2775 VGND.n2774 0.0083125
R28703 VGND.n2988 VGND.n2987 0.0083125
R28704 VGND.n2985 VGND.n2984 0.0083125
R28705 VGND.n8859 VGND.n8857 0.0083125
R28706 VGND.n8850 VGND.n8848 0.0083125
R28707 VGND.n8844 VGND.n8842 0.0083125
R28708 VGND.n8913 VGND.n8912 0.0083125
R28709 VGND.n9036 VGND.n9035 0.0083125
R28710 VGND.n9044 VGND.n9043 0.0083125
R28711 VGND.n3196 VGND.n3195 0.0083125
R28712 VGND.n3193 VGND.n3192 0.0083125
R28713 VGND.n3918 VGND.n3916 0.0083125
R28714 VGND.n3909 VGND.n3907 0.0083125
R28715 VGND.n3903 VGND.n3901 0.0083125
R28716 VGND.n160 VGND.n157 0.0083125
R28717 VGND.n8697 VGND.n8696 0.0083125
R28718 VGND.n8705 VGND.n8704 0.0083125
R28719 VGND.n8543 VGND.n8542 0.0083125
R28720 VGND.n8540 VGND.n8539 0.0083125
R28721 VGND.n8450 VGND.n271 0.0083125
R28722 VGND.n7760 VGND.n7759 0.0083125
R28723 VGND.n7752 VGND.n7751 0.0083125
R28724 VGND.n7749 VGND.n7747 0.0083125
R28725 VGND.n7818 VGND.n7817 0.0083125
R28726 VGND.n8083 VGND.n8082 0.0083125
R28727 VGND.n8090 VGND.n8089 0.0083125
R28728 VGND.n8425 VGND.n8424 0.0083125
R28729 VGND.n8422 VGND.n8421 0.0083125
R28730 VGND.n7633 VGND.n7631 0.0083125
R28731 VGND.n7624 VGND.n7622 0.0083125
R28732 VGND.n7618 VGND.n7615 0.0083125
R28733 VGND.n682 VGND.n681 0.0083125
R28734 VGND.n8198 VGND.n8197 0.0083125
R28735 VGND.n8195 VGND.n8194 0.0083125
R28736 VGND.n8330 VGND.n310 0.0083125
R28737 VGND.n326 VGND.n325 0.0083125
R28738 VGND.n407 VGND.n406 0.0083125
R28739 VGND.n7428 VGND.n787 0.0083125
R28740 VGND.n7340 VGND.n7335 0.0083125
R28741 VGND.n869 VGND.n868 0.0083125
R28742 VGND.n1019 VGND.n885 0.0083125
R28743 VGND.n1308 VGND.n1307 0.0083125
R28744 VGND.n1316 VGND.n1315 0.0083125
R28745 VGND.n7306 VGND.n890 0.0083125
R28746 VGND.n980 VGND.n979 0.0083125
R28747 VGND.n6216 VGND.n6214 0.0083125
R28748 VGND.n6276 VGND.n6275 0.0083125
R28749 VGND.n1679 VGND.n1678 0.0083125
R28750 VGND.n6340 VGND.n1687 0.0083125
R28751 VGND.n6814 VGND.n6813 0.0083125
R28752 VGND.n6818 VGND.n6817 0.0083125
R28753 VGND.n6971 VGND.n6970 0.0083125
R28754 VGND.n6968 VGND.n6967 0.0083125
R28755 VGND.n6055 VGND.n1767 0.0083125
R28756 VGND.n6574 VGND.n6573 0.0083125
R28757 VGND.n6566 VGND.n6562 0.0083125
R28758 VGND.n6558 VGND.n6556 0.0083125
R28759 VGND.n6634 VGND.n6633 0.0083125
R28760 VGND.n5357 VGND.n5356 0.0083125
R28761 VGND.n5367 VGND.n5366 0.0083125
R28762 VGND.n5331 VGND.n5330 0.0083125
R28763 VGND.n5334 VGND.n5333 0.0083125
R28764 VGND.n5222 VGND.n5211 0.0083125
R28765 VGND.n5974 VGND 0.0083125
R28766 VGND VGND.n5973 0.0083125
R28767 VGND.n5891 VGND.n5890 0.0083125
R28768 VGND.n5883 VGND.n5881 0.0083125
R28769 VGND.n5877 VGND.n5875 0.0083125
R28770 VGND.n5499 VGND.n5122 0.0083125
R28771 VGND.n5633 VGND.n5632 0.0083125
R28772 VGND.n5638 VGND.n5637 0.0083125
R28773 VGND.n5806 VGND.n5805 0.0083125
R28774 VGND.n5803 VGND.n5802 0.0083125
R28775 VGND.n9213 VGND 0.0083125
R28776 VGND VGND.n9212 0.0083125
R28777 VGND.n2245 VGND.n2244 0.0083125
R28778 VGND.n2255 VGND.n2253 0.0083125
R28779 VGND.n2260 VGND.n2259 0.0083125
R28780 VGND.n2622 VGND.n2621 0.0083125
R28781 VGND.n2507 VGND.n2506 0.0083125
R28782 VGND.n2512 VGND.n2511 0.0083125
R28783 VGND.n9173 VGND.n9172 0.0083125
R28784 VGND.n9170 VGND.n9169 0.0083125
R28785 VGND.n7296 VGND.n7295 0.00803709
R28786 VGND.n1000 VGND.n999 0.00803709
R28787 VGND.n1002 VGND.n1001 0.00762121
R28788 VGND.n899 VGND.n898 0.00762121
R28789 VGND.n798 VGND.n797 0.00762121
R28790 VGND.n820 VGND.n819 0.00762121
R28791 VGND.n4365 VGND.n4364 0.00735251
R28792 VGND.n1571 VGND.n1570 0.00735251
R28793 VGND.n4181 VGND.n4180 0.00735251
R28794 VGND.n4704 VGND.n4703 0.00735251
R28795 VGND.n1782 VGND.n1781 0.00725676
R28796 VGND.n1755 VGND.n1754 0.00725676
R28797 VGND.n5090 VGND.n5089 0.00725676
R28798 VGND.n4816 VGND.n4815 0.00725676
R28799 VGND.n4136 VGND.n4135 0.00725676
R28800 VGND.n2890 VGND.n2889 0.00725676
R28801 VGND.n2085 VGND.n2084 0.00725676
R28802 VGND.n3138 VGND.n3137 0.00725676
R28803 VGND.n3614 VGND.n3613 0.00725676
R28804 VGND.n8556 VGND.n8555 0.00725676
R28805 VGND.n3760 VGND.n3759 0.00725676
R28806 VGND.n301 VGND.n300 0.00725676
R28807 VGND.n1996 VGND.n1995 0.00725676
R28808 VGND.n7525 VGND.n7524 0.00725676
R28809 VGND.n1169 VGND.n1168 0.00725676
R28810 VGND.n7495 VGND.n7494 0.00725676
R28811 VGND.n1580 VGND.n1579 0.00725676
R28812 VGND.n6157 VGND.n6156 0.00725676
R28813 VGND.n5306 VGND.n5305 0.00725676
R28814 VGND.n5777 VGND.n5776 0.00725676
R28815 VGND.n2363 VGND.n2362 0.00725676
R28816 VGND.n3477 VGND.n3476 0.00725676
R28817 VGND VGND.n4800 0.00701042
R28818 VGND.n4853 VGND.n4850 0.00701042
R28819 VGND.n4968 VGND.n4967 0.00701042
R28820 VGND.n4971 VGND.n4970 0.00701042
R28821 VGND.n7211 VGND.n7209 0.00701042
R28822 VGND.n5095 VGND.n5094 0.00701042
R28823 VGND.n5094 VGND 0.00701042
R28824 VGND.n7083 VGND.n7082 0.00701042
R28825 VGND VGND.n7074 0.00701042
R28826 VGND VGND.n4158 0.00701042
R28827 VGND.n4159 VGND 0.00701042
R28828 VGND.n4726 VGND.n4724 0.00701042
R28829 VGND.n4356 VGND.n4355 0.00701042
R28830 VGND.n4353 VGND.n4308 0.00701042
R28831 VGND.n4502 VGND.n4500 0.00701042
R28832 VGND.n1473 VGND.n1472 0.00701042
R28833 VGND.n1472 VGND 0.00701042
R28834 VGND.n1470 VGND.n1469 0.00701042
R28835 VGND.n3565 VGND.n3564 0.00701042
R28836 VGND.n3376 VGND.n3375 0.00701042
R28837 VGND.n3373 VGND.n3372 0.00701042
R28838 VGND.n3226 VGND.n52 0.00701042
R28839 VGND.n9077 VGND 0.00701042
R28840 VGND.n2989 VGND 0.00701042
R28841 VGND.n2987 VGND.n2986 0.00701042
R28842 VGND.n8854 VGND.n8853 0.00701042
R28843 VGND.n8851 VGND.n8850 0.00701042
R28844 VGND.n9031 VGND.n9029 0.00701042
R28845 VGND.n3198 VGND.n3197 0.00701042
R28846 VGND.n3197 VGND 0.00701042
R28847 VGND.n3195 VGND.n3194 0.00701042
R28848 VGND.n3831 VGND.n3829 0.00701042
R28849 VGND.n3913 VGND.n3912 0.00701042
R28850 VGND.n3910 VGND.n3909 0.00701042
R28851 VGND.n8664 VGND.n8662 0.00701042
R28852 VGND VGND.n8679 0.00701042
R28853 VGND.n303 VGND.n302 0.00701042
R28854 VGND.n302 VGND 0.00701042
R28855 VGND.n8542 VGND.n8541 0.00701042
R28856 VGND.n8530 VGND 0.00701042
R28857 VGND.n1918 VGND 0.00701042
R28858 VGND.n7756 VGND.n7755 0.00701042
R28859 VGND.n7753 VGND.n7752 0.00701042
R28860 VGND.n8078 VGND.n8076 0.00701042
R28861 VGND.n8427 VGND.n8426 0.00701042
R28862 VGND.n8426 VGND 0.00701042
R28863 VGND.n8424 VGND.n8423 0.00701042
R28864 VGND.n7552 VGND.n7550 0.00701042
R28865 VGND.n7628 VGND.n7627 0.00701042
R28866 VGND.n7625 VGND.n7624 0.00701042
R28867 VGND.n8205 VGND.n8203 0.00701042
R28868 VGND.n8332 VGND.n8331 0.00701042
R28869 VGND.n8331 VGND 0.00701042
R28870 VGND.n324 VGND.n310 0.00701042
R28871 VGND.n408 VGND 0.00701042
R28872 VGND.n7439 VGND.n7437 0.00701042
R28873 VGND.n862 VGND.n861 0.00701042
R28874 VGND.n865 VGND.n864 0.00701042
R28875 VGND.n1303 VGND.n1302 0.00701042
R28876 VGND.n7308 VGND.n7307 0.00701042
R28877 VGND.n7307 VGND 0.00701042
R28878 VGND.n978 VGND.n890 0.00701042
R28879 VGND VGND.n986 0.00701042
R28880 VGND.n6112 VGND 0.00701042
R28881 VGND VGND.n6100 0.00701042
R28882 VGND.n6182 VGND.n6180 0.00701042
R28883 VGND.n1676 VGND.n1675 0.00701042
R28884 VGND.n6809 VGND.n6807 0.00701042
R28885 VGND.n6973 VGND.n6972 0.00701042
R28886 VGND.n6972 VGND 0.00701042
R28887 VGND.n6970 VGND.n6969 0.00701042
R28888 VGND.n6065 VGND.n6063 0.00701042
R28889 VGND.n6570 VGND.n6569 0.00701042
R28890 VGND.n6567 VGND.n6566 0.00701042
R28891 VGND.n5352 VGND.n5351 0.00701042
R28892 VGND.n5312 VGND.n5311 0.00701042
R28893 VGND.n5311 VGND 0.00701042
R28894 VGND.n5332 VGND.n5331 0.00701042
R28895 VGND.n5290 VGND 0.00701042
R28896 VGND VGND.n5289 0.00701042
R28897 VGND.n5994 VGND.n5992 0.00701042
R28898 VGND.n5887 VGND.n5886 0.00701042
R28899 VGND.n5884 VGND.n5883 0.00701042
R28900 VGND.n5592 VGND.n5590 0.00701042
R28901 VGND.n5808 VGND.n5807 0.00701042
R28902 VGND.n5807 VGND 0.00701042
R28903 VGND.n5805 VGND.n5804 0.00701042
R28904 VGND.n2249 VGND.n2248 0.00701042
R28905 VGND.n2253 VGND.n2251 0.00701042
R28906 VGND.n2502 VGND.n2500 0.00701042
R28907 VGND.n9175 VGND.n9174 0.00701042
R28908 VGND.n9174 VGND 0.00701042
R28909 VGND.n9172 VGND.n9171 0.00701042
R28910 VGND.n6197 VGND.n6196 0.00696227
R28911 VGND.n7292 VGND.n829 0.00657697
R28912 VGND.n7295 VGND.n7294 0.00657697
R28913 VGND.n7297 VGND.n1000 0.00657697
R28914 VGND.n6204 VGND.n6203 0.00657697
R28915 VGND.n6201 VGND.n6200 0.00657697
R28916 VGND.n6956 VGND.n1541 0.00648266
R28917 VGND.n6208 VGND.n1695 0.00648266
R28918 VGND.n6789 VGND.n6788 0.00648266
R28919 VGND.n6786 VGND.n6785 0.00648266
R28920 VGND.n1663 VGND.n1662 0.00648266
R28921 VGND.n6742 VGND.n6741 0.00619697
R28922 VGND.n6760 VGND.n6746 0.00619697
R28923 VGND.n6088 VGND.n6087 0.00619697
R28924 VGND.n6083 VGND.n6082 0.00619697
R28925 VGND.n7093 VGND.n7092 0.00619697
R28926 VGND.n7088 VGND.n7087 0.00619697
R28927 VGND.n7251 VGND.n7241 0.00619697
R28928 VGND.n7237 VGND.n7236 0.00619697
R28929 VGND.n4838 VGND.n4837 0.00619697
R28930 VGND.n4833 VGND.n4832 0.00619697
R28931 VGND.n5000 VGND.n4999 0.00619697
R28932 VGND.n4995 VGND.n4994 0.00619697
R28933 VGND.n4749 VGND.n4748 0.00619697
R28934 VGND.n4744 VGND.n4743 0.00619697
R28935 VGND.n4208 VGND.n4207 0.00619697
R28936 VGND.n4203 VGND.n4202 0.00619697
R28937 VGND.n6987 VGND.n1383 0.00619697
R28938 VGND.n1567 VGND.n1555 0.00619697
R28939 VGND.n4349 VGND.n4348 0.00619697
R28940 VGND.n4344 VGND.n4343 0.00619697
R28941 VGND.n3002 VGND.n3001 0.00619697
R28942 VGND.n2997 VGND.n2996 0.00619697
R28943 VGND.n3554 VGND.n3553 0.00619697
R28944 VGND.n3549 VGND.n3548 0.00619697
R28945 VGND.n9086 VGND.n9085 0.00619697
R28946 VGND.n9071 VGND.n56 0.00619697
R28947 VGND.n3348 VGND.n3347 0.00619697
R28948 VGND.n3353 VGND.n3352 0.00619697
R28949 VGND.n3157 VGND.n3156 0.00619697
R28950 VGND.n3152 VGND.n3151 0.00619697
R28951 VGND.n3610 VGND.n3609 0.00619697
R28952 VGND.n3605 VGND.n3604 0.00619697
R28953 VGND.n9064 VGND.n9063 0.00619697
R28954 VGND.n71 VGND.n59 0.00619697
R28955 VGND.n8826 VGND.n8825 0.00619697
R28956 VGND.n8831 VGND.n8830 0.00619697
R28957 VGND.n8552 VGND.n8551 0.00619697
R28958 VGND.n8547 VGND.n8546 0.00619697
R28959 VGND.n3756 VGND.n3755 0.00619697
R28960 VGND.n3751 VGND.n3750 0.00619697
R28961 VGND.n8673 VGND.n8672 0.00619697
R28962 VGND.n8691 VGND.n8688 0.00619697
R28963 VGND.n8810 VGND.n8809 0.00619697
R28964 VGND.n8805 VGND.n8804 0.00619697
R28965 VGND.n8434 VGND.n294 0.00619697
R28966 VGND.n290 VGND.n289 0.00619697
R28967 VGND.n2029 VGND.n2028 0.00619697
R28968 VGND.n2024 VGND.n2023 0.00619697
R28969 VGND.n475 VGND.n474 0.00619697
R28970 VGND.n8110 VGND.n8098 0.00619697
R28971 VGND.n7730 VGND.n7729 0.00619697
R28972 VGND.n7735 VGND.n7734 0.00619697
R28973 VGND.n747 VGND.n746 0.00619697
R28974 VGND.n742 VGND.n741 0.00619697
R28975 VGND.n8209 VGND.n8127 0.00619697
R28976 VGND.n8123 VGND.n8122 0.00619697
R28977 VGND.n426 VGND.n425 0.00619697
R28978 VGND.n8324 VGND.n316 0.00619697
R28979 VGND.n7714 VGND.n7713 0.00619697
R28980 VGND.n7709 VGND.n7708 0.00619697
R28981 VGND.n7271 VGND.n7262 0.00619697
R28982 VGND.n7290 VGND.n7279 0.00619697
R28983 VGND.n1180 VGND.n1179 0.00619697
R28984 VGND.n7300 VGND.n894 0.00619697
R28985 VGND.n7449 VGND.n772 0.00619697
R28986 VGND.n764 VGND.n753 0.00619697
R28987 VGND.n841 VGND.n831 0.00619697
R28988 VGND.n859 VGND.n855 0.00619697
R28989 VGND.n6953 VGND.n6952 0.00619697
R28990 VGND.n1553 VGND.n1543 0.00619697
R28991 VGND.n6166 VGND.n6165 0.00619697
R28992 VGND.n6194 VGND.n6095 0.00619697
R28993 VGND.n1611 VGND.n1603 0.00619697
R28994 VGND.n6779 VGND.n6766 0.00619697
R28995 VGND.n6491 VGND.n6481 0.00619697
R28996 VGND.n6475 VGND.n1666 0.00619697
R28997 VGND.n5844 VGND.n5843 0.00619697
R28998 VGND.n5851 VGND.n5848 0.00619697
R28999 VGND.n2161 VGND.n2149 0.00619697
R29000 VGND.n6537 VGND.n6536 0.00619697
R29001 VGND.n6542 VGND.n6541 0.00619697
R29002 VGND.n5320 VGND.n5319 0.00619697
R29003 VGND.n5325 VGND.n5324 0.00619697
R29004 VGND.n5771 VGND.n5770 0.00619697
R29005 VGND.n5788 VGND.n5775 0.00619697
R29006 VGND.n2376 VGND.n2375 0.00619697
R29007 VGND.n5484 VGND.n5483 0.00619697
R29008 VGND.n5623 VGND.n5488 0.00619697
R29009 VGND.n2535 VGND.n2525 0.00619697
R29010 VGND.n3533 VGND.n3474 0.00619697
R29011 VGND.n9225 VGND.n9219 0.00619697
R29012 VGND.n6004 VGND.n1791 0.00619697
R29013 VGND.n5983 VGND.n5982 0.00619697
R29014 VGND.n6954 VGND.n1571 0.00590801
R29015 VGND.n6195 VGND.n6092 0.00590801
R29016 VGND.n4814 VGND.n4813 0.00570833
R29017 VGND.n4011 VGND.n4008 0.00570833
R29018 VGND.n5096 VGND.n5093 0.00570833
R29019 VGND.n4134 VGND.n4133 0.00570833
R29020 VGND.n4480 VGND.n4213 0.00570833
R29021 VGND.n6982 VGND.n6981 0.00570833
R29022 VGND.n2083 VGND.n2082 0.00570833
R29023 VGND.n3460 VGND 0.00570833
R29024 VGND.n2894 VGND.n2893 0.00570833
R29025 VGND.n3702 VGND.n3701 0.00570833
R29026 VGND.n9020 VGND.n9018 0.00570833
R29027 VGND VGND.n9022 0.00570833
R29028 VGND.n3199 VGND.n2665 0.00570833
R29029 VGND.n3814 VGND.n3813 0.00570833
R29030 VGND.n8653 VGND.n196 0.00570833
R29031 VGND.n304 VGND.n257 0.00570833
R29032 VGND.n1994 VGND.n1993 0.00570833
R29033 VGND.n7919 VGND.n7918 0.00570833
R29034 VGND.n8429 VGND.n8428 0.00570833
R29035 VGND.n7531 VGND.n7530 0.00570833
R29036 VGND.n8129 VGND.n456 0.00570833
R29037 VGND VGND.n8131 0.00570833
R29038 VGND.n8333 VGND.n309 0.00570833
R29039 VGND.n7493 VGND.n7492 0.00570833
R29040 VGND VGND.n786 0.00570833
R29041 VGND.n1133 VGND.n1130 0.00570833
R29042 VGND.n7309 VGND.n889 0.00570833
R29043 VGND.n6155 VGND.n6154 0.00570833
R29044 VGND.n6798 VGND.n6795 0.00570833
R29045 VGND.n6974 VGND.n1476 0.00570833
R29046 VGND.n1757 VGND.n1756 0.00570833
R29047 VGND.n6726 VGND.n6723 0.00570833
R29048 VGND.n5314 VGND.n5313 0.00570833
R29049 VGND.n1835 VGND.n1834 0.00570833
R29050 VGND.n5605 VGND.n5602 0.00570833
R29051 VGND.n5809 VGND.n5126 0.00570833
R29052 VGND.n3519 VGND.n3518 0.00570833
R29053 VGND.n3526 VGND 0.00570833
R29054 VGND.n2318 VGND.n2317 0.00570833
R29055 VGND.n9176 VGND.n21 0.00570833
R29056 VGND.n6206 VGND.n6205 0.005649
R29057 VGND.n1781 VGND.n1780 0.00556757
R29058 VGND.n6003 VGND.n1796 0.00556757
R29059 VGND.n1755 VGND.n1747 0.00556757
R29060 VGND.n6074 VGND.n1704 0.00556757
R29061 VGND.n6016 VGND.n6015 0.00556757
R29062 VGND.n6498 VGND.n6497 0.00556757
R29063 VGND.n6519 VGND.n6511 0.00556757
R29064 VGND.n7073 VGND.n7072 0.00556757
R29065 VGND.n4815 VGND.n4764 0.00556757
R29066 VGND.n4839 VGND.n4091 0.00556757
R29067 VGND.n4050 VGND.n4049 0.00556757
R29068 VGND.n5008 VGND.n5007 0.00556757
R29069 VGND.n4135 VGND.n4096 0.00556757
R29070 VGND.n4735 VGND.n4146 0.00556757
R29071 VGND.n4299 VGND.n4232 0.00556757
R29072 VGND.n4373 VGND.n4372 0.00556757
R29073 VGND.n2084 VGND.n2040 0.00556757
R29074 VGND.n3555 VGND.n3463 0.00556757
R29075 VGND.n3339 VGND.n3338 0.00556757
R29076 VGND.n3331 VGND.n2641 0.00556757
R29077 VGND.n3613 VGND.n3612 0.00556757
R29078 VGND.n3596 VGND.n3591 0.00556757
R29079 VGND.n8817 VGND.n8816 0.00556757
R29080 VGND.n131 VGND.n126 0.00556757
R29081 VGND.n8528 VGND.n8527 0.00556757
R29082 VGND.n3759 VGND.n3758 0.00556757
R29083 VGND.n3742 VGND.n3737 0.00556757
R29084 VGND.n3897 VGND.n3896 0.00556757
R29085 VGND.n8789 VGND.n155 0.00556757
R29086 VGND.n1995 VGND.n1876 0.00556757
R29087 VGND.n2015 VGND.n2010 0.00556757
R29088 VGND.n7721 VGND.n7720 0.00556757
R29089 VGND.n568 VGND.n562 0.00556757
R29090 VGND.n7526 VGND.n7525 0.00556757
R29091 VGND.n733 VGND.n728 0.00556757
R29092 VGND.n409 VGND.n323 0.00556757
R29093 VGND.n576 VGND.n575 0.00556757
R29094 VGND.n7693 VGND.n604 0.00556757
R29095 VGND.n7494 VGND.n7452 0.00556757
R29096 VGND.n7448 VGND.n773 0.00556757
R29097 VGND.n759 VGND.n758 0.00556757
R29098 VGND.n802 VGND.n801 0.00556757
R29099 VGND.n818 VGND.n817 0.00556757
R29100 VGND.n7323 VGND.n847 0.00556757
R29101 VGND.n6156 VGND.n6116 0.00556757
R29102 VGND.n6167 VGND.n6114 0.00556757
R29103 VGND.n6099 VGND.n6098 0.00556757
R29104 VGND.n6218 VGND.n6217 0.00556757
R29105 VGND.n6271 VGND.n6270 0.00556757
R29106 VGND.n6466 VGND.n6465 0.00556757
R29107 VGND.n2240 VGND.n2239 0.00556757
R29108 VGND.n2627 VGND.n2168 0.00556757
R29109 VGND.n5288 VGND.n5287 0.00556757
R29110 VGND.n3476 VGND.n3475 0.00556757
R29111 VGND.n3532 VGND.n3529 0.00556757
R29112 VGND.n9204 VGND.n2 0.00556757
R29113 VGND.n5824 VGND.n5114 0.00556757
R29114 VGND.n5859 VGND.n5858 0.00556757
R29115 VGND.n4703 VGND.n1696 0.00554564
R29116 VGND.n6780 VGND.n6764 0.00500002
R29117 VGND.n4180 VGND.n1612 0.00500002
R29118 VGND.n6493 VGND.n6492 0.00495986
R29119 VGND.n6219 VGND 0.00490236
R29120 VGND.n4056 VGND.n842 0.00482801
R29121 VGND.n1361 VGND.n895 0.00482801
R29122 VGND.n7272 VGND.n7255 0.00482801
R29123 VGND.n7450 VGND.n765 0.00482801
R29124 VGND.n1321 VGND.n1142 0.00477273
R29125 VGND.n991 VGND.n897 0.00477273
R29126 VGND.n751 VGND.n750 0.00477273
R29127 VGND.n7328 VGND.n822 0.00477273
R29128 VGND.n6927 VGND.n6926 0.00477273
R29129 VGND.n6161 VGND.n6160 0.00477273
R29130 VGND.n2162 VGND.n2142 0.00460158
R29131 VGND.n3346 VGND.n2633 0.00460158
R29132 VGND.n8824 VGND.n118 0.00460158
R29133 VGND.n8812 VGND.n8811 0.00460158
R29134 VGND.n7728 VGND.n556 0.00460158
R29135 VGND.n7716 VGND.n7715 0.00460158
R29136 VGND.n5001 VGND.n4058 0.00460158
R29137 VGND.n4231 VGND.n4230 0.00460158
R29138 VGND.n5852 VGND.n5835 0.00460158
R29139 VGND.n2370 VGND.n2369 0.00460158
R29140 VGND.n5789 VGND.n5464 0.00460158
R29141 VGND.n2536 VGND.n2518 0.00460158
R29142 VGND.n9088 VGND.n9087 0.00460158
R29143 VGND.n9066 VGND.n9065 0.00460158
R29144 VGND.n203 VGND.n202 0.00460158
R29145 VGND.n2033 VGND.n476 0.00460158
R29146 VGND.n8210 VGND.n8113 0.00460158
R29147 VGND.n4209 VGND.n4184 0.00460158
R29148 VGND.n5620 VGND.n5489 0.00460158
R29149 VGND.n3534 VGND.n3466 0.00460158
R29150 VGND.n3540 VGND.n3539 0.00460158
R29151 VGND.n3611 VGND.n3584 0.00460158
R29152 VGND.n3757 VGND.n3730 0.00460158
R29153 VGND.n2031 VGND.n2030 0.00460158
R29154 VGND.n1873 VGND.n748 0.00460158
R29155 VGND.n4824 VGND.n4095 0.00460158
R29156 VGND.n4751 VGND.n4750 0.00460158
R29157 VGND.n6090 VGND.n6089 0.00460158
R29158 VGND.n4814 VGND.n4801 0.00440625
R29159 VGND.n4858 VGND.n4857 0.00440625
R29160 VGND.n4965 VGND.n4964 0.00440625
R29161 VGND.n4991 VGND.n4981 0.00440625
R29162 VGND.n4990 VGND 0.00440625
R29163 VGND.n5010 VGND.n5009 0.00440625
R29164 VGND.n7198 VGND.n7196 0.00440625
R29165 VGND.n7084 VGND 0.00440625
R29166 VGND.n7074 VGND.n1370 0.00440625
R29167 VGND.n4134 VGND.n4131 0.00440625
R29168 VGND.n4722 VGND 0.00440625
R29169 VGND.n4719 VGND.n4718 0.00440625
R29170 VGND.n4306 VGND.n4305 0.00440625
R29171 VGND VGND.n4329 0.00440625
R29172 VGND.n4340 VGND.n4334 0.00440625
R29173 VGND VGND.n4338 0.00440625
R29174 VGND.n4375 VGND.n4374 0.00440625
R29175 VGND.n4520 VGND.n4519 0.00440625
R29176 VGND VGND.n1471 0.00440625
R29177 VGND.n2083 VGND.n2080 0.00440625
R29178 VGND.n3569 VGND.n3568 0.00440625
R29179 VGND.n3379 VGND.n3378 0.00440625
R29180 VGND.n3358 VGND.n3357 0.00440625
R29181 VGND VGND.n2126 0.00440625
R29182 VGND.n3330 VGND.n3329 0.00440625
R29183 VGND.n2782 VGND.n2780 0.00440625
R29184 VGND.n2989 VGND 0.00440625
R29185 VGND VGND.n2988 0.00440625
R29186 VGND.n3701 VGND.n3700 0.00440625
R29187 VGND.n3721 VGND.n3720 0.00440625
R29188 VGND.n8857 VGND.n8856 0.00440625
R29189 VGND.n8836 VGND.n8835 0.00440625
R29190 VGND VGND.n102 0.00440625
R29191 VGND.n130 VGND.n129 0.00440625
R29192 VGND.n3040 VGND.n3039 0.00440625
R29193 VGND VGND.n3196 0.00440625
R29194 VGND.n3813 VGND.n3812 0.00440625
R29195 VGND.n3836 VGND.n3835 0.00440625
R29196 VGND.n3916 VGND.n3915 0.00440625
R29197 VGND VGND.n8799 0.00440625
R29198 VGND.n8788 VGND.n8787 0.00440625
R29199 VGND.n8650 VGND.n8649 0.00440625
R29200 VGND.n8543 VGND 0.00440625
R29201 VGND.n8529 VGND.n271 0.00440625
R29202 VGND.n1994 VGND.n1918 0.00440625
R29203 VGND.n1974 VGND.n1973 0.00440625
R29204 VGND.n7759 VGND.n7758 0.00440625
R29205 VGND.n7740 VGND.n7739 0.00440625
R29206 VGND VGND.n540 0.00440625
R29207 VGND.n567 VGND.n507 0.00440625
R29208 VGND.n8067 VGND.n8065 0.00440625
R29209 VGND VGND.n8425 0.00440625
R29210 VGND.n7530 VGND.n7529 0.00440625
R29211 VGND.n7557 VGND.n7556 0.00440625
R29212 VGND.n7631 VGND.n7630 0.00440625
R29213 VGND.n7705 VGND.n599 0.00440625
R29214 VGND.n7704 VGND 0.00440625
R29215 VGND.n7692 VGND.n7691 0.00440625
R29216 VGND.n8191 VGND.n8189 0.00440625
R29217 VGND VGND.n8330 0.00440625
R29218 VGND.n408 VGND.n407 0.00440625
R29219 VGND.n7493 VGND.n7491 0.00440625
R29220 VGND.n7431 VGND.n7430 0.00440625
R29221 VGND.n794 VGND.n787 0.00440625
R29222 VGND.n7335 VGND.n7334 0.00440625
R29223 VGND.n879 VGND.n876 0.00440625
R29224 VGND.n883 VGND 0.00440625
R29225 VGND.n7322 VGND.n7321 0.00440625
R29226 VGND.n1296 VGND.n1295 0.00440625
R29227 VGND VGND.n7306 0.00440625
R29228 VGND.n6155 VGND.n6153 0.00440625
R29229 VGND VGND.n6184 0.00440625
R29230 VGND.n6187 VGND.n6186 0.00440625
R29231 VGND.n6216 VGND.n6215 0.00440625
R29232 VGND.n6275 VGND.n6274 0.00440625
R29233 VGND VGND.n1684 0.00440625
R29234 VGND.n6467 VGND.n6458 0.00440625
R29235 VGND.n6825 VGND.n6824 0.00440625
R29236 VGND VGND.n6971 0.00440625
R29237 VGND.n1756 VGND.n1705 0.00440625
R29238 VGND.n6058 VGND.n6057 0.00440625
R29239 VGND.n1771 VGND.n1767 0.00440625
R29240 VGND.n6573 VGND.n6572 0.00440625
R29241 VGND.n6550 VGND.n6548 0.00440625
R29242 VGND VGND.n1654 0.00440625
R29243 VGND.n6518 VGND.n6517 0.00440625
R29244 VGND.n5372 VGND.n5370 0.00440625
R29245 VGND.n5330 VGND 0.00440625
R29246 VGND.n5289 VGND.n5211 0.00440625
R29247 VGND.n1834 VGND.n1833 0.00440625
R29248 VGND.n5990 VGND 0.00440625
R29249 VGND.n5975 VGND.n5974 0.00440625
R29250 VGND.n5890 VGND.n5889 0.00440625
R29251 VGND.n5869 VGND.n5867 0.00440625
R29252 VGND.n5862 VGND 0.00440625
R29253 VGND.n5860 VGND.n5818 0.00440625
R29254 VGND.n5645 VGND.n5643 0.00440625
R29255 VGND VGND.n5806 0.00440625
R29256 VGND.n3518 VGND.n3517 0.00440625
R29257 VGND VGND.n6 0.00440625
R29258 VGND.n9214 VGND.n9213 0.00440625
R29259 VGND.n2246 VGND.n2245 0.00440625
R29260 VGND.n2277 VGND.n2266 0.00440625
R29261 VGND VGND.n2278 0.00440625
R29262 VGND.n2282 VGND 0.00440625
R29263 VGND.n2626 VGND.n2625 0.00440625
R29264 VGND.n2492 VGND.n2487 0.00440625
R29265 VGND VGND.n9173 0.00440625
R29266 VGND.n6734 VGND.n1615 0.00406061
R29267 VGND.n6013 VGND.n6012 0.00406061
R29268 VGND.n6996 VGND.n6991 0.00406061
R29269 VGND.n4001 VGND.n3999 0.00406061
R29270 VGND.n4762 VGND.n4756 0.00406061
R29271 VGND.n4054 VGND.n4047 0.00406061
R29272 VGND.n4708 VGND.n4707 0.00406061
R29273 VGND.n4492 VGND.n4491 0.00406061
R29274 VGND.n4369 VGND.n4368 0.00406061
R29275 VGND.n3017 VGND.n2745 0.00406061
R29276 VGND.n3581 VGND.n2096 0.00406061
R29277 VGND.n3343 VGND.n3336 0.00406061
R29278 VGND.n3178 VGND.n3024 0.00406061
R29279 VGND.n3727 VGND.n3625 0.00406061
R29280 VGND.n8821 VGND.n8814 0.00406061
R29281 VGND.n8444 VGND.n8439 0.00406061
R29282 VGND.n3770 VGND.n3769 0.00406061
R29283 VGND.n3894 VGND.n3890 0.00406061
R29284 VGND.n7976 VGND.n7971 0.00406061
R29285 VGND.n1966 VGND.n1965 0.00406061
R29286 VGND.n7725 VGND.n7718 0.00406061
R29287 VGND.n7517 VGND.n7511 0.00406061
R29288 VGND.n8151 VGND.n8150 0.00406061
R29289 VGND.n580 VGND.n573 0.00406061
R29290 VGND.n1139 VGND.n1002 0.00406061
R29291 VGND.n1320 VGND.n1143 0.00406061
R29292 VGND.n1200 VGND.n1199 0.00406061
R29293 VGND.n990 VGND.n899 0.00406061
R29294 VGND.n7498 VGND.n7451 0.00406061
R29295 VGND.n799 VGND.n798 0.00406061
R29296 VGND.n7329 VGND.n820 0.00406061
R29297 VGND.n7325 VGND.n843 0.00406061
R29298 VGND.n6928 VGND.n6924 0.00406061
R29299 VGND.n6958 VGND.n6957 0.00406061
R29300 VGND.n6210 VGND.n6209 0.00406061
R29301 VGND.n6790 VGND.n1598 0.00406061
R29302 VGND.n6784 VGND.n6781 0.00406061
R29303 VGND.n6462 VGND.n6461 0.00406061
R29304 VGND.n5833 VGND.n5823 0.00406061
R29305 VGND.n2629 VGND.n2165 0.00406061
R29306 VGND.n6504 VGND.n6496 0.00406061
R29307 VGND.n5461 VGND.n5193 0.00406061
R29308 VGND.n5749 VGND.n5745 0.00406061
R29309 VGND.n9096 VGND.n9095 0.00406061
R29310 VGND.n5612 VGND.n5491 0.00406061
R29311 VGND.n2516 VGND.n2330 0.00406061
R29312 VGND.n9221 VGND.n9220 0.00406061
R29313 VGND.n1788 VGND.n1779 0.00406061
R29314 VGND.n3344 VGND.n3335 0.00393497
R29315 VGND.n8822 VGND.n8813 0.00393497
R29316 VGND.n3892 VGND.n3891 0.00393497
R29317 VGND.n7726 VGND.n7717 0.00393497
R29318 VGND.n581 VGND.n572 0.00393497
R29319 VGND.n4229 VGND.n4055 0.00393497
R29320 VGND.n6524 VGND.n1658 0.00393497
R29321 VGND.n2631 VGND.n2630 0.00393497
R29322 VGND.n5834 VGND.n5822 0.00393497
R29323 VGND.n4367 VGND.n4366 0.00393497
R29324 VGND.n6505 VGND.n6495 0.00393497
R29325 VGND.n2887 VGND.n44 0.00393497
R29326 VGND.n3019 VGND.n3018 0.00393497
R29327 VGND.n3021 VGND.n3020 0.00393497
R29328 VGND.n3179 VGND.n3023 0.00393497
R29329 VGND.n3022 VGND.n265 0.00393497
R29330 VGND.n8445 VGND.n8438 0.00393497
R29331 VGND.n8436 VGND.n8435 0.00393497
R29332 VGND.n7974 VGND.n7973 0.00393497
R29333 VGND.n8321 VGND.n317 0.00393497
R29334 VGND.n1364 VGND.n1363 0.00393497
R29335 VGND.n6997 VGND.n6990 0.00393497
R29336 VGND.n1569 VGND.n1568 0.00393497
R29337 VGND.n5299 VGND.n5298 0.00393497
R29338 VGND.n5463 VGND.n5462 0.00393497
R29339 VGND.n9094 VGND.n9093 0.00393497
R29340 VGND.n5191 VGND.n5190 0.00393497
R29341 VGND.n7972 VGND.n318 0.00393497
R29342 VGND.n6989 VGND.n6988 0.00393497
R29343 VGND.n7253 VGND.n7252 0.00393497
R29344 VGND.n4183 VGND.n1322 0.00393497
R29345 VGND.n4490 VGND.n4182 0.00393497
R29346 VGND.n2517 VGND.n46 0.00393497
R29347 VGND.n5613 VGND.n5490 0.00393497
R29348 VGND.n460 VGND.n459 0.00393497
R29349 VGND.n8112 VGND.n8111 0.00393497
R29350 VGND.n200 VGND.n199 0.00393497
R29351 VGND.n201 VGND.n72 0.00393497
R29352 VGND.n9068 VGND.n9067 0.00393497
R29353 VGND.n6735 VGND.n1614 0.00393497
R29354 VGND.n6762 VGND.n6761 0.00393497
R29355 VGND.n3583 VGND.n3582 0.00393497
R29356 VGND.n3729 VGND.n3728 0.00393497
R29357 VGND.n3768 VGND.n2039 0.00393497
R29358 VGND.n1875 VGND.n1874 0.00393497
R29359 VGND.n7518 VGND.n7507 0.00393497
R29360 VGND.n4763 VGND.n4752 0.00393497
R29361 VGND.n4706 VGND.n4705 0.00393497
R29362 VGND.n6011 VGND.n6010 0.00393497
R29363 VGND.n6006 VGND.n6005 0.00393497
R29364 VGND.n3537 VGND.n3536 0.00393497
R29365 VGND.n6009 VGND.n6008 0.00393497
R29366 VGND.n4800 VGND.n4798 0.00360244
R29367 VGND.n4130 VGND.n4128 0.00360244
R29368 VGND.n2079 VGND.n2077 0.00360244
R29369 VGND.n3699 VGND.n3698 0.00360244
R29370 VGND.n3811 VGND.n3809 0.00360244
R29371 VGND.n1917 VGND.n1915 0.00360244
R29372 VGND.n7528 VGND.n7527 0.00360244
R29373 VGND.n7490 VGND.n7488 0.00360244
R29374 VGND.n6152 VGND.n6150 0.00360244
R29375 VGND.n1746 VGND.n1745 0.00360244
R29376 VGND.n1832 VGND.n1830 0.00360244
R29377 VGND.n3516 VGND.n3514 0.00360244
R29378 VGND.n6494 VGND.n6493 0.00358437
R29379 VGND.n5297 VGND.n5296 0.00358437
R29380 VGND.n6764 VGND.n6763 0.00358437
R29381 VGND.n6092 VGND.n6091 0.00358437
R29382 VGND.n6159 VGND.n6115 0.0033671
R29383 VGND.n6268 VGND.n6267 0.0033671
R29384 VGND.n826 VGND.n825 0.0032017
R29385 VGND.n6476 VGND.n1659 0.0032017
R29386 VGND.n4364 VGND.n1659 0.0032017
R29387 VGND.n827 VGND.n826 0.0032017
R29388 VGND.n996 VGND.n995 0.0032017
R29389 VGND.n6955 VGND.n1542 0.0032017
R29390 VGND.n5296 VGND.n1542 0.0032017
R29391 VGND.n995 VGND.n994 0.0032017
R29392 VGND.n7276 VGND.n7275 0.0032017
R29393 VGND.n7277 VGND.n7276 0.0032017
R29394 VGND.n7503 VGND.n7502 0.0032017
R29395 VGND.n7504 VGND.n7503 0.0032017
R29396 VGND.n5822 VGND 0.00314375
R29397 VGND.n5190 VGND 0.00314375
R29398 VGND.n5490 VGND 0.00314375
R29399 VGND.n6005 VGND 0.00314375
R29400 VGND.n4802 VGND 0.00310417
R29401 VGND VGND.n5014 0.00310417
R29402 VGND VGND.n2895 0.00310417
R29403 VGND.n7816 VGND.n7815 0.00310417
R29404 VGND.n7981 VGND 0.00310417
R29405 VGND.n7690 VGND.n7688 0.00310417
R29406 VGND VGND.n8201 0.00310417
R29407 VGND.n7320 VGND.n7316 0.00310417
R29408 VGND.n6632 VGND.n1636 0.00310417
R29409 VGND.n5629 VGND 0.00310417
R29410 VGND.n2163 VGND.n2162 0.0028004
R29411 VGND.n7715 VGND.n582 0.0028004
R29412 VGND.n7728 VGND.n7727 0.0028004
R29413 VGND.n8811 VGND.n135 0.0028004
R29414 VGND.n8824 VGND.n8823 0.0028004
R29415 VGND.n3346 VGND.n3345 0.0028004
R29416 VGND.n5002 VGND.n5001 0.0028004
R29417 VGND.n4363 VGND.n4231 0.0028004
R29418 VGND.n2370 VGND.n43 0.0028004
R29419 VGND.n5790 VGND.n5789 0.0028004
R29420 VGND.n2537 VGND.n2536 0.0028004
R29421 VGND.n5620 VGND.n5619 0.0028004
R29422 VGND.n4489 VGND.n4209 0.0028004
R29423 VGND.n8096 VGND.n476 0.0028004
R29424 VGND.n8711 VGND.n203 0.0028004
R29425 VGND.n9065 VGND.n9050 0.0028004
R29426 VGND.n9087 VGND.n47 0.0028004
R29427 VGND.n8211 VGND.n8210 0.0028004
R29428 VGND.n3540 VGND.n2092 0.0028004
R29429 VGND.n3621 VGND.n3611 0.0028004
R29430 VGND.n3767 VGND.n3757 0.0028004
R29431 VGND.n2030 VGND.n2003 0.0028004
R29432 VGND.n7519 VGND.n748 0.0028004
R29433 VGND.n4824 VGND.n4823 0.0028004
R29434 VGND.n4750 VGND.n4143 0.0028004
R29435 VGND.n6089 VGND.n1697 0.0028004
R29436 VGND.n3535 VGND.n3534 0.0028004
R29437 VGND.n5853 VGND.n5852 0.0028004
R29438 VGND.n1752 VGND.n1750 0.00251462
R29439 VGND.n4822 VGND.n4821 0.00251462
R29440 VGND.n4142 VGND.n4141 0.00251462
R29441 VGND.n4488 VGND.n4487 0.00251462
R29442 VGND.n4584 VGND.n4582 0.00251462
R29443 VGND.n4362 VGND.n4361 0.00251462
R29444 VGND.n2091 VGND.n2090 0.00251462
R29445 VGND.n3241 VGND.n3239 0.00251462
R29446 VGND.n3620 VGND.n3619 0.00251462
R29447 VGND.n9011 VGND.n57 0.00251462
R29448 VGND.n3766 VGND.n3765 0.00251462
R29449 VGND.n8714 VGND.n8712 0.00251462
R29450 VGND.n2002 VGND.n2001 0.00251462
R29451 VGND.n7911 VGND.n461 0.00251462
R29452 VGND.n7522 VGND.n7520 0.00251462
R29453 VGND.n8214 VGND.n8212 0.00251462
R29454 VGND.n8319 VGND.n8318 0.00251462
R29455 VGND.n571 VGND.n570 0.00251462
R29456 VGND.n8794 VGND.n8793 0.00251462
R29457 VGND.n134 VGND.n133 0.00251462
R29458 VGND.n3334 VGND.n3333 0.00251462
R29459 VGND.n7698 VGND.n7697 0.00251462
R29460 VGND.n5004 VGND.n5003 0.00251462
R29461 VGND.n412 VGND.n411 0.00251462
R29462 VGND.n1458 VGND.n1457 0.00251462
R29463 VGND.n8095 VGND.n8094 0.00251462
R29464 VGND.n8710 VGND.n8709 0.00251462
R29465 VGND.n9049 VGND.n9048 0.00251462
R29466 VGND.n2762 VGND.n2761 0.00251462
R29467 VGND.n5344 VGND.n1613 0.00251462
R29468 VGND.n2630 VGND.n2163 0.00246749
R29469 VGND.n4367 VGND.n4363 0.00246749
R29470 VGND.n6523 VGND.n6505 0.00246749
R29471 VGND.n5853 VGND.n5834 0.00246749
R29472 VGND.n582 VGND.n581 0.00246749
R29473 VGND.n7727 VGND.n7726 0.00246749
R29474 VGND.n3892 VGND.n135 0.00246749
R29475 VGND.n8823 VGND.n8822 0.00246749
R29476 VGND.n3345 VGND.n3344 0.00246749
R29477 VGND.n5002 VGND.n4055 0.00246749
R29478 VGND.n6524 VGND.n6523 0.00246749
R29479 VGND.n9094 VGND.n43 0.00246749
R29480 VGND.n8320 VGND.n318 0.00246749
R29481 VGND.n6988 VGND.n1378 0.00246749
R29482 VGND.n5790 VGND.n5191 0.00246749
R29483 VGND.n5462 VGND.n5192 0.00246749
R29484 VGND.n3018 VGND.n2744 0.00246749
R29485 VGND.n3180 VGND.n3179 0.00246749
R29486 VGND.n8446 VGND.n8445 0.00246749
R29487 VGND.n7974 VGND.n279 0.00246749
R29488 VGND.n8435 VGND.n279 0.00246749
R29489 VGND.n8446 VGND.n265 0.00246749
R29490 VGND.n3180 VGND.n3021 0.00246749
R29491 VGND.n2887 VGND.n2744 0.00246749
R29492 VGND.n8321 VGND.n8320 0.00246749
R29493 VGND.n6998 VGND.n6997 0.00246749
R29494 VGND.n6998 VGND.n1364 0.00246749
R29495 VGND.n5299 VGND.n5192 0.00246749
R29496 VGND.n1568 VGND.n1378 0.00246749
R29497 VGND.n2537 VGND.n2517 0.00246749
R29498 VGND.n9068 VGND.n47 0.00246749
R29499 VGND.n9050 VGND.n72 0.00246749
R29500 VGND.n8711 VGND.n200 0.00246749
R29501 VGND.n8111 VGND.n8096 0.00246749
R29502 VGND.n8211 VGND.n460 0.00246749
R29503 VGND.n6761 VGND.n6736 0.00246749
R29504 VGND.n6736 VGND.n6735 0.00246749
R29505 VGND.n5619 VGND.n5613 0.00246749
R29506 VGND.n4490 VGND.n4489 0.00246749
R29507 VGND.n7227 VGND.n1322 0.00246749
R29508 VGND.n7252 VGND.n7227 0.00246749
R29509 VGND.n3536 VGND.n3535 0.00246749
R29510 VGND.n6008 VGND.n6007 0.00246749
R29511 VGND.n3582 VGND.n2092 0.00246749
R29512 VGND.n3728 VGND.n3621 0.00246749
R29513 VGND.n3768 VGND.n3767 0.00246749
R29514 VGND.n2003 VGND.n1875 0.00246749
R29515 VGND.n7519 VGND.n7518 0.00246749
R29516 VGND.n4823 VGND.n4763 0.00246749
R29517 VGND.n4706 VGND.n4143 0.00246749
R29518 VGND.n6011 VGND.n1697 0.00246749
R29519 VGND.n6007 VGND.n6006 0.00246749
R29520 VGND.n4377 VGND.n4376 0.00228056
R29521 VGND.n8786 VGND.n8785 0.00228056
R29522 VGND.n6457 VGND.n6456 0.00228056
R29523 VGND.n2624 VGND.n2623 0.00228056
R29524 VGND.n5012 VGND.n5011 0.00228056
R29525 VGND.n3328 VGND.n3327 0.00228056
R29526 VGND.n8911 VGND.n82 0.00228056
R29527 VGND.n5817 VGND.n5816 0.00228056
R29528 VGND.n1785 VGND.n1782 0.00218919
R29529 VGND.n1794 VGND.n1793 0.00218919
R29530 VGND.n5977 VGND.n5976 0.00218919
R29531 VGND.n5985 VGND.n5984 0.00218919
R29532 VGND.n1854 VGND.n1849 0.00218919
R29533 VGND.n1754 VGND.n1753 0.00218919
R29534 VGND.n1702 VGND.n1701 0.00218919
R29535 VGND.n6076 VGND.n6075 0.00218919
R29536 VGND.n6081 VGND.n6080 0.00218919
R29537 VGND.n6014 VGND.n1775 0.00218919
R29538 VGND.n6531 VGND.n6530 0.00218919
R29539 VGND.n1355 VGND.n1354 0.00218919
R29540 VGND.n7095 VGND.n1357 0.00218919
R29541 VGND.n4819 VGND.n4816 0.00218919
R29542 VGND.n4805 VGND.n4804 0.00218919
R29543 VGND.n4826 VGND.n4825 0.00218919
R29544 VGND.n4831 VGND.n4830 0.00218919
R29545 VGND.n4761 VGND.n4760 0.00218919
R29546 VGND.n4067 VGND.n4066 0.00218919
R29547 VGND.n4139 VGND.n4136 0.00218919
R29548 VGND.n4156 VGND.n4155 0.00218919
R29549 VGND.n4737 VGND.n4736 0.00218919
R29550 VGND.n4742 VGND.n4741 0.00218919
R29551 VGND.n4709 VGND.n4699 0.00218919
R29552 VGND.n1385 VGND.n1384 0.00218919
R29553 VGND.n1388 VGND.n1387 0.00218919
R29554 VGND.n4327 VGND.n4326 0.00218919
R29555 VGND.n2881 VGND.n2880 0.00218919
R29556 VGND.n3004 VGND.n2883 0.00218919
R29557 VGND.n2088 VGND.n2085 0.00218919
R29558 VGND.n3454 VGND.n3453 0.00218919
R29559 VGND.n3542 VGND.n3541 0.00218919
R29560 VGND.n3547 VGND.n3546 0.00218919
R29561 VGND.n3580 VGND.n2100 0.00218919
R29562 VGND.n2137 VGND.n2136 0.00218919
R29563 VGND.n3134 VGND.n3133 0.00218919
R29564 VGND.n3159 VGND.n3136 0.00218919
R29565 VGND.n3617 VGND.n3614 0.00218919
R29566 VGND.n3589 VGND.n3588 0.00218919
R29567 VGND.n3598 VGND.n3597 0.00218919
R29568 VGND.n3603 VGND.n3602 0.00218919
R29569 VGND.n3726 VGND.n3629 0.00218919
R29570 VGND.n113 VGND.n112 0.00218919
R29571 VGND.n259 VGND.n258 0.00218919
R29572 VGND.n262 VGND.n261 0.00218919
R29573 VGND.n3763 VGND.n3760 0.00218919
R29574 VGND.n3735 VGND.n3734 0.00218919
R29575 VGND.n3744 VGND.n3743 0.00218919
R29576 VGND.n3749 VGND.n3748 0.00218919
R29577 VGND.n3771 VGND.n1869 0.00218919
R29578 VGND.n144 VGND.n143 0.00218919
R29579 VGND.n296 VGND.n295 0.00218919
R29580 VGND.n299 VGND.n298 0.00218919
R29581 VGND.n1999 VGND.n1996 0.00218919
R29582 VGND.n2008 VGND.n2007 0.00218919
R29583 VGND.n2017 VGND.n2016 0.00218919
R29584 VGND.n2022 VGND.n2021 0.00218919
R29585 VGND.n1967 VGND.n1961 0.00218919
R29586 VGND.n551 VGND.n550 0.00218919
R29587 VGND.n7524 VGND.n7523 0.00218919
R29588 VGND.n726 VGND.n725 0.00218919
R29589 VGND.n735 VGND.n734 0.00218919
R29590 VGND.n740 VGND.n739 0.00218919
R29591 VGND.n7516 VGND.n7515 0.00218919
R29592 VGND.n414 VGND.n413 0.00218919
R29593 VGND.n428 VGND.n416 0.00218919
R29594 VGND.n591 VGND.n590 0.00218919
R29595 VGND.n1165 VGND.n1164 0.00218919
R29596 VGND.n1182 VGND.n1167 0.00218919
R29597 VGND.n7497 VGND.n7495 0.00218919
R29598 VGND.n783 VGND.n782 0.00218919
R29599 VGND.n755 VGND.n754 0.00218919
R29600 VGND.n762 VGND.n761 0.00218919
R29601 VGND.n800 VGND.n796 0.00218919
R29602 VGND.n849 VGND.n848 0.00218919
R29603 VGND.n1575 VGND.n1574 0.00218919
R29604 VGND.n1578 VGND.n1577 0.00218919
R29605 VGND.n6158 VGND.n6157 0.00218919
R29606 VGND.n6105 VGND.n6104 0.00218919
R29607 VGND.n6173 VGND.n6172 0.00218919
R29608 VGND.n6191 VGND.n6190 0.00218919
R29609 VGND.n6211 VGND.n1694 0.00218919
R29610 VGND.n1682 VGND.n1681 0.00218919
R29611 VGND.n2156 VGND.n2155 0.00218919
R29612 VGND.n5301 VGND.n5300 0.00218919
R29613 VGND.n5304 VGND.n5303 0.00218919
R29614 VGND.n5742 VGND.n5741 0.00218919
R29615 VGND.n5467 VGND.n5466 0.00218919
R29616 VGND.n2359 VGND.n2358 0.00218919
R29617 VGND.n2378 VGND.n2361 0.00218919
R29618 VGND.n3478 VGND.n3477 0.00218919
R29619 VGND.n3483 VGND.n3482 0.00218919
R29620 VGND.n9229 VGND.n9228 0.00218919
R29621 VGND.n9226 VGND.n9217 0.00218919
R29622 VGND.n9208 VGND.n9207 0.00218919
R29623 VGND.n5118 VGND.n5117 0.00218919
R29624 VGND.n5855 VGND.n5854 0.00218193
R29625 VGND.n2237 VGND.n2235 0.00218193
R29626 VGND.n6522 VGND.n6521 0.00218193
R29627 VGND.n5792 VGND.n5791 0.00218193
R29628 VGND.n2396 VGND.n2394 0.00218193
R29629 VGND.n8413 VGND.n8412 0.00218193
R29630 VGND.n8448 VGND.n8447 0.00218193
R29631 VGND.n3182 VGND.n3181 0.00218193
R29632 VGND.n2975 VGND.n2974 0.00218193
R29633 VGND.n7000 VGND.n6999 0.00218193
R29634 VGND.n5220 VGND.n5219 0.00218193
R29635 VGND.n5618 VGND.n5617 0.00218193
R29636 VGND.n2540 VGND.n2538 0.00218193
R29637 VGND.n7226 VGND.n7225 0.00218193
R29638 VGND.n3468 VGND.n3467 0.00218193
R29639 VGND.n1853 VGND.n1789 0.00218193
R29640 VGND.n6207 VGND.n1696 0.00185526
R29641 VGND.n4810 VGND.n4808 0.00180208
R29642 VGND.n4848 VGND.n4847 0.00180208
R29643 VGND.n4977 VGND.n4976 0.00180208
R29644 VGND.n7102 VGND.n7099 0.00180208
R29645 VGND.n7097 VGND.n7096 0.00180208
R29646 VGND.n4153 VGND.n4152 0.00180208
R29647 VGND.n4729 VGND.n4727 0.00180208
R29648 VGND.n4329 VGND.n4328 0.00180208
R29649 VGND.n4576 VGND.n4572 0.00180208
R29650 VGND.n4570 VGND.n4569 0.00180208
R29651 VGND.n3459 VGND.n3458 0.00180208
R29652 VGND.n3563 VGND.n3562 0.00180208
R29653 VGND.n3363 VGND.n3362 0.00180208
R29654 VGND VGND.n3230 0.00180208
R29655 VGND.n3009 VGND.n3008 0.00180208
R29656 VGND.n3006 VGND.n3005 0.00180208
R29657 VGND.n3709 VGND.n3708 0.00180208
R29658 VGND.n3716 VGND.n3715 0.00180208
R29659 VGND.n8841 VGND.n8840 0.00180208
R29660 VGND.n3165 VGND.n3163 0.00180208
R29661 VGND.n3161 VGND.n3160 0.00180208
R29662 VGND.n3819 VGND.n3818 0.00180208
R29663 VGND.n3827 VGND.n3826 0.00180208
R29664 VGND.n3900 VGND.n3899 0.00180208
R29665 VGND.n8657 VGND 0.00180208
R29666 VGND.n8564 VGND.n8562 0.00180208
R29667 VGND.n8560 VGND.n8559 0.00180208
R29668 VGND.n1990 VGND.n1988 0.00180208
R29669 VGND.n1982 VGND.n1981 0.00180208
R29670 VGND.n7746 VGND.n7745 0.00180208
R29671 VGND.n7983 VGND.n7982 0.00180208
R29672 VGND.n7980 VGND.n7979 0.00180208
R29673 VGND.n7538 VGND.n7537 0.00180208
R29674 VGND.n7548 VGND.n7547 0.00180208
R29675 VGND.n7614 VGND.n7613 0.00180208
R29676 VGND.n8134 VGND 0.00180208
R29677 VGND.n435 VGND.n432 0.00180208
R29678 VGND.n430 VGND.n429 0.00180208
R29679 VGND.n779 VGND.n778 0.00180208
R29680 VGND.n7442 VGND.n7440 0.00180208
R29681 VGND.n871 VGND.n870 0.00180208
R29682 VGND.n1188 VGND.n1186 0.00180208
R29683 VGND.n1184 VGND.n1183 0.00180208
R29684 VGND.n6111 VGND.n6110 0.00180208
R29685 VGND.n6178 VGND.n6177 0.00180208
R29686 VGND.n1684 VGND.n1683 0.00180208
R29687 VGND.n6941 VGND.n6940 0.00180208
R29688 VGND.n6944 VGND.n6943 0.00180208
R29689 VGND.n1762 VGND.n1761 0.00180208
R29690 VGND.n6068 VGND.n6066 0.00180208
R29691 VGND.n6555 VGND.n6554 0.00180208
R29692 VGND.n5307 VGND.n5196 0.00180208
R29693 VGND.n5310 VGND.n5309 0.00180208
R29694 VGND.n1841 VGND.n1840 0.00180208
R29695 VGND.n5997 VGND.n5995 0.00180208
R29696 VGND.n5874 VGND.n5873 0.00180208
R29697 VGND.n5762 VGND.n5761 0.00180208
R29698 VGND.n5765 VGND.n5764 0.00180208
R29699 VGND.n3525 VGND.n3524 0.00180208
R29700 VGND.n4 VGND.n0 0.00180208
R29701 VGND.n2262 VGND.n2261 0.00180208
R29702 VGND.n2384 VGND.n2382 0.00180208
R29703 VGND.n2380 VGND.n2379 0.00180208
R29704 VGND.n6955 VGND.n6954 0.0014919
R29705 VGND.n6207 VGND.n6195 0.0014919
R29706 VGND.n6492 VGND.n6476 0.00144128
R29707 VGND.n7327 VGND.n842 0.00142658
R29708 VGND.n7298 VGND.n895 0.00142658
R29709 VGND.n7291 VGND.n7272 0.00142658
R29710 VGND.n7500 VGND.n7450 0.00142658
R29711 VGND.n6787 VGND.n1612 0.00140106
R29712 VGND.n6787 VGND.n6780 0.00140106
R29713 VGND.n828 VGND.n827 0.00107355
R29714 VGND.n997 VGND.n996 0.00107355
R29715 VGND.n7278 VGND.n7277 0.00107355
R29716 VGND.n7502 VGND.n7501 0.00107355
R29717 VGND.n825 VGND.n824 0.00107344
R29718 VGND.n824 VGND.n823 0.00107344
R29719 VGND.n994 VGND.n993 0.00107344
R29720 VGND.n993 VGND.n992 0.00107344
R29721 VGND.n7274 VGND.n7273 0.00107344
R29722 VGND.n7275 VGND.n7274 0.00107344
R29723 VGND.n7505 VGND.n7504 0.00107344
R29724 VGND.n7506 VGND.n7505 0.00107344
R29725 VGND.n7327 VGND.n828 0.00107332
R29726 VGND.n7298 VGND.n997 0.00107332
R29727 VGND.n7291 VGND.n7278 0.00107332
R29728 VGND.n7501 VGND.n7500 0.00107332
R29729 trimb[4].n9 trimb[4].n8 349.738
R29730 trimb[4].n11 trimb[4].n10 292.5
R29731 trimb[4].n11 trimb[4].n4 292.5
R29732 trimb[4].n13 trimb[4].n3 193.387
R29733 trimb[4].n7 trimb[4].n5 151.127
R29734 trimb[4].n7 trimb[4].n6 107.763
R29735 trimb[4].n5 trimb[4].t5 40.0005
R29736 trimb[4].n5 trimb[4].t6 40.0005
R29737 trimb[4].n6 trimb[4].t7 40.0005
R29738 trimb[4].n6 trimb[4].t4 40.0005
R29739 trimb[4].n8 trimb[4].t0 27.5805
R29740 trimb[4].n8 trimb[4].t1 27.5805
R29741 trimb[4].n12 trimb[4].t2 23.6405
R29742 trimb[4].n3 trimb[4].t3 23.1644
R29743 trimb[4].n10 trimb[4].n9 14.7697
R29744 trimb[4].n4 trimb[4].n2 11.243
R29745 trimb[4] trimb[4].n7 10.4115
R29746 trimb[4].n13 trimb[4].n1 9.3005
R29747 trimb[4].n14 trimb[4].n13 9.3005
R29748 trimb[4].n13 trimb[4].n12 9.3005
R29749 trimb[4].n14 trimb[4].n0 9.04377
R29750 trimb[4].n1 trimb[4].n0 9.01973
R29751 trimb[4].n11 trimb[4].n3 4.23401
R29752 trimb[4].n15 trimb[4].n2 4.13041
R29753 trimb[4].n12 trimb[4].n11 3.9405
R29754 trimb[4].n13 trimb[4].n2 3.09077
R29755 trimb[4] trimb[4].n16 2.48707
R29756 trimb[4].n16 trimb[4].n15 2.24426
R29757 trimb[4].n9 trimb[4].n4 1.96973
R29758 trimb[4].n10 trimb[4] 0.246654
R29759 trimb[4].n15 trimb[4].n1 0.03175
R29760 trimb[4].n16 trimb[4].n0 0.0141816
R29761 trimb[4].n15 trimb[4].n14 0.0101154
R29762 clknet_2_1__leaf_clk.n35 clknet_2_1__leaf_clk.t33 294.557
R29763 clknet_2_1__leaf_clk.n51 clknet_2_1__leaf_clk.t39 294.557
R29764 clknet_2_1__leaf_clk.n37 clknet_2_1__leaf_clk.t45 294.557
R29765 clknet_2_1__leaf_clk.n39 clknet_2_1__leaf_clk.t54 294.557
R29766 clknet_2_1__leaf_clk.n41 clknet_2_1__leaf_clk.t56 294.557
R29767 clknet_2_1__leaf_clk.n33 clknet_2_1__leaf_clk.t49 294.557
R29768 clknet_2_1__leaf_clk.n27 clknet_2_1__leaf_clk.t36 294.557
R29769 clknet_2_1__leaf_clk.n30 clknet_2_1__leaf_clk.t43 294.557
R29770 clknet_2_1__leaf_clk.n43 clknet_2_1__leaf_clk.t42 292.704
R29771 clknet_2_1__leaf_clk.n45 clknet_2_1__leaf_clk.t47 292.704
R29772 clknet_2_1__leaf_clk.n17 clknet_2_1__leaf_clk.t52 292.704
R29773 clknet_2_1__leaf_clk.n15 clknet_2_1__leaf_clk.t34 292.704
R29774 clknet_2_1__leaf_clk.n21 clknet_2_1__leaf_clk.t40 292.704
R29775 clknet_2_1__leaf_clk.n43 clknet_2_1__leaf_clk.t48 211.56
R29776 clknet_2_1__leaf_clk.n45 clknet_2_1__leaf_clk.t51 211.56
R29777 clknet_2_1__leaf_clk.n17 clknet_2_1__leaf_clk.t35 211.56
R29778 clknet_2_1__leaf_clk.n15 clknet_2_1__leaf_clk.t44 211.56
R29779 clknet_2_1__leaf_clk.n21 clknet_2_1__leaf_clk.t46 211.56
R29780 clknet_2_1__leaf_clk.n35 clknet_2_1__leaf_clk.t41 211.01
R29781 clknet_2_1__leaf_clk.n51 clknet_2_1__leaf_clk.t50 211.01
R29782 clknet_2_1__leaf_clk.n37 clknet_2_1__leaf_clk.t55 211.01
R29783 clknet_2_1__leaf_clk.n39 clknet_2_1__leaf_clk.t37 211.01
R29784 clknet_2_1__leaf_clk.n41 clknet_2_1__leaf_clk.t38 211.01
R29785 clknet_2_1__leaf_clk.n33 clknet_2_1__leaf_clk.t57 211.01
R29786 clknet_2_1__leaf_clk.n27 clknet_2_1__leaf_clk.t53 211.01
R29787 clknet_2_1__leaf_clk.n30 clknet_2_1__leaf_clk.t32 211.01
R29788 clknet_2_1__leaf_clk.n67 clknet_2_1__leaf_clk.n65 187.052
R29789 clknet_2_1__leaf_clk.n3 clknet_2_1__leaf_clk.n1 156.138
R29790 clknet_2_1__leaf_clk.n67 clknet_2_1__leaf_clk.n66 155.052
R29791 clknet_2_1__leaf_clk.n69 clknet_2_1__leaf_clk.n68 155.052
R29792 clknet_2_1__leaf_clk.n71 clknet_2_1__leaf_clk.n70 155.052
R29793 clknet_2_1__leaf_clk.n73 clknet_2_1__leaf_clk.n72 155.052
R29794 clknet_2_1__leaf_clk.n75 clknet_2_1__leaf_clk.n74 155.052
R29795 clknet_2_1__leaf_clk.n77 clknet_2_1__leaf_clk.n76 155.052
R29796 clknet_2_1__leaf_clk clknet_2_1__leaf_clk.n64 151.438
R29797 clknet_2_1__leaf_clk.n3 clknet_2_1__leaf_clk.n2 110.963
R29798 clknet_2_1__leaf_clk.n5 clknet_2_1__leaf_clk.n4 110.963
R29799 clknet_2_1__leaf_clk.n9 clknet_2_1__leaf_clk.n8 110.963
R29800 clknet_2_1__leaf_clk.n11 clknet_2_1__leaf_clk.n10 110.963
R29801 clknet_2_1__leaf_clk.n7 clknet_2_1__leaf_clk.n6 109.956
R29802 clknet_2_1__leaf_clk.n63 clknet_2_1__leaf_clk.n62 107.712
R29803 clknet_2_1__leaf_clk clknet_2_1__leaf_clk.n35 80.2062
R29804 clknet_2_1__leaf_clk clknet_2_1__leaf_clk.n51 80.2062
R29805 clknet_2_1__leaf_clk clknet_2_1__leaf_clk.n37 80.2062
R29806 clknet_2_1__leaf_clk clknet_2_1__leaf_clk.n39 80.2062
R29807 clknet_2_1__leaf_clk clknet_2_1__leaf_clk.n27 80.2062
R29808 clknet_2_1__leaf_clk clknet_2_1__leaf_clk.n30 80.2062
R29809 clknet_2_1__leaf_clk.n42 clknet_2_1__leaf_clk.n41 76.0005
R29810 clknet_2_1__leaf_clk.n34 clknet_2_1__leaf_clk.n33 76.0005
R29811 clknet_2_1__leaf_clk.n5 clknet_2_1__leaf_clk.n3 45.177
R29812 clknet_2_1__leaf_clk.n11 clknet_2_1__leaf_clk.n9 45.177
R29813 clknet_2_1__leaf_clk.n61 clknet_2_1__leaf_clk.n11 45.177
R29814 clknet_2_1__leaf_clk.n7 clknet_2_1__leaf_clk.n5 44.0476
R29815 clknet_2_1__leaf_clk.n9 clknet_2_1__leaf_clk.n7 44.0476
R29816 clknet_2_1__leaf_clk.n12 clknet_2_1__leaf_clk.t26 40.2593
R29817 clknet_2_1__leaf_clk.n1 clknet_2_1__leaf_clk.t30 40.0005
R29818 clknet_2_1__leaf_clk.n1 clknet_2_1__leaf_clk.t27 40.0005
R29819 clknet_2_1__leaf_clk.n2 clknet_2_1__leaf_clk.t16 40.0005
R29820 clknet_2_1__leaf_clk.n2 clknet_2_1__leaf_clk.t18 40.0005
R29821 clknet_2_1__leaf_clk.n4 clknet_2_1__leaf_clk.t20 40.0005
R29822 clknet_2_1__leaf_clk.n4 clknet_2_1__leaf_clk.t21 40.0005
R29823 clknet_2_1__leaf_clk.n6 clknet_2_1__leaf_clk.t17 40.0005
R29824 clknet_2_1__leaf_clk.n6 clknet_2_1__leaf_clk.t19 40.0005
R29825 clknet_2_1__leaf_clk.n8 clknet_2_1__leaf_clk.t25 40.0005
R29826 clknet_2_1__leaf_clk.n8 clknet_2_1__leaf_clk.t22 40.0005
R29827 clknet_2_1__leaf_clk.n10 clknet_2_1__leaf_clk.t23 40.0005
R29828 clknet_2_1__leaf_clk.n10 clknet_2_1__leaf_clk.t24 40.0005
R29829 clknet_2_1__leaf_clk.n62 clknet_2_1__leaf_clk.t29 40.0005
R29830 clknet_2_1__leaf_clk.n62 clknet_2_1__leaf_clk.t31 40.0005
R29831 clknet_2_1__leaf_clk.n12 clknet_2_1__leaf_clk.t28 36.9737
R29832 clknet_2_1__leaf_clk.n69 clknet_2_1__leaf_clk.n67 32.0005
R29833 clknet_2_1__leaf_clk.n71 clknet_2_1__leaf_clk.n69 32.0005
R29834 clknet_2_1__leaf_clk.n75 clknet_2_1__leaf_clk.n73 32.0005
R29835 clknet_2_1__leaf_clk.n77 clknet_2_1__leaf_clk.n75 32.0005
R29836 clknet_2_1__leaf_clk.n73 clknet_2_1__leaf_clk.n71 31.2005
R29837 clknet_2_1__leaf_clk.n64 clknet_2_1__leaf_clk.t0 27.5805
R29838 clknet_2_1__leaf_clk.n64 clknet_2_1__leaf_clk.t2 27.5805
R29839 clknet_2_1__leaf_clk.n65 clknet_2_1__leaf_clk.t1 27.5805
R29840 clknet_2_1__leaf_clk.n65 clknet_2_1__leaf_clk.t14 27.5805
R29841 clknet_2_1__leaf_clk.n66 clknet_2_1__leaf_clk.t3 27.5805
R29842 clknet_2_1__leaf_clk.n66 clknet_2_1__leaf_clk.t5 27.5805
R29843 clknet_2_1__leaf_clk.n68 clknet_2_1__leaf_clk.t7 27.5805
R29844 clknet_2_1__leaf_clk.n68 clknet_2_1__leaf_clk.t8 27.5805
R29845 clknet_2_1__leaf_clk.n70 clknet_2_1__leaf_clk.t4 27.5805
R29846 clknet_2_1__leaf_clk.n70 clknet_2_1__leaf_clk.t6 27.5805
R29847 clknet_2_1__leaf_clk.n72 clknet_2_1__leaf_clk.t12 27.5805
R29848 clknet_2_1__leaf_clk.n72 clknet_2_1__leaf_clk.t9 27.5805
R29849 clknet_2_1__leaf_clk.n74 clknet_2_1__leaf_clk.t10 27.5805
R29850 clknet_2_1__leaf_clk.n74 clknet_2_1__leaf_clk.t11 27.5805
R29851 clknet_2_1__leaf_clk.n76 clknet_2_1__leaf_clk.t13 27.5805
R29852 clknet_2_1__leaf_clk.n76 clknet_2_1__leaf_clk.t15 27.5805
R29853 clknet_2_1__leaf_clk.n48 clknet_2_1__leaf_clk 19.1246
R29854 clknet_2_1__leaf_clk.n47 clknet_2_1__leaf_clk.n46 17.7668
R29855 clknet_2_1__leaf_clk.n53 clknet_2_1__leaf_clk.n50 14.1755
R29856 clknet_2_1__leaf_clk.n61 clknet_2_1__leaf_clk.n60 13.7535
R29857 clknet_2_1__leaf_clk.n63 clknet_2_1__leaf_clk.n61 13.177
R29858 clknet_2_1__leaf_clk.n19 clknet_2_1__leaf_clk.n16 11.993
R29859 clknet_2_1__leaf_clk.n55 clknet_2_1__leaf_clk.n54 11.353
R29860 clknet_2_1__leaf_clk.n49 clknet_2_1__leaf_clk.n40 10.6768
R29861 clknet_2_1__leaf_clk clknet_2_1__leaf_clk.n42 10.4234
R29862 clknet_2_1__leaf_clk clknet_2_1__leaf_clk.n34 10.4234
R29863 clknet_2_1__leaf_clk.n78 clknet_2_1__leaf_clk.n77 10.2022
R29864 clknet_2_1__leaf_clk.n36 clknet_2_1__leaf_clk 9.32621
R29865 clknet_2_1__leaf_clk.n52 clknet_2_1__leaf_clk 9.32621
R29866 clknet_2_1__leaf_clk.n38 clknet_2_1__leaf_clk 9.32621
R29867 clknet_2_1__leaf_clk.n40 clknet_2_1__leaf_clk 9.32621
R29868 clknet_2_1__leaf_clk.n28 clknet_2_1__leaf_clk 9.32621
R29869 clknet_2_1__leaf_clk.n31 clknet_2_1__leaf_clk 9.32621
R29870 clknet_2_1__leaf_clk.n32 clknet_2_1__leaf_clk.n29 9.28724
R29871 clknet_2_1__leaf_clk.n18 clknet_2_1__leaf_clk.n17 7.84669
R29872 clknet_2_1__leaf_clk.n16 clknet_2_1__leaf_clk.n15 7.84669
R29873 clknet_2_1__leaf_clk.n44 clknet_2_1__leaf_clk.n43 7.84584
R29874 clknet_2_1__leaf_clk.n46 clknet_2_1__leaf_clk.n45 7.84584
R29875 clknet_2_1__leaf_clk.n56 clknet_2_1__leaf_clk.n32 7.60918
R29876 clknet_2_1__leaf_clk.n19 clknet_2_1__leaf_clk.n18 7.26768
R29877 clknet_2_1__leaf_clk.n22 clknet_2_1__leaf_clk.n21 7.10009
R29878 clknet_2_1__leaf_clk.n13 clknet_2_1__leaf_clk.n12 6.93977
R29879 clknet_2_1__leaf_clk.n29 clknet_2_1__leaf_clk.n28 6.71896
R29880 clknet_2_1__leaf_clk.n47 clknet_2_1__leaf_clk.n44 6.60337
R29881 clknet_2_1__leaf_clk.n58 clknet_2_1__leaf_clk.n56 6.53553
R29882 clknet_2_1__leaf_clk.n54 clknet_2_1__leaf_clk.n53 6.20946
R29883 clknet_2_1__leaf_clk.n50 clknet_2_1__leaf_clk.n49 6.20769
R29884 clknet_2_1__leaf_clk.n54 clknet_2_1__leaf_clk.n36 6.06336
R29885 clknet_2_1__leaf_clk.n56 clknet_2_1__leaf_clk.n55 6.01149
R29886 clknet_2_1__leaf_clk.n26 clknet_2_1__leaf_clk.n19 5.94006
R29887 clknet_2_1__leaf_clk.n32 clknet_2_1__leaf_clk.n31 4.6505
R29888 clknet_2_1__leaf_clk.n53 clknet_2_1__leaf_clk.n52 4.58353
R29889 clknet_2_1__leaf_clk.n50 clknet_2_1__leaf_clk.n38 4.58312
R29890 clknet_2_1__leaf_clk.n29 clknet_2_1__leaf_clk.n26 4.5005
R29891 clknet_2_1__leaf_clk.n0 clknet_2_1__leaf_clk.n23 4.01346
R29892 clknet_2_1__leaf_clk.n60 clknet_2_1__leaf_clk.n14 3.98526
R29893 clknet_2_1__leaf_clk.n26 clknet_2_1__leaf_clk.n25 3.79018
R29894 clknet_2_1__leaf_clk clknet_2_1__leaf_clk.n78 3.68119
R29895 clknet_2_1__leaf_clk.n36 clknet_2_1__leaf_clk 3.10907
R29896 clknet_2_1__leaf_clk.n52 clknet_2_1__leaf_clk 3.10907
R29897 clknet_2_1__leaf_clk.n38 clknet_2_1__leaf_clk 3.10907
R29898 clknet_2_1__leaf_clk.n40 clknet_2_1__leaf_clk 3.10907
R29899 clknet_2_1__leaf_clk.n28 clknet_2_1__leaf_clk 3.10907
R29900 clknet_2_1__leaf_clk.n31 clknet_2_1__leaf_clk 3.10907
R29901 clknet_2_1__leaf_clk.n24 clknet_2_1__leaf_clk.n0 3.0059
R29902 clknet_2_1__leaf_clk.n60 clknet_2_1__leaf_clk.n13 2.63794
R29903 clknet_2_1__leaf_clk.n18 clknet_2_1__leaf_clk 2.3354
R29904 clknet_2_1__leaf_clk.n16 clknet_2_1__leaf_clk 2.3354
R29905 clknet_2_1__leaf_clk.n44 clknet_2_1__leaf_clk 2.3353
R29906 clknet_2_1__leaf_clk.n46 clknet_2_1__leaf_clk 2.3353
R29907 clknet_2_1__leaf_clk.n48 clknet_2_1__leaf_clk.n47 2.2972
R29908 clknet_2_1__leaf_clk.n14 clknet_2_1__leaf_clk.n58 2.24505
R29909 clknet_2_1__leaf_clk.n42 clknet_2_1__leaf_clk 2.01193
R29910 clknet_2_1__leaf_clk.n34 clknet_2_1__leaf_clk 2.01193
R29911 clknet_2_1__leaf_clk.n49 clknet_2_1__leaf_clk.n48 1.99363
R29912 clknet_2_1__leaf_clk.n23 clknet_2_1__leaf_clk 1.69089
R29913 clknet_2_1__leaf_clk.n23 clknet_2_1__leaf_clk.n22 1.65408
R29914 clknet_2_1__leaf_clk.n55 clknet_2_1__leaf_clk 1.37207
R29915 clknet_2_1__leaf_clk clknet_2_1__leaf_clk.n63 1.26402
R29916 clknet_2_1__leaf_clk.n78 clknet_2_1__leaf_clk 0.0554356
R29917 clknet_2_1__leaf_clk.n0 clknet_2_1__leaf_clk.n20 0.0405928
R29918 clknet_2_1__leaf_clk.n14 clknet_2_1__leaf_clk.n59 0.0365577
R29919 clknet_2_1__leaf_clk.n25 clknet_2_1__leaf_clk.n24 0.0262437
R29920 clknet_2_1__leaf_clk.n58 clknet_2_1__leaf_clk.n57 0.01396
R29921 _063_.n10 _063_.t19 260.394
R29922 _063_.n8 _063_.t15 239.651
R29923 _063_.n3 _063_.t11 228.304
R29924 _063_.n4 _063_.t10 212.081
R29925 _063_.n5 _063_.t14 212.081
R29926 _063_.n18 _063_.n16 201.645
R29927 _063_.n8 _063_.t18 169.826
R29928 _063_.n3 _063_.t16 157.667
R29929 _063_.n10 _063_.t13 156.441
R29930 _063_.n4 _063_.t12 139.78
R29931 _063_.n5 _063_.t17 139.78
R29932 _063_.n18 _063_.n17 108.608
R29933 _063_.n19 _063_.n15 108.606
R29934 _063_ _063_.n21 106.278
R29935 _063_.n7 _063_.n6 100.96
R29936 _063_.n19 _063_.n18 57.0187
R29937 _063_.n6 _063_.n4 30.6732
R29938 _063_.n6 _063_.n5 30.6732
R29939 _063_.n20 _063_.n19 29.6732
R29940 _063_.n16 _063_.t6 26.5955
R29941 _063_.n16 _063_.t7 26.5955
R29942 _063_.n21 _063_.t2 26.5955
R29943 _063_.n21 _063_.t3 26.5955
R29944 _063_.n15 _063_.t9 26.5955
R29945 _063_.n15 _063_.t8 26.5955
R29946 _063_.n17 _063_.t1 26.5955
R29947 _063_.n17 _063_.t0 26.5955
R29948 _063_.n2 _063_.t4 24.7093
R29949 _063_.n2 _063_.t5 23.9668
R29950 _063_.n13 _063_ 16.8563
R29951 _063_.n9 _063_.n7 14.5761
R29952 _063_.n20 _063_ 13.5267
R29953 _063_.n0 _063_ 1.84272
R29954 _063_.n12 _063_.n11 9.20785
R29955 _063_.n14 _063_.n2 8.78218
R29956 _063_.n11 _063_.n10 8.16569
R29957 _063_.n14 _063_.n13 7.64136
R29958 _063_.n0 _063_.n3 8.53199
R29959 _063_.n1 _063_.n8 9.57193
R29960 _063_.n7 _063_ 5.1205
R29961 _063_ _063_.n14 4.94071
R29962 _063_.n12 _063_.n9 4.52385
R29963 _063_.n13 _063_.n12 3.20792
R29964 _063_.n11 _063_ 2.60881
R29965 _063_ _063_.n20 2.32777
R29966 _063_.n1 _063_ 5.3328
R29967 _063_.n0 _063_ 3.0365
R29968 _063_.n9 _063_.n1 3.52964
R29969 _048_.n5 _048_.t14 471.289
R29970 _048_.n32 _048_.t13 405.416
R29971 _048_.n26 _048_.t35 241.536
R29972 _048_.n30 _048_.t19 239.986
R29973 _048_.n10 _048_.t37 239.986
R29974 _048_.n15 _048_.t18 229.036
R29975 _048_.n12 _048_.t23 221.72
R29976 _048_.n13 _048_.t32 221.72
R29977 _048_.n18 _048_.t34 212.081
R29978 _048_.n17 _048_.t27 212.081
R29979 _048_.n7 _048_.t21 212.081
R29980 _048_.n8 _048_.t29 212.081
R29981 _048_.n23 _048_.t24 206.751
R29982 _048_.n2 _048_.n0 197.595
R29983 _048_.n26 _048_.t25 169.237
R29984 _048_.n30 _048_.t17 167.685
R29985 _048_.n10 _048_.t33 167.685
R29986 _048_.n41 _048_.n3 165.219
R29987 _048_.n39 _048_.n38 165.218
R29988 _048_.n15 _048_.t22 158.464
R29989 _048_.n19 _048_ 153.024
R29990 _048_.n12 _048_.t30 149.421
R29991 _048_.n13 _048_.t20 149.421
R29992 _048_.n5 _048_.t12 148.35
R29993 _048_.n23 _048_.t26 146.494
R29994 _048_.n18 _048_.t16 139.78
R29995 _048_.n17 _048_.t31 139.78
R29996 _048_.n7 _048_.t28 139.78
R29997 _048_.n8 _048_.t36 139.78
R29998 _048_.n2 _048_.n1 138.054
R29999 _048_.n32 _048_.t15 135.496
R30000 _048_.n39 _048_.n37 105.677
R30001 _048_.n41 _048_.n4 105.677
R30002 _048_.n11 _048_.n10 88.244
R30003 _048_.n6 _048_.n5 85.775
R30004 _048_ _048_.n30 83.5135
R30005 _048_ _048_.n26 82.6735
R30006 _048_ _048_.n9 81.791
R30007 _048_ _048_.n14 76.9605
R30008 _048_.n33 _048_.n32 76.0005
R30009 _048_.n18 _048_.n17 61.346
R30010 _048_.n27 _048_ 60.3156
R30011 _048_.n9 _048_.n7 40.1672
R30012 _048_.n14 _048_.n12 37.4894
R30013 _048_.n14 _048_.n13 37.4894
R30014 _048_.n22 _048_ 32.3436
R30015 _048_.n29 _048_ 28.4511
R30016 _048_.n0 _048_.t1 26.5955
R30017 _048_.n0 _048_.t4 26.5955
R30018 _048_.n3 _048_.t3 26.5955
R30019 _048_.n3 _048_.t0 26.5955
R30020 _048_.n38 _048_.t2 26.5955
R30021 _048_.n38 _048_.t5 26.5955
R30022 _048_.n37 _048_.t11 24.9236
R30023 _048_.n37 _048_.t8 24.9236
R30024 _048_.n1 _048_.t10 24.9236
R30025 _048_.n1 _048_.t7 24.9236
R30026 _048_.n4 _048_.t6 24.9236
R30027 _048_.n4 _048_.t9 24.9236
R30028 _048_.n19 _048_.n18 21.1793
R30029 _048_.n9 _048_.n8 21.1793
R30030 _048_.n20 _048_.n19 19.9024
R30031 _048_.n31 _048_ 16.6802
R30032 _048_.n29 _048_.n28 14.9255
R30033 _048_.n25 _048_.n24 13.7051
R30034 _048_.n34 _048_ 12.3175
R30035 _048_.n41 _048_.n40 12.0732
R30036 _048_.n16 _048_.n15 8.71725
R30037 _048_ _048_.n33 8.45333
R30038 _048_.n28 _048_.n27 8.37682
R30039 _048_.n27 _048_.n25 8.1449
R30040 _048_.n24 _048_.n23 8.04894
R30041 _048_.n33 _048_ 7.97031
R30042 _048_.n36 _048_.n35 7.82565
R30043 _048_.n40 _048_ 7.36386
R30044 _048_.n22 _048_.n21 6.84518
R30045 _048_.n35 _048_.n31 6.45533
R30046 _048_.n36 _048_.n6 6.06336
R30047 _048_.n21 _048_.n16 5.63748
R30048 _048_.n11 _048_ 4.73093
R30049 _048_.n35 _048_.n34 4.6505
R30050 _048_.n28 _048_.n11 4.58368
R30051 _048_.n34 _048_ 4.10616
R30052 _048_.n6 _048_ 3.95686
R30053 _048_ _048_.n41 3.49141
R30054 _048_.n20 _048_ 3.17702
R30055 _048_.n21 _048_.n20 3.13776
R30056 _048_.n24 _048_ 2.94112
R30057 _048_.n31 _048_.n29 2.9222
R30058 _048_.n16 _048_ 2.90557
R30059 _048_.n25 _048_.n22 2.59528
R30060 _048_ _048_.n2 2.47323
R30061 _048_ _048_.n36 1.30284
R30062 _048_.n40 _048_.n39 0.145955
R30063 net34.n8 net34.t0 440.25
R30064 net34.n0 net34.t4 238.59
R30065 net34.n3 net34.t2 212.081
R30066 net34.n2 net34.t3 212.081
R30067 net34.n0 net34.t7 203.244
R30068 net34.n3 net34.t5 139.78
R30069 net34.n2 net34.t6 139.78
R30070 net34.t0 net34.n6 133.933
R30071 net34.n7 net34.t1 123.654
R30072 net34 net34.n7 78.8791
R30073 net34.n1 net34.n0 76.0005
R30074 net34.n3 net34.n2 61.346
R30075 net34.n5 net34.n4 57.9773
R30076 net34.n4 net34.n3 39.6822
R30077 net34 net34.n8 10.9042
R30078 net34.n5 net34 9.17193
R30079 net34 net34.n1 8.22907
R30080 net34.n8 net34 5.21532
R30081 net34.n7 net34 5.16973
R30082 net34.n1 net34 4.20621
R30083 net34.n10 net34.n9 4.14532
R30084 net34.n9 net34 3.00754
R30085 net34.n9 net34.n6 2.97937
R30086 net34.n4 net34 2.44789
R30087 net34.n11 net34.n10 2.24505
R30088 net34 net34.n5 0.999271
R30089 net34 net34.n11 0.985393
R30090 sample.n15 sample.n14 585
R30091 sample.n11 sample.n10 349.738
R30092 sample.n13 sample.n12 292.5
R30093 sample.n13 sample.n6 292.5
R30094 sample.n9 sample.n7 151.127
R30095 sample.n9 sample.n8 107.763
R30096 sample.n7 sample.t6 40.0005
R30097 sample.n7 sample.t7 40.0005
R30098 sample.n8 sample.t4 40.0005
R30099 sample.n8 sample.t5 40.0005
R30100 sample.n10 sample.t0 27.5805
R30101 sample.n10 sample.t1 27.5805
R30102 sample.n4 sample.t3 23.7598
R30103 sample.n14 sample.t2 14.7755
R30104 sample.n12 sample.n11 14.7697
R30105 sample.n14 sample.n13 12.8055
R30106 sample.n6 sample.n3 11.243
R30107 sample sample.n9 10.4115
R30108 sample.n15 sample.n5 9.3005
R30109 sample.n16 sample.n15 9.3005
R30110 sample.n5 sample.n0 9.0697
R30111 sample.n17 sample.n16 9.02214
R30112 sample.n15 sample.n4 8.9018
R30113 sample.n3 sample.n2 4.13041
R30114 sample.n13 sample.n4 3.77188
R30115 sample.n18 sample.n17 3.41895
R30116 sample.n15 sample.n3 3.09077
R30117 sample.n11 sample.n6 1.96973
R30118 sample.n2 sample.n1 1.35818
R30119 sample.n18 sample.n0 0.868169
R30120 sample.n12 sample 0.246654
R30121 sample sample.n18 0.129323
R30122 sample.n17 sample.n1 0.0376622
R30123 sample.n16 sample.n2 0.03175
R30124 sample.n1 sample.n0 0.0103621
R30125 sample.n5 sample.n2 0.0101154
R30126 ctlp[4].n4 ctlp[4].n1 292.5
R30127 ctlp[4].n3 ctlp[4].n2 92.5005
R30128 ctlp[4] ctlp[4].n3 81.3181
R30129 ctlp[4].n1 ctlp[4].t0 26.5955
R30130 ctlp[4].n0 ctlp[4].t1 25.8903
R30131 ctlp[4].n2 ctlp[4].t2 24.9236
R30132 ctlp[4].n2 ctlp[4].t3 24.9236
R30133 ctlp[4] ctlp[4].n4 15.5613
R30134 ctlp[4].n6 ctlp[4] 10.132
R30135 ctlp[4].n5 ctlp[4].n0 9.48617
R30136 ctlp[4].n3 ctlp[4] 5.27109
R30137 ctlp[4].n5 ctlp[4] 2.60833
R30138 ctlp[4] ctlp[4].n5 1.85252
R30139 ctlp[4].n4 ctlp[4] 1.50638
R30140 ctlp[4].n1 ctlp[4].n0 0.248635
R30141 ctlp[4].n6 ctlp[4] 0.0844286
R30142 ctlp[4] ctlp[4].n6 0.012146
R30143 net30.n12 net30.n0 328.209
R30144 net30.n5 net30.t4 256.887
R30145 net30.n8 net30.t10 238.59
R30146 net30.n1 net30.t8 212.081
R30147 net30.n2 net30.t5 212.081
R30148 net30.n8 net30.t6 203.244
R30149 net30.n5 net30.t9 178.756
R30150 net30.n1 net30.t11 139.78
R30151 net30.n2 net30.t7 139.78
R30152 net30 net30.n13 123.963
R30153 net30.n9 net30.n8 76.0005
R30154 net30.n4 net30.n3 76.0005
R30155 net30.n11 net30 66.4415
R30156 net30.n13 net30.t3 38.5719
R30157 net30.n13 net30.t2 38.5719
R30158 net30.n3 net30.n1 30.6732
R30159 net30.n3 net30.n2 30.6732
R30160 net30.n0 net30.t1 26.5955
R30161 net30.n0 net30.t0 26.5955
R30162 net30.n7 net30.n4 25.4856
R30163 net30.n7 net30.n6 24.9815
R30164 net30.n9 net30 8.22907
R30165 net30.n6 net30.n5 7.99568
R30166 net30.n11 net30.n7 7.00204
R30167 net30 net30.n10 4.74918
R30168 net30.n12 net30.n11 4.6505
R30169 net30 net30.n12 3.2005
R30170 net30.n10 net30 3.10907
R30171 net30.n6 net30 1.94261
R30172 net30.n10 net30.n9 1.09764
R30173 net30.n4 net30 0.5125
R30174 trim[1].n11 trim[1].n10 585
R30175 trim[1].n9 trim[1].n7 291.764
R30176 trim[1].n4 trim[1].n2 151.127
R30177 trim[1].n4 trim[1].n3 107.763
R30178 trim[1].n6 trim[1].n5 96.9298
R30179 trim[1].n7 trim[1].n6 60.6531
R30180 trim[1].n2 trim[1].t6 40.0005
R30181 trim[1].n2 trim[1].t7 40.0005
R30182 trim[1].n3 trim[1].t4 40.0005
R30183 trim[1].n3 trim[1].t5 40.0005
R30184 trim[1].n5 trim[1].t0 27.5805
R30185 trim[1].n5 trim[1].t1 27.5805
R30186 trim[1].n8 trim[1].t2 25.6105
R30187 trim[1].n10 trim[1].n9 14.7755
R30188 trim[1].n10 trim[1].t3 12.8055
R30189 trim[1] trim[1].n4 10.4115
R30190 trim[1].n6 trim[1] 9.6475
R30191 trim[1].n11 trim[1].n1 9.3005
R30192 trim[1].n11 trim[1].n8 9.3005
R30193 trim[1].n12 trim[1].n0 9.05196
R30194 trim[1].n1 trim[1].n0 9.01492
R30195 trim[1].n12 trim[1].n11 3.72602
R30196 trim[1].n11 trim[1].n7 2.70497
R30197 trim[1] trim[1].n14 2.52311
R30198 trim[1].n14 trim[1].n13 2.24426
R30199 trim[1].n9 trim[1].n8 1.9705
R30200 trim[1].n13 trim[1].n1 0.0365577
R30201 trim[1].n14 trim[1].n0 0.0141816
R30202 trim[1].n13 trim[1].n12 0.00292567
R30203 ctlp[6].n2 ctlp[6].n0 151.127
R30204 ctlp[6].n2 ctlp[6].n1 107.763
R30205 ctlp[6].n11 ctlp[6].n10 96.9298
R30206 ctlp[6].n11 ctlp[6].n9 60.5294
R30207 ctlp[6].n0 ctlp[6].t4 40.0005
R30208 ctlp[6].n0 ctlp[6].t6 40.0005
R30209 ctlp[6].n1 ctlp[6].t5 40.0005
R30210 ctlp[6].n1 ctlp[6].t7 40.0005
R30211 ctlp[6].n10 ctlp[6].t3 27.5805
R30212 ctlp[6].n10 ctlp[6].t1 27.5805
R30213 ctlp[6].n7 ctlp[6].t0 25.6105
R30214 ctlp[6].n12 ctlp[6] 19.2609
R30215 ctlp[6].n12 ctlp[6].n11 15.309
R30216 ctlp[6].n6 ctlp[6].n5 14.7755
R30217 ctlp[6].n5 ctlp[6].t2 12.8055
R30218 ctlp[6].n8 ctlp[6] 10.9647
R30219 ctlp[6].n8 ctlp[6].n7 9.3005
R30220 ctlp[6] ctlp[6].n3 9.00791
R30221 ctlp[6].n3 ctlp[6].n2 6.77697
R30222 ctlp[6] ctlp[6].n4 3.62598
R30223 ctlp[6] ctlp[6].n12 2.70819
R30224 ctlp[6].n9 ctlp[6].n8 2.58125
R30225 ctlp[6].n7 ctlp[6].n6 1.9705
R30226 ctlp[6].n3 ctlp[6] 1.73877
R30227 ctlp[6].n4 ctlp[6] 0.154033
R30228 ctlp[6].n4 ctlp[6] 0.00363333
R30229 result[3].n10 result[3].n7 185
R30230 result[3].n4 result[3].n3 143.643
R30231 result[3].n5 result[3] 81.5159
R30232 result[3].n3 result[3].t1 26.5955
R30233 result[3].n3 result[3].t0 26.5955
R30234 result[3].n6 result[3].t3 24.9236
R30235 result[3].n7 result[3].n6 15.6928
R30236 result[3].n10 result[3].n9 9.3005
R30237 result[3].n11 result[3].n10 9.3005
R30238 result[3].n7 result[3].t2 9.23127
R30239 result[3].n12 result[3].n11 9.05098
R30240 result[3].n9 result[3].n0 9.04085
R30241 result[3] result[3].n4 9.02598
R30242 result[3].n6 result[3].n5 8.25053
R30243 result[3].n4 result[3] 7.64268
R30244 result[3].n8 result[3].n2 3.79439
R30245 result[3].n13 result[3].n12 3.41895
R30246 result[3].n8 result[3] 2.08974
R30247 result[3].n10 result[3].n8 2.03855
R30248 result[3].n2 result[3].n1 1.35818
R30249 result[3].n13 result[3].n0 0.868169
R30250 result[3].n10 result[3].n5 0.214619
R30251 result[3] result[3].n13 0.129323
R30252 result[3].n9 result[3].n2 0.0389615
R30253 result[3].n12 result[3].n1 0.0376622
R30254 result[3].n1 result[3].n0 0.0103621
R30255 result[3].n11 result[3].n2 0.00290385
R30256 net43.n120 net43.t11 413.315
R30257 net43.n134 net43.t40 413.315
R30258 net43.n103 net43.t26 413.313
R30259 net43.n68 net43.t37 413.313
R30260 net43.n92 net43.t21 413.313
R30261 net43.n82 net43.t31 413.313
R30262 net43.n72 net43.t46 413.313
R30263 net43.n56 net43.t19 413.313
R30264 net43.n45 net43.t34 413.313
R30265 net43.n129 net43.t38 413.313
R30266 net43.n148 net43.n147 354.634
R30267 net43.n117 net43.t42 344.005
R30268 net43.n138 net43.t10 344.005
R30269 net43.n107 net43.t14 343.113
R30270 net43.n65 net43.t24 343.113
R30271 net43.n98 net43.t35 343.113
R30272 net43.n86 net43.t30 343.113
R30273 net43.n76 net43.t45 343.113
R30274 net43.n53 net43.t47 343.113
R30275 net43.n42 net43.t17 343.113
R30276 net43.n126 net43.t39 343.113
R30277 net43.n105 net43.t25 187.798
R30278 net43.n63 net43.t23 187.798
R30279 net43.n95 net43.t13 187.798
R30280 net43.n84 net43.t20 187.798
R30281 net43.n74 net43.t33 187.798
R30282 net43.n51 net43.t36 187.798
R30283 net43.n40 net43.t8 187.798
R30284 net43.n124 net43.t9 187.798
R30285 net43.n116 net43.t22 187.321
R30286 net43.n133 net43.t32 187.321
R30287 net43.n107 net43.n106 152
R30288 net43.n65 net43.n64 152
R30289 net43.n98 net43.n97 152
R30290 net43.n86 net43.n85 152
R30291 net43.n76 net43.n75 152
R30292 net43.n53 net43.n52 152
R30293 net43.n42 net43.n41 152
R30294 net43.n117 net43.n115 152
R30295 net43.n139 net43.n138 152
R30296 net43.n126 net43.n125 152
R30297 net43.n37 net43.n35 151.127
R30298 net43.n120 net43.t18 126.127
R30299 net43.n134 net43.t44 126.127
R30300 net43.n103 net43.t16 126.127
R30301 net43.n68 net43.t15 126.127
R30302 net43.n92 net43.t27 126.127
R30303 net43.n82 net43.t43 126.127
R30304 net43.n72 net43.t12 126.127
R30305 net43.n56 net43.t28 126.127
R30306 net43.n45 net43.t41 126.127
R30307 net43.n129 net43.t29 126.127
R30308 net43.n37 net43.n36 107.763
R30309 net43.n148 net43.n146 96.9298
R30310 net43.n105 net43.n104 73.4143
R30311 net43.n63 net43.n62 73.4143
R30312 net43.n96 net43.n95 73.4143
R30313 net43.n84 net43.n83 73.4143
R30314 net43.n74 net43.n73 73.4143
R30315 net43.n51 net43.n50 73.4143
R30316 net43.n40 net43.n39 73.4143
R30317 net43.n124 net43.n123 73.4143
R30318 net43.n116 net43.n113 73.2067
R30319 net43.n133 net43.n132 73.2067
R30320 net43.n35 net43.t6 40.0005
R30321 net43.n35 net43.t7 40.0005
R30322 net43.n36 net43.t4 40.0005
R30323 net43.n36 net43.t5 40.0005
R30324 net43.n142 net43 28.6268
R30325 net43.n143 net43.n142 27.962
R30326 net43.n146 net43.t1 27.5805
R30327 net43.n146 net43.t2 27.5805
R30328 net43.n147 net43.t3 27.5805
R30329 net43.n147 net43.t0 27.5805
R30330 net43 net43.n114 14.0185
R30331 net43.n140 net43 14.0185
R30332 net43.n100 net43 10.8576
R30333 net43.n69 net43.n68 10.648
R30334 net43.n93 net43.n92 10.648
R30335 net43.n57 net43.n56 10.648
R30336 net43.n46 net43.n45 10.648
R30337 net43.n130 net43.n129 10.648
R30338 net43.n121 net43.n120 10.647
R30339 net43.n135 net43.n134 10.647
R30340 net43 net43.n37 10.4115
R30341 net43 net43.n148 9.6475
R30342 net43.n107 net43.n105 9.63724
R30343 net43.n65 net43.n63 9.63724
R30344 net43.n98 net43.n95 9.63724
R30345 net43.n86 net43.n84 9.63724
R30346 net43.n76 net43.n74 9.63724
R30347 net43.n53 net43.n51 9.63724
R30348 net43.n42 net43.n40 9.63724
R30349 net43.n126 net43.n124 9.63724
R30350 net43.n145 net43.n144 9.44462
R30351 net43.n23 net43.n22 1.8618
R30352 net43.n108 net43.n107 9.3005
R30353 net43.n111 net43.n110 9.3005
R30354 net43.n25 net43.n26 2.84046
R30355 net43.n31 net43.n9 2.82124
R30356 net43.n66 net43.n65 9.3005
R30357 net43 net43.n67 9.3005
R30358 net43.n21 net43.n20 1.8618
R30359 net43.n87 net43.n86 9.3005
R30360 net43.n90 net43.n89 9.3005
R30361 net43.n27 net43.n28 2.84046
R30362 net43.n19 net43.n18 1.8618
R30363 net43.n77 net43.n76 9.3005
R30364 net43.n80 net43.n79 9.3005
R30365 net43.n29 net43.n30 2.84046
R30366 net43.n99 net43.n34 0.569404
R30367 net43.n99 net43.n98 9.3005
R30368 net43.n24 net43 2.75366
R30369 net43 net43.n34 4.3668
R30370 net43.n17 net43.n16 1.8618
R30371 net43.n54 net43.n53 9.3005
R30372 net43.n15 net43.n14 1.8618
R30373 net43.n43 net43.n42 9.3005
R30374 net43 net43.n119 9.3005
R30375 net43.n32 net43.n10 2.82124
R30376 net43.n118 net43.n117 9.3005
R30377 net43.n13 net43.n12 1.8618
R30378 net43.n138 net43.n137 9.3005
R30379 net43.n33 net43.n11 2.82124
R30380 net43.n127 net43.n126 9.3005
R30381 net43 net43.n128 9.3005
R30382 net43.n117 net43.n116 9.15991
R30383 net43.n138 net43.n133 9.15991
R30384 net43.n5 net43.n81 9.0005
R30385 net43 net43.n3 6.79444
R30386 net43.n2 net43.n102 9.0005
R30387 net43.n145 net43 8.05976
R30388 net43.n111 net43.n103 7.02742
R30389 net43.n90 net43.n82 7.02742
R30390 net43.n80 net43.n72 7.02742
R30391 net43 net43.n49 6.86314
R30392 net43.n143 net43 5.84528
R30393 net43.n101 net43.n100 5.66671
R30394 net43.n102 net43.n101 4.97887
R30395 net43.n144 net43.n0 5.01211
R30396 net43.n114 net43 4.7293
R30397 net43.n141 net43.n140 4.6505
R30398 net43.n114 net43 4.53383
R30399 net43.n140 net43 4.53383
R30400 net43.n61 net43.n60 4.5005
R30401 net43.n4 net43.n71 4.48961
R30402 net43.n1 net43.n38 4.48961
R30403 net43.n8 net43.n7 0.0199018
R30404 net43.n5 net43.n3 2.98419
R30405 net43.n2 net43.n0 2.98419
R30406 net43.n101 net43.n61 4.4222
R30407 net43.n144 net43.n143 3.20792
R30408 net43.n106 net43 3.11401
R30409 net43.n64 net43 3.11401
R30410 net43.n97 net43 3.11401
R30411 net43.n85 net43 3.11401
R30412 net43.n75 net43 3.11401
R30413 net43.n52 net43 3.11401
R30414 net43.n41 net43 3.11401
R30415 net43.n115 net43 3.11401
R30416 net43 net43.n139 3.11401
R30417 net43.n125 net43 3.11401
R30418 net43.n26 net43.n111 3.46381
R30419 net43.n28 net43.n90 3.46381
R30420 net43.n30 net43.n80 3.46381
R30421 net43 net43.n145 2.68692
R30422 net43.n109 net43 2.36657
R30423 net43 net43.n70 2.36657
R30424 net43.n88 net43 2.36657
R30425 net43.n78 net43 2.36657
R30426 net43 net43.n94 2.36657
R30427 net43 net43.n122 2.36657
R30428 net43 net43.n136 2.36657
R30429 net43 net43.n131 2.36657
R30430 net43.n61 net43 2.36314
R30431 net43.n55 net43 1.83532
R30432 net43.n44 net43 1.83532
R30433 net43.n106 net43.n104 1.55726
R30434 net43.n64 net43.n62 1.55726
R30435 net43.n67 net43.n31 1.97739
R30436 net43.n97 net43.n96 1.55726
R30437 net43.n85 net43.n83 1.55726
R30438 net43.n75 net43.n73 1.55726
R30439 net43.n52 net43.n50 1.55726
R30440 net43.n41 net43.n39 1.55726
R30441 net43.n115 net43.n113 1.55726
R30442 net43.n119 net43.n32 1.97739
R30443 net43.n139 net43.n132 1.55726
R30444 net43.n125 net43.n123 1.55726
R30445 net43.n128 net43.n33 1.97739
R30446 net43.n108 net43.n104 1.38428
R30447 net43.n23 net43.n108 1.23632
R30448 net43.n23 net43 2.68891
R30449 net43.n66 net43.n62 1.38428
R30450 net43.n31 net43.n66 0.84027
R30451 net43.n67 net43 1.38428
R30452 net43.n24 net43.n99 1.96578
R30453 net43.n87 net43.n83 1.38428
R30454 net43.n21 net43.n87 1.23632
R30455 net43.n21 net43 2.68891
R30456 net43.n77 net43.n73 1.38428
R30457 net43.n19 net43.n77 1.23632
R30458 net43.n19 net43 2.68891
R30459 net43.n54 net43.n50 1.38428
R30460 net43.n17 net43.n54 1.23632
R30461 net43.n17 net43 2.68891
R30462 net43.n43 net43.n39 1.38428
R30463 net43.n15 net43.n43 1.23632
R30464 net43.n15 net43 2.68891
R30465 net43.n118 net43.n113 1.38428
R30466 net43.n32 net43.n118 0.84027
R30467 net43.n119 net43 1.38428
R30468 net43.n137 net43.n132 1.38428
R30469 net43.n137 net43.n13 1.23632
R30470 net43.n13 net43 2.68891
R30471 net43.n127 net43.n123 1.38428
R30472 net43.n33 net43.n127 0.84027
R30473 net43.n128 net43 1.38428
R30474 net43.n2 net43.n26 22.5084
R30475 net43.n5 net43.n28 22.5084
R30476 net43.n8 net43.n30 22.5084
R30477 net43.n24 net43 2.22988
R30478 net43.n55 net43 1.11211
R30479 net43.n44 net43 1.11211
R30480 net43.n109 net43 0.580857
R30481 net43.n70 net43 0.580857
R30482 net43.n88 net43 0.580857
R30483 net43.n78 net43 0.580857
R30484 net43.n94 net43 0.580857
R30485 net43.n58 net43 0.580857
R30486 net43.n47 net43 0.580857
R30487 net43.n122 net43 0.580857
R30488 net43.n136 net43 0.580857
R30489 net43.n131 net43 0.580857
R30490 net43.n59 net43 0.445212
R30491 net43.n48 net43 0.445212
R30492 net43.n142 net43.n141 0.383906
R30493 net43.n69 net43 0.272889
R30494 net43.n93 net43 0.272889
R30495 net43.n57 net43 0.272889
R30496 net43.n46 net43 0.272889
R30497 net43.n121 net43 0.272889
R30498 net43.n135 net43 0.272889
R30499 net43.n130 net43 0.272889
R30500 net43.n59 net43.n58 0.246036
R30501 net43.n48 net43.n47 0.246036
R30502 net43.n100 net43 0.179071
R30503 net43.n112 net43 0.17713
R30504 net43.n91 net43 0.17713
R30505 net43.n6 net43 0.17713
R30506 net43.n96 net43.n34 0.742377
R30507 net43.n112 net43.n25 0.0847391
R30508 net43.n91 net43.n27 0.0847391
R30509 net43.n6 net43.n29 0.0847391
R30510 net43.n70 net43.n69 0.0827155
R30511 net43.n94 net43.n93 0.0827155
R30512 net43.n58 net43.n57 0.0827155
R30513 net43.n47 net43.n46 0.0827155
R30514 net43.n122 net43.n121 0.0827155
R30515 net43.n136 net43.n135 0.0827155
R30516 net43.n131 net43.n130 0.0827155
R30517 net43.n141 net43 0.0793043
R30518 net43.n60 net43.n55 0.0774231
R30519 net43.n60 net43.n59 0.0774231
R30520 net43.n49 net43.n44 0.0774231
R30521 net43.n49 net43.n48 0.0774231
R30522 net43.n7 net43.n6 0.0935116
R30523 net43.n1 net43.n112 0.0550287
R30524 net43.n4 net43.n91 0.0550287
R30525 net43.n3 net43.n71 0.0185295
R30526 net43.n0 net43.n38 0.0185295
R30527 net43.n81 net43.n71 0.0509808
R30528 net43.n102 net43.n38 0.0509808
R30529 net43 net43.n22 0.04675
R30530 net43 net43.n20 0.04675
R30531 net43 net43.n18 0.04675
R30532 net43 net43.n16 0.04675
R30533 net43 net43.n14 0.04675
R30534 net43.n12 net43 0.04675
R30535 net43 net43.n11 0.04675
R30536 net43 net43.n10 0.04675
R30537 net43 net43.n9 0.04675
R30538 net43.n110 net43.n109 0.0466957
R30539 net43.n89 net43.n88 0.0466957
R30540 net43.n79 net43.n78 0.0466957
R30541 net43.n79 net43.n29 0.0466957
R30542 net43.n89 net43.n27 0.0466957
R30543 net43.n110 net43.n25 0.0466957
R30544 net43.n8 net43 0.0442052
R30545 net43.n5 net43 0.0442052
R30546 net43.n2 net43 0.0442052
R30547 net43 net43.n11 0.0335068
R30548 net43.n12 net43 0.0335068
R30549 net43 net43.n10 0.0335068
R30550 net43 net43.n14 0.0335068
R30551 net43 net43.n16 0.0335068
R30552 net43 net43.n18 0.0335068
R30553 net43 net43.n20 0.0335068
R30554 net43 net43.n9 0.0335068
R30555 net43 net43.n22 0.0335068
R30556 net43.n81 net43.n7 6.1473
R30557 net43.n5 net43.n4 0.0578686
R30558 net43.n2 net43.n1 0.0578686
R30559 result[6].n2 result[6].n1 354.634
R30560 result[6].n6 result[6].n4 151.127
R30561 result[6].n6 result[6].n5 107.763
R30562 result[6].n2 result[6].n0 96.9298
R30563 result[6].n4 result[6].t6 40.0005
R30564 result[6].n4 result[6].t4 40.0005
R30565 result[6].n5 result[6].t5 40.0005
R30566 result[6].n5 result[6].t7 40.0005
R30567 result[6].n0 result[6].t0 27.5805
R30568 result[6].n0 result[6].t2 27.5805
R30569 result[6].n1 result[6].t1 27.5805
R30570 result[6].n1 result[6].t3 27.5805
R30571 result[6] result[6].n3 19.2609
R30572 result[6].n3 result[6].n2 15.309
R30573 result[6] result[6].n8 10.0086
R30574 result[6].n8 result[6] 8.05976
R30575 result[6].n7 result[6].n6 6.77697
R30576 result[6].n3 result[6] 2.70819
R30577 result[6].n7 result[6] 1.73877
R30578 result[6].n8 result[6].n7 0.948648
R30579 ctln[6].n2 ctln[6].n0 354.634
R30580 ctln[6].n12 ctln[6].n4 107.763
R30581 ctln[6].n2 ctln[6].n1 96.9298
R30582 ctln[6].n12 ctln[6].n11 58.6278
R30583 ctln[6].n10 ctln[6].t6 40.3946
R30584 ctln[6].n4 ctln[6].t4 40.0005
R30585 ctln[6].n4 ctln[6].t5 40.0005
R30586 ctln[6].n10 ctln[6].t7 36.871
R30587 ctln[6].n1 ctln[6].t3 27.5805
R30588 ctln[6].n1 ctln[6].t0 27.5805
R30589 ctln[6].n0 ctln[6].t1 27.5805
R30590 ctln[6].n0 ctln[6].t2 27.5805
R30591 ctln[6] ctln[6].n3 19.2609
R30592 ctln[6].n3 ctln[6].n2 15.309
R30593 ctln[6].n13 ctln[6] 9.00791
R30594 ctln[6].n11 ctln[6].n10 7.36486
R30595 ctln[6].n13 ctln[6].n12 6.77697
R30596 ctln[6].n11 ctln[6].n9 4.57357
R30597 ctln[6].n6 ctln[6] 4.21294
R30598 ctln[6].n3 ctln[6] 2.70819
R30599 ctln[6].n8 ctln[6].n6 2.24426
R30600 ctln[6] ctln[6].n13 1.73877
R30601 ctln[6].n8 ctln[6].n7 0.0365577
R30602 ctln[6].n6 ctln[6].n5 0.0141816
R30603 ctln[6].n9 ctln[6].n8 0.00336382
R30604 trimb[0].n12 trimb[0].n5 585
R30605 trimb[0].n4 trimb[0].n3 349.738
R30606 trimb[0].n10 trimb[0].n9 292.5
R30607 trimb[0].n10 trimb[0].n4 152.91
R30608 trimb[0].n8 trimb[0].n6 151.127
R30609 trimb[0].n8 trimb[0].n7 107.763
R30610 trimb[0].n6 trimb[0].t6 40.0005
R30611 trimb[0].n6 trimb[0].t4 40.0005
R30612 trimb[0].n7 trimb[0].t7 40.0005
R30613 trimb[0].n7 trimb[0].t5 40.0005
R30614 trimb[0].n3 trimb[0].t3 27.5805
R30615 trimb[0].n3 trimb[0].t1 27.5805
R30616 trimb[0].n11 trimb[0].t0 23.6405
R30617 trimb[0].n5 trimb[0].t2 14.7755
R30618 trimb[0].n10 trimb[0].n5 12.8055
R30619 trimb[0].n9 trimb[0].n2 11.243
R30620 trimb[0] trimb[0].n8 10.4115
R30621 trimb[0].n12 trimb[0].n1 9.3005
R30622 trimb[0].n13 trimb[0].n12 9.3005
R30623 trimb[0].n12 trimb[0].n11 9.3005
R30624 trimb[0].n13 trimb[0].n0 9.04377
R30625 trimb[0].n1 trimb[0].n0 9.01973
R30626 trimb[0].n14 trimb[0].n2 4.13041
R30627 trimb[0].n11 trimb[0].n10 3.9405
R30628 trimb[0].n12 trimb[0].n2 3.09077
R30629 trimb[0] trimb[0].n15 2.29709
R30630 trimb[0].n15 trimb[0].n14 2.24426
R30631 trimb[0].n9 trimb[0] 0.246654
R30632 trimb[0].n12 trimb[0].n4 0.246654
R30633 trimb[0].n14 trimb[0].n1 0.03175
R30634 trimb[0].n15 trimb[0].n0 0.0141816
R30635 trimb[0].n14 trimb[0].n13 0.0101154
R30636 _065_.n12 _065_.t10 471.289
R30637 _065_ _065_.n1 303.024
R30638 _065_.n2 _065_.t9 238.59
R30639 _065_.n5 _065_.t18 229.233
R30640 _065_.n9 _065_.t6 229.001
R30641 _065_.n18 _065_.t17 212.081
R30642 _065_.n19 _065_.t7 212.081
R30643 _065_.n26 _065_.t16 206.19
R30644 _065_.n2 _065_.t13 203.244
R30645 _065_.n6 _065_.t8 192.639
R30646 _065_.n5 _065_.t5 158.671
R30647 _065_.n9 _065_.t12 156.702
R30648 _065_.n26 _065_.t11 148.35
R30649 _065_.n12 _065_.t19 148.35
R30650 _065_.n18 _065_.t4 139.78
R30651 _065_.n19 _065_.t14 139.78
R30652 _065_.n6 _065_.t15 134.799
R30653 _065_ _065_.n29 112.127
R30654 _065_.n10 _065_.n9 90.6968
R30655 _065_ _065_.n12 81.8187
R30656 _065_.n7 _065_.n6 80.2291
R30657 _065_ _065_.n26 78.6571
R30658 _065_.n3 _065_.n2 76.0005
R30659 _065_.n22 _065_.n18 35.7853
R30660 _065_.n16 _065_ 27.5205
R30661 _065_.n1 _065_.t0 26.5955
R30662 _065_.n1 _065_.t1 26.5955
R30663 _065_.n29 _065_.t3 24.9236
R30664 _065_.n29 _065_.t2 24.9236
R30665 _065_.n27 _065_ 22.9285
R30666 _065_.n27 _065_.n25 19.0554
R30667 _065_.n13 _065_.n11 18.5184
R30668 _065_.n11 _065_.n8 16.9816
R30669 _065_.n28 _065_ 14.5072
R30670 _065_.n20 _065_.n19 13.146
R30671 _065_.n14 _065_.n4 13.1049
R30672 _065_.n28 _065_.n27 11.596
R30673 _065_.n13 _065_ 9.78835
R30674 _065_.n21 _065_.n20 9.49444
R30675 _065_.n23 _065_.n22 9.3005
R30676 _065_.n3 _065_ 8.22907
R30677 _065_.n24 _065_.n23 7.99801
R30678 _065_.n14 _065_.n13 7.48814
R30679 _065_.n0 _065_.n5 8.69361
R30680 _065_.n11 _065_.n10 5.01055
R30681 _065_ _065_.n28 4.83606
R30682 _065_.n8 _065_.n7 4.58184
R30683 _065_.n15 _065_.n14 4.37172
R30684 _065_.n17 _065_.n16 4.1605
R30685 _065_.n10 _065_ 4.03013
R30686 _065_.n0 _065_ 3.17119
R30687 _065_.n4 _065_ 3.10907
R30688 _065_.n22 _065_.n21 2.92171
R30689 _065_.n7 _065_ 1.94336
R30690 _065_.n23 _065_.n17 1.2805
R30691 _065_.n4 _065_.n3 1.09764
R30692 _065_.n8 _065_ 0.0802539
R30693 _065_.n25 _065_.n24 0.0533846
R30694 _065_.n24 _065_.n15 0.0509808
R30695 _065_.n0 _065_ 13.6983
R30696 ctlp[7].n2 ctlp[7].n0 151.127
R30697 ctlp[7].n2 ctlp[7].n1 107.763
R30698 ctlp[7].n11 ctlp[7].n10 96.9298
R30699 ctlp[7].n11 ctlp[7].n9 60.5294
R30700 ctlp[7].n0 ctlp[7].t5 40.0005
R30701 ctlp[7].n0 ctlp[7].t6 40.0005
R30702 ctlp[7].n1 ctlp[7].t7 40.0005
R30703 ctlp[7].n1 ctlp[7].t4 40.0005
R30704 ctlp[7].n10 ctlp[7].t3 27.5805
R30705 ctlp[7].n10 ctlp[7].t0 27.5805
R30706 ctlp[7].n7 ctlp[7].t2 25.6105
R30707 ctlp[7].n12 ctlp[7] 19.2609
R30708 ctlp[7].n12 ctlp[7].n11 15.309
R30709 ctlp[7].n6 ctlp[7].n5 14.7755
R30710 ctlp[7].n8 ctlp[7] 13.7751
R30711 ctlp[7].n5 ctlp[7].t1 12.8055
R30712 ctlp[7].n8 ctlp[7].n7 9.3005
R30713 ctlp[7] ctlp[7].n3 9.00791
R30714 ctlp[7].n3 ctlp[7].n2 6.77697
R30715 ctlp[7] ctlp[7].n12 2.70819
R30716 ctlp[7].n9 ctlp[7].n8 2.58125
R30717 ctlp[7].n7 ctlp[7].n6 1.9705
R30718 ctlp[7].n3 ctlp[7] 1.73877
R30719 ctlp[7] ctlp[7].n4 0.106146
R30720 ctlp[7].n4 ctlp[7] 0.0739375
R30721 ctlp[7].n4 ctlp[7] 0.0138097
R30722 result[4].n8 result[4].n7 185
R30723 result[4].n4 result[4].n3 143.643
R30724 result[4].n5 result[4] 81.5159
R30725 result[4].n3 result[4].t1 26.5955
R30726 result[4].n3 result[4].t0 26.5955
R30727 result[4].n6 result[4].t3 24.9236
R30728 result[4].n7 result[4].n6 15.6928
R30729 result[4].n8 result[4].n1 9.3005
R30730 result[4].n9 result[4].n8 9.3005
R30731 result[4].n7 result[4].t2 9.23127
R30732 result[4].n9 result[4].n0 9.05098
R30733 result[4] result[4].n4 9.02598
R30734 result[4].n1 result[4].n0 9.01252
R30735 result[4].n6 result[4].n5 8.25053
R30736 result[4].n4 result[4] 7.64268
R30737 result[4].n10 result[4].n2 3.79439
R30738 result[4] result[4].n11 2.45104
R30739 result[4].n11 result[4].n10 2.24426
R30740 result[4].n2 result[4] 2.08974
R30741 result[4].n8 result[4].n2 2.03855
R30742 result[4].n8 result[4].n5 0.214619
R30743 result[4].n10 result[4].n1 0.0389615
R30744 result[4].n11 result[4].n0 0.0141816
R30745 result[4].n10 result[4].n9 0.00290385
R30746 _123_.n8 _123_.t5 337.832
R30747 _123_.n6 _123_.t6 241.536
R30748 _123_.n11 _123_.t4 241.536
R30749 _123_.n5 _123_.n3 192.752
R30750 _123_.n6 _123_.t8 169.237
R30751 _123_.n11 _123_.t7 169.237
R30752 _123_.n8 _123_.t3 153.666
R30753 _123_.n15 _123_.n2 143.026
R30754 _123_.n7 _123_.n6 87.2645
R30755 _123_.n12 _123_.n11 87.2645
R30756 _123_.n0 _123_.t1 85.775
R30757 _123_ _123_.n15 29.0496
R30758 _123_.n4 _123_.t2 25.6105
R30759 _123_.n3 _123_.t0 21.126
R30760 _123_.n14 _123_.n13 17.2044
R30761 _123_.n10 _123_.n9 16.3826
R30762 _123_.n15 _123_.n14 15.2685
R30763 _123_.n9 _123_ 15.0071
R30764 _123_.n5 _123_.n4 9.3005
R30765 _123_.n13 _123_.n12 7.75331
R30766 _123_.n10 _123_.n7 6.06336
R30767 _123_.n3 _123_.n2 5.19377
R30768 _123_.n1 _123_.n0 4.13971
R30769 _123_ _123_.n1 3.76521
R30770 _123_.n7 _123_ 3.0725
R30771 _123_.n12 _123_ 3.0725
R30772 _123_ _123_.n10 2.36534
R30773 _123_.n9 _123_.n8 1.88374
R30774 _123_.n0 _123_ 1.18808
R30775 _123_.n14 _123_.n5 1.12307
R30776 _123_.n4 _123_.n2 0.9855
R30777 _123_.n1 _123_ 0.921363
R30778 _123_.n13 _123_ 0.541709
R30779 _051_.n21 _051_.t21 334.188
R30780 _051_.n8 _051_.t12 327.507
R30781 _051_.n6 _051_.t20 293.969
R30782 _051_.n19 _051_.t15 233.989
R30783 _051_.n11 _051_.t14 204.656
R30784 _051_.n8 _051_.t16 201.119
R30785 _051_ _051_.n1 197.595
R30786 _051_.n5 _051_.n3 165.219
R30787 _051_.n27 _051_.n26 165.218
R30788 _051_.n18 _051_.t19 158.602
R30789 _051_.n6 _051_.t13 138.338
R30790 _051_ _051_.n0 138.054
R30791 _051_.n21 _051_.t18 131.748
R30792 _051_.n10 _051_.t17 121.109
R30793 _051_.n27 _051_.n2 105.677
R30794 _051_.n5 _051_.n4 105.677
R30795 _051_.n22 _051_.n21 90.6325
R30796 _051_.n10 _051_ 80.3299
R30797 _051_ _051_.n6 78.065
R30798 _051_.n12 _051_.n11 76.0005
R30799 _051_.n11 _051_.n10 40.9982
R30800 _051_.n3 _051_.t1 26.5955
R30801 _051_.n3 _051_.t0 26.5955
R30802 _051_.n1 _051_.t2 26.5955
R30803 _051_.n1 _051_.t4 26.5955
R30804 _051_.n26 _051_.t3 26.5955
R30805 _051_.n26 _051_.t5 26.5955
R30806 _051_.n2 _051_.t11 24.9236
R30807 _051_.n2 _051_.t7 24.9236
R30808 _051_.n4 _051_.t9 24.9236
R30809 _051_.n4 _051_.t8 24.9236
R30810 _051_.n0 _051_.t10 24.9236
R30811 _051_.n0 _051_.t6 24.9236
R30812 _051_.n24 _051_.n23 21.002
R30813 _051_.n23 _051_.n20 17.4031
R30814 _051_.n7 _051_ 15.4844
R30815 _051_.n24 _051_ 15.1152
R30816 _051_.n16 _051_ 14.1338
R30817 _051_.n14 _051_.n9 12.5079
R30818 _051_.n27 _051_.n25 12.0732
R30819 _051_.n15 _051_.n14 10.7295
R30820 _051_.n25 _051_.n24 10.1118
R30821 _051_.n12 _051_ 9.6005
R30822 _051_.n13 _051_ 9.6005
R30823 _051_.n9 _051_.n8 9.47703
R30824 _051_.n14 _051_.n13 9.44462
R30825 _051_.n20 _051_.n19 9.3005
R30826 _051_.n19 _051_.n18 7.13769
R30827 _051_ _051_.n27 5.96414
R30828 _051_.n9 _051_ 5.25872
R30829 _051_.n23 _051_.n22 4.6505
R30830 _051_.n15 _051_.n7 4.58328
R30831 _051_.n7 _051_ 3.51018
R30832 _051_ _051_.n12 3.2005
R30833 _051_.n13 _051_ 3.2005
R30834 _051_ _051_.n15 2.78292
R30835 _051_.n17 _051_.n16 2.4005
R30836 _051_.n20 _051_.n17 2.13383
R30837 _051_.n22 _051_ 1.23686
R30838 _051_.n25 _051_.n5 0.145955
R30839 trimb[2].n9 trimb[2].n8 349.738
R30840 trimb[2].n11 trimb[2].n10 292.5
R30841 trimb[2].n11 trimb[2].n4 292.5
R30842 trimb[2].n13 trimb[2].n3 193.387
R30843 trimb[2].n7 trimb[2].n5 151.127
R30844 trimb[2].n7 trimb[2].n6 107.763
R30845 trimb[2].n5 trimb[2].t4 40.0005
R30846 trimb[2].n5 trimb[2].t6 40.0005
R30847 trimb[2].n6 trimb[2].t5 40.0005
R30848 trimb[2].n6 trimb[2].t7 40.0005
R30849 trimb[2].n8 trimb[2].t2 27.5805
R30850 trimb[2].n8 trimb[2].t0 27.5805
R30851 trimb[2].n12 trimb[2].t3 23.6405
R30852 trimb[2].n3 trimb[2].t1 23.1644
R30853 trimb[2].n10 trimb[2].n9 14.7697
R30854 trimb[2].n4 trimb[2].n2 11.243
R30855 trimb[2] trimb[2].n7 10.4115
R30856 trimb[2].n13 trimb[2].n1 9.3005
R30857 trimb[2].n14 trimb[2].n13 9.3005
R30858 trimb[2].n13 trimb[2].n12 9.3005
R30859 trimb[2].n14 trimb[2].n0 9.04377
R30860 trimb[2].n1 trimb[2].n0 9.01973
R30861 trimb[2].n11 trimb[2].n3 4.23401
R30862 trimb[2].n15 trimb[2].n2 4.13041
R30863 trimb[2].n12 trimb[2].n11 3.9405
R30864 trimb[2].n13 trimb[2].n2 3.09077
R30865 trimb[2] trimb[2].n16 2.48707
R30866 trimb[2].n16 trimb[2].n15 2.24426
R30867 trimb[2].n9 trimb[2].n4 1.96973
R30868 trimb[2].n10 trimb[2] 0.246654
R30869 trimb[2].n15 trimb[2].n1 0.03175
R30870 trimb[2].n16 trimb[2].n0 0.0141816
R30871 trimb[2].n15 trimb[2].n14 0.0101154
R30872 trimb[1].n9 trimb[1].n8 349.738
R30873 trimb[1].n11 trimb[1].n10 292.5
R30874 trimb[1].n11 trimb[1].n4 292.5
R30875 trimb[1].n13 trimb[1].n3 193.387
R30876 trimb[1].n7 trimb[1].n5 151.127
R30877 trimb[1].n7 trimb[1].n6 107.763
R30878 trimb[1].n5 trimb[1].t4 40.0005
R30879 trimb[1].n5 trimb[1].t6 40.0005
R30880 trimb[1].n6 trimb[1].t5 40.0005
R30881 trimb[1].n6 trimb[1].t7 40.0005
R30882 trimb[1].n8 trimb[1].t1 27.5805
R30883 trimb[1].n8 trimb[1].t2 27.5805
R30884 trimb[1].n12 trimb[1].t3 23.6405
R30885 trimb[1].n3 trimb[1].t0 23.1644
R30886 trimb[1].n10 trimb[1].n9 14.7697
R30887 trimb[1].n4 trimb[1].n2 11.243
R30888 trimb[1] trimb[1].n7 10.4115
R30889 trimb[1].n13 trimb[1].n1 9.3005
R30890 trimb[1].n14 trimb[1].n13 9.3005
R30891 trimb[1].n13 trimb[1].n12 9.3005
R30892 trimb[1].n14 trimb[1].n0 9.04377
R30893 trimb[1].n1 trimb[1].n0 9.01973
R30894 trimb[1].n11 trimb[1].n3 4.23401
R30895 trimb[1].n15 trimb[1].n2 4.13041
R30896 trimb[1].n12 trimb[1].n11 3.9405
R30897 trimb[1].n13 trimb[1].n2 3.09077
R30898 trimb[1] trimb[1].n16 2.48707
R30899 trimb[1].n16 trimb[1].n15 2.24426
R30900 trimb[1].n9 trimb[1].n4 1.96973
R30901 trimb[1].n10 trimb[1] 0.246654
R30902 trimb[1].n15 trimb[1].n1 0.03175
R30903 trimb[1].n16 trimb[1].n0 0.0141816
R30904 trimb[1].n15 trimb[1].n14 0.0101154
R30905 ctln[0].n3 ctln[0].n2 143.643
R30906 ctln[0].n4 ctln[0] 81.5159
R30907 ctln[0].n2 ctln[0].t1 26.5955
R30908 ctln[0].n2 ctln[0].t0 26.5955
R30909 ctln[0].n1 ctln[0].t3 24.9236
R30910 ctln[0].n1 ctln[0].n0 15.6928
R30911 ctln[0].n0 ctln[0].t2 9.23127
R30912 ctln[0] ctln[0].n3 9.02598
R30913 ctln[0].n4 ctln[0].n1 8.25053
R30914 ctln[0].n3 ctln[0] 7.64268
R30915 ctln[0].n8 ctln[0] 4.18004
R30916 ctln[0].n11 ctln[0].n10 3.79439
R30917 ctln[0].n10 ctln[0].n8 2.24426
R30918 ctln[0] ctln[0].n11 2.08974
R30919 ctln[0].n11 ctln[0].n5 2.03855
R30920 ctln[0].n5 ctln[0].n4 0.214619
R30921 ctln[0].n10 ctln[0].n6 0.0389615
R30922 ctln[0].n8 ctln[0].n7 0.0141816
R30923 ctln[0].n10 ctln[0].n9 0.00290385
R30924 trim[4].n9 trim[4].n8 349.738
R30925 trim[4].n11 trim[4].n10 292.5
R30926 trim[4].n11 trim[4].n4 292.5
R30927 trim[4].n13 trim[4].n3 193.387
R30928 trim[4].n7 trim[4].n5 151.127
R30929 trim[4].n7 trim[4].n6 107.763
R30930 trim[4].n5 trim[4].t7 40.0005
R30931 trim[4].n5 trim[4].t4 40.0005
R30932 trim[4].n6 trim[4].t5 40.0005
R30933 trim[4].n6 trim[4].t6 40.0005
R30934 trim[4].n8 trim[4].t3 27.5805
R30935 trim[4].n8 trim[4].t0 27.5805
R30936 trim[4].n12 trim[4].t1 23.6405
R30937 trim[4].n3 trim[4].t2 23.1644
R30938 trim[4].n10 trim[4].n9 14.7697
R30939 trim[4].n4 trim[4].n2 11.243
R30940 trim[4] trim[4].n7 10.4115
R30941 trim[4].n13 trim[4].n1 9.3005
R30942 trim[4].n14 trim[4].n13 9.3005
R30943 trim[4].n13 trim[4].n12 9.3005
R30944 trim[4].n14 trim[4].n0 9.04377
R30945 trim[4].n1 trim[4].n0 9.01973
R30946 trim[4].n11 trim[4].n3 4.23401
R30947 trim[4].n15 trim[4].n2 4.13041
R30948 trim[4].n12 trim[4].n11 3.9405
R30949 trim[4].n13 trim[4].n2 3.09077
R30950 trim[4] trim[4].n16 2.48707
R30951 trim[4].n16 trim[4].n15 2.24426
R30952 trim[4].n9 trim[4].n4 1.96973
R30953 trim[4].n10 trim[4] 0.246654
R30954 trim[4].n15 trim[4].n1 0.03175
R30955 trim[4].n16 trim[4].n0 0.0141816
R30956 trim[4].n15 trim[4].n14 0.0101154
R30957 valid.n5 valid.n4 354.634
R30958 valid.n7 valid.n6 151.127
R30959 valid.n5 valid.n3 96.9298
R30960 valid.n2 valid.t4 41.7262
R30961 valid.n6 valid.t6 40.0005
R30962 valid.n6 valid.t7 40.0005
R30963 valid.n2 valid.t5 35.4961
R30964 valid.n3 valid.t0 27.5805
R30965 valid.n3 valid.t1 27.5805
R30966 valid.n4 valid.t2 27.5805
R30967 valid.n4 valid.t3 27.5805
R30968 valid.n8 valid.n7 15.262
R30969 valid.n7 valid 10.4115
R30970 valid valid.n5 9.6475
R30971 valid.n9 valid.n8 9.3005
R30972 valid.n9 valid.n0 9.01973
R30973 valid.n11 valid.n10 9.0005
R30974 valid.n8 valid.n2 7.31891
R30975 valid.n8 valid.n1 4.5765
R30976 valid valid.n11 4.23171
R30977 valid.n1 valid.n0 2.25706
R30978 valid.n11 valid.n0 0.0509808
R30979 valid.n10 valid.n9 0.0341538
R30980 valid.n10 valid.n1 0.00200872
R30981 trim[3].n9 trim[3].n8 349.738
R30982 trim[3].n11 trim[3].n10 292.5
R30983 trim[3].n11 trim[3].n4 292.5
R30984 trim[3].n13 trim[3].n3 193.387
R30985 trim[3].n7 trim[3].n5 151.127
R30986 trim[3].n7 trim[3].n6 107.763
R30987 trim[3].n5 trim[3].t7 40.0005
R30988 trim[3].n5 trim[3].t4 40.0005
R30989 trim[3].n6 trim[3].t5 40.0005
R30990 trim[3].n6 trim[3].t6 40.0005
R30991 trim[3].n8 trim[3].t0 27.5805
R30992 trim[3].n8 trim[3].t1 27.5805
R30993 trim[3].n12 trim[3].t2 23.6405
R30994 trim[3].n3 trim[3].t3 23.1644
R30995 trim[3].n10 trim[3].n9 14.7697
R30996 trim[3].n4 trim[3].n2 11.243
R30997 trim[3] trim[3].n7 10.4115
R30998 trim[3].n13 trim[3].n1 9.3005
R30999 trim[3].n14 trim[3].n13 9.3005
R31000 trim[3].n13 trim[3].n12 9.3005
R31001 trim[3].n14 trim[3].n0 9.04377
R31002 trim[3].n1 trim[3].n0 9.01973
R31003 trim[3].n11 trim[3].n3 4.23401
R31004 trim[3].n15 trim[3].n2 4.13041
R31005 trim[3].n12 trim[3].n11 3.9405
R31006 trim[3].n13 trim[3].n2 3.09077
R31007 trim[3] trim[3].n16 2.48707
R31008 trim[3].n16 trim[3].n15 2.24426
R31009 trim[3].n9 trim[3].n4 1.96973
R31010 trim[3].n10 trim[3] 0.246654
R31011 trim[3].n15 trim[3].n1 0.03175
R31012 trim[3].n16 trim[3].n0 0.0141816
R31013 trim[3].n15 trim[3].n14 0.0101154
R31014 result[0].n6 result[0] 585.251
R31015 result[0].n8 result[0].n7 585
R31016 result[0].n6 result[0].n5 292.5
R31017 result[0] result[0].n4 95.7632
R31018 result[0].n5 result[0] 79.5613
R31019 result[0].n6 result[0].t0 26.5955
R31020 result[0].n4 result[0].t3 24.9236
R31021 result[0].n4 result[0].t2 24.9236
R31022 result[0].n7 result[0].n6 16.7455
R31023 result[0] result[0].n2 10.4588
R31024 result[0].n7 result[0].t1 9.8505
R31025 result[0].n8 result[0].n1 9.3005
R31026 result[0].n9 result[0].n8 9.3005
R31027 result[0].n6 result[0].n3 9.1516
R31028 result[0].n9 result[0].n0 9.05098
R31029 result[0].n1 result[0].n0 9.01252
R31030 result[0].n5 result[0] 7.02795
R31031 result[0] result[0].n3 4.01265
R31032 result[0].n10 result[0].n2 3.75172
R31033 result[0] result[0].n11 2.45104
R31034 result[0].n11 result[0].n10 2.24426
R31035 result[0].n8 result[0].n2 1.87152
R31036 result[0].n10 result[0].n1 0.0389615
R31037 result[0].n11 result[0].n0 0.0141816
R31038 result[0].n8 result[0].n3 0.00492585
R31039 result[0].n10 result[0].n9 0.00290385
R31040 ctln[5].n1 ctln[5].n0 143.643
R31041 ctln[5].n2 ctln[5] 79.4173
R31042 ctln[5].n0 ctln[5].t1 26.5955
R31043 ctln[5].n0 ctln[5].t0 26.5955
R31044 ctln[5].n5 ctln[5].t3 24.0005
R31045 ctln[5].n4 ctln[5].n3 14.7697
R31046 ctln[5].n3 ctln[5].t2 10.1543
R31047 ctln[5].n6 ctln[5].n5 9.3005
R31048 ctln[5] ctln[5].n1 9.02598
R31049 ctln[5].n1 ctln[5] 7.64268
R31050 ctln[5].n7 ctln[5] 7.373
R31051 ctln[5] ctln[5].n7 2.82782
R31052 ctln[5].n6 ctln[5].n2 2.36635
R31053 ctln[5].n5 ctln[5].n4 0.923577
R31054 ctln[5].n7 ctln[5].n6 0.905693
R31055 ctlp[5].n4 ctlp[5].n1 292.5
R31056 ctlp[5].n3 ctlp[5].n2 92.5005
R31057 ctlp[5] ctlp[5].n3 81.3181
R31058 ctlp[5].n1 ctlp[5].t0 26.5955
R31059 ctlp[5].n0 ctlp[5].t1 25.8903
R31060 ctlp[5].n2 ctlp[5].t2 24.9236
R31061 ctlp[5].n2 ctlp[5].t3 24.9236
R31062 ctlp[5] ctlp[5].n4 15.5613
R31063 ctlp[5].n6 ctlp[5] 10.1093
R31064 ctlp[5].n5 ctlp[5].n0 9.48617
R31065 ctlp[5].n3 ctlp[5] 5.27109
R31066 ctlp[5].n5 ctlp[5] 2.60833
R31067 ctlp[5] ctlp[5].n5 1.85252
R31068 ctlp[5].n4 ctlp[5] 1.50638
R31069 ctlp[5].n1 ctlp[5].n0 0.248635
R31070 ctlp[5].n6 ctlp[5] 0.0788333
R31071 ctlp[5] ctlp[5].n6 0.0129779
R31072 ctln[2].n1 ctln[2].n0 143.643
R31073 ctln[2].n2 ctln[2] 79.4173
R31074 ctln[2].n0 ctln[2].t1 26.5955
R31075 ctln[2].n0 ctln[2].t0 26.5955
R31076 ctln[2].n5 ctln[2].t2 24.0005
R31077 ctln[2].n4 ctln[2].n3 14.7697
R31078 ctln[2].n7 ctln[2] 10.7299
R31079 ctln[2].n3 ctln[2].t3 10.1543
R31080 ctln[2].n6 ctln[2].n5 9.3005
R31081 ctln[2] ctln[2].n1 9.02598
R31082 ctln[2].n1 ctln[2] 7.64268
R31083 ctln[2] ctln[2].n7 2.82364
R31084 ctln[2].n6 ctln[2].n2 2.36635
R31085 ctln[2].n5 ctln[2].n4 0.923577
R31086 ctln[2].n7 ctln[2].n6 0.910763
R31087 ctln[7].n2 ctln[7].n0 354.634
R31088 ctln[7].n7 ctln[7].n4 107.763
R31089 ctln[7].n2 ctln[7].n1 96.9298
R31090 ctln[7].n7 ctln[7].n6 58.6278
R31091 ctln[7].n5 ctln[7].t4 40.3946
R31092 ctln[7].n4 ctln[7].t6 40.0005
R31093 ctln[7].n4 ctln[7].t7 40.0005
R31094 ctln[7].n5 ctln[7].t5 36.871
R31095 ctln[7].n1 ctln[7].t0 27.5805
R31096 ctln[7].n1 ctln[7].t1 27.5805
R31097 ctln[7].n0 ctln[7].t2 27.5805
R31098 ctln[7].n0 ctln[7].t3 27.5805
R31099 ctln[7] ctln[7].n3 19.2609
R31100 ctln[7].n3 ctln[7].n2 15.309
R31101 ctln[7].n6 ctln[7] 12.9442
R31102 ctln[7].n8 ctln[7] 9.00791
R31103 ctln[7].n6 ctln[7].n5 7.36486
R31104 ctln[7].n8 ctln[7].n7 6.77697
R31105 ctln[7].n3 ctln[7] 2.70819
R31106 ctln[7] ctln[7].n8 1.73877
R31107 net37.n0 net37.t4 238.59
R31108 net37.n0 net37.t5 203.244
R31109 net37.n7 net37.n6 111.322
R31110 net37.n1 net37.n0 76.0005
R31111 net37 net37.n2 38.4012
R31112 net37.n6 net37.t0 26.5955
R31113 net37.n6 net37.t1 26.5955
R31114 net37.n3 net37.t3 24.9236
R31115 net37.n3 net37.t2 24.9236
R31116 net37 net37.n5 11.2645
R31117 net37 net37.n4 8.65445
R31118 net37.n4 net37.n3 8.343
R31119 net37.n1 net37 8.22907
R31120 net37.n5 net37 6.1445
R31121 net37.n5 net37 4.65505
R31122 net37.n4 net37 3.69206
R31123 net37.n2 net37 3.10907
R31124 net37.n7 net37 2.0485
R31125 net37 net37.n7 1.55202
R31126 net37.n2 net37.n1 1.09764
R31127 ctlp[0].n16 ctlp[0].n4 349.738
R31128 ctlp[0].n2 ctlp[0].n0 151.127
R31129 ctlp[0].n2 ctlp[0].n1 107.763
R31130 ctlp[0].n0 ctlp[0].t6 40.0005
R31131 ctlp[0].n0 ctlp[0].t4 40.0005
R31132 ctlp[0].n1 ctlp[0].t5 40.0005
R31133 ctlp[0].n1 ctlp[0].t7 40.0005
R31134 ctlp[0].n4 ctlp[0].t2 27.5805
R31135 ctlp[0].n4 ctlp[0].t0 27.5805
R31136 ctlp[0].n7 ctlp[0].t3 23.6405
R31137 ctlp[0].n5 ctlp[0].t1 23.1644
R31138 ctlp[0].n18 ctlp[0] 19.2609
R31139 ctlp[0].n17 ctlp[0].n16 14.7697
R31140 ctlp[0].n15 ctlp[0].n14 11.243
R31141 ctlp[0].n8 ctlp[0].n7 9.3005
R31142 ctlp[0] ctlp[0].n3 9.00791
R31143 ctlp[0].n3 ctlp[0].n2 6.77697
R31144 ctlp[0].n18 ctlp[0].n17 5.90819
R31145 ctlp[0].n6 ctlp[0].n5 4.23401
R31146 ctlp[0].n14 ctlp[0].n13 4.13041
R31147 ctlp[0].n7 ctlp[0].n6 3.9405
R31148 ctlp[0].n9 ctlp[0] 3.38228
R31149 ctlp[0].n14 ctlp[0].n8 3.09077
R31150 ctlp[0] ctlp[0].n18 2.70819
R31151 ctlp[0].n11 ctlp[0].n10 2.25561
R31152 ctlp[0].n16 ctlp[0].n15 1.96973
R31153 ctlp[0].n3 ctlp[0] 1.73877
R31154 ctlp[0].n10 ctlp[0].n9 0.0509808
R31155 ctlp[0].n13 ctlp[0].n12 0.03175
R31156 ctlp[0].n13 ctlp[0].n11 0.00339788
R31157 _062_.n24 _062_.t15 471.289
R31158 _062_.n28 _062_.t12 334.723
R31159 _062_.n21 _062_.t17 238.858
R31160 _062_.n15 _062_.t9 232.446
R31161 _062_.n10 _062_.t10 212.081
R31162 _062_.n11 _062_.t18 212.081
R31163 _062_.n28 _062_.t16 206.19
R31164 _062_.n7 _062_.n6 183.22
R31165 _062_.n14 _062_.t11 159.381
R31166 _062_.n19 _062_.t19 156.739
R31167 _062_.n9 _062_.n8 153.805
R31168 _062_.n7 _062_.n5 153.548
R31169 _062_.n19 _062_ 152.785
R31170 _062_.n20 _062_.n18 152
R31171 _062_.n24 _062_.t13 148.35
R31172 _062_ _062_.n4 141.07
R31173 _062_.n10 _062_.t14 139.78
R31174 _062_.n11 _062_.t8 139.78
R31175 _062_.n13 _062_.n12 102.561
R31176 _062_.n9 _062_.n7 79.8031
R31177 _062_.n29 _062_.n28 76.0005
R31178 _062_.n25 _062_.n24 76.0005
R31179 _062_.n14 _062_ 48.5769
R31180 _062_.n12 _062_.n10 38.7066
R31181 _062_.n26 _062_.n25 36.5315
R31182 _062_.n5 _062_.t7 26.5955
R31183 _062_.n5 _062_.t6 26.5955
R31184 _062_.n8 _062_.t2 26.5955
R31185 _062_.n8 _062_.t3 26.5955
R31186 _062_.n6 _062_.t1 26.5955
R31187 _062_.n6 _062_.t0 26.5955
R31188 _062_.n4 _062_.t4 24.9236
R31189 _062_.n4 _062_.t5 24.9236
R31190 _062_.n31 _062_.n9 23.2732
R31191 _062_.n12 _062_.n11 22.6399
R31192 _062_.n30 _062_.n29 20.2667
R31193 _062_.n29 _062_ 14.4462
R31194 _062_.n25 _062_ 13.7314
R31195 _062_ _062_.n31 13.2078
R31196 _062_.n20 _062_.n19 12.4968
R31197 _062_.n23 _062_ 11.2153
R31198 _062_.n3 _062_.n2 0.0138153
R31199 _062_.n22 _062_.n3 4.64889
R31200 _062_.n16 _062_.n15 9.3005
R31201 _062_.n27 _062_.n17 9.1834
R31202 _062_.n2 _062_.n26 9.0005
R31203 _062_.n30 _062_.n27 8.97028
R31204 _062_.n22 _062_.n21 8.76429
R31205 _062_.n27 _062_.n1 7.39146
R31206 _062_.n13 _062_ 5.1205
R31207 _062_.n31 _062_.n30 4.83846
R31208 _062_.n17 _062_.n13 4.58329
R31209 _062_.n15 _062_.n14 4.36393
R31210 _062_ _062_.n16 4.288
R31211 _062_.n2 _062_.n23 3.81297
R31212 _062_.n2 _062_.n1 2.24013
R31213 _062_ _062_.n18 2.87397
R31214 _062_.n21 _062_.n20 2.67828
R31215 _062_.n17 _062_ 2.5166
R31216 _062_.n23 _062_.n22 2.2837
R31217 _062_.n16 _062_ 1.55202
R31218 _062_.n22 _062_.n18 0.784173
R31219 _062_.n1 _062_.n0 0.0141573
R31220 _062_.n26 _062_.n0 0.0509808
R31221 _062_.n3 _062_.n0 9.04985
R31222 net20.t0 net20 459.913
R31223 net20.n1 net20.t0 440.25
R31224 net20.n2 net20.t5 238.59
R31225 net20.n4 net20.t3 212.081
R31226 net20.n5 net20.t4 212.081
R31227 net20.n2 net20.t2 203.244
R31228 net20.n4 net20.t6 139.78
R31229 net20.n5 net20.t7 139.78
R31230 net20 net20.n8 79.0438
R31231 net20 net20.n2 78.0119
R31232 net20.n5 net20.n4 61.346
R31233 net20.n0 net20.n5 40.2726
R31234 net20.n8 net20.t1 38.6168
R31235 net20.n1 net20 10.9042
R31236 net20.n3 net20 9.32621
R31237 net20.n6 net20.n3 5.50712
R31238 net20 net20.n1 5.21532
R31239 net20.n0 net20 3.17119
R31240 net20.n3 net20 3.10907
R31241 net20.n7 net20 2.78389
R31242 net20.n7 net20 2.77331
R31243 net20.n8 net20.n7 1.13595
R31244 net20 net20.n6 0.858673
R31245 net20.n0 net20.n6 12.0761
R31246 _110_.n4 _110_.t4 260.384
R31247 _110_.n11 _110_.t2 256.07
R31248 _110_.n1 _110_.t5 256.07
R31249 _110_.n6 _110_.t6 256.07
R31250 _110_.n14 _110_.t0 188.135
R31251 _110_.n4 _110_.t8 156.468
R31252 _110_.n11 _110_.t9 150.03
R31253 _110_.n1 _110_.t7 150.03
R31254 _110_.n6 _110_.t3 150.03
R31255 _110_.n0 _110_.t1 130.641
R31256 _110_.n12 _110_.n11 76.0005
R31257 _110_.n2 _110_.n1 76.0005
R31258 _110_.n7 _110_.n6 76.0005
R31259 _110_.n14 _110_.n13 28.0855
R31260 _110_.n9 _110_.n8 27.6795
R31261 _110_.n13 _110_ 25.7725
R31262 _110_.n10 _110_.n3 20.5235
R31263 _110_.n13 _110_ 16.8988
R31264 _110_.n7 _110_ 16.3845
R31265 _110_.n10 _110_.n9 10.7607
R31266 _110_.n9 _110_.n5 9.19185
R31267 _110_ _110_.n12 8.23114
R31268 _110_.n5 _110_.n4 7.99433
R31269 _110_.n12 _110_ 7.6805
R31270 _110_.n2 _110_ 7.6805
R31271 _110_.n3 _110_.n2 4.6085
R31272 _110_.n8 _110_.n7 4.6085
R31273 _110_.n3 _110_ 4.58918
R31274 _110_.n8 _110_ 4.58918
R31275 _110_.n0 _110_ 4.47034
R31276 _110_ _110_.n14 3.55533
R31277 _110_ _110_.n0 2.63228
R31278 _110_.n5 _110_ 2.39384
R31279 _110_ _110_.n10 1.77494
R31280 ctlp[2].n7 ctlp[2].n6 92.5005
R31281 ctlp[2] ctlp[2].n7 81.3181
R31282 ctlp[2].n2 ctlp[2].t0 25.6105
R31283 ctlp[2].n6 ctlp[2].t3 24.9236
R31284 ctlp[2].n6 ctlp[2].t2 24.9236
R31285 ctlp[2].n0 ctlp[2].t1 21.1429
R31286 ctlp[2] ctlp[2].n8 15.5613
R31287 ctlp[2].n3 ctlp[2].n2 9.3005
R31288 ctlp[2].n7 ctlp[2] 5.27109
R31289 ctlp[2].n1 ctlp[2].n0 5.17648
R31290 ctlp[2].n5 ctlp[2] 5.02021
R31291 ctlp[2] ctlp[2].n4 3.63219
R31292 ctlp[2] ctlp[2].n5 2.60941
R31293 ctlp[2].n8 ctlp[2] 1.50638
R31294 ctlp[2].n2 ctlp[2].n1 0.9855
R31295 ctlp[2].n5 ctlp[2].n3 0.84894
R31296 ctlp[2].n4 ctlp[2] 0.0788333
R31297 ctlp[2].n4 ctlp[2] 0.0129779
R31298 trimb[3].n2 trimb[3].n0 585
R31299 trimb[3].n11 trimb[3].n4 349.738
R31300 trimb[3].n10 trimb[3].n3 292.5
R31301 trimb[3].n12 trimb[3].n3 292.5
R31302 trimb[3].n7 trimb[3].n5 151.127
R31303 trimb[3].n7 trimb[3].n6 107.763
R31304 trimb[3].n5 trimb[3].t4 40.0005
R31305 trimb[3].n5 trimb[3].t6 40.0005
R31306 trimb[3].n6 trimb[3].t5 40.0005
R31307 trimb[3].n6 trimb[3].t7 40.0005
R31308 trimb[3].n4 trimb[3].t2 27.5805
R31309 trimb[3].n4 trimb[3].t0 27.5805
R31310 trimb[3].n1 trimb[3].t3 23.7598
R31311 trimb[3].n9 trimb[3] 19.2609
R31312 trimb[3].n2 trimb[3].t1 14.7755
R31313 trimb[3].n11 trimb[3].n10 14.7697
R31314 trimb[3].n3 trimb[3].n2 12.8055
R31315 trimb[3].n13 trimb[3].n12 12.3259
R31316 trimb[3] trimb[3].n8 9.00791
R31317 trimb[3].n1 trimb[3].n0 8.9018
R31318 trimb[3].n8 trimb[3].n7 6.77697
R31319 trimb[3].n10 trimb[3].n9 5.90819
R31320 trimb[3].n3 trimb[3].n1 3.77188
R31321 trimb[3].n9 trimb[3] 2.70819
R31322 trimb[3].n12 trimb[3].n11 1.96973
R31323 trimb[3] trimb[3].n13 1.77665
R31324 trimb[3].n8 trimb[3] 1.73877
R31325 trimb[3].n13 trimb[3].n0 1.20582
R31326 clk.n0 clk.t4 184.768
R31327 clk.n1 clk.t2 184.768
R31328 clk.n2 clk.t1 184.768
R31329 clk.n3 clk.t0 184.768
R31330 clk.n0 clk.t7 146.208
R31331 clk.n1 clk.t6 146.208
R31332 clk.n2 clk.t5 146.208
R31333 clk.n3 clk.t3 146.208
R31334 clk clk.n3 97.6099
R31335 clk clk.n4 60.0555
R31336 clk.n1 clk.n0 40.6397
R31337 clk.n2 clk.n1 40.6397
R31338 clk.n3 clk.n2 40.6397
R31339 clk.n4 clk 10.3624
R31340 clk.n4 clk 3.45447
R31341 ctln[1].n1 ctln[1].n0 143.643
R31342 ctln[1].n2 ctln[1] 79.4173
R31343 ctln[1].n0 ctln[1].t0 26.5955
R31344 ctln[1].n0 ctln[1].t1 26.5955
R31345 ctln[1].n5 ctln[1].t2 24.0005
R31346 ctln[1].n4 ctln[1].n3 14.7697
R31347 ctln[1].n3 ctln[1].t3 10.1543
R31348 ctln[1].n6 ctln[1].n5 9.3005
R31349 ctln[1] ctln[1].n1 9.02598
R31350 ctln[1].n1 ctln[1] 7.64268
R31351 ctln[1].n7 ctln[1] 7.38553
R31352 ctln[1] ctln[1].n7 2.82782
R31353 ctln[1].n6 ctln[1].n2 2.36635
R31354 ctln[1].n5 ctln[1].n4 0.923577
R31355 ctln[1].n7 ctln[1].n6 0.905693
R31356 ctlp[3].n6 ctlp[3].n5 92.5005
R31357 ctlp[3] ctlp[3].n6 81.3181
R31358 ctlp[3].n2 ctlp[3].t0 25.6105
R31359 ctlp[3].n5 ctlp[3].t3 24.9236
R31360 ctlp[3].n5 ctlp[3].t2 24.9236
R31361 ctlp[3].n0 ctlp[3].t1 21.1429
R31362 ctlp[3] ctlp[3].n7 15.5613
R31363 ctlp[3].n3 ctlp[3].n2 9.3005
R31364 ctlp[3].n4 ctlp[3] 5.32379
R31365 ctlp[3].n6 ctlp[3] 5.27109
R31366 ctlp[3].n1 ctlp[3].n0 5.17648
R31367 ctlp[3] ctlp[3].n4 2.60941
R31368 ctlp[3].n7 ctlp[3] 1.50638
R31369 ctlp[3].n2 ctlp[3].n1 0.9855
R31370 ctlp[3].n4 ctlp[3].n3 0.84894
R31371 _042_.n2 _042_.t2 259.027
R31372 _042_.n3 _042_.t0 188.135
R31373 _042_.n2 _042_.t3 175.782
R31374 _042_.n1 _042_.t1 130.641
R31375 _042_.n3 _042_ 13.9349
R31376 _042_ _042_.n0 57.1727
R31377 _042_.n0 _042_.n2 8.25129
R31378 _042_.n1 _042_ 4.47034
R31379 _042_ _042_.n3 3.55533
R31380 _042_ _042_.n1 2.63228
R31381 _042_ _042_.n0 2.2524
R31382 ctln[4].n8 ctln[4].n7 185
R31383 ctln[4].n4 ctln[4].n3 143.643
R31384 ctln[4].n5 ctln[4] 81.5159
R31385 ctln[4].n3 ctln[4].t1 26.5955
R31386 ctln[4].n3 ctln[4].t0 26.5955
R31387 ctln[4].n6 ctln[4].t3 24.9236
R31388 ctln[4].n7 ctln[4].n6 15.6928
R31389 ctln[4].n8 ctln[4].n1 9.3005
R31390 ctln[4].n9 ctln[4].n8 9.3005
R31391 ctln[4].n7 ctln[4].t2 9.23127
R31392 ctln[4].n9 ctln[4].n0 9.05098
R31393 ctln[4] ctln[4].n4 9.02598
R31394 ctln[4].n1 ctln[4].n0 9.01252
R31395 ctln[4].n6 ctln[4].n5 8.25053
R31396 ctln[4].n4 ctln[4] 7.64268
R31397 ctln[4].n10 ctln[4].n2 3.79439
R31398 ctln[4] ctln[4].n11 3.17386
R31399 ctln[4].n11 ctln[4].n10 2.24426
R31400 ctln[4].n2 ctln[4] 2.08974
R31401 ctln[4].n8 ctln[4].n2 2.03855
R31402 ctln[4].n8 ctln[4].n5 0.214619
R31403 ctln[4].n12 ctln[4] 0.0747105
R31404 ctln[4].n10 ctln[4].n1 0.0389615
R31405 ctln[4].n11 ctln[4].n0 0.0141816
R31406 ctln[4] ctln[4].n12 0.0105337
R31407 ctln[4].n12 ctln[4] 0.00842135
R31408 ctln[4].n10 ctln[4].n9 0.00290385
R31409 net4.t0 net4.n10 440.25
R31410 net4.n12 net4.t7 275.267
R31411 net4.n2 net4.t5 238.59
R31412 net4.n7 net4.t3 222.725
R31413 net4.n2 net4.t2 203.244
R31414 net4.n12 net4.t4 196.74
R31415 net4.n5 net4.t6 177.171
R31416 net4.n5 net4.n4 152
R31417 net4.n6 net4.n3 152
R31418 net4.n11 net4.t0 135.105
R31419 net4.n9 net4.t1 123.654
R31420 net4 net4.n9 78.8791
R31421 net4 net4.n2 78.0119
R31422 net4.n16 net4.n0 28.5515
R31423 net4.n0 net4.n11 29.3078
R31424 net4.n10 net4 10.9042
R31425 net4.n16 net4 10.8096
R31426 net4.n6 net4.n5 10.5442
R31427 net4.n17 net4 9.32621
R31428 net4.n1 net4 24.4766
R31429 net4 net4.n1 2.27879
R31430 net4.n8 net4.n7 8.76429
R31431 net4.n17 net4.n16 7.40891
R31432 net4.n13 net4.n12 7.35429
R31433 net4.n4 net4 5.51161
R31434 net4.n10 net4 5.21532
R31435 net4.n9 net4 5.16973
R31436 net4.n0 net4.n15 4.56795
R31437 net4.n11 net4 4.06431
R31438 net4 net4.n17 3.10907
R31439 net4.n4 net4.n3 2.48939
R31440 net4.n7 net4.n6 2.25988
R31441 net4.n15 net4.n14 2.24915
R31442 net4.n8 net4.n1 0.729716
R31443 net4.n15 net4.n13 0.692392
R31444 net4.n14 net4 0.692392
R31445 net4.n8 net4.n3 0.533833
R31446 clkc.t0 clkc.n3 440.25
R31447 clkc.n4 clkc.t0 133.882
R31448 clkc clkc.t1 126.855
R31449 clkc.n3 clkc 80.894
R31450 clkc clkc.n2 11.0668
R31451 clkc.n5 clkc.n1 9.3005
R31452 clkc.n6 clkc.n5 9.3005
R31453 clkc.n6 clkc.n0 9.04617
R31454 clkc.n1 clkc.n0 9.01733
R31455 clkc.n7 clkc.n2 4.14532
R31456 clkc.n5 clkc.n2 2.97937
R31457 clkc.n3 clkc 2.84494
R31458 clkc clkc.n8 2.45104
R31459 clkc.n8 clkc.n7 2.24426
R31460 clkc.n4 clkc 1.83668
R31461 clkc.n5 clkc.n4 0.0512129
R31462 clkc.n7 clkc.n1 0.0341538
R31463 clkc.n8 clkc.n0 0.0141816
R31464 clkc.n7 clkc.n6 0.00771154
R31465 ctln[3].n1 ctln[3].n0 143.643
R31466 ctln[3].n2 ctln[3] 79.4173
R31467 ctln[3].n0 ctln[3].t1 26.5955
R31468 ctln[3].n0 ctln[3].t0 26.5955
R31469 ctln[3].n5 ctln[3].t2 24.0005
R31470 ctln[3].n4 ctln[3].n3 14.7697
R31471 ctln[3].n3 ctln[3].t3 10.1543
R31472 ctln[3].n6 ctln[3].n5 9.3005
R31473 ctln[3] ctln[3].n1 9.02598
R31474 ctln[3].n1 ctln[3] 7.64268
R31475 ctln[3].n7 ctln[3] 7.38553
R31476 ctln[3] ctln[3].n7 2.82782
R31477 ctln[3].n6 ctln[3].n2 2.36635
R31478 ctln[3].n5 ctln[3].n4 0.923577
R31479 ctln[3].n7 ctln[3].n6 0.905693
R31480 ctlp[1].n4 ctlp[1].n1 292.5
R31481 ctlp[1].n3 ctlp[1].n2 92.5005
R31482 ctlp[1] ctlp[1].n3 81.3181
R31483 ctlp[1].n1 ctlp[1].t1 26.5955
R31484 ctlp[1].n0 ctlp[1].t0 25.8903
R31485 ctlp[1].n2 ctlp[1].t3 24.9236
R31486 ctlp[1].n2 ctlp[1].t2 24.9236
R31487 ctlp[1] ctlp[1].n4 15.5613
R31488 ctlp[1].n6 ctlp[1] 10.1205
R31489 ctlp[1].n5 ctlp[1].n0 9.48617
R31490 ctlp[1].n3 ctlp[1] 5.27109
R31491 ctlp[1].n5 ctlp[1] 2.60833
R31492 ctlp[1] ctlp[1].n5 1.85252
R31493 ctlp[1].n4 ctlp[1] 1.50638
R31494 ctlp[1].n1 ctlp[1].n0 0.248635
R31495 ctlp[1].n6 ctlp[1] 0.131056
R31496 ctlp[1] ctlp[1].n6 0.00798673
R31497 result[2].n2 result[2].n1 354.634
R31498 result[2].n6 result[2].n4 151.127
R31499 result[2].n6 result[2].n5 107.763
R31500 result[2].n2 result[2].n0 96.9298
R31501 result[2].n4 result[2].t6 40.0005
R31502 result[2].n4 result[2].t7 40.0005
R31503 result[2].n5 result[2].t4 40.0005
R31504 result[2].n5 result[2].t5 40.0005
R31505 result[2].n0 result[2].t0 27.5805
R31506 result[2].n0 result[2].t1 27.5805
R31507 result[2].n1 result[2].t2 27.5805
R31508 result[2].n1 result[2].t3 27.5805
R31509 result[2] result[2].n3 19.2609
R31510 result[2].n3 result[2].n2 15.309
R31511 result[2].n8 result[2] 8.05976
R31512 result[2].n7 result[2].n6 6.77697
R31513 result[2] result[2].n8 6.41086
R31514 result[2].n3 result[2] 2.70819
R31515 result[2].n7 result[2] 1.73877
R31516 result[2].n8 result[2].n7 0.948648
R31517 trim[2].n9 trim[2].n8 349.738
R31518 trim[2].n11 trim[2].n10 292.5
R31519 trim[2].n11 trim[2].n4 292.5
R31520 trim[2].n13 trim[2].n3 193.387
R31521 trim[2].n7 trim[2].n5 151.127
R31522 trim[2].n7 trim[2].n6 107.763
R31523 trim[2].n5 trim[2].t7 40.0005
R31524 trim[2].n5 trim[2].t4 40.0005
R31525 trim[2].n6 trim[2].t5 40.0005
R31526 trim[2].n6 trim[2].t6 40.0005
R31527 trim[2].n8 trim[2].t3 27.5805
R31528 trim[2].n8 trim[2].t0 27.5805
R31529 trim[2].n12 trim[2].t1 23.6405
R31530 trim[2].n3 trim[2].t2 23.1644
R31531 trim[2].n10 trim[2].n9 14.7697
R31532 trim[2].n4 trim[2].n2 11.243
R31533 trim[2] trim[2].n7 10.4115
R31534 trim[2].n13 trim[2].n1 9.3005
R31535 trim[2].n14 trim[2].n13 9.3005
R31536 trim[2].n13 trim[2].n12 9.3005
R31537 trim[2].n14 trim[2].n0 9.04377
R31538 trim[2].n1 trim[2].n0 9.01973
R31539 trim[2].n11 trim[2].n3 4.23401
R31540 trim[2].n15 trim[2].n2 4.13041
R31541 trim[2].n12 trim[2].n11 3.9405
R31542 trim[2].n13 trim[2].n2 3.09077
R31543 trim[2] trim[2].n16 2.48707
R31544 trim[2].n16 trim[2].n15 2.24426
R31545 trim[2].n9 trim[2].n4 1.96973
R31546 trim[2].n10 trim[2] 0.246654
R31547 trim[2].n15 trim[2].n1 0.03175
R31548 trim[2].n16 trim[2].n0 0.0141816
R31549 trim[2].n15 trim[2].n14 0.0101154
R31550 result[7].n6 result[7].n5 585
R31551 result[7].n2 result[7].n0 585
R31552 result[7] result[7].n6 297.269
R31553 result[7].n4 result[7].n3 92.5005
R31554 result[7].n5 result[7].n4 79.8123
R31555 result[7].n6 result[7].t0 26.5955
R31556 result[7].n3 result[7].t2 24.9236
R31557 result[7].n3 result[7].t3 24.9236
R31558 result[7].n6 result[7].n2 16.7455
R31559 result[7].n7 result[7] 12.2035
R31560 result[7].n2 result[7].t1 9.8505
R31561 result[7].n6 result[7].n1 9.13618
R31562 result[7].n4 result[7] 5.27109
R31563 result[7] result[7].n7 3.45106
R31564 result[7] result[7].n1 2.73954
R31565 result[7].n5 result[7] 1.50638
R31566 result[7].n7 result[7].n0 1.10628
R31567 result[7].n1 result[7].n0 0.0205962
R31568 result[5].n8 result[5].n7 185
R31569 result[5].n4 result[5].n3 143.643
R31570 result[5].n5 result[5] 81.5159
R31571 result[5].n3 result[5].t1 26.5955
R31572 result[5].n3 result[5].t0 26.5955
R31573 result[5].n6 result[5].t3 24.9236
R31574 result[5].n7 result[5].n6 15.6928
R31575 result[5].n8 result[5].n1 9.3005
R31576 result[5].n9 result[5].n8 9.3005
R31577 result[5].n7 result[5].t2 9.23127
R31578 result[5].n9 result[5].n0 9.05098
R31579 result[5] result[5].n4 9.02598
R31580 result[5].n1 result[5].n0 9.01252
R31581 result[5].n6 result[5].n5 8.25053
R31582 result[5].n4 result[5] 7.64268
R31583 result[5].n10 result[5].n2 3.79439
R31584 result[5] result[5].n11 3.05818
R31585 result[5].n11 result[5].n10 2.24426
R31586 result[5].n2 result[5] 2.08974
R31587 result[5].n8 result[5].n2 2.03855
R31588 result[5].n8 result[5].n5 0.214619
R31589 result[5].n10 result[5].n1 0.0389615
R31590 result[5].n11 result[5].n0 0.0141816
R31591 result[5].n10 result[5].n9 0.00290385
R31592 result[1].n6 result[1] 585.251
R31593 result[1].n8 result[1].n7 585
R31594 result[1].n6 result[1].n5 292.5
R31595 result[1] result[1].n4 95.7632
R31596 result[1].n5 result[1] 79.5613
R31597 result[1].n6 result[1].t0 26.5955
R31598 result[1].n4 result[1].t3 24.9236
R31599 result[1].n4 result[1].t2 24.9236
R31600 result[1].n7 result[1].n6 16.7455
R31601 result[1] result[1].n2 10.4588
R31602 result[1].n7 result[1].t1 9.8505
R31603 result[1].n8 result[1].n1 9.3005
R31604 result[1].n9 result[1].n8 9.3005
R31605 result[1].n6 result[1].n3 9.1516
R31606 result[1].n9 result[1].n0 9.05098
R31607 result[1].n1 result[1].n0 9.01252
R31608 result[1].n5 result[1] 7.02795
R31609 result[1] result[1].n3 4.01265
R31610 result[1].n10 result[1].n2 3.75172
R31611 result[1] result[1].n11 3.05818
R31612 result[1].n11 result[1].n10 2.24426
R31613 result[1].n8 result[1].n2 1.87152
R31614 result[1].n10 result[1].n1 0.0389615
R31615 result[1].n11 result[1].n0 0.0141816
R31616 result[1].n8 result[1].n3 0.00492585
R31617 result[1].n10 result[1].n9 0.00290385
R31618 trim[0].n2 trim[0].n0 585
R31619 trim[0].n11 trim[0].n4 349.738
R31620 trim[0].n10 trim[0].n3 292.5
R31621 trim[0].n12 trim[0].n3 292.5
R31622 trim[0].n7 trim[0].n5 151.127
R31623 trim[0].n7 trim[0].n6 107.763
R31624 trim[0].n5 trim[0].t7 40.0005
R31625 trim[0].n5 trim[0].t4 40.0005
R31626 trim[0].n6 trim[0].t5 40.0005
R31627 trim[0].n6 trim[0].t6 40.0005
R31628 trim[0].n4 trim[0].t3 27.5805
R31629 trim[0].n4 trim[0].t0 27.5805
R31630 trim[0].n1 trim[0].t1 23.7598
R31631 trim[0].n9 trim[0] 19.2609
R31632 trim[0].n2 trim[0].t2 14.7755
R31633 trim[0].n11 trim[0].n10 14.7697
R31634 trim[0].n3 trim[0].n2 12.8055
R31635 trim[0].n13 trim[0].n12 12.3259
R31636 trim[0] trim[0].n8 9.00791
R31637 trim[0].n1 trim[0].n0 8.9018
R31638 trim[0].n8 trim[0].n7 6.77697
R31639 trim[0].n10 trim[0].n9 5.90819
R31640 trim[0].n3 trim[0].n1 3.77188
R31641 trim[0].n9 trim[0] 2.70819
R31642 trim[0].n12 trim[0].n11 1.96973
R31643 trim[0] trim[0].n13 1.77665
R31644 trim[0].n8 trim[0] 1.73877
R31645 trim[0].n13 trim[0].n0 1.20582
R31646 net3.t0 net3.n5 440.25
R31647 net3.n0 net3.t2 323.342
R31648 net3.n1 net3.t3 309.017
R31649 net3.n1 net3.t5 231.897
R31650 net3.n0 net3.t4 194.809
R31651 net3.n6 net3.t0 135.105
R31652 net3.n4 net3.t1 123.654
R31653 net3.n2 net3.n1 92.3677
R31654 net3 net3.n4 82.2255
R31655 net3 net3.n0 78.9338
R31656 net3 net3.n3 29.2625
R31657 net3.n3 net3 23.4732
R31658 net3.n2 net3 17.8366
R31659 net3.n5 net3 10.9042
R31660 net3 net3.n6 6.41453
R31661 net3.n3 net3.n2 5.35533
R31662 net3.n5 net3 5.21532
R31663 net3.n4 net3 5.16973
R31664 net3.n6 net3 4.06431
R31665 comp.n7 comp.t0 222.725
R31666 comp.n5 comp.t1 177.171
R31667 comp.n5 comp.n4 152
R31668 comp.n6 comp.n3 152
R31669 comp.n6 comp.n5 10.5442
R31670 comp.n9 comp.n8 9.3005
R31671 comp.n8 comp.n1 9.3005
R31672 comp.n9 comp.n0 9.05098
R31673 comp.n1 comp.n0 9.01252
R31674 comp.n8 comp.n7 8.76429
R31675 comp.n4 comp 5.51161
R31676 comp.n10 comp.n2 4.02719
R31677 comp comp.n11 3.39779
R31678 comp.n4 comp.n3 2.48939
R31679 comp.n7 comp.n6 2.25988
R31680 comp.n11 comp.n10 2.24426
R31681 comp.n2 comp 1.64775
R31682 comp.n8 comp.n2 1.61183
R31683 comp.n8 comp.n3 0.533833
R31684 comp.n10 comp.n1 0.0389615
R31685 comp.n11 comp.n0 0.0141816
R31686 comp.n10 comp.n9 0.00290385
R31687 cal.n3 cal.t0 259.022
R31688 cal.n3 cal.t1 175.798
R31689 cal.n6 cal.n4 9.3005
R31690 cal.n7 cal.n6 9.3005
R31691 cal.n4 cal.n0 9.04669
R31692 cal.n8 cal.n7 9.04377
R31693 cal.n6 cal.n3 7.31035
R31694 cal.n5 cal.n2 3.98384
R31695 cal.n9 cal.n8 3.41895
R31696 cal.n5 cal 1.78438
R31697 cal.n6 cal.n5 1.74562
R31698 cal.n2 cal.n1 1.35824
R31699 cal.n9 cal.n0 0.867979
R31700 cal cal.n9 0.381556
R31701 cal.n8 cal.n1 0.0376622
R31702 cal.n4 cal.n2 0.03175
R31703 cal.n7 cal.n2 0.0101154
R31704 cal.n1 cal.n0 0.00974356
R31705 rstn.n3 rstn.t0 259.027
R31706 rstn.n3 rstn.t1 175.782
R31707 rstn.n5 rstn.n4 9.3005
R31708 rstn.n8 rstn.n7 9.3005
R31709 rstn.n4 rstn.n0 9.0697
R31710 rstn.n9 rstn.n8 9.02214
R31711 rstn.n5 rstn.n3 7.31533
R31712 rstn.n6 rstn.n2 4.57427
R31713 rstn.n10 rstn.n9 3.41895
R31714 rstn.n7 rstn.n6 2.24915
R31715 rstn.n2 rstn.n1 1.35818
R31716 rstn.n10 rstn.n0 0.868169
R31717 rstn.n6 rstn.n5 0.692392
R31718 rstn.n7 rstn 0.692392
R31719 rstn rstn.n10 0.0932894
R31720 rstn.n9 rstn.n1 0.0376622
R31721 rstn.n8 rstn.n2 0.03175
R31722 rstn.n1 rstn.n0 0.0103621
R31723 rstn.n4 rstn.n2 0.0101154
R31724 en.n2 en.t0 259.027
R31725 en.n2 en.t1 175.782
R31726 en.n3 en.n1 9.3005
R31727 en.n6 en.n5 9.3005
R31728 en.n1 en.n0 9.04136
R31729 en.n6 en.n0 9.02214
R31730 en.n3 en.n2 7.31533
R31731 en.n7 en.n4 4.57427
R31732 en en.n8 3.02215
R31733 en.n5 en.n4 2.24915
R31734 en.n8 en.n7 2.24426
R31735 en.n4 en.n3 0.692392
R31736 en.n5 en 0.692392
R31737 en.n7 en.n6 0.03175
R31738 en.n8 en.n0 0.0141816
R31739 en.n7 en.n1 0.0101154
C0 _013_ a_995_3530# 2.53e-20
C1 a_4512_11305# a_4655_10071# 4.4e-20
C2 a_561_6031# a_2313_6183# 1.18e-19
C3 net53 a_3868_10217# 4.72e-19
C4 a_10699_3311# a_11343_3317# 2.44e-19
C5 net44 _083_ 0.00381f
C6 net9 a_11987_8757# 0.0159f
C7 _048_ a_3847_4438# 3.1e-19
C8 _081_ _039_ 9.79e-21
C9 net15 _099_ 0.0134f
C10 a_9839_3615# VPWR 0.371f
C11 a_10699_3311# a_11149_3017# 1.18e-19
C12 _004_ a_1129_6273# 0.00175f
C13 a_14347_9480# _128_ 0.167f
C14 _063_ a_7088_7119# 9.17e-21
C15 _101_ a_3053_8207# 0.00183f
C16 _129_ _130_ 0.292f
C17 net46 _027_ 0.283f
C18 _024_ _058_ 0.047f
C19 _110_ a_10111_1679# 0.00158f
C20 _065_ a_8083_8181# 0.0512f
C21 _128_ a_13142_7271# 1.32e-20
C22 net40 a_13607_4943# 7.76e-19
C23 a_395_6031# a_1476_4777# 4.72e-21
C24 net13 a_4805_8207# 1.84e-20
C25 net43 _081_ 0.00795f
C26 a_1476_6031# a_395_4405# 4.72e-21
C27 a_8298_5487# a_10699_5487# 2.93e-20
C28 _059_ _093_ 9.99e-21
C29 net4 a_9459_7895# 0.0121f
C30 clknet_2_2__leaf_clk a_10543_2455# 5.1e-19
C31 a_9734_2223# VPWR 9.76e-19
C32 _078_ result[1] 4.11e-20
C33 cal_itt\[2\] a_9460_6807# 5.23e-21
C34 net15 a_3053_8457# 0.00523f
C35 a_1476_10217# a_1844_9129# 1.55e-20
C36 a_1651_10143# net24 3.61e-22
C37 mask\[7\] a_3133_11247# 9.47e-19
C38 _059_ a_5166_5193# 5.19e-20
C39 a_8745_4943# _107_ 3.06e-19
C40 a_10781_5487# VPWR 0.192f
C41 net12 a_5878_9295# 3.73e-19
C42 a_4993_6273# a_5502_6397# 2.6e-19
C43 a_4425_6031# a_4871_6031# 2.28e-19
C44 _040_ a_4349_8449# 0.0242f
C45 net19 _119_ 0.442f
C46 clknet_2_0__leaf_clk a_561_4405# 0.0103f
C47 trim_mask\[4\] a_7223_2465# 2.7e-19
C48 _036_ cal_count\[1\] 2.79e-20
C49 _066_ trim_mask\[1\] 1.32e-21
C50 a_4443_9295# a_5423_9011# 0.0117f
C51 net14 a_395_2767# 0.00162f
C52 net12 _054_ 2.18e-21
C53 _042_ a_561_9845# 2.53e-20
C54 _007_ _006_ 0.00117f
C55 net26 _008_ 0.317f
C56 _136_ a_10138_5807# 1.49e-19
C57 cal_itt\[0\] a_9957_7663# 0.114f
C58 net18 a_10005_6031# 1.49e-19
C59 net14 a_455_3571# 0.00326f
C60 _067_ a_11016_6691# 4.38e-19
C61 net47 clknet_2_3__leaf_clk 0.481f
C62 net44 a_3303_7119# 2.16e-20
C63 net44 a_8360_10383# 0.00175f
C64 mask\[4\] a_2953_9845# 2.97e-20
C65 net13 a_5067_2045# 0.00247f
C66 a_12231_6005# a_13111_6031# 2.14e-19
C67 net52 a_5423_9011# 6.74e-22
C68 a_15054_5193# _047_ 4.96e-19
C69 a_9207_3311# VPWR 0.144f
C70 _065_ a_11709_6273# 4.41e-19
C71 net46 a_12870_2589# 0.00339f
C72 clknet_2_1__leaf_clk a_4043_10143# 0.0101f
C73 _065_ mask\[0\] 6.95e-19
C74 _047_ trim_val\[1\] 0.00257f
C75 a_5691_7637# a_6835_7669# 5.84e-21
C76 net4 clk 0.0808f
C77 a_2815_9447# a_2857_7637# 1.56e-20
C78 _010_ net27 1.37e-19
C79 net4 en_co_clk 0.125f
C80 trim_mask\[4\] a_9099_3689# 0.0358f
C81 a_13393_1707# VPWR 5.67e-19
C82 _074_ result[3] 6.03e-19
C83 _019_ a_3615_8207# 1.79e-19
C84 a_15023_6031# clkc 7.28e-19
C85 net23 a_1476_7119# 0.00198f
C86 _002_ VPWR 0.414f
C87 a_4687_12319# mask\[6\] 1.6e-20
C88 mask\[1\] clknet_0_clk 1.17e-19
C89 net23 mask\[0\] 0.241f
C90 net13 a_5363_591# 0.241f
C91 cal_itt\[2\] _107_ 5.64e-19
C92 a_8307_4943# a_8473_5193# 0.144f
C93 clknet_2_3__leaf_clk a_8820_6005# 0.00128f
C94 net4 a_9084_4515# 0.00574f
C95 _032_ a_10016_1679# 0.16f
C96 a_9595_1679# a_10219_2045# 9.73e-19
C97 _050_ VPWR 1.82f
C98 calibrate net41 0.0278f
C99 _030_ a_13625_3317# 0.329f
C100 a_13459_3317# a_14193_3285# 0.0701f
C101 _037_ a_11622_7485# 2.13e-19
C102 net24 result[2] 0.0288f
C103 _036_ a_12612_8725# 2.56e-19
C104 a_11987_8757# a_12436_9129# 0.198f
C105 net46 a_11955_3689# 0.00181f
C106 a_10055_5487# trim_mask\[4\] 1.81e-20
C107 net15 a_4259_6031# 2.65e-20
C108 net22 _121_ 7.52e-21
C109 mask\[6\] net13 0.015f
C110 a_2787_9845# a_3303_10217# 0.106f
C111 _018_ a_3521_9813# 1.1e-20
C112 _051_ net42 0.00681f
C113 _051_ a_4901_2773# 3.97e-19
C114 a_7916_8041# a_8078_7663# 0.00645f
C115 net46 _117_ 5.03e-19
C116 clknet_2_1__leaf_clk a_2787_7119# 0.00309f
C117 _066_ a_10781_5807# 3.82e-20
C118 _052_ VPWR 0.357f
C119 net37 a_15299_6575# 6.9e-20
C120 a_1099_12533# result[7] 0.0905f
C121 a_5055_1679# VPWR 0.001f
C122 net3 _013_ 1.05e-19
C123 clknet_2_2__leaf_clk a_13607_1513# 7.44e-19
C124 a_8307_6575# a_8389_5193# 8.03e-21
C125 clknet_0_clk _015_ 2e-20
C126 a_561_6031# VPWR 0.581f
C127 _029_ _058_ 0.00671f
C128 _098_ VPWR 0.184f
C129 a_10593_9295# a_10774_9661# 8.75e-19
C130 trim_mask\[4\] a_10018_3677# 0.00226f
C131 a_1867_3317# a_2479_3689# 3.82e-19
C132 _110_ a_13519_4007# 0.132f
C133 a_2033_3317# a_2288_3677# 0.0642f
C134 _077_ a_6056_8359# 0.105f
C135 a_9602_6614# VPWR 1.7e-19
C136 _076_ _072_ 0.00276f
C137 cal_itt\[1\] a_10383_7093# 0.0627f
C138 cal_itt\[2\] a_8495_6895# 0.12f
C139 a_3615_8207# VPWR 0.429f
C140 mask\[0\] a_2225_7663# 0.00641f
C141 state\[2\] a_4815_3031# 0.0739f
C142 a_2953_9845# a_2815_9447# 1.24e-19
C143 net54 state\[1\] 0.201f
C144 net52 a_2489_7983# 0.00236f
C145 net49 a_13975_3689# 0.00704f
C146 _016_ a_1476_7119# 6.48e-19
C147 _088_ trim_mask\[4\] 1.03e-19
C148 net31 a_13459_3317# 1.1e-20
C149 net43 result[5] 7.57e-19
C150 a_8455_10383# _041_ 7.81e-21
C151 cal_count\[0\] trimb[4] 5.67e-20
C152 mask\[0\] _016_ 0.0328f
C153 _026_ a_12625_2601# 7.86e-21
C154 a_12056_6031# a_13349_6031# 8.66e-20
C155 _104_ a_7184_2339# 1.36e-22
C156 net51 a_6419_8207# 4.69e-19
C157 state\[0\] a_4815_3031# 0.216f
C158 _108_ a_14702_3311# 2.09e-19
C159 clknet_2_3__leaf_clk net5 7.24e-20
C160 clknet_2_1__leaf_clk a_3208_10205# 1.61e-19
C161 net15 a_4043_7093# 8.76e-19
C162 clknet_2_1__leaf_clk a_2689_8751# 2.91e-20
C163 _128_ a_13562_8751# 0.00794f
C164 net14 a_1129_4373# 0.0127f
C165 a_14931_591# ctln[2] 0.00504f
C166 a_4443_9295# a_4871_8181# 0.00137f
C167 mask\[0\] a_1019_6397# 1.44e-20
C168 _062_ _105_ 2.74e-19
C169 net50 a_10219_2045# 0.0012f
C170 a_4512_12393# _046_ 6.99e-20
C171 a_10872_1455# VPWR 1.33e-19
C172 a_14422_7093# a_14788_7369# 0.00519f
C173 _092_ a_3461_5193# 0.00685f
C174 _075_ a_5625_4943# 0.00123f
C175 _060_ a_4576_3427# 0.132f
C176 trim_val\[4\] trim_mask\[4\] 0.336f
C177 a_8583_3317# a_8298_2767# 0.0189f
C178 _065_ net54 0.0165f
C179 a_13783_6183# _061_ 5.51e-19
C180 _135_ a_14564_6397# 4.37e-19
C181 net4 ctln[0] 0.0219f
C182 net9 cal_count\[3\] 0.129f
C183 a_15259_7637# a_14377_7983# 7.66e-20
C184 a_6375_12021# a_7456_12393# 0.102f
C185 _101_ a_6743_10933# 2.95e-20
C186 net52 a_4871_8181# 2.4e-19
C187 a_10207_1679# trim_val\[3\] 2.33e-20
C188 net52 _076_ 0.0165f
C189 a_8154_11721# VPWR 0.00224f
C190 _112_ trim_mask\[2\] 6.44e-20
C191 a_4993_6273# a_5340_6031# 0.0512f
C192 _053_ _038_ 0.0563f
C193 _082_ a_1677_9545# 0.1f
C194 _123_ a_13279_8207# 0.025f
C195 net15 a_1660_12393# 1.64e-20
C196 a_11343_3317# a_11955_3689# 0.00188f
C197 _025_ a_11764_3677# 0.158f
C198 _104_ a_9839_3615# 0.0587f
C199 net4 _059_ 3.63e-20
C200 net9 a_12586_3311# 1.5e-19
C201 net54 a_5054_4399# 0.003f
C202 net45 a_5363_7369# 6.53e-19
C203 _028_ a_6906_2355# 0.00379f
C204 a_11764_3677# _026_ 2.79e-19
C205 mask\[4\] mask\[3\] 0.0432f
C206 a_9125_4943# VPWR 1.32e-19
C207 a_929_8757# a_1497_8725# 0.181f
C208 net55 _107_ 0.116f
C209 _132_ a_14788_7369# 0.0139f
C210 net19 a_9225_2197# 0.00452f
C211 a_6633_9845# a_7201_9813# 0.181f
C212 a_1137_5487# calibrate 2.18e-19
C213 _042_ a_11803_10383# 0.222f
C214 a_8820_12533# ctlp[5] 0.168f
C215 _014_ a_2479_3689# 8.45e-19
C216 a_11233_4405# a_10699_3311# 2.21e-20
C217 _073_ _062_ 5.27e-20
C218 a_13783_6183# a_13257_4943# 9.75e-21
C219 net33 a_14788_7369# 0.00445f
C220 clknet_2_0__leaf_clk result[0] 0.152f
C221 net12 a_6181_10383# 8.77e-19
C222 _101_ net45 0.349f
C223 _092_ a_12231_6005# 1.81e-21
C224 _120_ net30 1.38e-19
C225 cal_itt\[0\] a_10903_7261# 2.9e-21
C226 net23 a_448_6549# 3.74e-20
C227 _023_ a_1660_11305# 1.26e-19
C228 a_579_10933# net52 3.61e-19
C229 a_8381_9295# _041_ 1.89e-19
C230 a_7019_4407# a_7527_4631# 0.011f
C231 net19 a_8215_9295# 0.015f
C232 a_1019_6397# _079_ 4.5e-20
C233 _049_ net55 0.0429f
C234 clk ctln[1] 0.00132f
C235 _024_ a_11488_4765# 0.168f
C236 state\[2\] a_5087_3855# 9.29e-19
C237 a_9084_4515# a_9166_4515# 0.00477f
C238 a_11067_4405# a_11679_4777# 0.00188f
C239 _107_ a_7715_3285# 0.0022f
C240 a_7689_2589# clk 0.00121f
C241 _029_ a_13607_4943# 5.32e-19
C242 _104_ a_9207_3311# 5.97e-19
C243 _100_ a_4815_3031# 3.01e-21
C244 _084_ a_5997_10927# 1.14e-19
C245 trim_mask\[0\] a_13512_4943# 5.1e-19
C246 state\[2\] a_4443_1679# 6.3e-19
C247 a_4471_4007# state\[1\] 3.97e-19
C248 _127_ a_14467_8751# 2.03e-20
C249 _040_ net2 1.61e-21
C250 a_10747_8970# VPWR 0.209f
C251 a_448_7637# result[3] 0.00101f
C252 cal_count\[3\] a_10188_4105# 1.25e-21
C253 state\[0\] a_4443_1679# 0.00104f
C254 a_14564_6397# a_14649_6031# 0.00539f
C255 _061_ a_14181_6031# 2.39e-19
C256 a_11753_6031# _136_ 4.9e-19
C257 clknet_2_3__leaf_clk _068_ 1.16e-19
C258 _064_ a_10270_4105# 4.36e-20
C259 _069_ _071_ 4.41e-20
C260 _013_ valid 6.4e-21
C261 a_1129_9813# a_911_10217# 0.21f
C262 net16 a_14552_9071# 2.61e-19
C263 _041_ clknet_0_clk 2.41e-20
C264 _050_ _104_ 0.0258f
C265 _049_ a_7715_3285# 0.00139f
C266 a_7456_12393# a_7824_11305# 4.89e-20
C267 net44 _000_ 0.024f
C268 _065_ a_4471_4007# 1.46e-19
C269 _101_ a_3868_10217# 0.0581f
C270 clknet_0_clk a_7184_2339# 0.00248f
C271 _071_ a_8022_7119# 0.0217f
C272 a_4498_4373# a_4576_3427# 1.12e-19
C273 _122_ a_13111_6031# 3.83e-19
C274 a_5177_9537# a_5055_9295# 3.16e-19
C275 net16 clknet_2_2__leaf_clk 1.2e-19
C276 a_13091_4943# a_13519_4007# 7.88e-19
C277 clknet_2_1__leaf_clk _011_ 0.185f
C278 a_13459_3317# a_14083_3311# 9.73e-19
C279 net27 a_8154_11721# 3.75e-19
C280 net47 a_8827_9295# 9.59e-19
C281 mask\[3\] a_2815_9447# 0.197f
C282 _094_ _092_ 0.105f
C283 a_4259_6031# a_5449_6031# 2.56e-19
C284 a_9007_2601# clk 1.65e-19
C285 net45 a_6703_2197# 0.338f
C286 _125_ net2 0.0333f
C287 cal_count\[0\] _130_ 7.12e-22
C288 _058_ trim_mask\[1\] 0.00544f
C289 a_8301_8207# cal_itt\[3\] 1.98e-21
C290 a_2877_2197# net7 4.61e-20
C291 _052_ _104_ 0.434f
C292 a_5423_9011# _065_ 0.246f
C293 a_3303_7119# a_3565_7119# 0.00171f
C294 _015_ net41 0.00932f
C295 a_3868_7119# a_4030_7485# 0.00645f
C296 _110_ a_9839_3615# 0.00565f
C297 _074_ a_3947_12393# 2.34e-20
C298 a_2953_7119# a_5363_7369# 3.22e-20
C299 clknet_2_3__leaf_clk net46 0.375f
C300 net22 a_816_6031# 1.88e-19
C301 a_6375_12021# a_6743_10933# 1.9e-20
C302 a_13825_6031# a_13825_5185# 8.57e-20
C303 trim_mask\[0\] _103_ 0.232f
C304 _048_ _106_ 0.275f
C305 a_13919_8751# trimb[4] 4.07e-21
C306 a_1660_12393# a_1822_12015# 0.00645f
C307 _050_ a_7200_3631# 8.98e-19
C308 net52 a_395_9845# 5.43e-22
C309 _098_ _104_ 8.66e-21
C310 net19 a_8298_5487# 0.018f
C311 net24 _040_ 1.22e-19
C312 mask\[7\] a_1476_10217# 1.79e-19
C313 _093_ _107_ 1.73e-19
C314 _110_ a_9734_2223# 1.46e-19
C315 net26 a_8949_9537# 0.00133f
C316 clknet_2_2__leaf_clk a_10699_3311# 0.0282f
C317 _074_ a_3425_11721# 1.18e-19
C318 _062_ cal_count\[3\] 0.0484f
C319 _101_ a_2953_7119# 0.00234f
C320 net14 a_1660_12393# 0.00242f
C321 net45 _060_ 1.14e-19
C322 a_11369_7119# VPWR 3.32e-19
C323 _090_ a_6197_4399# 3.4e-19
C324 a_11116_8983# a_11258_9117# 0.00783f
C325 net49 trim_val\[1\] 0.115f
C326 _052_ a_7200_3631# 0.00403f
C327 a_14715_3615# a_15023_1679# 1.3e-19
C328 net43 a_3781_8207# 0.00113f
C329 mask\[3\] _081_ 2.32e-20
C330 trim_val\[2\] a_14471_591# 1.29e-20
C331 _100_ a_5087_3855# 0.0701f
C332 a_14972_5193# trim_val\[0\] 0.215f
C333 a_3597_12021# a_5496_12131# 5.89e-21
C334 net8 a_14931_591# 0.00169f
C335 a_8389_5193# VPWR 0.16f
C336 _122_ a_11622_7485# 0.0014f
C337 _037_ a_14422_7093# 5.48e-21
C338 a_4687_11231# mask\[4\] 3.75e-20
C339 net18 a_10864_7387# 0.0092f
C340 net31 a_15023_1135# 1.78e-19
C341 _049_ _093_ 0.0979f
C342 _048_ a_3667_3829# 0.315f
C343 a_10864_7387# a_10820_7485# 1.46e-19
C344 net44 mask\[4\] 0.42f
C345 a_3388_4631# _093_ 4.41e-19
C346 _099_ a_5363_4719# 0.0373f
C347 _065_ a_9677_8457# 0.00221f
C348 a_4227_8207# VPWR 8.7e-19
C349 cal_itt\[1\] a_8298_5487# 0.0102f
C350 trim_mask\[0\] a_11845_4765# 3.21e-21
C351 a_1651_7093# net22 8.92e-21
C352 _074_ _008_ 0.0504f
C353 net31 _125_ 0.00536f
C354 _048_ _033_ 3.33e-21
C355 _089_ _054_ 6.64e-21
C356 a_10699_5487# a_10781_5487# 0.171f
C357 net15 _097_ 0.211f
C358 a_10781_5807# _058_ 6.13e-20
C359 net4 a_9802_4007# 5.29e-20
C360 _123_ _069_ 5.86e-20
C361 a_579_10933# a_1679_10633# 9.57e-19
C362 net16 ctln[2] 1.33e-20
C363 net31 trimb[0] 0.00722f
C364 _029_ _113_ 5.19e-19
C365 net4 a_3399_2527# 0.0129f
C366 net43 a_1579_11471# 1.59e-19
C367 net40 a_13783_6183# 0.00154f
C368 net44 a_7447_8041# 7.55e-19
C369 net47 a_12664_8029# 0.00187f
C370 net4 _108_ 0.0253f
C371 _078_ a_1660_11305# 0.00364f
C372 _078_ a_1476_7119# 0.0125f
C373 a_3411_9839# mask\[2\] 1.94e-19
C374 cal_itt\[0\] a_9889_6873# 0.265f
C375 net23 a_1125_7663# 0.00889f
C376 clknet_0_clk _050_ 0.783f
C377 trim_val\[2\] a_13825_1109# 0.00131f
C378 _078_ mask\[0\] 0.177f
C379 a_4043_7093# a_4222_7119# 0.0074f
C380 net20 net44 0.0362f
C381 a_6007_7119# a_7088_7119# 0.102f
C382 _003_ a_7263_7093# 1.29e-20
C383 a_3868_7119# a_3977_7119# 0.00742f
C384 _133_ a_13356_7369# 0.00556f
C385 net53 a_2787_9845# 2.51e-22
C386 net8 a_13607_1513# 0.00525f
C387 a_13233_4737# VPWR 3.29e-19
C388 result[2] result[1] 0.0367f
C389 net23 a_2489_7983# 0.00101f
C390 _021_ a_7999_11231# 6.94e-21
C391 a_4687_12319# ctlp[7] 0.00107f
C392 net19 a_7902_10205# 5.5e-20
C393 a_6743_10933# a_7824_11305# 0.102f
C394 _074_ a_5524_9295# 6.87e-19
C395 a_7891_3617# VPWR 0.235f
C396 _034_ _049_ 0.0137f
C397 en_co_clk _064_ 3.22e-20
C398 net46 a_14715_3615# 0.277f
C399 a_7939_10383# a_7548_10217# 5.58e-19
C400 a_8105_10383# a_7723_10143# 1.72e-19
C401 a_745_10933# a_1822_10927# 1.46e-19
C402 a_9459_7895# _053_ 3.78e-20
C403 net18 a_7939_10383# 6.31e-21
C404 a_2019_9055# VPWR 0.392f
C405 net4 a_10655_2932# 3.38e-19
C406 _065_ a_4871_8181# 0.00212f
C407 a_561_4405# a_1585_4777# 2.36e-20
C408 a_395_2767# VPWR 0.283f
C409 clknet_0_clk _052_ 1.9e-20
C410 _065_ _076_ 0.669f
C411 clknet_2_2__leaf_clk _027_ 0.0294f
C412 a_455_3571# VPWR 0.437f
C413 _012_ a_1476_4777# 1.26e-19
C414 net55 trim_mask\[4\] 6.4e-20
C415 _108_ a_14172_4943# 8.3e-20
C416 mask\[7\] a_1357_11293# 9e-20
C417 net4 a_9460_6807# 0.0136f
C418 clknet_0_clk _098_ 4.99e-20
C419 a_9595_5193# _107_ 9.44e-19
C420 trim_val\[2\] a_13307_1707# 6.49e-19
C421 net45 a_4864_1679# 2.45e-19
C422 a_14347_9480# net40 2.3e-20
C423 mask\[6\] a_5915_10927# 0.121f
C424 a_7088_7119# _092_ 1.92e-19
C425 a_13881_1653# net8 0.00281f
C426 a_3615_8207# clknet_0_clk 3.01e-19
C427 a_3781_8207# a_2857_7637# 0.00198f
C428 a_12153_8757# a_12341_8751# 0.149f
C429 net26 a_3303_10217# 6.88e-20
C430 net53 a_7657_10217# 5.17e-20
C431 _074_ sample 0.0136f
C432 net5 _047_ 4.5e-19
C433 net44 a_7091_9839# 0.0134f
C434 a_4259_6031# a_5363_4719# 1.6e-20
C435 state\[2\] a_6822_4105# 1.95e-19
C436 _040_ a_4677_7882# 0.193f
C437 _063_ _092_ 0.367f
C438 a_1660_11305# a_3597_10933# 1.29e-20
C439 _078_ _079_ 0.0139f
C440 _094_ a_5547_5603# 3.47e-19
C441 _053_ clk 0.00574f
C442 _048_ _054_ 1.46e-19
C443 a_12520_7637# a_12249_7663# 7.79e-20
C444 a_12061_7669# a_12454_8041# 0.00206f
C445 _016_ a_1125_7663# 5.52e-20
C446 a_7939_10383# a_9129_10383# 2.56e-19
C447 _110_ a_10872_1455# 7.91e-21
C448 clknet_2_1__leaf_clk a_2368_9955# 0.0653f
C449 net43 a_561_9845# 0.0404f
C450 net47 a_9182_10749# 1.7e-19
C451 a_8673_10625# a_8551_10383# 3.16e-19
C452 _053_ en_co_clk 0.014f
C453 a_10005_6031# VPWR 0.582f
C454 a_855_4105# a_1201_3855# 0.0134f
C455 net50 net10 0.0105f
C456 net4 a_9004_3677# 2.01e-20
C457 a_8731_9295# _035_ 2.78e-21
C458 a_9471_9269# a_10239_9295# 7.36e-19
C459 a_763_8757# a_455_8181# 8.25e-19
C460 a_929_8757# a_1129_7361# 2.21e-21
C461 a_13142_8359# net2 0.0528f
C462 _005_ a_845_7663# 0.0125f
C463 trim_mask\[4\] a_7715_3285# 0.0619f
C464 clknet_2_2__leaf_clk a_12870_2589# 4.85e-19
C465 a_2489_7983# _016_ 1.97e-19
C466 net30 _051_ 0.705f
C467 _038_ a_11425_5487# 0.00313f
C468 net18 _111_ 7.79e-21
C469 _060_ a_4905_3855# 0.00527f
C470 _119_ trim_mask\[3\] 0.0315f
C471 net31 trim[1] 0.0412f
C472 _049_ a_3830_6281# 2.91e-19
C473 net30 _014_ 1.8e-20
C474 a_8307_4943# _103_ 2.31e-19
C475 net34 a_14788_7369# 3.27e-20
C476 net4 _107_ 0.0857f
C477 _122_ a_12992_8751# 0.00357f
C478 net32 a_14649_3689# 7.32e-20
C479 a_7088_7119# cal_itt\[3\] 0.00238f
C480 _062_ _119_ 1.74e-19
C481 net8 a_14334_1135# 1.46e-19
C482 net6 net7 0.00138f
C483 _087_ VPWR 0.506f
C484 a_5363_12559# _045_ 0.0124f
C485 _041_ a_6523_7119# 1.18e-21
C486 a_12424_3689# a_13183_3311# 4.38e-19
C487 a_12599_3615# a_13459_3317# 8.44e-21
C488 a_11859_3689# _030_ 2.04e-20
C489 a_8839_9661# VPWR 0.143f
C490 _042_ a_3977_10217# 1.61e-19
C491 net18 a_12631_591# 5.56e-21
C492 a_561_6031# a_2476_6281# 5.99e-20
C493 _092_ _096_ 0.276f
C494 a_8827_9295# _068_ 2.23e-19
C495 a_6519_3829# VPWR 0.256f
C496 _063_ cal_itt\[3\] 0.0056f
C497 mask\[4\] a_4801_9839# 0.0105f
C498 net47 a_13184_9117# 4.9e-19
C499 net14 _097_ 1.49e-20
C500 a_5340_6031# net3 6.9e-20
C501 net15 a_3748_6281# 0.00169f
C502 clknet_2_2__leaf_clk a_11955_3689# 5.75e-19
C503 net46 a_14099_1929# 0.00102f
C504 _108_ a_14099_3017# 9.71e-20
C505 _095_ a_4863_4917# 0.111f
C506 _099_ VPWR 0.234f
C507 net4 _049_ 2.26e-19
C508 _129_ a_13356_7369# 2.17e-20
C509 clknet_2_2__leaf_clk _117_ 8.95e-22
C510 net44 a_6987_12393# 9.54e-19
C511 _037_ _136_ 0.00132f
C512 net4 a_3388_4631# 5.62e-20
C513 a_8389_5193# _104_ 4.63e-19
C514 a_6927_591# VPWR 0.487f
C515 _062_ _095_ 4.99e-20
C516 a_6906_2355# ctln[6] 3.54e-20
C517 a_1129_4373# VPWR 0.222f
C518 a_4871_8181# a_4696_8207# 0.234f
C519 a_4349_8449# _077_ 4.25e-20
C520 _074_ a_6891_12393# 3.22e-20
C521 cal_itt\[0\] a_11141_6031# 0.00165f
C522 a_9761_1679# a_10787_1135# 6.67e-20
C523 a_7210_5807# _103_ 2.68e-19
C524 clknet_2_3__leaf_clk _065_ 0.305f
C525 _076_ a_4696_8207# 0.00196f
C526 a_3303_7119# _049_ 8.73e-19
C527 _078_ a_6099_10633# 9.33e-19
C528 a_3339_2767# a_2309_2229# 1.34e-19
C529 a_3053_8457# VPWR 0.196f
C530 _111_ trim_val\[0\] 4.54e-20
C531 net21 _084_ 1.92e-20
C532 trim_mask\[1\] _113_ 0.0392f
C533 _130_ en_co_clk 3.39e-20
C534 _072_ a_6835_7669# 0.0117f
C535 a_8083_8181# a_7001_7669# 2.48e-19
C536 _112_ a_14193_3285# 4.82e-19
C537 mask\[4\] a_8992_9955# 0.195f
C538 state\[0\] a_1867_3317# 2.65e-19
C539 net16 a_14335_2442# 0.0176f
C540 net40 a_14870_7369# 4.26e-19
C541 a_12231_6005# _136_ 0.00872f
C542 a_6906_2355# a_7181_2589# 0.00742f
C543 _048_ a_5731_4943# 0.00242f
C544 net43 a_4393_8207# 7.98e-21
C545 _100_ a_6822_4105# 6.54e-20
C546 a_14649_3689# VPWR 3.36e-20
C547 net16 net8 0.103f
C548 _128_ _036_ 0.0109f
C549 net13 a_4655_10071# 0.0128f
C550 clknet_2_1__leaf_clk a_6485_8181# 0.00601f
C551 _050_ net41 1.45e-20
C552 _024_ a_10975_4105# 0.121f
C553 mask\[0\] _004_ 8.96e-20
C554 clknet_2_0__leaf_clk a_3521_7361# 0.0526f
C555 a_3933_2767# a_4815_3031# 7.46e-19
C556 a_12061_7669# a_12430_7663# 4.45e-20
C557 state\[1\] a_2564_2589# 7.84e-20
C558 _053_ _059_ 4.32e-20
C559 a_6763_5193# _107_ 0.00349f
C560 _092_ a_5455_4943# 0.0669f
C561 _136_ a_13697_4373# 8.24e-20
C562 _104_ a_7891_3617# 7.15e-20
C563 clknet_2_0__leaf_clk a_1129_7361# 6.24e-20
C564 net52 a_6835_7669# 5.39e-21
C565 net46 _047_ 6.63e-19
C566 _041_ a_14249_8725# 0.00233f
C567 a_13562_8751# net40 1.88e-20
C568 _052_ net41 0.00169f
C569 net18 a_10676_1679# 0.00662f
C570 clknet_2_3__leaf_clk a_11233_4405# 4.14e-19
C571 net19 _041_ 0.013f
C572 a_10877_7983# VPWR 7.03e-20
C573 a_5537_4943# VPWR 1.4e-19
C574 cal_itt\[2\] a_8761_7983# 2.46e-19
C575 net19 a_7184_2339# 0.00104f
C576 _122_ a_14422_7093# 1.63e-20
C577 net9 a_11292_1251# 2.97e-19
C578 _083_ _008_ 0.129f
C579 a_13257_4943# a_14281_4943# 2.36e-20
C580 net31 _112_ 1.19e-20
C581 _045_ ctlp[6] 6.87e-19
C582 mask\[4\] a_9374_10383# 0.00237f
C583 _051_ state\[2\] 0.601f
C584 net46 _116_ 3.1e-19
C585 clknet_2_1__leaf_clk a_6007_7119# 5.04e-20
C586 net43 a_1844_9129# 0.221f
C587 a_7263_7093# a_7262_5461# 5.38e-22
C588 a_8105_10383# _042_ 0.545f
C589 _049_ a_6763_5193# 0.012f
C590 a_4259_6031# VPWR 0.413f
C591 en_co_clk a_3891_4943# 0.0534f
C592 a_10688_9295# _053_ 9.6e-21
C593 _051_ state\[0\] 0.205f
C594 a_579_10933# _023_ 0.166f
C595 mask\[7\] a_3597_12021# 2.26e-19
C596 net43 _006_ 0.00128f
C597 _095_ a_3817_4697# 0.00165f
C598 a_7010_3311# _028_ 0.0854f
C599 _078_ a_5423_9011# 0.0386f
C600 _014_ state\[0\] 1.06e-20
C601 _122_ _132_ 7.95e-21
C602 a_11023_5108# _111_ 1.05e-21
C603 net37 _135_ 1.53e-20
C604 trim_mask\[3\] a_9225_2197# 8.58e-21
C605 a_8298_2767# a_9572_2601# 0.00167f
C606 a_10055_2767# a_9747_2527# 0.00774f
C607 _004_ _079_ 0.149f
C608 _107_ a_9166_4515# 1.6e-19
C609 _036_ a_11895_7669# 0.00113f
C610 a_11987_8757# _037_ 2.81e-20
C611 net33 _122_ 9.06e-21
C612 _083_ a_5524_9295# 0.00198f
C613 _063_ a_9003_3829# 2.43e-20
C614 _093_ a_3123_3615# 9.52e-20
C615 clknet_2_0__leaf_clk _095_ 0.0837f
C616 a_9572_2601# a_9681_2601# 0.00742f
C617 a_9007_2601# a_9115_2223# 0.0572f
C618 a_9747_2527# a_9926_2589# 0.0074f
C619 clknet_0_clk a_8389_5193# 0.00374f
C620 a_7548_10217# a_7710_9839# 0.00645f
C621 cal_count\[1\] trimb[4] 5.25e-20
C622 _066_ _058_ 0.00225f
C623 _074_ a_1173_4765# 6.43e-19
C624 a_14199_7369# comp 2.03e-19
C625 _108_ net48 0.00244f
C626 net40 a_10055_5487# 6.94e-19
C627 mask\[3\] a_3781_8207# 9.22e-21
C628 _088_ a_6737_3855# 0.0482f
C629 _001_ a_13279_7119# 2.78e-21
C630 a_8022_7119# a_8935_6895# 0.00389f
C631 net17 net47 1.8e-20
C632 a_13783_6183# a_13349_6031# 1.53e-19
C633 a_13111_6031# a_13825_6031# 1.53e-19
C634 clknet_2_3__leaf_clk _067_ 0.0407f
C635 net3 a_2309_2229# 8.87e-20
C636 a_4043_7093# VPWR 0.368f
C637 a_7456_12393# a_6743_10933# 7.23e-19
C638 cal_count\[2\] _130_ 0.15f
C639 a_8563_10749# VPWR 0.134f
C640 a_9020_10383# a_9296_9295# 1.46e-20
C641 a_8455_10383# a_8839_9661# 4.92e-20
C642 a_1476_10217# a_1677_9545# 0.00151f
C643 _101_ a_2787_9845# 0.457f
C644 _060_ a_6210_4989# 1.71e-19
C645 a_4863_4917# calibrate 1.35e-20
C646 clknet_2_1__leaf_clk result[4] 0.0505f
C647 _007_ a_1677_9545# 2.9e-19
C648 _104_ a_6519_3829# 0.0025f
C649 net9 _135_ 4.07e-19
C650 net19 a_9207_3311# 0.00269f
C651 a_8820_6005# a_9443_6059# 0.0212f
C652 net43 result[7] 9.52e-20
C653 a_7379_2197# clk 0.00889f
C654 net37 _127_ 0.00111f
C655 a_14972_5193# VPWR 0.167f
C656 net13 _095_ 0.00928f
C657 _062_ calibrate 3.45e-19
C658 a_1660_11305# a_1651_10143# 3.09e-21
C659 a_1835_11231# a_1476_10217# 3.98e-19
C660 a_11435_2229# a_11601_2229# 0.906f
C661 a_1184_9117# _081_ 2.48e-21
C662 _110_ a_13233_4737# 5.4e-19
C663 a_5363_591# ctln[6] 1.71e-19
C664 _096_ a_5536_4399# 5.63e-20
C665 net47 a_12061_7669# 0.203f
C666 _041_ _001_ 8.1e-20
C667 a_1660_12393# VPWR 0.325f
C668 net40 _131_ 0.0122f
C669 mask\[1\] a_4995_7119# 9.97e-21
C670 a_1203_10927# a_1461_10357# 6.67e-19
C671 net19 _002_ 1.69e-20
C672 _078_ a_1125_7663# 0.0661f
C673 _136_ a_13825_5185# 2.34e-20
C674 net3 a_5691_2741# 3.74e-21
C675 _064_ a_9802_4007# 1.42e-20
C676 a_1095_12393# a_1203_12015# 0.0572f
C677 net14 a_1095_11305# 0.00717f
C678 a_1835_12319# a_2014_12381# 0.0074f
C679 a_1660_12393# a_1769_12393# 0.00742f
C680 _051_ _100_ 0.00624f
C681 clknet_0_clk a_7891_3617# 0.00165f
C682 clknet_2_3__leaf_clk clknet_2_2__leaf_clk 1.6e-20
C683 _023_ a_395_9845# 6.27e-19
C684 a_448_6549# _004_ 0.00117f
C685 net22 a_395_6031# 0.175f
C686 mask\[0\] a_1830_7119# 4.24e-19
C687 a_3565_10205# VPWR 1.18e-19
C688 net4 trim_mask\[4\] 0.0156f
C689 a_12341_8751# VPWR 0.104f
C690 _057_ ctln[4] 1.27e-19
C691 net24 a_2143_7663# 0.00126f
C692 _064_ _108_ 0.06f
C693 net20 a_7618_12015# 4.33e-20
C694 a_5363_12559# _078_ 1.82e-19
C695 net40 trim_val\[4\] 1.61e-20
C696 cal_count\[0\] _124_ 0.0173f
C697 net45 a_4576_3427# 3.5e-20
C698 _101_ a_2092_8457# 0.00187f
C699 trim_mask\[0\] net42 3.74e-20
C700 net46 a_14334_5309# 7.94e-19
C701 net12 net54 3.08e-20
C702 trim_mask\[3\] a_11292_1251# 0.103f
C703 mask\[2\] a_4443_9295# 0.0965f
C704 _035_ _122_ 3.09e-20
C705 _123_ a_13142_7271# 0.094f
C706 _112_ a_14083_3311# 8.3e-19
C707 net53 net26 0.132f
C708 a_561_9845# a_1585_10217# 2.36e-20
C709 net19 _052_ 2.02e-21
C710 a_12516_2601# net48 2.35e-20
C711 _078_ a_4871_8181# 4.8e-19
C712 a_3461_5193# a_3365_4943# 0.00219f
C713 a_7393_5193# VPWR 0.0075f
C714 a_561_7119# a_1129_7361# 0.186f
C715 a_395_9845# a_816_10205# 0.0931f
C716 _078_ _076_ 0.0104f
C717 a_8381_9295# a_8839_9661# 0.0346f
C718 a_8731_9295# a_9296_9295# 7.99e-20
C719 _064_ a_10655_2932# 0.0176f
C720 _077_ net2 8.99e-20
C721 net51 a_5363_7369# 0.049f
C722 net52 mask\[2\] 0.407f
C723 _035_ _063_ 8.42e-20
C724 a_3388_4631# a_3057_4719# 7.48e-20
C725 a_5547_5603# a_5455_4943# 6.99e-19
C726 _072_ a_6428_7119# 1.94e-20
C727 _074_ a_3303_10217# 4.42e-20
C728 clknet_2_1__leaf_clk _009_ 0.113f
C729 a_5340_6031# net54 1.55e-20
C730 _062_ a_8298_5487# 0.159f
C731 a_9460_6807# _064_ 1.78e-19
C732 a_10864_7387# VPWR 0.597f
C733 a_12077_3285# VPWR 0.215f
C734 _101_ a_2198_9117# 4.66e-20
C735 _133_ a_14377_7983# 0.0439f
C736 a_14686_3017# VPWR 0.00191f
C737 _122_ _136_ 0.00727f
C738 net12 a_6099_10633# 0.00691f
C739 _101_ net51 0.426f
C740 trim_val\[0\] a_14981_4020# 6.71e-21
C741 cal_count\[2\] a_13821_7119# 5.18e-19
C742 mask\[3\] a_5686_9661# 3.65e-19
C743 a_10990_7485# a_11396_6031# 1.91e-20
C744 _053_ _108_ 0.00353f
C745 trim_mask\[3\] a_10111_1679# 4.03e-20
C746 _012_ _014_ 1.56e-20
C747 a_561_9845# mask\[3\] 1.41e-20
C748 a_5455_4943# a_5536_4399# 2.58e-19
C749 calibrate a_3817_4697# 5.7e-20
C750 mask\[6\] a_4209_11293# 0.00211f
C751 _078_ a_579_10933# 0.00987f
C752 cal_count\[1\] _130_ 0.00126f
C753 a_5363_7369# _003_ 9.28e-20
C754 net2 a_10975_6031# 1.15e-20
C755 _114_ a_13257_1141# 5.54e-20
C756 _022_ a_2787_9845# 7.92e-21
C757 a_13881_1653# trim[2] 2e-19
C758 a_9503_4399# VPWR 0.651f
C759 a_5915_10927# _021_ 0.119f
C760 net45 a_1638_4399# 1.7e-19
C761 a_14422_7093# comp 4.35e-19
C762 cal_itt\[1\] a_9602_6614# 9.79e-19
C763 clknet_2_1__leaf_clk a_448_10357# 0.0227f
C764 a_1651_4703# a_1476_4777# 0.234f
C765 net46 a_13183_3311# 0.0424f
C766 a_1129_4373# a_1007_4777# 3.16e-19
C767 _002_ _001_ 2.75e-20
C768 net19 a_8154_11721# 1.13e-19
C769 net13 a_4866_11293# 4.27e-19
C770 clknet_2_0__leaf_clk calibrate 0.0216f
C771 a_745_10933# a_1203_10927# 0.0346f
C772 _037_ cal_count\[3\] 4.07e-20
C773 net4 a_3123_3615# 0.00105f
C774 _074_ a_1173_7119# 6.63e-19
C775 net43 a_4425_6031# 3.14e-20
C776 a_6763_5193# trim_mask\[4\] 1.85e-21
C777 net44 a_3781_8207# 0.0241f
C778 net15 _090_ 7.61e-19
C779 _108_ trim[0] 9.39e-20
C780 _074_ a_455_8181# 0.0126f
C781 net22 net30 0.0562f
C782 clknet_0_clk _099_ 2.05e-20
C783 _101_ _003_ 5.74e-19
C784 _064_ _107_ 0.00119f
C785 net19 a_9125_4943# 1.68e-19
C786 a_9369_3855# VPWR 9.97e-19
C787 a_14236_8457# a_14377_7983# 2.98e-19
C788 a_7942_2223# VPWR 0.0844f
C789 _053_ a_9460_6807# 0.00262f
C790 _051_ _118_ 2.39e-21
C791 a_9195_10357# net4 5.5e-20
C792 _065_ a_6835_7669# 8.53e-20
C793 _133_ a_10903_7261# 0.00172f
C794 a_7939_10383# VPWR 0.484f
C795 _132_ comp 0.00448f
C796 _024_ trim_val\[4\] 1.29e-20
C797 a_15023_1135# a_14931_591# 4.2e-19
C798 net45 a_1830_4765# 0.00342f
C799 net46 a_11691_4399# 0.0133f
C800 a_11394_9509# _041_ 8.03e-20
C801 _042_ a_1677_9545# 4.09e-19
C802 a_12231_6005# cal_count\[3\] 0.108f
C803 _017_ a_2857_7637# 0.0101f
C804 net33 comp 3.24e-19
C805 trim_mask\[1\] a_10975_4105# 0.0717f
C806 _015_ a_3224_2601# 5.52e-19
C807 a_7259_11305# mask\[4\] 1.92e-20
C808 a_929_8757# mask\[1\] 9.34e-20
C809 _095_ a_4091_4943# 1.24e-19
C810 net13 calibrate 0.00629f
C811 _074_ a_1019_9839# 0.00464f
C812 net16 a_13459_3317# 0.0152f
C813 a_9919_6614# en_co_clk 0.00124f
C814 a_8455_10383# a_8563_10749# 0.0572f
C815 net9 a_13279_7119# 2.06e-20
C816 net12 a_5423_9011# 0.00291f
C817 net46 net49 0.0204f
C818 net46 a_9269_2589# 0.0019f
C819 _076_ a_5502_6397# 3.59e-20
C820 _020_ a_6181_10383# 6.05e-20
C821 cal_itt\[1\] a_9125_4943# 2.8e-20
C822 _108_ a_14335_4020# 0.196f
C823 a_5997_11247# VPWR 6.5e-19
C824 a_9747_2527# VPWR 0.384f
C825 net43 a_3868_7119# 0.219f
C826 _010_ a_4209_12381# 2.14e-19
C827 net1 _013_ 0.00186f
C828 _078_ a_395_9845# 0.00749f
C829 a_8745_6895# a_8298_5487# 1.07e-20
C830 _053_ _107_ 0.0484f
C831 a_11116_8983# _041_ 0.0591f
C832 _097_ VPWR 0.461f
C833 net2 a_6173_7119# 1.04e-20
C834 net18 trim_mask\[2\] 0.00588f
C835 _074_ ctlp[0] 0.00279f
C836 _002_ a_7916_8041# 0.0343f
C837 net16 _109_ 0.0017f
C838 _122_ a_11987_8757# 6.27e-21
C839 a_9369_4105# a_9662_3855# 5.08e-20
C840 _058_ a_14071_3689# 4.87e-19
C841 _065_ a_5515_6005# 5.5e-21
C842 a_6007_7119# cal_itt\[3\] 1.84e-19
C843 trim_mask\[4\] a_7689_2589# 2.12e-19
C844 a_11803_10383# cal_count\[0\] 2.04e-19
C845 a_1129_6273# a_1007_6031# 3.16e-19
C846 a_14347_1439# a_14172_1513# 0.234f
C847 _111_ VPWR 0.369f
C848 _129_ a_14377_7983# 0.0619f
C849 _041_ a_4995_7119# 4.69e-21
C850 _025_ a_12424_3689# 7.13e-20
C851 a_11343_3317# a_13183_3311# 1.35e-20
C852 trim_mask\[1\] a_13881_2741# 0.118f
C853 net26 a_6007_9839# 0.0486f
C854 _048_ net3 1.05f
C855 net9 _041_ 0.00973f
C856 a_929_8757# a_1387_8751# 0.0276f
C857 net41 a_455_3571# 0.223f
C858 net43 mask\[7\] 0.0343f
C859 clknet_2_1__leaf_clk mask\[6\] 0.125f
C860 a_14347_9480# a_14565_9295# 0.00723f
C861 net46 a_11601_2229# 0.0283f
C862 mask\[1\] a_6198_8534# 1.34e-19
C863 _053_ _049_ 0.402f
C864 a_2564_2589# a_2755_2601# 4.61e-19
C865 _095_ a_2948_3689# 9.99e-20
C866 net42 a_8307_4943# 0.0928f
C867 mask\[5\] a_8105_10383# 6.07e-19
C868 a_12631_591# VPWR 0.268f
C869 net43 a_3977_10217# 0.00134f
C870 net16 trim[2] 4.03e-19
C871 clknet_0_clk a_4259_6031# 0.0239f
C872 _063_ _105_ 0.127f
C873 _125_ trimb[1] 0.00521f
C874 a_8563_10749# a_8381_9295# 1.92e-21
C875 _103_ a_8307_4719# 0.0945f
C876 _119_ _028_ 2.08e-20
C877 net27 a_7939_10383# 4.72e-19
C878 cal_itt\[3\] _092_ 4.32e-20
C879 net44 a_5686_9661# 1.67e-20
C880 trimb[0] trimb[1] 0.0464f
C881 net18 a_11045_3631# 1.51e-19
C882 net2 a_15023_5487# 4.69e-19
C883 a_5535_8181# a_5691_7637# 0.0197f
C884 _093_ a_1201_3855# 0.00193f
C885 net18 a_9719_1473# 4.1e-19
C886 a_7088_7119# _073_ 1.09e-19
C887 mask\[5\] a_6261_11247# 2.82e-19
C888 a_1651_7093# a_1476_6031# 1.05e-20
C889 mask\[4\] _008_ 0.0966f
C890 net33 trim[3] 0.00119f
C891 _064_ a_10838_2045# 6.72e-20
C892 _076_ a_7001_7669# 6.5e-19
C893 mask\[0\] a_1651_6005# 0.00278f
C894 a_6835_7669# _067_ 1.18e-20
C895 _063_ _073_ 1.41e-19
C896 a_13257_1141# VPWR 0.601f
C897 _087_ net41 1.99e-19
C898 mask\[1\] clknet_2_0__leaf_clk 7.16e-19
C899 a_816_4765# valid 0.00102f
C900 a_995_3530# a_2033_3317# 1.11e-19
C901 a_2857_7637# a_3868_7119# 0.00376f
C902 clknet_0_clk a_4043_7093# 0.0256f
C903 a_14347_9480# a_14335_7895# 1.75e-19
C904 _074_ a_579_12021# 0.00141f
C905 a_6519_3829# net41 9.74e-20
C906 net12 _076_ 0.619f
C907 a_10329_1921# a_10373_1679# 3.69e-19
C908 a_10111_1679# a_10207_1679# 0.0138f
C909 _101_ a_763_8757# 5.47e-20
C910 a_9761_1679# trim_val\[3\] 8.29e-19
C911 _104_ a_9503_4399# 6.77e-21
C912 _123_ _131_ 2.67e-19
C913 a_14715_3615# a_14540_3689# 0.234f
C914 a_13975_3689# _055_ 1.88e-20
C915 mask\[4\] a_5524_9295# 1.63e-20
C916 mask\[2\] _065_ 1.79e-20
C917 a_13142_8725# a_13562_8751# 0.144f
C918 a_12436_9129# _041_ 0.043f
C919 cal_itt\[0\] net30 3.6e-20
C920 net45 a_2953_7119# 2.36e-19
C921 _015_ a_5524_1679# 1.26e-19
C922 _025_ a_11435_2229# 1.44e-20
C923 net18 a_9595_1679# 2.82e-20
C924 net20 _008_ 7.12e-22
C925 a_6703_2197# a_7223_2465# 0.0435f
C926 cal_itt\[1\] a_11369_7119# 1.4e-19
C927 a_2828_12131# net52 8.6e-20
C928 _026_ a_11435_2229# 0.174f
C929 a_4043_10143# a_4655_10071# 0.0186f
C930 _095_ a_3461_5193# 0.00915f
C931 _029_ a_14281_4943# 2.47e-21
C932 a_845_7663# VPWR 0.00725f
C933 mask\[2\] net23 2.03e-20
C934 _104_ a_9369_3855# 0.00142f
C935 net46 a_14172_1513# 0.237f
C936 net31 a_15023_5487# 0.00667f
C937 a_9471_9269# _069_ 4.45e-19
C938 _076_ a_5340_6031# 0.00105f
C939 a_1467_7923# a_1129_7361# 0.00118f
C940 a_455_8181# a_448_7637# 0.0217f
C941 a_10676_1679# VPWR 0.305f
C942 net13 mask\[1\] 0.0277f
C943 a_7939_10383# a_8455_10383# 0.115f
C944 a_4995_7119# _050_ 1.33e-21
C945 net18 a_11098_6691# 4.94e-19
C946 clknet_2_2__leaf_clk _116_ 2.26e-20
C947 _101_ net26 0.261f
C948 clknet_2_0__leaf_clk _015_ 0.0843f
C949 trim_mask\[1\] a_9099_3689# 5.37e-21
C950 a_10188_4105# a_9839_3615# 0.00107f
C951 a_9802_4007# a_9664_3689# 7.96e-19
C952 a_1493_11721# a_1095_11305# 2.12e-19
C953 a_13607_4943# _058_ 0.00456f
C954 net43 _121_ 0.0321f
C955 a_3748_6281# VPWR 0.157f
C956 a_10593_9295# a_10798_9295# 3.7e-19
C957 net35 a_14172_4943# 0.00429f
C958 state\[1\] a_2143_2229# 1.28e-19
C959 net14 a_1211_7983# 3.92e-19
C960 trim_val\[3\] a_10787_1135# 0.00937f
C961 net44 a_4393_8207# 0.0019f
C962 a_9296_9295# _063_ 1.29e-21
C963 a_8298_2767# a_8491_2229# 0.0293f
C964 _037_ a_10383_7093# 1.58e-20
C965 a_6056_8359# VPWR 0.117f
C966 _108_ a_9664_3689# 2.38e-19
C967 _051_ a_3933_2767# 0.311f
C968 net22 a_1585_6031# 1.27e-19
C969 _065_ a_6428_7119# 2.9e-20
C970 _097_ a_2383_3689# 3.7e-19
C971 _010_ a_3431_10933# 5.33e-19
C972 _028_ a_7617_2589# 6.71e-19
C973 a_8491_2229# a_9681_2601# 2.56e-19
C974 trim_val\[2\] a_15023_2223# 0.00947f
C975 _008_ a_7091_9839# 2.01e-20
C976 _064_ trim_mask\[4\] 0.254f
C977 _092_ a_6737_4719# 2.32e-20
C978 net54 _089_ 4.07e-20
C979 cal_itt\[2\] _071_ 0.447f
C980 net46 a_10016_1679# 0.0054f
C981 _074_ net53 0.0143f
C982 _104_ a_9747_2527# 0.00112f
C983 a_7569_7637# net30 1.72e-20
C984 _049_ a_3891_4943# 9.03e-19
C985 _092_ a_5547_5603# 5.28e-20
C986 _102_ a_763_8757# 4.1e-21
C987 net16 a_14655_4399# 7.97e-19
C988 net32 a_14981_4020# 5.19e-19
C989 a_4165_11989# a_4674_12015# 2.6e-19
C990 a_14422_7093# a_14199_7369# 0.00498f
C991 net13 _015_ 0.171f
C992 a_1045_9545# VPWR 0.00478f
C993 _122_ cal_count\[3\] 4.88e-19
C994 state\[1\] a_4815_3031# 0.0651f
C995 a_8749_3317# a_9099_3689# 0.224f
C996 a_448_10357# result[4] 0.158f
C997 _110_ a_12077_3285# 5.43e-20
C998 net16 _125_ 0.0151f
C999 trim_mask\[2\] a_10055_2767# 0.00289f
C1000 a_13111_6031# _136_ 0.0118f
C1001 _086_ net26 6.86e-21
C1002 net45 a_2857_5461# 9.16e-19
C1003 clknet_0_clk a_10864_7387# 5.02e-20
C1004 a_7710_9839# VPWR 4.91e-19
C1005 net18 net50 1.09f
C1006 a_1129_9813# _082_ 0.00213f
C1007 a_9020_10383# a_8215_9295# 4.49e-21
C1008 _106_ a_7800_4631# 3.64e-19
C1009 mask\[2\] _016_ 2.53e-20
C1010 _096_ a_3365_4943# 2.32e-19
C1011 a_1095_11305# VPWR 0.212f
C1012 trim_mask\[1\] a_10018_3677# 1.97e-21
C1013 trim_mask\[4\] a_10851_1653# 7.62e-19
C1014 _063_ cal_count\[3\] 0.168f
C1015 net16 trimb[0] 1.1e-19
C1016 a_4443_9295# a_4609_9295# 0.737f
C1017 _062_ a_9839_3615# 3.55e-19
C1018 a_11509_3317# a_11967_3311# 0.0276f
C1019 a_7939_10383# a_8381_9295# 9.08e-21
C1020 _092_ a_5536_4399# 0.00326f
C1021 _035_ a_11814_9295# 6.62e-21
C1022 _028_ a_9225_2197# 5.82e-23
C1023 _122_ a_14981_8235# 5.55e-20
C1024 _023_ a_911_10217# 7.13e-19
C1025 _132_ a_14199_7369# 8.29e-19
C1026 a_13470_7663# a_13279_7119# 3.17e-21
C1027 _102_ net26 0.408f
C1028 net22 a_911_6031# 0.015f
C1029 a_579_10933# a_1651_10143# 3.63e-19
C1030 net46 a_11396_6031# 2.46e-19
C1031 a_2953_9845# a_3977_10217# 2.36e-20
C1032 a_3521_9813# a_3565_10205# 3.69e-19
C1033 a_11709_6273# a_11599_6397# 0.0977f
C1034 _110_ a_9503_4399# 0.109f
C1035 _084_ a_7109_11989# 2.17e-20
C1036 _042_ a_3840_8867# 7.6e-19
C1037 net52 a_4609_9295# 5.82e-23
C1038 a_10864_7387# a_10699_5487# 3.45e-21
C1039 net30 trim_mask\[0\] 0.0433f
C1040 net3 a_2033_3317# 1.57e-20
C1041 a_2787_7119# a_3521_7361# 0.0535f
C1042 _053_ trim_mask\[4\] 0.0186f
C1043 mask\[2\] a_4696_8207# 5.22e-21
C1044 _069_ a_9693_8029# 6.92e-19
C1045 _076_ a_6197_6281# 0.0142f
C1046 net22 _012_ 9.79e-21
C1047 trim_val\[4\] trim_mask\[1\] 0.00357f
C1048 _110_ a_9369_3855# 1.61e-20
C1049 net19 a_8839_9661# 0.00477f
C1050 a_911_7119# a_1173_7119# 0.00171f
C1051 a_9099_3689# a_9361_3677# 0.00171f
C1052 a_9317_3285# a_9773_3689# 4.2e-19
C1053 _094_ _095_ 0.0016f
C1054 net34 comp 0.108f
C1055 a_8583_3317# clk 2.69e-21
C1056 trim_mask\[2\] a_12691_2527# 0.0687f
C1057 a_10688_9295# _124_ 0.00285f
C1058 a_14981_4020# VPWR 0.279f
C1059 mask\[1\] a_561_7119# 6.5e-20
C1060 a_7939_3855# a_7223_2465# 3.56e-21
C1061 a_2857_7637# _121_ 5.11e-19
C1062 trim_mask\[2\] _114_ 0.154f
C1063 a_911_10217# a_816_10205# 0.0498f
C1064 a_1129_9813# a_1007_10217# 3.16e-19
C1065 calibrate _028_ 1.24e-19
C1066 a_11233_4405# a_11691_4399# 0.0346f
C1067 _058_ a_11488_4765# 0.00438f
C1068 cal_itt\[1\] a_10005_6031# 3.16e-19
C1069 a_11622_7485# _136_ 4.81e-19
C1070 _049_ a_7379_2197# 1.15e-19
C1071 a_9084_4515# a_8583_3317# 5.87e-21
C1072 _107_ a_9664_3689# 0.00111f
C1073 _022_ net26 8.91e-20
C1074 a_13091_4943# a_14972_5193# 5.68e-21
C1075 net44 a_4680_6031# 2.85e-19
C1076 _060_ _088_ 5.91e-21
C1077 a_13257_4943# a_14172_4943# 0.117f
C1078 a_4674_12015# VPWR 7.57e-19
C1079 a_11435_2229# _031_ 8.51e-20
C1080 a_11601_2229# a_12059_2223# 0.0346f
C1081 a_11067_3017# trim_val\[3\] 1.39e-19
C1082 net45 a_3386_2223# 1.7e-19
C1083 _046_ a_4055_12015# 4.33e-19
C1084 _050_ a_4863_4917# 2.2e-19
C1085 _048_ net54 0.0101f
C1086 _000_ a_8949_9537# 3.71e-19
C1087 a_8215_9295# a_8731_9295# 0.111f
C1088 clknet_2_1__leaf_clk a_1497_8725# 9.01e-21
C1089 mask\[4\] a_9195_10357# 0.122f
C1090 state\[1\] a_5087_3855# 0.214f
C1091 _058_ _113_ 0.00723f
C1092 trim_val\[4\] a_8749_3317# 0.0128f
C1093 a_9003_3829# a_9317_3285# 1.09e-19
C1094 net43 _080_ 0.00453f
C1095 _136_ a_13825_6031# 0.0495f
C1096 net47 a_13356_8457# 4.05e-19
C1097 a_1651_4703# _014_ 6.06e-19
C1098 _041_ clknet_2_0__leaf_clk 4.53e-21
C1099 net2 a_7351_8041# 1.86e-19
C1100 _110_ a_9747_2527# 0.0103f
C1101 _062_ _050_ 0.504f
C1102 _090_ a_5363_4719# 1.29e-19
C1103 net20 a_6891_12393# 0.00959f
C1104 net44 a_5633_9295# 0.00148f
C1105 state\[1\] a_4443_1679# 4.72e-21
C1106 a_1387_8751# a_561_7119# 2.17e-21
C1107 a_4709_2773# VPWR 0.138f
C1108 net15 a_3667_3829# 0.00151f
C1109 net24 _005_ 0.00456f
C1110 cal_count\[0\] a_14377_7983# 2.37e-20
C1111 a_8298_2767# _032_ 1.45e-19
C1112 cal_count\[2\] a_13356_7369# 7.38e-20
C1113 _055_ trim_val\[1\] 0.125f
C1114 a_10055_2767# a_9595_1679# 7.43e-20
C1115 a_2953_7119# a_2857_5461# 5.02e-20
C1116 net27 a_1095_11305# 5.3e-20
C1117 _134_ trim_mask\[0\] 1.05e-19
C1118 net16 trim[1] 5.53e-20
C1119 a_4680_6031# en_co_clk 5.36e-19
C1120 a_395_9845# a_1651_10143# 0.0436f
C1121 _065_ a_12061_7669# 1.53e-20
C1122 _010_ a_4687_12319# 2.58e-19
C1123 mask\[1\] a_4239_8573# 0.0278f
C1124 _078_ a_5915_11721# 0.0637f
C1125 _111_ _110_ 0.00413f
C1126 net45 a_8657_2229# 5.82e-23
C1127 a_4308_4917# VPWR 0.329f
C1128 net48 _056_ 0.0137f
C1129 _062_ _052_ 2.54e-20
C1130 _104_ a_10676_1679# 7.7e-20
C1131 net15 net24 0.00618f
C1132 a_14099_1929# net8 6.57e-19
C1133 _108_ _057_ 2.53e-21
C1134 a_11059_7356# a_10975_6031# 8.14e-19
C1135 _039_ a_816_6031# 1.22e-19
C1136 a_10903_7261# _038_ 1.35e-20
C1137 _062_ _098_ 3.97e-19
C1138 net13 _041_ 0.0129f
C1139 net46 _025_ 0.00717f
C1140 a_579_10933# a_1191_11305# 0.00188f
C1141 _023_ a_1000_11293# 0.16f
C1142 _074_ a_6007_9839# 1.16e-20
C1143 _101_ a_2961_9295# 0.00199f
C1144 net46 _026_ 0.0054f
C1145 a_3388_4631# a_3530_4438# 0.00557f
C1146 a_9460_6807# a_9919_6614# 6.64e-19
C1147 _062_ a_9602_6614# 2.49e-20
C1148 a_455_5747# sample 0.338f
C1149 net44 _017_ 2.51e-19
C1150 clknet_2_2__leaf_clk a_13183_3311# 0.0696f
C1151 net40 a_9595_5193# 1.45e-19
C1152 mask\[7\] mask\[3\] 5.1e-19
C1153 clknet_2_1__leaf_clk ctlp[7] 1.53e-19
C1154 trim_mask\[0\] a_13975_3689# 1.73e-19
C1155 _078_ a_7201_9813# 1.33e-20
C1156 net34 trim[3] 0.0749f
C1157 mask\[4\] a_8949_9537# 5.88e-19
C1158 _092_ _136_ 0.222f
C1159 a_14282_7119# VPWR 3.78e-19
C1160 _111_ a_12148_4777# 0.00162f
C1161 trim_mask\[3\] a_10872_1455# 0.0101f
C1162 trim_mask\[0\] state\[2\] 0.00126f
C1163 _108_ a_10245_5193# 1.2e-19
C1164 a_11023_5108# net50 0.109f
C1165 a_15023_8751# net2 0.0013f
C1166 a_1276_565# rstn 4.51e-19
C1167 _052_ a_9195_3689# 4.96e-21
C1168 net18 net2 0.0112f
C1169 _088_ a_7939_3855# 5.46e-19
C1170 a_7800_4631# _054_ 7.34e-20
C1171 mask\[6\] _009_ 4.05e-19
C1172 _134_ a_13933_6281# 0.00106f
C1173 _048_ a_7019_4407# 0.0259f
C1174 _132_ a_14422_7093# 0.0119f
C1175 a_14335_7895# _131_ 3.37e-19
C1176 a_7824_11305# net26 1.04e-19
C1177 a_561_4405# cal 0.00305f
C1178 a_395_4405# en 1.21e-19
C1179 net16 a_13142_8359# 5.04e-19
C1180 clknet_2_2__leaf_clk a_11691_4399# 9.04e-19
C1181 _013_ a_2143_2229# 2.38e-19
C1182 a_395_9845# result[2] 7.53e-20
C1183 a_2033_3317# valid 8.33e-20
C1184 _048_ a_4471_4007# 1.73e-20
C1185 trim_mask\[0\] a_13915_4399# 0.0595f
C1186 net33 a_14422_7093# 1.21e-19
C1187 a_5547_5603# a_5536_4399# 4.86e-19
C1188 _050_ a_3817_4697# 0.00133f
C1189 net50 a_10055_2767# 1.66e-20
C1190 net43 a_1677_9545# 3.67e-19
C1191 clknet_2_1__leaf_clk _021_ 0.143f
C1192 _053_ a_7320_3631# 0.00107f
C1193 a_2288_3677# VPWR 0.0846f
C1194 a_15299_6575# comp 0.00409f
C1195 a_1476_7119# a_1549_6794# 1.9e-19
C1196 a_1651_7093# _039_ 0.0101f
C1197 _072_ _051_ 8.19e-19
C1198 _110_ a_13257_1141# 0.00154f
C1199 a_7310_2223# VPWR 0.232f
C1200 net47 a_12522_8751# 2.38e-19
C1201 clknet_2_2__leaf_clk a_9269_2589# 0.00252f
C1202 clknet_2_2__leaf_clk net49 3.7e-21
C1203 _067_ a_9443_6059# 8.66e-19
C1204 _078_ a_1585_7119# 3.07e-19
C1205 trim_val\[1\] trim_val\[2\] 0.0161f
C1206 net43 a_1835_11231# 0.278f
C1207 net43 a_1651_7093# 0.294f
C1208 net30 a_8307_4943# 0.00193f
C1209 _123_ _036_ 0.012f
C1210 net18 _033_ 1.37e-20
C1211 _015_ a_2948_3689# 3.41e-20
C1212 clknet_2_0__leaf_clk _050_ 0.115f
C1213 net7 clk 0.0053f
C1214 net33 _132_ 0.00629f
C1215 _070_ VPWR 0.673f
C1216 a_1497_8725# a_1953_9129# 4.2e-19
C1217 a_1279_9129# a_1541_9117# 0.00171f
C1218 net44 a_4425_6031# 0.0282f
C1219 _065_ _120_ 0.123f
C1220 net53 _083_ 0.0625f
C1221 a_11343_3317# _025_ 0.389f
C1222 a_6891_12393# a_6987_12393# 0.0138f
C1223 net31 a_15023_8751# 0.00659f
C1224 _006_ a_1184_9117# 0.158f
C1225 _011_ a_1095_12393# 0.00291f
C1226 trim_mask\[2\] VPWR 1.14f
C1227 a_579_12021# a_1835_12319# 0.0436f
C1228 a_11343_3317# _026_ 8.37e-20
C1229 net19 a_8563_10749# 0.00193f
C1230 a_395_6031# a_1476_6031# 0.102f
C1231 a_8636_9295# _071_ 6.22e-20
C1232 _063_ a_10383_7093# 0.00322f
C1233 a_11149_3017# _026_ 0.00169f
C1234 net30 a_8298_2767# 5.18e-19
C1235 _053_ a_11895_7669# 0.00282f
C1236 net16 _112_ 0.0667f
C1237 _110_ a_10676_1679# 1.75e-19
C1238 net46 _051_ 1.84e-21
C1239 net40 a_14172_4943# 7.08e-20
C1240 clknet_2_2__leaf_clk a_11601_2229# 0.00202f
C1241 _078_ mask\[2\] 0.208f
C1242 a_12213_2589# VPWR 1.87e-19
C1243 clknet_2_0__leaf_clk a_561_6031# 0.00805f
C1244 net25 net24 1.32e-20
C1245 a_7723_6807# net30 0.0435f
C1246 net13 _050_ 0.00894f
C1247 _090_ VPWR 1.24f
C1248 _074_ _101_ 0.969f
C1249 _065_ a_11396_6031# 0.00802f
C1250 a_4775_6031# a_4871_6031# 0.0138f
C1251 a_4993_6273# a_5037_6031# 3.69e-19
C1252 a_4425_6031# en_co_clk 0.0293f
C1253 _095_ _096_ 0.136f
C1254 clknet_2_0__leaf_clk a_3615_8207# 0.264f
C1255 trim_mask\[0\] _100_ 1.03e-20
C1256 _040_ a_4871_8181# 0.00258f
C1257 net14 net24 0.00633f
C1258 trim_mask\[4\] a_7379_2197# 3.65e-19
C1259 a_9871_10383# clknet_2_3__leaf_clk 6.4e-22
C1260 a_5177_9537# a_5423_9011# 0.00152f
C1261 a_10219_2045# _117_ 1.39e-19
C1262 net15 a_4677_7882# 0.109f
C1263 _126_ net2 0.0842f
C1264 _076_ _040_ 3.91e-20
C1265 a_3847_4438# VPWR 8.37e-19
C1266 _053_ a_11491_6031# 3.23e-19
C1267 _136_ a_11045_5807# 3.16e-19
C1268 _111_ a_13091_4943# 2.22e-19
C1269 trim_val\[0\] a_14000_4719# 3.13e-19
C1270 cal_itt\[0\] _118_ 0.0023f
C1271 net53 a_8360_10383# 1.6e-21
C1272 _075_ _100_ 1.35e-20
C1273 net44 a_3868_7119# 1.96e-19
C1274 _051_ a_5931_4105# 6.43e-21
C1275 net16 ctlp[3] 2.35e-19
C1276 a_6007_7119# _073_ 2.64e-20
C1277 _003_ a_6515_6794# 0.109f
C1278 _092_ _105_ 2.75e-20
C1279 net46 a_10752_565# 1.46e-20
C1280 net13 a_5055_1679# 0.00132f
C1281 a_2143_2229# a_2755_2601# 0.00188f
C1282 a_2309_2229# a_2564_2589# 0.0594f
C1283 a_12056_6031# a_13783_6183# 4.46e-20
C1284 cal_count\[3\] a_13111_6031# 0.0717f
C1285 a_12231_6005# _135_ 1.09e-19
C1286 net42 a_8307_4719# 5.16e-19
C1287 a_11045_3631# VPWR 5.17e-20
C1288 net46 _031_ 0.438f
C1289 net29 a_579_10933# 1.88e-19
C1290 a_7019_4407# a_7021_4105# 4.68e-19
C1291 _097_ net41 3.65e-19
C1292 clknet_2_1__leaf_clk a_4655_10071# 2.24e-20
C1293 a_6835_7669# a_7001_7669# 0.578f
C1294 _101_ a_1279_9129# 3.1e-20
C1295 net13 _098_ 2.72e-21
C1296 trim_mask\[4\] a_9664_3689# 0.0389f
C1297 a_6056_8359# a_6198_8207# 0.00783f
C1298 net31 trim_val\[0\] 1.55e-19
C1299 a_9719_1473# VPWR 0.237f
C1300 _019_ a_4349_8449# 1.17e-19
C1301 _092_ a_7010_3311# 1.12e-20
C1302 net24 a_395_7119# 8.97e-21
C1303 a_11016_6691# a_10975_6031# 3.15e-19
C1304 net13 a_3615_8207# 0.00721f
C1305 calibrate a_4617_3855# 1.78e-19
C1306 a_12153_8757# net2 4.56e-20
C1307 clknet_2_3__leaf_clk _091_ 0.0011f
C1308 net39 VPWR 0.307f
C1309 a_4866_12381# ctlp[7] 1.98e-20
C1310 _085_ _078_ 0.00491f
C1311 _074_ _086_ 0.0915f
C1312 trim_mask\[4\] a_10689_2223# 0.00151f
C1313 a_3597_10933# mask\[2\] 9.95e-20
C1314 _135_ a_13697_4373# 2.87e-21
C1315 a_13783_6183# _058_ 2.94e-19
C1316 mask\[0\] a_2143_7663# 0.0739f
C1317 _030_ a_13975_3689# 5.3e-19
C1318 a_13459_3317# a_14715_3615# 0.0436f
C1319 a_3868_7119# en_co_clk 3.26e-22
C1320 net12 a_6835_7669# 5.89e-19
C1321 _036_ a_13142_8725# 9.37e-20
C1322 mask\[1\] a_1467_7923# 0.0536f
C1323 a_11987_8757# a_12992_8751# 0.178f
C1324 a_2092_8457# net45 3.35e-20
C1325 _073_ _092_ 4.32e-20
C1326 net46 a_10781_3311# 5.48e-21
C1327 _076_ _048_ 1.71e-19
C1328 _018_ a_4043_10143# 4.83e-21
C1329 a_2787_9845# a_3868_10217# 0.102f
C1330 _108_ a_13625_3317# 0.00776f
C1331 _060_ a_5081_4943# 1.12e-19
C1332 net31 _126_ 0.00137f
C1333 a_1211_7983# VPWR 3.44e-19
C1334 _074_ _102_ 0.415f
C1335 a_448_6549# a_1549_6794# 1.07e-20
C1336 clknet_2_1__leaf_clk a_3521_7361# 1.4e-19
C1337 _066_ a_10055_5487# 0.00936f
C1338 a_1476_6031# net30 1.86e-19
C1339 trim_mask\[0\] trim_val\[1\] 8.27e-22
C1340 net12 a_6090_10159# 1.39e-19
C1341 a_9595_1679# VPWR 0.519f
C1342 a_6210_4989# a_6316_5193# 0.0922f
C1343 net46 a_11801_4373# 0.17f
C1344 clknet_2_2__leaf_clk a_14172_1513# 8.02e-20
C1345 net55 _060_ 0.168f
C1346 net34 a_12992_8751# 4.15e-21
C1347 _095_ a_5455_4943# 3.66e-19
C1348 a_9802_4007# a_8583_3317# 1.13e-20
C1349 a_6099_10633# _020_ 0.119f
C1350 clknet_2_3__leaf_clk a_12520_7637# 9.5e-21
C1351 _110_ a_14981_4020# 9.22e-20
C1352 net19 a_9503_4399# 2.68e-19
C1353 a_1867_3317# a_3057_3689# 2.56e-19
C1354 a_2601_3285# a_2479_3689# 3.16e-19
C1355 a_2383_3689# a_2288_3677# 0.0498f
C1356 net33 _136_ 3.56e-20
C1357 a_11098_6691# VPWR 0.00135f
C1358 a_8215_9295# _063_ 4.53e-21
C1359 trim_mask\[1\] a_14702_3311# 1.17e-20
C1360 net28 a_5363_12559# 0.00665f
C1361 cal_itt\[2\] a_8935_6895# 4.48e-19
C1362 cal_itt\[1\] a_10864_7387# 3.34e-19
C1363 a_4349_8449# VPWR 0.206f
C1364 _108_ a_8583_3317# 6.55e-19
C1365 clknet_2_1__leaf_clk a_1095_12393# 6.19e-19
C1366 cal_itt\[0\] a_10137_4943# 6.48e-20
C1367 net14 a_1129_6273# 0.00982f
C1368 net51 net45 1.03e-19
C1369 net49 a_14540_3689# 0.00521f
C1370 cal_itt\[3\] _073_ 0.0366f
C1371 net19 a_7942_2223# 5.77e-19
C1372 a_15023_2767# _056_ 1.1e-19
C1373 _083_ a_6007_9839# 0.0912f
C1374 trim_mask\[0\] _118_ 0.202f
C1375 a_4425_6031# _059_ 3.64e-19
C1376 a_6633_9845# a_7079_10217# 2.28e-19
C1377 net12 a_5515_6005# 8.78e-19
C1378 _074_ _022_ 1.49e-19
C1379 clknet_2_1__leaf_clk a_1638_9839# 6.5e-19
C1380 net15 a_3208_7119# 0.00961f
C1381 a_15023_9839# _125_ 0.0117f
C1382 a_4609_9295# a_4696_8207# 5.87e-21
C1383 a_5177_9537# a_4871_8181# 1.22e-19
C1384 net4 _071_ 1.18e-21
C1385 _074_ a_6375_12021# 7.4e-19
C1386 net19 a_7939_10383# 0.0156f
C1387 net16 a_13557_8457# 6.13e-20
C1388 clknet_2_2__leaf_clk a_10016_1679# 2.28e-19
C1389 a_13697_4373# a_13519_4007# 0.00111f
C1390 _058_ a_10975_4105# 0.0068f
C1391 _103_ clk 0.00537f
C1392 _092_ a_3365_4943# 0.0386f
C1393 en_co_clk _103_ 1.3e-20
C1394 a_7527_4631# a_7677_4759# 0.0026f
C1395 _033_ a_10055_2767# 0.0622f
C1396 a_15023_9839# trimb[0] 0.00178f
C1397 net52 a_5535_8181# 8.83e-19
C1398 a_8473_5193# _107_ 0.00229f
C1399 _005_ result[1] 0.077f
C1400 a_3511_11471# VPWR 3.71e-19
C1401 a_5515_6005# a_5340_6031# 0.234f
C1402 net34 a_15111_9295# 1.65e-19
C1403 a_561_7119# a_561_6031# 0.0016f
C1404 _119_ a_9761_1679# 1.36e-20
C1405 a_14181_6031# _058_ 7.04e-20
C1406 _104_ trim_mask\[2\] 0.553f
C1407 a_1000_12381# _023_ 1.94e-20
C1408 a_10903_7261# en_co_clk 7.65e-20
C1409 net54 a_6197_4399# 1.28e-21
C1410 net45 _003_ 1.36e-21
C1411 _028_ a_7184_2339# 0.547f
C1412 net50 VPWR 0.429f
C1413 calibrate a_7104_3855# 7.93e-19
C1414 a_929_8757# a_2019_9055# 0.0424f
C1415 _037_ a_13279_7119# 0.00228f
C1416 calibrate a_7181_2589# 6.96e-20
C1417 clknet_0_clk a_4308_4917# 0.0127f
C1418 a_6633_9845# a_7723_10143# 0.0424f
C1419 a_2787_9845# a_3399_10217# 3.82e-19
C1420 a_7201_9813# a_6983_10217# 0.21f
C1421 _096_ calibrate 0.00876f
C1422 _018_ a_3208_10205# 0.158f
C1423 _001_ a_10864_7387# 0.236f
C1424 net28 a_579_10933# 9.15e-20
C1425 net44 _121_ 2.33e-20
C1426 _014_ a_3057_3689# 7.1e-20
C1427 a_11233_4405# _025_ 8.86e-20
C1428 a_13783_6183# a_13607_4943# 1.61e-20
C1429 _135_ a_13825_5185# 3.35e-21
C1430 _058_ a_13881_2741# 3.09e-19
C1431 state\[0\] a_4658_3427# 0.00186f
C1432 net44 a_8105_10383# 0.00488f
C1433 _051_ a_7527_4631# 0.00701f
C1434 a_14172_1513# ctln[2] 1.72e-20
C1435 a_395_4405# sample 0.00261f
C1436 _092_ cal_count\[3\] 0.0602f
C1437 net55 a_7939_3855# 4.04e-19
C1438 clknet_2_3__leaf_clk _048_ 2.42e-19
C1439 a_8731_9295# _041_ 3.11e-20
C1440 a_8583_3317# a_9004_3677# 0.0897f
C1441 net2 a_13050_7637# 3.27e-20
C1442 _063_ a_8298_5487# 0.0504f
C1443 a_10975_6031# a_11709_6273# 0.0531f
C1444 a_7262_5461# a_7571_4943# 4.96e-20
C1445 _038_ a_11141_6031# 0.207f
C1446 _051_ state\[1\] 0.355f
C1447 a_1644_12533# _078_ 1.41e-19
C1448 net55 a_4498_4373# 0.0307f
C1449 _078_ a_1476_4777# 1.81e-19
C1450 _041_ _037_ 1.72e-20
C1451 _014_ state\[1\] 1.65e-20
C1452 _105_ a_9003_3829# 9.38e-20
C1453 _107_ a_8583_3317# 0.00341f
C1454 net21 a_5363_12559# 0.201f
C1455 a_3597_10933# a_4674_10927# 1.46e-19
C1456 a_4995_7119# a_4259_6031# 8.93e-21
C1457 a_7140_2223# clk 5.04e-20
C1458 _029_ a_14172_4943# 5.34e-21
C1459 a_8381_9295# _070_ 1.44e-19
C1460 _060_ _093_ 0.00231f
C1461 net49 a_14335_2442# 2.47e-19
C1462 _104_ a_11045_3631# 6.81e-19
C1463 _121_ en_co_clk 0.00168f
C1464 _062_ a_10005_6031# 7.77e-21
C1465 net26 _043_ 9.81e-19
C1466 _078_ a_2174_8457# 1.95e-19
C1467 trim_mask\[0\] a_10137_4943# 6.4e-21
C1468 a_2689_8751# mask\[1\] 0.0423f
C1469 state\[2\] a_5177_1921# 0.00114f
C1470 _065_ _051_ 8.6e-23
C1471 a_3615_8207# a_4239_8573# 9.73e-19
C1472 clknet_2_0__leaf_clk a_4227_8207# 3.68e-19
C1473 a_3781_8207# a_4036_8207# 0.0605f
C1474 a_14099_1929# trim[2] 1.59e-19
C1475 a_5055_9295# VPWR 4.88e-19
C1476 net34 _132_ 0.0169f
C1477 a_6885_8372# a_6741_7361# 2.69e-21
C1478 mask\[5\] a_5998_11471# 0.0103f
C1479 net37 a_14972_5193# 0.00916f
C1480 net53 _000_ 0.00139f
C1481 a_1129_9813# a_1476_10217# 0.0512f
C1482 net34 net33 0.433f
C1483 clknet_2_3__leaf_clk a_11599_6397# 0.00499f
C1484 _101_ _083_ 0.0013f
C1485 _122_ _135_ 2.59e-19
C1486 _007_ a_1129_9813# 0.00229f
C1487 a_4959_9295# a_5221_9295# 0.00171f
C1488 a_5524_9295# a_5686_9661# 0.00645f
C1489 a_4863_4917# _099_ 6.65e-20
C1490 _030_ trim_val\[1\] 1.15e-19
C1491 net27 a_3511_11471# 0.00143f
C1492 mask\[3\] a_1677_9545# 0.0523f
C1493 a_5455_4943# calibrate 8.89e-21
C1494 net47 cal_itt\[0\] 0.28f
C1495 a_4993_6273# a_5449_6031# 4.2e-19
C1496 _015_ a_4617_3855# 7.21e-19
C1497 net45 a_7223_2465# 0.298f
C1498 _081_ a_2006_8751# 2.96e-20
C1499 _070_ clknet_0_clk 0.00135f
C1500 _108_ a_14894_3677# 3.59e-19
C1501 net15 a_3339_2767# 0.00307f
C1502 a_12059_2223# _031_ 1.38e-19
C1503 _062_ _099_ 2.25e-21
C1504 a_13562_8751# a_13279_8207# 9.75e-21
C1505 _104_ a_9595_1679# 1.78e-19
C1506 _009_ _021_ 2.08e-20
C1507 _110_ trim_mask\[2\] 0.515f
C1508 _074_ a_4512_12393# 6.62e-20
C1509 a_3208_7119# a_3399_7119# 4.61e-19
C1510 net32 a_14193_3285# 1.34e-19
C1511 net40 trimb[4] 0.0167f
C1512 mask\[7\] a_2910_12131# 9.44e-19
C1513 net12 a_6428_7119# 0.00883f
C1514 _047_ _109_ 6.2e-21
C1515 _050_ _028_ 0.182f
C1516 net40 _064_ 0.347f
C1517 net30 a_9369_4105# 2.29e-19
C1518 mask\[0\] a_6173_7119# 7.13e-21
C1519 clknet_2_0__leaf_clk a_395_2767# 1.56e-19
C1520 cal_itt\[0\] a_8820_6005# 0.066f
C1521 _039_ a_395_6031# 7.99e-19
C1522 a_1019_4399# cal 5.19e-19
C1523 net45 a_855_4105# 2.35e-19
C1524 clknet_2_0__leaf_clk a_455_3571# 1.81e-20
C1525 clknet_2_2__leaf_clk _025_ 0.149f
C1526 trim_mask\[0\] a_12424_3689# 5.76e-19
C1527 a_3840_8867# a_2857_7637# 5.14e-19
C1528 clknet_2_2__leaf_clk _026_ 0.0985f
C1529 a_14604_2339# VPWR 0.147f
C1530 a_13557_7369# VPWR 0.00254f
C1531 _123_ a_11479_9117# 0.00504f
C1532 _111_ a_11067_4405# 1.77e-19
C1533 _049_ a_4680_6031# 0.009f
C1534 a_1651_6005# a_1830_6031# 0.0074f
C1535 a_1476_6031# a_1585_6031# 0.00742f
C1536 net43 a_395_6031# 4.95e-19
C1537 cal_count\[3\] a_11045_5807# 0.00137f
C1538 _105_ a_8485_4943# 1.74e-20
C1539 _052_ _028_ 0.207f
C1540 a_395_7119# a_3208_7119# 6.41e-22
C1541 clknet_0_clk _090_ 9.53e-21
C1542 _055_ a_15023_1679# 3.12e-22
C1543 net43 a_4131_8207# 1.01e-19
C1544 _107_ a_7190_3855# 0.00403f
C1545 a_13715_5309# trim_val\[0\] 4.58e-20
C1546 a_2971_8457# a_2857_7637# 0.0105f
C1547 net43 a_6793_8970# 9.98e-21
C1548 net14 result[1] 5.96e-20
C1549 a_10861_7119# _136_ 1.02e-19
C1550 trim_val\[2\] a_14686_2339# 7.85e-19
C1551 _035_ a_11987_8757# 2.25e-20
C1552 _106_ VPWR 0.516f
C1553 _119_ a_11067_3017# 9.01e-19
C1554 _122_ a_14063_7093# 1.87e-19
C1555 net53 mask\[4\] 0.646f
C1556 a_3521_7361# _092_ 2.39e-20
C1557 net18 a_11059_7356# 0.00332f
C1558 net9 a_12341_8751# 0.00292f
C1559 a_4043_10143# _041_ 9.15e-20
C1560 _098_ _028_ 1.39e-20
C1561 net21 ctlp[6] 3.56e-20
C1562 a_4498_4373# _093_ 0.37f
C1563 a_763_8757# net45 2.73e-20
C1564 net31 net32 0.0992f
C1565 net2 VPWR 2.05f
C1566 trim_mask\[0\] a_12502_4765# 5.41e-21
C1567 a_9889_6873# en_co_clk 0.0307f
C1568 en_co_clk a_3273_4943# 0.171f
C1569 net40 _053_ 0.00149f
C1570 a_14193_3285# VPWR 0.215f
C1571 _110_ a_9719_1473# 0.134f
C1572 _078_ a_4609_9295# 0.0036f
C1573 net4 trim_mask\[1\] 2.12e-21
C1574 _049_ a_7190_3855# 0.105f
C1575 a_4308_4917# net41 2.68e-21
C1576 _003_ a_6316_5193# 7.81e-21
C1577 net29 result[6] 5.77e-20
C1578 a_4259_6031# a_4863_4917# 5.73e-21
C1579 _062_ a_5537_4943# 0.00153f
C1580 net18 a_12257_4777# 5.39e-20
C1581 a_395_7119# result[1] 0.0203f
C1582 trim_mask\[0\] a_11321_3855# 0.00145f
C1583 net50 _104_ 0.363f
C1584 _011_ a_745_10933# 0.00135f
C1585 a_1313_11989# a_579_10933# 4.89e-21
C1586 net47 a_13092_8029# 8.78e-19
C1587 _013_ a_1867_3317# 0.218f
C1588 _074_ _046_ 5.07e-20
C1589 net35 trim[4] 0.0161f
C1590 _085_ a_3852_12381# 1.78e-19
C1591 a_911_6031# a_1476_6031# 7.99e-20
C1592 a_11488_4765# a_10975_4105# 6.81e-19
C1593 _099_ a_3817_4697# 0.0337f
C1594 a_3667_3829# VPWR 0.613f
C1595 net20 net53 3.24e-20
C1596 trim_val\[2\] a_14347_1439# 0.0646f
C1597 a_14335_2442# a_14172_1513# 3.8e-20
C1598 _133_ _134_ 0.00631f
C1599 net8 a_14172_1513# 0.0184f
C1600 net9 a_10864_7387# 0.0014f
C1601 a_14000_4719# VPWR 2.76e-19
C1602 mask\[6\] ctlp[7] 5.34e-19
C1603 net9 a_12077_3285# 0.00368f
C1604 _074_ a_5067_9661# 0.00182f
C1605 cal_count\[3\] a_9003_3829# 9.29e-19
C1606 _033_ VPWR 0.844f
C1607 net18 a_11057_3855# 4.58e-20
C1608 a_15259_7637# net5 0.00102f
C1609 net47 a_10405_9295# 0.509f
C1610 _000_ _071_ 1.61e-20
C1611 net34 _136_ 2.33e-20
C1612 _096_ _015_ 2.48e-19
C1613 _002_ a_8301_8207# 0.00166f
C1614 net46 _055_ 0.00649f
C1615 net52 a_3133_11247# 0.00166f
C1616 a_8105_10383# a_8992_9955# 1.55e-20
C1617 net4 a_8749_3317# 0.0115f
C1618 _034_ a_4498_4373# 1.16e-19
C1619 _106_ a_9478_4105# 0.00183f
C1620 a_11233_4405# a_11801_4373# 0.186f
C1621 _110_ a_9595_1679# 0.0268f
C1622 clknet_2_1__leaf_clk a_1461_10357# 6.49e-21
C1623 net4 _060_ 1.05e-19
C1624 a_2143_7663# a_2489_7983# 0.0134f
C1625 net24 VPWR 1.61f
C1626 clknet_2_0__leaf_clk _099_ 3.7e-20
C1627 net44 a_6885_8372# 0.00187f
C1628 a_561_4405# a_1019_4399# 0.0311f
C1629 _065_ a_5535_8181# 0.0703f
C1630 _064_ _024_ 1.83e-19
C1631 _092_ a_6566_5193# 0.0588f
C1632 net31 VPWR 1.38f
C1633 _084_ VPWR 0.346f
C1634 _092_ _095_ 0.533f
C1635 a_8820_6005# trim_mask\[0\] 1.5e-19
C1636 a_14715_3615# trim[1] 3.74e-20
C1637 _051_ clknet_2_2__leaf_clk 5.36e-19
C1638 net15 net3 0.0611f
C1639 _039_ net30 9.56e-19
C1640 net30 a_8307_4719# 0.0396f
C1641 _108_ a_13512_4943# 0.0154f
C1642 mask\[7\] a_2014_11293# 0.00136f
C1643 clknet_2_0__leaf_clk a_1129_4373# 0.00145f
C1644 a_4443_1679# ctln[7] 2.13e-19
C1645 _058_ trim_val\[4\] 0.0193f
C1646 trim_val\[2\] a_15023_1679# 0.0044f
C1647 _042_ a_1129_9813# 2.1e-20
C1648 net45 a_5686_2045# 1.7e-19
C1649 a_3053_8457# clknet_2_0__leaf_clk 1.16e-20
C1650 net14 a_995_3530# 0.00531f
C1651 mask\[6\] _021_ 0.0173f
C1652 a_10329_1921# a_10569_1109# 0.00132f
C1653 _056_ _057_ 8.97e-20
C1654 a_10383_7093# _092_ 4.48e-20
C1655 net43 net30 0.156f
C1656 a_4131_8207# a_2857_7637# 4.44e-19
C1657 a_12436_9129# a_12341_8751# 0.0356f
C1658 a_4349_8449# clknet_0_clk 0.00358f
C1659 net41 a_2288_3677# 0.0212f
C1660 net12 a_5087_3855# 1.4e-20
C1661 net53 a_7091_9839# 0.00167f
C1662 clknet_2_1__leaf_clk a_7256_8029# 4.84e-20
C1663 _122_ a_13279_7119# 0.0601f
C1664 net18 a_10543_2455# 0.00703f
C1665 a_1467_7923# a_561_6031# 1.71e-21
C1666 net40 _130_ 0.0102f
C1667 _020_ clknet_2_3__leaf_clk 0.00112f
C1668 net33 a_14981_8235# 6.02e-19
C1669 clknet_2_3__leaf_clk a_11352_9661# 9.56e-19
C1670 net52 a_4165_10901# 1.3e-20
C1671 net11 a_6927_591# 0.00102f
C1672 a_6191_12559# clknet_2_1__leaf_clk 5.37e-20
C1673 net13 _099_ 0.00749f
C1674 net12 a_4443_1679# 8.01e-19
C1675 a_15023_10927# a_14983_9269# 2.71e-21
C1676 _094_ _050_ 0.00885f
C1677 _014_ _013_ 0.0694f
C1678 a_12520_7637# a_12664_8029# 0.00196f
C1679 clknet_2_1__leaf_clk _018_ 0.0945f
C1680 a_12344_8041# a_12454_8041# 0.00807f
C1681 net47 a_8717_10383# 0.00316f
C1682 a_8673_10625# a_9129_10383# 4.2e-19
C1683 _049_ a_5625_4943# 7.09e-20
C1684 a_4883_6397# VPWR 0.143f
C1685 net4 a_9361_3677# 4.25e-19
C1686 a_9296_9295# _035_ 7.31e-20
C1687 a_14807_8359# net2 0.138f
C1688 a_10785_1679# VPWR 6.15e-20
C1689 trim_mask\[4\] a_8583_3317# 0.229f
C1690 clknet_2_2__leaf_clk _031_ 0.0711f
C1691 mask\[7\] a_2787_10927# 0.0953f
C1692 _053_ _024_ 5.87e-20
C1693 _049_ a_4425_6031# 0.0219f
C1694 _047_ a_14655_4399# 4.27e-20
C1695 a_14281_4943# _058_ 9.77e-20
C1696 a_9761_1679# a_10111_1679# 0.23f
C1697 _122_ _041_ 0.0417f
C1698 _019_ a_4677_7882# 4.93e-20
C1699 cal_itt\[0\] _072_ 0.00264f
C1700 trim_mask\[1\] a_11509_3317# 0.554f
C1701 a_15083_4659# trim_val\[1\] 1.5e-19
C1702 a_13257_1141# a_13512_1501# 0.0642f
C1703 a_11292_1251# a_10787_1135# 0.00615f
C1704 net50 _110_ 0.0487f
C1705 trim_mask\[1\] a_14099_3017# 0.0595f
C1706 a_13183_3311# a_13459_3317# 1.15e-19
C1707 a_12424_3689# _030_ 0.00135f
C1708 _042_ a_3411_9839# 0.00176f
C1709 a_5878_9295# VPWR 0.00178f
C1710 net55 a_7571_4943# 0.00638f
C1711 a_11545_9049# _036_ 0.00106f
C1712 cal_itt\[0\] _068_ 0.0535f
C1713 _054_ VPWR 0.243f
C1714 en_co_clk a_11141_6031# 5.4e-20
C1715 a_2143_2229# a_2309_2229# 0.9f
C1716 a_1191_12393# result[6] 3.88e-19
C1717 a_1000_11293# a_1191_11305# 4.61e-19
C1718 mask\[4\] a_6007_9839# 0.0526f
C1719 a_2368_9955# _018_ 0.00373f
C1720 a_13257_4943# trim[4] 1.01e-20
C1721 net46 trim_val\[2\] 0.00547f
C1722 _041_ _063_ 1.61e-20
C1723 net4 a_7939_3855# 1.45e-20
C1724 _019_ a_4801_10159# 1.97e-19
C1725 _090_ net41 0.00615f
C1726 clknet_2_2__leaf_clk a_10781_3311# 2.86e-20
C1727 clknet_2_0__leaf_clk a_4259_6031# 0.404f
C1728 clknet_2_1__leaf_clk mask\[1\] 0.00928f
C1729 a_5524_9295# a_5633_9295# 0.00742f
C1730 a_5699_9269# a_5878_9295# 0.0074f
C1731 _129_ _134_ 0.0297f
C1732 a_2787_7119# _050_ 1.58e-21
C1733 net28 result[6] 0.0457f
C1734 net18 a_11016_6691# 0.00837f
C1735 a_1129_6273# VPWR 0.207f
C1736 net55 a_4576_3427# 3.84e-19
C1737 clknet_2_1__leaf_clk a_745_10933# 0.0253f
C1738 _084_ net27 0.14f
C1739 net4 a_4498_4373# 2.27e-21
C1740 _101_ a_4055_10927# 2.38e-19
C1741 net4 a_4864_1679# 1.7e-19
C1742 net9 _111_ 0.174f
C1743 a_8072_11721# a_8154_11721# 0.00477f
C1744 clknet_2_2__leaf_clk a_11801_4373# 5.58e-19
C1745 _106_ _104_ 0.00183f
C1746 a_4871_8181# _077_ 2.48e-19
C1747 a_4696_8207# a_5535_8181# 2.12e-19
C1748 net29 a_911_10217# 4.49e-22
C1749 _108_ a_11845_4765# 1.45e-19
C1750 _076_ _077_ 0.0132f
C1751 a_10655_2932# a_11149_2767# 3.49e-20
C1752 a_3868_7119# _049_ 0.00215f
C1753 _003_ a_6210_4989# 3.62e-21
C1754 _078_ a_6181_10633# 1.15e-19
C1755 a_8820_6005# a_8949_6281# 0.0626f
C1756 _063_ a_9839_3615# 4.46e-19
C1757 mask\[3\] a_3840_8867# 3.51e-21
C1758 a_9802_4007# a_9662_3855# 0.00106f
C1759 net4 a_8935_6895# 0.00167f
C1760 net9 a_12631_591# 0.172f
C1761 _072_ a_7569_7637# 0.0264f
C1762 net49 a_13459_3317# 0.0136f
C1763 a_2857_7637# net30 3.38e-20
C1764 a_745_12021# _078_ 0.00266f
C1765 _005_ a_1476_7119# 1.51e-19
C1766 net15 a_2961_9545# 0.00362f
C1767 VPWR ctln[5] 0.195f
C1768 net5 a_13933_6281# 5.38e-20
C1769 a_14063_7093# comp 3.56e-19
C1770 state\[0\] a_2601_3285# 2.3e-19
C1771 _071_ _053_ 0.00497f
C1772 mask\[0\] _005_ 3.99e-20
C1773 a_7184_2339# a_7181_2589# 2.36e-20
C1774 a_4677_7882# VPWR 0.258f
C1775 cal_count\[3\] _136_ 0.258f
C1776 a_2368_9955# mask\[1\] 1.08e-21
C1777 net13 a_4259_6031# 0.0153f
C1778 a_14083_3311# VPWR 0.144f
C1779 state\[2\] a_8307_4719# 3.59e-21
C1780 net1 a_2033_3317# 6.22e-20
C1781 _108_ a_9662_3855# 0.0318f
C1782 a_15023_8751# trimb[1] 0.00214f
C1783 net14 net3 0.0121f
C1784 a_3116_12533# net52 1.33e-21
C1785 _014_ a_2755_2601# 9.32e-19
C1786 net15 a_1660_11305# 2.21e-20
C1787 net33 a_14347_4917# 5.11e-20
C1788 a_9003_3829# _119_ 0.309f
C1789 a_7190_3855# trim_mask\[4\] 1.48e-20
C1790 clknet_2_0__leaf_clk a_4043_7093# 0.0582f
C1791 a_13111_6031# _135_ 0.149f
C1792 net15 mask\[0\] 0.124f
C1793 a_12520_7637# a_12824_7663# 3.11e-19
C1794 a_4801_10159# VPWR 3.11e-19
C1795 a_12344_8041# a_12430_7663# 0.00972f
C1796 a_12900_7663# a_14377_7983# 4.99e-20
C1797 state\[1\] a_2921_2589# 9.25e-20
C1798 _103_ _107_ 0.0467f
C1799 clknet_2_1__leaf_clk a_6796_12381# 4.56e-19
C1800 _092_ calibrate 0.0617f
C1801 _104_ _033_ 0.0252f
C1802 a_9802_4007# a_9572_2601# 5.98e-21
C1803 net42 clk 0.0128f
C1804 clknet_2_3__leaf_clk a_11583_4777# 1.94e-19
C1805 a_12599_3615# a_12691_2527# 1.06e-19
C1806 a_12249_7663# VPWR 0.104f
C1807 en_co_clk net42 2.04e-20
C1808 _065_ net22 8.97e-21
C1809 a_5731_4943# VPWR 3.86e-19
C1810 state\[2\] a_7010_3631# 0.00134f
C1811 net9 a_13257_1141# 0.00121f
C1812 a_7223_2465# a_8657_2229# 0.00133f
C1813 _002_ a_7088_7119# 8.81e-19
C1814 net12 a_4609_9295# 3.45e-20
C1815 _108_ a_9572_2601# 5.54e-22
C1816 _047_ trim[1] 0.122f
C1817 a_8381_9295# net2 1.18e-20
C1818 net23 net22 0.00148f
C1819 a_7088_7119# _050_ 5.7e-20
C1820 a_15023_6031# trim_mask\[0\] 3.43e-20
C1821 net47 _042_ 0.0705f
C1822 en_co_clk a_4091_5309# 0.0229f
C1823 _049_ _103_ 0.0125f
C1824 a_4993_6273# VPWR 0.206f
C1825 net13 a_4043_7093# 5.1e-19
C1826 mask\[2\] _040_ 0.0363f
C1827 net19 _070_ 0.0709f
C1828 a_6316_5193# a_6519_4631# 1.54e-19
C1829 _012_ a_937_3855# 3.65e-20
C1830 net47 a_11008_9295# 0.00291f
C1831 _053_ a_11204_7485# 0.00352f
C1832 a_7891_3617# _028_ 4.62e-19
C1833 _101_ mask\[4\] 0.366f
C1834 trim_mask\[3\] a_9747_2527# 0.0628f
C1835 trim_mask\[1\] net48 1.98e-20
C1836 net46 trim_mask\[0\] 0.352f
C1837 calibrate a_6906_2355# 7.33e-19
C1838 _093_ a_4576_3427# 7.18e-20
C1839 _106_ _110_ 0.0828f
C1840 clknet_0_clk _106_ 5.55e-20
C1841 a_8992_9955# a_9074_9955# 0.00477f
C1842 _108_ a_14471_591# 9.16e-20
C1843 net2 _110_ 1.31e-20
C1844 _123_ _053_ 0.181f
C1845 _017_ a_4036_8207# 0.158f
C1846 mask\[1\] a_6485_8181# 5.76e-20
C1847 _092_ a_8298_5487# 0.00248f
C1848 _070_ cal_itt\[1\] 1.5e-19
C1849 net2 clknet_0_clk 1.8e-20
C1850 net29 _085_ 1.86e-19
C1851 _118_ a_9369_4105# 0.0157f
C1852 a_4167_11471# a_5915_11721# 1.62e-21
C1853 a_13783_6183# a_14181_6031# 0.00369f
C1854 _135_ a_13825_6031# 0.0675f
C1855 a_6793_8970# a_6741_7361# 3.83e-20
C1856 _076_ a_6173_7119# 0.0151f
C1857 a_1461_10357# result[4] 9.76e-20
C1858 _050_ _096_ 0.0653f
C1859 _126_ trimb[1] 4.36e-19
C1860 a_3208_7119# VPWR 0.0846f
C1861 state\[2\] a_6822_4399# 2.81e-19
C1862 net28 a_911_10217# 1.51e-20
C1863 a_6181_10383# VPWR 6.87e-19
C1864 a_11016_6691# a_11023_5108# 2.15e-21
C1865 net40 trim[4] 0.00188f
C1866 net45 net55 1.01e-19
C1867 a_7256_8029# _092_ 4.12e-20
C1868 cal_count\[3\] _105_ 0.0584f
C1869 net25 a_448_9269# 0.179f
C1870 a_4815_3031# a_4609_1679# 2.81e-20
C1871 _104_ _054_ 0.0343f
C1872 trim_mask\[1\] a_13091_1141# 1.41e-20
C1873 a_8491_2229# clk 0.00365f
C1874 a_9443_6059# _091_ 0.128f
C1875 _035_ a_11258_9117# 6.37e-20
C1876 net34 a_15299_6575# 0.00396f
C1877 a_13715_5309# VPWR 0.142f
C1878 _005_ a_448_6549# 1.31e-20
C1879 a_11601_2229# a_12169_2197# 0.186f
C1880 a_11435_2229# a_11951_2601# 0.115f
C1881 _121_ _049_ 0.0172f
C1882 a_11709_6273# a_12165_6031# 4.2e-19
C1883 a_1660_11305# net25 8.95e-20
C1884 a_816_10205# a_1007_10217# 4.61e-19
C1885 net22 a_1019_6397# 0.00352f
C1886 net52 a_1476_10217# 9.14e-20
C1887 net19 a_9719_1473# 5.08e-21
C1888 a_1313_11989# result[6] 4.99e-19
C1889 net47 a_12344_8041# 0.205f
C1890 _085_ a_3431_12021# 0.00843f
C1891 _036_ a_13279_8207# 0.00228f
C1892 _110_ _033_ 0.00853f
C1893 clknet_2_3__leaf_clk a_10975_6031# 0.8f
C1894 _039_ a_911_6031# 6.6e-19
C1895 _074_ net45 0.0117f
C1896 _064_ trim_mask\[1\] 0.273f
C1897 a_561_9845# a_455_8181# 5.71e-21
C1898 net37 a_14981_4020# 0.0246f
C1899 a_14733_7983# VPWR 2.02e-19
C1900 clknet_0_clk _033_ 0.00723f
C1901 clknet_2_1__leaf_clk _041_ 0.0101f
C1902 net14 a_1476_7119# 4.01e-19
C1903 _010_ clknet_2_1__leaf_clk 0.0338f
C1904 net14 mask\[0\] 0.00272f
C1905 net44 a_2971_8457# 2.21e-20
C1906 a_7999_11231# a_7939_10383# 0.00384f
C1907 _096_ _098_ 4.83e-19
C1908 mask\[0\] a_3399_7119# 0.00449f
C1909 a_4222_10205# VPWR 2.24e-19
C1910 calibrate cal 0.0111f
C1911 a_12756_9117# VPWR 1.16e-19
C1912 net14 valid 0.00598f
C1913 _101_ a_2815_9447# 0.132f
C1914 VPWR result[1] 0.361f
C1915 net43 a_911_6031# 1.29e-20
C1916 net31 _110_ 6.29e-20
C1917 _078_ a_1638_6397# 1.06e-19
C1918 _070_ _001_ 0.105f
C1919 _101_ a_7091_9839# 2.69e-21
C1920 trim_mask\[0\] a_11343_3317# 1.21e-20
C1921 net4 _066_ 2.22e-19
C1922 net46 a_13869_4943# 0.00316f
C1923 trim_mask\[0\] a_11149_3017# 3.49e-20
C1924 trim_mask\[1\] a_10851_1653# 1.15e-20
C1925 _063_ a_9125_4943# 5.07e-19
C1926 mask\[2\] a_5177_9537# 1.89e-19
C1927 a_1493_5487# a_395_4405# 3.34e-20
C1928 a_1279_9129# net45 1.49e-19
C1929 a_561_9845# a_1019_9839# 0.0276f
C1930 _035_ a_10383_7093# 1.83e-21
C1931 net19 a_9595_1679# 0.00104f
C1932 _115_ net48 0.0183f
C1933 _134_ a_14379_6397# 6.26e-19
C1934 a_13279_7119# a_13111_6031# 1.54e-20
C1935 _078_ a_5535_8181# 0.223f
C1936 a_6191_12559# a_6927_12559# 5.42e-20
C1937 _064_ a_8749_3317# 3.71e-20
C1938 a_395_7119# a_1476_7119# 0.102f
C1939 a_6909_10933# a_7355_11305# 2.28e-19
C1940 _031_ net8 0.00114f
C1941 calibrate a_6737_4719# 0.0509f
C1942 a_8731_9295# a_8839_9661# 0.0572f
C1943 _058_ a_14702_3311# 3.76e-21
C1944 net51 _003_ 0.00476f
C1945 net18 a_10699_3311# 0.00956f
C1946 mask\[0\] a_395_7119# 6.38e-21
C1947 net43 a_5691_7637# 0.0504f
C1948 _099_ a_3751_4765# 0.00174f
C1949 a_3817_4697# _097_ 2.46e-19
C1950 _058_ a_13693_3883# 3.85e-20
C1951 mask\[5\] a_6445_10383# 9.24e-19
C1952 _050_ a_5455_4943# 6.6e-19
C1953 cal_itt\[2\] _069_ 1.61e-19
C1954 en_co_clk a_4886_4399# 1.27e-19
C1955 _064_ a_10977_2543# 0.00153f
C1956 a_5087_3855# _089_ 8.68e-20
C1957 a_11059_7356# VPWR 0.207f
C1958 a_11425_5487# _024_ 1.86e-19
C1959 a_12599_3615# VPWR 0.353f
C1960 cal_itt\[2\] a_8022_7119# 0.0416f
C1961 net2 a_14564_6397# 1.13e-20
C1962 _078_ _082_ 0.055f
C1963 _101_ _081_ 0.024f
C1964 cal_itt\[0\] _065_ 0.0235f
C1965 net12 a_6181_10633# 0.00238f
C1966 net3 a_5363_4719# 2.03e-19
C1967 a_10747_8970# _122_ 8.88e-21
C1968 net14 _079_ 0.0167f
C1969 net16 trim_val\[0\] 0.0338f
C1970 net50 a_11057_4105# 0.0024f
C1971 a_12061_7669# a_12520_7637# 0.0849f
C1972 cal_count\[2\] a_15289_7119# 2.23e-20
C1973 mask\[3\] a_5221_9295# 4.33e-20
C1974 clknet_2_0__leaf_clk _097_ 1.42e-19
C1975 trim_mask\[3\] a_10676_1679# 0.00393f
C1976 calibrate a_5536_4399# 3.97e-19
C1977 mask\[6\] a_4866_11293# 0.00198f
C1978 _086_ a_1313_10901# 6.54e-20
C1979 a_1585_4777# _099_ 2.14e-20
C1980 a_4443_1679# a_4609_1679# 0.887f
C1981 _115_ a_13091_1141# 0.00138f
C1982 _092_ _015_ 4.53e-21
C1983 net20 a_6375_12021# 0.0263f
C1984 a_6191_12559# _009_ 1.44e-19
C1985 _045_ a_6541_12021# 3.32e-19
C1986 a_4167_6575# a_4259_6031# 1.36e-19
C1987 a_5455_4943# _098_ 1.11e-20
C1988 net28 _085_ 0.127f
C1989 a_1644_12533# net29 0.173f
C1990 a_12257_4777# VPWR 1.49e-19
C1991 _070_ a_7916_8041# 0.00102f
C1992 trim_mask\[1\] trim[0] 7.26e-19
C1993 net45 _093_ 0.0295f
C1994 net2 a_13091_4943# 2.97e-19
C1995 clknet_0_clk _054_ 3.05e-19
C1996 _049_ a_3273_4943# 0.00104f
C1997 a_1129_4373# a_1585_4777# 4.2e-19
C1998 net46 _030_ 0.0539f
C1999 a_911_4777# a_1173_4765# 0.00171f
C2000 a_10405_9295# a_10774_9661# 4.45e-20
C2001 a_10864_9269# a_10593_9295# 7.79e-20
C2002 a_1095_11305# a_1203_10927# 0.0572f
C2003 mask\[0\] a_4222_7119# 0.00198f
C2004 a_1313_10901# _102_ 1.46e-19
C2005 a_14063_7093# a_14199_7369# 0.0718f
C2006 a_1660_11305# a_1769_11305# 0.00742f
C2007 a_3339_2767# VPWR 0.289f
C2008 a_1835_11231# a_2014_11293# 0.0074f
C2009 net4 a_4576_3427# 5.8e-20
C2010 calibrate a_561_4405# 0.26f
C2011 a_3273_4943# a_3388_4631# 4.52e-20
C2012 _136_ a_11679_4777# 3.85e-19
C2013 net43 a_4775_6031# 3.35e-20
C2014 a_995_3530# VPWR 0.259f
C2015 net12 _051_ 0.23f
C2016 net16 _126_ 0.00142f
C2017 net44 a_4131_8207# 0.152f
C2018 net18 a_10593_9295# 0.00126f
C2019 clknet_2_1__leaf_clk _002_ 0.00753f
C2020 a_13257_4943# a_13625_3317# 5.9e-22
C2021 _072_ a_7723_6807# 0.149f
C2022 net40 a_10245_5193# 0.0105f
C2023 VPWR rstn 0.198f
C2024 a_11141_6031# _108_ 1.06e-19
C2025 net44 a_6793_8970# 0.00106f
C2026 a_11057_3855# VPWR 6.98e-20
C2027 a_14471_12559# a_15023_12559# 8.52e-19
C2028 a_8912_2589# VPWR 0.0851f
C2029 cal_itt\[0\] a_9761_8457# 3.23e-19
C2030 net55 a_4905_3855# 8.55e-19
C2031 _043_ net4 1.61e-20
C2032 _053_ a_10781_5807# 0.00306f
C2033 a_8673_10625# VPWR 0.215f
C2034 net45 a_2865_4460# 9.84e-19
C2035 trim_mask\[0\] a_7527_4631# 0.228f
C2036 a_11814_9295# _041_ 2.1e-19
C2037 net29 a_2828_12131# 0.105f
C2038 a_2174_8457# _040_ 4.96e-19
C2039 trim_mask\[4\] a_11149_2767# 1.17e-19
C2040 a_13881_1653# _114_ 0.118f
C2041 _042_ a_4443_9295# 4.43e-19
C2042 a_5340_6031# _051_ 1.6e-19
C2043 a_8298_5487# a_9003_3829# 6.1e-19
C2044 a_1679_10633# a_1476_10217# 6.39e-20
C2045 net26 a_2787_9845# 4.33e-20
C2046 net46 a_8298_2767# 0.0262f
C2047 _122_ a_11369_7119# 0.00166f
C2048 _041_ a_6485_8181# 3.19e-20
C2049 trim_mask\[1\] a_14335_4020# 1.16e-20
C2050 net18 _027_ 1.1e-19
C2051 _095_ a_4266_4943# 2.62e-21
C2052 net14 a_448_6549# 1.67e-19
C2053 net43 a_1129_9813# 0.174f
C2054 a_4043_7093# a_4167_6575# 8.51e-19
C2055 net16 a_12153_8757# 1.92e-21
C2056 _043_ a_8360_10383# 7.3e-22
C2057 clknet_0_clk a_4677_7882# 0.0326f
C2058 net52 _042_ 0.0113f
C2059 _048_ a_5087_3855# 2.01e-20
C2060 _006_ a_455_8181# 0.00974f
C2061 net46 a_9681_2601# 6.54e-19
C2062 _005_ a_1125_7663# 6.78e-19
C2063 a_2857_5461# net55 6.68e-20
C2064 a_3667_3829# net41 1.53e-19
C2065 state\[0\] a_4617_4105# 1.27e-19
C2066 a_10543_2455# VPWR 0.277f
C2067 a_7164_11293# VPWR 0.0859f
C2068 a_8215_9295# _035_ 1.88e-19
C2069 net43 a_3411_7485# 0.0122f
C2070 a_6056_8359# a_6198_8534# 0.00557f
C2071 _010_ a_4866_12381# 4.67e-20
C2072 _046_ a_4055_10927# 4.66e-20
C2073 clknet_2_1__leaf_clk a_3615_8207# 0.00248f
C2074 net49 trim[1] 1.86e-19
C2075 a_2828_12131# a_3431_12021# 4.15e-19
C2076 net2 a_6523_7119# 2.27e-20
C2077 _063_ a_8389_5193# 8.95e-19
C2078 net24 a_2775_9071# 4.81e-19
C2079 _094_ _099_ 5.11e-20
C2080 a_1844_9129# a_2006_8751# 0.00645f
C2081 trim_mask\[4\] a_9662_3855# 0.00114f
C2082 _058_ a_14237_3677# 2.61e-19
C2083 a_395_7119# a_448_6549# 0.0131f
C2084 a_14172_1513# a_15023_1135# 5.37e-19
C2085 a_911_6031# a_1173_6031# 0.00171f
C2086 a_10405_9295# _065_ 1.8e-20
C2087 a_448_7637# net45 6.32e-21
C2088 trim_mask\[1\] a_15023_2767# 0.00105f
C2089 a_11343_3317# _030_ 2.88e-20
C2090 a_7723_10143# _065_ 2.03e-21
C2091 net47 _133_ 1.57e-19
C2092 a_1019_9839# _006_ 1.1e-20
C2093 _053_ a_7939_3855# 0.0358f
C2094 a_9471_9269# net4 0.00105f
C2095 _127_ a_15111_9295# 8.17e-20
C2096 cal_itt\[0\] _067_ 0.942f
C2097 a_9296_9295# a_9463_8725# 0.0021f
C2098 _085_ net21 8.48e-20
C2099 a_7109_11989# ctlp[6] 0.00104f
C2100 a_11023_5108# a_10699_3311# 9.43e-22
C2101 a_6835_7669# a_8025_8041# 2.56e-19
C2102 net46 a_11951_2601# 0.153f
C2103 net43 a_3411_9839# 0.0122f
C2104 a_14931_591# VPWR 0.244f
C2105 clknet_0_clk a_4993_6273# 2.53e-20
C2106 net44 net30 0.0123f
C2107 a_15159_9269# _125_ 0.243f
C2108 _009_ a_6796_12381# 0.158f
C2109 clknet_2_0__leaf_clk a_3748_6281# 0.0127f
C2110 a_8767_591# VPWR 0.276f
C2111 a_6375_12021# a_6987_12393# 0.00188f
C2112 _078_ net22 0.0116f
C2113 net29 a_1000_12381# 8.96e-20
C2114 net50 a_11067_4405# 0.00315f
C2115 net9 trim_mask\[2\] 0.0102f
C2116 trim_mask\[0\] a_11233_4405# 0.00497f
C2117 net33 _135_ 2.17e-20
C2118 a_6191_12559# mask\[6\] 7.31e-22
C2119 trim_mask\[4\] a_9572_2601# 1.95e-22
C2120 a_2033_3317# a_2143_2229# 1.35e-20
C2121 a_1867_3317# a_2309_2229# 6.94e-21
C2122 net44 a_5221_9295# 0.0043f
C2123 trim_val\[3\] a_11292_1251# 0.191f
C2124 a_11016_6691# VPWR 0.165f
C2125 net3 VPWR 2.8f
C2126 a_455_12533# net29 2.96e-19
C2127 mask\[6\] _018_ 3.93e-20
C2128 a_14377_9545# a_14236_8457# 6.54e-21
C2129 _112_ a_13183_3311# 7.61e-19
C2130 mask\[5\] a_7355_11305# 1.48e-19
C2131 net18 _117_ 8.86e-19
C2132 net9 a_12213_2589# 4.44e-19
C2133 mask\[0\] a_2313_6183# 0.163f
C2134 _086_ result[5] 3.98e-19
C2135 _007_ net23 3.02e-20
C2136 _100_ a_4617_4105# 0.00161f
C2137 _104_ a_11413_2767# 6.81e-19
C2138 net16 _114_ 8.85e-19
C2139 a_13142_7271# _131_ 0.00179f
C2140 a_14063_7093# a_14422_7093# 0.141f
C2141 net14 a_1229_8457# 0.00101f
C2142 a_4609_9295# _040_ 1.3e-20
C2143 net30 clk 1.03f
C2144 en_co_clk net30 0.00826f
C2145 net15 a_579_10933# 6.55e-22
C2146 a_13607_1513# VPWR 0.226f
C2147 net4 net45 0.179f
C2148 net19 _106_ 0.159f
C2149 _120_ _048_ 0.0423f
C2150 a_2857_7637# a_3411_7485# 9.92e-19
C2151 net12 a_5535_8181# 0.0021f
C2152 net30 a_9084_4515# 0.0328f
C2153 a_14249_8725# net2 5.27e-19
C2154 net28 a_2828_12131# 0.0184f
C2155 net4 _058_ 4.91e-20
C2156 a_10111_1679# trim_val\[3\] 1.48e-20
C2157 net19 net2 0.00927f
C2158 a_12341_8751# _037_ 1.56e-19
C2159 VPWR trimb[1] 0.537f
C2160 a_3529_6281# a_4425_6031# 9.28e-20
C2161 net6 a_395_591# 0.00163f
C2162 a_10872_1455# a_10787_1135# 1.48e-19
C2163 _094_ a_4259_6031# 0.222f
C2164 a_13715_5309# _110_ 2.02e-20
C2165 a_2857_5461# _093_ 2.69e-21
C2166 a_15023_6031# a_15083_4659# 2.58e-19
C2167 trim_val\[4\] a_10975_4105# 5.6e-20
C2168 _132_ a_14063_7093# 0.00272f
C2169 a_14335_7895# _130_ 5.4e-20
C2170 a_14540_3689# _055_ 0.00518f
C2171 net33 _127_ 0.0235f
C2172 a_12992_8751# _041_ 0.044f
C2173 ctlp[0] result[7] 0.144f
C2174 net45 a_3303_7119# 6.88e-20
C2175 a_2491_3311# a_2143_2229# 2.78e-20
C2176 net16 a_13050_7637# 7.99e-19
C2177 _136_ a_8298_5487# 8.86e-19
C2178 _019_ a_2961_9545# 6.51e-21
C2179 a_6906_2355# a_7184_2339# 0.125f
C2180 _026_ a_12169_2197# 7.06e-19
C2181 clknet_2_1__leaf_clk a_3249_9295# 3.7e-19
C2182 mask\[6\] a_745_10933# 4.14e-20
C2183 _095_ a_3365_4943# 0.0543f
C2184 a_3868_10217# _083_ 4.68e-23
C2185 net4 a_9693_8029# 1.92e-19
C2186 _113_ a_13693_3883# 0.00141f
C2187 _112_ net49 5.7e-19
C2188 _002_ a_6007_7119# 0.00358f
C2189 _063_ a_10005_6031# 0.00133f
C2190 _092_ a_10781_5487# 0.00303f
C2191 _104_ a_11057_3855# 0.00354f
C2192 _067_ trim_mask\[0\] 0.0937f
C2193 trim_val\[2\] ctln[2] 1.8e-20
C2194 cal_count\[3\] _119_ 3.29e-21
C2195 net42 _107_ 0.0111f
C2196 _014_ a_2309_2229# 0.217f
C2197 a_6007_7119# _050_ 3.23e-20
C2198 a_13881_1653# VPWR 0.239f
C2199 cal_itt\[1\] _106_ 8.72e-20
C2200 a_8673_10625# a_8455_10383# 0.21f
C2201 a_7939_10383# a_9020_10383# 0.102f
C2202 a_8105_10383# a_9195_10357# 0.0424f
C2203 a_10239_9295# _053_ 1.98e-21
C2204 net47 _129_ 1.66e-19
C2205 trim_mask\[1\] a_9664_3689# 2.78e-19
C2206 _078_ a_4165_10901# 1.14e-21
C2207 net14 a_1125_7663# 0.0087f
C2208 net47 a_9405_9295# 8.66e-19
C2209 a_14172_4943# _058_ 0.00185f
C2210 net2 cal_itt\[1\] 5.03e-19
C2211 state\[1\] a_2877_2197# 2.01e-19
C2212 net55 a_6210_4989# 1.38e-19
C2213 net54 a_5363_4719# 0.0492f
C2214 net19 _033_ 0.00928f
C2215 _016_ a_4030_7485# 1.55e-20
C2216 a_11895_7669# a_10903_7261# 0.00162f
C2217 _037_ a_10864_7387# 8.53e-19
C2218 a_10055_2767# _027_ 2.72e-19
C2219 a_8083_8181# VPWR 0.266f
C2220 _051_ a_5691_2741# 0.0551f
C2221 trim_mask\[1\] a_10689_2223# 1.38e-20
C2222 _018_ a_1763_9295# 3.21e-20
C2223 _049_ net42 0.0459f
C2224 _097_ a_2948_3689# 9.37e-19
C2225 _028_ a_7942_2223# 0.17f
C2226 a_4043_7093# _094_ 1.33e-20
C2227 _034_ a_2857_5461# 4.34e-20
C2228 a_8491_2229# a_9115_2223# 9.73e-19
C2229 _134_ en_co_clk 0.0584f
C2230 trim_mask\[0\] clknet_2_2__leaf_clk 0.0931f
C2231 _051_ a_7524_2223# 2.87e-19
C2232 _104_ a_10543_2455# 0.201f
C2233 a_1000_12381# a_1191_12393# 4.61e-19
C2234 net33 a_14604_3017# 0.00219f
C2235 _049_ a_4091_5309# 0.00495f
C2236 _092_ _050_ 0.882f
C2237 mask\[6\] a_6796_12381# 2.83e-21
C2238 a_8749_3317# a_9664_3689# 0.125f
C2239 net16 net32 1.21e-20
C2240 a_14334_1135# VPWR 7.7e-19
C2241 a_2961_9545# VPWR 0.177f
C2242 _051_ a_5726_5807# 5.53e-21
C2243 _064_ _066_ 6.91e-19
C2244 _110_ a_12599_3615# 5.34e-21
C2245 net28 a_1000_12381# 0.0037f
C2246 trim_mask\[2\] trim_mask\[3\] 0.0993f
C2247 _135_ _136_ 0.189f
C2248 _070_ _062_ 3.11e-20
C2249 a_448_9269# VPWR 0.3f
C2250 mask\[3\] a_5691_7637# 1.65e-21
C2251 calibrate a_7010_3311# 0.0711f
C2252 a_1651_10143# _082_ 3.18e-19
C2253 _096_ _087_ 3.13e-20
C2254 a_1660_11305# VPWR 0.328f
C2255 a_455_12533# net28 0.225f
C2256 trim_mask\[1\] a_10781_3631# 8.34e-19
C2257 a_6835_7669# a_6173_7119# 1.92e-19
C2258 trim_mask\[2\] a_10689_2543# 2.72e-20
C2259 a_4609_9295# a_5177_9537# 0.173f
C2260 a_1476_7119# VPWR 0.323f
C2261 net30 _059_ 1.8e-20
C2262 a_4443_9295# a_4959_9295# 0.114f
C2263 a_11709_6273# VPWR 0.213f
C2264 a_12424_3689# a_12533_3689# 0.00742f
C2265 trim_mask\[3\] a_12213_2589# 4.63e-20
C2266 a_11859_3689# a_11967_3311# 0.0572f
C2267 a_12599_3615# a_12778_3677# 0.0074f
C2268 a_7939_10383# a_8731_9295# 1.23e-20
C2269 mask\[0\] VPWR 1.44f
C2270 a_8105_10383# a_8949_9537# 4e-21
C2271 a_8673_10625# a_8381_9295# 1.8e-21
C2272 _092_ _052_ 3.03e-19
C2273 net2 _001_ 0.148f
C2274 VPWR valid 0.59f
C2275 a_3597_10933# a_4165_10901# 0.186f
C2276 clknet_2_0__leaf_clk a_4308_4917# 3.69e-20
C2277 a_579_12021# result[7] 0.00352f
C2278 _101_ a_3781_8207# 3.1e-20
C2279 a_6927_591# ctln[6] 0.342f
C2280 state\[2\] clk 0.0574f
C2281 a_579_10933# net25 2.09e-19
C2282 a_15023_9839# a_15023_8751# 0.00222f
C2283 _090_ a_4863_4917# 0.001f
C2284 a_11709_6273# a_12218_6397# 2.6e-19
C2285 a_2953_9845# a_3411_9839# 0.0346f
C2286 mask\[3\] a_5089_10159# 4.58e-19
C2287 a_11141_6031# a_11587_6031# 2.28e-19
C2288 _002_ cal_itt\[3\] 1.29e-19
C2289 net17 ctlp[3] 0.00723f
C2290 a_11059_7356# a_10699_5487# 8.26e-20
C2291 _092_ _098_ 0.0892f
C2292 a_3273_4943# a_3123_3615# 4.66e-21
C2293 _096_ _099_ 0.28f
C2294 a_12323_4703# a_12424_3689# 2.15e-22
C2295 _058_ a_11509_3317# 0.00399f
C2296 _014_ a_3110_3311# 5.82e-20
C2297 a_7019_4407# a_6927_3311# 7.24e-21
C2298 _023_ _007_ 2.04e-20
C2299 net22 _004_ 0.00877f
C2300 a_2953_7119# a_3303_7119# 0.22f
C2301 a_2787_7119# a_4043_7093# 0.0436f
C2302 _058_ a_14099_3017# 6.04e-19
C2303 net14 a_579_10933# 0.0078f
C2304 state\[0\] clk 2.86e-19
C2305 a_11008_9295# _065_ 1.61e-20
C2306 en_co_clk state\[0\] 0.00123f
C2307 _069_ a_10043_7983# 0.00189f
C2308 net15 a_2564_2589# 0.00169f
C2309 _050_ a_6906_2355# 7.7e-19
C2310 net13 a_4709_2773# 0.00396f
C2311 net29 a_745_12021# 0.00662f
C2312 a_5537_4105# VPWR 0.00469f
C2313 a_9317_3285# a_9207_3311# 0.0977f
C2314 _053_ _066_ 0.0928f
C2315 a_8298_5487# _105_ 0.00233f
C2316 trim_mask\[2\] a_13415_2442# 0.036f
C2317 net16 VPWR 2.18f
C2318 a_911_10217# a_1173_10205# 0.00171f
C2319 a_1129_9813# a_1585_10217# 4.2e-19
C2320 clknet_2_3__leaf_clk a_10864_9269# 0.0268f
C2321 _051_ _089_ 0.00231f
C2322 a_12148_4777# a_12257_4777# 0.00742f
C2323 a_12323_4703# a_12502_4765# 0.0074f
C2324 _024_ a_12310_4399# 4.33e-20
C2325 a_11583_4777# a_11691_4399# 0.0572f
C2326 _058_ a_9166_4515# 4.73e-20
C2327 a_10055_2767# _117_ 5.57e-19
C2328 trim_mask\[3\] a_9719_1473# 2e-20
C2329 a_15023_5487# _047_ 0.00251f
C2330 net18 clknet_2_3__leaf_clk 0.0822f
C2331 _007_ a_816_10205# 0.158f
C2332 a_13257_4943# a_13512_4943# 0.0564f
C2333 a_13607_4943# a_14172_4943# 7.99e-20
C2334 a_13091_4943# a_13715_5309# 9.73e-19
C2335 clknet_2_2__leaf_clk a_13869_4943# 2.34e-19
C2336 _052_ a_6906_2355# 2.8e-19
C2337 a_6197_12015# VPWR 0.00572f
C2338 a_12516_2601# a_12625_2601# 0.00742f
C2339 a_12691_2527# a_12870_2589# 0.0074f
C2340 a_12169_2197# _031_ 1.76e-19
C2341 a_11951_2601# a_12059_2223# 0.0572f
C2342 net45 a_7689_2589# 9.54e-19
C2343 _051_ a_4609_1679# 2.52e-19
C2344 a_5915_10927# a_5997_11247# 0.00393f
C2345 a_8215_9295# a_9296_9295# 0.102f
C2346 _000_ a_9471_9269# 9.79e-21
C2347 calibrate a_3148_4399# 9.09e-20
C2348 _079_ VPWR 0.122f
C2349 mask\[4\] _043_ 0.0799f
C2350 clknet_2_1__leaf_clk a_2019_9055# 5.21e-21
C2351 net26 a_763_8757# 4.53e-21
C2352 trim_val\[4\] a_9099_3689# 1.05e-19
C2353 _074_ a_2787_9845# 2.72e-20
C2354 _136_ a_14649_6031# 1.17e-19
C2355 clknet_2_0__leaf_clk a_2288_3677# 9.35e-19
C2356 a_5455_4943# _087_ 0.0764f
C2357 net4 _069_ 0.0991f
C2358 a_816_4765# _014_ 1.1e-21
C2359 net2 a_7916_8041# 1.43e-20
C2360 _124_ _123_ 0.0129f
C2361 a_10699_3311# VPWR 0.22f
C2362 clknet_2_3__leaf_clk a_12165_6031# 0.00112f
C2363 net20 a_7456_12393# 0.00215f
C2364 net4 a_8022_7119# 0.0159f
C2365 a_4973_2773# VPWR 1.08e-19
C2366 net19 ctln[5] 0.00146f
C2367 _118_ a_10270_4105# 8.55e-19
C2368 _053_ a_7571_4943# 1.84e-20
C2369 trim_mask\[3\] a_9595_1679# 0.002f
C2370 cal_count\[2\] _134_ 0.0359f
C2371 a_395_9845# net25 0.00131f
C2372 _048_ a_7677_4759# 3.75e-19
C2373 a_5455_4943# _099_ 2.83e-19
C2374 calibrate a_1019_4399# 0.0256f
C2375 mask\[1\] a_3317_8207# 1.91e-20
C2376 _010_ mask\[6\] 3.7e-19
C2377 a_14335_2442# trim_val\[2\] 0.00255f
C2378 _086_ a_1579_11471# 0.00151f
C2379 net54 VPWR 0.751f
C2380 trim_val\[2\] net8 0.179f
C2381 a_6822_4105# a_7021_4105# 3.58e-19
C2382 _045_ _042_ 1.83e-21
C2383 net14 a_395_9845# 0.00725f
C2384 _121_ a_3529_6281# 3.7e-19
C2385 en_co_clk _100_ 8.95e-19
C2386 a_4259_6031# _096_ 0.00163f
C2387 net45 a_3057_4719# 1.02e-19
C2388 a_15023_9839# _126_ 0.0104f
C2389 _090_ a_3817_4697# 0.147f
C2390 a_10990_7485# _038_ 0.00102f
C2391 clknet_2_3__leaf_clk trim_val\[0\] 3.62e-22
C2392 _049_ a_4886_4399# 0.014f
C2393 net34 _135_ 1.32e-20
C2394 a_11622_7485# a_11369_7119# 4.61e-19
C2395 a_579_10933# a_1769_11305# 2.56e-19
C2396 _074_ a_2092_8457# 1.04e-20
C2397 _101_ a_5686_9661# 1.37e-19
C2398 a_6099_10633# a_6467_9845# 0.0111f
C2399 _059_ state\[2\] 3.46e-20
C2400 clknet_2_2__leaf_clk _030_ 0.179f
C2401 a_9003_3829# a_9207_3311# 6.53e-20
C2402 trim_mask\[0\] a_14540_3689# 3.4e-19
C2403 a_7262_5461# _088_ 8.22e-20
C2404 a_448_6549# VPWR 0.311f
C2405 _111_ a_13697_4373# 3.52e-20
C2406 clknet_2_0__leaf_clk _090_ 0.00154f
C2407 a_5547_5603# _050_ 0.137f
C2408 net4 a_3386_2223# 1.46e-19
C2409 net44 a_5691_7637# 6.17e-19
C2410 _051_ _048_ 0.486f
C2411 clknet_2_3__leaf_clk a_11575_8790# 2.46e-19
C2412 net37 net2 0.61f
C2413 a_8307_4943# clknet_2_2__leaf_clk 7.63e-20
C2414 a_6099_10633# VPWR 0.226f
C2415 a_10593_9295# VPWR 0.104f
C2416 net43 _072_ 0.0964f
C2417 a_13279_7119# _136_ 0.00109f
C2418 _048_ _014_ 1.92e-19
C2419 _035_ _041_ 0.126f
C2420 _123_ a_13356_7369# 0.00285f
C2421 clknet_0_clk net3 8.51e-19
C2422 a_8993_9295# cal_itt\[0\] 8.9e-20
C2423 a_745_12021# a_1191_12393# 2.28e-19
C2424 net43 _068_ 1.05e-19
C2425 _052_ a_6737_4719# 0.00891f
C2426 a_6519_4631# _088_ 1.81e-20
C2427 a_6316_5193# a_6763_5193# 0.0551f
C2428 net14 a_2564_2589# 1.74e-19
C2429 a_4043_12393# _078_ 1.01e-19
C2430 a_6743_10933# mask\[4\] 9.76e-21
C2431 a_6099_10633# a_5699_9269# 1.05e-20
C2432 a_6191_12559# ctlp[7] 3.27e-19
C2433 VPWR trimb[3] 0.553f
C2434 _050_ a_5536_4399# 5.24e-20
C2435 clknet_2_2__leaf_clk a_8298_2767# 1.71f
C2436 a_6541_12021# net12 8.37e-19
C2437 net28 a_745_12021# 0.0133f
C2438 net50 trim_mask\[3\] 0.158f
C2439 _078_ a_1476_10217# 0.0108f
C2440 _074_ net51 5.04e-19
C2441 net30 a_9802_4007# 7.15e-20
C2442 _098_ a_6737_4719# 0.0523f
C2443 net34 _127_ 1.73e-19
C2444 net2 a_13193_6031# 0.00236f
C2445 _110_ a_13607_1513# 3.4e-20
C2446 a_11116_8983# net2 2.09e-21
C2447 a_5455_4943# a_5537_4943# 0.00578f
C2448 _027_ VPWR 0.706f
C2449 _078_ _007_ 1.77e-19
C2450 a_11016_6691# a_10699_5487# 5.22e-19
C2451 net47 a_13100_8751# 6.59e-19
C2452 net13 _090_ 0.0117f
C2453 net47 _038_ 4.05e-20
C2454 a_3615_8207# a_4805_8207# 2.56e-19
C2455 clknet_2_2__leaf_clk a_9681_2601# 4.62e-19
C2456 _085_ ctlp[1] 0.0037f
C2457 _062_ net50 1.8e-19
C2458 net4 a_8657_2229# 2.27e-19
C2459 net43 net52 0.151f
C2460 net30 _108_ 0.0409f
C2461 clknet_2_1__leaf_clk a_3053_8457# 0.00544f
C2462 net43 a_816_7119# 5.45e-19
C2463 a_7019_4407# VPWR 0.26f
C2464 cal_count\[3\] a_8298_5487# 0.0047f
C2465 net9 net2 0.0285f
C2466 clknet_2_3__leaf_clk a_12153_8757# 0.00203f
C2467 net41 a_3339_2767# 5.27e-20
C2468 _122_ a_10864_7387# 0.00922f
C2469 _115_ _057_ 1.61e-20
C2470 _056_ a_13307_1707# 8.32e-21
C2471 net44 a_4775_6031# 0.153f
C2472 a_1497_8725# a_1387_8751# 0.0977f
C2473 net41 a_995_3530# 0.0639f
C2474 a_6173_7119# a_6428_7119# 0.0642f
C2475 a_8022_7119# a_10586_7371# 4.44e-19
C2476 a_3891_4943# a_4175_4943# 8.61e-19
C2477 a_9719_1473# net11 9.67e-20
C2478 a_4471_4007# VPWR 0.176f
C2479 net20 a_6743_10933# 0.0134f
C2480 clknet_2_3__leaf_clk a_11023_5108# 1.9e-19
C2481 net44 a_6633_9845# 0.0334f
C2482 net31 net37 0.249f
C2483 _098_ a_5536_4399# 4.91e-19
C2484 a_579_12021# mask\[7\] 1.54e-19
C2485 cal_count\[1\] _134_ 2.26e-21
C2486 _011_ a_1660_12393# 1.26e-19
C2487 net47 cal_count\[0\] 0.268f
C2488 cal_count\[0\] a_14377_9545# 0.0075f
C2489 cal_itt\[0\] a_7001_7669# 4.7e-21
C2490 _063_ a_10864_7387# 0.00209f
C2491 _110_ a_13881_1653# 4.04e-19
C2492 net40 a_13512_4943# 6.16e-19
C2493 a_8949_6031# _106_ 1.13e-19
C2494 _092_ a_8389_5193# 1.19e-19
C2495 _064_ _058_ 0.12f
C2496 _059_ _100_ 0.0368f
C2497 clknet_2_2__leaf_clk a_11951_2601# 2.28e-19
C2498 a_12870_2589# VPWR 2.5e-19
C2499 a_5423_9011# VPWR 0.475f
C2500 net14 net1 0.0299f
C2501 a_9460_6807# net30 8.82e-21
C2502 a_561_6031# a_561_4405# 2.34e-19
C2503 mask\[7\] a_2869_10927# 0.0111f
C2504 net40 a_14377_7983# 0.00447f
C2505 net27 a_6099_10633# 4e-20
C2506 a_1229_8457# VPWR 0.00533f
C2507 a_4775_6031# en_co_clk 0.003f
C2508 _040_ a_5535_8181# 3.4e-19
C2509 clknet_2_0__leaf_clk a_4349_8449# 4.81e-19
C2510 _045_ a_3597_12021# 1.48e-20
C2511 trim_mask\[4\] a_8491_2229# 1.35e-21
C2512 a_5699_9269# a_5423_9011# 0.00472f
C2513 _063_ a_9503_4399# 3.05e-19
C2514 a_4970_4399# VPWR 0.00569f
C2515 clknet_2_3__leaf_clk a_8307_6575# 3.8e-20
C2516 a_8083_8181# clknet_0_clk 2.29e-19
C2517 _136_ a_10781_5487# 0.0131f
C2518 net44 a_3411_7485# 2.61e-20
C2519 clknet_2_3__leaf_clk a_11268_9295# 2.82e-19
C2520 _113_ a_11509_3317# 8.33e-20
C2521 net5 a_14379_6397# 1.94e-19
C2522 mask\[4\] a_3868_10217# 1.5e-19
C2523 _104_ a_10699_3311# 0.242f
C2524 a_2659_2601# a_2564_2589# 0.0498f
C2525 a_2877_2197# a_2755_2601# 3.16e-19
C2526 a_2143_2229# a_3333_2601# 2.56e-19
C2527 cal_count\[3\] _135_ 0.00333f
C2528 a_11955_3689# VPWR 3.07e-19
C2529 VPWR clkc 0.367f
C2530 a_7001_7669# a_7569_7637# 0.172f
C2531 a_6835_7669# a_7351_8041# 0.106f
C2532 net45 _053_ 5.85e-20
C2533 _108_ a_15023_2223# 6.33e-19
C2534 _134_ _108_ 3.3e-20
C2535 _101_ a_1844_9129# 0.00106f
C2536 a_1867_3317# a_2033_3317# 0.904f
C2537 _117_ VPWR 0.231f
C2538 _053_ _058_ 0.00145f
C2539 a_9677_8457# VPWR 0.00273f
C2540 net54 _104_ 0.00148f
C2541 net30 _107_ 0.239f
C2542 net13 a_4349_8449# 0.00446f
C2543 a_12436_9129# net2 1.28e-19
C2544 a_9595_1679# a_10207_1679# 4.78e-19
C2545 net52 a_2857_7637# 0.241f
C2546 a_11141_6031# a_11491_6031# 0.206f
C2547 trim_mask\[1\] a_13625_3317# 0.00414f
C2548 a_2857_5461# a_3057_4719# 1.08e-19
C2549 mask\[0\] clknet_0_clk 0.00866f
C2550 _030_ a_14540_3689# 1.61e-19
C2551 a_13459_3317# _055_ 3.54e-19
C2552 a_4995_7119# a_4883_6397# 5.72e-20
C2553 net12 a_7569_7637# 7.74e-20
C2554 a_11987_8757# _041_ 0.0381f
C2555 _036_ a_13562_8751# 1.37e-20
C2556 a_3748_6281# _094_ 0.0449f
C2557 a_1125_7663# VPWR 0.241f
C2558 net46 a_12533_3689# 0.00112f
C2559 a_455_8181# _080_ 8.56e-20
C2560 _108_ a_13975_3689# 0.0112f
C2561 a_6888_10205# a_7079_10217# 4.61e-19
C2562 a_2489_7983# VPWR 6.3e-19
C2563 _049_ net30 0.0182f
C2564 clknet_2_1__leaf_clk a_4043_7093# 0.0013f
C2565 _066_ a_11425_5487# 0.0125f
C2566 a_1644_12533# ctlp[1] 1.47e-19
C2567 calibrate a_6566_5193# 0.024f
C2568 net46 a_12323_4703# 0.294f
C2569 net3 net41 0.00983f
C2570 a_3667_3829# a_3224_2601# 8.6e-20
C2571 a_5363_12559# VPWR 0.455f
C2572 _095_ calibrate 0.00101f
C2573 trim_mask\[1\] a_8583_3317# 4.07e-20
C2574 a_10188_4105# _033_ 3.76e-22
C2575 net14 result[6] 4.91e-20
C2576 net13 a_3511_11471# 3.31e-21
C2577 a_6181_10633# _020_ 0.00169f
C2578 a_1493_11721# a_579_10933# 2.65e-20
C2579 _062_ _106_ 0.0208f
C2580 a_2383_3689# a_2645_3677# 0.00171f
C2581 a_2601_3285# a_3057_3689# 4.2e-19
C2582 net16 _110_ 0.0575f
C2583 a_1867_3317# a_2491_3311# 9.73e-19
C2584 _078_ _042_ 0.0121f
C2585 a_7715_3285# a_7223_2465# 1.17e-19
C2586 a_7010_3311# a_7184_2339# 5.77e-21
C2587 net43 a_1679_10633# 6.99e-20
C2588 _090_ a_4091_4943# 1.09e-19
C2589 trim_val\[3\] a_10872_1455# 3.91e-19
C2590 a_3840_8867# a_4036_8207# 9.86e-19
C2591 _108_ a_13915_4399# 0.0687f
C2592 net2 _062_ 1.3e-20
C2593 _074_ a_855_4105# 0.096f
C2594 cal_itt\[1\] a_11059_7356# 1.58e-19
C2595 a_4871_8181# VPWR 0.366f
C2596 a_10005_6031# _092_ 0.368f
C2597 _081_ net45 6.44e-20
C2598 net12 trim_mask\[0\] 5.52e-21
C2599 clknet_2_1__leaf_clk a_1660_12393# 4.87e-19
C2600 a_745_12021# a_1313_11989# 0.186f
C2601 _076_ VPWR 1.44f
C2602 _014_ a_2033_3317# 0.0222f
C2603 _101_ a_5633_9295# 2.21e-19
C2604 net18 _116_ 0.0016f
C2605 net19 a_8912_2589# 0.00495f
C2606 a_4775_6031# _059_ 4.42e-20
C2607 a_6983_10217# a_7079_10217# 0.0138f
C2608 _055_ trim[2] 1.84e-20
C2609 net12 _075_ 0.057f
C2610 a_8298_5487# _119_ 2.64e-20
C2611 _104_ _027_ 0.146f
C2612 a_2787_7119# a_3748_6281# 7.58e-19
C2613 a_2828_12131# ctlp[1] 3.63e-19
C2614 clknet_2_1__leaf_clk a_3565_10205# 4.26e-19
C2615 net47 a_13919_8751# 4.17e-20
C2616 _051_ a_7758_4759# 1.93e-20
C2617 net19 a_8673_10625# 0.00947f
C2618 mask\[0\] a_2476_6281# 0.00141f
C2619 net52 a_2953_9845# 0.0131f
C2620 _058_ a_14335_4020# 0.005f
C2621 net50 a_10207_1679# 3.14e-19
C2622 a_8583_3317# a_8749_3317# 0.735f
C2623 _092_ _087_ 0.0261f
C2624 _096_ _097_ 0.0117f
C2625 a_7019_4407# _104_ 1.3e-19
C2626 _033_ trim_mask\[3\] 4.38e-20
C2627 _074_ a_763_8757# 0.0189f
C2628 a_579_10933# VPWR 0.466f
C2629 a_5340_6031# _075_ 0.00231f
C2630 _119_ a_10111_1679# 1.05e-20
C2631 a_11343_3317# a_12533_3689# 2.56e-19
C2632 _025_ a_12121_3677# 1.11e-19
C2633 net22 a_1651_6005# 0.136f
C2634 _092_ _099_ 0.341f
C2635 a_13142_8359# a_13356_8457# 0.013f
C2636 _028_ a_7310_2223# 0.0322f
C2637 net55 _088_ 0.044f
C2638 _101_ _017_ 8.39e-20
C2639 a_929_8757# net24 0.551f
C2640 a_8657_2229# a_9007_2601# 0.22f
C2641 net46 a_14379_6397# 3.5e-19
C2642 a_10975_6031# a_11396_6031# 0.0866f
C2643 clknet_0_clk net54 4.49e-20
C2644 a_3597_10933# _042_ 2.83e-19
C2645 a_7201_9813# a_7548_10217# 0.0512f
C2646 trim_val\[0\] _047_ 0.039f
C2647 _045_ mask\[5\] 3.91e-21
C2648 a_561_6031# result[0] 0.001f
C2649 a_395_6031# sample 0.00361f
C2650 a_5496_12131# a_6375_12021# 2.1e-21
C2651 _001_ a_11059_7356# 0.0119f
C2652 net15 mask\[2\] 0.291f
C2653 net13 a_5055_9295# 0.00121f
C2654 net55 a_7262_5461# 8.85e-21
C2655 net47 a_9459_7895# 1.02e-19
C2656 a_763_8757# a_1279_9129# 0.115f
C2657 _014_ a_2491_3311# 0.00325f
C2658 _074_ net26 1.16f
C2659 a_11583_4777# _025_ 9.83e-21
C2660 net53 a_8105_10383# 0.00126f
C2661 a_11583_4777# _026_ 4.33e-20
C2662 net44 net47 6.3e-19
C2663 state\[2\] _107_ 0.0225f
C2664 _078_ a_1476_6031# 0.0138f
C2665 a_15023_9839# VPWR 0.457f
C2666 a_5363_12559# net27 6.42e-21
C2667 net23 _039_ 1.96e-19
C2668 net43 _065_ 0.0751f
C2669 a_395_2767# cal 0.00459f
C2670 a_9296_9295# _041_ 4.03e-20
C2671 mask\[1\] a_1129_7361# 5.96e-19
C2672 net2 a_13470_7663# 4.96e-19
C2673 _038_ net46 0.0265f
C2674 a_455_3571# cal 0.0251f
C2675 net9 a_12249_7663# 0.003f
C2676 VPWR ctlp[6] 0.774f
C2677 _078_ a_6909_10933# 1.08e-20
C2678 _035_ a_10747_8970# 0.12f
C2679 a_3933_2767# clk 0.00238f
C2680 net55 a_6519_4631# 0.048f
C2681 a_10239_9295# _124_ 2.26e-20
C2682 net43 net23 0.0439f
C2683 a_11067_4405# a_12257_4777# 2.56e-19
C2684 _093_ a_855_4105# 0.205f
C2685 a_1095_12393# a_745_10933# 2.28e-19
C2686 a_4995_7119# a_4993_6273# 4.89e-20
C2687 a_5363_7369# a_4425_6031# 2.43e-20
C2688 net53 a_6261_11247# 0.00193f
C2689 _049_ state\[2\] 0.00628f
C2690 _029_ a_13512_4943# 0.158f
C2691 net16 a_14564_6397# 0.00604f
C2692 net44 a_7355_11305# 0.00198f
C2693 mask\[2\] a_4030_9839# 6e-20
C2694 trim_mask\[0\] a_13703_4943# 0.00131f
C2695 _050_ a_7010_3311# 0.0243f
C2696 a_3852_12381# a_4043_12393# 4.61e-19
C2697 state\[2\] a_5699_1653# 0.0638f
C2698 net19 a_8767_591# 2.97e-19
C2699 trim_val\[2\] trim[2] 0.00257f
C2700 a_4131_8207# a_4036_8207# 0.0498f
C2701 net47 en_co_clk 1.35e-19
C2702 a_4349_8449# a_4239_8573# 0.0977f
C2703 _104_ _117_ 8.64e-20
C2704 net52 a_1585_10217# 9.61e-21
C2705 _049_ state\[0\] 4.22e-19
C2706 _069_ _053_ 0.00188f
C2707 cal_count\[2\] a_12430_7663# 6.34e-21
C2708 net15 a_2143_2229# 0.0147f
C2709 clknet_2_3__leaf_clk VPWR 3.33f
C2710 a_3817_4697# a_3667_3829# 0.00601f
C2711 clknet_2_2__leaf_clk a_9369_4105# 6e-20
C2712 _072_ a_6741_7361# 1.19e-19
C2713 _094_ a_4308_4917# 3.55e-19
C2714 net15 _085_ 0.46f
C2715 a_3597_12021# _078_ 8.12e-19
C2716 _110_ _027_ 0.00725f
C2717 _053_ a_8022_7119# 8.73e-19
C2718 net41 valid 0.0214f
C2719 net16 a_14467_8751# 0.00195f
C2720 a_911_10217# net25 8.59e-19
C2721 a_1651_10143# a_1476_10217# 0.234f
C2722 _073_ _050_ 3.44e-20
C2723 _090_ a_3751_4765# 0.00553f
C2724 clknet_2_1__leaf_clk a_7939_10383# 0.243f
C2725 clknet_2_3__leaf_clk a_12218_6397# 8.2e-20
C2726 a_395_9845# VPWR 0.488f
C2727 a_9871_10383# cal_itt\[0\] 4.47e-22
C2728 _052_ a_7010_3311# 0.22f
C2729 a_4864_9295# a_5055_9295# 4.61e-19
C2730 net16 a_13091_4943# 0.0122f
C2731 net27 a_579_10933# 0.00215f
C2732 net14 a_911_10217# 0.00416f
C2733 _062_ _054_ 1.53e-22
C2734 mask\[3\] a_4443_9295# 0.309f
C2735 clknet_2_0__leaf_clk a_3667_3829# 4.38e-20
C2736 a_8820_6005# en_co_clk 0.0268f
C2737 clknet_0_clk a_7019_4407# 1.68e-20
C2738 a_4259_6031# _092_ 0.00189f
C2739 a_10752_565# net10 0.184f
C2740 _098_ a_7010_3311# 2.07e-21
C2741 net45 a_7379_2197# 0.155f
C2742 _108_ trim_val\[1\] 0.139f
C2743 net41 a_5537_4105# 0.0113f
C2744 a_3868_7119# a_5363_7369# 4.17e-20
C2745 net32 a_14715_3615# 0.00146f
C2746 _039_ a_1019_6397# 6.5e-19
C2747 _114_ a_14099_1929# 2.49e-19
C2748 net52 mask\[3\] 0.261f
C2749 net43 _016_ 8.35e-19
C2750 net30 sample 0.017f
C2751 net55 a_8745_4943# 2.93e-19
C2752 net24 clknet_2_0__leaf_clk 1.23e-19
C2753 _064_ a_8657_2229# 2.68e-21
C2754 net30 trim_mask\[4\] 1.57e-19
C2755 _118_ a_9802_4007# 0.0492f
C2756 _107_ _100_ 0.0129f
C2757 cal_itt\[0\] _091_ 0.134f
C2758 a_561_4405# a_455_3571# 5.23e-20
C2759 _070_ a_8301_8207# 0.0486f
C2760 _101_ a_3868_7119# 7.56e-20
C2761 trim_mask\[0\] a_13459_3317# 4.34e-20
C2762 _065_ a_2857_7637# 6.09e-19
C2763 a_2564_2589# VPWR 0.0794f
C2764 _095_ _015_ 1.44e-20
C2765 net13 a_3667_3829# 4.35e-19
C2766 a_10055_2767# _116_ 9.48e-21
C2767 _108_ _118_ 0.445f
C2768 _105_ a_9125_4943# 0.0096f
C2769 cal_count\[3\] a_10781_5487# 0.0172f
C2770 a_7001_7669# a_7723_6807# 6.15e-20
C2771 a_3597_12021# a_3597_10933# 1.55e-20
C2772 a_395_7119# a_1585_7119# 2.56e-19
C2773 net46 ctln[4] 1.77e-19
C2774 net43 a_4696_8207# 5.92e-19
C2775 a_1129_4373# cal 6.15e-19
C2776 _050_ a_3365_4943# 8.07e-19
C2777 net23 a_2857_7637# 0.00115f
C2778 a_4512_12393# a_5496_12131# 2.65e-19
C2779 a_11369_7119# _136_ 2.96e-19
C2780 a_9747_2527# a_9761_1679# 0.00203f
C2781 _070_ a_9621_8029# 2.89e-20
C2782 net9 a_12756_9117# 2.99e-19
C2783 _007_ result[2] 4.52e-19
C2784 _049_ _100_ 0.0119f
C2785 a_10864_7387# a_11622_7485# 0.0604f
C2786 a_10903_7261# a_11204_7485# 9.73e-19
C2787 net43 _067_ 0.00265f
C2788 _099_ a_6737_4719# 4.21e-19
C2789 mask\[7\] _101_ 0.132f
C2790 net13 net24 2.64e-19
C2791 trim_mask\[0\] _109_ 0.103f
C2792 cal_itt\[2\] net55 1.23e-20
C2793 a_10975_4105# a_11509_3317# 3.43e-19
C2794 net5 en_co_clk 6.94e-19
C2795 _060_ a_5625_4943# 1.78e-19
C2796 _084_ net13 5.3e-20
C2797 clknet_2_0__leaf_clk a_4883_6397# 1.08e-20
C2798 net12 _042_ 0.00452f
C2799 net45 a_3530_4438# 8.89e-20
C2800 _087_ a_5536_4399# 0.00945f
C2801 a_11425_5487# _058_ 2.5e-19
C2802 net12 a_7723_6807# 2.86e-19
C2803 a_14715_3615# VPWR 0.359f
C2804 _110_ _117_ 0.0389f
C2805 _078_ a_4959_9295# 7.59e-21
C2806 _053_ a_8657_2229# 1.33e-19
C2807 net54 net41 0.407f
C2808 a_9463_8725# _041_ 0.0425f
C2809 net12 a_7210_5807# 4.34e-22
C2810 net4 a_7223_2465# 1.01e-19
C2811 _123_ a_10903_7261# 1.94e-19
C2812 clknet_2_2__leaf_clk a_8307_4719# 4.21e-20
C2813 a_11116_8983# a_11059_7356# 3.01e-20
C2814 net43 _023_ 0.00545f
C2815 _124_ a_11545_9049# 1.38e-20
C2816 net47 cal_count\[2\] 0.00129f
C2817 a_10747_8970# a_11987_8757# 2.52e-21
C2818 _013_ a_2601_3285# 3.21e-20
C2819 _099_ a_5536_4399# 0.0441f
C2820 trim_val\[2\] a_15023_1135# 0.0717f
C2821 _058_ a_10781_3631# 1.22e-19
C2822 _004_ a_1476_6031# 5.47e-21
C2823 net1 VPWR 0.177f
C2824 net14 a_2143_2229# 8.86e-19
C2825 net9 a_12599_3615# 0.0067f
C2826 a_2857_5461# a_3891_4943# 0.00268f
C2827 net15 a_4443_1679# 7.97e-21
C2828 net47 a_10688_9295# 0.254f
C2829 _075_ a_5726_5807# 0.00673f
C2830 _094_ _090_ 2.67e-20
C2831 a_10405_9295# a_10798_9295# 0.00127f
C2832 _072_ a_9459_7895# 8.68e-20
C2833 net13 a_4883_6397# 0.00431f
C2834 a_1644_12533# net15 1.16e-20
C2835 net29 a_3116_12533# 8.41e-19
C2836 mask\[7\] _086_ 0.0853f
C2837 a_13881_2741# a_14099_3017# 0.0821f
C2838 net4 a_9099_3689# 0.0072f
C2839 a_1660_11305# a_1822_10927# 0.00645f
C2840 net47 a_8992_9955# 0.00372f
C2841 _136_ a_13233_4737# 1.14e-19
C2842 a_13512_4943# trim_mask\[1\] 1.91e-20
C2843 a_11801_4373# a_11583_4777# 0.21f
C2844 a_11233_4405# a_12323_4703# 0.0424f
C2845 _064_ a_10569_1109# 1.27e-19
C2846 a_2857_7637# _016_ 0.0198f
C2847 a_14335_4020# _113_ 3.36e-21
C2848 net44 _072_ 0.477f
C2849 a_561_4405# _099_ 7.61e-21
C2850 clknet_2_0__leaf_clk a_1129_6273# 2.62e-19
C2851 net43 a_816_10205# 5.45e-19
C2852 _092_ a_7393_5193# 0.00184f
C2853 a_5691_7637# _049_ 4.88e-19
C2854 _091_ trim_mask\[0\] 7.39e-20
C2855 _055_ trim[1] 0.00585f
C2856 net44 _068_ 0.0278f
C2857 cal_count\[3\] _098_ 1.22e-20
C2858 a_5363_591# a_6927_591# 5.8e-21
C2859 _108_ a_10137_4943# 3.51e-19
C2860 _078_ mask\[5\] 0.281f
C2861 mask\[7\] _102_ 0.206f
C2862 a_5177_1921# ctln[7] 8.2e-20
C2863 _118_ _107_ 0.0151f
C2864 a_561_4405# a_1129_4373# 0.181f
C2865 a_4687_11231# a_4443_9295# 1.42e-20
C2866 _042_ a_1651_10143# 2.13e-19
C2867 _079_ a_1137_5487# 1.66e-20
C2868 net45 a_5221_1679# 0.00316f
C2869 net28 a_6541_12021# 1.5e-20
C2870 net44 a_4443_9295# 0.301f
C2871 a_8455_10383# clknet_2_3__leaf_clk 2.78e-20
C2872 _041_ a_11258_9117# 0.0019f
C2873 a_12436_9129# a_12756_9117# 0.00184f
C2874 a_12612_8725# a_13016_9117# 3.94e-19
C2875 state\[2\] trim_mask\[4\] 0.168f
C2876 net41 a_2645_3677# 0.00208f
C2877 net2 a_14788_7369# 0.177f
C2878 clknet_2_3__leaf_clk _104_ 1.02e-19
C2879 net26 _083_ 0.256f
C2880 net15 a_2828_12131# 8.23e-19
C2881 net18 a_11601_2229# 5.13e-20
C2882 a_5515_6005# a_5363_4719# 1.43e-21
C2883 clknet_2_0__leaf_clk a_4677_7882# 3.11e-19
C2884 a_11057_4105# a_10699_3311# 8.48e-20
C2885 net16 a_14249_8725# 0.00959f
C2886 a_1679_10633# mask\[3\] 1.23e-21
C2887 _072_ clk 0.207f
C2888 net18 net17 0.0821f
C2889 net44 net52 0.0125f
C2890 _072_ en_co_clk 1.19e-19
C2891 net12 a_5177_1921# 9.81e-19
C2892 net55 a_5081_4943# 0.0563f
C2893 _096_ a_4709_2773# 8.02e-19
C2894 a_3781_8207# net45 4.53e-20
C2895 net12 a_6909_10933# 3.78e-20
C2896 _065_ _038_ 0.243f
C2897 a_12520_7637# a_13092_8029# 1.57e-19
C2898 net47 a_9374_10383# 0.00223f
C2899 a_1830_6031# VPWR 2.57e-19
C2900 net23 a_1638_7485# 5.16e-20
C2901 _068_ clk 2.05e-20
C2902 net24 a_561_7119# 5.52e-22
C2903 a_8083_8181# _001_ 3.4e-20
C2904 trim_val\[0\] net49 4.74e-20
C2905 a_14099_1929# VPWR 0.276f
C2906 _068_ en_co_clk 0.0292f
C2907 net45 a_395_4405# 0.298f
C2908 _075_ _089_ 5.41e-22
C2909 net11 ctln[5] 0.0102f
C2910 a_4471_4007# net41 2.57e-19
C2911 state\[1\] a_4617_4105# 9.96e-21
C2912 _076_ a_6198_8207# 0.00129f
C2913 a_14564_6397# clkc 7.77e-19
C2914 mask\[7\] _022_ 0.00132f
C2915 clknet_2_1__leaf_clk a_6056_8359# 0.00533f
C2916 en_co_clk a_15023_6031# 0.00106f
C2917 _096_ a_4308_4917# 4.47e-19
C2918 a_763_8757# a_911_7119# 3.47e-19
C2919 _049_ a_4775_6031# 0.0111f
C2920 a_395_591# clk 0.00296f
C2921 _105_ a_8389_5193# 0.00736f
C2922 _047_ net32 0.147f
C2923 _068_ a_8386_8457# 4e-19
C2924 a_9761_1679# a_10676_1679# 0.125f
C2925 a_4425_6031# a_4498_4373# 3.63e-22
C2926 trim_mask\[1\] a_11859_3689# 0.03f
C2927 a_13825_1109# a_13703_1513# 3.16e-19
C2928 net18 a_12061_7669# 1.81e-20
C2929 a_13607_1513# a_13512_1501# 0.0498f
C2930 calibrate _015_ 0.0209f
C2931 a_8827_9295# VPWR 4.33e-19
C2932 a_13459_3317# _030_ 0.381f
C2933 net13 a_4677_7882# 0.00464f
C2934 mask\[5\] a_3597_10933# 3.3e-20
C2935 a_4167_11471# a_4165_10901# 0.00118f
C2936 VPWR result[6] 0.49f
C2937 net15 _120_ 0.0591f
C2938 a_13257_1141# trim[3] 1.78e-19
C2939 a_2143_2229# a_2659_2601# 0.115f
C2940 a_2309_2229# a_2877_2197# 0.181f
C2941 net22 a_1549_6794# 0.0015f
C2942 a_13607_4943# trim[4] 7.31e-20
C2943 mask\[4\] a_7657_10217# 8.37e-19
C2944 clknet_2_1__leaf_clk a_1045_9545# 8.92e-19
C2945 net47 cal_count\[1\] 4.73e-19
C2946 _067_ a_8270_8029# 1.46e-21
C2947 net4 trim_val\[4\] 0.0023f
C2948 _060_ _103_ 8.17e-21
C2949 clknet_2_2__leaf_clk a_12533_3689# 1.2e-21
C2950 clknet_2_0__leaf_clk a_4993_6273# 6.55e-19
C2951 a_745_10933# a_1461_10357# 2.09e-19
C2952 clknet_2_3__leaf_clk a_8381_9295# 0.588f
C2953 net13 a_4801_10159# 5.63e-19
C2954 net46 a_9084_4515# 2.34e-20
C2955 _126_ a_14733_9545# 7.6e-19
C2956 a_3868_10217# a_3781_8207# 4.8e-21
C2957 net55 a_7715_3285# 1.95e-21
C2958 a_7109_11989# a_7565_12393# 4.2e-19
C2959 net44 a_7153_12381# 0.00316f
C2960 clknet_2_1__leaf_clk a_1095_11305# 6.62e-19
C2961 a_10137_4943# _107_ 9.64e-19
C2962 clknet_2_2__leaf_clk a_12323_4703# 0.00475f
C2963 _070_ _063_ 0.0225f
C2964 _078_ _039_ 0.2f
C2965 trim_mask\[0\] a_14655_4399# 2.95e-19
C2966 a_5535_8181# _077_ 0.326f
C2967 _108_ a_12502_4765# 4.2e-20
C2968 a_3339_2767# a_3224_2601# 6.5e-20
C2969 a_3411_7485# _049_ 2.26e-19
C2970 mask\[3\] _065_ 2.22e-20
C2971 net21 a_6541_12021# 2.49e-21
C2972 net4 a_9823_6941# 4.03e-19
C2973 a_2787_9845# a_2815_9447# 0.00133f
C2974 net28 a_3116_12533# 2.54e-19
C2975 net14 a_1644_12533# 0.0211f
C2976 _072_ a_8091_7967# 0.0404f
C2977 a_8083_8181# a_7916_8041# 6.84e-19
C2978 _065_ a_6741_7361# 1.3e-21
C2979 a_1099_12533# net29 0.00225f
C2980 net15 a_4609_9295# 1.58e-21
C2981 net43 _078_ 2.59f
C2982 state\[0\] a_3123_3615# 0.062f
C2983 _047_ VPWR 0.374f
C2984 net14 a_1476_4777# 0.00637f
C2985 a_7223_2465# a_7689_2589# 0.00188f
C2986 _074_ a_1279_9129# 0.00391f
C2987 net12 a_5633_1679# 9.9e-20
C2988 a_7310_2223# a_7181_2589# 4.2e-19
C2989 a_6835_7669# VPWR 0.48f
C2990 _092_ _097_ 0.0631f
C2991 mask\[3\] net23 2.04e-20
C2992 _050_ _119_ 2.53e-20
C2993 net13 a_4993_6273# 0.00672f
C2994 clknet_2_3__leaf_clk _110_ 1.07e-20
C2995 _048_ trim_mask\[0\] 0.124f
C2996 a_15159_9269# a_15023_8751# 0.0126f
C2997 net47 a_12612_8725# 0.158f
C2998 net1 a_2383_3689# 1.71e-20
C2999 _068_ a_8091_7967# 6.01e-19
C3000 clknet_2_3__leaf_clk clknet_0_clk 0.00541f
C3001 net37 trimb[1] 0.0164f
C3002 _116_ VPWR 0.299f
C3003 a_3597_12021# a_3852_12381# 0.0612f
C3004 a_3431_12021# a_4043_12393# 3.82e-19
C3005 net33 a_14972_5193# 0.00612f
C3006 clknet_2_0__leaf_clk a_3208_7119# 0.0139f
C3007 net43 a_2869_11247# 3.35e-21
C3008 _075_ _048_ 0.0203f
C3009 a_5524_9295# a_5691_7637# 2.12e-19
C3010 _064_ a_10975_4105# 0.0912f
C3011 _084_ a_7631_12319# 1.03e-21
C3012 a_14335_7895# a_14377_7983# 0.0175f
C3013 a_6090_10159# VPWR 5.72e-19
C3014 a_561_7119# a_1129_6273# 6.96e-20
C3015 state\[1\] a_3578_2589# 6.42e-19
C3016 _052_ _119_ 2.32e-21
C3017 a_5915_11721# VPWR 0.254f
C3018 clknet_2_1__leaf_clk a_4674_12015# 3.05e-19
C3019 a_395_591# ctln[0] 3.49e-19
C3020 net51 a_7447_8041# 3.68e-19
C3021 _050_ a_6566_5193# 7.3e-19
C3022 _067_ _038_ 3.04e-20
C3023 a_12424_3689# a_12516_2601# 4.15e-21
C3024 clknet_2_3__leaf_clk a_10699_5487# 0.0472f
C3025 a_12664_8029# VPWR 3.86e-19
C3026 a_4801_9839# a_4443_9295# 2.38e-19
C3027 _095_ _050_ 0.501f
C3028 a_5166_5193# a_5081_4943# 8.13e-19
C3029 net55 _093_ 0.0155f
C3030 net19 _027_ 0.0148f
C3031 _008_ a_6633_9845# 0.301f
C3032 net27 result[6] 9.45e-21
C3033 net9 a_13607_1513# 4.91e-19
C3034 a_6467_9845# a_7201_9813# 0.0701f
C3035 a_14347_4917# a_14526_4943# 0.0074f
C3036 a_14172_4943# a_14281_4943# 0.00742f
C3037 net17 a_12153_8757# 1.07e-20
C3038 a_15023_2223# _056_ 0.171f
C3039 a_9871_10383# _042_ 0.0295f
C3040 _103_ a_7939_3855# 1.75e-19
C3041 a_11067_4405# a_10699_3311# 0.00109f
C3042 _012_ sample 3.98e-19
C3043 net55 a_5166_5193# 0.00112f
C3044 a_5515_6005# VPWR 0.36f
C3045 clknet_2_0__leaf_clk result[1] 0.0172f
C3046 net43 a_3597_10933# 0.044f
C3047 _096_ _090_ 0.372f
C3048 mask\[3\] a_2225_7663# 2.59e-20
C3049 a_6566_5193# _052_ 2.72e-19
C3050 _074_ _093_ 3.37e-19
C3051 a_7201_9813# VPWR 0.215f
C3052 net47 a_11436_9295# 0.00173f
C3053 a_8215_9295# _041_ 2.19e-19
C3054 net2 _037_ 1.05e-19
C3055 _033_ _028_ 7.86e-20
C3056 _096_ a_3847_4438# 0.00526f
C3057 trim_mask\[3\] a_10543_2455# 0.172f
C3058 _038_ clknet_2_2__leaf_clk 1.8e-20
C3059 _095_ _098_ 2.5e-20
C3060 a_12153_8757# a_12061_7669# 4.41e-21
C3061 calibrate a_7184_2339# 1.61e-19
C3062 cal_count\[3\] a_8389_5193# 2.87e-19
C3063 mask\[2\] _019_ 0.3f
C3064 a_10543_2455# a_10689_2543# 0.0134f
C3065 a_11067_3017# a_10676_1679# 3.02e-20
C3066 a_9225_2197# a_9734_2223# 2.6e-19
C3067 net4 cal_itt\[2\] 1.64e-21
C3068 _081_ a_2092_8457# 0.0504f
C3069 cal_count\[0\] a_14552_9071# 0.00958f
C3070 _078_ a_2857_7637# 0.0012f
C3071 _122_ a_11098_6691# 4.96e-19
C3072 _108_ a_14686_2339# 5.09e-19
C3073 net2 a_12231_6005# 0.00641f
C3074 a_911_10217# VPWR 0.197f
C3075 trim_mask\[0\] trim[1] 6.55e-19
C3076 net13 a_4222_10205# 2.3e-19
C3077 a_9463_8725# a_10747_8970# 1.92e-20
C3078 a_6056_8359# a_6007_7119# 1.43e-20
C3079 _118_ trim_mask\[4\] 0.0192f
C3080 net28 a_4043_12393# 0.00432f
C3081 mask\[5\] net12 0.318f
C3082 _126_ a_15159_9269# 0.0944f
C3083 a_14983_9269# _125_ 0.0677f
C3084 net3 a_3224_2601# 1.46e-20
C3085 _076_ a_6523_7119# 0.00105f
C3086 a_1585_7119# VPWR 5.6e-20
C3087 clknet_2_3__leaf_clk a_14564_6397# 0.00159f
C3088 a_9182_10749# VPWR 5.68e-19
C3089 a_9003_3829# a_9369_3855# 0.0245f
C3090 a_4815_3031# a_4959_1679# 4.71e-20
C3091 net27 a_5915_11721# 0.00977f
C3092 a_13625_3317# a_14071_3689# 2.28e-19
C3093 net28 a_1099_12533# 0.0464f
C3094 net2 a_8301_8207# 0.0404f
C3095 _035_ a_12341_8751# 9.09e-21
C3096 net15 a_1867_3317# 2.99e-20
C3097 a_14334_5309# VPWR 5.43e-19
C3098 _065_ a_9459_7895# 2.44e-19
C3099 a_12169_2197# a_11951_2601# 0.21f
C3100 a_11601_2229# a_12691_2527# 0.0424f
C3101 a_11435_2229# a_12516_2601# 0.102f
C3102 net22 a_1007_6031# 9.4e-19
C3103 net46 a_12410_6031# 0.00225f
C3104 net19 _117_ 5.71e-21
C3105 net44 _065_ 0.752f
C3106 net47 a_12900_7663# 0.217f
C3107 _058_ a_13625_3317# 0.00218f
C3108 _084_ a_5915_10927# 4.16e-19
C3109 a_7527_4631# clk 5.87e-19
C3110 a_8820_6005# _107_ 9.99e-19
C3111 net3 a_4863_4917# 0.0348f
C3112 _090_ a_5455_4943# 8.61e-20
C3113 _108_ a_14347_1439# 4.38e-19
C3114 mask\[7\] _046_ 0.0168f
C3115 net16 net37 2.55e-20
C3116 a_12824_7663# VPWR 0.00403f
C3117 clknet_2_0__leaf_clk a_3339_2767# 4.69e-20
C3118 _051_ a_7800_4631# 0.122f
C3119 a_7824_11305# a_8105_10383# 7.71e-20
C3120 _039_ _004_ 1.08e-19
C3121 clknet_2_0__leaf_clk a_995_3530# 6.32e-20
C3122 net45 a_2283_4020# 0.0324f
C3123 _074_ a_448_7637# 0.00436f
C3124 net9 a_11709_6273# 7.52e-19
C3125 mask\[0\] a_4995_7119# 4.45e-19
C3126 mask\[2\] VPWR 0.609f
C3127 a_13184_9117# VPWR 8.97e-20
C3128 a_13881_2741# trim[0] 1.8e-19
C3129 state\[1\] clk 0.00418f
C3130 en_co_clk state\[1\] 6.36e-19
C3131 net26 _000_ 5.23e-20
C3132 a_395_6031# a_1493_5487# 7.96e-20
C3133 _062_ net3 0.0875f
C3134 _078_ a_2953_9845# 3.45e-20
C3135 _058_ a_12310_4399# 1.09e-19
C3136 a_15083_4659# _109_ 4.83e-20
C3137 a_13697_4373# a_14000_4719# 0.00138f
C3138 a_15023_10927# trimb[2] 0.00188f
C3139 _063_ net50 2.42e-20
C3140 mask\[2\] a_5699_9269# 8.98e-21
C3141 _048_ a_8307_4943# 0.101f
C3142 net16 a_13193_6031# 4.35e-20
C3143 _065_ clk 2.07e-20
C3144 _065_ en_co_clk 0.198f
C3145 _134_ _061_ 0.0033f
C3146 a_7259_11305# a_7355_11305# 0.0138f
C3147 a_6909_10933# a_5997_10927# 4.14e-19
C3148 a_8949_9537# a_9458_9661# 2.6e-19
C3149 a_8381_9295# a_8827_9295# 2.28e-19
C3150 net15 a_3302_3677# 2.71e-19
C3151 net18 _025_ 0.00262f
C3152 _104_ _116_ 1.8e-20
C3153 net43 a_7001_7669# 0.639f
C3154 _099_ a_3148_4399# 0.00421f
C3155 _065_ a_8386_8457# 0.00191f
C3156 net32 net49 1.42e-20
C3157 net27 a_911_10217# 1.76e-21
C3158 net15 _051_ 2.07e-20
C3159 _050_ calibrate 0.573f
C3160 a_10137_4943# trim_mask\[4\] 2.53e-20
C3161 _074_ _083_ 0.0735f
C3162 net16 net9 0.00341f
C3163 en_co_clk a_5054_4399# 4.78e-19
C3164 net4 net55 1.05e-20
C3165 a_6428_7119# VPWR 0.0849f
C3166 a_10005_6031# cal_count\[3\] 0.0022f
C3167 net21 a_4043_12393# 1.32e-19
C3168 a_13183_3311# VPWR 0.201f
C3169 net15 _014_ 0.0791f
C3170 _048_ a_8298_2767# 3.38e-21
C3171 _110_ a_14099_1929# 1.47e-19
C3172 a_7263_7093# net30 2.19e-20
C3173 a_561_7119# result[1] 0.00876f
C3174 a_2143_2229# VPWR 0.476f
C3175 a_1000_11293# VPWR 0.0859f
C3176 trim_mask\[2\] a_9761_1679# 1.44e-20
C3177 _034_ _093_ 1.2e-21
C3178 _064_ a_10055_5487# 0.0518f
C3179 a_12061_7669# a_13050_7637# 0.0728f
C3180 a_12520_7637# a_12344_8041# 0.26f
C3181 _134_ a_13257_4943# 4.73e-20
C3182 a_1651_6005# a_1476_6031# 0.234f
C3183 a_10864_7387# _136_ 0.00208f
C3184 trim_mask\[0\] _112_ 1.56e-19
C3185 _078_ a_1638_7485# 1.46e-19
C3186 _085_ VPWR 0.278f
C3187 net43 net12 0.00841f
C3188 a_7723_6807# _048_ 1.4e-20
C3189 trim_mask\[0\] a_7758_4759# 4.03e-19
C3190 calibrate _052_ 0.233f
C3191 mask\[6\] a_5997_11247# 0.00348f
C3192 net28 a_1357_11293# 2.68e-20
C3193 a_4609_1679# a_5177_1921# 0.181f
C3194 a_4443_1679# a_4959_1679# 0.115f
C3195 _102_ a_1677_9545# 3.99e-20
C3196 _048_ a_7210_5807# 2.21e-19
C3197 _045_ net44 2.82e-20
C3198 net26 mask\[4\] 0.718f
C3199 a_3597_10933# a_2953_9845# 1.07e-20
C3200 calibrate _098_ 0.382f
C3201 _041_ mask\[1\] 0.0171f
C3202 a_11691_4399# VPWR 0.144f
C3203 a_4674_10927# _019_ 8.1e-21
C3204 net46 a_9802_4007# 0.00143f
C3205 net2 a_13825_5185# 1.86e-20
C3206 a_1129_4373# a_1019_4399# 0.0977f
C3207 a_10688_9295# a_10774_9661# 0.00972f
C3208 a_10864_9269# a_11168_9661# 3.11e-19
C3209 _001_ a_9677_8457# 0.0121f
C3210 a_4815_3031# VPWR 0.268f
C3211 a_1835_11231# _102_ 0.00375f
C3212 _130_ a_14870_7369# 0.00145f
C3213 net4 a_7715_3285# 8.59e-22
C3214 _020_ a_7723_10143# 6.17e-19
C3215 net3 a_3817_4697# 0.0158f
C3216 net18 a_11168_9661# 7.18e-19
C3217 net27 mask\[2\] 4.53e-21
C3218 net44 a_4696_8207# 0.234f
C3219 net53 a_6793_8970# 0.12f
C3220 net46 _108_ 0.0945f
C3221 _067_ a_9459_7895# 0.248f
C3222 net49 VPWR 0.357f
C3223 _078_ a_1585_10217# 3.02e-19
C3224 a_9269_2589# VPWR 2.28e-19
C3225 net30 a_1493_5487# 0.0281f
C3226 _074_ a_911_7119# 0.0157f
C3227 _068_ a_9460_6807# 0.0783f
C3228 _065_ a_8091_7967# 6.43e-20
C3229 a_14733_9545# VPWR 0.0085f
C3230 _053_ a_10055_5487# 2.1e-19
C3231 trim_val\[1\] _056_ 5.31e-19
C3232 _059_ state\[1\] 0.00785f
C3233 clknet_2_0__leaf_clk net3 0.0115f
C3234 _115_ a_13307_1707# 0.119f
C3235 _094_ a_4883_6397# 8.78e-22
C3236 net29 a_3597_12021# 0.0017f
C3237 _002_ a_7256_8029# 0.183f
C3238 clknet_2_3__leaf_clk a_11057_4105# 1.28e-20
C3239 a_9761_1679# a_9719_1473# 1.13e-21
C3240 _064_ trim_val\[4\] 0.0378f
C3241 a_11987_8757# a_12341_8751# 0.0675f
C3242 a_745_12021# a_1822_12015# 1.46e-19
C3243 net43 a_3852_12381# 0.00219f
C3244 net34 a_14972_5193# 0.0078f
C3245 net11 a_8767_591# 0.178f
C3246 a_10903_7261# _066_ 2.59e-21
C3247 net46 a_10655_2932# 0.00431f
C3248 a_13257_4943# a_13915_4399# 4.56e-20
C3249 _047_ _110_ 2.45e-20
C3250 _122_ a_13557_7369# 0.0108f
C3251 a_10864_7387# a_10861_7119# 2.36e-20
C3252 net52 a_2787_10927# 0.245f
C3253 net43 a_1651_10143# 0.337f
C3254 a_1660_11305# a_3431_10933# 3.16e-20
C3255 net19 ctlp[6] 1.79e-21
C3256 net45 a_911_4777# 0.153f
C3257 a_395_591# en 1.99e-20
C3258 _065_ _059_ 0.00213f
C3259 a_7843_3677# VPWR 1.7e-19
C3260 a_929_8757# a_1476_7119# 7.29e-21
C3261 net46 a_9115_2223# 0.0122f
C3262 _037_ a_12249_7663# 0.149f
C3263 a_1279_9129# a_911_7119# 5.29e-20
C3264 a_1644_12533# a_1493_11721# 1.79e-20
C3265 _110_ _116_ 0.503f
C3266 _092_ a_4308_4917# 0.0198f
C3267 a_9443_6059# VPWR 0.205f
C3268 net14 a_745_12021# 0.0067f
C3269 a_1099_12533# a_1313_11989# 0.00321f
C3270 a_11601_2229# VPWR 0.612f
C3271 _078_ mask\[3\] 0.248f
C3272 net40 net30 0.0489f
C3273 a_4674_10927# VPWR 8.1e-19
C3274 net43 a_1830_7119# 0.00384f
C3275 _070_ a_6485_8181# 5.95e-22
C3276 _067_ en_co_clk 0.0436f
C3277 _122_ net2 0.244f
C3278 net1 net41 0.0625f
C3279 net17 VPWR 1.33f
C3280 _091_ a_9529_6059# 5.76e-19
C3281 _053_ _088_ 0.00465f
C3282 a_3431_12021# a_3597_12021# 0.582f
C3283 net13 net3 0.0105f
C3284 _085_ net27 0.0174f
C3285 _063_ _106_ 0.0377f
C3286 a_2313_6183# _120_ 2.11e-20
C3287 a_7571_4943# _103_ 0.0649f
C3288 net19 clknet_2_3__leaf_clk 0.0276f
C3289 net4 _093_ 2.32e-20
C3290 _053_ a_7262_5461# 2.5e-19
C3291 a_4609_1679# a_5633_1679# 2.36e-20
C3292 a_9595_1679# a_9761_1679# 0.906f
C3293 net24 a_2689_8751# 0.0111f
C3294 net45 net7 1.3e-20
C3295 trim_mask\[4\] a_11321_3855# 2.84e-19
C3296 net35 trim_val\[1\] 0.00225f
C3297 a_10569_1109# _057_ 1.13e-19
C3298 a_10688_9295# _065_ 4.08e-20
C3299 net2 _063_ 1.05e-19
C3300 net18 a_10752_565# 0.00701f
C3301 net26 a_7091_9839# 0.0265f
C3302 _000_ cal_itt\[2\] 0.00363f
C3303 net46 a_9004_3677# 2.46e-19
C3304 a_5087_3855# VPWR 0.24f
C3305 net36 a_15023_10927# 0.218f
C3306 _072_ _049_ 1.81e-20
C3307 a_1313_10901# net26 7.11e-20
C3308 _136_ _111_ 0.0028f
C3309 a_763_8757# _081_ 0.00169f
C3310 net46 a_12516_2601# 0.266f
C3311 a_7569_7637# a_8025_8041# 4.2e-19
C3312 a_6835_7669# a_7459_7663# 9.73e-19
C3313 a_7351_8041# a_7613_8029# 0.00171f
C3314 a_14655_4399# a_15083_4659# 0.0126f
C3315 net14 _014_ 3.31e-19
C3316 a_12061_7669# VPWR 0.311f
C3317 clknet_2_2__leaf_clk clk 0.0052f
C3318 a_14199_7369# a_14282_7119# 1.58e-20
C3319 clknet_0_clk a_5515_6005# 2.34e-19
C3320 a_4443_1679# VPWR 0.518f
C3321 net46 _107_ 0.00233f
C3322 a_1644_12533# VPWR 0.294f
C3323 clknet_2_1__leaf_clk a_3511_11471# 4.52e-19
C3324 net43 result[2] 5.53e-20
C3325 a_1476_4777# VPWR 0.299f
C3326 clknet_2_3__leaf_clk cal_itt\[1\] 0.00118f
C3327 trim_mask\[0\] a_11583_4777# 5.05e-19
C3328 cal_itt\[0\] a_10975_6031# 1.88e-19
C3329 _078_ a_1579_5807# 0.00106f
C3330 a_2383_3689# a_2143_2229# 1.37e-20
C3331 trim_mask\[4\] a_11435_2229# 4.49e-19
C3332 a_2601_3285# a_2309_2229# 1.78e-20
C3333 trim_mask\[2\] a_11067_3017# 0.172f
C3334 a_10699_3311# trim_mask\[3\] 3.91e-19
C3335 net45 a_4425_6031# 2.77e-20
C3336 a_9595_1679# a_10787_1135# 1.03e-19
C3337 net37 clkc 5.01e-19
C3338 net18 a_10781_3311# 0.0056f
C3339 a_10055_2767# _026_ 4.89e-21
C3340 _063_ _033_ 1.18e-21
C3341 _013_ clk 1.58e-19
C3342 a_2174_8457# VPWR 0.00335f
C3343 _068_ a_8495_6895# 0.00289f
C3344 net21 _042_ 4.64e-20
C3345 net52 _049_ 2.01e-19
C3346 _112_ _030_ 0.0213f
C3347 _113_ a_13625_3317# 6.65e-20
C3348 mask\[5\] a_5997_10927# 0.0136f
C3349 net40 _134_ 1.8e-19
C3350 net16 a_13415_2442# 6.84e-19
C3351 net54 a_4863_4917# 0.201f
C3352 a_4091_5309# _060_ 2.07e-20
C3353 net18 a_11801_4373# 7.42e-19
C3354 _107_ a_5931_4105# 7.58e-19
C3355 state\[2\] a_6737_3855# 3.69e-19
C3356 _130_ _131_ 0.203f
C3357 a_8091_7967# _067_ 2.17e-19
C3358 a_2828_12131# VPWR 0.178f
C3359 _050_ _015_ 6.2e-21
C3360 net50 a_9761_1679# 0.00563f
C3361 a_14172_1513# VPWR 0.303f
C3362 mask\[1\] a_3615_8207# 0.00686f
C3363 net43 a_1191_11305# 9.54e-19
C3364 a_2948_3689# a_3339_2767# 0.00133f
C3365 _101_ a_3840_8867# 1.1e-20
C3366 _096_ a_3667_3829# 0.00593f
C3367 a_11895_7669# a_12430_7663# 6.02e-19
C3368 _078_ a_4043_11305# 1.55e-19
C3369 net30 _024_ 1.38e-20
C3370 net28 a_3597_12021# 0.0255f
C3371 clknet_2_0__leaf_clk a_1476_7119# 0.00133f
C3372 a_15159_9269# VPWR 0.219f
C3373 a_10676_1679# trim_val\[3\] 0.00159f
C3374 clknet_2_0__leaf_clk mask\[0\] 0.0635f
C3375 _094_ a_4993_6273# 0.0133f
C3376 _057_ a_11374_1251# 4.96e-19
C3377 _101_ a_2971_8457# 0.147f
C3378 clknet_2_0__leaf_clk valid 0.00553f
C3379 a_10383_7093# a_10005_6031# 0.00128f
C3380 clknet_2_3__leaf_clk _001_ 0.381f
C3381 net45 a_3868_7119# 0.00151f
C3382 clknet_2_3__leaf_clk a_11067_4405# 3.43e-20
C3383 _053_ a_8745_4943# 0.00116f
C3384 net16 a_13470_7663# 0.00324f
C3385 _019_ a_4609_9295# 0.253f
C3386 _026_ a_12691_2527# 1.29e-20
C3387 a_6906_2355# a_7310_2223# 0.0512f
C3388 a_7223_2465# a_7379_2197# 0.112f
C3389 mask\[6\] a_1095_11305# 1.16e-21
C3390 _095_ _087_ 3.83e-20
C3391 a_13091_4943# _047_ 1.63e-20
C3392 net28 a_1137_11721# 3.5e-19
C3393 net4 a_9595_5193# 8.17e-19
C3394 _092_ _090_ 0.187f
C3395 net33 a_14981_4020# 0.00588f
C3396 a_15023_12015# trimb[2] 0.337f
C3397 _014_ a_2659_2601# 0.00234f
C3398 _012_ a_1201_3855# 1.97e-19
C3399 net47 a_9195_10357# 0.294f
C3400 a_8673_10625# a_9020_10383# 0.0512f
C3401 a_10016_1679# VPWR 0.1f
C3402 a_8105_10383# _043_ 7e-20
C3403 _020_ _042_ 0.0462f
C3404 _120_ VPWR 0.327f
C3405 net50 a_10787_1135# 0.0493f
C3406 mask\[2\] clknet_0_clk 1.5e-19
C3407 a_1644_12533# net27 1.35e-21
C3408 a_3116_12533# ctlp[1] 0.166f
C3409 _078_ a_4687_11231# 1.76e-20
C3410 net47 _128_ 0.0987f
C3411 a_13512_4943# _058_ 0.00217f
C3412 a_13715_5309# a_13697_4373# 2.18e-21
C3413 _095_ _099_ 0.0338f
C3414 _128_ a_14377_9545# 0.072f
C3415 a_2601_3285# a_3110_3311# 2.6e-19
C3416 net44 _078_ 0.0366f
C3417 state\[1\] a_3399_2527# 0.0668f
C3418 a_2033_3317# a_4658_3427# 1.56e-20
C3419 net13 mask\[0\] 0.00197f
C3420 a_15083_4659# trim[1] 0.343f
C3421 _037_ a_11059_7356# 2.7e-19
C3422 trim_mask\[3\] _027_ 0.0622f
C3423 a_1651_10143# a_2953_9845# 3.21e-20
C3424 net3 a_4091_4943# 0.00452f
C3425 _095_ a_1129_4373# 1.86e-20
C3426 a_3597_12021# a_4167_11471# 6.61e-20
C3427 cal_itt\[2\] _053_ 3.35e-19
C3428 a_3597_10933# a_4043_11305# 2.28e-19
C3429 _028_ a_8912_2589# 1.13e-20
C3430 a_561_9845# a_2787_9845# 1.7e-22
C3431 a_2755_2601# clk 5.58e-19
C3432 _125_ _133_ 4.17e-21
C3433 a_1000_12381# VPWR 0.0836f
C3434 _027_ a_10689_2543# 1.97e-19
C3435 clknet_2_0__leaf_clk _079_ 0.0308f
C3436 net46 a_10838_2045# 2.76e-19
C3437 _104_ a_11601_2229# 5.06e-20
C3438 _071_ net30 1.26e-19
C3439 a_11396_6031# VPWR 0.0776f
C3440 _065_ _108_ 8.54e-20
C3441 _101_ a_2225_7983# 0.00145f
C3442 a_4863_4917# a_4471_4007# 9.24e-21
C3443 a_9317_3285# trim_mask\[2\] 1.41e-21
C3444 a_455_12533# VPWR 0.402f
C3445 a_9099_3689# a_9664_3689# 7.99e-20
C3446 _131_ a_13821_7119# 0.00951f
C3447 a_4609_9295# VPWR 0.407f
C3448 _062_ a_7019_4407# 1.74e-19
C3449 _051_ a_7460_5807# 0.00187f
C3450 net54 a_3817_4697# 1.53e-19
C3451 a_4091_5309# a_4498_4373# 0.0237f
C3452 a_4871_8181# a_4995_7119# 2.76e-20
C3453 net28 a_1357_12381# 7.38e-19
C3454 _110_ a_13183_3311# 0.00989f
C3455 mask\[5\] a_8767_11471# 0.00284f
C3456 a_2288_3677# cal 3.68e-20
C3457 net25 _082_ 0.415f
C3458 a_6835_7669# a_6523_7119# 0.00347f
C3459 trim_mask\[1\] a_11764_3677# 0.0164f
C3460 trim_mask\[2\] a_11856_2589# 8.76e-20
C3461 a_2815_9447# a_2961_9295# 0.0134f
C3462 a_5177_9537# a_4959_9295# 0.21f
C3463 a_4609_9295# a_5699_9269# 0.0424f
C3464 a_4443_9295# a_5524_9295# 0.102f
C3465 net2 comp 0.0198f
C3466 _054_ a_7104_3855# 1.88e-20
C3467 net21 a_3597_12021# 8.73e-19
C3468 _005_ net22 0.00141f
C3469 a_12077_3285# a_12586_3311# 2.6e-19
C3470 net47 a_8949_9537# 0.171f
C3471 a_8298_5487# a_8389_5193# 9e-20
C3472 _104_ a_5087_3855# 2.64e-21
C3473 a_4165_10901# a_3947_11305# 0.21f
C3474 a_3597_10933# a_4687_11231# 0.0424f
C3475 net14 _082_ 0.00888f
C3476 _051_ a_6927_3311# 2.34e-19
C3477 a_1549_6794# a_1476_6031# 8.52e-19
C3478 _039_ a_1651_6005# 0.0346f
C3479 a_11141_6031# a_13441_6281# 1.22e-20
C3480 net37 a_15023_9839# 0.218f
C3481 a_3521_9813# mask\[2\] 2.7e-19
C3482 a_3303_10217# a_3411_9839# 0.0572f
C3483 net46 a_11587_6031# 0.00108f
C3484 a_11709_6273# a_11753_6031# 3.69e-19
C3485 a_3868_10217# a_3977_10217# 0.00742f
C3486 a_4043_10143# a_4222_10205# 0.0074f
C3487 clknet_2_1__leaf_clk net2 0.0109f
C3488 _101_ a_6793_8970# 3.72e-21
C3489 _125_ a_14236_8457# 0.00518f
C3490 _110_ a_11691_4399# 6.5e-21
C3491 _129_ a_12520_7637# 2.33e-21
C3492 a_6541_12021# a_7109_11989# 0.186f
C3493 net3 a_2948_3689# 9.66e-19
C3494 net47 a_11895_7669# 0.0445f
C3495 _041_ _002_ 3.63e-20
C3496 a_2953_7119# a_3868_7119# 0.125f
C3497 a_2787_7119# a_3208_7119# 0.0867f
C3498 _058_ a_11859_3689# 0.0026f
C3499 _065_ a_9460_6807# 8.83e-20
C3500 net12 mask\[3\] 0.011f
C3501 net15 net22 4.98e-20
C3502 _088_ a_7379_2197# 1.96e-21
C3503 net43 a_1651_6005# 2.34e-20
C3504 ctln[6] ctln[5] 0.00305f
C3505 net12 a_6741_7361# 0.00389f
C3506 _069_ a_9957_7663# 0.1f
C3507 net15 a_2921_2589# 5.85e-19
C3508 a_6909_10933# _020_ 3.29e-20
C3509 _074_ mask\[4\] 0.189f
C3510 _004_ a_1579_5807# 1.84e-21
C3511 _108_ a_11233_4405# 0.00281f
C3512 _050_ a_7184_2339# 0.00139f
C3513 net13 a_4973_2773# 6.93e-19
C3514 _097_ a_3148_4399# 0.0012f
C3515 a_7527_4631# _107_ 0.00952f
C3516 _110_ net49 8.81e-19
C3517 net29 net43 0.0617f
C3518 a_6822_4105# VPWR 0.00468f
C3519 net34 a_13257_1141# 2.5e-19
C3520 net19 a_8827_9295# 0.00129f
C3521 a_4259_6031# _095_ 0.00525f
C3522 clknet_2_0__leaf_clk a_448_6549# 0.0311f
C3523 net50 a_11067_3017# 0.00128f
C3524 _053_ a_11297_7119# 6.41e-19
C3525 clknet_2_3__leaf_clk a_11394_9509# 0.0623f
C3526 a_1129_9813# a_1019_9839# 0.0977f
C3527 _058_ a_11845_4765# 4.69e-19
C3528 a_12323_4703# _109_ 1.29e-19
C3529 net13 net54 0.0449f
C3530 a_3365_4943# _097_ 2.12e-19
C3531 trim_mask\[3\] _117_ 6.22e-19
C3532 a_561_7119# a_1476_7119# 0.125f
C3533 net43 _040_ 8.69e-20
C3534 a_13607_4943# a_13512_4943# 0.0498f
C3535 a_14347_4917# a_14972_5193# 0.00113f
C3536 net44 a_5502_6397# 2.59e-19
C3537 a_13825_5185# a_13715_5309# 0.0977f
C3538 mask\[0\] a_561_7119# 3.45e-20
C3539 a_12691_2527# _031_ 0.00166f
C3540 a_11601_2229# a_12678_2223# 1.46e-19
C3541 net45 a_7140_2223# 3.47e-19
C3542 net45 _121_ 2.82e-20
C3543 _021_ a_5997_11247# 6.05e-20
C3544 _031_ _114_ 0.00585f
C3545 net31 comp 0.149f
C3546 _000_ a_8636_9295# 0.16f
C3547 a_8215_9295# a_8839_9661# 9.73e-19
C3548 _049_ a_7527_4631# 0.0102f
C3549 net46 trim_mask\[4\] 0.468f
C3550 clknet_2_1__leaf_clk net24 0.0488f
C3551 a_2865_4460# a_3057_4719# 0.00424f
C3552 net15 a_3133_11247# 5.93e-19
C3553 _074_ net20 0.00949f
C3554 _053_ net55 0.0461f
C3555 clknet_2_1__leaf_clk _084_ 0.277f
C3556 a_1095_12393# a_1660_12393# 7.99e-20
C3557 trim_val\[4\] a_9664_3689# 0.00135f
C3558 a_455_12533# net27 1.41e-19
C3559 net43 a_3431_12021# 0.311f
C3560 a_1099_12533# ctlp[1] 5.95e-22
C3561 a_11141_6031# _066_ 1.06e-20
C3562 calibrate _087_ 0.0116f
C3563 _049_ state\[1\] 6.95e-20
C3564 _041_ a_3615_8207# 7.84e-19
C3565 _110_ a_11601_2229# 2.48e-19
C3566 _125_ _129_ 0.0064f
C3567 _025_ VPWR 0.333f
C3568 clknet_2_3__leaf_clk a_13193_6031# 0.00307f
C3569 net2 a_13111_6031# 0.398f
C3570 clknet_2_3__leaf_clk a_11116_8983# 0.00387f
C3571 calibrate a_6519_3829# 0.0432f
C3572 _026_ VPWR 0.389f
C3573 _033_ a_9761_1679# 6.71e-22
C3574 _044_ a_8105_10383# 1.39e-21
C3575 a_1651_10143# mask\[3\] 0.00292f
C3576 a_5363_4719# a_5445_4399# 8.13e-19
C3577 a_929_8757# a_1125_7663# 2.38e-20
C3578 net38 a_15023_10927# 0.0398f
C3579 a_3868_7119# a_2857_5461# 1.63e-20
C3580 net33 trim_mask\[2\] 0.00626f
C3581 a_745_12021# a_1493_11721# 1.97e-19
C3582 a_5502_6397# en_co_clk 7.91e-20
C3583 trim_mask\[0\] a_15023_5487# 9.4e-19
C3584 mask\[1\] a_4227_8207# 7.19e-21
C3585 _048_ a_8307_4719# 0.00344f
C3586 calibrate _099_ 4.75e-19
C3587 _065_ _049_ 0.339f
C3588 _131_ trim[4] 3.48e-21
C3589 a_448_11445# a_579_10933# 3.72e-19
C3590 _067_ _108_ 2.97e-19
C3591 a_3273_4943# a_3557_5193# 0.0148f
C3592 net9 clknet_2_3__leaf_clk 0.162f
C3593 mask\[2\] a_2775_9071# 0.0105f
C3594 _056_ a_14686_2339# 4.96e-19
C3595 net19 _116_ 0.00268f
C3596 net52 a_4036_8207# 5.81e-19
C3597 cal_count\[3\] _111_ 0.00281f
C3598 a_2368_9955# net24 0.00108f
C3599 _101_ net30 4.32e-20
C3600 _090_ a_5536_4399# 0.022f
C3601 a_395_4405# a_855_4105# 1.81e-19
C3602 calibrate a_1129_4373# 0.0238f
C3603 a_1867_3317# VPWR 0.522f
C3604 net4 a_9166_4515# 1.65e-19
C3605 _049_ a_5054_4399# 2.35e-19
C3606 clknet_0_clk a_5087_3855# 4.43e-21
C3607 a_12153_8757# a_12522_8751# 4.45e-20
C3608 a_13142_7271# a_13356_7369# 0.013f
C3609 a_579_10933# a_1203_10927# 9.73e-19
C3610 a_4498_4373# a_4886_4399# 0.00167f
C3611 _107_ a_11233_4405# 5.4e-21
C3612 net16 a_14788_7369# 2.83e-19
C3613 net4 ctln[1] 0.0343f
C3614 _074_ a_1313_10901# 0.00387f
C3615 trim_val\[4\] a_10781_3631# 4.68e-19
C3616 net40 _118_ 0.129f
C3617 a_13142_8359# _133_ 1.09e-20
C3618 a_7001_7669# a_9459_7895# 6.08e-20
C3619 _078_ a_1184_9117# 3.69e-19
C3620 a_7677_4759# VPWR 1.14e-19
C3621 net44 a_7001_7669# 0.0117f
C3622 _108_ clknet_2_2__leaf_clk 0.124f
C3623 a_6181_10633# VPWR 0.178f
C3624 _067_ a_9460_6807# 0.187f
C3625 a_11168_9661# VPWR 0.0046f
C3626 net2 a_6485_8181# 0.147f
C3627 trim_mask\[4\] a_11343_3317# 9.71e-19
C3628 net13 a_4471_4007# 0.00819f
C3629 trim_mask\[4\] a_11149_3017# 0.00592f
C3630 _123_ _134_ 2.37e-20
C3631 a_745_12021# VPWR 0.59f
C3632 net37 a_14715_3615# 9e-19
C3633 net14 net22 0.467f
C3634 a_9761_1679# a_10785_1679# 2.36e-20
C3635 a_2019_9055# mask\[1\] 0.00327f
C3636 a_1844_9129# a_2092_8457# 1.48e-19
C3637 _040_ a_2857_7637# 0.00524f
C3638 a_745_12021# a_1769_12393# 2.36e-20
C3639 a_1313_11989# a_1357_12381# 3.69e-19
C3640 net43 a_1191_12393# 9.54e-19
C3641 net53 a_5089_10159# 0.00321f
C3642 net41 a_2143_2229# 1.11e-20
C3643 net44 a_6888_10205# 8.11e-19
C3644 _043_ a_9074_9955# 4.96e-19
C3645 _006_ a_2092_8457# 4.01e-20
C3646 _074_ _081_ 0.0746f
C3647 a_2953_7119# _121_ 3.72e-20
C3648 _050_ _052_ 0.349f
C3649 net44 net12 0.0433f
C3650 clknet_2_2__leaf_clk a_10655_2932# 0.0284f
C3651 net39 net33 1.61e-20
C3652 net28 net43 0.435f
C3653 net45 a_3273_4943# 4.61e-20
C3654 a_3302_3677# VPWR 6.13e-20
C3655 net2 a_13825_6031# 3.31e-19
C3656 a_5455_4943# a_5731_4943# 0.00119f
C3657 mask\[0\] a_4167_6575# 4.16e-20
C3658 trim_mask\[2\] trim_val\[3\] 3.18e-19
C3659 _050_ _098_ 0.201f
C3660 _051_ VPWR 2.08f
C3661 a_13091_4943# net49 5.23e-20
C3662 a_4349_8449# a_4805_8207# 4.2e-19
C3663 a_7001_7669# clk 0.00448f
C3664 clknet_2_2__leaf_clk a_9115_2223# 0.00252f
C3665 a_7001_7669# en_co_clk 3.91e-21
C3666 net4 a_9007_2601# 3.94e-19
C3667 _076_ a_6198_8534# 0.00733f
C3668 clk ctln[7] 1.18e-20
C3669 clknet_2_3__leaf_clk a_10188_4105# 3.62e-21
C3670 a_10747_8970# _041_ 0.0515f
C3671 _014_ VPWR 1f
C3672 _074_ a_6987_12393# 5.75e-21
C3673 net34 a_14981_4020# 2.42e-20
C3674 net13 a_4970_4399# 9.18e-19
C3675 a_561_7119# a_448_6549# 2.68e-19
C3676 a_395_7119# net22 1.73e-19
C3677 net41 a_4815_3031# 3.77e-20
C3678 _122_ a_11059_7356# 0.0129f
C3679 _080_ net45 0.00397f
C3680 _056_ a_15023_1679# 0.208f
C3681 a_1279_9129# _081_ 6.06e-19
C3682 _074_ a_455_5747# 0.0204f
C3683 net44 a_5340_6031# 0.263f
C3684 a_10383_7093# a_10864_7387# 0.0424f
C3685 _119_ a_9369_3855# 3.7e-19
C3686 a_6741_7361# a_6631_7485# 0.0977f
C3687 a_6523_7119# a_6428_7119# 0.0498f
C3688 a_8022_7119# a_10903_7261# 8.33e-21
C3689 net53 a_6633_9845# 0.0181f
C3690 a_4091_5309# a_4175_4943# 0.00101f
C3691 clknet_2_1__leaf_clk a_4677_7882# 4.73e-19
C3692 _117_ net11 1.72e-19
C3693 a_6891_12393# a_7153_12381# 0.00171f
C3694 net44 a_6983_10217# 0.156f
C3695 _048_ a_6822_4399# 0.0158f
C3696 _098_ _052_ 0.141f
C3697 a_13625_3317# a_13881_2741# 0.00164f
C3698 net19 a_9182_10749# 1.39e-19
C3699 net12 clk 0.0267f
C3700 net30 a_8749_3317# 5.93e-22
C3701 net12 en_co_clk 0.013f
C3702 _091_ _038_ 1.84e-20
C3703 _110_ a_10016_1679# 0.00206f
C3704 net42 a_7571_4943# 0.147f
C3705 _094_ net3 0.0127f
C3706 _125_ a_14318_8457# 2.24e-19
C3707 a_3116_12533# net15 0.191f
C3708 net40 a_10137_4943# 0.039f
C3709 mask\[5\] _020_ 0.00752f
C3710 a_10752_565# VPWR 0.297f
C3711 _092_ _106_ 2.91e-20
C3712 clknet_2_2__leaf_clk a_12516_2601# 0.00393f
C3713 clknet_0_clk _120_ 8.5e-19
C3714 _031_ VPWR 0.426f
C3715 net43 a_4167_11471# 0.0159f
C3716 _108_ ctln[2] 1.05e-19
C3717 a_8563_10749# a_8215_9295# 2.28e-20
C3718 clknet_2_2__leaf_clk _107_ 0.00487f
C3719 _118_ _024_ 1.14e-20
C3720 _121_ a_2857_5461# 0.00357f
C3721 a_5340_6031# en_co_clk 0.05f
C3722 net46 a_12723_4943# 0.0145f
C3723 trim_mask\[0\] a_7800_4631# 0.0225f
C3724 clknet_2_0__leaf_clk a_4871_8181# 2.89e-20
C3725 _119_ a_9747_2527# 4.21e-20
C3726 _033_ a_11067_3017# 9.34e-20
C3727 _078_ result[3] 3.52e-19
C3728 _064_ a_9595_5193# 0.195f
C3729 trim_val\[3\] a_9719_1473# 2.68e-19
C3730 a_5524_9295# _065_ 3.11e-20
C3731 _076_ clknet_2_0__leaf_clk 0.00551f
C3732 clknet_2_3__leaf_clk _062_ 0.177f
C3733 a_5445_4399# VPWR 0.00532f
C3734 a_745_12021# net27 8.02e-20
C3735 net2 a_14199_7369# 3.72e-20
C3736 net45 a_816_6031# 2.47e-19
C3737 net53 a_6445_10383# 0.00204f
C3738 clknet_2_3__leaf_clk a_11508_9295# 3.98e-19
C3739 a_7527_4631# trim_mask\[4\] 8.9e-21
C3740 clknet_2_3__leaf_clk a_10138_5807# 5.14e-19
C3741 net44 a_8551_10383# 4.2e-19
C3742 mask\[4\] _083_ 0.365f
C3743 net5 _061_ 0.00366f
C3744 net39 ctlp[2] 0.0015f
C3745 a_561_9845# a_763_8757# 0.00127f
C3746 a_395_9845# a_929_8757# 6.43e-21
C3747 net54 a_2948_3689# 2.02e-20
C3748 _104_ _025_ 0.00198f
C3749 a_2877_2197# a_3333_2601# 4.2e-19
C3750 a_2659_2601# a_2921_2589# 0.00171f
C3751 a_2143_2229# a_2767_2223# 9.73e-19
C3752 net46 _056_ 4.84e-20
C3753 a_10781_3311# VPWR 0.196f
C3754 _104_ _026_ 0.00621f
C3755 net21 net43 0.0469f
C3756 a_7569_7637# a_7351_8041# 0.21f
C3757 a_6835_7669# a_7916_8041# 0.102f
C3758 a_7001_7669# a_8091_7967# 0.0424f
C3759 a_8083_8181# a_8301_8207# 0.0326f
C3760 a_2033_3317# a_2601_3285# 0.186f
C3761 a_1867_3317# a_2383_3689# 0.111f
C3762 mask\[1\] a_3053_8457# 0.00164f
C3763 net18 cal_itt\[0\] 4.6e-19
C3764 a_13356_8457# VPWR 0.00902f
C3765 a_11801_4373# VPWR 0.221f
C3766 a_5633_9295# net51 1.93e-20
C3767 net2 cal_itt\[3\] 2.98e-22
C3768 net13 a_4871_8181# 0.0124f
C3769 mask\[4\] net4 1.18e-20
C3770 net6 a_1276_565# 0.211f
C3771 a_12992_8751# net2 2.56e-20
C3772 a_5087_3855# net41 0.00163f
C3773 _032_ a_10373_1679# 1.01e-19
C3774 a_9595_1679# trim_val\[3\] 0.0124f
C3775 net13 _076_ 1.04e-20
C3776 net46 a_11491_6031# 0.153f
C3777 a_11141_6031# a_12056_6031# 0.119f
C3778 trim_mask\[1\] a_13975_3689# 7.04e-19
C3779 a_4512_11305# mask\[2\] 4.31e-20
C3780 net26 a_561_9845# 8.49e-20
C3781 _074_ result[5] 2.8e-19
C3782 _095_ _097_ 9.72e-19
C3783 a_15023_6031# net35 1.73e-19
C3784 _072_ a_8761_7983# 0.0096f
C3785 net4 _064_ 0.0666f
C3786 _096_ a_3339_2767# 5.43e-19
C3787 net44 a_6197_6281# 2.44e-19
C3788 _099_ _015_ 3.09e-20
C3789 net41 a_4443_1679# 1.75e-20
C3790 a_7613_8029# VPWR 1.7e-19
C3791 net46 a_11967_3311# 0.0122f
C3792 mask\[6\] a_3511_11471# 0.00965f
C3793 net30 a_7939_3855# 0.185f
C3794 _106_ a_9317_3285# 6.44e-20
C3795 _068_ a_8761_7983# 1.96e-19
C3796 _108_ a_14540_3689# 0.0171f
C3797 state\[2\] a_6703_2197# 6.97e-19
C3798 net45 a_1651_7093# 0.0158f
C3799 a_1467_7923# a_1476_7119# 0.00423f
C3800 mask\[4\] a_8360_10383# 1.8e-19
C3801 net3 a_4617_3855# 1.2e-19
C3802 a_1467_7923# mask\[0\] 0.00867f
C3803 a_1549_6794# _039_ 0.194f
C3804 a_1638_6397# VPWR 6.74e-19
C3805 net46 net35 0.00522f
C3806 a_6210_4989# _103_ 4.25e-20
C3807 net46 a_13059_4631# 2.04e-20
C3808 net12 _059_ 4.92e-20
C3809 net43 a_1549_6794# 0.0341f
C3810 a_2601_3285# a_2491_3311# 0.0977f
C3811 net37 _047_ 0.454f
C3812 net16 a_12231_6005# 2.94e-20
C3813 a_7715_3285# a_7379_2197# 3.65e-21
C3814 a_7010_3311# a_7310_2223# 7.97e-21
C3815 a_5535_8181# VPWR 0.396f
C3816 a_7999_11231# clknet_2_3__leaf_clk 5.51e-21
C3817 en_co_clk a_6197_6281# 0.00235f
C3818 _060_ state\[2\] 1.84e-19
C3819 a_1313_11989# net43 0.176f
C3820 net44 a_6631_7485# 0.013f
C3821 a_855_4105# a_2283_4020# 5.09e-20
C3822 a_11233_4405# trim_mask\[4\] 0.00205f
C3823 _014_ a_2383_3689# 0.0124f
C3824 net16 a_13880_3677# 0.00323f
C3825 a_2787_10927# a_2869_11247# 0.00393f
C3826 a_11098_6691# _136_ 1.5e-19
C3827 a_2857_5461# a_3273_4943# 0.0142f
C3828 a_2971_8457# a_3053_8207# 0.00393f
C3829 net4 _053_ 1.21f
C3830 net19 a_9269_2589# 3.89e-19
C3831 a_14099_3017# net48 1.06e-19
C3832 net45 a_937_4105# 0.00122f
C3833 cal_count\[0\] _125_ 0.504f
C3834 a_5340_6031# _059_ 4.98e-19
C3835 _111_ a_11679_4777# 1.76e-19
C3836 _060_ state\[0\] 0.0791f
C3837 net34 trim_mask\[2\] 2.69e-19
C3838 net38 a_15023_12015# 0.215f
C3839 net47 net40 1.13e-20
C3840 a_5699_9269# a_5535_8181# 9.72e-19
C3841 a_4864_9295# a_4871_8181# 2.48e-20
C3842 _051_ _104_ 0.00947f
C3843 _122_ a_11016_6691# 0.111f
C3844 mask\[0\] _094_ 0.0519f
C3845 mask\[3\] _040_ 3.21e-20
C3846 net16 a_13697_4373# 0.0035f
C3847 net50 trim_val\[3\] 0.0617f
C3848 a_8583_3317# a_9099_3689# 0.109f
C3849 _082_ VPWR 0.403f
C3850 net12 a_7197_7119# 8.28e-20
C3851 _061_ a_15023_6031# 0.212f
C3852 _110_ _026_ 4.25e-20
C3853 net18 trim_mask\[0\] 0.0149f
C3854 a_5691_7637# a_5363_7369# 8.58e-19
C3855 _119_ a_10676_1679# 1.34e-21
C3856 a_12522_8751# VPWR 0.00343f
C3857 a_11343_3317# a_11967_3311# 9.73e-19
C3858 a_7939_10383# a_8215_9295# 1.62e-20
C3859 net22 a_2313_6183# 0.174f
C3860 a_10405_9295# a_10864_9269# 0.078f
C3861 net2 a_14422_7093# 9.13e-19
C3862 _028_ _027_ 0.00438f
C3863 a_2309_2229# clk 0.00965f
C3864 a_7723_10143# a_7548_10217# 0.234f
C3865 net18 a_10405_9295# 0.0121f
C3866 a_8657_2229# a_9572_2601# 0.125f
C3867 a_3947_11305# _042_ 0.00153f
C3868 a_2787_9845# a_3977_10217# 2.56e-19
C3869 _084_ _009_ 0.189f
C3870 a_763_8757# a_1844_9129# 0.102f
C3871 _108_ a_14335_2442# 0.188f
C3872 _106_ a_9003_3829# 0.00425f
C3873 a_10752_12533# net18 0.172f
C3874 mask\[1\] a_4043_7093# 9.46e-20
C3875 net33 a_14604_2339# 0.0158f
C3876 a_448_11445# result[6] 7.93e-20
C3877 _136_ net50 0.00145f
C3878 _101_ a_5691_7637# 0.0034f
C3879 _108_ net8 4.46e-19
C3880 a_763_8757# _006_ 0.169f
C3881 net44 a_5726_5807# 1.57e-19
C3882 a_1651_7093# a_2953_7119# 1.03e-19
C3883 a_1476_7119# a_2787_7119# 1.09e-19
C3884 a_5915_10927# a_6099_10633# 8.82e-20
C3885 mask\[0\] a_2787_7119# 0.23f
C3886 a_1007_10217# VPWR 7.41e-19
C3887 _067_ trim_mask\[4\] 6.2e-21
C3888 net2 _132_ 0.00922f
C3889 _096_ net3 0.027f
C3890 clknet_2_0__leaf_clk a_2564_2589# 0.017f
C3891 net9 a_12664_8029# 5.14e-19
C3892 _101_ a_5089_10159# 0.00145f
C3893 a_3748_6281# _095_ 4.78e-19
C3894 net33 net2 0.612f
C3895 net46 a_13257_4943# 0.595f
C3896 a_11067_4405# a_11691_4399# 9.73e-19
C3897 net39 net34 0.147f
C3898 cal_itt\[1\] a_9443_6059# 9.72e-19
C3899 a_1095_12393# a_1095_11305# 0.00139f
C3900 a_1660_12393# a_745_10933# 3.21e-21
C3901 a_4512_11305# a_4674_10927# 0.00645f
C3902 _060_ _100_ 0.312f
C3903 a_8298_5487# a_9503_4399# 4.03e-20
C3904 a_9296_9295# _070_ 2.47e-19
C3905 a_7524_2223# clk 0.00269f
C3906 _104_ a_10781_3311# 0.0322f
C3907 trim_mask\[0\] trim_val\[0\] 0.551f
C3908 _050_ a_7891_3617# 0.236f
C3909 a_4498_4373# state\[2\] 1.3e-19
C3910 state\[2\] a_4864_1679# 3.21e-21
C3911 calibrate _097_ 0.0132f
C3912 net15 a_3977_7119# 6.04e-20
C3913 a_3781_8207# a_4858_8573# 1.46e-19
C3914 a_3615_8207# a_4227_8207# 3.82e-19
C3915 en_co_clk a_5726_5807# 2.33e-19
C3916 _024_ a_11321_3855# 1.97e-19
C3917 net15 a_2877_2197# 0.0136f
C3918 a_15023_5487# a_15083_4659# 0.003f
C3919 a_4498_4373# state\[0\] 8.12e-19
C3920 clknet_2_2__leaf_clk trim_mask\[4\] 0.559f
C3921 _072_ a_7263_7093# 0.00214f
C3922 a_9003_3829# _033_ 0.00101f
C3923 net40 net5 1.96e-19
C3924 trim_val\[4\] a_8583_3317# 6.67e-19
C3925 _094_ net54 0.0691f
C3926 _081_ a_911_7119# 7.83e-20
C3927 _053_ a_10586_7371# 7.74e-19
C3928 a_3947_12393# _078_ 0.0015f
C3929 a_1476_10217# net25 0.0523f
C3930 _090_ a_3148_4399# 3.97e-19
C3931 _051_ _110_ 3.65e-20
C3932 clknet_2_3__leaf_clk a_11753_6031# 8.08e-19
C3933 _045_ a_6891_12393# 1.35e-19
C3934 clknet_2_1__leaf_clk a_8673_10625# 2.53e-19
C3935 _101_ a_6633_9845# 4.59e-21
C3936 _052_ a_7891_3617# 0.00112f
C3937 cal_itt\[0\] a_8307_6575# 2.61e-20
C3938 clknet_0_clk _051_ 1.46f
C3939 trim_mask\[1\] trim_val\[1\] 0.32f
C3940 _007_ net25 0.0825f
C3941 net16 a_13825_5185# 0.00716f
C3942 _093_ a_3530_4438# 1.07e-19
C3943 net14 a_1476_10217# 4.01e-19
C3944 mask\[3\] a_5177_9537# 0.0506f
C3945 a_3110_3311# clk 2.55e-20
C3946 _090_ a_3365_4943# 0.00432f
C3947 a_4993_6273# _092_ 1.3e-19
C3948 _091_ en_co_clk 0.00219f
C3949 net45 a_2479_3689# 5.93e-19
C3950 net31 _132_ 0.00487f
C3951 _074_ a_395_4405# 0.0275f
C3952 a_911_4777# a_855_4105# 0.00338f
C3953 _078_ a_3425_11721# 0.05f
C3954 net14 _007_ 7.62e-19
C3955 a_12516_2601# a_14335_2442# 2.03e-20
C3956 net45 a_8491_2229# 7.48e-21
C3957 a_1099_12533# net14 0.201f
C3958 trim_val\[2\] _114_ 0.0134f
C3959 _031_ a_12678_2223# 3.59e-20
C3960 clknet_2_0__leaf_clk net1 1.47e-19
C3961 net18 a_11258_8790# 7.07e-19
C3962 net43 a_8025_8041# 6.59e-20
C3963 _106_ a_8485_4943# 6.6e-20
C3964 net32 _055_ 0.0157f
C3965 net33 net31 0.485f
C3966 _024_ a_11435_2229# 1.74e-20
C3967 net12 a_7250_7485# 3.74e-20
C3968 _125_ a_13919_8751# 0.00216f
C3969 a_14983_9269# a_15023_8751# 9.59e-19
C3970 clknet_2_1__leaf_clk a_7164_11293# 8.22e-19
C3971 net15 _042_ 0.00595f
C3972 net3 a_5455_4943# 0.155f
C3973 _064_ a_9007_2601# 1.16e-21
C3974 _110_ a_10752_565# 4.1e-20
C3975 a_14099_3017# trim[0] 1.79e-19
C3976 _118_ trim_mask\[1\] 4.41e-20
C3977 _110_ _031_ 0.188f
C3978 net44 _040_ 0.284f
C3979 net22 VPWR 0.751f
C3980 _123_ a_12430_7663# 0.00221f
C3981 _065_ a_11491_6031# 0.00413f
C3982 a_2921_2589# VPWR 5.66e-20
C3983 _101_ a_6445_10383# 5.79e-19
C3984 _078_ _008_ 0.165f
C3985 mask\[4\] _000_ 3.63e-20
C3986 _035_ net2 4.55e-20
C3987 cal_count\[0\] a_13142_8359# 1.96e-20
C3988 _049_ a_5502_6397# 1.04e-19
C3989 trim_mask\[3\] _116_ 6.05e-19
C3990 a_3597_12021# a_3947_11305# 3.45e-20
C3991 a_7351_8041# a_7723_6807# 7.48e-19
C3992 a_3947_12393# a_3597_10933# 2.85e-21
C3993 a_4165_11989# a_4165_10901# 3.75e-20
C3994 trim_mask\[0\] a_11023_5108# 3.37e-21
C3995 net9 a_12824_7663# 3.42e-19
C3996 a_4609_1679# clk 0.546f
C3997 _050_ _087_ 6.6e-20
C3998 _088_ a_7190_3855# 0.0285f
C3999 mask\[6\] _084_ 0.0364f
C4000 a_13557_7369# _136_ 1.66e-20
C4001 a_9747_2527# a_10111_1679# 4.14e-19
C4002 a_10543_2455# a_9761_1679# 3.27e-19
C4003 _001_ a_12061_7669# 5.65e-20
C4004 net48 a_13091_1141# 0.00996f
C4005 cal_itt\[2\] a_8473_5193# 2.71e-19
C4006 a_7262_5461# a_7190_3855# 1.01e-20
C4007 a_11059_7356# a_11622_7485# 0.0498f
C4008 a_10990_7485# a_11204_7485# 0.0977f
C4009 a_10903_7261# a_13142_7271# 6.77e-20
C4010 net16 _122_ 0.0236f
C4011 a_4498_4373# _100_ 1.42e-20
C4012 a_2143_7663# a_2857_7637# 0.0172f
C4013 _065_ a_6419_8207# 0.00369f
C4014 _042_ a_4030_9839# 2.02e-19
C4015 _118_ a_8749_3317# 3.81e-21
C4016 _050_ _099_ 2.42e-19
C4017 _086_ a_1129_9813# 1.59e-22
C4018 _087_ _052_ 3.07e-19
C4019 net2 _136_ 0.0141f
C4020 _055_ VPWR 0.517f
C4021 _078_ a_5524_9295# 0.0161f
C4022 _101_ a_3411_9839# 8.49e-19
C4023 a_3133_11247# VPWR 3.06e-19
C4024 net43 a_1019_7485# 0.0122f
C4025 a_11801_4373# _110_ 1.61e-20
C4026 _052_ a_6519_3829# 0.0101f
C4027 _071_ a_8820_6005# 0.0776f
C4028 net4 a_7379_2197# 1.41e-19
C4029 _098_ _087_ 0.105f
C4030 net42 a_6316_5193# 3.84e-19
C4031 net44 _048_ 2e-20
C4032 net30 a_7571_4943# 1.1e-19
C4033 net41 a_1867_3317# 0.19f
C4034 net21 mask\[3\] 9.79e-21
C4035 a_1203_10927# a_911_10217# 3.01e-20
C4036 a_395_4405# _093_ 8.32e-20
C4037 _099_ _052_ 1.41e-19
C4038 trim_mask\[0\] a_7460_5807# 8.43e-21
C4039 _058_ a_11764_3677# 0.00115f
C4040 _065_ a_3529_6281# 2.4e-19
C4041 _062_ a_5515_6005# 4.43e-19
C4042 en_co_clk a_14655_4399# 6.91e-20
C4043 a_9463_8725# _070_ 1.46e-19
C4044 net14 a_1357_11293# 6.71e-19
C4045 net37 net49 1.62e-19
C4046 net14 a_2877_2197# 6.77e-20
C4047 a_2857_5461# a_4091_5309# 4.98e-19
C4048 _095_ a_4308_4917# 0.151f
C4049 _098_ _099_ 0.0998f
C4050 a_3868_10217# a_3840_8867# 5.65e-20
C4051 _074_ a_561_9845# 0.015f
C4052 net18 _042_ 0.169f
C4053 net47 a_11244_9661# 0.245f
C4054 _075_ a_7460_5807# 4.95e-20
C4055 a_10864_9269# a_11008_9295# 0.00196f
C4056 a_10688_9295# a_10798_9295# 0.00807f
C4057 a_11067_3017# a_11413_2767# 0.0134f
C4058 net40 net46 0.33f
C4059 a_14604_3017# a_14686_3017# 0.00477f
C4060 net52 a_2869_10927# 0.0474f
C4061 net4 a_9664_3689# 0.00131f
C4062 a_11801_4373# a_12148_4777# 0.0512f
C4063 _078_ sample 1.76e-19
C4064 net18 a_11008_9295# 4.63e-19
C4065 a_14983_9269# _126_ 0.194f
C4066 result[3] result[2] 0.037f
C4067 trim_val\[0\] _030_ 0.00101f
C4068 net47 a_11204_7485# 0.0122f
C4069 a_4165_10901# VPWR 0.207f
C4070 net43 a_1173_10205# 0.00368f
C4071 a_6541_12021# VPWR 0.574f
C4072 net12 _107_ 0.0371f
C4073 a_1467_7923# a_1125_7663# 7.26e-19
C4074 _048_ clk 0.137f
C4075 en_co_clk _048_ 0.0131f
C4076 a_395_4405# a_2865_4460# 2.24e-21
C4077 trim_mask\[0\] a_12691_2527# 5.88e-20
C4078 a_6515_6794# net30 0.0371f
C4079 _108_ a_13703_4943# 0.00129f
C4080 _010_ a_1660_12393# 1.93e-21
C4081 net53 a_4443_9295# 2.38e-20
C4082 _042_ net25 9.06e-19
C4083 a_4512_11305# a_4609_9295# 2.21e-19
C4084 _048_ a_9084_4515# 0.206f
C4085 net44 a_5177_9537# 0.186f
C4086 _059_ _089_ 0.0142f
C4087 _041_ a_12341_8751# 0.0194f
C4088 net41 a_3302_3677# 0.00184f
C4089 net47 _123_ 0.192f
C4090 a_12723_4943# clknet_2_2__leaf_clk 0.0215f
C4091 a_14931_591# trim[3] 7.28e-19
C4092 net15 a_3597_12021# 1.11e-19
C4093 net20 mask\[4\] 1.68e-22
C4094 net14 _042_ 1.65e-20
C4095 net12 _049_ 0.214f
C4096 _051_ net41 0.116f
C4097 _064_ a_10851_1653# 0.00209f
C4098 _118_ a_7939_3855# 1.86e-20
C4099 net45 a_395_6031# 0.298f
C4100 net12 a_5699_1653# 0.00577f
C4101 a_4259_6031# _050_ 1.51e-19
C4102 net55 a_8473_5193# 0.00126f
C4103 _014_ net41 0.00917f
C4104 a_4131_8207# net45 4.02e-20
C4105 a_12520_7637# cal_count\[2\] 1.56e-19
C4106 a_12900_7663# a_12924_8029# 0.0016f
C4107 _057_ ctln[3] 0.0412f
C4108 a_4871_6031# VPWR 2.44e-19
C4109 a_4471_4007# a_4617_3855# 0.0134f
C4110 trim_val\[2\] VPWR 0.557f
C4111 net43 a_6173_7119# 5.95e-20
C4112 _119_ trim_mask\[2\] 0.104f
C4113 net19 a_7565_12393# 3.38e-20
C4114 a_4801_9839# _040_ 4.45e-20
C4115 a_455_8181# net23 0.0138f
C4116 _076_ a_8301_8207# 6.01e-21
C4117 _096_ net54 0.376f
C4118 net34 a_14604_2339# 0.00256f
C4119 _049_ a_5340_6031# 0.0107f
C4120 _105_ _106_ 0.14f
C4121 a_11987_8757# net2 1.57e-19
C4122 _053_ _064_ 0.0826f
C4123 a_10111_1679# a_10676_1679# 7.99e-20
C4124 a_4775_6031# a_4498_4373# 5.02e-21
C4125 trim_mask\[1\] a_12424_3689# 0.049f
C4126 a_6428_7119# a_6619_7119# 4.61e-19
C4127 a_15023_12559# a_15023_12015# 0.0523f
C4128 a_3431_10933# mask\[2\] 1.68e-19
C4129 net11 _116_ 5.63e-20
C4130 a_13091_1141# a_14281_1513# 2.56e-19
C4131 cal_itt\[0\] VPWR 2.46f
C4132 trim_mask\[1\] a_14184_2767# 0.0103f
C4133 a_3840_8867# a_3922_8867# 0.00477f
C4134 cal_count\[3\] net50 0.0229f
C4135 a_6909_10933# a_7548_10217# 7.02e-21
C4136 a_7477_10901# a_7723_10143# 5.29e-20
C4137 net26 a_1764_10383# 0.00117f
C4138 net9 a_11601_2229# 0.0159f
C4139 a_13607_1513# trim[3] 2.57e-20
C4140 clknet_2_1__leaf_clk a_2961_9545# 0.00436f
C4141 a_14172_4943# trim[4] 5.6e-19
C4142 a_2309_2229# a_3399_2527# 0.0418f
C4143 a_2143_2229# a_3224_2601# 0.102f
C4144 a_2877_2197# a_2659_2601# 0.21f
C4145 _067_ a_8761_7983# 2.18e-20
C4146 _108_ a_13459_3317# 0.00562f
C4147 net17 net9 0.111f
C4148 net34 net2 0.0237f
C4149 a_15259_7637# VPWR 0.407f
C4150 clknet_2_2__leaf_clk a_11967_3311# 0.00165f
C4151 clknet_2_1__leaf_clk a_448_9269# 0.0196f
C4152 a_1095_11305# a_1461_10357# 0.00344f
C4153 clknet_2_3__leaf_clk a_8731_9295# 0.0335f
C4154 _076_ _094_ 5.86e-20
C4155 net27 a_4165_10901# 3.28e-20
C4156 net46 _024_ 0.0203f
C4157 a_6541_12021# net27 2.95e-19
C4158 net44 a_7810_12381# 0.00288f
C4159 a_7109_11989# a_6999_12015# 0.0977f
C4160 clknet_2_1__leaf_clk a_1660_11305# 0.00135f
C4161 net29 a_2910_12131# 2.03e-19
C4162 mask\[7\] net26 0.0661f
C4163 clknet_2_1__leaf_clk mask\[0\] 1.88e-19
C4164 clknet_2_3__leaf_clk _037_ 0.0387f
C4165 clknet_2_2__leaf_clk a_13059_4631# 0.0181f
C4166 _074_ a_2283_4020# 1.47e-21
C4167 a_3116_12533# VPWR 0.242f
C4168 a_9664_3689# a_11509_3317# 2.05e-20
C4169 _125_ cal_count\[2\] 2.52e-20
C4170 _108_ _109_ 0.00222f
C4171 net14 a_1476_6031# 0.00335f
C4172 _119_ a_9719_1473# 6.99e-22
C4173 net21 a_4687_11231# 0.0015f
C4174 a_8820_6005# a_9043_6031# 0.0115f
C4175 _048_ _059_ 0.0919f
C4176 _095_ _090_ 0.132f
C4177 net9 a_12061_7669# 0.0212f
C4178 _105_ _033_ 1.58e-21
C4179 net4 a_9919_6614# 2.01e-19
C4180 a_13625_3317# a_14702_3311# 1.46e-19
C4181 a_6210_4989# net42 1.79e-19
C4182 _072_ _071_ 0.0822f
C4183 state\[0\] a_4576_3427# 0.167f
C4184 a_7310_2223# a_7617_2589# 3.69e-19
C4185 a_7184_2339# a_7942_2223# 0.0612f
C4186 a_7379_2197# a_7689_2589# 0.0138f
C4187 _008_ a_6888_10205# 0.158f
C4188 a_7569_7637# VPWR 0.22f
C4189 a_6467_9845# a_7079_10217# 3.82e-19
C4190 net13 a_5515_6005# 2.47e-19
C4191 net16 comp 3e-20
C4192 net47 a_13142_8725# 0.116f
C4193 net37 a_15159_9269# 3.35e-19
C4194 clknet_2_3__leaf_clk a_12231_6005# 0.0722f
C4195 a_9503_4399# a_9839_3615# 1.04e-19
C4196 _074_ a_5496_12131# 0.0534f
C4197 _068_ _071_ 0.319f
C4198 _074_ _006_ 0.274f
C4199 net12 _008_ 0.00728f
C4200 a_8307_6575# a_8307_4943# 2.9e-21
C4201 a_4308_4917# calibrate 2.36e-20
C4202 _108_ trim[2] 4.34e-20
C4203 a_4165_11989# a_4043_12393# 3.16e-19
C4204 net45 net30 0.0259f
C4205 a_3947_12393# a_3852_12381# 0.0498f
C4206 a_7715_3285# a_8583_3317# 3.37e-21
C4207 mask\[3\] a_2143_7663# 1.03e-19
C4208 net10 ctln[4] 0.0067f
C4209 mask\[1\] a_6056_8359# 3.42e-19
C4210 net43 a_3852_11293# 0.00323f
C4211 net34 net31 0.966f
C4212 a_12900_7663# a_13008_7663# 0.00523f
C4213 a_395_7119# a_1476_6031# 4.25e-21
C4214 _132_ a_14733_7983# 0.0018f
C4215 a_7079_10217# VPWR 2.33e-19
C4216 a_8298_2767# a_10055_2767# 0.0029f
C4217 net30 _058_ 0.00133f
C4218 _096_ a_4471_4007# 0.0924f
C4219 _103_ _088_ 0.121f
C4220 clknet_2_1__leaf_clk a_6197_12015# 0.00422f
C4221 _119_ a_9595_1679# 1.68e-19
C4222 _049_ a_6197_6281# 0.00121f
C4223 a_1497_8725# net24 0.0191f
C4224 a_1279_9129# a_1844_9129# 7.99e-20
C4225 trim_mask\[1\] a_11435_2229# 8.3e-22
C4226 a_7262_5461# _103_ 1.28e-19
C4227 _050_ a_7393_5193# 1.84e-20
C4228 a_1129_6273# result[0] 5.27e-19
C4229 _004_ sample 0.0175f
C4230 net14 net6 0.0991f
C4231 clknet_2_3__leaf_clk a_13697_4373# 3.16e-21
C4232 a_13092_8029# VPWR 9.06e-20
C4233 a_14334_1135# trim[3] 1.63e-20
C4234 _006_ a_1279_9129# 5.1e-19
C4235 a_8491_2229# a_8657_2229# 0.614f
C4236 a_455_3571# a_395_2767# 0.0101f
C4237 net9 a_14172_1513# 2.52e-20
C4238 _008_ a_6983_10217# 5.01e-19
C4239 a_6467_9845# a_7723_10143# 0.0436f
C4240 trim_mask\[0\] VPWR 3.23f
C4241 net19 _051_ 7.23e-20
C4242 net12 a_5524_9295# 0.00241f
C4243 _091_ _108_ 3.2e-20
C4244 a_11067_4405# _025_ 5.29e-19
C4245 net46 a_13703_1513# 0.00418f
C4246 _024_ a_11343_3317# 0.00115f
C4247 a_7723_6807# a_8307_6575# 0.0134f
C4248 a_9296_9295# net2 4.77e-21
C4249 net14 a_1137_11721# 5.22e-19
C4250 _024_ a_11149_3017# 6.81e-20
C4251 a_11067_4405# _026_ 2.01e-20
C4252 net44 _020_ 0.0153f
C4253 _092_ net3 0.0901f
C4254 mask\[2\] clknet_2_0__leaf_clk 8.35e-19
C4255 _075_ VPWR 0.573f
C4256 a_10405_9295# VPWR 0.273f
C4257 net43 a_3947_11305# 0.164f
C4258 a_995_3530# cal 0.196f
C4259 net55 a_7190_3855# 1.88e-19
C4260 _103_ a_6519_4631# 7.62e-20
C4261 net20 a_6987_12393# 0.00117f
C4262 a_6885_8372# net51 0.111f
C4263 a_745_10933# a_1095_11305# 0.23f
C4264 a_7723_10143# VPWR 0.362f
C4265 net47 a_14565_9295# 1.21e-20
C4266 trim_val\[0\] a_15083_4659# 0.00905f
C4267 a_10752_12533# VPWR 0.291f
C4268 a_10975_6031# _038_ 0.218f
C4269 a_2033_3317# clk 6.05e-19
C4270 a_7210_5807# a_7460_5807# 0.097f
C4271 _093_ a_2283_4020# 0.0377f
C4272 a_9839_3615# a_9747_2527# 7.1e-20
C4273 _074_ result[7] 1.76e-20
C4274 _098_ a_7393_5193# 0.002f
C4275 a_6631_7485# _049_ 5.46e-20
C4276 trim_mask\[3\] a_11601_2229# 0.003f
C4277 net46 _029_ 0.0415f
C4278 a_12153_8757# a_12344_8041# 3.29e-21
C4279 a_12436_9129# a_12061_7669# 5.41e-19
C4280 a_10699_3311# a_9761_1679# 3.18e-22
C4281 a_14540_3689# _056_ 1.92e-19
C4282 cal_count\[3\] _106_ 0.00111f
C4283 a_8215_9295# _070_ 8.05e-20
C4284 net16 a_13111_6031# 2.14e-19
C4285 _065_ net40 1.05e-19
C4286 clknet_2_2__leaf_clk a_13257_4943# 0.00303f
C4287 _107_ a_5691_2741# 1.77e-19
C4288 _062_ a_9443_6059# 0.00845f
C4289 net2 a_15299_6575# 9.38e-19
C4290 net12 trim_mask\[4\] 0.0958f
C4291 a_13933_6281# VPWR 0.00924f
C4292 _125_ cal_count\[1\] 0.0748f
C4293 a_1476_10217# VPWR 0.286f
C4294 net2 cal_count\[3\] 0.29f
C4295 net13 mask\[2\] 0.0636f
C4296 net26 a_8105_10383# 0.00549f
C4297 mask\[3\] _077_ 6.46e-21
C4298 _134_ _058_ 4.45e-19
C4299 net4 _124_ 0.00181f
C4300 net50 _119_ 0.00107f
C4301 net28 a_2910_12131# 3.76e-19
C4302 _054_ a_7010_3311# 0.00149f
C4303 a_7800_4631# a_8307_4719# 2.21e-19
C4304 clknet_2_0__leaf_clk a_6428_7119# 1.99e-19
C4305 _007_ VPWR 0.791f
C4306 trim_mask\[0\] a_9478_4105# 0.0551f
C4307 a_1099_12533# VPWR 0.432f
C4308 clknet_2_0__leaf_clk a_2143_2229# 0.323f
C4309 a_4030_7485# VPWR 7.67e-19
C4310 net14 a_1357_12381# 6.71e-19
C4311 _074_ a_911_4777# 0.016f
C4312 a_8717_10383# VPWR 3.81e-19
C4313 a_2953_7119# net30 9.05e-20
C4314 clknet_2_1__leaf_clk a_6099_10633# 0.058f
C4315 trim_val\[4\] a_9662_3855# 0.00235f
C4316 a_13975_3689# a_14071_3689# 0.0138f
C4317 a_2491_3311# clk 1.11e-19
C4318 cal_itt\[0\] a_9650_9295# 5.1e-19
C4319 net2 a_14981_8235# 0.00219f
C4320 a_13869_4943# VPWR 0.00186f
C4321 _013_ a_1201_3855# 5.79e-20
C4322 a_11601_2229# a_13415_2442# 1.35e-19
C4323 a_12169_2197# a_12516_2601# 0.0512f
C4324 net22 a_2476_6281# 1.11e-20
C4325 net53 _065_ 1.47e-19
C4326 net29 a_2787_10927# 5.81e-21
C4327 net21 a_4801_9839# 2.6e-21
C4328 net45 state\[2\] 0.0716f
C4329 net47 a_14335_7895# 1.21e-19
C4330 net35 a_14540_3689# 3.91e-20
C4331 net32 _030_ 3.33e-21
C4332 _058_ a_13975_3689# 0.00144f
C4333 net40 a_11233_4405# 2.47e-20
C4334 _049_ a_5726_5807# 2.08e-19
C4335 _091_ _107_ 0.00135f
C4336 _090_ calibrate 0.0169f
C4337 a_14485_7663# VPWR 0.00559f
C4338 net43 _005_ 9e-19
C4339 a_13142_8359# cal_count\[2\] 1.5e-19
C4340 clknet_2_3__leaf_clk a_13825_5185# 1.75e-20
C4341 net45 state\[0\] 0.00525f
C4342 net15 _039_ 8.96e-21
C4343 _108_ a_14655_4399# 0.00233f
C4344 mask\[0\] a_6007_7119# 4.4e-20
C4345 _101_ a_4443_9295# 0.0181f
C4346 a_4425_6031# a_5081_4943# 6.67e-21
C4347 a_15023_2767# trim[0] 0.337f
C4348 a_11258_8790# VPWR 0.00203f
C4349 net31 a_15299_6575# 0.00676f
C4350 a_8949_6281# VPWR 0.191f
C4351 net27 a_7723_10143# 2.42e-19
C4352 a_7723_6807# a_7897_6913# 0.00658f
C4353 _085_ net13 6.8e-21
C4354 net15 net43 0.0355f
C4355 a_561_7119# a_1585_7119# 2.36e-20
C4356 a_14983_9269# VPWR 0.166f
C4357 trim_mask\[2\] a_11292_1251# 4.08e-20
C4358 a_4425_6031# net55 1.84e-19
C4359 _048_ a_3399_2527# 1.69e-19
C4360 _058_ a_13915_4399# 0.00973f
C4361 net52 _101_ 0.874f
C4362 mask\[2\] a_4864_9295# 0.00264f
C4363 _048_ _108_ 0.00102f
C4364 a_561_9845# a_2450_9955# 1.9e-20
C4365 net16 a_13825_6031# 0.00322f
C4366 _107_ _089_ 0.00335f
C4367 net3 cal 0.00534f
C4368 _027_ a_9761_1679# 9.9e-20
C4369 _064_ a_9664_3689# 1.31e-19
C4370 net14 a_937_3855# 9.7e-20
C4371 a_6909_10933# a_7933_11305# 2.36e-20
C4372 a_7477_10901# a_7521_11293# 3.69e-19
C4373 _056_ net8 0.00123f
C4374 a_395_9845# a_3208_10205# 6.41e-22
C4375 a_8731_9295# a_8827_9295# 0.0138f
C4376 a_8381_9295# cal_itt\[0\] 3.26e-19
C4377 a_8949_9537# a_8993_9295# 3.69e-19
C4378 net13 a_4815_3031# 0.0132f
C4379 net30 a_2857_5461# 0.0321f
C4380 a_3852_11293# a_2953_9845# 6.78e-20
C4381 net43 a_7351_8041# 0.187f
C4382 a_763_8757# _080_ 5.04e-20
C4383 _087_ a_6519_3829# 0.0111f
C4384 _065_ _024_ 3.21e-19
C4385 _015_ a_4709_2773# 0.00193f
C4386 _042_ _019_ 7.08e-19
C4387 _092_ a_11709_6273# 1.29e-21
C4388 a_8083_8181# cal_itt\[3\] 4.21e-22
C4389 _034_ a_4680_6031# 0.157f
C4390 mask\[0\] _092_ 2e-19
C4391 a_9463_8725# net2 5.94e-20
C4392 _064_ a_10689_2223# 0.0116f
C4393 _110_ trim_val\[2\] 2.39e-19
C4394 net27 _007_ 2.83e-20
C4395 a_3977_7119# VPWR 4.45e-20
C4396 _087_ _099_ 0.153f
C4397 _030_ VPWR 0.405f
C4398 a_455_12533# a_448_11445# 0.00249f
C4399 a_1099_12533# net27 2.42e-20
C4400 a_8022_7119# net30 0.00164f
C4401 _066_ a_10137_4943# 3.47e-20
C4402 a_911_4777# _093_ 1.44e-19
C4403 a_448_9269# result[4] 0.0022f
C4404 _053_ a_7379_2197# 1.42e-21
C4405 _049_ _089_ 0.00246f
C4406 a_4308_4917# _015_ 3.58e-20
C4407 a_1357_11293# VPWR 6.77e-19
C4408 a_2877_2197# VPWR 0.216f
C4409 a_12520_7637# a_12900_7663# 0.00971f
C4410 a_12061_7669# a_13470_7663# 4.25e-19
C4411 net40 _067_ 3.32e-19
C4412 clknet_2_2__leaf_clk a_6941_2589# 3.64e-20
C4413 a_1651_6005# _049_ 1.66e-19
C4414 a_1476_6031# a_2313_6183# 3.43e-19
C4415 a_11059_7356# _136_ 0.00126f
C4416 _134_ a_13607_4943# 1.86e-19
C4417 clknet_2_3__leaf_clk _122_ 0.15f
C4418 a_8307_4943# VPWR 0.222f
C4419 _011_ a_579_10933# 1.73e-19
C4420 trim_mask\[0\] _104_ 0.348f
C4421 net45 a_1585_6031# 6.92e-19
C4422 mask\[6\] a_7164_11293# 2.48e-21
C4423 a_1313_10901# result[5] 9.44e-20
C4424 comp clkc 0.0375f
C4425 result[1] result[0] 0.0489f
C4426 a_395_4405# a_3057_4719# 1.52e-21
C4427 _045_ net53 1.02e-19
C4428 a_5177_1921# a_4959_1679# 0.21f
C4429 a_4443_1679# a_5524_1679# 0.102f
C4430 a_4609_1679# a_5699_1653# 0.0424f
C4431 a_10689_2223# a_10851_1653# 3.4e-19
C4432 a_6173_7119# a_6741_7361# 0.186f
C4433 a_3597_10933# a_3303_10217# 8.89e-21
C4434 clknet_2_3__leaf_clk _063_ 0.0185f
C4435 cal_itt\[0\] clknet_0_clk 0.00304f
C4436 a_6909_10933# a_7477_10901# 0.186f
C4437 net9 _025_ 9.33e-19
C4438 _042_ a_6467_9845# 3.4e-21
C4439 _064_ a_10781_3631# 0.00489f
C4440 net46 trim_mask\[1\] 0.046f
C4441 a_10699_3311# a_11067_3017# 8.59e-20
C4442 net9 _026_ 0.0184f
C4443 a_15299_3311# trim[0] 2.73e-19
C4444 net47 a_10239_9295# 0.101f
C4445 a_15023_8751# _129_ 2.28e-19
C4446 _040_ _049_ 2.28e-19
C4447 a_8298_2767# VPWR 1.25f
C4448 net13 a_4674_10927# 1.29e-19
C4449 net52 _102_ 0.17f
C4450 a_14063_7093# a_14282_7119# 0.0105f
C4451 net4 a_8583_3317# 0.00723f
C4452 a_11067_4405# a_11801_4373# 0.0701f
C4453 _024_ a_11233_4405# 0.303f
C4454 _106_ _119_ 0.00412f
C4455 _136_ a_12257_4777# 7.17e-20
C4456 net44 _077_ 0.00501f
C4457 clknet_2_0__leaf_clk a_4443_1679# 0.248f
C4458 net16 a_14199_7369# 0.00289f
C4459 a_14172_4943# a_13625_3317# 1.42e-21
C4460 net40 clknet_2_2__leaf_clk 0.0226f
C4461 a_9681_2601# VPWR 8.79e-20
C4462 clknet_2_0__leaf_clk a_1476_4777# 0.016f
C4463 _042_ VPWR 6.5f
C4464 a_7723_6807# VPWR 0.222f
C4465 _078_ a_2006_8751# 9.62e-20
C4466 _065_ _071_ 6.44e-20
C4467 cal_count\[1\] a_13142_8359# 0.00316f
C4468 mask\[2\] a_4239_8573# 4.21e-20
C4469 _053_ a_11425_5487# 1.93e-19
C4470 net15 a_2857_7637# 0.11f
C4471 a_7210_5807# VPWR 0.00334f
C4472 net28 a_2787_10927# 0.00115f
C4473 _108_ trim[1] 3.27e-19
C4474 a_10543_2455# trim_val\[3\] 7.23e-21
C4475 _048_ _107_ 0.176f
C4476 _074_ mask\[7\] 0.156f
C4477 net29 a_3947_12393# 1.85e-22
C4478 net45 a_911_6031# 0.153f
C4479 a_10329_1921# a_10195_1354# 7.23e-19
C4480 _031_ a_13512_1501# 0.156f
C4481 a_9761_1679# _117_ 8.94e-20
C4482 _032_ a_10569_1109# 6.04e-19
C4483 net46 a_8749_3317# 0.0247f
C4484 _126_ a_14236_8457# 0.106f
C4485 a_14983_9269# a_14807_8359# 1.16e-19
C4486 net43 a_1822_12015# 3.18e-19
C4487 net13 a_5087_3855# 0.00466f
C4488 clknet_2_1__leaf_clk a_2489_7983# 1.69e-19
C4489 a_13607_4943# a_13915_4399# 9.16e-20
C4490 a_1677_9545# a_763_8757# 2.65e-20
C4491 net14 _039_ 0.00319f
C4492 net52 _022_ 0.00375f
C4493 net43 net25 0.261f
C4494 a_10864_7387# a_11369_7119# 2.28e-19
C4495 net16 a_12992_8751# 0.00115f
C4496 a_9020_10383# a_9182_10749# 0.00645f
C4497 a_8455_10383# a_8717_10383# 0.00171f
C4498 a_5363_12559# clknet_2_1__leaf_clk 7.72e-20
C4499 net13 a_4443_1679# 0.0199f
C4500 net55 _103_ 0.0766f
C4501 a_4658_3427# VPWR 0.00214f
C4502 a_11895_7669# a_12924_8029# 0.00248f
C4503 a_3513_12809# ctlp[1] 8.48e-19
C4504 net45 _012_ 6.1e-19
C4505 _092_ net54 0.204f
C4506 net33 trimb[1] 6.99e-19
C4507 net9 a_11168_9661# 1.21e-19
C4508 a_2092_8457# a_2971_8457# 7.2e-21
C4509 net14 net43 2.29f
C4510 a_11951_2601# VPWR 0.229f
C4511 a_7521_11293# VPWR 4.08e-19
C4512 net43 a_3399_7119# 4.36e-19
C4513 a_3748_6281# _050_ 1.25e-19
C4514 _049_ _048_ 0.598f
C4515 a_763_8757# a_1651_7093# 6.42e-21
C4516 _119_ _033_ 0.728f
C4517 _006_ a_911_7119# 8.48e-20
C4518 mask\[7\] a_1279_9129# 8.38e-21
C4519 _048_ a_3388_4631# 0.0676f
C4520 a_1276_565# clk 0.00421f
C4521 net45 a_5691_7637# 3.93e-19
C4522 a_9478_4105# a_8298_2767# 6.65e-21
C4523 a_3431_12021# a_3947_12393# 0.106f
C4524 a_3597_12021# a_4165_11989# 0.176f
C4525 clknet_2_1__leaf_clk _076_ 0.0855f
C4526 a_855_4105# a_937_4105# 0.171f
C4527 a_4259_6031# _099_ 8.76e-22
C4528 _120_ a_3817_4697# 0.00182f
C4529 a_9595_1679# a_10111_1679# 0.113f
C4530 _032_ a_10329_1921# 2.11e-19
C4531 _058_ trim_val\[1\] 7.73e-19
C4532 trim_mask\[1\] a_11343_3317# 0.0506f
C4533 a_13091_1141# _057_ 9.67e-20
C4534 _117_ a_10787_1135# 2.22e-19
C4535 cal valid 0.0947f
C4536 net26 a_9074_9955# 1.05e-19
C4537 a_448_10357# a_448_9269# 5.69e-19
C4538 trim_mask\[0\] _110_ 0.0683f
C4539 _095_ a_3667_3829# 5.12e-19
C4540 a_15299_3311# a_15023_2767# 0.00944f
C4541 net46 a_9361_3677# 0.0019f
C4542 a_3431_12021# a_3425_11721# 2.2e-19
C4543 _065_ a_11204_7485# 9.08e-20
C4544 a_1835_11231# net26 2.13e-20
C4545 clknet_0_clk trim_mask\[0\] 0.00637f
C4546 net43 a_395_7119# 0.313f
C4547 en_co_clk a_10975_6031# 2.39e-19
C4548 net46 _115_ 0.241f
C4549 _128_ a_13256_9117# 3.98e-19
C4550 a_15083_4659# net32 0.237f
C4551 a_7569_7637# a_7459_7663# 0.0977f
C4552 net15 a_2953_9845# 0.0117f
C4553 _034_ a_4425_6031# 0.293f
C4554 a_12344_8041# VPWR 0.296f
C4555 a_1476_6031# VPWR 0.298f
C4556 _090_ _015_ 6.44e-20
C4557 clknet_2_0__leaf_clk _120_ 0.0431f
C4558 trim_mask\[0\] a_12778_3677# 8.3e-20
C4559 _126_ _129_ 0.0109f
C4560 clknet_0_clk _075_ 0.261f
C4561 a_5177_1921# VPWR 0.217f
C4562 net47 a_10621_7119# 0.00288f
C4563 _009_ a_6197_12015# 0.0113f
C4564 net50 a_11292_1251# 8.75e-19
C4565 clknet_2_1__leaf_clk a_579_10933# 0.397f
C4566 a_6909_10933# VPWR 0.6f
C4567 net27 _042_ 9.12e-20
C4568 net29 a_2014_12381# 4.31e-19
C4569 _118_ _058_ 0.00858f
C4570 clknet_2_2__leaf_clk _024_ 0.153f
C4571 trim_mask\[0\] a_10699_5487# 4.91e-21
C4572 _078_ a_1493_5487# 0.0496f
C4573 a_3615_8207# a_6056_8359# 3.03e-21
C4574 trim_mask\[0\] a_12148_4777# 0.00583f
C4575 _065_ _123_ 0.0142f
C4576 _130_ trim[4] 2.59e-20
C4577 trim_mask\[2\] a_14604_3017# 1.33e-19
C4578 a_3123_3615# a_2309_2229# 1.12e-20
C4579 net45 a_4775_6031# 3.42e-20
C4580 a_2948_3689# a_2143_2229# 1.69e-20
C4581 _064_ a_10245_5193# 5.72e-19
C4582 mask\[1\] a_1211_7983# 0.00963f
C4583 cal_itt\[2\] a_9889_6873# 3.68e-21
C4584 trim_mask\[3\] _026_ 0.00645f
C4585 _068_ a_8935_6895# 0.0412f
C4586 net44 a_6173_7119# 0.0299f
C4587 a_10043_7983# a_9957_7663# 2.42e-19
C4588 _100_ a_4905_3855# 4.58e-19
C4589 _113_ a_13975_3689# 3.51e-20
C4590 a_579_12021# _078_ 9.87e-19
C4591 _065_ a_5363_7369# 0.0937f
C4592 mask\[5\] a_7933_11305# 1.52e-19
C4593 a_11016_6691# _136_ 0.00218f
C4594 net9 _031_ 7.5e-19
C4595 a_2953_9845# a_4030_9839# 1.46e-19
C4596 _092_ a_7019_4407# 1.19e-19
C4597 a_4655_10071# a_4801_10159# 0.0134f
C4598 trimb[2] trimb[0] 0.0503f
C4599 _107_ a_7021_4105# 0.00161f
C4600 net18 a_12323_4703# 2.81e-19
C4601 net47 a_11545_9049# 0.0104f
C4602 _108_ _112_ 0.00294f
C4603 a_3597_12021# VPWR 0.593f
C4604 _071_ _067_ 0.0665f
C4605 _102_ a_1679_10633# 0.0476f
C4606 net43 a_4222_7119# 0.00223f
C4607 net16 a_14422_7093# 0.00306f
C4608 a_8307_4943# _104_ 8.47e-20
C4609 net50 a_10111_1679# 0.00214f
C4610 net6 VPWR 0.495f
C4611 mask\[1\] a_4349_8449# 0.0192f
C4612 _054_ _119_ 0.00224f
C4613 net43 a_1769_11305# 6.03e-19
C4614 _101_ _065_ 0.722f
C4615 net4 net7 0.0774f
C4616 a_15083_4659# VPWR 0.499f
C4617 a_13050_7637# _133_ 9.84e-20
C4618 clknet_0_clk a_4030_7485# 9.87e-20
C4619 a_1276_565# ctln[0] 0.156f
C4620 net28 a_3947_12393# 0.0358f
C4621 mask\[6\] a_2961_9545# 5.16e-21
C4622 a_10016_1679# a_10207_1679# 4.61e-19
C4623 a_1137_11721# VPWR 0.00508f
C4624 a_3830_6281# a_4425_6031# 1.24e-19
C4625 a_7891_3617# a_7942_2223# 2.27e-21
C4626 _094_ a_5515_6005# 6.51e-19
C4627 _101_ net23 0.0393f
C4628 _049_ a_7021_4105# 0.0588f
C4629 a_6173_7119# clk 2.25e-19
C4630 a_561_4405# valid 0.00582f
C4631 _104_ a_8298_2767# 0.0012f
C4632 net16 _132_ 4.18e-20
C4633 _019_ a_4959_9295# 3.53e-19
C4634 mask\[6\] a_1660_11305# 6.58e-20
C4635 a_3852_11293# a_4043_11305# 4.61e-19
C4636 a_7223_2465# a_8491_2229# 0.0967f
C4637 a_7184_2339# a_7310_2223# 0.18f
C4638 net28 a_3425_11721# 0.00758f
C4639 mask\[5\] a_7477_10901# 2.14e-19
C4640 net13 a_4609_9295# 0.0153f
C4641 a_9195_10357# a_9871_10383# 2.18e-19
C4642 a_8455_10383# _042_ 0.0296f
C4643 net16 net33 0.11f
C4644 net42 _088_ 0.00164f
C4645 _014_ a_3224_2601# 5.47e-21
C4646 _009_ a_6099_10633# 4.03e-20
C4647 net47 _043_ 0.0686f
C4648 a_5633_1679# VPWR 2.19e-19
C4649 clknet_2_1__leaf_clk a_395_9845# 0.324f
C4650 _041_ _070_ 6.58e-20
C4651 a_7262_5461# net42 1.7e-19
C4652 _050_ a_4709_2773# 3.88e-20
C4653 net27 a_6909_10933# 2.33e-19
C4654 _078_ net53 0.229f
C4655 a_10005_6031# a_9503_4399# 3.44e-21
C4656 _076_ a_6485_8181# 0.254f
C4657 trim_val\[0\] a_12323_4703# 2.3e-20
C4658 a_6793_8970# net51 3.53e-19
C4659 a_13142_8359# a_12900_7663# 6.61e-19
C4660 a_8827_9295# _063_ 3.94e-20
C4661 _050_ a_4308_4917# 8.37e-19
C4662 _051_ a_4863_4917# 1.18e-20
C4663 net25 a_2953_9845# 6.82e-20
C4664 net3 a_4266_4943# 9.36e-19
C4665 a_3947_12393# a_4167_11471# 9.58e-20
C4666 a_13625_3317# net48 4.16e-21
C4667 a_4043_7093# a_4259_6031# 1.4e-19
C4668 a_3947_11305# a_4043_11305# 0.0138f
C4669 a_3333_2601# clk 5.25e-20
C4670 _029_ clknet_2_2__leaf_clk 0.0802f
C4671 cal_count\[1\] a_13557_8457# 0.00124f
C4672 a_1357_12381# VPWR 2.69e-19
C4673 net19 a_6541_12021# 4.79e-20
C4674 net15 mask\[3\] 0.00596f
C4675 _027_ a_11856_2589# 2e-20
C4676 _101_ a_2225_7663# 0.0116f
C4677 _079_ a_561_4405# 7.45e-20
C4678 trim_mask\[0\] a_13091_4943# 0.00555f
C4679 _111_ a_13233_4737# 7.45e-19
C4680 net46 a_10373_1679# 0.00447f
C4681 a_395_9845# a_2368_9955# 4.56e-21
C4682 _062_ _051_ 0.0941f
C4683 _124_ _053_ 1.67e-20
C4684 _040_ a_4036_8207# 0.0214f
C4685 a_9529_6059# VPWR 1.91e-19
C4686 _101_ _016_ 0.0162f
C4687 _060_ state\[1\] 0.0926f
C4688 _126_ a_14318_8457# 4.96e-19
C4689 calibrate a_3667_3829# 0.0444f
C4690 a_9839_3615# trim_mask\[2\] 0.00755f
C4691 a_3597_12021# net27 5.06e-22
C4692 _131_ a_15289_7119# 7.51e-19
C4693 a_4959_9295# VPWR 0.197f
C4694 net18 _038_ 0.0268f
C4695 _123_ _067_ 5.69e-19
C4696 _107_ a_7758_4759# 9.57e-20
C4697 net54 a_5536_4399# 0.00361f
C4698 net28 a_2014_12381# 7.77e-20
C4699 _110_ _030_ 0.00981f
C4700 a_11059_7356# cal_count\[3\] 3.03e-21
C4701 net34 a_14931_591# 0.12f
C4702 _048_ trim_mask\[4\] 2.84e-20
C4703 _045_ _101_ 7.28e-21
C4704 _076_ a_6007_7119# 0.0196f
C4705 clknet_2_3__leaf_clk a_13111_6031# 0.0435f
C4706 _042_ a_8381_9295# 2.78e-21
C4707 a_6835_7669# a_7088_7119# 1.65e-19
C4708 a_7001_7669# a_7263_7093# 0.00444f
C4709 trim_mask\[1\] a_9826_3311# 1.19e-20
C4710 trim_mask\[3\] a_10752_565# 0.0104f
C4711 a_4609_9295# a_4864_9295# 0.0594f
C4712 a_4443_9295# a_5067_9661# 9.73e-19
C4713 a_5177_9537# a_5524_9295# 0.0512f
C4714 a_7010_3631# a_6927_3311# 2.43e-19
C4715 _065_ _060_ 5.79e-21
C4716 net21 a_3947_12393# 0.00136f
C4717 _046_ net52 1.65e-19
C4718 clknet_0_clk a_8307_4943# 0.00311f
C4719 a_8298_5487# _106_ 0.00664f
C4720 net47 a_9471_9269# 0.344f
C4721 a_7939_10383# a_8839_9661# 4.77e-20
C4722 a_10864_9269# cal_count\[0\] 2.2e-20
C4723 a_4165_10901# a_4512_11305# 0.0512f
C4724 _101_ a_4696_8207# 1.13e-19
C4725 cal_count\[0\] a_15023_8751# 3.06e-19
C4726 a_6835_7669# _063_ 4.88e-21
C4727 net18 cal_count\[0\] 0.00559f
C4728 _039_ a_2313_6183# 0.106f
C4729 a_4043_10143# mask\[2\] 0.062f
C4730 a_11709_6273# _136_ 0.00384f
C4731 _049_ a_7758_4759# 1.28e-19
C4732 _038_ a_12165_6031# 1.94e-20
C4733 a_11233_4405# trim_mask\[1\] 9.96e-21
C4734 _129_ a_13050_7637# 5.56e-20
C4735 a_7109_11989# net44 0.17f
C4736 net16 ctlp[2] 0.00725f
C4737 _011_ result[6] 0.0016f
C4738 _058_ a_12424_3689# 0.00215f
C4739 a_3303_7119# a_3868_7119# 7.99e-20
C4740 a_2953_7119# a_3411_7485# 0.0346f
C4741 a_1313_10901# a_561_9845# 6.88e-21
C4742 _056_ trim[2] 0.00662f
C4743 clknet_2_0__leaf_clk a_1867_3317# 0.268f
C4744 _074_ _080_ 0.235f
C4745 a_14379_6397# trim_val\[0\] 9.02e-21
C4746 net21 a_3425_11721# 4.04e-19
C4747 _110_ a_8298_2767# 0.0083f
C4748 _133_ VPWR 1.11f
C4749 net12 a_7263_7093# 0.00158f
C4750 a_9369_4105# VPWR 0.0647f
C4751 a_7259_11305# _020_ 7.24e-20
C4752 clknet_0_clk a_8298_2767# 0.326f
C4753 net9 a_12522_8751# 4.34e-19
C4754 _050_ a_7310_2223# 0.00234f
C4755 _108_ a_11583_4777# 5.7e-19
C4756 _076_ _092_ 4.94e-20
C4757 a_7019_4407# a_6737_4719# 0.0382f
C4758 a_8749_3317# a_9826_3311# 1.46e-19
C4759 _110_ a_9681_2601# 4.53e-19
C4760 a_937_3855# VPWR 1.28e-19
C4761 net19 cal_itt\[0\] 0.0181f
C4762 net34 a_13607_1513# 3.03e-21
C4763 _121_ _034_ 0.0165f
C4764 _070_ _002_ 9.91e-19
C4765 mask\[5\] VPWR 1.68f
C4766 net51 net30 8.47e-20
C4767 a_10781_3311# trim_mask\[3\] 1.15e-19
C4768 net36 trimb[0] 0.0182f
C4769 clknet_0_clk a_7723_6807# 0.00228f
C4770 trim_mask\[2\] a_13393_1707# 0.00278f
C4771 clknet_2_3__leaf_clk a_11814_9295# 0.0097f
C4772 net45 a_3933_2767# 0.00532f
C4773 net35 _109_ 3.95e-20
C4774 _058_ a_12502_4765# 2.66e-19
C4775 a_13059_4631# _109_ 0.0986f
C4776 net7 ctln[1] 0.0117f
C4777 net34 trimb[1] 0.0785f
C4778 clknet_0_clk a_7210_5807# 0.0319f
C4779 a_13825_5185# a_14334_5309# 2.6e-19
C4780 a_13257_4943# a_13703_4943# 2.28e-19
C4781 net16 _136_ 0.0255f
C4782 clknet_2_3__leaf_clk a_11622_7485# 0.0162f
C4783 net44 a_5037_6031# 0.0019f
C4784 a_6999_12015# VPWR 0.142f
C4785 a_13415_2442# _031_ 0.11f
C4786 _053_ a_8473_5193# 0.018f
C4787 mask\[5\] a_5699_9269# 5.3e-21
C4788 _134_ a_13783_6183# 0.0393f
C4789 mask\[2\] a_2787_7119# 7.21e-21
C4790 _064_ a_8583_3317# 8.59e-21
C4791 a_5363_12559# a_6927_12559# 4.46e-21
C4792 _051_ a_5524_1679# 2.53e-19
C4793 a_6743_10933# a_7355_11305# 0.00188f
C4794 _021_ a_7164_11293# 0.158f
C4795 a_6210_4989# _100_ 0.0016f
C4796 mask\[6\] a_6099_10633# 6.45e-20
C4797 a_6173_7119# a_7197_7119# 2.36e-20
C4798 _065_ a_6515_8534# 0.00104f
C4799 _099_ _097_ 0.0211f
C4800 a_3817_4697# _014_ 2.65e-20
C4801 _058_ a_11321_3855# 2.63e-19
C4802 a_14236_8457# VPWR 0.176f
C4803 net43 a_4165_11989# 0.166f
C4804 a_1835_12319# mask\[7\] 0.00165f
C4805 _074_ a_816_6031# 0.00471f
C4806 net46 _066_ 2.54e-19
C4807 net47 a_13279_8207# 1.11e-19
C4808 cal_itt\[0\] cal_itt\[1\] 0.944f
C4809 a_1129_7361# result[1] 0.00102f
C4810 a_455_8181# result[2] 0.332f
C4811 _110_ a_11951_2601# 9.34e-19
C4812 _076_ cal_itt\[3\] 1.53e-20
C4813 net12 a_6737_3855# 8.49e-19
C4814 a_4498_4373# state\[1\] 8.56e-19
C4815 clknet_2_0__leaf_clk _051_ 3.44e-19
C4816 net2 _135_ 0.0394f
C4817 clknet_2_3__leaf_clk a_13825_6031# 0.0449f
C4818 _003_ net30 0.0681f
C4819 _125_ _128_ 8.35e-19
C4820 calibrate _054_ 6.74e-19
C4821 net4 a_10903_7261# 1.42e-21
C4822 net43 _019_ 0.0021f
C4823 _033_ a_10111_1679# 1.35e-19
C4824 net18 ctln[4] 0.00336f
C4825 mask\[7\] a_2450_9955# 1.25e-20
C4826 net25 mask\[3\] 0.199f
C4827 a_9839_3615# a_9595_1679# 6.38e-21
C4828 _050_ _090_ 0.0666f
C4829 _107_ a_6197_4399# 2.8e-19
C4830 a_11895_7669# a_12520_7637# 0.185f
C4831 _037_ a_12061_7669# 0.0834f
C4832 a_9369_4105# a_9478_4105# 0.14f
C4833 _078_ a_6007_9839# 0.0791f
C4834 clknet_2_0__leaf_clk _014_ 0.0967f
C4835 trim_mask\[0\] a_11057_4105# 0.0828f
C4836 net43 a_1493_11721# 0.0107f
C4837 a_5037_6031# en_co_clk 2.38e-19
C4838 cal_count\[0\] a_11575_8790# 0.00526f
C4839 mask\[1\] net2 3.22e-20
C4840 net14 mask\[3\] 2.84e-21
C4841 net3 a_3365_4943# 2.32e-20
C4842 a_1579_11471# result[5] 5.81e-21
C4843 a_1129_6273# calibrate 3.2e-20
C4844 a_3208_10205# mask\[2\] 6.41e-20
C4845 mask\[2\] a_2689_8751# 0.0502f
C4846 _065_ a_4498_4373# 0.00109f
C4847 a_6191_12559# _084_ 0.00229f
C4848 net20 a_5496_12131# 2.23e-19
C4849 _045_ a_6375_12021# 6.75e-19
C4850 _121_ a_3830_6281# 4.96e-19
C4851 a_7800_4631# clk 0.00819f
C4852 en_co_clk a_7800_4631# 2.05e-21
C4853 cal_count\[0\] _126_ 0.239f
C4854 a_1476_4777# a_1585_4777# 0.00742f
C4855 a_1651_4703# a_1830_4765# 0.0074f
C4856 _042_ a_3521_9813# 0.00526f
C4857 _053_ a_8583_3317# 0.00136f
C4858 _090_ _052_ 1.32e-19
C4859 a_2601_3285# VPWR 0.213f
C4860 net15 net44 2.1e-21
C4861 _049_ a_6197_4399# 5.97e-22
C4862 _035_ a_10593_9295# 0.144f
C4863 a_10239_9295# a_10774_9661# 0.0018f
C4864 a_12612_8725# a_12916_8751# 3.11e-19
C4865 a_12436_9129# a_12522_8751# 0.00972f
C4866 _010_ a_3511_11471# 1.01e-19
C4867 _023_ _102_ 2.21e-19
C4868 _020_ _008_ 3.4e-20
C4869 a_13142_7271# _134_ 2.16e-19
C4870 a_4498_4373# a_5054_4399# 0.0139f
C4871 clknet_2_2__leaf_clk trim_mask\[1\] 0.374f
C4872 net13 _051_ 0.0111f
C4873 net34 a_14334_1135# 5.17e-20
C4874 _090_ _098_ 1.75e-19
C4875 a_13257_4943# a_13459_3317# 7.12e-22
C4876 _074_ a_1835_11231# 5.88e-20
C4877 _072_ a_6515_6794# 2.13e-20
C4878 a_10975_6031# _108_ 5.19e-20
C4879 clknet_2_2__leaf_clk a_6703_2197# 5.33e-20
C4880 net27 mask\[5\] 0.816f
C4881 _039_ VPWR 0.68f
C4882 _078_ a_1541_9117# 0.00136f
C4883 net19 trim_mask\[0\] 0.287f
C4884 cal_itt\[0\] _001_ 0.0135f
C4885 ctlp[2] trimb[3] 0.00996f
C4886 _122_ a_12824_7663# 3.06e-19
C4887 a_8307_4719# VPWR 0.00295f
C4888 _129_ VPWR 0.627f
C4889 net4 a_9662_3855# 3.06e-19
C4890 net44 a_7351_8041# 0.00943f
C4891 clknet_2_3__leaf_clk _092_ 0.0956f
C4892 a_9405_9295# VPWR 1.15e-19
C4893 a_1677_9545# a_1279_9129# 2.12e-19
C4894 net31 _135_ 6.2e-21
C4895 net2 a_14063_7093# 0.0259f
C4896 a_11016_6691# cal_count\[3\] 2.16e-19
C4897 clknet_2_1__leaf_clk result[6] 0.0373f
C4898 cal_count\[0\] a_12153_8757# 0.498f
C4899 _048_ a_3530_4765# 1.16e-19
C4900 net33 clkc 2.25e-19
C4901 a_6999_12015# net27 2.35e-19
C4902 net43 VPWR 4.71f
C4903 _056_ a_15023_1135# 7.29e-19
C4904 net37 _055_ 0.0027f
C4905 _067_ a_10781_5807# 1.47e-19
C4906 net24 mask\[1\] 0.00304f
C4907 a_13919_8751# a_15023_8751# 2.19e-20
C4908 net43 a_1769_12393# 6.03e-19
C4909 a_745_12021# a_1203_12015# 0.0346f
C4910 net45 a_1651_4703# 0.344f
C4911 net19 a_7723_10143# 0.00189f
C4912 net53 a_6888_10205# 0.00818f
C4913 net15 clk 0.0472f
C4914 net15 en_co_clk 0.00947f
C4915 a_6763_5193# _103_ 7.91e-19
C4916 a_13257_4943# _109_ 0.00209f
C4917 net14 a_1579_5807# 1.81e-19
C4918 clknet_2_2__leaf_clk a_8749_3317# 0.00584f
C4919 a_14335_4020# a_13625_3317# 3.4e-20
C4920 net16 a_11987_8757# 6.15e-20
C4921 net12 net53 0.0178f
C4922 a_6927_12559# ctlp[6] 0.372f
C4923 a_14604_3017# a_14604_2339# 0.0129f
C4924 a_7010_3631# VPWR 4.8e-20
C4925 a_8105_10383# a_8360_10383# 0.0594f
C4926 a_7939_10383# a_8563_10749# 9.73e-19
C4927 _120_ a_3461_5193# 8.29e-19
C4928 a_3667_3829# _015_ 0.0142f
C4929 _074_ a_937_4105# 0.0159f
C4930 cal_itt\[1\] trim_mask\[0\] 7.2e-20
C4931 a_395_9845# result[4] 0.0131f
C4932 a_14236_8457# a_14807_8359# 0.00852f
C4933 _040_ a_6419_8207# 2.37e-20
C4934 a_7351_8041# en_co_clk 4.11e-21
C4935 clknet_2_2__leaf_clk a_10977_2543# 3.13e-21
C4936 _078_ a_5363_7369# 4.42e-20
C4937 net4 a_9572_2601# 9.85e-20
C4938 net16 net34 0.0142f
C4939 _074_ a_5578_12131# 5.4e-19
C4940 a_5515_6005# a_5455_4943# 0.00132f
C4941 trim_val\[2\] a_13512_1501# 7.84e-20
C4942 net55 net42 0.163f
C4943 a_1844_9129# _081_ 0.00126f
C4944 net24 a_1387_8751# 0.0265f
C4945 a_10586_7371# a_10903_7261# 0.102f
C4946 _119_ a_8912_2589# 4.88e-19
C4947 a_6173_7119# a_7250_7485# 1.46e-19
C4948 net53 a_6983_10217# 0.00637f
C4949 clknet_2_1__leaf_clk a_6835_7669# 0.26f
C4950 net31 _127_ 3.67e-20
C4951 a_10239_9295# _065_ 1.44e-20
C4952 net8 a_13703_1513# 7.53e-19
C4953 _104_ a_9369_4105# 6.76e-19
C4954 a_448_7637# _080_ 0.00498f
C4955 a_11509_3317# a_11859_3689# 0.207f
C4956 net44 a_7548_10217# 0.235f
C4957 _006_ _081_ 0.117f
C4958 _078_ _101_ 1.01f
C4959 net19 a_8717_10383# 5.15e-19
C4960 a_448_6549# result[0] 0.158f
C4961 cal_count\[0\] a_11268_9295# 4.68e-20
C4962 _053_ a_7190_3855# 0.186f
C4963 net30 a_9099_3689# 3.34e-21
C4964 cal_itt\[0\] a_7916_8041# 7.11e-20
C4965 a_579_10933# a_448_10357# 3.9e-19
C4966 mask\[5\] a_8455_10383# 4.63e-19
C4967 _009_ ctlp[6] 2.05e-20
C4968 net35 a_14655_4399# 0.11f
C4969 net31 a_13519_4007# 2.36e-20
C4970 a_13557_7369# a_13279_7119# 3.25e-19
C4971 clknet_2_2__leaf_clk _115_ 8.04e-20
C4972 _084_ a_6796_12381# 4.93e-20
C4973 clknet_2_1__leaf_clk a_5915_11721# 0.00345f
C4974 _101_ a_2869_11247# 0.00145f
C4975 net30 a_10055_5487# 7.16e-19
C4976 trim_mask\[0\] a_11067_4405# 8.88e-19
C4977 clknet_2_0__leaf_clk a_5535_8181# 3.24e-21
C4978 net42 a_7715_3285# 2.09e-21
C4979 a_3615_8207# a_4349_8449# 0.0701f
C4980 a_5363_12559# mask\[6\] 0.00634f
C4981 _119_ a_10543_2455# 4.94e-19
C4982 _045_ a_4512_12393# 7.2e-20
C4983 _032_ a_9805_1473# 0.00138f
C4984 trim_val\[3\] _117_ 0.00648f
C4985 a_9761_1679# _116_ 3.56e-20
C4986 a_6822_4399# VPWR 0.00464f
C4987 net43 net27 0.021f
C4988 net2 a_13279_7119# 0.00118f
C4989 net18 en_co_clk 0.00801f
C4990 net19 a_8949_6281# 0.00228f
C4991 _067_ a_8935_6895# 6.58e-21
C4992 net4 a_9889_6873# 7.28e-19
C4993 a_2857_7637# VPWR 1.22f
C4994 net47 _069_ 3.22e-19
C4995 _128_ a_13142_8359# 0.233f
C4996 _113_ a_12424_3689# 0.00303f
C4997 clknet_2_3__leaf_clk a_11045_5807# 0.00164f
C4998 _126_ a_13919_8751# 6.56e-22
C4999 _086_ _078_ 0.00406f
C5000 a_11491_6031# a_11599_6397# 0.0572f
C5001 net31 a_14604_3017# 0.0148f
C5002 a_2953_9845# _019_ 1.38e-19
C5003 a_2877_2197# a_2767_2223# 0.0977f
C5004 net47 a_8022_7119# 3.95e-19
C5005 a_12533_3689# VPWR 1.2e-20
C5006 clknet_2_1__leaf_clk a_7201_9813# 7.33e-21
C5007 a_7569_7637# a_7916_8041# 0.0512f
C5008 a_7001_7669# _071_ 1.05e-19
C5009 a_1019_4399# valid 7.82e-19
C5010 _093_ a_937_4105# 0.00717f
C5011 _101_ a_3597_10933# 5.62e-19
C5012 a_2601_3285# a_2383_3689# 0.21f
C5013 a_2033_3317# a_3123_3615# 0.0424f
C5014 a_1867_3317# a_2948_3689# 0.102f
C5015 _011_ a_1000_11293# 2.6e-20
C5016 _136_ clkc 5.39e-20
C5017 a_14318_8457# VPWR 0.00246f
C5018 a_12323_4703# VPWR 0.411f
C5019 _078_ _102_ 0.00123f
C5020 net30 _088_ 2.51e-19
C5021 cal_count\[0\] a_13050_7637# 1.02e-20
C5022 net46 a_12056_6031# 0.227f
C5023 a_11709_6273# cal_count\[3\] 0.0186f
C5024 trim_mask\[4\] net10 5.9e-22
C5025 net37 a_15259_7637# 4.62e-20
C5026 trim_mask\[1\] a_14540_3689# 4.23e-19
C5027 cal_itt\[1\] a_8949_6281# 0.0437f
C5028 net14 clk 0.0521f
C5029 _094_ _120_ 0.0625f
C5030 net38 _125_ 1.01e-19
C5031 _116_ a_10787_1135# 5.83e-20
C5032 net30 a_7262_5461# 0.00307f
C5033 a_13625_3317# a_15299_3311# 1.92e-19
C5034 a_8022_7119# a_8820_6005# 1.35e-20
C5035 _096_ a_4815_3031# 6.38e-21
C5036 a_12153_8757# a_13919_8751# 3.33e-21
C5037 net44 a_5449_6031# 6.03e-19
C5038 clknet_2_1__leaf_clk a_911_10217# 0.0364f
C5039 net41 a_5177_1921# 2.4e-20
C5040 _053_ a_9957_7663# 3.07e-19
C5041 net33 a_15023_9839# 0.0101f
C5042 a_3748_6281# a_4259_6031# 6.09e-19
C5043 a_448_10357# a_395_9845# 0.0131f
C5044 a_8270_8029# VPWR 3.12e-19
C5045 net46 a_14071_3689# 0.00328f
C5046 mask\[6\] a_579_10933# 5.74e-21
C5047 _065_ _066_ 0.107f
C5048 net38 trimb[0] 0.00705f
C5049 net30 trim_val\[4\] 6.05e-20
C5050 net52 net45 0.356f
C5051 state\[2\] a_7223_2465# 1.55e-21
C5052 _063_ a_9443_6059# 0.185f
C5053 _110_ a_9369_4105# 0.004f
C5054 net19 a_8307_4943# 0.00233f
C5055 _065_ a_10621_7119# 4.06e-19
C5056 net34 trimb[3] 0.00164f
C5057 en_co_clk trim_val\[0\] 7.78e-20
C5058 a_8307_4719# _104_ 0.096f
C5059 net12 a_6007_9839# 0.00206f
C5060 a_1173_6031# VPWR 2.38e-19
C5061 net46 _058_ 0.0779f
C5062 _008_ _077_ 1.23e-20
C5063 _101_ a_5502_6397# 8.97e-21
C5064 _081_ _017_ 8.78e-21
C5065 net50 a_10872_1455# 3.6e-19
C5066 clknet_2_3__leaf_clk a_9003_3829# 4.93e-20
C5067 a_7571_4943# a_7527_4631# 7.99e-20
C5068 _078_ _022_ 2.81e-20
C5069 _065_ a_4175_4943# 1.74e-20
C5070 a_2953_9845# VPWR 0.585f
C5071 net29 ctlp[0] 4.27e-19
C5072 a_10239_9295# _067_ 1.25e-19
C5073 a_7109_11989# a_7618_12015# 2.6e-19
C5074 net16 cal_count\[3\] 2.33e-19
C5075 a_4091_5309# _093_ 8.93e-19
C5076 _122_ a_12061_7669# 0.00197f
C5077 net35 trim[1] 0.0359f
C5078 net51 a_5691_7637# 0.293f
C5079 net19 a_8298_2767# 0.0269f
C5080 en_co_clk a_5449_6031# 3.92e-19
C5081 a_6173_7119# _049_ 4.22e-19
C5082 net24 _041_ 0.0067f
C5083 _014_ a_2948_3689# 0.00182f
C5084 a_7019_4407# a_7010_3311# 2.25e-20
C5085 a_2787_7119# _120_ 1.8e-20
C5086 _095_ net3 0.193f
C5087 net23 a_3053_8207# 3.31e-21
C5088 _063_ a_12061_7669# 3.52e-20
C5089 net19 _042_ 0.0106f
C5090 _104_ a_7010_3631# 0.00332f
C5091 a_7201_9813# a_7245_10205# 3.69e-19
C5092 a_6633_9845# a_7657_10217# 2.36e-20
C5093 a_8657_2229# a_9103_2601# 2.28e-19
C5094 clknet_2_1__leaf_clk mask\[2\] 0.387f
C5095 net15 a_3565_7119# 3.43e-19
C5096 net55 a_4886_4399# 4.17e-20
C5097 a_5524_9295# _077_ 5.29e-19
C5098 a_14379_6397# VPWR 0.217f
C5099 state\[1\] a_4576_3427# 2.14e-19
C5100 _074_ a_3840_8867# 2.68e-20
C5101 _033_ a_9839_3615# 2.48e-20
C5102 a_8583_3317# a_9664_3689# 0.102f
C5103 _131_ _134_ 0.0982f
C5104 a_4308_4917# _099_ 3.79e-20
C5105 a_1638_7485# VPWR 8.34e-19
C5106 net37 trim_mask\[0\] 0.00301f
C5107 calibrate a_3339_2767# 1.6e-20
C5108 a_5691_7637# _003_ 2.29e-19
C5109 a_13100_8751# VPWR 0.00296f
C5110 _038_ VPWR 0.377f
C5111 _118_ a_10975_4105# 2.6e-19
C5112 calibrate a_995_3530# 0.00115f
C5113 trim_mask\[1\] a_14335_2442# 2.07e-19
C5114 _034_ a_4091_5309# 6.52e-19
C5115 a_8673_10625# a_8215_9295# 9.42e-21
C5116 a_8105_10383# _000_ 2.54e-19
C5117 _096_ a_5087_3855# 0.00608f
C5118 a_10405_9295# a_11394_9509# 0.0728f
C5119 a_9296_9295# a_10593_9295# 5.79e-20
C5120 a_8381_9295# a_9405_9295# 2.36e-20
C5121 a_10864_9269# a_10688_9295# 0.26f
C5122 net2 _002_ 0.0574f
C5123 trim_val\[1\] a_13881_2741# 0.184f
C5124 _022_ a_3597_10933# 0.329f
C5125 a_3431_10933# a_4165_10901# 0.0701f
C5126 net4 a_11141_6031# 1.23e-21
C5127 a_2659_2601# clk 0.00437f
C5128 net14 ctln[0] 0.00137f
C5129 _051_ _028_ 0.156f
C5130 cal_itt\[1\] a_7723_6807# 5.31e-20
C5131 a_7548_10217# a_8992_9955# 4.14e-20
C5132 a_4512_11305# _042_ 1.08e-19
C5133 a_9007_2601# a_9572_2601# 7.99e-20
C5134 net18 a_10688_9295# 0.00994f
C5135 mask\[3\] _019_ 0.0342f
C5136 a_10975_6031# a_11587_6031# 0.00188f
C5137 a_2787_9845# a_3411_9839# 9.73e-19
C5138 a_1651_6005# a_1493_5487# 3.48e-20
C5139 result[7] result[5] 7.15e-19
C5140 net1 cal 0.0211f
C5141 en_co_clk a_11023_5108# 1.38e-21
C5142 _058_ a_11343_3317# 0.00513f
C5143 _065_ a_6515_6794# 1.15e-19
C5144 clknet_2_1__leaf_clk a_6428_7119# 2.39e-19
C5145 _058_ a_11149_3017# 2.93e-19
C5146 net52 a_2953_7119# 8.1e-20
C5147 _096_ a_1476_4777# 4.88e-19
C5148 net44 a_7460_5807# 2.22e-22
C5149 state\[2\] _088_ 0.00635f
C5150 _061_ trim[1] 6.73e-21
C5151 clknet_2_1__leaf_clk a_1000_11293# 0.00313f
C5152 cal_count\[0\] VPWR 1.12f
C5153 a_5915_10927# a_6181_10633# 1.58e-19
C5154 _021_ a_6099_10633# 7.91e-20
C5155 net34 clkc 0.00407f
C5156 _064_ a_11149_2767# 0.00344f
C5157 clknet_2_0__leaf_clk net22 0.0104f
C5158 a_1585_10217# VPWR 5.52e-20
C5159 mask\[0\] a_3521_7361# 0.0221f
C5160 _085_ clknet_2_1__leaf_clk 0.196f
C5161 net29 a_579_12021# 0.00205f
C5162 a_4617_4105# VPWR 0.178f
C5163 net9 a_13092_8029# 1.72e-20
C5164 a_7263_7093# _048_ 3.18e-20
C5165 _101_ a_6888_10205# 2.57e-21
C5166 a_10405_9295# a_11116_8983# 0.00114f
C5167 net9 trim_mask\[0\] 0.0947f
C5168 _054_ a_7184_2339# 1.63e-22
C5169 a_1129_7361# a_1476_7119# 0.0512f
C5170 clknet_0_clk a_8307_4719# 9.47e-19
C5171 _067_ _066_ 0.155f
C5172 net46 a_13607_4943# 0.183f
C5173 clknet_2_3__leaf_clk _035_ 0.107f
C5174 _050_ a_3667_3829# 5.94e-19
C5175 net12 _101_ 0.0151f
C5176 mask\[7\] a_1313_10901# 0.00354f
C5177 _067_ a_10621_7119# 4.31e-19
C5178 net53 a_5997_10927# 0.0106f
C5179 _029_ a_13703_4943# 2.29e-19
C5180 a_8307_6575# clk 1.17e-19
C5181 net33 a_14715_3615# 0.00975f
C5182 net44 a_7933_11305# 8.4e-19
C5183 cal_itt\[2\] net30 0.00218f
C5184 _053_ _103_ 9.49e-19
C5185 a_8307_6575# en_co_clk 1.15e-19
C5186 net43 clknet_0_clk 0.152f
C5187 net14 a_1184_9117# 0.00314f
C5188 net9 a_10405_9295# 5.19e-20
C5189 a_6519_4631# state\[2\] 0.00202f
C5190 _050_ _033_ 9.69e-19
C5191 net19 a_6909_10933# 5.02e-19
C5192 state\[2\] a_5686_2045# 8.41e-20
C5193 a_1191_12393# ctlp[0] 3.92e-20
C5194 a_4349_8449# a_4227_8207# 3.16e-19
C5195 _072_ _069_ 4.94e-20
C5196 a_7460_5807# clk 0.00292f
C5197 a_5449_6031# _059_ 1.23e-19
C5198 net52 a_3922_8867# 1.32e-19
C5199 mask\[3\] VPWR 1.86f
C5200 _072_ a_8022_7119# 0.0135f
C5201 net28 ctlp[0] 0.0759f
C5202 mask\[4\] a_8105_10383# 0.00152f
C5203 a_4259_6031# a_4308_4917# 3.85e-20
C5204 _101_ a_5340_6031# 1.38e-19
C5205 _128_ a_13557_8457# 6.9e-20
C5206 _068_ _069_ 1.84e-20
C5207 _053_ a_10903_7261# 0.0108f
C5208 a_6741_7361# VPWR 0.219f
C5209 clknet_2_3__leaf_clk _136_ 0.181f
C5210 _045_ a_7456_12393# 9.55e-21
C5211 _101_ a_6983_10217# 3.18e-21
C5212 _074_ a_395_6031# 0.0166f
C5213 _066_ clknet_2_2__leaf_clk 6.69e-19
C5214 a_9471_9269# _065_ 2.22e-20
C5215 _068_ a_8022_7119# 0.0139f
C5216 cal_itt\[0\] _062_ 0.266f
C5217 _122_ a_11396_6031# 3.67e-19
C5218 net16 a_14347_4917# 0.00684f
C5219 _093_ a_4886_4399# 5.61e-19
C5220 _074_ a_6793_8970# 7.09e-21
C5221 mask\[3\] a_5699_9269# 0.101f
C5222 _090_ _087_ 0.0952f
C5223 _048_ a_6737_3855# 0.00637f
C5224 cal_itt\[0\] a_10138_5807# 2.4e-19
C5225 a_5515_6005# _092_ 7.91e-20
C5226 net45 a_3057_3689# 4.56e-19
C5227 a_13415_2442# trim_val\[2\] 1.82e-19
C5228 _115_ a_14335_2442# 9.01e-19
C5229 _090_ a_6519_3829# 1.96e-20
C5230 mask\[0\] _095_ 0.00186f
C5231 VPWR ctln[4] 0.193f
C5232 _115_ net8 2.98e-19
C5233 _106_ a_9125_4943# 7.22e-21
C5234 net43 a_7459_7663# 0.0135f
C5235 a_561_4405# net1 0.00824f
C5236 _012_ a_855_4105# 0.152f
C5237 a_14467_8751# a_14236_8457# 0.00117f
C5238 net44 a_7477_10901# 0.177f
C5239 _039_ a_2476_6281# 4.96e-19
C5240 en_co_clk a_5363_4719# 8.37e-19
C5241 net15 a_2787_10927# 0.0133f
C5242 _090_ _099_ 0.07f
C5243 net12 a_6785_7119# 4.47e-19
C5244 _125_ net40 0.227f
C5245 net37 a_14983_9269# 0.0104f
C5246 net3 calibrate 0.00995f
C5247 net24 a_3615_8207# 1.18e-19
C5248 _064_ a_9572_2601# 8.48e-20
C5249 net12 a_6703_2197# 0.00486f
C5250 _100_ _088_ 3.2e-19
C5251 _107_ a_7800_4631# 0.00575f
C5252 net45 state\[1\] 0.105f
C5253 trim_mask\[0\] a_10188_4105# 0.0193f
C5254 _029_ a_13459_3317# 2.08e-20
C5255 _123_ a_13008_7663# 0.00163f
C5256 net43 a_3521_9813# 0.182f
C5257 _076_ _073_ 7.03e-20
C5258 a_10270_4105# VPWR 0.00144f
C5259 a_3578_2589# VPWR 7.03e-20
C5260 a_11116_8983# a_11258_8790# 0.00557f
C5261 a_1579_5807# VPWR 1.43e-19
C5262 _049_ a_5037_6031# 3.28e-19
C5263 a_3947_12393# a_3947_11305# 0.00153f
C5264 a_4959_1679# clk 0.0298f
C5265 _119_ a_10699_3311# 1.41e-19
C5266 a_4687_12319# a_6541_12021# 9.64e-21
C5267 a_10543_2455# a_10111_1679# 0.00351f
C5268 net46 a_11488_4765# 8.97e-19
C5269 _065_ net45 6.92e-19
C5270 _129_ a_14564_6397# 7.67e-22
C5271 _094_ _051_ 9.78e-22
C5272 _050_ _054_ 0.0156f
C5273 net25 result[3] 0.00624f
C5274 _049_ a_7800_4631# 0.00546f
C5275 net12 _060_ 2.45e-20
C5276 a_579_12021# a_1191_12393# 0.00188f
C5277 _011_ a_1000_12381# 0.16f
C5278 a_4687_11231# _019_ 9.46e-20
C5279 a_2857_7637# clknet_0_clk 0.345f
C5280 a_6519_4631# _100_ 0.109f
C5281 _029_ _109_ 7.06e-19
C5282 net44 _019_ 5.55e-19
C5283 _046_ _078_ 0.357f
C5284 _065_ _058_ 8.88e-19
C5285 a_911_10217# result[4] 0.00118f
C5286 a_7897_6913# clk 9.6e-19
C5287 _118_ a_9099_3689# 0.0115f
C5288 net23 net45 0.0169f
C5289 a_15299_6575# clkc 0.11f
C5290 net13 a_4165_10901# 0.00324f
C5291 net30 net55 0.0559f
C5292 a_5363_12559# ctlp[7] 0.373f
C5293 net14 result[3] 8.01e-20
C5294 a_455_12533# _011_ 0.00175f
C5295 net18 _108_ 0.192f
C5296 net28 a_579_12021# 0.0118f
C5297 a_6375_12021# net12 1.3e-19
C5298 net27 mask\[3\] 1.52e-20
C5299 net46 _113_ 0.14f
C5300 trim_mask\[0\] trim_mask\[3\] 3.32e-21
C5301 a_13919_8751# VPWR 0.242f
C5302 _129_ a_14467_8751# 0.00178f
C5303 a_3513_12809# VPWR 0.00643f
C5304 a_4043_11305# VPWR 5.51e-19
C5305 a_448_11445# _007_ 8.94e-20
C5306 net34 a_15023_9839# 0.0167f
C5307 net43 a_1007_7119# 0.00168f
C5308 _052_ _054_ 3.87e-19
C5309 a_12323_4703# _110_ 4.67e-19
C5310 a_13257_4943# _112_ 0.00101f
C5311 a_561_7119# net22 8.85e-20
C5312 a_5340_6031# _060_ 3.21e-21
C5313 net4 a_8491_2229# 2.28e-19
C5314 net42 a_6763_5193# 0.00125f
C5315 a_9889_6873# _064_ 1.39e-19
C5316 _062_ trim_mask\[0\] 0.245f
C5317 _074_ net30 0.0754f
C5318 net41 a_2601_3285# 0.0219f
C5319 _102_ a_1651_10143# 4.63e-19
C5320 a_10055_5487# _118_ 3.83e-19
C5321 clknet_2_3__leaf_clk a_11987_8757# 0.22f
C5322 net18 a_10655_2932# 6.73e-20
C5323 _015_ a_3339_2767# 6.02e-20
C5324 net48 a_13307_1707# 4.38e-19
C5325 a_8949_6281# a_8949_6031# 6.96e-20
C5326 trim_mask\[0\] a_10138_5807# 0.00917f
C5327 a_6007_7119# a_6428_7119# 0.0931f
C5328 a_13091_1141# a_13825_1109# 0.0701f
C5329 _062_ _075_ 0.442f
C5330 net15 _049_ 0.0163f
C5331 a_1099_12533# a_1203_10927# 1.35e-20
C5332 net9 _030_ 3.65e-20
C5333 net44 a_6467_9845# 0.304f
C5334 _095_ net54 0.173f
C5335 _126_ cal_count\[1\] 0.095f
C5336 net15 a_3388_4631# 0.00477f
C5337 clknet_2_1__leaf_clk a_2828_12131# 0.00905f
C5338 net47 a_14347_9480# 8.66e-20
C5339 a_4259_6031# _090_ 5.41e-22
C5340 a_561_6031# a_1129_6273# 0.18f
C5341 net13 a_4871_6031# 0.00101f
C5342 a_9471_9269# _067_ 2.4e-21
C5343 a_10864_9269# a_11436_9295# 1.57e-19
C5344 a_14347_9480# a_14377_9545# 0.025f
C5345 a_13881_2741# a_14184_2767# 0.00138f
C5346 mask\[7\] result[5] 0.00214f
C5347 net46 a_8657_2229# 0.024f
C5348 a_12323_4703# a_12148_4777# 0.234f
C5349 a_10975_4105# a_11321_3855# 0.0134f
C5350 a_11233_4405# _058_ 0.042f
C5351 a_9459_7895# VPWR 0.222f
C5352 net18 a_11436_9295# 1.57e-19
C5353 net47 a_13142_7271# 8.16e-19
C5354 a_4687_11231# VPWR 0.382f
C5355 net43 a_1830_10205# 0.00413f
C5356 net43 a_2775_9071# 1.37e-20
C5357 _059_ a_5363_4719# 0.0535f
C5358 _101_ a_6631_7485# 7.37e-21
C5359 net45 a_2225_7663# 0.0535f
C5360 net44 VPWR 3.87f
C5361 _046_ a_3597_10933# 6.44e-20
C5362 _108_ trim_val\[0\] 0.37f
C5363 a_11488_4765# a_11343_3317# 9.89e-21
C5364 net45 _016_ 0.0528f
C5365 net33 _047_ 0.0023f
C5366 a_4864_1679# ctln[7] 5.95e-20
C5367 a_14249_8725# _133_ 1.84e-20
C5368 net53 a_5177_9537# 4.45e-21
C5369 net19 a_9369_4105# 0.00139f
C5370 _017_ a_3781_8207# 0.316f
C5371 _119_ _027_ 6.44e-20
C5372 net45 a_1019_6397# 0.0122f
C5373 a_13307_1707# a_13091_1141# 0.00722f
C5374 net44 a_5699_9269# 0.337f
C5375 a_12153_8757# cal_count\[1\] 6.28e-20
C5376 _041_ a_12756_9117# 0.00181f
C5377 a_13142_8725# a_13256_9117# 1.84e-19
C5378 a_12992_8751# a_13184_9117# 0.00536f
C5379 a_395_4405# a_911_4777# 0.115f
C5380 net26 a_6633_9845# 0.555f
C5381 a_561_9845# _006_ 1.06e-20
C5382 a_395_9845# a_1497_8725# 1.76e-19
C5383 a_1313_11989# ctlp[0] 9.95e-19
C5384 a_8389_5193# _106_ 3.99e-19
C5385 _065_ a_2953_7119# 5.84e-19
C5386 a_3615_8207# a_4677_7882# 3.45e-19
C5387 net19 mask\[5\] 0.033f
C5388 _042_ net9 3.59e-19
C5389 net5 a_13783_6183# 7.27e-20
C5390 clknet_2_1__leaf_clk _120_ 8.85e-21
C5391 _118_ trim_val\[4\] 0.385f
C5392 a_10975_4105# a_11435_2229# 1.23e-19
C5393 a_5515_6005# a_5547_5603# 0.00185f
C5394 a_4696_8207# net45 1.03e-19
C5395 net18 _107_ 2.1e-20
C5396 a_12900_7663# a_13164_8029# 0.00384f
C5397 a_13050_7637# cal_count\[2\] 0.00355f
C5398 calibrate valid 0.00353f
C5399 net14 en 0.0186f
C5400 VPWR clk 4.31f
C5401 en_co_clk VPWR 6.66f
C5402 net23 a_2953_7119# 8.7e-20
C5403 state\[1\] a_4905_3855# 1.67e-19
C5404 net43 a_6523_7119# 1.25e-19
C5405 ctlp[7] ctlp[6] 0.0358f
C5406 net15 a_3425_11721# 2.39e-19
C5407 net6 a_3063_591# 3.17e-21
C5408 _121_ a_3891_4943# 9.37e-20
C5409 a_8386_8457# VPWR 0.00587f
C5410 a_9084_4515# VPWR 0.174f
C5411 a_14249_8725# a_14236_8457# 5.27e-19
C5412 _092_ a_4815_3031# 1.18e-21
C5413 net30 _093_ 9.79e-21
C5414 a_10975_6031# a_11491_6031# 0.111f
C5415 a_9761_1679# a_10016_1679# 0.0642f
C5416 a_5515_6005# a_5536_4399# 7.38e-22
C5417 clknet_2_1__leaf_clk a_1000_12381# 0.00142f
C5418 trim_mask\[1\] a_13459_3317# 0.0168f
C5419 a_6428_7119# cal_itt\[3\] 1.38e-19
C5420 a_13825_1109# a_14281_1513# 4.2e-19
C5421 a_13607_1513# a_13869_1501# 0.00171f
C5422 a_13091_1141# a_13715_1135# 9.73e-19
C5423 net55 state\[2\] 0.0135f
C5424 a_6210_4989# a_5931_4105# 8.56e-21
C5425 calibrate a_5537_4105# 0.00292f
C5426 _065_ a_3922_8867# 8.49e-22
C5427 a_12153_8757# a_12612_8725# 0.078f
C5428 mask\[5\] a_4512_11305# 1.74e-20
C5429 a_7999_11231# a_7723_10143# 3.86e-20
C5430 net9 a_11951_2601# 0.00535f
C5431 _062_ a_8949_6281# 0.0075f
C5432 a_14172_1513# trim[3] 4.32e-19
C5433 a_455_12533# clknet_2_1__leaf_clk 0.0131f
C5434 a_2877_2197# a_3224_2601# 0.0512f
C5435 clknet_2_1__leaf_clk a_4609_9295# 0.00174f
C5436 a_11067_3017# a_11601_2229# 3.43e-19
C5437 mask\[6\] a_5915_11721# 0.00553f
C5438 mask\[4\] a_9074_9955# 5.78e-19
C5439 a_2953_9845# a_3521_9813# 0.176f
C5440 net55 state\[0\] 0.00109f
C5441 _095_ a_4471_4007# 8.62e-21
C5442 _067_ a_9693_8029# 0.00165f
C5443 _019_ a_4801_9839# 0.00891f
C5444 net46 a_10569_1109# 1.21e-19
C5445 _063_ _051_ 7.4e-20
C5446 clknet_2_0__leaf_clk _075_ 0.00194f
C5447 clknet_2_3__leaf_clk a_9296_9295# 0.0604f
C5448 net27 a_4687_11231# 6.09e-20
C5449 net45 clknet_2_2__leaf_clk 0.00335f
C5450 _038_ a_10699_5487# 0.111f
C5451 net3 _015_ 0.0538f
C5452 a_11023_5108# _108_ 0.221f
C5453 _109_ trim_mask\[1\] 1.61e-20
C5454 net44 net27 0.105f
C5455 net34 a_14715_3615# 0.00138f
C5456 _101_ a_5997_10927# 0.0119f
C5457 net4 _032_ 3.38e-21
C5458 _123_ a_12520_7637# 0.0316f
C5459 clknet_2_2__leaf_clk _058_ 0.0751f
C5460 _065_ a_2857_5461# 0.0331f
C5461 trim_val\[3\] _116_ 0.00305f
C5462 _065_ _069_ 0.131f
C5463 _016_ a_2953_7119# 0.289f
C5464 net21 net53 1.58e-20
C5465 a_9443_6059# _092_ 0.0421f
C5466 _034_ net30 0.0547f
C5467 net9 a_12344_8041# 0.0153f
C5468 a_579_12021# a_1313_11989# 0.0701f
C5469 _001_ _133_ 5.05e-20
C5470 _011_ a_745_12021# 0.26f
C5471 _018_ a_2961_9545# 0.00249f
C5472 net45 _013_ 0.0723f
C5473 a_7800_4631# trim_mask\[4\] 3.9e-21
C5474 _108_ a_10055_2767# 1.48e-20
C5475 _065_ a_8022_7119# 1.79e-20
C5476 a_1125_7663# a_1129_7361# 0.00133f
C5477 a_10137_4943# trim_val\[4\] 3.3e-19
C5478 net37 a_15083_4659# 0.00802f
C5479 a_8091_7967# VPWR 0.349f
C5480 net13 _075_ 2.54e-20
C5481 a_14249_8725# _129_ 0.115f
C5482 net46 a_10329_1921# 0.189f
C5483 _051_ _096_ 4.33e-21
C5484 net47 a_13562_8751# 0.00217f
C5485 _127_ trimb[1] 6.52e-19
C5486 clknet_2_3__leaf_clk cal_count\[3\] 0.519f
C5487 net19 a_9405_9295# 1.84e-19
C5488 net52 a_2787_9845# 0.0211f
C5489 _062_ a_8307_4943# 3.41e-21
C5490 net54 calibrate 0.0341f
C5491 a_3431_12021# a_4621_12393# 2.56e-19
C5492 a_7891_3617# _033_ 2.41e-20
C5493 VPWR ctln[0] 0.194f
C5494 _096_ _014_ 7.19e-19
C5495 net19 net43 4.36e-20
C5496 clknet_2_0__leaf_clk a_4030_7485# 4.01e-19
C5497 a_3781_8207# a_3868_7119# 9.6e-21
C5498 net43 a_1822_10927# 2.06e-19
C5499 a_14379_6397# a_14564_6397# 0.183f
C5500 a_6541_12021# a_7631_12319# 0.0424f
C5501 a_7109_11989# a_6891_12393# 0.21f
C5502 a_10055_2767# a_10655_2932# 0.0197f
C5503 a_8298_2767# trim_mask\[3\] 1.5e-20
C5504 a_4801_9839# VPWR 0.199f
C5505 _092_ a_5087_3855# 2.66e-19
C5506 _059_ VPWR 0.816f
C5507 _053_ a_11141_6031# 0.0171f
C5508 _049_ a_5449_6031# 1.93e-19
C5509 a_2019_9055# net24 0.133f
C5510 trim_mask\[3\] a_9681_2601# 1.1e-19
C5511 a_11509_3317# a_11764_3677# 0.0564f
C5512 a_3273_4943# a_3891_4943# 0.00113f
C5513 a_8215_9295# a_10593_9295# 7.45e-21
C5514 _069_ a_9761_8457# 0.0012f
C5515 _110_ ctln[4] 1.91e-19
C5516 _101_ _040_ 0.0781f
C5517 cal_count\[2\] VPWR 0.615f
C5518 _122_ a_13356_8457# 4.41e-20
C5519 a_2961_9545# mask\[1\] 1.12e-20
C5520 net55 _100_ 0.253f
C5521 _125_ _123_ 1.37e-21
C5522 _006_ a_1844_9129# 1.26e-19
C5523 a_3431_10933# _042_ 1.4e-19
C5524 _027_ a_9225_2197# 0.0431f
C5525 a_8491_2229# a_9007_2601# 0.106f
C5526 net30 a_9595_5193# 0.00331f
C5527 _008_ a_7548_10217# 1.09e-19
C5528 net46 a_13783_6183# 3.11e-20
C5529 a_6467_9845# a_8992_9955# 1.72e-21
C5530 a_11709_6273# _135_ 1.11e-20
C5531 net44 a_8455_10383# 0.00197f
C5532 net53 _020_ 0.156f
C5533 a_7723_6807# _062_ 6.02e-20
C5534 net43 cal_itt\[1\] 6.61e-21
C5535 mask\[1\] a_1476_7119# 1.87e-20
C5536 net43 a_4512_11305# 0.226f
C5537 a_10688_9295# VPWR 0.267f
C5538 _062_ a_7210_5807# 0.0985f
C5539 _072_ net51 2.5e-20
C5540 mask\[1\] mask\[0\] 0.0883f
C5541 a_745_10933# a_1660_11305# 0.125f
C5542 a_1184_9117# VPWR 0.0791f
C5543 a_8992_9955# VPWR 0.179f
C5544 a_2383_3689# clk 4.67e-19
C5545 a_7197_7119# VPWR 7.1e-20
C5546 _093_ state\[0\] 0.0554f
C5547 net29 _086_ 0.162f
C5548 a_9664_3689# a_9572_2601# 6.38e-21
C5549 trim_mask\[3\] a_11951_2601# 0.00103f
C5550 mask\[6\] mask\[2\] 1.18e-20
C5551 a_4222_7119# _049_ 9.02e-20
C5552 a_12992_8751# a_12061_7669# 1.02e-20
C5553 a_12436_9129# a_12344_8041# 0.00255f
C5554 a_12153_8757# a_12900_7663# 2.36e-20
C5555 a_11233_4405# a_11488_4765# 0.0604f
C5556 mask\[7\] a_1579_11471# 0.0106f
C5557 a_1467_7923# net22 4.37e-22
C5558 a_1095_12393# a_579_10933# 1.17e-20
C5559 mask\[3\] a_3521_9813# 5.12e-21
C5560 _051_ a_5455_4943# 0.0397f
C5561 net16 _135_ 0.00779f
C5562 a_4443_9295# net51 3.21e-20
C5563 clknet_2_2__leaf_clk a_13607_4943# 0.00121f
C5564 a_2910_12131# VPWR 0.00213f
C5565 _107_ a_10055_2767# 1.45e-20
C5566 a_11435_2229# a_12047_2601# 0.00188f
C5567 a_11601_2229# a_11856_2589# 0.0642f
C5568 _104_ clk 0.00692f
C5569 a_9572_2601# a_10689_2223# 1.52e-19
C5570 net45 a_2755_2601# 9.54e-19
C5571 net4 net30 0.0619f
C5572 _046_ a_3852_12381# 1.64e-19
C5573 net29 _102_ 2.32e-20
C5574 a_12410_6031# VPWR 6.25e-20
C5575 calibrate a_7019_4407# 0.0484f
C5576 cal_count\[0\] a_14467_8751# 0.0903f
C5577 net26 net47 0.00334f
C5578 _074_ a_911_6031# 0.0152f
C5579 net35 a_15023_5487# 0.265f
C5580 net52 net51 0.229f
C5581 _099_ a_3667_3829# 6.81e-20
C5582 a_9084_4515# _104_ 0.00161f
C5583 _072_ _003_ 6.33e-20
C5584 net28 a_4621_12393# 8.92e-19
C5585 _054_ a_7891_3617# 0.00299f
C5586 _060_ _089_ 3.49e-19
C5587 calibrate a_4471_4007# 0.0313f
C5588 clknet_2_3__leaf_clk a_9463_8725# 1.9e-20
C5589 _069_ _067_ 0.0468f
C5590 clknet_2_0__leaf_clk a_2877_2197# 0.0196f
C5591 a_3565_7119# VPWR 1.2e-19
C5592 _078_ net45 0.412f
C5593 net46 a_10975_4105# 7.71e-19
C5594 a_7460_5807# _107_ 6.77e-19
C5595 _090_ _097_ 7.45e-19
C5596 net14 a_2014_12381# 2.52e-19
C5597 a_1099_12533# a_1203_12015# 1.74e-19
C5598 net44 a_8381_9295# 0.00334f
C5599 _053_ net42 0.0279f
C5600 a_9374_10383# VPWR 1.98e-19
C5601 clknet_2_1__leaf_clk a_6181_10633# 0.00341f
C5602 _067_ a_8022_7119# 0.00733f
C5603 _097_ a_3847_4438# 1.33e-19
C5604 _074_ _012_ 0.0814f
C5605 _060_ a_4609_1679# 9.79e-21
C5606 clknet_2_1__leaf_clk a_745_12021# 0.0242f
C5607 a_14193_3285# a_14649_3689# 4.2e-19
C5608 a_4815_3031# a_5067_2045# 8.32e-20
C5609 _055_ a_13880_3677# 8.27e-22
C5610 a_13975_3689# a_14237_3677# 0.00171f
C5611 net37 _133_ 2.9e-20
C5612 _120_ _092_ 0.0763f
C5613 net15 a_3123_3615# 0.0144f
C5614 net18 trim_mask\[4\] 0.366f
C5615 net22 _094_ 0.00156f
C5616 a_12691_2527# a_12516_2601# 0.234f
C5617 a_9747_2527# a_9719_1473# 7.73e-20
C5618 _058_ a_14540_3689# 3.95e-19
C5619 _085_ mask\[6\] 0.104f
C5620 _107_ a_6927_3311# 0.0013f
C5621 a_7999_11231# _042_ 2.73e-20
C5622 net33 net49 1.57e-20
C5623 net16 _127_ 0.00342f
C5624 net34 _047_ 0.103f
C5625 _125_ a_13142_8725# 9.71e-21
C5626 a_14807_8359# cal_count\[2\] 8.42e-19
C5627 clknet_2_3__leaf_clk a_14347_4917# 1.26e-21
C5628 net33 a_14733_9545# 0.00159f
C5629 net16 a_14063_7093# 0.0116f
C5630 _108_ net32 2.14e-19
C5631 _064_ a_8491_2229# 5.22e-21
C5632 net28 _101_ 5.23e-20
C5633 _074_ a_5089_10159# 4.39e-19
C5634 cal_count\[1\] VPWR 1.03f
C5635 a_4775_6031# a_5081_4943# 1.22e-20
C5636 _101_ a_5177_9537# 0.00355f
C5637 a_5694_6031# VPWR 2.55e-19
C5638 net46 a_13881_2741# 2.74e-20
C5639 a_5363_4719# _107_ 2.06e-19
C5640 clknet_0_clk a_9459_7895# 1.31e-19
C5641 net16 a_13519_4007# 0.00339f
C5642 a_8307_6575# a_8495_6895# 0.0716f
C5643 _042_ clknet_2_0__leaf_clk 1.44e-20
C5644 a_3781_8207# _121_ 1.99e-19
C5645 net44 clknet_0_clk 0.00545f
C5646 _078_ a_3868_10217# 1.62e-20
C5647 trim_mask\[2\] a_13257_1141# 0.00989f
C5648 a_4775_6031# net55 0.00186f
C5649 _092_ a_11396_6031# 5.82e-21
C5650 _049_ a_6927_3311# 0.033f
C5651 a_8298_2767# net11 2.35e-20
C5652 trim_val\[1\] a_14702_3311# 1.87e-19
C5653 net14 sample 8.01e-20
C5654 VPWR result[3] 0.268f
C5655 clknet_2_3__leaf_clk a_11258_9117# 2.48e-19
C5656 net16 a_14649_6031# 4.92e-19
C5657 net9 _133_ 1.33e-19
C5658 _027_ a_10111_1679# 5.87e-19
C5659 a_9747_2527# a_9595_1679# 0.011f
C5660 _061_ a_15023_5487# 7.29e-19
C5661 a_6909_10933# a_7367_10927# 0.0346f
C5662 a_8731_9295# cal_itt\[0\] 1.64e-19
C5663 a_7618_12015# VPWR 7.19e-19
C5664 a_3852_11293# a_3303_10217# 1.3e-20
C5665 net43 a_7916_8041# 0.258f
C5666 clknet_2_2__leaf_clk a_11488_4765# 0.00253f
C5667 a_10975_4105# a_11343_3317# 0.0111f
C5668 _041_ a_8083_8181# 4.47e-20
C5669 a_6519_3829# _054_ 1.26e-20
C5670 net16 a_14604_3017# 0.00115f
C5671 a_9802_4007# VPWR 0.238f
C5672 net13 _042_ 0.0188f
C5673 _048_ _060_ 0.392f
C5674 a_7250_7485# VPWR 7.67e-19
C5675 clknet_0_clk clk 0.191f
C5676 net12 a_6515_6794# 0.00856f
C5677 net21 a_4621_12393# 5.32e-20
C5678 net28 _086_ 0.106f
C5679 clknet_0_clk en_co_clk 0.0377f
C5680 a_12612_8725# VPWR 0.247f
C5681 _053_ a_8491_2229# 9.79e-21
C5682 _123_ a_13142_8359# 0.0968f
C5683 net54 _015_ 0.00246f
C5684 a_2014_11293# VPWR 0.00178f
C5685 a_3399_2527# VPWR 0.353f
C5686 _131_ net5 0.00988f
C5687 trim_mask\[2\] a_10676_1679# 5.98e-21
C5688 net44 a_7459_7663# 0.00382f
C5689 clknet_2_2__leaf_clk _113_ 0.174f
C5690 a_9084_4515# _110_ 0.106f
C5691 a_13050_7637# a_12900_7663# 0.344f
C5692 a_2313_6183# _049_ 1.37e-19
C5693 _012_ _093_ 0.0256f
C5694 _078_ a_2953_7119# 1.47e-21
C5695 _108_ VPWR 1.68f
C5696 net4 state\[2\] 0.325f
C5697 _050_ net3 0.148f
C5698 clknet_2_3__leaf_clk a_10383_7093# 4.73e-20
C5699 a_1835_11231# result[5] 1.47e-19
C5700 a_9761_1679# a_10752_565# 2.95e-19
C5701 a_4443_1679# a_5067_2045# 9.73e-19
C5702 a_4609_1679# a_4864_1679# 0.0594f
C5703 a_5177_1921# a_5524_1679# 0.0512f
C5704 _074_ a_1129_9813# 0.0091f
C5705 net4 state\[0\] 0.0129f
C5706 a_6741_7361# a_6523_7119# 0.21f
C5707 a_6173_7119# a_7263_7093# 0.0424f
C5708 a_3597_10933# a_3868_10217# 3.1e-20
C5709 _117_ a_11292_1251# 7.35e-20
C5710 _000_ a_6793_8970# 2.8e-20
C5711 a_7477_10901# a_7259_11305# 0.21f
C5712 a_6909_10933# a_7999_11231# 0.0424f
C5713 net30 a_9166_4515# 0.00133f
C5714 net18 a_9195_10357# 3.42e-19
C5715 net13 a_4658_3427# 3.34e-19
C5716 _025_ a_11067_3017# 0.00121f
C5717 a_11244_9661# a_11352_9661# 0.00523f
C5718 net37 _129_ 1.3e-19
C5719 a_13919_8751# a_14467_8751# 3.09e-19
C5720 a_10655_2932# VPWR 0.209f
C5721 net40 a_10975_6031# 4.38e-21
C5722 clknet_2_0__leaf_clk a_1476_6031# 3.1e-19
C5723 a_11067_3017# _026_ 0.11f
C5724 a_11067_4405# a_12323_4703# 0.0435f
C5725 _024_ a_11583_4777# 0.00409f
C5726 a_3748_6281# _090_ 3.1e-19
C5727 net21 _101_ 3.33e-21
C5728 a_2787_10927# VPWR 0.259f
C5729 clknet_2_3__leaf_clk a_11679_4777# 3.69e-20
C5730 net43 a_1375_9129# 0.00156f
C5731 a_9115_2223# VPWR 0.145f
C5732 clknet_2_2__leaf_clk a_8657_2229# 0.0446f
C5733 a_9460_6807# VPWR 0.103f
C5734 _078_ a_3922_8867# 0.00132f
C5735 a_561_4405# a_1476_4777# 0.119f
C5736 mask\[2\] a_3317_8207# 0.00122f
C5737 cal_count\[1\] a_14807_8359# 0.17f
C5738 a_9802_4007# a_9478_4105# 0.0153f
C5739 a_10781_3311# a_9761_1679# 5.17e-22
C5740 a_4725_5487# VPWR 0.0042f
C5741 net28 _022_ 8.53e-19
C5742 VPWR en 0.243f
C5743 _094_ a_4871_6031# 0.00511f
C5744 a_4259_6031# a_4883_6397# 9.73e-19
C5745 a_4425_6031# a_4680_6031# 0.0642f
C5746 clknet_2_1__leaf_clk a_7613_8029# 1.33e-20
C5747 a_10787_1135# a_10752_565# 4.68e-19
C5748 _057_ a_14471_591# 0.0648f
C5749 a_6927_591# ctln[5] 2.68e-20
C5750 cal_count\[0\] a_14249_8725# 0.115f
C5751 a_10111_1679# _117_ 1.78e-19
C5752 _042_ a_4864_9295# 2.87e-20
C5753 a_3891_4943# a_4091_5309# 0.145f
C5754 net46 a_9099_3689# 0.152f
C5755 a_11987_8757# a_13184_9117# 1.63e-19
C5756 net43 a_4209_12381# 0.00191f
C5757 _125_ a_14335_7895# 0.001f
C5758 cal_itt\[0\] a_9621_8029# 4.2e-20
C5759 _087_ a_5731_4943# 9.6e-20
C5760 _108_ a_9478_4105# 0.0111f
C5761 a_11023_5108# trim_mask\[4\] 1.36e-21
C5762 net45 _004_ 0.00493f
C5763 net27 a_7618_12015# 8.03e-20
C5764 a_5423_9011# mask\[1\] 9.85e-20
C5765 a_10990_7485# a_11297_7119# 3.69e-19
C5766 a_11059_7356# a_11369_7119# 0.0138f
C5767 net16 _041_ 0.0115f
C5768 _078_ a_2857_5461# 1.16e-19
C5769 clknet_0_clk a_8091_7967# 0.00155f
C5770 net13 a_5177_1921# 0.00583f
C5771 net26 _072_ 1.07e-20
C5772 net36 _126_ 6.86e-20
C5773 _048_ a_7939_3855# 0.00273f
C5774 net46 a_12047_2601# 9.54e-19
C5775 a_9004_3677# VPWR 0.0833f
C5776 net12 a_6743_10933# 5.32e-19
C5777 a_2092_8457# net23 0.17f
C5778 a_8178_11293# VPWR 3.61e-19
C5779 cal_itt\[2\] a_8820_6005# 0.137f
C5780 a_12516_2601# VPWR 0.307f
C5781 net43 a_4995_7119# 0.0499f
C5782 a_763_8757# a_816_7119# 5.28e-21
C5783 a_8083_8181# _002_ 0.107f
C5784 net31 a_14972_5193# 4.7e-19
C5785 net26 _068_ 3.89e-20
C5786 a_8992_9955# a_8381_9295# 1.58e-19
C5787 _048_ a_4498_4373# 4.6e-19
C5788 trim_mask\[4\] a_10055_2767# 0.00133f
C5789 _135_ clkc 2.25e-19
C5790 a_4471_4007# _015_ 0.113f
C5791 en_co_clk a_14564_6397# 0.195f
C5792 _107_ VPWR 1.04f
C5793 net45 ctln[7] 3.98e-19
C5794 a_6763_5193# state\[2\] 3.98e-20
C5795 a_2828_12131# mask\[6\] 6.03e-19
C5796 a_3431_12021# a_4512_12393# 0.102f
C5797 net2 a_10864_7387# 1.14e-20
C5798 a_4165_11989# a_3947_12393# 0.21f
C5799 a_3597_12021# a_4687_12319# 0.0423f
C5800 _072_ a_7262_5461# 5.62e-20
C5801 net30 a_3057_4719# 7.26e-20
C5802 a_13142_8725# a_13142_8359# 0.0121f
C5803 clknet_0_clk _059_ 0.0276f
C5804 _101_ _020_ 0.00744f
C5805 net26 a_4443_9295# 1.42e-20
C5806 _032_ a_10851_1653# 1.97e-20
C5807 a_5524_1679# a_5633_1679# 0.00742f
C5808 a_5699_1653# a_5878_1679# 0.0074f
C5809 a_9595_1679# a_10676_1679# 0.102f
C5810 _131_ a_15023_6031# 7.53e-22
C5811 a_5363_12559# a_6191_12559# 1.13e-19
C5812 mask\[5\] a_3431_10933# 2.2e-21
C5813 net15 a_3529_6281# 0.00108f
C5814 _065_ net51 0.153f
C5815 _106_ a_9503_4399# 0.206f
C5816 net46 a_10018_3677# 0.00196f
C5817 net52 net26 0.0105f
C5818 clknet_2_1__leaf_clk _082_ 0.00131f
C5819 net12 net45 0.0673f
C5820 net15 a_3303_10217# 0.00541f
C5821 _034_ a_4775_6031# 0.00142f
C5822 a_12900_7663# VPWR 0.427f
C5823 _049_ VPWR 1.51f
C5824 _081_ a_2971_8457# 2.76e-19
C5825 a_579_10933# a_1461_10357# 1.02e-19
C5826 clknet_2_3__leaf_clk a_8215_9295# 0.851f
C5827 a_3388_4631# VPWR 0.107f
C5828 a_5699_1653# VPWR 0.405f
C5829 net27 a_2787_10927# 2.01e-19
C5830 _126_ _128_ 3.32e-19
C5831 _038_ a_11067_4405# 2.98e-20
C5832 net47 a_11297_7119# 0.00316f
C5833 a_7259_11305# VPWR 0.214f
C5834 net29 _046_ 0.00419f
C5835 _044_ net12 4.19e-20
C5836 trim_mask\[4\] a_6927_3311# 0.11f
C5837 a_9839_3615# a_10699_3311# 1.8e-20
C5838 mask\[1\] a_1125_7663# 0.0552f
C5839 a_2092_8457# a_2225_7663# 5.91e-20
C5840 mask\[0\] _050_ 9.79e-21
C5841 trim_mask\[0\] a_13697_4373# 0.112f
C5842 a_8495_6895# VPWR 0.00277f
C5843 mask\[1\] a_2489_7983# 9.32e-19
C5844 net41 clk 3.86e-20
C5845 net46 trim_val\[4\] 0.00883f
C5846 net14 a_1173_4765# 5.85e-19
C5847 en_co_clk net41 3.57e-19
C5848 trim_mask\[1\] _112_ 0.216f
C5849 net21 a_6375_12021# 2.25e-21
C5850 net44 a_6523_7119# 0.154f
C5851 _092_ _051_ 0.0918f
C5852 _107_ a_9478_4105# 0.00129f
C5853 _104_ a_9802_4007# 1.94e-19
C5854 cal_count\[0\] _001_ 4.97e-19
C5855 a_455_8181# _005_ 7.02e-19
C5856 _113_ a_14540_3689# 3.38e-21
C5857 a_1313_11989# _086_ 1.62e-19
C5858 _065_ _003_ 0.0016f
C5859 a_9595_5193# _118_ 7.13e-19
C5860 net40 a_15023_5487# 0.0147f
C5861 _026_ a_11856_2589# 0.16f
C5862 net13 a_5633_1679# 1.14e-19
C5863 _092_ _014_ 0.00462f
C5864 _088_ a_5931_4105# 1.01e-19
C5865 clknet_2_1__leaf_clk a_1007_10217# 9.94e-19
C5866 a_1095_12393# result[6] 8.65e-19
C5867 net47 _036_ 0.0224f
C5868 _128_ a_12153_8757# 8.08e-20
C5869 a_3947_12393# VPWR 0.227f
C5870 a_8072_11721# a_7723_10143# 6.2e-22
C5871 _108_ _104_ 0.0175f
C5872 a_11233_4405# a_10975_4105# 2.86e-20
C5873 net50 a_10676_1679# 0.0118f
C5874 a_3431_12021# _046_ 0.0294f
C5875 clknet_2_2__leaf_clk a_10329_1921# 2.9e-19
C5876 a_1476_7119# a_561_6031# 5.24e-20
C5877 a_911_7119# a_911_6031# 8.87e-19
C5878 a_561_7119# a_1476_6031# 6.41e-22
C5879 mask\[1\] a_4871_8181# 0.0914f
C5880 net43 a_1203_10927# 0.0139f
C5881 mask\[0\] a_561_6031# 0.00201f
C5882 _076_ mask\[1\] 2.4e-19
C5883 a_13470_7663# _133_ 0.00808f
C5884 net28 a_4512_12393# 0.044f
C5885 mask\[6\] a_4609_9295# 5.57e-22
C5886 _090_ a_4308_4917# 5.02e-20
C5887 a_3425_11721# VPWR 0.261f
C5888 a_4259_6031# a_4993_6273# 0.0701f
C5889 _094_ _075_ 1.22e-19
C5890 net30 _064_ 0.184f
C5891 _123_ a_13557_8457# 4.54e-20
C5892 a_6523_7119# clk 3.57e-21
C5893 net9 a_12533_3689# 1.84e-20
C5894 net46 a_14281_4943# 2.95e-19
C5895 a_13919_8751# a_14249_8725# 0.0184f
C5896 net45 a_1830_7119# 5.4e-19
C5897 a_455_3571# a_995_3530# 0.00329f
C5898 _104_ a_10655_2932# 0.0245f
C5899 cal_itt\[3\] _051_ 3.84e-20
C5900 a_7184_2339# _027_ 1.93e-19
C5901 _101_ a_2143_7663# 0.142f
C5902 _083_ a_6633_9845# 5.05e-19
C5903 a_6467_9845# _008_ 0.279f
C5904 a_14347_4917# _047_ 1.23e-20
C5905 clknet_2_3__leaf_clk a_8298_5487# 1.62f
C5906 a_6191_12559# ctlp[6] 0.001f
C5907 net4 _118_ 0.00759f
C5908 a_9020_10383# _042_ 0.0531f
C5909 VPWR trimb[2] 0.581f
C5910 a_1461_10357# a_395_9845# 0.0015f
C5911 _043_ a_9871_10383# 0.194f
C5912 net13 a_4959_9295# 0.00836f
C5913 mask\[5\] a_7999_11231# 0.0652f
C5914 _103_ a_7190_3855# 3.65e-19
C5915 _104_ a_9115_2223# 6.03e-20
C5916 net9 a_12323_4703# 0.0171f
C5917 a_1867_3317# cal 8.2e-19
C5918 cal_count\[2\] a_14564_6397# 3.89e-19
C5919 a_10838_2045# VPWR 8.38e-19
C5920 cal_itt\[0\] _122_ 6.25e-20
C5921 net43 a_3431_10933# 0.313f
C5922 _008_ VPWR 0.534f
C5923 net43 a_929_8757# 0.031f
C5924 a_579_10933# a_745_10933# 0.883f
C5925 net27 a_7259_11305# 2e-19
C5926 net35 trim_val\[0\] 0.138f
C5927 a_13703_4943# _058_ 8.33e-19
C5928 trim_val\[0\] a_13059_4631# 3.87e-19
C5929 _097_ a_3667_3829# 0.00108f
C5930 _033_ a_9747_2527# 1.15e-20
C5931 trim_val\[4\] a_11343_3317# 3.04e-21
C5932 cal_itt\[0\] _063_ 0.357f
C5933 _051_ a_9317_3285# 1.05e-20
C5934 a_561_6031# _079_ 4.88e-19
C5935 net25 a_3303_10217# 2.89e-20
C5936 _050_ net54 2.65e-19
C5937 a_11987_8757# a_12061_7669# 0.00126f
C5938 a_12153_8757# a_11895_7669# 0.00117f
C5939 a_395_4405# a_937_4105# 1.46e-19
C5940 _072_ cal_itt\[2\] 0.145f
C5941 net16 a_14526_4943# 2.04e-19
C5942 net19 a_9459_7895# 0.00225f
C5943 _008_ a_5699_9269# 4.31e-20
C5944 a_3597_10933# a_4621_11305# 2.36e-20
C5945 a_4165_10901# a_4209_11293# 3.69e-19
C5946 _053_ net30 0.173f
C5947 a_395_6031# a_455_5747# 0.0123f
C5948 a_2767_2223# clk 0.00154f
C5949 a_5423_9011# _041_ 0.0753f
C5950 _104_ a_9004_3677# 2.61e-19
C5951 a_2014_12381# VPWR 0.00178f
C5952 _112_ _115_ 0.00388f
C5953 _093_ a_3933_2767# 2.98e-20
C5954 net19 net44 0.0822f
C5955 _027_ a_9734_2223# 3.05e-19
C5956 trim_mask\[0\] a_13825_5185# 0.0255f
C5957 _068_ cal_itt\[2\] 0.0725f
C5958 a_395_9845# _018_ 2.75e-21
C5959 _040_ a_3053_8207# 0.00443f
C5960 net26 a_1679_10633# 6.75e-19
C5961 _059_ net41 0.174f
C5962 _110_ a_9802_4007# 0.00639f
C5963 a_3947_12393# net27 2.25e-20
C5964 a_5524_9295# VPWR 0.31f
C5965 net54 _052_ 1.63e-20
C5966 _107_ _104_ 0.0234f
C5967 net28 _046_ 0.389f
C5968 mask\[5\] net13 9.08e-20
C5969 a_11396_6031# _136_ 0.00158f
C5970 calibrate net1 0.00394f
C5971 a_7631_12319# a_6909_10933# 1.08e-19
C5972 clknet_2_3__leaf_clk _135_ 0.194f
C5973 net54 _098_ 1.04e-19
C5974 _108_ _110_ 0.0421f
C5975 a_7001_7669# a_8022_7119# 0.00157f
C5976 trim_mask\[1\] a_12121_3677# 4.53e-21
C5977 _071_ a_6173_7119# 6.82e-21
C5978 a_7351_8041# a_7263_7093# 1.1e-19
C5979 trim_mask\[2\] a_12213_2589# 9.76e-20
C5980 a_5177_9537# a_5067_9661# 0.0977f
C5981 a_5699_9269# a_5524_9295# 0.234f
C5982 a_4959_9295# a_4864_9295# 0.0498f
C5983 clknet_2_2__leaf_clk a_10975_4105# 0.0116f
C5984 _030_ a_13880_3677# 0.158f
C5985 net21 a_4512_12393# 0.00661f
C5986 net27 a_3425_11721# 2.1e-19
C5987 a_9459_7895# cal_itt\[1\] 0.215f
C5988 clknet_0_clk _108_ 1.25e-20
C5989 _014_ cal 3e-20
C5990 a_11394_9509# cal_count\[0\] 0.00246f
C5991 net47 a_8636_9295# 2.48e-19
C5992 net12 a_6316_5193# 0.0104f
C5993 trim_val\[1\] a_14099_3017# 0.0585f
C5994 a_4687_11231# a_4512_11305# 0.234f
C5995 net19 clk 0.039f
C5996 net37 cal_count\[0\] 2.9e-19
C5997 _101_ _077_ 0.00277f
C5998 net19 en_co_clk 0.00479f
C5999 a_7569_7637# _063_ 4.1e-20
C6000 a_10975_6031# a_13349_6031# 6.92e-21
C6001 net45 a_2309_2229# 0.0265f
C6002 _049_ _104_ 0.307f
C6003 a_4655_10071# mask\[2\] 0.00222f
C6004 net25 a_455_8181# 2.02e-20
C6005 _123_ a_12916_8751# 0.00243f
C6006 _129_ a_13470_7663# 4.04e-19
C6007 net52 a_2961_9295# 7e-19
C6008 a_11856_2589# _031_ 3.97e-20
C6009 net14 a_1173_7119# 5.85e-19
C6010 _128_ a_13050_7637# 3.45e-20
C6011 a_13697_4373# _030_ 2.45e-19
C6012 _107_ a_7200_3631# 2.81e-19
C6013 _058_ a_13459_3317# 0.00266f
C6014 a_3303_7119# a_3411_7485# 0.0572f
C6015 clknet_2_0__leaf_clk a_2601_3285# 6.07e-21
C6016 a_5915_10927# _042_ 5.22e-20
C6017 _048_ a_4175_4943# 0.00535f
C6018 net19 a_9084_4515# 0.00778f
C6019 _110_ a_10655_2932# 7.08e-22
C6020 VPWR sample 0.531f
C6021 _051_ a_6737_4719# 1.36e-20
C6022 trim_mask\[4\] VPWR 1.13f
C6023 a_7824_11305# _020_ 0.00287f
C6024 a_448_6549# a_561_6031# 2.18e-19
C6025 a_745_10933# a_395_9845# 1.33e-20
C6026 a_10699_5487# _108_ 6.25e-19
C6027 net3 a_395_2767# 0.108f
C6028 _108_ a_12148_4777# 1.55e-19
C6029 net9 _038_ 1.21e-20
C6030 _122_ a_13092_8029# 7.52e-20
C6031 _051_ a_5547_5603# 0.2f
C6032 a_7527_4631# _088_ 0.0915f
C6033 net3 a_455_3571# 9.02e-19
C6034 a_1129_7361# a_1585_7119# 4.2e-19
C6035 net34 a_14172_1513# 0.00409f
C6036 net27 _008_ 9.66e-23
C6037 a_763_8757# net23 3.7e-20
C6038 clknet_2_0__leaf_clk _039_ 0.00324f
C6039 a_7262_5461# a_7527_4631# 4.59e-21
C6040 _050_ a_7019_4407# 0.00933f
C6041 cal_count\[0\] a_11116_8983# 0.319f
C6042 clknet_0_clk a_9460_6807# 1.29e-19
C6043 _046_ a_4167_11471# 0.203f
C6044 net15 a_579_12021# 1.97e-21
C6045 a_1476_10217# a_3208_10205# 2e-21
C6046 a_6796_12381# ctlp[6] 7.83e-20
C6047 _078_ a_2787_9845# 6.69e-19
C6048 _049_ a_7200_3631# 0.00256f
C6049 _090_ a_3847_4438# 0.00106f
C6050 _058_ _109_ 0.0221f
C6051 cal_itt\[1\] clk 1.25e-20
C6052 cal_itt\[1\] en_co_clk 0.133f
C6053 net34 a_15159_9269# 0.0108f
C6054 mask\[7\] a_1764_10383# 0.00918f
C6055 net14 a_1201_3855# 7.15e-19
C6056 net43 clknet_2_0__leaf_clk 0.373f
C6057 _063_ trim_mask\[0\] 0.271f
C6058 _048_ a_7571_4943# 0.0537f
C6059 a_13607_4943# a_13703_4943# 0.0138f
C6060 a_13825_5185# a_13869_4943# 3.69e-19
C6061 a_13257_4943# trim_val\[0\] 1.93e-19
C6062 net14 a_1019_9839# 0.00145f
C6063 a_12516_2601# a_12678_2223# 0.00645f
C6064 net26 _065_ 2.68e-20
C6065 net45 a_7524_2223# 0.0135f
C6066 net9 cal_count\[0\] 0.045f
C6067 _051_ a_5536_4399# 0.0135f
C6068 _006_ _080_ 9.8e-20
C6069 a_455_8181# a_395_7119# 3.92e-20
C6070 _056_ _114_ 1.67e-19
C6071 cal_itt\[1\] a_9084_4515# 8.13e-20
C6072 a_8215_9295# a_8827_9295# 0.00188f
C6073 a_395_9845# a_1387_8751# 6.14e-21
C6074 a_6056_8359# net2 0.188f
C6075 mask\[6\] a_6181_10633# 1.44e-19
C6076 a_455_5747# net30 0.246f
C6077 _052_ a_7019_4407# 4.47e-19
C6078 net15 a_2869_10927# 0.00109f
C6079 clknet_2_1__leaf_clk a_4165_10901# 6.93e-20
C6080 a_4036_8207# VPWR 0.0828f
C6081 net43 a_4687_12319# 0.272f
C6082 clknet_2_1__leaf_clk a_6541_12021# 0.0256f
C6083 _048_ a_4576_3427# 8.76e-22
C6084 _041_ a_4871_8181# 1.05e-19
C6085 _110_ a_12516_2601# 2.85e-19
C6086 a_8072_11721# _042_ 1.02e-20
C6087 a_9443_6059# cal_count\[3\] 3.92e-20
C6088 _098_ a_7019_4407# 0.0229f
C6089 a_15023_2223# trim[0] 9.86e-19
C6090 _076_ _041_ 0.0928f
C6091 net21 _046_ 0.0125f
C6092 net14 ctlp[0] 0.0159f
C6093 net36 VPWR 0.383f
C6094 trim_mask\[2\] a_9595_1679# 3.11e-19
C6095 a_9664_3689# _032_ 3.86e-21
C6096 _053_ state\[2\] 0.13f
C6097 _107_ _110_ 0.0146f
C6098 a_9478_4105# trim_mask\[4\] 5.72e-20
C6099 a_11895_7669# a_13050_7637# 0.0608f
C6100 _037_ a_12344_8041# 0.00265f
C6101 _078_ a_2092_8457# 0.00199f
C6102 a_561_4405# _014_ 0.00248f
C6103 net43 net13 0.127f
C6104 clknet_0_clk _107_ 0.039f
C6105 net45 a_3110_3311# 3.67e-19
C6106 _053_ state\[0\] 0.0174f
C6107 a_2787_7119# a_3977_7119# 2.56e-19
C6108 a_6891_12393# VPWR 0.195f
C6109 a_5363_7369# a_6173_7119# 3.15e-19
C6110 _001_ en_co_clk 6.44e-20
C6111 _075_ _096_ 5.91e-20
C6112 a_3597_10933# a_2787_9845# 5.65e-19
C6113 net33 _031_ 2.32e-21
C6114 _121_ a_4425_6031# 7.28e-19
C6115 a_3431_10933# a_2953_9845# 2.01e-19
C6116 _042_ a_4043_10143# 0.0066f
C6117 _074_ a_4443_9295# 0.00841f
C6118 a_5915_10927# a_6909_10933# 2.84e-19
C6119 a_3123_3615# VPWR 0.375f
C6120 a_8386_8457# _001_ 1.78e-20
C6121 a_12061_7669# cal_count\[3\] 1.07e-20
C6122 _130_ _134_ 0.00574f
C6123 a_6927_591# a_8767_591# 4.72e-21
C6124 net3 _099_ 0.0116f
C6125 a_5536_4399# a_5445_4399# 0.00145f
C6126 clknet_0_clk _049_ 0.0925f
C6127 net4 a_3933_2767# 0.0493f
C6128 a_1007_10217# result[4] 3.91e-19
C6129 a_13607_4943# a_13459_3317# 2.44e-21
C6130 a_3840_8867# a_3781_8207# 0.00162f
C6131 _074_ net52 0.0103f
C6132 _101_ a_6173_7119# 0.00382f
C6133 _074_ a_816_7119# 0.00411f
C6134 clknet_2_2__leaf_clk a_7223_2465# 0.274f
C6135 a_9195_10357# VPWR 0.364f
C6136 a_7916_8041# a_9459_7895# 5.62e-20
C6137 _078_ a_2198_9117# 0.00213f
C6138 _108_ a_13091_4943# 0.445f
C6139 _078_ net51 0.00111f
C6140 net44 a_7916_8041# 9.86e-21
C6141 a_1467_7923# a_1476_6031# 4.94e-22
C6142 net45 a_1651_6005# 0.291f
C6143 _128_ VPWR 0.684f
C6144 trim_val\[1\] net48 9.98e-21
C6145 _122_ a_11258_8790# 7.33e-19
C6146 a_15259_7637# comp 0.233f
C6147 net55 a_5931_4105# 6.38e-20
C6148 net47 net4 0.0335f
C6149 cal_count\[0\] a_12436_9129# 0.0503f
C6150 net45 a_4609_1679# 0.026f
C6151 clknet_0_clk a_8495_6895# 2.56e-19
C6152 a_10851_1653# a_11030_1679# 0.0074f
C6153 a_10676_1679# a_10785_1679# 0.00742f
C6154 a_9595_1679# a_9719_1473# 0.00105f
C6155 _067_ a_10055_5487# 0.103f
C6156 net37 a_13919_8751# 1.83e-21
C6157 clknet_2_0__leaf_clk a_2857_7637# 0.0448f
C6158 net40 a_15023_8751# 0.246f
C6159 clknet_2_3__leaf_clk a_13279_7119# 1.91e-20
C6160 net43 a_1203_12015# 0.0139f
C6161 net19 a_8992_9955# 0.013f
C6162 a_4512_11305# a_4801_9839# 5.3e-21
C6163 net45 a_816_4765# 2.47e-19
C6164 net18 net40 0.0116f
C6165 a_4055_12015# _078_ 4.99e-19
C6166 clknet_2_2__leaf_clk a_9099_3689# 0.00149f
C6167 net12 a_6210_4989# 0.0098f
C6168 net50 trim_mask\[2\] 0.00675f
C6169 net14 a_1493_5487# 0.00505f
C6170 _063_ a_8949_6281# 0.0069f
C6171 a_3868_7119# _121_ 1.8e-19
C6172 a_14335_4020# a_13975_3689# 0.00125f
C6173 net46 a_14702_3311# 2.06e-19
C6174 a_2019_9055# mask\[0\] 1.94e-19
C6175 a_15023_2767# a_15023_2223# 0.0523f
C6176 _040_ net45 0.0264f
C6177 a_7320_3631# VPWR 1.63e-19
C6178 a_395_2767# valid 9.25e-19
C6179 net47 a_8360_10383# 2.46e-19
C6180 a_8673_10625# a_8563_10749# 0.0977f
C6181 _120_ a_3365_4943# 3.38e-19
C6182 a_3063_591# clk 0.00341f
C6183 net14 a_579_12021# 0.00552f
C6184 a_1099_12533# _011_ 1.29e-19
C6185 _023_ a_763_8757# 1.73e-22
C6186 a_455_3571# valid 0.336f
C6187 _077_ a_6515_8534# 2.83e-20
C6188 a_14347_4917# net49 1.28e-21
C6189 a_7916_8041# clk 0.00238f
C6190 net4 a_8820_6005# 0.00116f
C6191 VPWR ctlp[5] 0.353f
C6192 net42 a_8473_5193# 0.0041f
C6193 _076_ _002_ 1.23e-19
C6194 a_855_4105# _013_ 2.65e-19
C6195 a_7631_12319# mask\[5\] 5.46e-20
C6196 a_3530_4765# VPWR 4.61e-20
C6197 _074_ a_7153_12381# 2.48e-21
C6198 a_561_7119# _039_ 4.38e-19
C6199 _075_ a_5455_4943# 0.0637f
C6200 trim_val\[3\] a_10752_565# 0.0101f
C6201 a_1476_6031# _094_ 3.31e-23
C6202 clknet_2_3__leaf_clk _041_ 0.011f
C6203 a_4863_4917# a_4617_4105# 2.02e-20
C6204 net13 a_2857_7637# 2.91e-19
C6205 a_10864_7387# a_11059_7356# 0.23f
C6206 a_6741_7361# a_6619_7119# 3.16e-19
C6207 a_10586_7371# a_10990_7485# 0.0512f
C6208 a_10195_1354# _057_ 6.35e-20
C6209 a_11292_1251# _116_ 3.67e-20
C6210 net53 a_7548_10217# 0.00102f
C6211 clknet_2_1__leaf_clk a_7569_7637# 3.05e-20
C6212 _104_ trim_mask\[4\] 0.297f
C6213 a_12723_4943# VPWR 0.257f
C6214 a_6891_12393# net27 2.14e-19
C6215 a_11509_3317# a_12424_3689# 0.119f
C6216 a_8949_9537# VPWR 0.213f
C6217 _042_ a_3208_10205# 2.86e-19
C6218 net43 a_561_7119# 0.0431f
C6219 trim_val\[2\] trim[3] 8.5e-19
C6220 a_14715_3615# a_14604_3017# 2.46e-19
C6221 net44 a_7442_7119# 0.00288f
C6222 cal_count\[0\] a_11508_9295# 9.23e-20
C6223 a_14099_3017# a_14184_2767# 1.48e-19
C6224 mask\[4\] a_5089_10159# 0.00184f
C6225 _023_ net26 0.0652f
C6226 net35 net32 2.58e-19
C6227 a_816_10205# a_763_8757# 1.58e-20
C6228 a_13697_4373# a_15083_4659# 2.75e-20
C6229 _058_ a_14655_4399# 0.196f
C6230 net31 a_14981_4020# 0.149f
C6231 a_11895_7669# VPWR 0.437f
C6232 _067_ trim_val\[4\] 0.00182f
C6233 a_4259_6031# net3 6.19e-19
C6234 net50 a_11045_3631# 1.65e-19
C6235 net40 trim_val\[0\] 3.63e-20
C6236 _134_ a_13821_7119# 1.68e-19
C6237 a_1173_4765# VPWR 4.89e-19
C6238 _056_ VPWR 0.517f
C6239 a_6835_7669# a_7256_8029# 0.0867f
C6240 _129_ a_14788_7369# 4.36e-19
C6241 _063_ a_8307_4943# 0.171f
C6242 a_2953_9845# clknet_2_0__leaf_clk 9.79e-21
C6243 _065_ cal_itt\[2\] 0.00575f
C6244 net50 a_9719_1473# 4.67e-19
C6245 net45 _048_ 4.74e-19
C6246 a_5496_12131# a_5578_12131# 0.00477f
C6247 _101_ a_3852_11293# 2e-19
C6248 _044_ a_8767_11471# 0.195f
C6249 trim_mask\[4\] a_7200_3631# 3.96e-19
C6250 _048_ _058_ 2.11e-19
C6251 a_3781_8207# a_4131_8207# 0.217f
C6252 a_3615_8207# a_4871_8181# 0.0436f
C6253 a_10111_1679# _116_ 0.00144f
C6254 _032_ _057_ 3.05e-20
C6255 _064_ _118_ 0.0875f
C6256 _076_ a_3615_8207# 2.2e-21
C6257 a_14249_8725# cal_count\[1\] 0.00317f
C6258 a_3891_4943# state\[0\] 3.6e-21
C6259 net37 en_co_clk 1.95e-19
C6260 a_395_6031# a_395_4405# 2.09e-19
C6261 a_11491_6031# VPWR 0.204f
C6262 mask\[3\] a_929_8757# 1.96e-19
C6263 a_10188_4105# a_10270_4105# 0.00477f
C6264 _067_ a_9823_6941# 0.0061f
C6265 net44 a_4995_7119# 0.156f
C6266 a_10688_9295# _001_ 2.17e-20
C6267 clknet_2_3__leaf_clk a_10781_5487# 7.57e-20
C6268 _113_ a_13459_3317# 0.0141f
C6269 mask\[4\] a_6633_9845# 0.0256f
C6270 _126_ net40 0.234f
C6271 clknet_2_2__leaf_clk trim_val\[4\] 1.6e-19
C6272 net43 a_4239_8573# 2.97e-20
C6273 a_2309_2229# a_3386_2223# 1.46e-19
C6274 cal_count\[3\] a_11396_6031# 0.0163f
C6275 net47 a_10586_7371# 0.254f
C6276 net18 _024_ 0.029f
C6277 clknet_2_1__leaf_clk a_7723_10143# 0.00123f
C6278 a_11967_3311# VPWR 0.133f
C6279 trim_mask\[3\] ctln[4] 1.69e-19
C6280 _108_ a_11057_4105# 7.11e-19
C6281 a_8091_7967# a_7916_8041# 0.234f
C6282 _063_ a_7723_6807# 3.84e-19
C6283 net13 a_2953_9845# 1.73e-20
C6284 _101_ a_3947_11305# 2.6e-19
C6285 a_2601_3285# a_2948_3689# 0.0512f
C6286 a_2033_3317# a_4576_3427# 2.13e-20
C6287 net50 a_9595_1679# 0.00398f
C6288 _074_ a_1679_10633# 0.0564f
C6289 a_6419_8207# VPWR 7.04e-19
C6290 net35 VPWR 0.519f
C6291 a_13059_4631# VPWR 0.22f
C6292 _037_ _133_ 0.0115f
C6293 _109_ _113_ 3.58e-19
C6294 a_1129_4373# valid 9.39e-19
C6295 net46 ctln[3] 4.12e-20
C6296 trim_mask\[2\] a_14604_2339# 0.101f
C6297 a_7456_12393# _020_ 6.99e-22
C6298 _049_ net41 0.0018f
C6299 _136_ a_11801_4373# 9.25e-19
C6300 a_4995_7119# en_co_clk 1.91e-21
C6301 net9 en_co_clk 0.0171f
C6302 a_11509_3317# a_11435_2229# 9.64e-20
C6303 clknet_2_1__leaf_clk a_1476_10217# 0.0679f
C6304 trim_val\[1\] trim[0] 0.00247f
C6305 _053_ _118_ 1.98e-19
C6306 a_8761_7983# VPWR 1.33e-19
C6307 net55 a_7527_4631# 0.0971f
C6308 net46 a_14237_3677# 0.00322f
C6309 a_5081_4943# state\[1\] 4.89e-22
C6310 _070_ net2 0.38f
C6311 clknet_2_1__leaf_clk _007_ 0.233f
C6312 mask\[5\] a_5915_10927# 0.101f
C6313 net40 a_11023_5108# 0.0347f
C6314 _110_ trim_mask\[4\] 0.0431f
C6315 net19 _108_ 8.39e-19
C6316 _065_ a_11297_7119# 3.02e-20
C6317 net55 state\[1\] 0.0176f
C6318 _020_ _043_ 2.16e-21
C6319 clknet_0_clk trim_mask\[4\] 0.0177f
C6320 a_3529_6281# VPWR 0.00643f
C6321 _111_ a_12599_3615# 2.19e-19
C6322 a_3303_10217# VPWR 0.216f
C6323 a_7939_10383# a_8673_10625# 0.0701f
C6324 net43 a_4167_6575# 0.0336f
C6325 trim_mask\[2\] a_14193_3285# 4.36e-20
C6326 _122_ a_12344_8041# 0.00178f
C6327 a_8583_3317# a_8491_2229# 4.35e-20
C6328 _058_ trim[1] 0.00145f
C6329 _095_ a_1476_4777# 7.61e-19
C6330 _064_ a_10137_4943# 0.00201f
C6331 net42 a_7190_3855# 7.65e-19
C6332 _051_ a_7010_3311# 0.00143f
C6333 net51 a_7001_7669# 0.00359f
C6334 _065_ net55 7.5e-20
C6335 a_6523_7119# _049_ 3.01e-20
C6336 net19 a_10655_2932# 1.78e-22
C6337 _078_ a_763_8757# 0.0158f
C6338 a_1651_10143# a_2787_9845# 5.37e-21
C6339 a_1476_10217# a_2368_9955# 3.64e-19
C6340 a_4655_10071# a_4609_9295# 3.05e-19
C6341 net44 a_6619_7119# 9.54e-19
C6342 net54 _087_ 9.31e-20
C6343 a_7527_4631# a_7715_3285# 3.67e-21
C6344 calibrate a_2143_2229# 4.43e-22
C6345 a_10699_5487# trim_mask\[4\] 1.27e-19
C6346 a_3521_7361# _120_ 2.43e-20
C6347 a_3431_10933# a_4043_11305# 3.82e-19
C6348 _022_ a_3852_11293# 0.158f
C6349 a_14335_4020# trim_val\[1\] 1.75e-20
C6350 _104_ a_7320_3631# 4.85e-19
C6351 a_6927_12559# a_6541_12021# 0.00122f
C6352 net38 VPWR 0.411f
C6353 _097_ a_3339_2767# 2.22e-19
C6354 net19 a_9115_2223# 0.00323f
C6355 a_6633_9845# a_7091_9839# 0.0276f
C6356 a_9007_2601# a_9103_2601# 0.0138f
C6357 a_9225_2197# a_9269_2589# 3.69e-19
C6358 net30 a_395_4405# 8.1e-21
C6359 net19 a_9460_6807# 7.11e-20
C6360 _111_ a_12257_4777# 1.58e-19
C6361 a_455_5747# _012_ 1.46e-19
C6362 cal_itt\[2\] _067_ 3.46e-19
C6363 net55 a_5054_4399# 0.00257f
C6364 _061_ VPWR 0.248f
C6365 _068_ net4 0.00707f
C6366 mask\[0\] a_4259_6031# 7.17e-20
C6367 _074_ _065_ 0.0585f
C6368 _101_ _005_ 2.24e-20
C6369 mask\[3\] clknet_2_0__leaf_clk 1.61e-20
C6370 net13 a_4617_4105# 0.00326f
C6371 _033_ trim_mask\[2\] 0.00893f
C6372 a_10864_7387# a_11016_6691# 7.13e-21
C6373 net12 net51 0.0437f
C6374 net54 _099_ 0.0742f
C6375 clknet_2_0__leaf_clk a_6741_7361# 2.53e-19
C6376 cal_itt\[0\] _092_ 0.0807f
C6377 mask\[5\] a_8072_11721# 0.231f
C6378 net4 a_395_591# 0.109f
C6379 net37 cal_count\[2\] 1.17e-19
C6380 net34 _031_ 7.71e-23
C6381 _078_ net26 0.062f
C6382 _074_ net23 0.211f
C6383 a_1173_7119# VPWR 4.2e-19
C6384 a_9195_10357# a_8381_9295# 3.34e-19
C6385 a_8455_10383# a_8949_9537# 4.73e-19
C6386 _090_ a_3667_3829# 0.00462f
C6387 calibrate a_4815_3031# 1.25e-21
C6388 net15 _101_ 0.749f
C6389 a_455_8181# VPWR 0.438f
C6390 _082_ a_1763_9295# 0.00151f
C6391 net47 _000_ 0.00829f
C6392 a_10405_9295# a_11814_9295# 4.3e-19
C6393 a_10864_9269# a_11244_9661# 0.00971f
C6394 a_13142_8359# a_13279_8207# 0.0907f
C6395 net4 net46 0.0382f
C6396 a_3431_10933# a_4687_11231# 0.0436f
C6397 net19 a_9004_3677# 0.00617f
C6398 _022_ a_3947_11305# 5.3e-19
C6399 a_1638_6397# result[0] 7.73e-21
C6400 trim_val\[1\] a_15023_2767# 0.00829f
C6401 a_3224_2601# clk 0.00521f
C6402 a_1844_9129# a_3840_8867# 1.04e-20
C6403 a_13257_4943# VPWR 0.275f
C6404 a_9747_2527# a_10543_2455# 0.00828f
C6405 a_9459_7895# _062_ 6.55e-20
C6406 cal_itt\[1\] a_9460_6807# 0.0366f
C6407 net51 a_5340_6031# 5.9e-20
C6408 _038_ a_11753_6031# 7.31e-19
C6409 _018_ mask\[2\] 4.03e-19
C6410 a_745_10933# a_911_10217# 1.44e-20
C6411 net18 a_11244_9661# 0.00919f
C6412 a_1184_9117# a_1375_9129# 4.61e-19
C6413 net30 a_10245_5193# 8.41e-21
C6414 _009_ a_6541_12021# 0.234f
C6415 a_6375_12021# a_7109_11989# 0.0701f
C6416 net44 _062_ 5.01e-19
C6417 net13 mask\[3\] 0.109f
C6418 net18 a_11204_7485# 9.07e-20
C6419 _048_ a_6316_5193# 0.0991f
C6420 net19 _107_ 0.0393f
C6421 a_1095_12393# a_1000_12381# 0.0498f
C6422 a_4995_7119# _059_ 1.22e-21
C6423 a_2857_5461# _048_ 0.012f
C6424 a_13825_6031# trim_mask\[0\] 1.56e-19
C6425 net12 _003_ 0.181f
C6426 net52 a_3303_7119# 6.98e-19
C6427 a_1201_3855# VPWR 4.86e-19
C6428 a_6743_10933# _020_ 6.39e-20
C6429 _108_ a_11067_4405# 0.03f
C6430 cal_itt\[0\] cal_itt\[3\] 0.00179f
C6431 mask\[0\] a_4043_7093# 0.109f
C6432 a_1019_9839# VPWR 0.134f
C6433 net22 a_561_4405# 0.00108f
C6434 a_2006_8751# VPWR 9.56e-19
C6435 _014_ a_3148_4399# 0.00855f
C6436 mask\[7\] a_1677_9545# 1.54e-19
C6437 net43 a_5915_10927# 4.17e-21
C6438 _120_ _095_ 0.0356f
C6439 net9 cal_count\[2\] 1.69e-20
C6440 net45 a_2033_3317# 0.0342f
C6441 _101_ a_4030_9839# 3.07e-19
C6442 en_co_clk a_4863_4917# 0.00618f
C6443 a_10688_9295# a_11116_8983# 0.00437f
C6444 a_2857_7637# a_4167_6575# 2.04e-21
C6445 a_561_7119# a_1638_7485# 1.46e-19
C6446 a_911_7119# a_816_7119# 0.0498f
C6447 net46 a_14172_4943# 0.286f
C6448 _093_ state\[1\] 3.64e-20
C6449 trim_mask\[0\] a_11067_3017# 6.41e-20
C6450 net18 _123_ 0.00946f
C6451 net19 _049_ 1.21e-20
C6452 _112_ a_14071_3689# 6.26e-19
C6453 mask\[7\] a_1835_11231# 0.0788f
C6454 a_3597_10933# net26 4.29e-20
C6455 _046_ ctlp[1] 0.00205f
C6456 _062_ clk 0.0102f
C6457 net44 a_7367_10927# 0.0154f
C6458 net33 _055_ 0.0246f
C6459 _062_ en_co_clk 0.114f
C6460 VPWR ctlp[0] 0.42f
C6461 net9 a_10688_9295# 7.29e-20
C6462 mask\[2\] mask\[1\] 0.014f
C6463 net19 a_7259_11305# 6.58e-20
C6464 a_1467_7923# _039_ 2.5e-19
C6465 state\[2\] a_5221_1679# 1.41e-19
C6466 net45 a_1549_6794# 0.0027f
C6467 cal_itt\[1\] _107_ 3.8e-19
C6468 a_8381_9295# a_8949_9537# 0.176f
C6469 a_4696_8207# a_4858_8573# 0.00645f
C6470 a_4131_8207# a_4393_8207# 0.00171f
C6471 a_1019_4399# _014_ 7.28e-21
C6472 _074_ a_1019_6397# 0.00467f
C6473 _058_ _112_ 0.0036f
C6474 _074_ _045_ 0.158f
C6475 net15 _102_ 7.88e-20
C6476 _065_ _093_ 0.0062f
C6477 _062_ a_9084_4515# 3.65e-20
C6478 clknet_2_1__leaf_clk _042_ 0.665f
C6479 a_4259_6031# net54 0.00143f
C6480 net43 a_1467_7923# 0.35f
C6481 mask\[4\] net47 0.243f
C6482 a_10975_6031# _066_ 0.0126f
C6483 _064_ a_11321_3855# 2.84e-19
C6484 _053_ a_10990_7485# 0.00917f
C6485 a_7263_7093# VPWR 0.377f
C6486 _099_ a_4471_4007# 9.67e-21
C6487 _092_ trim_mask\[0\] 0.00122f
C6488 cal_count\[3\] _051_ 1.48e-20
C6489 calibrate a_5087_3855# 0.0232f
C6490 a_6210_4989# _089_ 1.88e-19
C6491 clknet_2_3__leaf_clk a_10747_8970# 4.39e-22
C6492 _044_ _020_ 1.01e-19
C6493 _033_ a_9595_1679# 5.24e-22
C6494 net3 _097_ 5.88e-20
C6495 _041_ a_6835_7669# 1.2e-20
C6496 a_15299_3311# trim_val\[1\] 0.1f
C6497 mask\[3\] a_4864_9295# 0.0168f
C6498 net9 a_12410_6031# 4.41e-20
C6499 _011_ a_1137_11721# 0.0157f
C6500 a_579_12021# a_1493_11721# 0.00106f
C6501 net45 a_2491_3311# 0.0138f
C6502 _075_ _092_ 0.0268f
C6503 mask\[6\] a_3133_11247# 0.00286f
C6504 net37 cal_count\[1\] 6.29e-19
C6505 _063_ a_9529_6059# 6.66e-19
C6506 net53 a_7477_10901# 5.65e-19
C6507 _106_ net50 2.39e-21
C6508 calibrate a_1476_4777# 0.0542f
C6509 net44 a_7999_11231# 0.284f
C6510 _039_ _094_ 1.23e-20
C6511 net15 _022_ 0.00821f
C6512 _042_ a_2368_9955# 0.106f
C6513 a_10903_7261# a_11141_6031# 5.81e-21
C6514 cal_itt\[1\] a_8495_6895# 7.48e-20
C6515 clknet_2_1__leaf_clk a_7521_11293# 1.32e-19
C6516 _101_ net25 1.56e-20
C6517 a_9443_6059# a_8298_5487# 0.0067f
C6518 net46 a_11509_3317# 0.0269f
C6519 a_11987_8757# a_12522_8751# 6.02e-19
C6520 _064_ a_11435_2229# 3.82e-21
C6521 net12 a_7223_2465# 1.36e-19
C6522 a_745_10933# a_1000_11293# 0.0642f
C6523 net43 _094_ 2.06e-20
C6524 _107_ a_11067_4405# 0.00192f
C6525 net46 a_14099_3017# 0.00155f
C6526 _065_ _034_ 0.148f
C6527 net44 clknet_2_0__leaf_clk 0.173f
C6528 a_3840_8867# _017_ 3.47e-19
C6529 net43 a_4043_10143# 0.3f
C6530 _074_ _023_ 0.175f
C6531 a_6737_3855# VPWR 0.00397f
C6532 a_6941_2589# VPWR 7.03e-20
C6533 _123_ a_11575_8790# 0.00177f
C6534 a_1493_5487# VPWR 0.252f
C6535 _122_ _133_ 0.11f
C6536 a_13470_7663# en_co_clk 5.5e-22
C6537 net47 _053_ 0.0146f
C6538 a_2971_8457# _017_ 0.117f
C6539 a_4687_12319# a_4687_11231# 9.75e-19
C6540 _071_ a_8307_6575# 0.00405f
C6541 mask\[6\] a_4165_10901# 0.0219f
C6542 a_5524_1679# clk 0.0526f
C6543 en_co_clk a_3817_4697# 5.93e-19
C6544 _082_ a_1497_8725# 5.07e-21
C6545 mask\[6\] a_6541_12021# 3.48e-20
C6546 a_10543_2455# a_10676_1679# 0.00164f
C6547 _126_ _123_ 2.34e-21
C6548 net18 trim_mask\[1\] 0.204f
C6549 a_579_12021# VPWR 0.459f
C6550 _119_ _026_ 2.56e-20
C6551 net33 trim_val\[2\] 0.00704f
C6552 a_9595_1679# a_10785_1679# 2.56e-19
C6553 net30 a_8473_5193# 6.47e-19
C6554 clknet_2_3__leaf_clk a_11369_7119# 2.64e-19
C6555 net51 a_6631_7485# 3.67e-19
C6556 a_579_12021# a_1769_12393# 2.56e-19
C6557 net53 _019_ 0.00889f
C6558 _015_ a_2143_2229# 9.18e-22
C6559 a_1476_10217# result[4] 2.85e-19
C6560 clknet_2_2__leaf_clk a_7715_3285# 4.38e-20
C6561 net50 _033_ 2.07e-20
C6562 net37 _108_ 1.02e-19
C6563 _118_ a_9664_3689# 8.28e-20
C6564 net13 a_4687_11231# 0.0175f
C6565 _074_ a_816_10205# 0.00248f
C6566 trim_mask\[0\] a_9317_3285# 1.49e-20
C6567 clknet_2_0__leaf_clk clk 0.0705f
C6568 _074_ _013_ 1.14e-20
C6569 net44 net13 0.217f
C6570 clknet_2_1__leaf_clk a_6909_10933# 0.0064f
C6571 clknet_2_0__leaf_clk en_co_clk 0.0128f
C6572 _062_ _059_ 0.102f
C6573 _007_ result[4] 7.64e-20
C6574 net23 a_448_7637# 0.181f
C6575 _053_ a_8820_6005# 0.0384f
C6576 net40 VPWR 2.22f
C6577 _078_ a_2961_9295# 1.2e-20
C6578 net45 a_2143_7663# 0.0631f
C6579 a_1467_7923# a_2857_7637# 1.43e-20
C6580 a_2869_10927# VPWR 0.181f
C6581 _048_ a_6210_4989# 0.111f
C6582 net43 a_2787_7119# 0.298f
C6583 _132_ a_15259_7637# 0.00127f
C6584 a_13059_4631# _110_ 0.17f
C6585 net14 _086_ 0.0147f
C6586 a_13607_4943# _112_ 1.87e-20
C6587 net42 _103_ 0.127f
C6588 a_12231_6005# a_12323_4703# 1.03e-20
C6589 _122_ a_14236_8457# 1.55e-19
C6590 _123_ a_12153_8757# 0.017f
C6591 net18 a_8749_3317# 8.89e-21
C6592 net41 a_3123_3615# 0.0673f
C6593 _102_ net25 2.7e-20
C6594 _002_ a_6835_7669# 0.284f
C6595 cal_itt\[0\] a_9602_6941# 2.23e-19
C6596 _015_ a_4815_3031# 5.91e-19
C6597 net4 a_7527_4631# 2.66e-21
C6598 _000_ _072_ 6.76e-22
C6599 _058_ a_12121_3677# 2.61e-19
C6600 net22 result[0] 0.00496f
C6601 trim_mask\[4\] a_11057_4105# 0.00264f
C6602 _065_ a_3830_6281# 2.58e-19
C6603 a_1137_5487# sample 3.96e-19
C6604 a_13257_1141# a_13607_1513# 0.23f
C6605 a_13091_1141# a_14347_1439# 0.0436f
C6606 net53 a_6467_9845# 0.0225f
C6607 net14 _102_ 1.21e-20
C6608 a_11343_3317# a_11509_3317# 0.578f
C6609 net26 a_6888_10205# 0.0163f
C6610 net9 a_12612_8725# 0.0048f
C6611 a_929_8757# a_1184_9117# 0.0594f
C6612 clknet_2_1__leaf_clk a_3597_12021# 0.597f
C6613 a_745_12021# a_1095_12393# 0.23f
C6614 a_13459_3317# a_13881_2741# 0.00145f
C6615 net18 a_10977_2543# 3.1e-19
C6616 net4 state\[1\] 0.483f
C6617 net13 clk 0.015f
C6618 net30 a_8583_3317# 6.14e-21
C6619 a_11244_9661# a_11268_9295# 0.0016f
C6620 _000_ _068_ 0.101f
C6621 net13 en_co_clk 0.0537f
C6622 _127_ a_14733_9545# 0.00787f
C6623 a_13557_8457# a_13279_8207# 3.25e-19
C6624 net12 net26 0.102f
C6625 net9 _108_ 0.0117f
C6626 a_13519_4007# net49 3.31e-19
C6627 a_11583_4777# _058_ 0.0112f
C6628 a_12148_4777# a_13059_4631# 3.19e-19
C6629 net46 a_9007_2601# 0.152f
C6630 _095_ a_1867_3317# 1.61e-19
C6631 net53 VPWR 0.629f
C6632 net43 a_3208_10205# 0.0251f
C6633 a_13356_7369# _134_ 6.3e-20
C6634 net12 _088_ 3.71e-19
C6635 a_2857_7637# _094_ 2.84e-21
C6636 _046_ a_3947_11305# 1.31e-19
C6637 a_2787_9845# _040_ 1.17e-21
C6638 net50 a_10785_1679# 1.51e-19
C6639 clknet_2_1__leaf_clk a_1137_11721# 4.44e-19
C6640 _065_ net4 0.0126f
C6641 net53 a_5699_9269# 3.23e-20
C6642 trim_mask\[0\] a_6737_4719# 2.27e-21
C6643 net19 trim_mask\[4\] 0.00699f
C6644 _017_ a_4131_8207# 5.03e-19
C6645 net44 a_4864_9295# 7.6e-19
C6646 net45 a_1007_6031# 9.54e-19
C6647 a_13881_1653# a_13257_1141# 4.54e-19
C6648 _041_ a_13184_9117# 0.00127f
C6649 _051_ _119_ 4.4e-20
C6650 mask\[2\] _041_ 0.284f
C6651 net2 a_13557_7369# 2.43e-20
C6652 a_579_12021# net27 0.00152f
C6653 a_1651_10143# a_763_8757# 1.17e-19
C6654 net26 a_6983_10217# 0.0301f
C6655 a_12723_4943# a_13091_4943# 5.61e-20
C6656 a_3116_12533# mask\[6\] 5.65e-21
C6657 a_395_4405# _012_ 0.17f
C6658 _122_ _129_ 0.00432f
C6659 a_6173_7119# a_6515_6794# 5.35e-19
C6660 _092_ a_8307_4943# 8.22e-20
C6661 _059_ a_3817_4697# 7.37e-21
C6662 net12 a_6519_4631# 0.00775f
C6663 net49 a_14604_3017# 0.00295f
C6664 _075_ a_5547_5603# 0.159f
C6665 a_5515_6005# _050_ 0.00416f
C6666 trim_mask\[0\] a_9003_3829# 0.0296f
C6667 a_13470_7663# cal_count\[2\] 0.132f
C6668 _093_ _013_ 0.0321f
C6669 net46 net48 9.52e-19
C6670 net43 a_7088_7119# 1.11e-19
C6671 cal_itt\[0\] _035_ 0.0171f
C6672 a_2092_8457# _040_ 0.106f
C6673 mask\[1\] a_2174_8457# 2.2e-19
C6674 _121_ a_4091_5309# 7.67e-21
C6675 _051_ a_6566_5193# 1.67e-19
C6676 net33 trim_mask\[0\] 0.0121f
C6677 a_2857_7637# a_2787_7119# 0.0219f
C6678 _024_ VPWR 0.523f
C6679 clknet_2_0__leaf_clk _059_ 2.05e-19
C6680 net26 a_1651_10143# 6.96e-20
C6681 _095_ _051_ 6.97e-20
C6682 mask\[4\] _068_ 3.07e-20
C6683 net43 _063_ 0.00244f
C6684 net40 a_14807_8359# 0.00443f
C6685 net16 _111_ 7.22e-22
C6686 net4 a_9761_8457# 4.24e-19
C6687 cal_count\[0\] _037_ 2.17e-20
C6688 clknet_2_3__leaf_clk a_10005_6031# 0.00105f
C6689 a_9802_4007# a_10188_4105# 0.0158f
C6690 a_15023_12559# VPWR 0.407f
C6691 net23 a_911_7119# 6.34e-19
C6692 a_10111_1679# a_10016_1679# 0.0498f
C6693 a_10975_6031# a_12056_6031# 0.102f
C6694 _075_ a_5536_4399# 0.00358f
C6695 a_10329_1921# a_10219_2045# 0.0977f
C6696 _038_ a_12231_6005# 1.39e-19
C6697 net37 a_12900_7663# 9.31e-37
C6698 _074_ _078_ 0.166f
C6699 a_13257_1141# a_14334_1135# 1.46e-19
C6700 a_13825_1109# a_13715_1135# 0.0977f
C6701 a_14564_6397# net35 0.025f
C6702 a_448_10357# _007_ 0.00126f
C6703 a_13257_4943# _110_ 0.00146f
C6704 calibrate a_6822_4105# 0.00142f
C6705 _095_ _014_ 0.123f
C6706 a_13625_3317# a_13975_3689# 0.23f
C6707 mask\[4\] a_4443_9295# 5.48e-19
C6708 a_12612_8725# a_12436_9129# 0.26f
C6709 a_12153_8757# a_13142_8725# 0.0728f
C6710 net9 a_12516_2601# 0.0115f
C6711 _015_ a_4443_1679# 0.17f
C6712 _108_ a_10188_4105# 0.0216f
C6713 a_11023_5108# trim_mask\[1\] 8.85e-19
C6714 a_3399_2527# a_3224_2601# 0.234f
C6715 a_3521_9813# a_3303_10217# 0.21f
C6716 a_2953_9845# a_4043_10143# 0.0424f
C6717 net30 a_7190_3855# 2.4e-19
C6718 _113_ _112_ 0.11f
C6719 _106_ _033_ 6.82e-20
C6720 _067_ a_10043_7983# 6.92e-19
C6721 _092_ a_7210_5807# 0.00778f
C6722 net46 a_13091_1141# 0.502f
C6723 _085_ _010_ 0.19f
C6724 _104_ a_6737_3855# 0.03f
C6725 clknet_2_3__leaf_clk a_8839_9661# 8.49e-19
C6726 _076_ a_4259_6031# 8.74e-20
C6727 net13 a_4801_9839# 0.00833f
C6728 net27 net53 1.42e-19
C6729 a_14983_9269# a_15111_9295# 0.00476f
C6730 net34 _055_ 0.161f
C6731 _130_ net5 2.21e-19
C6732 _078_ a_1279_9129# 0.00886f
C6733 a_2689_8751# a_2857_7637# 1.49e-19
C6734 net13 _059_ 0.00434f
C6735 _040_ net51 0.00283f
C6736 _123_ a_13050_7637# 0.0391f
C6737 net46 _064_ 0.0173f
C6738 net35 a_13091_4943# 7.94e-19
C6739 a_13091_4943# a_13059_4631# 0.00126f
C6740 _119_ a_10781_3311# 1.08e-19
C6741 trim_mask\[2\] a_12599_3615# 6.44e-20
C6742 net15 _046_ 0.135f
C6743 trim_mask\[2\] a_11413_2767# 0.00175f
C6744 net44 a_4239_8573# 0.0122f
C6745 net30 a_911_4777# 4.91e-21
C6746 net31 net2 0.00231f
C6747 _016_ a_3303_7119# 0.00139f
C6748 _133_ comp 5.22e-20
C6749 a_4995_7119# _049_ 0.0028f
C6750 net9 a_12900_7663# 0.00332f
C6751 _011_ net43 6.44e-19
C6752 a_14540_3689# a_14702_3311# 0.00645f
C6753 a_11067_4405# trim_mask\[4\] 0.00152f
C6754 _024_ a_9478_4105# 6.23e-22
C6755 _065_ a_10586_7371# 0.00918f
C6756 cal_itt\[3\] a_7723_6807# 0.14f
C6757 _068_ _053_ 0.00191f
C6758 _118_ a_10245_5193# 5.24e-19
C6759 net19 a_9195_10357# 0.00502f
C6760 _027_ a_7942_2223# 9.25e-21
C6761 a_7223_2465# a_7524_2223# 9.73e-19
C6762 a_6467_9845# a_6007_9839# 3e-20
C6763 _008_ a_5829_9839# 0.0125f
C6764 _071_ VPWR 0.473f
C6765 a_14347_9480# _125_ 0.023f
C6766 a_8949_6031# _107_ 1.42e-19
C6767 _127_ a_15159_9269# 6.21e-19
C6768 _074_ a_3597_10933# 9.03e-20
C6769 cal_itt\[2\] a_7001_7669# 0.00182f
C6770 net46 a_10851_1653# 0.367f
C6771 net16 a_13257_1141# 3.08e-20
C6772 net4 _067_ 0.0556f
C6773 _128_ a_14249_8725# 3.86e-19
C6774 _062_ _108_ 0.0054f
C6775 a_3431_12021# a_4055_12015# 9.73e-19
C6776 clknet_2_1__leaf_clk mask\[5\] 0.0811f
C6777 a_4165_11989# a_4621_12393# 4.2e-19
C6778 a_3947_12393# a_4209_12381# 0.00171f
C6779 a_13703_1513# VPWR 0.00447f
C6780 en_co_clk a_4091_4943# 1.02e-19
C6781 net43 a_4209_11293# 0.00237f
C6782 a_9317_3285# a_8298_2767# 0.00792f
C6783 mask\[0\] a_3748_6281# 3.54e-19
C6784 a_14564_6397# _061_ 0.16f
C6785 net44 a_7631_12319# 0.287f
C6786 _132_ a_14485_7663# 0.00372f
C6787 a_7109_11989# a_7456_12393# 0.0512f
C6788 net3 a_4709_2773# 4.79e-20
C6789 a_6007_9839# VPWR 0.178f
C6790 a_10655_2932# trim_mask\[3\] 6.83e-19
C6791 calibrate a_1867_3317# 2.84e-20
C6792 net1 a_455_3571# 0.189f
C6793 cal_count\[1\] a_13470_7663# 0.00724f
C6794 _053_ net46 6.57e-19
C6795 ctln[3] ctln[2] 0.00303f
C6796 _078_ _093_ 4.53e-21
C6797 a_11859_3689# a_11764_3677# 0.0498f
C6798 a_12077_3285# a_11955_3689# 3.16e-19
C6799 trim_mask\[1\] a_12691_2527# 1.09e-19
C6800 a_10239_9295# a_10864_9269# 0.185f
C6801 net3 a_4308_4917# 0.0394f
C6802 _035_ a_10405_9295# 0.173f
C6803 net45 a_6173_7119# 4.54e-22
C6804 a_2787_10927# a_3431_10933# 0.00122f
C6805 a_6007_9839# a_5699_9269# 1.4e-19
C6806 a_4609_9295# mask\[1\] 2e-21
C6807 _029_ VPWR 0.411f
C6808 a_8491_2229# a_9572_2601# 0.102f
C6809 _027_ a_9747_2527# 0.0413f
C6810 net18 a_10239_9295# 0.016f
C6811 a_2953_9845# a_3208_10205# 0.0604f
C6812 _107_ a_10188_4105# 2.75e-20
C6813 net4 clknet_2_2__leaf_clk 0.744f
C6814 _009_ _042_ 5.83e-21
C6815 net52 a_2815_9447# 0.177f
C6816 net44 a_9020_10383# 5.49e-20
C6817 net17 _041_ 1.18e-20
C6818 net19 ctlp[5] 0.00847f
C6819 net44 a_4167_6575# 3.92e-21
C6820 a_11233_4405# a_11509_3317# 4e-20
C6821 net46 a_14281_1513# 6.14e-19
C6822 a_9460_6807# _062_ 0.109f
C6823 net33 a_14983_9269# 0.00314f
C6824 _136_ trim_mask\[0\] 0.00162f
C6825 _064_ a_11343_3317# 3.82e-21
C6826 mask\[2\] a_3615_8207# 0.00131f
C6827 a_11244_9661# VPWR 0.433f
C6828 a_4425_6031# net30 7.21e-20
C6829 _064_ a_11149_3017# 0.0106f
C6830 net20 a_7153_12381# 4.97e-19
C6831 a_1541_9117# VPWR 2.95e-19
C6832 net34 trim_val\[2\] 0.0981f
C6833 a_1313_10901# net52 2.03e-19
C6834 a_1095_11305# a_1660_11305# 7.99e-20
C6835 a_7459_7663# a_7263_7093# 8.82e-19
C6836 net19 a_8949_9537# 0.00894f
C6837 _133_ a_13111_6031# 4.7e-21
C6838 a_2948_3689# clk 5.5e-19
C6839 a_11204_7485# VPWR 0.143f
C6840 _101_ _019_ 0.0725f
C6841 trim_mask\[2\] a_10543_2455# 9.79e-20
C6842 trim_mask\[3\] a_12516_2601# 1.06e-19
C6843 a_11801_4373# a_11679_4777# 3.16e-19
C6844 a_11583_4777# a_11488_4765# 0.0498f
C6845 _130_ a_15023_6031# 5.13e-22
C6846 a_1660_12393# a_579_10933# 6.19e-20
C6847 a_10699_3311# a_10676_1679# 4.52e-21
C6848 mask\[3\] a_4043_10143# 5.87e-20
C6849 _051_ calibrate 0.00542f
C6850 net15 a_3053_8207# 5.78e-20
C6851 _060_ a_5363_4719# 0.00436f
C6852 a_10245_5193# a_10137_4943# 5.37e-19
C6853 a_13091_4943# a_13257_4943# 0.685f
C6854 clknet_2_2__leaf_clk a_14172_4943# 2.43e-21
C6855 a_4621_12393# VPWR 3.99e-20
C6856 a_15023_2767# a_15023_1679# 8.27e-21
C6857 net33 _030_ 1.44e-20
C6858 a_12169_2197# a_12047_2601# 3.16e-19
C6859 a_11951_2601# a_11856_2589# 0.0498f
C6860 net45 a_3333_2601# 6.92e-19
C6861 calibrate _014_ 0.00963f
C6862 a_13349_6031# VPWR 0.00701f
C6863 _050_ a_4815_3031# 3.11e-19
C6864 _123_ VPWR 3.25f
C6865 net52 _081_ 1.28e-19
C6866 _091_ a_10055_5487# 3.02e-20
C6867 _129_ comp 0.00337f
C6868 _062_ _107_ 0.0161f
C6869 net34 a_15259_7637# 0.00866f
C6870 _024_ _104_ 0.00874f
C6871 net40 _110_ 1.8e-20
C6872 _074_ _004_ 0.136f
C6873 _136_ a_13933_6281# 0.00188f
C6874 a_9003_3829# a_8298_2767# 0.00226f
C6875 _125_ a_14870_7369# 2.38e-20
C6876 clknet_2_0__leaf_clk a_3399_2527# 0.0495f
C6877 a_5363_7369# VPWR 0.404f
C6878 net46 a_14335_4020# 2.15e-19
C6879 a_745_12021# a_1461_10357# 2.75e-22
C6880 a_3868_7119# net30 1.04e-20
C6881 net44 a_8731_9295# 5.09e-19
C6882 _101_ a_6467_9845# 6.71e-21
C6883 _049_ a_4863_4917# 0.00169f
C6884 _000_ _065_ 6.57e-20
C6885 _067_ a_10586_7371# 0.0051f
C6886 a_561_9845# a_1129_9813# 0.181f
C6887 clknet_2_1__leaf_clk net43 0.305f
C6888 a_9004_3677# a_9195_3689# 4.61e-19
C6889 a_14193_3285# a_14083_3311# 0.0977f
C6890 a_13625_3317# trim_val\[1\] 6.71e-19
C6891 cal_count\[2\] a_14788_7369# 0.101f
C6892 _028_ clk 0.0679f
C6893 _012_ a_2283_4020# 1.22e-19
C6894 _010_ a_2828_12131# 2.42e-19
C6895 mask\[6\] a_1357_11293# 1.94e-21
C6896 _062_ _049_ 0.0151f
C6897 a_12516_2601# a_13415_2442# 0.00253f
C6898 a_5997_10927# net26 5.73e-20
C6899 _133_ a_11622_7485# 8.76e-21
C6900 _086_ a_1493_11721# 0.0985f
C6901 _101_ VPWR 1.68f
C6902 _115_ _114_ 0.142f
C6903 net12 net55 0.00863f
C6904 _107_ a_9195_3689# 2.69e-19
C6905 a_6541_12021# _021_ 1.23e-20
C6906 net44 a_5915_10927# 9.27e-20
C6907 net40 a_10699_5487# 1.71e-19
C6908 net18 _066_ 0.0344f
C6909 _122_ _038_ 0.00538f
C6910 _125_ a_13562_8751# 1.71e-20
C6911 _050_ a_7843_3677# 0.00186f
C6912 calibrate a_5445_4399# 8.7e-21
C6913 _101_ a_5699_9269# 1.38e-19
C6914 _051_ a_8298_5487# 0.00607f
C6915 en_co_clk a_3461_5193# 0.00424f
C6916 a_9043_6031# VPWR 1.45e-19
C6917 _062_ a_8495_6895# 7.64e-19
C6918 clknet_2_2__leaf_clk a_11509_3317# 0.596f
C6919 a_4131_8207# _121_ 5.22e-20
C6920 _074_ net12 4.02e-19
C6921 net43 a_2368_9955# 0.0294f
C6922 a_4055_12015# a_4167_11471# 8.84e-19
C6923 _078_ _083_ 0.147f
C6924 trim_mask\[2\] a_13607_1513# 2.23e-19
C6925 _092_ a_9529_6059# 0.00232f
C6926 _090_ net3 0.0948f
C6927 _037_ en_co_clk 3.09e-20
C6928 clknet_2_0__leaf_clk a_4725_5487# 1.15e-20
C6929 mask\[2\] a_3249_9295# 8.74e-19
C6930 clknet_2_3__leaf_clk a_12341_8751# 6.75e-19
C6931 cal_count\[0\] _122_ 0.0604f
C6932 clknet_2_0__leaf_clk en 6.3e-20
C6933 a_8307_4943# a_8485_4943# 0.00762f
C6934 a_7569_7637# _073_ 2.27e-20
C6935 a_3947_12393# a_3431_10933# 3.71e-21
C6936 _052_ a_7843_3677# 0.00101f
C6937 mask\[3\] a_3208_10205# 1.66e-20
C6938 trim_mask\[0\] _105_ 0.00879f
C6939 net3 a_3847_4438# 2.81e-19
C6940 _088_ _089_ 5.01e-19
C6941 a_13142_8359# a_13142_7271# 8.87e-19
C6942 mask\[6\] _042_ 1.95e-19
C6943 net9 trim_mask\[4\] 2.61e-20
C6944 a_10543_2455# a_9595_1679# 2.31e-19
C6945 a_9572_2601# _032_ 0.00731f
C6946 _001_ a_11895_7669# 1.09e-19
C6947 net29 net26 2.24e-20
C6948 a_7999_11231# a_8178_11293# 0.0074f
C6949 a_7259_11305# a_7367_10927# 0.0572f
C6950 a_7824_11305# a_7933_11305# 0.00742f
C6951 a_7477_10901# a_7986_10927# 2.6e-19
C6952 a_9296_9295# cal_itt\[0\] 0.00177f
C6953 net30 _103_ 0.102f
C6954 _050_ a_5087_3855# 5.91e-21
C6955 _086_ VPWR 0.158f
C6956 net5 trim[4] 2.79e-19
C6957 net18 a_11545_9049# 4.43e-19
C6958 net36 net37 0.00645f
C6959 _118_ a_8583_3317# 1.22e-19
C6960 a_3425_11721# a_3431_10933# 1.15e-19
C6961 _034_ a_5502_6397# 1.66e-20
C6962 net44 a_8072_11721# 0.00258f
C6963 trim_mask\[1\] VPWR 1.98f
C6964 a_6785_7119# VPWR 6.92e-20
C6965 a_9459_7895# a_9621_8029# 0.00401f
C6966 net21 a_4055_12015# 2.12e-19
C6967 a_1129_7361# net22 1.74e-19
C6968 a_13142_8725# VPWR 0.248f
C6969 net8 ctln[3] 2.28e-19
C6970 _123_ a_14807_8359# 2.1e-21
C6971 _102_ VPWR 0.508f
C6972 a_6703_2197# VPWR 0.391f
C6973 trim_mask\[2\] a_13881_1653# 0.111f
C6974 _040_ a_5050_8207# 6.31e-19
C6975 net50 a_11057_3855# 2.29e-19
C6976 _024_ _110_ 1.51e-21
C6977 net13 a_4725_5487# 1.33e-19
C6978 _052_ a_5087_3855# 2.83e-37
C6979 clknet_2_2__leaf_clk a_7689_2589# 2.44e-19
C6980 a_12900_7663# a_13470_7663# 0.111f
C6981 _001_ a_11491_6031# 2.66e-19
C6982 a_745_12021# a_745_10933# 6.68e-19
C6983 net40 a_14564_6397# 0.0142f
C6984 _053_ a_7527_4631# 6.7e-20
C6985 _049_ a_3817_4697# 8.24e-19
C6986 a_8083_8181# _070_ 0.0951f
C6987 clknet_2_3__leaf_clk a_10864_7387# 0.161f
C6988 _015_ a_1867_3317# 3.05e-21
C6989 net45 a_5037_6031# 5.61e-21
C6990 a_4609_9295# _041_ 1.44e-20
C6991 clknet_2_1__leaf_clk a_2857_7637# 1.63f
C6992 a_4443_1679# a_5055_1679# 0.00188f
C6993 a_4609_1679# a_5686_2045# 1.46e-19
C6994 a_4959_1679# a_4864_1679# 0.0498f
C6995 a_5177_1921# a_5067_2045# 0.0977f
C6996 a_11435_2229# _057_ 1.44e-20
C6997 a_5699_1653# a_5524_1679# 0.234f
C6998 net44 _094_ 0.14f
C6999 cal_itt\[0\] cal_count\[3\] 8.11e-20
C7000 a_6173_7119# a_8022_7119# 2.77e-19
C7001 net27 _101_ 1.61e-19
C7002 _074_ a_1651_10143# 0.0107f
C7003 _133_ a_14199_7369# 1.4e-21
C7004 a_6741_7361# a_7088_7119# 0.0512f
C7005 _053_ state\[1\] 0.0276f
C7006 _078_ a_911_7119# 0.00147f
C7007 _042_ _035_ 2.32e-20
C7008 a_7477_10901# a_7824_11305# 0.0512f
C7009 _043_ a_7548_10217# 2.32e-20
C7010 net41 a_6737_3855# 4.1e-20
C7011 a_8749_3317# VPWR 0.591f
C7012 cal_count\[1\] a_14788_7369# 4.41e-21
C7013 a_15259_7637# a_15299_6575# 4.01e-20
C7014 net18 _043_ 0.0211f
C7015 a_10239_9295# a_11268_9295# 0.00248f
C7016 _060_ VPWR 0.535f
C7017 net46 a_15299_3311# 5.03e-19
C7018 _096_ a_4617_4105# 0.016f
C7019 net40 a_14467_8751# 0.0103f
C7020 clknet_2_0__leaf_clk _049_ 0.221f
C7021 a_8386_8457# a_8301_8207# 8.13e-19
C7022 a_561_6031# a_1476_4777# 5.53e-21
C7023 a_1476_6031# a_561_4405# 5.53e-21
C7024 a_11067_4405# a_13059_4631# 5.67e-21
C7025 _024_ a_12148_4777# 0.00102f
C7026 clknet_2_0__leaf_clk a_3388_4631# 4.11e-20
C7027 net16 a_14282_7119# 4.83e-19
C7028 _125_ _131_ 3e-21
C7029 _022_ VPWR 0.439f
C7030 net43 a_1953_9129# 2.95e-19
C7031 net40 a_13091_4943# 0.0196f
C7032 _065_ _053_ 0.352f
C7033 net50 a_10543_2455# 0.0102f
C7034 net13 _107_ 5.96e-20
C7035 clknet_2_2__leaf_clk a_9007_2601# 0.0413f
C7036 net2 a_14733_7983# 5.79e-19
C7037 a_10977_2543# VPWR 6e-20
C7038 a_6375_12021# VPWR 0.43f
C7039 net54 a_4709_2773# 3.91e-19
C7040 _121_ net30 0.0346f
C7041 a_1651_10143# a_1279_9129# 9.43e-19
C7042 a_10188_4105# trim_mask\[4\] 0.135f
C7043 net45 _005_ 8.46e-20
C7044 a_11016_6691# a_11098_6691# 0.00477f
C7045 a_8495_6895# a_8745_6895# 0.089f
C7046 a_14565_9295# VPWR 8.6e-19
C7047 a_395_4405# a_1651_4703# 0.0435f
C7048 _012_ a_911_4777# 0.00484f
C7049 a_12992_8751# _133_ 7.58e-21
C7050 _094_ en_co_clk 0.112f
C7051 a_4993_6273# a_4883_6397# 0.0977f
C7052 a_4775_6031# a_4680_6031# 0.0498f
C7053 a_1129_9813# _006_ 2.15e-19
C7054 _048_ _088_ 0.283f
C7055 mask\[6\] a_6909_10933# 6.26e-20
C7056 a_4308_4917# net54 0.142f
C7057 net46 a_9664_3689# 0.223f
C7058 net43 a_4866_12381# 0.00196f
C7059 net47 _124_ 0.0145f
C7060 a_7262_5461# _048_ 0.0893f
C7061 net27 _086_ 0.193f
C7062 a_7939_10383# clknet_2_3__leaf_clk 1.16e-20
C7063 net44 a_2787_7119# 3.16e-20
C7064 net15 net45 1.2f
C7065 net13 _049_ 0.127f
C7066 _051_ _015_ 0.0399f
C7067 net33 a_15083_4659# 0.00242f
C7068 clknet_0_clk _071_ 0.0306f
C7069 _112_ a_13881_2741# 0.115f
C7070 a_448_7637# _004_ 9.22e-20
C7071 net13 a_5699_1653# 0.00214f
C7072 _120_ _050_ 0.0965f
C7073 _066_ a_11023_5108# 1.04e-19
C7074 net46 a_10689_2223# 0.00236f
C7075 _037_ cal_count\[2\] 2.99e-19
C7076 a_9361_3677# VPWR 2.92e-19
C7077 _074_ result[2] 0.00705f
C7078 clknet_2_1__leaf_clk a_2953_9845# 0.131f
C7079 net9 _128_ 0.00665f
C7080 a_7986_10927# VPWR 7.73e-19
C7081 _115_ VPWR 0.452f
C7082 mask\[4\] a_4696_8207# 8.26e-21
C7083 a_9296_9295# a_10405_9295# 9.13e-19
C7084 net43 a_6007_7119# 1.21e-19
C7085 clknet_2_2__leaf_clk net48 2.26e-20
C7086 a_6927_12559# a_6999_12015# 2.85e-19
C7087 a_9478_4105# a_8749_3317# 7.53e-21
C7088 a_8992_9955# a_8731_9295# 0.00374f
C7089 _048_ a_6519_4631# 0.124f
C7090 net46 a_11425_5487# 1.51e-19
C7091 trim_mask\[4\] trim_mask\[3\] 0.352f
C7092 net18 a_9471_9269# 6.47e-19
C7093 a_6515_8534# VPWR 7.28e-19
C7094 a_2092_8457# a_2143_7663# 7.94e-19
C7095 _103_ state\[2\] 0.00629f
C7096 a_4165_11989# a_4512_12393# 0.0512f
C7097 net2 a_11059_7356# 3.56e-20
C7098 a_3597_12021# mask\[6\] 1.19e-20
C7099 net34 a_14983_9269# 0.0122f
C7100 net28 net26 1.3e-20
C7101 a_8301_8207# a_8091_7967# 3e-19
C7102 mask\[2\] a_2019_9055# 1.21e-20
C7103 a_5515_6005# _099_ 1.09e-21
C7104 net16 trim_mask\[2\] 0.0178f
C7105 _062_ trim_mask\[4\] 1.19e-20
C7106 a_14347_1439# _057_ 1.12e-19
C7107 _029_ _110_ 1.78e-19
C7108 net46 trim[4] 5.7e-19
C7109 _045_ net20 0.014f
C7110 a_12424_3689# a_13625_3317# 6.92e-20
C7111 _067_ _064_ 0.0254f
C7112 a_11545_9049# a_12153_8757# 1.07e-19
C7113 a_6743_10933# a_7548_10217# 2.8e-21
C7114 cal_itt\[0\] a_9463_8725# 0.00255f
C7115 cal_count\[3\] trim_mask\[0\] 2.78e-19
C7116 a_7939_3855# VPWR 0.344f
C7117 net46 a_10781_3631# 1.94e-21
C7118 _009_ mask\[5\] 1.37e-19
C7119 a_2368_9955# a_2953_9845# 4.27e-20
C7120 net14 a_1638_4399# 1.25e-19
C7121 a_7569_7637# a_8078_7663# 2.6e-19
C7122 _034_ a_5340_6031# 1.97e-19
C7123 a_14335_7895# VPWR 0.376f
C7124 _081_ net23 0.0986f
C7125 net46 a_14184_1679# 1.37e-19
C7126 _074_ a_1191_11305# 0.00132f
C7127 clknet_2_3__leaf_clk _111_ 2.64e-20
C7128 net43 _092_ 2.25e-20
C7129 a_4498_4373# VPWR 0.367f
C7130 _129_ a_14199_7369# 0.0763f
C7131 a_4864_1679# VPWR 0.0829f
C7132 a_395_6031# a_816_6031# 0.0931f
C7133 _105_ a_8307_4943# 0.165f
C7134 a_6375_12021# net27 2.6e-19
C7135 clknet_2_2__leaf_clk a_13091_1141# 0.254f
C7136 a_7824_11305# VPWR 0.303f
C7137 a_937_3855# cal 1.54e-19
C7138 net9 a_12723_4943# 0.00327f
C7139 a_4471_4007# a_4709_2773# 6.94e-21
C7140 a_9664_3689# a_11343_3317# 3.63e-20
C7141 a_9839_3615# _025_ 6.6e-21
C7142 trim_mask\[2\] a_10699_3311# 0.0648f
C7143 trim_mask\[4\] a_9195_3689# 0.00435f
C7144 en_co_clk a_4617_3855# 7.94e-20
C7145 a_3123_3615# a_3224_2601# 3.54e-22
C7146 a_8935_6895# VPWR 0.00379f
C7147 _064_ clknet_2_2__leaf_clk 0.246f
C7148 a_6793_8970# a_6885_8372# 1.62e-19
C7149 _076_ a_6056_8359# 0.342f
C7150 net43 result[4] 7.88e-19
C7151 net9 a_11895_7669# 0.019f
C7152 _133_ a_14422_7093# 3.3e-19
C7153 net44 a_7088_7119# 0.249f
C7154 _018_ _082_ 9.07e-20
C7155 _104_ trim_mask\[1\] 0.212f
C7156 a_9459_7895# _063_ 0.0778f
C7157 _067_ _053_ 0.0272f
C7158 net37 net35 0.0143f
C7159 _094_ _059_ 0.0451f
C7160 a_12056_6031# a_12165_6031# 0.00742f
C7161 cal_count\[3\] a_13933_6281# 6.02e-20
C7162 a_3868_10217# a_4030_9839# 0.00645f
C7163 _083_ a_6888_10205# 4.21e-20
C7164 a_12231_6005# a_12410_6031# 0.0074f
C7165 net18 _058_ 0.0388f
C7166 _088_ a_7021_4105# 0.0463f
C7167 a_12992_8751# _129_ 6.61e-20
C7168 a_1660_12393# result[6] 1.96e-19
C7169 a_11204_7485# a_10699_5487# 9.19e-21
C7170 net44 _063_ 1.71e-20
C7171 net15 a_2953_7119# 0.0179f
C7172 net4 a_7001_7669# 6.04e-21
C7173 a_4512_12393# VPWR 0.31f
C7174 net12 _083_ 0.00879f
C7175 net43 cal_itt\[3\] 1.33e-20
C7176 a_4165_11989# _046_ 0.00279f
C7177 clknet_2_2__leaf_clk a_10851_1653# 4.35e-20
C7178 net27 a_7986_10927# 1.8e-20
C7179 mask\[1\] a_5535_8181# 0.00518f
C7180 a_9003_3829# a_9369_4105# 0.12f
C7181 net16 net39 0.0166f
C7182 _065_ a_3891_4943# 0.00195f
C7183 a_7460_5807# a_7571_4943# 8.25e-21
C7184 net9 a_11491_6031# 1.97e-19
C7185 _132_ _133_ 0.00744f
C7186 _078_ a_4055_10927# 2.26e-19
C7187 net52 a_3781_8207# 0.00316f
C7188 _090_ net54 0.259f
C7189 _103_ _100_ 3.7e-20
C7190 a_1476_6031# result[0] 3.43e-19
C7191 _033_ a_8912_2589# 6.61e-19
C7192 _122_ en_co_clk 0.465f
C7193 a_4425_6031# a_4775_6031# 0.23f
C7194 a_4259_6031# a_5515_6005# 0.0435f
C7195 net33 _133_ 5.06e-20
C7196 _104_ a_8749_3317# 0.287f
C7197 a_10699_3311# a_11045_3631# 0.0134f
C7198 a_7088_7119# clk 0.00192f
C7199 net21 net26 2.96e-20
C7200 net12 net4 0.00967f
C7201 net14 net45 0.0278f
C7202 net22 calibrate 1.75e-20
C7203 net9 a_11967_3311# 0.00125f
C7204 _052_ a_6822_4105# 0.00165f
C7205 a_14249_8725# net40 0.00278f
C7206 a_14236_8457# a_14422_7093# 6.12e-19
C7207 _053_ clknet_2_2__leaf_clk 0.00227f
C7208 _083_ a_6983_10217# 5.28e-20
C7209 _101_ clknet_0_clk 0.00175f
C7210 a_14972_5193# _047_ 0.11f
C7211 _051_ a_7184_2339# 0.00143f
C7212 _063_ clk 7.88e-20
C7213 net15 a_3399_10217# 1.49e-19
C7214 _063_ en_co_clk 0.0175f
C7215 cal_itt\[2\] _048_ 2.04e-20
C7216 clknet_2_1__leaf_clk mask\[3\] 0.737f
C7217 net46 _057_ 1.95e-19
C7218 clknet_2_0__leaf_clk sample 0.236f
C7219 _074_ a_5997_10927# 9.52e-21
C7220 net9 a_13059_4631# 3.47e-19
C7221 a_2601_3285# cal 2.1e-20
C7222 _073_ a_7723_6807# 0.111f
C7223 clknet_2_1__leaf_clk a_6741_7361# 1.63e-19
C7224 _093_ a_2309_2229# 3.73e-21
C7225 a_10373_1679# VPWR 3.65e-19
C7226 _049_ a_4091_4943# 2.36e-20
C7227 mask\[2\] a_3053_8457# 0.0456f
C7228 _063_ a_9084_4515# 1.54e-20
C7229 a_10239_9295# VPWR 0.697f
C7230 _077_ net51 1.67e-19
C7231 net55 _089_ 3.16e-19
C7232 _045_ a_6987_12393# 1.15e-19
C7233 net27 a_7824_11305# 0.00103f
C7234 _023_ a_1313_10901# 8.7e-19
C7235 a_579_10933# a_1095_11305# 0.115f
C7236 clk ctln[6] 1.18e-20
C7237 a_14807_8359# a_14335_7895# 0.00179f
C7238 a_14236_8457# _132_ 0.00342f
C7239 trim_val\[0\] _058_ 0.0634f
C7240 a_816_6031# net30 4.57e-19
C7241 _033_ a_10543_2455# 4.61e-19
C7242 net45 a_395_7119# 2.93e-20
C7243 net37 _061_ 0.00617f
C7244 _097_ net1 3.15e-20
C7245 a_12436_9129# a_11895_7669# 1.06e-20
C7246 a_11987_8757# a_12344_8041# 8.3e-21
C7247 net15 a_2857_5461# 0.0194f
C7248 mask\[6\] mask\[5\] 0.017f
C7249 mask\[3\] a_2368_9955# 0.173f
C7250 a_10699_3311# a_9595_1679# 2.3e-20
C7251 a_3597_10933# a_4055_10927# 0.0346f
C7252 _029_ a_13091_4943# 0.285f
C7253 _104_ a_9361_3677# 4.96e-19
C7254 _046_ VPWR 0.782f
C7255 en_co_clk _096_ 0.0308f
C7256 trim_mask\[0\] a_14347_4917# 0.107f
C7257 a_13441_6281# VPWR 0.00591f
C7258 clknet_2_0__leaf_clk a_4036_8207# 0.00139f
C7259 a_448_7637# result[2] 7.83e-19
C7260 net26 _020_ 3.23e-19
C7261 _110_ trim_mask\[1\] 0.0802f
C7262 net29 _074_ 3.58e-19
C7263 _024_ a_11057_4105# 0.00732f
C7264 a_5067_9661# VPWR 0.138f
C7265 _074_ a_816_4765# 0.00471f
C7266 _088_ a_7758_4759# 1.25e-20
C7267 _129_ a_14422_7093# 0.0652f
C7268 a_9761_1679# ctln[4] 3.05e-19
C7269 trim_mask\[0\] _119_ 0.0387f
C7270 a_7631_12319# a_7259_11305# 0.00141f
C7271 _101_ a_3521_9813# 0.0432f
C7272 trim_mask\[2\] a_12870_2589# 5.43e-19
C7273 _078_ mask\[4\] 0.174f
C7274 _074_ _040_ 4.02e-21
C7275 cal_count\[3\] a_8307_4943# 4.56e-19
C7276 a_12231_6005# _108_ 1.43e-20
C7277 _099_ a_4815_3031# 1.08e-21
C7278 _028_ a_9004_3677# 4.1e-20
C7279 a_11814_9295# cal_count\[0\] 0.0857f
C7280 _090_ a_4471_4007# 8.83e-19
C7281 net12 a_6763_5193# 0.00146f
C7282 _104_ a_7939_3855# 0.0483f
C7283 net3 a_3667_3829# 0.0238f
C7284 a_4512_11305# net53 2.71e-20
C7285 _094_ a_5694_6031# 2.57e-19
C7286 net44 a_5455_4943# 4.7e-21
C7287 _051_ a_9207_3311# 7.37e-21
C7288 a_8091_7967# _063_ 3.38e-19
C7289 a_4167_6575# _049_ 0.0032f
C7290 net45 a_2659_2601# 0.153f
C7291 _129_ _132_ 0.319f
C7292 a_10699_5487# trim_mask\[1\] 1.57e-21
C7293 _027_ a_9719_1473# 1.64e-21
C7294 net39 trimb[3] 0.0254f
C7295 net13 a_4036_8207# 3.09e-19
C7296 _110_ a_8749_3317# 0.0134f
C7297 _107_ _028_ 7.9e-19
C7298 _128_ a_13470_7663# 7.48e-19
C7299 a_2953_7119# a_3399_7119# 2.28e-19
C7300 a_3521_7361# a_4030_7485# 2.6e-19
C7301 _074_ a_3431_12021# 0.0119f
C7302 net40 a_11067_4405# 8.8e-20
C7303 clknet_2_0__leaf_clk a_3123_3615# 3.04e-21
C7304 _048_ a_5081_4943# 0.0341f
C7305 a_8360_10383# a_8551_10383# 4.61e-19
C7306 net33 _129_ 2.66e-19
C7307 clknet_0_clk a_8749_3317# 7.24e-19
C7308 clknet_2_1__leaf_clk a_4043_11305# 3.39e-19
C7309 a_1095_11305# a_395_9845# 9.08e-19
C7310 clknet_0_clk _060_ 1.05e-20
C7311 _122_ cal_count\[2\] 0.224f
C7312 _108_ a_13697_4373# 0.00934f
C7313 a_11023_5108# _058_ 0.0034f
C7314 _051_ _050_ 0.567f
C7315 net55 _048_ 0.907f
C7316 a_10787_1135# ctln[4] 0.00151f
C7317 a_9664_3689# a_9826_3311# 0.00645f
C7318 _133_ _136_ 7.12e-19
C7319 _075_ _095_ 8.5e-20
C7320 _066_ VPWR 0.621f
C7321 net50 a_10699_3311# 0.00549f
C7322 _070_ a_9677_8457# 1.38e-19
C7323 net20 _078_ 1.54e-19
C7324 net9 a_13257_4943# 2.35e-19
C7325 a_1099_12533# a_1095_12393# 0.00343f
C7326 net34 a_15083_4659# 0.0191f
C7327 a_1476_10217# a_1638_9839# 0.00645f
C7328 _090_ a_4970_4399# 0.0146f
C7329 _049_ _028_ 0.00101f
C7330 a_8912_2589# ctln[5] 4.12e-20
C7331 en_co_clk a_5455_4943# 0.00555f
C7332 net49 a_14649_3689# 1.84e-19
C7333 a_395_7119# a_2953_7119# 1.77e-21
C7334 net18 _069_ 1.21e-20
C7335 a_13607_4943# trim_val\[0\] 1.9e-19
C7336 _058_ a_10055_2767# 1.08e-19
C7337 a_14335_2442# net48 0.109f
C7338 _027_ a_9595_1679# 6.08e-20
C7339 _051_ _052_ 0.0393f
C7340 a_4175_4943# VPWR 6.97e-20
C7341 _046_ net27 0.0365f
C7342 _021_ a_7521_11293# 7.78e-20
C7343 a_6743_10933# a_7933_11305# 2.56e-19
C7344 _031_ a_13393_1707# 6.16e-19
C7345 net48 net8 0.0209f
C7346 a_8215_9295# cal_itt\[0\] 1.43e-19
C7347 _000_ a_8993_9295# 3.81e-19
C7348 _049_ a_3751_4765# 7.78e-20
C7349 a_8083_8181# net2 0.0392f
C7350 a_6485_8181# a_6741_7361# 8.62e-21
C7351 a_7263_7093# a_7442_7119# 0.0074f
C7352 mask\[1\] net22 1.8e-20
C7353 net51 a_6173_7119# 0.00189f
C7354 a_7088_7119# a_7197_7119# 0.00742f
C7355 clknet_2_1__leaf_clk a_4687_11231# 5.54e-20
C7356 _092_ _038_ 0.00841f
C7357 a_3053_8207# VPWR 2.99e-19
C7358 trim_mask\[0\] a_11679_4777# 5.51e-21
C7359 _051_ _098_ 0.00409f
C7360 clknet_2_1__leaf_clk net44 0.0466f
C7361 net43 mask\[6\] 0.414f
C7362 _041_ a_5535_8181# 3.39e-20
C7363 _048_ a_7715_3285# 2.41e-23
C7364 a_5087_3855# a_6519_3829# 2.84e-20
C7365 _110_ _115_ 0.00253f
C7366 net31 trimb[1] 0.109f
C7367 _096_ _059_ 0.0162f
C7368 a_10699_5487# a_10781_5807# 0.00393f
C7369 a_11545_9049# VPWR 0.149f
C7370 _078_ a_2815_9447# 0.0114f
C7371 _101_ a_2775_9071# 3.77e-19
C7372 net14 a_2857_5461# 7.11e-22
C7373 net30 net42 0.00662f
C7374 a_6737_4719# a_6822_4399# 8.13e-19
C7375 _099_ a_5087_3855# 7.04e-20
C7376 _118_ a_9662_3855# 3.03e-20
C7377 a_11895_7669# a_13470_7663# 4.5e-20
C7378 _037_ a_12900_7663# 1.39e-19
C7379 net19 _071_ 4.17e-19
C7380 net4 a_2309_2229# 0.0134f
C7381 net18 a_11488_4765# 0.0021f
C7382 a_7571_4943# VPWR 0.205f
C7383 _078_ a_1313_10901# 0.0108f
C7384 _023_ result[5] 8.38e-19
C7385 _076_ _070_ 2.23e-20
C7386 a_9747_2527# _116_ 1.78e-20
C7387 a_7456_12393# VPWR 0.302f
C7388 net2 a_11709_6273# 1.57e-22
C7389 a_6007_7119# a_6741_7361# 0.0701f
C7390 _003_ a_6173_7119# 0.221f
C7391 _104_ a_10373_1679# 1.17e-20
C7392 a_3521_7361# a_3977_7119# 4.2e-19
C7393 a_14099_1929# a_13257_1141# 4.55e-20
C7394 a_9719_1473# _117_ 0.114f
C7395 _022_ a_3521_9813# 7.48e-20
C7396 net8 a_13091_1141# 0.013f
C7397 a_1476_4777# _099_ 1.31e-19
C7398 net28 _074_ 0.0147f
C7399 _021_ a_6909_10933# 0.234f
C7400 _074_ a_5177_9537# 0.0107f
C7401 a_6743_10933# a_7477_10901# 0.0694f
C7402 _042_ a_4655_10071# 5.2e-19
C7403 _043_ a_6467_9845# 8.03e-22
C7404 a_4576_3427# VPWR 0.176f
C7405 clknet_0_clk a_7939_3855# 0.00186f
C7406 a_12992_8751# a_13100_8751# 0.00523f
C7407 net46 a_13625_3317# 0.0553f
C7408 a_12344_8041# cal_count\[3\] 1.54e-19
C7409 _065_ a_9919_6614# 1.25e-20
C7410 a_11067_4405# _024_ 0.213f
C7411 net16 a_14604_2339# 0.00422f
C7412 net4 a_5691_2741# 0.0367f
C7413 a_1585_10217# result[4] 6.14e-21
C7414 net16 a_13557_7369# 3.42e-20
C7415 _065_ a_3781_8207# 4.41e-20
C7416 a_1129_4373# a_1476_4777# 0.0512f
C7417 clknet_0_clk a_4498_4373# 2.86e-21
C7418 _091_ a_9595_5193# 1.14e-19
C7419 _101_ a_6523_7119# 4.44e-21
C7420 net50 _027_ 0.002f
C7421 clknet_2_2__leaf_clk a_7379_2197# 3.85e-19
C7422 _071_ cal_itt\[1\] 6.15e-19
C7423 _043_ VPWR 0.484f
C7424 _078_ _081_ 0.0714f
C7425 a_6515_6794# VPWR 0.263f
C7426 a_8767_591# ctln[5] 0.16f
C7427 _108_ a_13825_5185# 0.0315f
C7428 _002_ a_7613_8029# 0.0023f
C7429 net23 a_3781_8207# 6.01e-21
C7430 net45 a_2313_6183# 0.00161f
C7431 _122_ cal_count\[1\] 0.201f
C7432 cal_itt\[0\] a_8298_5487# 0.00811f
C7433 _048_ _093_ 0.153f
C7434 net46 a_12310_4399# 3.35e-19
C7435 cal_count\[0\] a_12992_8751# 0.0796f
C7436 net45 a_4959_1679# 0.153f
C7437 _085_ a_1660_12393# 1.44e-20
C7438 _032_ a_10195_1354# 0.109f
C7439 net16 net2 0.203f
C7440 a_9595_1679# _117_ 0.00205f
C7441 _067_ a_11425_5487# 4.22e-21
C7442 net37 net40 0.016f
C7443 net46 a_8583_3317# 0.296f
C7444 net53 a_5829_9839# 8.05e-19
C7445 net44 a_7245_10205# 0.00215f
C7446 _059_ a_5455_4943# 0.00764f
C7447 clknet_2_2__leaf_clk a_9664_3689# 0.00144f
C7448 net24 a_1476_7119# 3.38e-21
C7449 a_14981_4020# a_14715_3615# 0.00139f
C7450 net16 a_14193_3285# 0.00842f
C7451 net24 mask\[0\] 3.77e-20
C7452 net34 _133_ 2.23e-20
C7453 a_1211_7983# a_1125_7663# 2.42e-19
C7454 a_12061_7669# a_10877_7983# 5.7e-21
C7455 _074_ a_4167_11471# 1.62e-19
C7456 trim_mask\[0\] calibrate 4.16e-20
C7457 a_8215_9295# a_10405_9295# 7.98e-21
C7458 a_8381_9295# a_10239_9295# 0.00228f
C7459 net30 a_8491_2229# 6.12e-20
C7460 net4 _091_ 0.0128f
C7461 clknet_2_2__leaf_clk a_10689_2223# 6.37e-21
C7462 _038_ a_11045_5807# 1.97e-19
C7463 _119_ a_8298_2767# 0.151f
C7464 en_co_clk a_13111_6031# 1.4e-19
C7465 a_1638_4399# VPWR 5.74e-19
C7466 _075_ calibrate 1.61e-20
C7467 _049_ _094_ 0.166f
C7468 net16 a_14000_4719# 8.6e-20
C7469 _036_ a_13142_8359# 0.106f
C7470 _060_ net41 0.161f
C7471 trim_val\[2\] a_13869_1501# 9.25e-20
C7472 net32 a_14071_3689# 1.09e-19
C7473 a_7088_7119# a_7250_7485# 0.00645f
C7474 a_6523_7119# a_6785_7119# 0.00171f
C7475 a_6741_7361# cal_itt\[3\] 3.97e-19
C7476 a_10903_7261# a_10990_7485# 0.0701f
C7477 net8 a_14281_1513# 5.59e-19
C7478 a_3557_5193# VPWR 0.00217f
C7479 a_9471_9269# VPWR 0.453f
C7480 a_11343_3317# a_13625_3317# 2.74e-21
C7481 a_7456_12393# net27 0.00276f
C7482 a_11859_3689# a_12424_3689# 7.99e-20
C7483 _034_ _048_ 2.06e-21
C7484 a_929_8757# a_2006_8751# 1.46e-19
C7485 net9 net40 0.0692f
C7486 net47 a_14377_7983# 1.15e-19
C7487 _039_ result[0] 2.93e-19
C7488 _055_ a_14604_3017# 0.105f
C7489 _122_ _108_ 4.53e-21
C7490 _063_ a_9802_4007# 3.67e-19
C7491 a_911_6031# a_816_6031# 0.0498f
C7492 a_5915_10927# _008_ 2.07e-21
C7493 a_561_6031# a_1638_6397# 1.46e-19
C7494 net44 a_6485_8181# 2.17e-19
C7495 cal_count\[0\] a_15111_9295# 5.23e-19
C7496 _074_ net21 0.474f
C7497 mask\[4\] a_6888_10205# 0.0249f
C7498 net47 a_12546_9129# 1.16e-19
C7499 clknet_2_3__leaf_clk _070_ 2.49e-20
C7500 state\[2\] a_4901_2773# 1.57e-21
C7501 _058_ net32 0.00353f
C7502 net16 net31 4.4e-20
C7503 net15 a_2787_9845# 0.0128f
C7504 clknet_2_0__leaf_clk a_3529_6281# 1.76e-21
C7505 clknet_2_1__leaf_clk a_4801_9839# 6.27e-22
C7506 net12 mask\[4\] 0.105f
C7507 net43 result[0] 6.17e-20
C7508 a_4443_9295# a_5633_9295# 2.56e-19
C7509 a_7001_7669# a_7447_8041# 2.28e-19
C7510 a_1830_4765# VPWR 4.59e-19
C7511 _063_ _108_ 6.65e-19
C7512 cal_count\[2\] comp 8.28e-20
C7513 a_6541_12021# a_6796_12381# 0.0642f
C7514 a_6743_10933# VPWR 0.455f
C7515 net50 _117_ 9.65e-19
C7516 state\[0\] a_4901_2773# 1.53e-19
C7517 _084_ a_6197_12015# 0.00265f
C7518 net4 a_4609_1679# 1.57e-19
C7519 _123_ cal_itt\[1\] 4.01e-20
C7520 trim_mask\[4\] _028_ 0.0918f
C7521 a_8583_3317# a_11343_3317# 1.59e-21
C7522 _065_ _124_ 5.23e-20
C7523 net45 a_5878_1679# 0.00288f
C7524 a_3781_8207# a_4696_8207# 0.119f
C7525 a_3615_8207# a_5535_8181# 2.73e-21
C7526 a_2971_8457# net30 7.56e-21
C7527 a_4091_5309# state\[0\] 1.68e-21
C7528 _076_ a_4349_8449# 3.49e-21
C7529 a_2787_7119# _049_ 0.0011f
C7530 mask\[6\] a_2953_9845# 7.54e-20
C7531 a_8298_5487# trim_mask\[0\] 0.127f
C7532 net19 a_9043_6031# 0.00109f
C7533 a_12056_6031# VPWR 0.297f
C7534 trim_mask\[1\] a_11057_4105# 0.00342f
C7535 a_11244_9661# _001_ 2.61e-19
C7536 net44 a_6007_7119# 0.304f
C7537 cal_count\[0\] a_14422_7093# 4.7e-20
C7538 a_579_12021# a_448_11445# 3.9e-19
C7539 a_8022_7119# a_8307_6575# 0.012f
C7540 net18 a_10569_1109# 0.00275f
C7541 mask\[4\] a_6983_10217# 0.0356f
C7542 net17 a_12341_8751# 8.46e-20
C7543 a_11436_9295# _122_ 1.73e-19
C7544 a_14335_4020# a_14335_2442# 5.35e-19
C7545 net49 a_14686_3017# 3.05e-19
C7546 a_3868_10217# _019_ 4.75e-19
C7547 a_12056_6031# a_12218_6397# 0.00645f
C7548 _078_ result[5] 4.73e-20
C7549 a_11491_6031# a_11753_6031# 0.00171f
C7550 net47 a_10903_7261# 0.301f
C7551 a_11987_8757# _129_ 4.2e-20
C7552 net20 net12 0.103f
C7553 a_14071_3689# VPWR 8.68e-19
C7554 _001_ a_11204_7485# 1.44e-20
C7555 clknet_2_1__leaf_clk a_1184_9117# 2.63e-20
C7556 a_7916_8041# _071_ 2.83e-19
C7557 _063_ a_9460_6807# 5.74e-19
C7558 mask\[0\] a_1129_6273# 7.07e-20
C7559 net45 VPWR 4.53f
C7560 _105_ a_8307_4719# 1.18e-19
C7561 _101_ a_4512_11305# 2.63e-19
C7562 a_3123_3615# a_2948_3689# 0.234f
C7563 a_13279_8207# VPWR 0.00846f
C7564 _058_ VPWR 1.27f
C7565 net52 _017_ 0.0168f
C7566 _049_ a_4617_3855# 1.84e-19
C7567 a_6519_3829# a_6822_4105# 0.00145f
C7568 cal_count\[0\] _132_ 8.08e-21
C7569 net29 a_1835_12319# 0.0966f
C7570 a_1644_12533# a_1660_12393# 7.19e-19
C7571 net34 _129_ 9.43e-20
C7572 net12 _053_ 0.00965f
C7573 a_455_3571# a_1867_3317# 1.6e-21
C7574 _044_ VPWR 0.512f
C7575 clknet_2_1__leaf_clk a_2910_12131# 6.18e-21
C7576 a_1461_10357# a_1476_10217# 4.33e-19
C7577 _120_ a_4259_6031# 6.92e-19
C7578 a_13512_1501# a_13703_1513# 4.61e-19
C7579 net40 a_10188_4105# 4.36e-20
C7580 _136_ a_12323_4703# 0.00212f
C7581 a_6007_7119# clk 1.37e-20
C7582 _123_ _001_ 0.0103f
C7583 a_14540_3689# a_15299_3311# 4.54e-19
C7584 net33 cal_count\[0\] 0.00507f
C7585 a_12992_8751# a_13919_8751# 4.27e-19
C7586 net44 _092_ 7.09e-20
C7587 a_4498_4373# net41 4.77e-21
C7588 a_9693_8029# VPWR 1.68e-19
C7589 cal_itt\[2\] a_8025_8041# 1.19e-20
C7590 net46 a_14894_3677# 0.00288f
C7591 a_14604_3017# trim_val\[2\] 5.43e-19
C7592 _102_ a_1822_10927# 5.01e-20
C7593 _112_ a_13693_3883# 6.69e-19
C7594 mask\[5\] _021_ 9.18e-20
C7595 a_5829_9839# a_6007_9839# 1.95e-20
C7596 a_9195_10357# a_9020_10383# 0.234f
C7597 mask\[4\] a_8551_10383# 4.1e-19
C7598 a_8455_10383# _043_ 1.57e-20
C7599 net9 _024_ 2.6e-20
C7600 net4 _048_ 0.00405f
C7601 cal_count\[2\] a_13111_6031# 8.29e-19
C7602 _097_ a_2143_2229# 4.22e-21
C7603 _084_ a_6099_10633# 1.18e-20
C7604 net43 a_1497_8725# 0.166f
C7605 _135_ trim_mask\[0\] 2.05e-20
C7606 clknet_2_2__leaf_clk _057_ 2.3e-19
C7607 _063_ _107_ 0.019f
C7608 _096_ a_4725_5487# 0.0114f
C7609 net1 a_2288_3677# 1.29e-20
C7610 a_1660_12393# a_2828_12131# 7.54e-20
C7611 net27 a_6743_10933# 2.02e-19
C7612 a_6999_12015# _021_ 6.03e-21
C7613 a_3868_10217# VPWR 0.304f
C7614 a_8105_10383# net47 0.0258f
C7615 net43 _073_ 1.23e-19
C7616 a_7010_3311# a_7010_3631# 0.00278f
C7617 a_1129_6273# _079_ 3.2e-19
C7618 _122_ a_12900_7663# 0.0353f
C7619 net19 a_8749_3317# 0.014f
C7620 _012_ a_937_4105# 0.0526f
C7621 _033_ _027_ 2.18e-19
C7622 _051_ a_7891_3617# 0.13f
C7623 net51 a_7351_8041# 0.00137f
C7624 a_8298_2767# a_9225_2197# 0.00656f
C7625 _092_ clk 0.034f
C7626 a_1476_10217# _018_ 5.62e-19
C7627 net25 a_2787_9845# 9.67e-20
C7628 _004_ a_455_5747# 0.0445f
C7629 a_395_6031# net30 1.97e-19
C7630 en_co_clk _092_ 0.274f
C7631 _047_ a_14981_4020# 0.191f
C7632 net44 cal_itt\[3\] 0.0612f
C7633 _093_ a_2033_3317# 6.32e-20
C7634 net18 a_11374_1251# 3.05e-19
C7635 net16 a_14083_3311# 0.0056f
C7636 net40 _062_ 0.122f
C7637 a_6927_12559# net44 0.00394f
C7638 net19 a_6375_12021# 6.86e-20
C7639 _063_ _049_ 9.1e-20
C7640 a_7201_9813# a_7710_9839# 2.6e-19
C7641 a_6983_10217# a_7091_9839# 0.0572f
C7642 a_7548_10217# a_7657_10217# 0.00742f
C7643 a_9225_2197# a_9681_2601# 4.2e-19
C7644 a_7723_10143# a_7902_10205# 0.0074f
C7645 _066_ a_10699_5487# 0.278f
C7646 net55 a_6197_4399# 0.00361f
C7647 a_8949_6281# a_8298_5487# 2.65e-19
C7648 _107_ a_7104_3855# 8.79e-20
C7649 a_11059_7356# a_11016_6691# 4.89e-19
C7650 _131_ a_15023_5487# 4.38e-22
C7651 _096_ _107_ 3.94e-19
C7652 clknet_2_0__leaf_clk a_7263_7093# 1.09e-20
C7653 a_14379_6397# _136_ 1.29e-19
C7654 _135_ a_13933_6281# 0.00605f
C7655 clknet_2_1__leaf_clk result[3] 0.0234f
C7656 a_2953_7119# VPWR 0.561f
C7657 net2 clkc 3.18e-19
C7658 _063_ a_8495_6895# 0.131f
C7659 _043_ a_8381_9295# 5.52e-19
C7660 a_9195_10357# a_8731_9295# 3.62e-19
C7661 mask\[6\] mask\[3\] 8.02e-19
C7662 net43 ctlp[7] 1.17e-19
C7663 cal_itt\[3\] clk 0.0472f
C7664 net27 _044_ 0.00619f
C7665 clknet_0_clk a_7571_4943# 8.82e-22
C7666 cal_itt\[3\] en_co_clk 1.08e-19
C7667 a_9296_9295# a_9405_9295# 0.00742f
C7668 _035_ cal_count\[0\] 2.29e-19
C7669 a_11394_9509# a_11244_9661# 0.344f
C7670 a_9471_9269# a_9650_9295# 0.0074f
C7671 trim_mask\[0\] a_13519_4007# 2.23e-19
C7672 _022_ a_4512_11305# 1.61e-19
C7673 a_6906_2355# clk 9.3e-19
C7674 _049_ a_7104_3855# 0.0101f
C7675 a_13607_4943# VPWR 0.207f
C7676 a_9572_2601# a_11435_2229# 2.73e-20
C7677 a_1313_10901# a_1651_10143# 1.09e-20
C7678 a_745_10933# a_1476_10217# 4.77e-21
C7679 net19 a_7986_10927# 3.32e-20
C7680 a_1095_11305# a_911_10217# 1.3e-20
C7681 _049_ _096_ 0.0741f
C7682 _038_ _136_ 0.0457f
C7683 a_11067_4405# trim_mask\[1\] 6.42e-19
C7684 _024_ a_10188_4105# 9.19e-21
C7685 _009_ net44 0.0049f
C7686 _096_ a_3388_4631# 0.318f
C7687 mask\[1\] a_4030_7485# 8.1e-21
C7688 net22 a_561_6031# 0.21f
C7689 a_745_10933# _007_ 1.42e-19
C7690 _023_ a_561_9845# 4.6e-19
C7691 net48 trim[2] 2.08e-19
C7692 a_1844_9129# net23 0.00161f
C7693 a_13783_6183# trim_val\[0\] 2.33e-21
C7694 _048_ a_6763_5193# 2.69e-19
C7695 a_1099_12533# a_745_10933# 3.39e-21
C7696 a_1095_12393# a_1357_12381# 0.00171f
C7697 net3 a_3339_2767# 0.0249f
C7698 _057_ ctln[2] 0.0674f
C7699 a_4905_3855# VPWR 1.97e-19
C7700 net18 a_10975_4105# 0.0106f
C7701 net52 a_1764_10383# 8.16e-20
C7702 a_1476_7119# a_3208_7119# 4.21e-21
C7703 clknet_2_3__leaf_clk net50 3.78e-21
C7704 _006_ net23 0.00178f
C7705 mask\[0\] a_3208_7119# 0.0264f
C7706 a_3399_10217# VPWR 2.07e-19
C7707 a_3922_8867# VPWR 0.00128f
C7708 cal_itt\[0\] _041_ 0.0129f
C7709 net28 a_1835_12319# 2.21e-19
C7710 _051_ _087_ 0.316f
C7711 a_8298_5487# a_8307_4943# 0.00344f
C7712 net9 _029_ 0.00231f
C7713 clknet_2_0__leaf_clk a_1493_5487# 0.0654f
C7714 _071_ a_8949_6031# 9.76e-19
C7715 _101_ a_5829_9839# 9.22e-19
C7716 net45 a_2383_3689# 0.156f
C7717 a_11394_9509# _123_ 3.03e-20
C7718 trim_mask\[2\] a_14099_1929# 0.0586f
C7719 net46 a_13512_4943# 0.0165f
C7720 a_14249_8725# a_14335_7895# 2.03e-20
C7721 a_11233_4405# a_12310_4399# 1.46e-19
C7722 a_9084_4515# a_9317_3285# 4.53e-19
C7723 a_455_8181# a_561_7119# 1.55e-19
C7724 mask\[7\] net52 0.199f
C7725 net53 a_7367_10927# 6.01e-19
C7726 a_561_9845# a_816_10205# 0.0594f
C7727 net31 clkc 0.146f
C7728 _065_ a_4680_6031# 1.52e-19
C7729 net9 a_11244_9661# 0.00191f
C7730 _078_ a_3781_8207# 3.94e-19
C7731 a_6316_5193# VPWR 0.136f
C7732 _051_ _099_ 0.012f
C7733 net19 a_7824_11305# 0.00166f
C7734 a_8949_9537# a_8731_9295# 0.21f
C7735 a_8381_9295# a_9471_9269# 0.0425f
C7736 net45 _104_ 2.79e-21
C7737 a_2857_5461# VPWR 1.3f
C7738 a_5455_4943# _107_ 0.00327f
C7739 a_6007_7119# a_7197_7119# 2.56e-19
C7740 mask\[4\] a_9871_10383# 0.049f
C7741 _092_ _059_ 0.289f
C7742 net44 a_4805_8207# 6.59e-20
C7743 _099_ _014_ 0.0885f
C7744 _076_ net2 0.44f
C7745 _074_ a_1007_6031# 0.00166f
C7746 a_1476_7119# result[1] 3.76e-19
C7747 a_3116_12533# _010_ 0.0629f
C7748 _078_ a_395_4405# 6.64e-20
C7749 clknet_2_1__leaf_clk a_2787_10927# 0.0348f
C7750 _069_ VPWR 0.288f
C7751 _048_ a_9166_4515# 5.59e-19
C7752 _058_ _104_ 0.00402f
C7753 a_4993_6273# net54 1.02e-19
C7754 net19 a_8935_6895# 0.00661f
C7755 a_1476_4777# _097_ 2.42e-20
C7756 trim_val\[3\] ctln[4] 0.00181f
C7757 net44 a_5547_5603# 2.28e-19
C7758 clk cal 2.95e-20
C7759 a_8022_7119# VPWR 1.33f
C7760 a_11116_8983# _123_ 0.202f
C7761 a_1844_9129# a_2225_7663# 6.06e-22
C7762 cal_itt\[2\] a_6173_7119# 8.89e-21
C7763 a_1129_4373# _014_ 1.89e-20
C7764 a_8091_7967# cal_itt\[3\] 1.82e-20
C7765 net16 a_13715_5309# 0.00193f
C7766 a_11895_7669# _037_ 0.151f
C7767 _119_ a_9369_4105# 0.0111f
C7768 a_10655_2932# a_9761_1679# 5.89e-20
C7769 cal_count\[2\] a_14199_7369# 3.59e-19
C7770 a_10055_2767# a_10329_1921# 0.00111f
C7771 _049_ a_5455_4943# 6.98e-19
C7772 mask\[3\] a_1763_9295# 0.0105f
C7773 net9 a_13349_6031# 8.04e-19
C7774 net9 _123_ 0.0156f
C7775 mask\[6\] a_4043_11305# 0.00432f
C7776 _078_ a_1579_11471# 7.62e-19
C7777 net44 a_5536_4399# 9.65e-21
C7778 net53 a_7999_11231# 2.43e-21
C7779 net43 a_8078_7663# 2.53e-19
C7780 a_763_8757# _005_ 9.51e-20
C7781 _045_ a_5496_12131# 0.106f
C7782 a_5997_10927# mask\[4\] 3.11e-19
C7783 a_14422_7093# en_co_clk 1.69e-19
C7784 a_4995_7119# a_5363_7369# 2.31e-19
C7785 net8 a_14184_1679# 3.26e-19
C7786 _081_ result[2] 5.8e-19
C7787 _127_ a_14983_9269# 0.0902f
C7788 a_14347_9480# _126_ 0.00393f
C7789 a_11488_4765# VPWR 0.0851f
C7790 _070_ a_6835_7669# 3.36e-21
C7791 _042_ _018_ 0.172f
C7792 a_10990_7485# a_11141_6031# 1.36e-20
C7793 cal_itt\[1\] a_8935_6895# 0.134f
C7794 en_co_clk a_5547_5603# 0.00658f
C7795 _091_ _064_ 0.003f
C7796 net46 a_11859_3689# 0.155f
C7797 _053_ a_5691_2741# 0.0314f
C7798 a_1313_10901# a_1191_11305# 3.16e-19
C7799 net12 a_7379_2197# 5.19e-20
C7800 a_1095_11305# a_1000_11293# 0.0498f
C7801 _074_ a_1019_7485# 0.00538f
C7802 _088_ a_7800_4631# 4e-20
C7803 net10 ctln[3] 3.57e-21
C7804 _065_ _017_ 6.2e-21
C7805 clknet_2_2__leaf_clk a_13625_3317# 8.94e-19
C7806 a_12992_8751# cal_count\[2\] 3.38e-21
C7807 net43 a_4655_10071# 0.00243f
C7808 a_7262_5461# a_7800_4631# 2.21e-20
C7809 _101_ a_4995_7119# 8.89e-19
C7810 trim_val\[0\] a_13881_2741# 2.93e-19
C7811 _113_ VPWR 0.355f
C7812 a_3386_2223# VPWR 5.3e-19
C7813 _132_ en_co_clk 1.15e-19
C7814 a_15023_9839# net2 3.29e-20
C7815 net23 _017_ 1.83e-20
C7816 mask\[6\] a_4687_11231# 0.129f
C7817 _071_ _062_ 2.92e-19
C7818 a_5067_2045# clk 0.0263f
C7819 en_co_clk a_5536_4399# 3.16e-19
C7820 mask\[6\] net44 2.19e-21
C7821 a_9084_4515# a_9003_3829# 0.00121f
C7822 a_8105_10383# _068_ 2.08e-22
C7823 a_14347_1439# a_14471_591# 9.9e-19
C7824 net45 a_1007_4777# 9.54e-19
C7825 net46 a_11845_4765# 0.00343f
C7826 a_10405_9295# _041_ 1.06e-19
C7827 net33 en_co_clk 4.99e-19
C7828 cal_count\[0\] a_11987_8757# 0.491f
C7829 a_3565_7119# _092_ 2.63e-21
C7830 a_579_12021# a_1203_12015# 9.73e-19
C7831 cal_itt\[3\] a_7197_7119# 1.52e-19
C7832 _063_ trim_mask\[4\] 1.61e-20
C7833 clknet_2_1__leaf_clk _049_ 5.62e-19
C7834 clknet_2_2__leaf_clk a_12310_4399# 2.27e-20
C7835 net15 net26 0.0071f
C7836 _042_ mask\[1\] 0.00296f
C7837 clknet_2_2__leaf_clk a_8583_3317# 0.252f
C7838 a_14335_4020# a_13459_3317# 4.72e-20
C7839 a_13519_4007# _030_ 3.44e-19
C7840 net13 net53 0.0143f
C7841 a_395_6031# a_1585_6031# 2.56e-19
C7842 _074_ a_1173_10205# 7.09e-19
C7843 trim_mask\[0\] a_9839_3615# 5.37e-20
C7844 clknet_2_1__leaf_clk a_7259_11305# 8.78e-19
C7845 clknet_2_3__leaf_clk _106_ 4.29e-19
C7846 a_995_3530# valid 1.27e-19
C7847 net47 a_9074_9955# 2.47e-19
C7848 net52 _121_ 2.08e-20
C7849 _076_ a_4883_6397# 1.38e-19
C7850 _053_ _091_ 3.98e-19
C7851 _020_ a_8360_10383# 0.158f
C7852 _078_ a_5686_9661# 1.91e-19
C7853 a_6099_10633# a_6181_10383# 0.00393f
C7854 net34 cal_count\[0\] 1.94e-19
C7855 a_1679_10633# a_1764_10383# 1.48e-19
C7856 a_11023_5108# a_10975_4105# 4.76e-21
C7857 trim[0] trim[2] 0.0391f
C7858 a_4621_11305# VPWR 1.19e-19
C7859 net45 clknet_0_clk 0.0745f
C7860 a_2283_4020# _013_ 0.109f
C7861 a_8657_2229# VPWR 0.589f
C7862 _078_ a_561_9845# 0.00812f
C7863 net43 a_3521_7361# 0.16f
C7864 clknet_2_3__leaf_clk net2 0.106f
C7865 _058_ _110_ 0.0486f
C7866 _010_ a_4043_12393# 5e-19
C7867 _074_ ctlp[1] 5.89e-19
C7868 net30 state\[2\] 9.58e-20
C7869 _123_ a_12436_9129# 0.0325f
C7870 net41 a_4576_3427# 0.0201f
C7871 cal_itt\[0\] a_9602_6614# 0.00697f
C7872 _002_ a_7569_7637# 0.0231f
C7873 net43 a_1129_7361# 0.175f
C7874 a_5694_6031# _092_ 3.4e-20
C7875 _115_ a_13512_1501# 5.13e-19
C7876 _065_ a_4425_6031# 0.00349f
C7877 _058_ a_12778_3677# 1.06e-19
C7878 mask\[7\] a_1679_10633# 0.0671f
C7879 net9 trim_mask\[1\] 0.00869f
C7880 trim_mask\[4\] a_7181_2589# 2.58e-19
C7881 a_9719_1473# _116_ 0.185f
C7882 net8 _057_ 0.159f
C7883 a_13257_1141# a_14172_1513# 0.125f
C7884 a_13091_1141# a_15023_1135# 4.36e-20
C7885 a_11343_3317# a_11859_3689# 0.111f
C7886 _025_ a_12077_3285# 1.82e-19
C7887 net31 a_15023_9839# 0.0146f
C7888 a_448_6549# result[1] 0.00288f
C7889 a_745_12021# a_1660_12393# 0.125f
C7890 net43 a_1095_12393# 0.157f
C7891 clknet_2_1__leaf_clk a_3947_12393# 0.0347f
C7892 cal_count\[1\] a_14199_7369# 6.02e-20
C7893 a_11244_9661# a_11508_9295# 0.00384f
C7894 a_12148_4777# _058_ 0.0142f
C7895 a_13059_4631# a_13697_4373# 0.00147f
C7896 a_10699_5487# _058_ 0.00216f
C7897 net46 a_9572_2601# 0.231f
C7898 a_14981_4020# net49 5.55e-21
C7899 _053_ a_12520_7637# 2.67e-20
C7900 a_395_6031# a_911_6031# 0.114f
C7901 _095_ a_2601_3285# 9.69e-20
C7902 a_6210_4989# VPWR 0.194f
C7903 net43 a_1638_9839# 1.09e-19
C7904 _125_ trimb[4] 0.00214f
C7905 net14 a_855_4105# 0.00997f
C7906 clknet_2_1__leaf_clk a_3425_11721# 0.0129f
C7907 a_5547_5603# _059_ 0.00252f
C7908 cal_count\[2\] a_14422_7093# 0.0242f
C7909 a_5221_1679# ctln[7] 2.48e-20
C7910 result[4] result[3] 0.0472f
C7911 _004_ a_395_4405# 1.61e-20
C7912 mask\[3\] a_1497_8725# 9.58e-19
C7913 net53 a_4864_9295# 5.51e-21
C7914 _017_ a_4696_8207# 1.49e-19
C7915 net45 a_2476_6281# 1.59e-19
C7916 a_7250_7485# _092_ 5.17e-21
C7917 a_9595_1679# _116_ 4.14e-20
C7918 a_13881_1653# a_13607_1513# 6.99e-19
C7919 a_12992_8751# cal_count\[1\] 0.0161f
C7920 _041_ a_11258_8790# 9.13e-19
C7921 _015_ a_4658_3427# 5.02e-19
C7922 a_10655_2932# a_11067_3017# 0.02f
C7923 a_4815_3031# a_4709_2773# 0.179f
C7924 net26 a_7548_10217# 0.0587f
C7925 _048_ _064_ 7.4e-21
C7926 _050_ trim_mask\[0\] 3.24e-20
C7927 net25 a_763_8757# 2.54e-19
C7928 a_395_9845# net24 2.97e-21
C7929 _071_ a_8745_6895# 0.00198f
C7930 a_9650_9295# _069_ 7.35e-20
C7931 net19 _066_ 8.99e-21
C7932 _065_ a_3868_7119# 8.33e-19
C7933 a_6523_7119# a_6515_6794# 3.36e-19
C7934 a_4167_11471# a_4055_10927# 1.26e-19
C7935 a_14715_3615# a_14604_2339# 1.68e-20
C7936 _092_ _108_ 7.49e-20
C7937 _059_ a_5536_4399# 0.0912f
C7938 _128_ _122_ 0.0325f
C7939 net40 a_14788_7369# 0.0078f
C7940 net46 a_14471_591# 8.79e-19
C7941 a_15023_8751# _131_ 3.38e-21
C7942 a_448_11445# _086_ 8.35e-19
C7943 net14 a_763_8757# 0.0121f
C7944 net12 a_5221_1679# 1.31e-19
C7945 _112_ a_14099_3017# 0.00116f
C7946 a_2787_9845# _019_ 7.83e-21
C7947 _075_ _050_ 0.059f
C7948 _132_ cal_count\[2\] 0.00622f
C7949 net29 a_1313_10901# 7.76e-20
C7950 clknet_2_1__leaf_clk _008_ 0.116f
C7951 a_15023_2767# trim[2] 0.00245f
C7952 a_2815_9447# _040_ 4.86e-21
C7953 _101_ a_3431_10933# 0.00168f
C7954 a_10569_1109# VPWR 0.209f
C7955 net33 cal_count\[2\] 3.22e-19
C7956 en_co_clk _136_ 0.00657f
C7957 _101_ a_929_8757# 2.73e-19
C7958 _101_ _062_ 3.72e-20
C7959 clknet_0_clk a_2953_7119# 0.00163f
C7960 a_2857_7637# a_3521_7361# 0.00668f
C7961 net26 net25 0.00158f
C7962 net18 trim_val\[4\] 1.73e-21
C7963 _038_ cal_count\[3\] 0.0219f
C7964 _134_ a_13915_4399# 7.39e-21
C7965 trim_mask\[0\] _098_ 0.00401f
C7966 a_9761_1679# a_10838_2045# 1.46e-19
C7967 _103_ a_7527_4631# 0.046f
C7968 a_3529_6281# _094_ 0.0129f
C7969 a_14564_6397# _058_ 7.15e-20
C7970 a_13607_4943# _110_ 1.5e-20
C7971 _096_ a_3123_3615# 6.93e-20
C7972 a_13625_3317# a_14540_3689# 0.125f
C7973 a_13050_7637# a_13142_7271# 0.00134f
C7974 net14 net26 0.00702f
C7975 a_13459_3317# a_15299_3311# 1.35e-20
C7976 mask\[4\] a_5177_9537# 2.91e-20
C7977 a_12153_8757# a_13562_8751# 4.25e-19
C7978 a_12612_8725# a_12992_8751# 0.00971f
C7979 a_11987_8757# a_13919_8751# 1.08e-19
C7980 a_763_8757# a_395_7119# 6.48e-21
C7981 net9 _115_ 2.05e-20
C7982 _015_ a_5177_1921# 6.55e-19
C7983 _062_ a_9043_6031# 3.3e-19
C7984 a_3748_6281# _120_ 0.103f
C7985 cal_itt\[1\] a_10621_7119# 4.99e-19
C7986 clknet_2_1__leaf_clk a_5524_9295# 1.12e-19
C7987 a_1203_10927# _102_ 1.19e-19
C7988 _053_ _048_ 0.0572f
C7989 net52 _080_ 2.07e-22
C7990 a_3521_9813# a_3868_10217# 0.0512f
C7991 a_2953_9845# a_4655_10071# 1.67e-19
C7992 _080_ a_816_7119# 7.37e-19
C7993 _067_ a_9957_7663# 0.0492f
C7994 _092_ a_4725_5487# 0.00351f
C7995 cal_itt\[0\] a_10747_8970# 0.00199f
C7996 net19 a_7571_4943# 4.1e-22
C7997 trim_mask\[0\] a_14526_4943# 0.00222f
C7998 net46 a_13825_1109# 0.168f
C7999 _076_ a_4993_6273# 1.76e-19
C8000 a_10329_1921# VPWR 0.212f
C8001 _083_ _077_ 5.66e-20
C8002 _081_ _040_ 0.165f
C8003 net50 _116_ 0.00151f
C8004 net34 a_13919_8751# 3.57e-21
C8005 _078_ a_1844_9129# 0.0499f
C8006 a_911_6031# net30 1.21e-19
C8007 _123_ a_13470_7663# 0.00883f
C8008 state\[2\] state\[0\] 0.0763f
C8009 net19 a_7456_12393# 6.62e-19
C8010 a_2787_9845# VPWR 0.445f
C8011 a_13091_4943# _058_ 0.00986f
C8012 a_13257_4943# a_13697_4373# 0.00351f
C8013 trim_mask\[1\] trim_mask\[3\] 1.44e-19
C8014 trim_mask\[2\] a_13183_3311# 8.82e-19
C8015 a_5496_12131# _078_ 0.00101f
C8016 _078_ _006_ 3.87e-19
C8017 _122_ a_11895_7669# 0.00249f
C8018 a_6885_8372# _072_ 8.44e-21
C8019 _051_ a_9503_4399# 1.79e-20
C8020 a_8949_9537# _063_ 7.96e-20
C8021 _016_ a_3868_7119# 1.93e-19
C8022 a_6007_7119# _049_ 8.61e-19
C8023 _108_ a_9317_3285# 0.00893f
C8024 net45 net41 0.413f
C8025 _097_ a_1867_3317# 0.00526f
C8026 _065_ a_10903_7261# 0.0109f
C8027 net31 a_14715_3615# 0.0177f
C8028 _028_ a_6941_2589# 2.52e-19
C8029 cal_itt\[3\] a_9460_6807# 4.72e-20
C8030 a_3431_10933# _102_ 3.99e-21
C8031 _042_ _041_ 4.99e-19
C8032 cal_count\[1\] a_14422_7093# 4.98e-21
C8033 a_7379_2197# a_7524_2223# 0.0572f
C8034 a_8491_2229# a_9103_2601# 3.82e-19
C8035 _027_ a_8912_2589# 0.17f
C8036 net19 _043_ 0.0119f
C8037 a_6467_9845# a_7657_10217# 2.56e-19
C8038 _092_ _107_ 0.0107f
C8039 a_15299_3311# trim[2] 8.78e-19
C8040 a_8298_5487# a_9369_4105# 2.66e-21
C8041 _104_ a_8657_2229# 1.8e-20
C8042 net46 a_13307_1707# 0.0121f
C8043 cal_itt\[2\] a_7351_8041# 9.12e-20
C8044 clknet_0_clk a_2857_5461# 0.346f
C8045 a_448_10357# result[3] 1.88e-20
C8046 _066_ a_11067_4405# 1.59e-20
C8047 a_13783_6183# VPWR 0.341f
C8048 _074_ a_7109_11989# 1.75e-20
C8049 net4 a_1276_565# 0.0302f
C8050 mask\[6\] a_2910_12131# 1.07e-19
C8051 a_4165_11989# a_4055_12015# 0.0977f
C8052 _125_ _130_ 4.49e-21
C8053 a_11374_1251# VPWR 0.00204f
C8054 _003_ a_7897_6913# 5.24e-20
C8055 en_co_clk a_4266_4943# 1.07e-19
C8056 clknet_2_0__leaf_clk a_5363_7369# 0.0417f
C8057 a_9839_3615# a_8298_2767# 0.0067f
C8058 net43 a_4866_11293# 0.00204f
C8059 a_11045_5807# _108_ 8.63e-21
C8060 a_4863_4917# _060_ 7.13e-20
C8061 clknet_0_clk a_8022_7119# 1.74f
C8062 a_7657_10217# VPWR 4.26e-20
C8063 a_2092_8457# VPWR 0.196f
C8064 net16 trimb[1] 4.04e-20
C8065 calibrate a_2601_3285# 6.54e-20
C8066 net49 trim_mask\[2\] 1.51e-19
C8067 cal_count\[1\] _132_ 1.61e-19
C8068 _049_ _092_ 0.291f
C8069 trim_mask\[1\] a_13415_2442# 1.93e-19
C8070 trim_mask\[3\] a_10977_2543# 0.00453f
C8071 a_8215_9295# a_9405_9295# 2.56e-19
C8072 net3 net54 0.195f
C8073 _035_ a_10688_9295# 0.0103f
C8074 _092_ a_3388_4631# 0.0622f
C8075 _062_ _060_ 0.0644f
C8076 a_10239_9295# a_11394_9509# 0.0608f
C8077 net45 a_6523_7119# 1e-21
C8078 a_13625_3317# a_14335_2442# 1.72e-20
C8079 a_3431_10933# _022_ 0.396f
C8080 _101_ clknet_2_0__leaf_clk 0.137f
C8081 net33 cal_count\[1\] 0.0109f
C8082 a_4959_9295# mask\[1\] 1.91e-19
C8083 net55 a_7800_4631# 0.0976f
C8084 net21 mask\[4\] 2.5e-19
C8085 _027_ a_10543_2455# 0.118f
C8086 a_14193_3285# a_14099_1929# 9.29e-21
C8087 a_3521_9813# a_3399_10217# 3.16e-19
C8088 _078_ result[7] 2.78e-20
C8089 a_3303_10217# a_3208_10205# 0.0498f
C8090 net30 _118_ 0.222f
C8091 trim_val\[0\] a_14281_4943# 3.85e-20
C8092 _090_ a_4815_3031# 2.65e-21
C8093 a_6191_12559# mask\[5\] 2.11e-21
C8094 net28 a_1313_10901# 9.18e-19
C8095 _078_ a_5633_9295# 1.61e-19
C8096 net16 a_13881_1653# 0.00258f
C8097 net44 _073_ 6.49e-20
C8098 a_11545_9049# _001_ 1.03e-19
C8099 _097_ a_3302_3677# 1.03e-19
C8100 net46 a_13715_1135# 0.0122f
C8101 _065_ _121_ 0.273f
C8102 cal_count\[2\] _136_ 9.64e-19
C8103 a_14379_6397# a_14347_4917# 1.11e-19
C8104 net22 a_1129_4373# 9.38e-20
C8105 state\[2\] _100_ 0.00152f
C8106 clknet_2_3__leaf_clk a_12249_7663# 0.00224f
C8107 mask\[2\] a_4349_8449# 1.96e-19
C8108 a_14347_9480# VPWR 0.179f
C8109 a_4775_6031# net30 1.27e-19
C8110 net34 en_co_clk 1.13e-19
C8111 net20 a_7810_12381# 1.27e-19
C8112 a_2198_9117# VPWR 3.65e-19
C8113 a_1835_11231# net52 0.0128f
C8114 _053_ a_7021_4105# 0.00863f
C8115 _014_ _097_ 0.0205f
C8116 cal_count\[0\] a_9463_8725# 1.46e-20
C8117 a_8749_3317# a_9195_3689# 2.28e-19
C8118 _110_ _113_ 0.255f
C8119 a_9003_3829# a_9802_4007# 0.00537f
C8120 a_1129_7361# a_1638_7485# 2.6e-19
C8121 a_911_7119# a_1019_7485# 0.0572f
C8122 a_15289_7119# net5 1.24e-19
C8123 a_7010_3311# clk 2.46e-19
C8124 net19 a_9471_9269# 1.08e-19
C8125 a_13142_7271# VPWR 0.298f
C8126 a_11141_6031# net46 0.0241f
C8127 net51 VPWR 0.641f
C8128 mask\[0\] a_1476_7119# 0.00229f
C8129 a_9207_3311# a_8298_2767# 0.00129f
C8130 net29 result[5] 6.48e-20
C8131 trim_mask\[2\] a_11601_2229# 4.46e-19
C8132 a_10239_9295# a_11116_8983# 1.64e-19
C8133 a_10405_9295# a_10747_8970# 0.00801f
C8134 a_10975_4105# VPWR 0.259f
C8135 cal_itt\[3\] _049_ 2.9e-21
C8136 a_12992_8751# a_12900_7663# 7.46e-19
C8137 net40 _037_ 3.14e-19
C8138 clknet_2_1__leaf_clk a_6891_12393# 2.56e-19
C8139 net13 _101_ 0.0171f
C8140 _108_ a_9003_3829# 0.333f
C8141 cal en 0.0365f
C8142 trim[1] trim[0] 0.0363f
C8143 net21 net20 0.00154f
C8144 _107_ a_9317_3285# 0.00133f
C8145 a_7800_4631# a_7715_3285# 2.38e-20
C8146 mask\[7\] _023_ 4.85e-19
C8147 mask\[3\] a_4655_10071# 0.0669f
C8148 net15 net55 1.07e-20
C8149 a_13257_4943# a_13825_5185# 0.175f
C8150 a_13091_4943# a_13607_4943# 0.112f
C8151 clknet_2_2__leaf_clk a_13512_4943# 0.00155f
C8152 _073_ clk 0.00414f
C8153 a_4055_12015# VPWR 0.143f
C8154 a_11435_2229# a_12625_2601# 2.56e-19
C8155 net9 a_10239_9295# 2.21e-19
C8156 _078_ _017_ 1.16e-19
C8157 net45 a_2767_2223# 0.0122f
C8158 _074_ _005_ 0.124f
C8159 net19 a_6743_10933# 3.72e-19
C8160 net16 a_14334_1135# 1.15e-20
C8161 _048_ a_3891_4943# 0.155f
C8162 a_14181_6031# VPWR 1.83e-19
C8163 _104_ a_10569_1109# 6.99e-22
C8164 a_12341_8751# a_12522_8751# 8.75e-19
C8165 _058_ a_11057_4105# 0.00327f
C8166 _002_ a_7723_6807# 5.1e-20
C8167 net33 _108_ 0.34f
C8168 cal_itt\[3\] a_8495_6895# 0.00223f
C8169 mask\[4\] _020_ 1.22e-19
C8170 clknet_2_1__leaf_clk a_9195_10357# 1.09e-20
C8171 _136_ a_12410_6031# 1.99e-19
C8172 _098_ a_8307_4943# 1.07e-20
C8173 a_9471_9269# cal_itt\[1\] 4.78e-20
C8174 a_9296_9295# a_9459_7895# 5.29e-21
C8175 net2 a_6835_7669# 1.9e-19
C8176 _110_ a_8657_2229# 0.00736f
C8177 trim_val\[4\] a_10055_2767# 0.00159f
C8178 net15 _074_ 0.00832f
C8179 net40 a_12231_6005# 1.69e-20
C8180 _072_ net42 1.06e-20
C8181 _003_ VPWR 0.418f
C8182 a_8298_5487# a_8307_4719# 1.92e-20
C8183 a_7460_5807# _088_ 1.17e-19
C8184 net44 a_9296_9295# 1.56e-20
C8185 net43 a_1461_10357# 0.0109f
C8186 _067_ a_10903_7261# 1.01e-19
C8187 a_13881_2741# VPWR 0.27f
C8188 a_561_9845# a_1651_10143# 0.0418f
C8189 _050_ a_7210_5807# 0.042f
C8190 a_7262_5461# a_7460_5807# 0.00788f
C8191 a_4863_4917# a_4498_4373# 3.62e-19
C8192 a_13975_3689# trim_val\[1\] 0.00171f
C8193 net9 a_13441_6281# 5.89e-20
C8194 a_14335_4020# trim[1] 2.73e-19
C8195 _010_ a_3597_12021# 0.217f
C8196 _133_ a_14063_7093# 4.06e-19
C8197 a_13415_2442# _115_ 0.187f
C8198 net30 a_10137_4943# 0.00632f
C8199 _090_ a_5087_3855# 6.18e-19
C8200 net3 a_4471_4007# 0.00209f
C8201 net53 a_5915_10927# 0.196f
C8202 mask\[0\] _079_ 0.111f
C8203 net44 _021_ 0.0069f
C8204 _104_ a_10329_1921# 0.00234f
C8205 net40 a_13697_4373# 1.62e-20
C8206 net19 _058_ 2.29e-20
C8207 net43 a_7256_8029# 0.0148f
C8208 net20 _020_ 2.56e-22
C8209 calibrate a_6822_4399# 4.65e-19
C8210 net19 _044_ 0.00813f
C8211 _122_ a_13257_4943# 8.3e-20
C8212 en_co_clk a_3365_4943# 0.0136f
C8213 _107_ a_6737_4719# 0.00311f
C8214 _065_ a_9889_6873# 2.68e-19
C8215 cal_itt\[0\] a_10005_6031# 0.0693f
C8216 a_9460_6807# a_9602_6941# 0.00783f
C8217 _062_ a_8935_6895# 0.0401f
C8218 clknet_2_2__leaf_clk a_11859_3689# 0.0363f
C8219 a_9003_3829# a_9004_3677# 6.19e-19
C8220 _085_ a_3511_11471# 0.00151f
C8221 net43 _018_ 0.193f
C8222 a_5547_5603# _107_ 1.04e-19
C8223 clknet_2_2__leaf_clk a_11149_2767# 0.00309f
C8224 trim_mask\[2\] a_14172_1513# 8.01e-19
C8225 a_14870_7369# VPWR 0.00127f
C8226 _095_ a_4617_4105# 8.87e-21
C8227 _111_ a_11801_4373# 2.55e-19
C8228 net31 _047_ 0.105f
C8229 mask\[2\] a_5055_9295# 4.73e-19
C8230 net4 a_3333_2601# 5.18e-19
C8231 a_15023_2767# trim[1] 0.00179f
C8232 mask\[6\] a_2787_10927# 0.132f
C8233 _107_ a_9003_3829# 0.0111f
C8234 a_14236_8457# a_14063_7093# 6.49e-20
C8235 a_11394_9509# a_11545_9049# 6.11e-20
C8236 trim_mask\[4\] a_11067_3017# 0.0102f
C8237 _129_ _135_ 7.86e-20
C8238 _031_ a_13257_1141# 0.222f
C8239 _049_ a_6737_4719# 0.00675f
C8240 net34 cal_count\[2\] 7.97e-20
C8241 net13 _060_ 0.202f
C8242 a_1763_9295# result[3] 5.04e-20
C8243 a_5536_4399# _107_ 0.112f
C8244 net9 _066_ 2.45e-20
C8245 _049_ a_5547_5603# 0.00282f
C8246 trim_mask\[0\] a_13233_4737# 0.0029f
C8247 net23 _080_ 0.299f
C8248 mask\[1\] _039_ 1.8e-20
C8249 a_15299_6575# en_co_clk 2.25e-19
C8250 net13 _022_ 1.44e-20
C8251 trim_mask\[0\] a_7891_3617# 1.5e-20
C8252 _084_ a_5915_11721# 0.0981f
C8253 cal_count\[3\] clk 1.09e-20
C8254 _112_ trim[0] 1.79e-20
C8255 en_co_clk cal_count\[3\] 0.00244f
C8256 net15 _093_ 0.00808f
C8257 _110_ a_10569_1109# 0.0625f
C8258 cal_itt\[1\] a_9693_8029# 0.00108f
C8259 a_13562_8751# VPWR 0.199f
C8260 _049_ a_9003_3829# 1.43e-19
C8261 net54 a_5537_4105# 1.18e-20
C8262 a_7223_2465# VPWR 0.449f
C8263 a_8820_12533# VPWR 0.298f
C8264 net43 mask\[1\] 0.15f
C8265 a_1835_11231# a_1679_10633# 0.00155f
C8266 a_13091_4943# _113_ 1.61e-20
C8267 a_12900_7663# _132_ 6.76e-20
C8268 a_10655_2932# trim_val\[3\] 4.87e-21
C8269 cal_count\[3\] a_9084_4515# 8.9e-19
C8270 a_1313_11989# a_1313_10901# 0.00117f
C8271 net43 a_745_10933# 0.0348f
C8272 a_745_12021# a_1095_11305# 1.97e-20
C8273 _078_ a_1764_10383# 5.45e-19
C8274 _049_ a_5536_4399# 9.78e-19
C8275 _092_ trim_mask\[4\] 2.7e-22
C8276 clknet_2_3__leaf_clk a_11059_7356# 0.00312f
C8277 a_10676_1679# a_10752_565# 2.48e-20
C8278 a_1173_6031# calibrate 3.52e-21
C8279 a_5177_1921# a_5055_1679# 3.16e-19
C8280 _136_ _108_ 0.008f
C8281 a_7263_7093# a_7088_7119# 0.234f
C8282 _074_ net25 0.123f
C8283 _133_ a_13279_7119# 0.0104f
C8284 a_561_6031# a_1476_6031# 0.125f
C8285 net53 a_4043_10143# 0.00285f
C8286 a_855_4105# VPWR 0.242f
C8287 net26 _019_ 6.44e-20
C8288 a_7999_11231# a_7824_11305# 0.234f
C8289 net9 a_11545_9049# 2.47e-19
C8290 _048_ a_3530_4438# 7.33e-19
C8291 _127_ _129_ 1.48e-19
C8292 net15 a_2865_4460# 0.00353f
C8293 a_9099_3689# VPWR 0.209f
C8294 a_11814_9295# _128_ 3.23e-20
C8295 _120_ _090_ 0.027f
C8296 net14 _074_ 0.926f
C8297 mask\[7\] _078_ 0.362f
C8298 a_11067_4405# _058_ 0.033f
C8299 net46 a_8491_2229# 0.296f
C8300 _129_ a_14063_7093# 0.12f
C8301 _110_ a_10329_1921# 1.39e-20
C8302 a_14335_4020# _112_ 1.37e-19
C8303 clknet_2_1__leaf_clk a_6419_8207# 5.61e-19
C8304 _104_ a_10975_4105# 0.226f
C8305 _065_ a_6885_8372# 0.0332f
C8306 net43 a_1387_8751# 0.0149f
C8307 net40 a_13825_5185# 3.26e-19
C8308 a_9463_8725# a_9459_7895# 2.81e-20
C8309 _046_ a_3431_10933# 7.78e-20
C8310 a_12047_2601# VPWR 2.96e-19
C8311 net50 a_11601_2229# 3.78e-20
C8312 clknet_2_2__leaf_clk a_9572_2601# 0.0234f
C8313 a_15299_3311# trim[1] 0.00392f
C8314 net15 _034_ 1.23e-19
C8315 a_10005_6031# trim_mask\[0\] 0.0047f
C8316 cal_itt\[2\] a_8307_6575# 0.0929f
C8317 net25 a_1279_9129# 3.39e-19
C8318 mask\[7\] a_2869_11247# 0.00419f
C8319 _080_ _016_ 8.64e-21
C8320 a_10781_3311# a_10676_1679# 1.11e-20
C8321 a_763_8757# VPWR 0.486f
C8322 a_8745_6895# a_8935_6895# 0.0905f
C8323 a_395_4405# a_816_4765# 0.0931f
C8324 a_8485_4943# _107_ 1.29e-19
C8325 a_10055_5487# VPWR 0.235f
C8326 a_4259_6031# a_4871_6031# 3.82e-19
C8327 a_4425_6031# a_5502_6397# 1.46e-19
C8328 _040_ a_3781_8207# 0.0404f
C8329 a_448_7637# _005_ 0.0668f
C8330 trim_mask\[4\] a_6906_2355# 0.0036f
C8331 mask\[6\] a_7259_11305# 7.79e-22
C8332 a_10016_1679# a_9719_1473# 4.67e-19
C8333 net14 a_1279_9129# 0.0113f
C8334 a_11987_8757# cal_count\[1\] 1.09e-19
C8335 _066_ a_10188_4105# 1.06e-20
C8336 net16 trimb[3] 3.69e-19
C8337 _011_ ctlp[0] 4.62e-19
C8338 net26 a_6467_9845# 0.0437f
C8339 _074_ a_395_7119# 0.0183f
C8340 cal_itt\[0\] a_10877_7983# 6.84e-20
C8341 _067_ a_9889_6873# 0.138f
C8342 trim_mask\[0\] _087_ 3.44e-21
C8343 net44 a_3521_7361# 5.86e-20
C8344 net13 a_4498_4373# 0.00856f
C8345 net13 a_4864_1679# 0.00562f
C8346 net52 a_3840_8867# 0.00329f
C8347 net46 a_12625_2601# 6.97e-19
C8348 net29 a_1579_11471# 5.38e-19
C8349 _065_ a_11141_6031# 0.0116f
C8350 a_10018_3677# VPWR 8.89e-19
C8351 _110_ a_11374_1251# 0.00108f
C8352 clknet_2_1__leaf_clk a_3303_10217# 0.0142f
C8353 _075_ _087_ 0.00266f
C8354 net26 VPWR 2.42f
C8355 net34 cal_count\[1\] 1.15e-20
C8356 trim_mask\[4\] a_9317_3285# 0.0221f
C8357 a_9478_4105# a_9099_3689# 4.32e-20
C8358 trim_mask\[0\] _099_ 8.74e-21
C8359 net52 a_2971_8457# 0.191f
C8360 net23 a_1651_7093# 0.0612f
C8361 mask\[7\] a_3597_10933# 1.79e-19
C8362 a_5050_8207# VPWR 6.24e-19
C8363 _131_ VPWR 0.563f
C8364 mask\[1\] a_2857_7637# 0.0121f
C8365 _088_ VPWR 0.704f
C8366 _092_ a_3123_3615# 4.55e-19
C8367 a_4687_12319# a_4512_12393# 0.234f
C8368 a_3947_12393# mask\[6\] 8.25e-21
C8369 a_8307_4943# a_8389_5193# 0.0961f
C8370 net19 _069_ 2.78e-20
C8371 net4 a_7800_4631# 1.04e-21
C8372 net26 a_5699_9269# 0.00125f
C8373 a_9595_1679# a_10016_1679# 0.0931f
C8374 _075_ _099_ 3.69e-19
C8375 mask\[2\] net24 0.725f
C8376 a_7262_5461# VPWR 0.327f
C8377 _122_ net40 5.85e-20
C8378 calibrate a_4617_4105# 0.0473f
C8379 _037_ a_11204_7485# 2.26e-19
C8380 a_13459_3317# a_13625_3317# 0.845f
C8381 net19 a_8022_7119# 0.0206f
C8382 _036_ a_12153_8757# 0.0549f
C8383 a_11987_8757# a_12612_8725# 0.181f
C8384 _055_ a_14686_3017# 4.96e-19
C8385 net15 a_3830_6281# 1.95e-19
C8386 net46 a_11764_3677# 6.55e-19
C8387 trim_val\[4\] VPWR 0.311f
C8388 a_4512_12393# net13 0.00232f
C8389 mask\[6\] a_3425_11721# 0.0504f
C8390 _062_ _066_ 0.0114f
C8391 _018_ a_2953_9845# 0.223f
C8392 a_2787_9845# a_3521_9813# 0.0535f
C8393 _006_ result[2] 8.61e-19
C8394 _051_ a_4709_2773# 0.0198f
C8395 net40 _063_ 4.59e-19
C8396 net14 _093_ 0.0132f
C8397 a_6737_3855# a_7104_3855# 2.15e-20
C8398 net46 a_10195_1354# 0.00127f
C8399 trim[4] trim[1] 0.0419f
C8400 net42 a_7527_4631# 7.88e-20
C8401 en_co_clk a_14347_4917# 3.21e-19
C8402 a_6519_4631# VPWR 0.236f
C8403 a_5686_2045# VPWR 6.47e-19
C8404 clknet_2_2__leaf_clk a_13825_1109# 5.11e-19
C8405 clknet_2_1__leaf_clk a_455_8181# 2.58e-19
C8406 net18 ctln[3] 2.83e-20
C8407 _051_ a_4308_4917# 3.56e-21
C8408 _081_ a_2143_7663# 1.53e-19
C8409 _123_ _037_ 0.0116f
C8410 a_6927_12559# a_6891_12393# 0.0111f
C8411 _038_ a_8298_5487# 7.24e-21
C8412 net51 clknet_0_clk 1.07e-20
C8413 _069_ cal_itt\[1\] 0.208f
C8414 trim_mask\[2\] _025_ 1.26e-19
C8415 a_1867_3317# a_2288_3677# 0.0859f
C8416 trim_mask\[4\] a_9773_3689# 9.77e-19
C8417 _119_ clk 2.39e-20
C8418 net34 _108_ 0.00839f
C8419 a_5535_8181# a_6056_8359# 5.06e-20
C8420 trim_mask\[2\] _026_ 0.0595f
C8421 net15 net4 0.384f
C8422 a_9823_6941# VPWR 0.00127f
C8423 _076_ a_8083_8181# 9.14e-20
C8424 cal_itt\[1\] a_8022_7119# 0.0143f
C8425 mask\[6\] _008_ 6.33e-21
C8426 a_579_12021# _011_ 0.167f
C8427 net29 a_561_9845# 9.97e-20
C8428 state\[2\] a_3933_2767# 7.2e-19
C8429 net52 a_2225_7983# 3.87e-21
C8430 net54 a_4471_4007# 0.00149f
C8431 a_6737_4719# trim_mask\[4\] 4.81e-21
C8432 _016_ a_1651_7093# 1.83e-20
C8433 net49 a_14193_3285# 0.0106f
C8434 net16 clkc 3e-20
C8435 a_14281_4943# VPWR 1.35e-19
C8436 net37 _058_ 3.24e-19
C8437 _026_ a_12213_2589# 3.24e-19
C8438 a_4655_10071# a_4801_9839# 0.171f
C8439 _092_ a_3530_4765# 9.49e-19
C8440 a_2953_9845# mask\[1\] 4.19e-21
C8441 net51 a_6198_8207# 1.68e-19
C8442 clknet_2_3__leaf_clk a_11016_6691# 0.002f
C8443 _041_ _129_ 0.00225f
C8444 net46 _032_ 0.0299f
C8445 _005_ a_911_7119# 0.00362f
C8446 _104_ a_7223_2465# 1.07e-19
C8447 state\[0\] a_3933_2767# 0.00282f
C8448 clknet_2_1__leaf_clk a_1019_9839# 0.0278f
C8449 a_14471_591# ctln[2] 0.16f
C8450 _128_ a_12992_8751# 0.0126f
C8451 net15 a_3303_7119# 0.00861f
C8452 _062_ a_7571_4943# 4.31e-19
C8453 a_15023_9839# trimb[1] 0.337f
C8454 a_10699_5487# a_10975_4105# 3.29e-21
C8455 net50 a_10016_1679# 7.97e-20
C8456 clknet_2_2__leaf_clk a_13307_1707# 0.00184f
C8457 a_9805_1473# VPWR 0.00228f
C8458 net27 net26 1.42e-19
C8459 net43 _041_ 5.66e-19
C8460 _075_ a_5537_4943# 1.72e-20
C8461 _060_ a_2948_3689# 1.92e-20
C8462 net1 a_995_3530# 0.11f
C8463 trim_val\[4\] a_9478_4105# 0.0098f
C8464 a_9003_3829# trim_mask\[4\] 6.28e-19
C8465 _065_ a_4091_5309# 0.122f
C8466 _010_ net43 0.015f
C8467 en_co_clk _095_ 0.648f
C8468 _135_ a_14379_6397# 0.00107f
C8469 a_13111_6031# _061_ 2.52e-20
C8470 net9 a_12056_6031# 0.00738f
C8471 _009_ a_6891_12393# 2.71e-19
C8472 clknet_0_clk _003_ 1.8e-20
C8473 a_6375_12021# a_7631_12319# 0.0435f
C8474 _110_ a_13881_2741# 0.00291f
C8475 _101_ a_5915_10927# 0.0912f
C8476 net52 a_4131_8207# 4.37e-19
C8477 net18 a_9595_5193# 1.36e-19
C8478 net51 a_7459_7663# 7.46e-20
C8479 _053_ a_10975_6031# 0.017f
C8480 a_4425_6031# a_5340_6031# 0.123f
C8481 _082_ a_1045_9545# 3.1e-19
C8482 _104_ a_9099_3689# 0.0247f
C8483 _046_ net13 7.78e-20
C8484 a_11343_3317# a_11764_3677# 0.0902f
C8485 _025_ a_11045_3631# 1.8e-19
C8486 a_10383_7093# en_co_clk 6.54e-20
C8487 _069_ _001_ 0.216f
C8488 net54 a_4970_4399# 0.00188f
C8489 net45 a_4995_7119# 0.165f
C8490 _028_ a_6703_2197# 0.00204f
C8491 _067_ a_11141_6031# 2.28e-20
C8492 net55 a_5363_4719# 0.00256f
C8493 a_8745_4943# VPWR 3.05e-19
C8494 net19 a_8657_2229# 0.0203f
C8495 _083_ a_7548_10217# 1.65e-20
C8496 net31 net49 0.00371f
C8497 _001_ a_8022_7119# 6.44e-21
C8498 a_6927_12559# ctlp[5] 5.22e-20
C8499 net13 a_5067_9661# 0.00105f
C8500 _014_ a_2288_3677# 0.00439f
C8501 net9 _058_ 0.0376f
C8502 a_13783_6183# a_13091_4943# 7.08e-21
C8503 _049_ a_4266_4943# 1.44e-19
C8504 _092_ a_11491_6031# 4.93e-21
C8505 _105_ _107_ 0.00862f
C8506 _101_ a_1467_7923# 0.00344f
C8507 cal_itt\[0\] a_10864_7387# 2.67e-20
C8508 _023_ a_1835_11231# 4.1e-20
C8509 _045_ a_5578_12131# 4.96e-19
C8510 a_579_10933# a_1660_11305# 0.102f
C8511 net2 a_12061_7669# 1.9e-19
C8512 a_8749_3317# _028_ 6.93e-20
C8513 _134_ net5 0.00203f
C8514 net18 net4 4.59e-22
C8515 a_11067_4405# a_11488_4765# 0.0894f
C8516 a_11987_8757# a_12900_7663# 4.51e-20
C8517 a_12992_8751# a_11895_7669# 2.42e-20
C8518 _036_ a_13050_7637# 7.23e-19
C8519 a_448_7637# a_395_7119# 0.0112f
C8520 _072_ net30 0.00455f
C8521 _107_ a_7010_3311# 0.00214f
C8522 cal_itt\[2\] VPWR 0.738f
C8523 mask\[3\] _018_ 0.163f
C8524 a_4512_11305# a_4621_11305# 0.00742f
C8525 a_3947_11305# a_4055_10927# 0.0572f
C8526 a_4687_11231# a_4866_11293# 0.0074f
C8527 a_7617_2589# clk 5.18e-19
C8528 _118_ a_10137_4943# 0.068f
C8529 _029_ a_13825_5185# 9.46e-20
C8530 _049_ _105_ 0.00221f
C8531 net26 a_8455_10383# 8.13e-19
C8532 trim_mask\[0\] a_14972_5193# 0.102f
C8533 _068_ net30 0.00285f
C8534 net33 net36 0.157f
C8535 a_14604_2339# a_14172_1513# 2.85e-20
C8536 a_14347_9480# a_14467_8751# 6.34e-20
C8537 _040_ a_4393_8207# 0.00258f
C8538 _051_ _090_ 0.202f
C8539 _088_ _104_ 0.102f
C8540 mask\[5\] a_8154_11721# 9.54e-19
C8541 _061_ a_13825_6031# 2.07e-19
C8542 a_11587_6031# _136_ 9.98e-19
C8543 _069_ a_7916_8041# 3.66e-20
C8544 _078_ _080_ 0.0018f
C8545 _049_ a_7010_3311# 0.11f
C8546 a_7262_5461# _104_ 6.3e-22
C8547 _090_ _014_ 0.00256f
C8548 net44 a_8215_9295# 0.00597f
C8549 net14 net4 1.54e-19
C8550 net43 _002_ 0.311f
C8551 _101_ a_4043_10143# 0.0616f
C8552 clknet_0_clk a_7223_2465# 0.0133f
C8553 trim_mask\[4\] trim_val\[3\] 3.15e-20
C8554 trim_mask\[1\] a_13880_3677# 4.06e-19
C8555 a_7916_8041# a_8022_7119# 0.00789f
C8556 trim_mask\[2\] _031_ 0.12f
C8557 _071_ a_7088_7119# 1.73e-20
C8558 cal_count\[3\] _108_ 0.00102f
C8559 a_4609_9295# a_5055_9295# 2.28e-19
C8560 a_5177_9537# a_5686_9661# 2.6e-19
C8561 _014_ a_3847_4438# 1.51e-20
C8562 net52 net30 1.74e-20
C8563 clknet_2_1__leaf_clk a_579_12021# 0.395f
C8564 net47 a_9458_9661# 1.81e-19
C8565 net46 net30 3.76e-21
C8566 _127_ cal_count\[0\] 0.286f
C8567 net43 _050_ 1.75e-20
C8568 _104_ trim_val\[4\] 0.0488f
C8569 net12 _103_ 8.81e-21
C8570 trim_val\[1\] a_14184_2767# 1.99e-19
C8571 a_3529_6281# _092_ 3.9e-19
C8572 _095_ _059_ 7.45e-19
C8573 _071_ _063_ 0.0685f
C8574 _073_ _049_ 6.44e-20
C8575 mask\[3\] mask\[1\] 9.14e-20
C8576 net40 comp 2.43e-19
C8577 net3 net1 8.1e-20
C8578 net45 a_3224_2601# 0.245f
C8579 _058_ a_10188_4105# 0.107f
C8580 a_15159_9269# net2 5.47e-21
C8581 net19 a_10569_1109# 2.46e-21
C8582 net15 ctln[1] 0.00218f
C8583 _027_ _117_ 1.84e-20
C8584 a_2309_2229# net7 1.8e-20
C8585 a_15023_2223# a_15023_1679# 0.00817f
C8586 net18 a_11479_9117# 2.47e-19
C8587 a_3840_8867# _065_ 8.62e-20
C8588 clknet_2_3__leaf_clk a_11709_6273# 0.0701f
C8589 _074_ a_4165_11989# 2.01e-20
C8590 _110_ a_9099_3689# 0.00179f
C8591 _015_ a_4617_4105# 0.00189f
C8592 a_2953_7119# a_4995_7119# 1.05e-19
C8593 a_3303_7119# a_3399_7119# 0.0138f
C8594 a_3521_7361# a_3565_7119# 3.69e-19
C8595 a_395_9845# a_448_9269# 0.0112f
C8596 net22 a_3748_6281# 1.48e-20
C8597 a_745_10933# mask\[3\] 2.68e-20
C8598 _048_ a_8473_5193# 0.0224f
C8599 mask\[7\] a_3852_12381# 4.96e-21
C8600 _050_ a_7010_3631# 1.85e-20
C8601 clknet_2_1__leaf_clk a_2869_10927# 1.3e-19
C8602 _039_ a_561_6031# 0.00143f
C8603 net33 _128_ 0.00162f
C8604 _074_ _019_ 7.53e-20
C8605 mask\[7\] a_1651_10143# 0.00273f
C8606 net14 a_911_7119# 0.00542f
C8607 trim_mask\[2\] a_10781_3311# 0.00203f
C8608 a_1173_4765# cal 4.66e-20
C8609 net26 a_8381_9295# 4.16e-20
C8610 _006_ _040_ 1e-19
C8611 net50 _025_ 9.84e-20
C8612 a_7939_3855# _028_ 4.32e-20
C8613 net9 a_13607_4943# 5.4e-20
C8614 _101_ a_2787_7119# 6.81e-20
C8615 net43 a_561_6031# 2.76e-19
C8616 net14 a_1835_12319# 0.00117f
C8617 a_2971_8457# net23 5.34e-20
C8618 net25 a_2450_9955# 2.14e-19
C8619 _090_ a_5445_4399# 0.00164f
C8620 a_11297_7119# VPWR 1.82e-19
C8621 calibrate clk 6.08e-20
C8622 en_co_clk calibrate 0.00117f
C8623 a_11244_9661# _122_ 0.0012f
C8624 _052_ a_7010_3631# 0.00318f
C8625 net49 a_14083_3311# 0.00301f
C8626 net43 a_3615_8207# 2.28e-20
C8627 a_13512_4943# a_13703_4943# 4.61e-19
C8628 a_14172_4943# trim_val\[0\] 0.0019f
C8629 _058_ trim_mask\[3\] 4.79e-21
C8630 a_3431_12021# a_5496_12131# 3.73e-21
C8631 _134_ a_15023_6031# 3.59e-21
C8632 net8 a_14471_591# 0.17f
C8633 _122_ a_11204_7485# 0.00442f
C8634 a_929_8757# net45 2.05e-19
C8635 a_5081_4943# VPWR 0.00571f
C8636 net13 a_4576_3427# 0.00304f
C8637 a_6743_10933# a_7367_10927# 9.73e-19
C8638 net16 clknet_2_3__leaf_clk 0.016f
C8639 net18 a_10586_7371# 6.42e-19
C8640 net51 a_6523_7119# 1.5e-19
C8641 a_10586_7371# a_10820_7485# 0.00645f
C8642 a_395_7119# a_911_7119# 0.115f
C8643 clknet_2_1__leaf_clk net53 0.87f
C8644 net34 trimb[2] 0.0773f
C8645 a_4858_8573# VPWR 5.58e-19
C8646 trim_mask\[0\] a_9503_4399# 5.26e-21
C8647 net55 VPWR 1.78f
C8648 _110_ a_10018_3677# 2.04e-19
C8649 _049_ a_3365_4943# 8.9e-20
C8650 net31 a_15159_9269# 0.00589f
C8651 _120_ a_3667_3829# 5.12e-20
C8652 a_3365_4943# a_3388_4631# 9.7e-19
C8653 net15 a_3057_4719# 0.00587f
C8654 _036_ VPWR 0.975f
C8655 net29 result[7] 0.00528f
C8656 _078_ a_1677_9545# 0.0784f
C8657 _134_ net46 6.57e-20
C8658 _101_ a_3208_10205# 0.0198f
C8659 _101_ a_2689_8751# 0.00483f
C8660 _122_ a_13349_6031# 9.84e-21
C8661 _123_ _122_ 0.941f
C8662 clknet_2_0__leaf_clk a_1638_4399# 1.67e-19
C8663 net4 a_2659_2601# 3.81e-19
C8664 _094_ _060_ 1.56e-20
C8665 result[0] sample 0.0473f
C8666 cal_count\[3\] _107_ 0.00455f
C8667 _074_ VPWR 3.7f
C8668 trim_mask\[0\] a_9369_3855# 3.36e-19
C8669 net40 a_13111_6031# 0.00196f
C8670 clknet_0_clk _088_ 5.9e-20
C8671 net44 a_7256_8029# 0.00192f
C8672 net47 a_12454_8041# 1.54e-19
C8673 a_9595_1679# a_10752_565# 3.61e-19
C8674 _078_ a_1651_7093# 0.00166f
C8675 clknet_0_clk a_7262_5461# 0.0512f
C8676 trim_val\[2\] a_13257_1141# 4.18e-19
C8677 _123_ _063_ 0.0556f
C8678 net20 a_7109_11989# 0.0042f
C8679 a_6007_7119# a_7263_7093# 0.0436f
C8680 _003_ a_6523_7119# 3.12e-19
C8681 net33 _056_ 0.0733f
C8682 a_3431_10933# a_3868_10217# 8.37e-21
C8683 a_14099_1929# a_13607_1513# 1.49e-19
C8684 net8 a_13825_1109# 0.00805f
C8685 net23 a_2225_7983# 0.00378f
C8686 _110_ trim_val\[4\] 0.0123f
C8687 _074_ a_5699_9269# 0.00292f
C8688 a_6743_10933# a_7999_11231# 0.0436f
C8689 _021_ a_7259_11305# 5.07e-19
C8690 a_7715_3285# VPWR 0.166f
C8691 en_co_clk a_8298_5487# 6.9e-19
C8692 net46 a_13975_3689# 0.174f
C8693 net12 a_6261_11247# 0.00129f
C8694 _130_ a_15023_5487# 0.00105f
C8695 _049_ cal_count\[3\] 5.13e-20
C8696 a_7939_10383# a_7723_10143# 9.27e-19
C8697 a_10975_4105# a_11057_4105# 0.171f
C8698 _052_ a_6822_4399# 0.00147f
C8699 net4 a_10055_2767# 0.208f
C8700 a_1279_9129# VPWR 0.195f
C8701 a_911_4777# a_816_4765# 0.0498f
C8702 _065_ a_4131_8207# 8.11e-20
C8703 a_14702_3311# VPWR 7.19e-19
C8704 a_8298_5487# a_9084_4515# 9.54e-19
C8705 a_5423_9011# _076_ 3.4e-20
C8706 _065_ a_6793_8970# 3.73e-19
C8707 a_13693_3883# VPWR 0.00207f
C8708 clknet_2_2__leaf_clk a_8491_2229# 0.514f
C8709 _012_ a_1651_4703# 4.1e-20
C8710 a_9802_4007# _119_ 3.79e-19
C8711 _002_ a_8270_8029# 7.49e-19
C8712 mask\[7\] a_1191_11305# 1.47e-19
C8713 _057_ net10 8.16e-19
C8714 net45 a_5524_1679# 0.242f
C8715 cal_count\[0\] _041_ 0.419f
C8716 net46 a_13915_4399# 3.28e-19
C8717 a_14347_9480# a_14249_8725# 6.66e-19
C8718 a_13279_8207# a_13470_7663# 6.57e-19
C8719 _040_ _017_ 0.0831f
C8720 net28 a_5496_12131# 0.105f
C8721 a_7263_7093# _092_ 1.19e-19
C8722 a_13881_1653# a_14099_1929# 0.0821f
C8723 a_13307_1707# net8 7.89e-20
C8724 ctlp[4] ctlp[3] 0.00165f
C8725 a_3615_8207# a_2857_7637# 0.013f
C8726 net1 valid 0.0364f
C8727 net53 a_7245_10205# 2.96e-19
C8728 _108_ _119_ 0.00869f
C8729 net44 a_7902_10205# 0.00222f
C8730 net44 mask\[1\] 0.145f
C8731 trim_mask\[0\] _111_ 0.226f
C8732 clknet_2_3__leaf_clk a_10593_9295# 0.0159f
C8733 _059_ calibrate 0.0092f
C8734 a_14981_4020# _055_ 1.54e-20
C8735 net33 net35 0.415f
C8736 net9 _113_ 3.21e-20
C8737 _063_ a_9043_6031# 0.00116f
C8738 _042_ a_8563_10749# 0.0262f
C8739 _048_ a_7190_3855# 2.47e-19
C8740 clknet_2_0__leaf_clk net45 0.854f
C8741 _110_ a_9805_1473# 0.00165f
C8742 a_8072_11721# a_7824_11305# 4.78e-20
C8743 a_12061_7669# a_12249_7663# 0.157f
C8744 _044_ a_7999_11231# 5.4e-19
C8745 a_8673_10625# a_9182_10749# 2.6e-19
C8746 a_8105_10383# a_8551_10383# 2.28e-19
C8747 net50 a_10752_565# 0.00167f
C8748 a_8949_9537# _035_ 7.91e-22
C8749 trim_mask\[4\] a_7010_3311# 0.0854f
C8750 _038_ a_10781_5487# 0.0017f
C8751 a_8992_9955# a_8215_9295# 5.08e-21
C8752 a_855_4105# net41 2.45e-20
C8753 _060_ a_4617_3855# 0.0045f
C8754 _119_ a_10655_2932# 0.207f
C8755 _053_ a_7800_4631# 8.89e-20
C8756 en_co_clk _135_ 0.00293f
C8757 _074_ net27 0.119f
C8758 _093_ VPWR 1.07f
C8759 net30 a_7527_4631# 1.72e-20
C8760 trim_val\[2\] a_14526_1501# 6.42e-19
C8761 _094_ a_4498_4373# 1.95e-21
C8762 mask\[3\] _041_ 8.1e-20
C8763 _122_ a_13142_8725# 2.09e-19
C8764 net32 a_14237_3677# 6.64e-20
C8765 a_7263_7093# cal_itt\[3\] 0.0644f
C8766 net8 a_13715_1135# 0.00203f
C8767 a_5166_5193# VPWR 0.00496f
C8768 a_8636_9295# VPWR 0.0834f
C8769 a_12077_3285# _030_ 7.31e-20
C8770 a_12599_3615# a_13183_3311# 2.79e-19
C8771 _042_ a_3565_10205# 2.51e-19
C8772 _136_ a_12723_4943# 0.0029f
C8773 net47 a_13016_9117# 7.28e-19
C8774 net13 net45 0.226f
C8775 mask\[0\] a_1830_6031# 3.18e-19
C8776 _004_ a_816_6031# 0.16f
C8777 net28 result[7] 0.11f
C8778 a_395_6031# a_1019_6397# 9.73e-19
C8779 a_5515_6005# net3 6.01e-19
C8780 net50 a_10781_3311# 0.00363f
C8781 net46 a_11030_1679# 0.00414f
C8782 clknet_2_2__leaf_clk a_11764_3677# 0.0164f
C8783 _040_ a_4425_6031# 4.4e-20
C8784 clknet_2_1__leaf_clk a_6007_9839# 5.24e-19
C8785 a_5177_9537# a_5633_9295# 4.2e-19
C8786 a_2865_4460# VPWR 0.151f
C8787 a_7351_8041# a_7447_8041# 0.0138f
C8788 net44 a_6796_12381# 5.97e-19
C8789 _065_ net30 0.634f
C8790 a_7109_11989# a_6987_12393# 3.16e-19
C8791 net4 a_4959_1679# 1.8e-20
C8792 net34 net36 0.206f
C8793 net38 net33 0.126f
C8794 _119_ a_9004_3677# 0.0083f
C8795 a_6703_2197# ctln[6] 1.83e-21
C8796 a_3781_8207# _077_ 0.00176f
C8797 net33 _061_ 0.0164f
C8798 a_4131_8207# a_4696_8207# 7.99e-20
C8799 _076_ a_4871_8181# 5.33e-20
C8800 _034_ VPWR 0.596f
C8801 _108_ a_11679_4777# 3.69e-19
C8802 net40 _092_ 1.05e-19
C8803 a_3339_2767# a_2143_2229# 9.76e-20
C8804 a_3521_7361# _049_ 9.8e-19
C8805 _015_ clk 0.0298f
C8806 _095_ a_4725_5487# 5.38e-19
C8807 _063_ a_8749_3317# 1.36e-19
C8808 VPWR ctln[3] 0.189f
C8809 net55 _104_ 0.0665f
C8810 en_co_clk _015_ 6.27e-19
C8811 net21 a_5496_12131# 0.00231f
C8812 _112_ a_13625_3317# 0.0105f
C8813 _107_ _119_ 0.0048f
C8814 _072_ a_5691_7637# 4.08e-21
C8815 cal_itt\[2\] clknet_0_clk 0.186f
C8816 net15 a_2815_9447# 0.00809f
C8817 a_8022_7119# _062_ 0.00163f
C8818 a_7631_12319# a_7456_12393# 0.234f
C8819 _011_ _086_ 0.184f
C8820 mask\[4\] a_7548_10217# 0.0402f
C8821 net40 a_14199_7369# 0.00128f
C8822 a_2283_4020# a_2033_3317# 2.94e-19
C8823 a_3224_2601# a_3386_2223# 0.00645f
C8824 net18 mask\[4\] 0.00596f
C8825 net43 a_4227_8207# 5.05e-20
C8826 a_11491_6031# _136_ 0.0067f
C8827 net47 a_10990_7485# 0.166f
C8828 _048_ a_5625_4943# 0.00231f
C8829 a_15023_8751# trimb[4] 0.337f
C8830 a_14237_3677# VPWR 4.56e-19
C8831 _100_ a_5931_4105# 0.0509f
C8832 _088_ net41 1.32e-20
C8833 net16 a_14099_1929# 0.00392f
C8834 _001_ a_13142_7271# 9.76e-20
C8835 _128_ a_11987_8757# 6.99e-19
C8836 net13 a_3868_10217# 0.00106f
C8837 net18 _064_ 0.0288f
C8838 a_2948_3689# a_4576_3427# 3.02e-20
C8839 a_9503_4399# a_8298_2767# 5.39e-21
C8840 clknet_2_2__leaf_clk _032_ 0.0022f
C8841 a_11067_4405# a_10975_4105# 5.24e-19
C8842 clknet_2_0__leaf_clk a_2953_7119# 0.606f
C8843 a_4425_6031# _048_ 1.59e-20
C8844 a_448_7637# VPWR 0.252f
C8845 en_co_clk a_14649_6031# 6.97e-19
C8846 _051_ _106_ 5.03e-19
C8847 net12 a_6885_8372# -2.1e-36
C8848 _049_ _119_ 1.08e-19
C8849 clknet_2_3__leaf_clk clkc 1.48e-19
C8850 net29 mask\[7\] 1.16f
C8851 a_7190_3855# a_7021_4105# 0.0821f
C8852 a_6566_5193# _107_ 5.69e-19
C8853 _136_ net35 4.2e-19
C8854 _136_ a_13059_4631# 7.02e-19
C8855 _041_ a_13919_8751# 0.207f
C8856 net52 a_5691_7637# 0.306f
C8857 a_12992_8751# net40 2.31e-19
C8858 net46 a_15054_5193# 1.6e-19
C8859 _096_ _060_ 0.0589f
C8860 net18 a_10851_1653# 0.00776f
C8861 a_10043_7983# VPWR 9.94e-19
C8862 net46 trim_val\[1\] 0.0319f
C8863 a_9595_5193# VPWR 0.459f
C8864 _010_ a_3513_12809# 0.0124f
C8865 a_8820_12533# net19 0.172f
C8866 net19 a_7223_2465# 0.00294f
C8867 _083_ a_6467_9845# 0.0291f
C8868 a_13091_4943# a_14281_4943# 2.56e-19
C8869 a_5363_12559# ctlp[6] 4.08e-19
C8870 a_9020_10383# _043_ 0.00275f
C8871 net15 _081_ 4.63e-20
C8872 mask\[4\] a_9129_10383# 5.2e-19
C8873 cal_count\[2\] _135_ 7.17e-20
C8874 _016_ net30 1.45e-19
C8875 cal_count\[3\] trim_mask\[4\] 1.55e-20
C8876 _024_ a_11067_3017# 8.17e-20
C8877 _084_ a_6181_10633# 5e-20
C8878 a_8105_10383# a_9871_10383# 1.52e-19
C8879 _049_ a_6566_5193# 0.0076f
C8880 net43 a_2019_9055# 0.271f
C8881 a_7939_10383# _042_ 0.05f
C8882 state\[2\] a_7527_4631# 4.33e-19
C8883 a_10864_9269# _053_ 9.89e-22
C8884 a_3830_6281# VPWR 0.00193f
C8885 net13 a_2953_7119# 1.73e-20
C8886 _049_ _095_ 0.0214f
C8887 a_1660_12393# a_3597_12021# 7.01e-21
C8888 net45 a_561_7119# 9.57e-19
C8889 mask\[7\] a_3431_12021# 6.7e-19
C8890 _083_ VPWR 0.172f
C8891 net18 _053_ 0.829f
C8892 a_2857_5461# a_3817_4697# 0.00244f
C8893 _095_ a_3388_4631# 0.00196f
C8894 a_14972_5193# a_15083_4659# 0.00593f
C8895 a_7010_3311# a_7320_3631# 0.0114f
C8896 _078_ a_3840_8867# 0.0426f
C8897 state\[2\] state\[1\] 0.204f
C8898 net19 a_9099_3689# 0.00765f
C8899 _051_ _033_ 4.8e-20
C8900 clknet_2_1__leaf_clk _101_ 1.01f
C8901 trim_mask\[3\] a_8657_2229# 1.89e-19
C8902 a_8298_2767# a_9747_2527# 0.0109f
C8903 net46 _118_ 6.17e-20
C8904 a_11987_8757# a_11895_7669# 3.88e-20
C8905 a_15023_5487# trim[4] 0.337f
C8906 _083_ a_5699_9269# 4.82e-19
C8907 state\[0\] state\[1\] 0.215f
C8908 _093_ a_2383_3689# 5.04e-20
C8909 a_3431_10933# a_4621_11305# 2.56e-19
C8910 net44 _041_ 0.0236f
C8911 _125_ a_14377_7983# 1.08e-20
C8912 clknet_2_0__leaf_clk a_2857_5461# 1.83f
C8913 net4 VPWR 4.24f
C8914 a_9225_2197# a_9115_2223# 0.0977f
C8915 net52 a_4775_6031# 3.49e-21
C8916 net13 a_4905_3855# 0.00167f
C8917 net55 _110_ 8.54e-21
C8918 _074_ a_1007_4777# 0.00164f
C8919 a_3365_4943# a_3123_3615# 1.96e-20
C8920 net13 a_3922_8867# 5.75e-20
C8921 clknet_0_clk net55 0.344f
C8922 a_8022_7119# a_8745_6895# 0.00282f
C8923 _126_ trimb[4] 0.00797f
C8924 _065_ state\[0\] 2.46e-21
C8925 a_13111_6031# a_13349_6031# 0.0175f
C8926 _061_ _136_ 0.00202f
C8927 _123_ a_13111_6031# 7.17e-20
C8928 net3 a_2143_2229# 1.33e-19
C8929 net34 _056_ 0.0887f
C8930 a_3303_7119# VPWR 0.223f
C8931 state\[2\] a_5054_4399# 2.02e-19
C8932 a_6891_12393# _021_ 2.75e-20
C8933 a_8360_10383# VPWR 0.0807f
C8934 cal_count\[2\] a_14063_7093# 0.0799f
C8935 a_7631_12319# a_6743_10933# 1.2e-19
C8936 _063_ a_8935_6895# 0.0339f
C8937 _043_ a_8731_9295# 7.66e-19
C8938 a_1651_10143# a_1677_9545# 0.00123f
C8939 _060_ a_5455_4943# 0.127f
C8940 _071_ a_6007_7119# 1.97e-21
C8941 trim_val\[4\] a_11057_4105# 9.23e-20
C8942 _007_ a_1045_9545# 0.0154f
C8943 trim_mask\[0\] a_14981_4020# 0.00115f
C8944 a_11244_9661# a_11814_9295# 0.111f
C8945 net9 a_13783_6183# 4.82e-20
C8946 clknet_2_1__leaf_clk _086_ 0.00107f
C8947 a_911_7119# VPWR 0.23f
C8948 a_7184_2339# clk 0.0195f
C8949 a_14172_4943# VPWR 0.292f
C8950 a_1313_10901# net25 1.58e-19
C8951 _009_ net53 1.32e-20
C8952 net19 net26 0.0105f
C8953 a_10543_2455# a_11601_2229# 3.28e-19
C8954 a_1095_11305# a_1476_10217# 1.16e-20
C8955 a_1835_11231# a_1651_10143# 1.51e-20
C8956 net9 a_11374_1251# 6.58e-20
C8957 net30 clknet_2_2__leaf_clk 0.00237f
C8958 _096_ a_4498_4373# 0.0796f
C8959 net40 a_14422_7093# 0.00526f
C8960 a_1835_12319# VPWR 0.408f
C8961 a_15023_8751# _130_ 5.69e-21
C8962 _136_ a_13257_4943# 0.00381f
C8963 _048_ _103_ 0.481f
C8964 a_1099_12533# a_1095_11305# 1.43e-20
C8965 net14 a_1313_10901# 0.00502f
C8966 net3 a_4815_3031# 5.43e-20
C8967 clknet_0_clk a_7715_3285# 2.23e-19
C8968 net52 a_3411_7485# 3.39e-19
C8969 a_1651_7093# a_1830_7119# 0.0074f
C8970 clknet_2_1__leaf_clk _102_ 1.34e-19
C8971 a_6909_10933# a_7939_10383# 0.00123f
C8972 a_579_10933# a_395_9845# 9.43e-22
C8973 a_1476_7119# a_1585_7119# 0.00742f
C8974 net12 net42 2.81e-20
C8975 a_2450_9955# VPWR 0.00131f
C8976 a_11479_9117# VPWR 6.47e-20
C8977 net4 a_9478_4105# 0.00404f
C8978 a_1844_9129# a_2143_7663# 3.74e-22
C8979 net28 mask\[7\] 0.0586f
C8980 _110_ a_13693_3883# 0.00123f
C8981 net27 _083_ 2.92e-21
C8982 _064_ a_11023_5108# 0.00294f
C8983 a_8298_5487# _108_ 1.24e-19
C8984 clknet_2_0__leaf_clk a_3386_2223# 6.2e-19
C8985 _040_ _121_ 2.96e-20
C8986 trim_mask\[2\] trim_val\[2\] 0.319f
C8987 _071_ _092_ 0.0264f
C8988 net45 a_2948_3689# 0.236f
C8989 a_1493_5487# a_561_4405# 3.16e-20
C8990 a_11814_9295# _123_ 4.3e-20
C8991 cal_count\[0\] a_10747_8970# 4.82e-19
C8992 net34 net35 0.00132f
C8993 a_561_7119# a_2953_7119# 0.00148f
C8994 _051_ _054_ 0.0162f
C8995 _100_ state\[1\] 0.0265f
C8996 net40 _132_ 0.201f
C8997 trim_mask\[3\] a_10569_1109# 0.062f
C8998 mask\[2\] a_2961_9545# 0.00166f
C8999 a_10239_9295# _122_ 0.00155f
C9000 a_4512_11305# net26 7.08e-20
C9001 cal_itt\[0\] _070_ 0.00994f
C9002 _078_ a_395_6031# 0.00861f
C9003 net14 _081_ 0.0112f
C9004 net33 net40 0.994f
C9005 _078_ a_4131_8207# 7.94e-20
C9006 a_6763_5193# VPWR 0.274f
C9007 a_8381_9295# a_8636_9295# 0.0612f
C9008 a_8949_9537# a_9296_9295# 0.0512f
C9009 _078_ a_6793_8970# 9.27e-20
C9010 net48 _114_ 0.00155f
C9011 calibrate _107_ 0.0534f
C9012 _064_ a_10055_2767# 0.00164f
C9013 a_5535_8181# net2 9.21e-20
C9014 _102_ a_2368_9955# 1.65e-19
C9015 net44 _002_ 0.0123f
C9016 net9 a_13142_7271# 0.00188f
C9017 clknet_2_1__leaf_clk _022_ 0.144f
C9018 mask\[2\] mask\[0\] 1.12e-19
C9019 clknet_2_1__leaf_clk a_6375_12021# 0.303f
C9020 a_9889_6873# _091_ 0.00583f
C9021 a_13349_6031# a_13825_6031# 0.00178f
C9022 net44 _050_ 4.63e-19
C9023 a_9460_6807# a_8298_5487# 1.49e-19
C9024 a_10586_7371# VPWR 0.307f
C9025 a_11509_3317# VPWR 0.269f
C9026 _101_ a_1953_9129# 9.27e-21
C9027 _071_ cal_itt\[3\] 1.65e-19
C9028 a_14099_3017# VPWR 0.237f
C9029 net16 a_14334_5309# 1.39e-19
C9030 a_14733_9545# trimb[1] 2.67e-19
C9031 _119_ trim_mask\[4\] 0.00837f
C9032 trim_mask\[3\] a_10329_1921# 5.63e-20
C9033 cal_count\[2\] a_13279_7119# 0.072f
C9034 a_15023_12015# a_15023_10927# 0.00249f
C9035 _053_ a_11023_5108# 1.3e-19
C9036 _049_ calibrate 0.236f
C9037 net9 a_14181_6031# 9.57e-21
C9038 _121_ _048_ 1.12e-20
C9039 net45 _028_ 0.0288f
C9040 clknet_0_clk _093_ 3.8e-20
C9041 _127_ cal_count\[1\] 1.22e-19
C9042 _078_ a_5998_11471# 1.28e-19
C9043 mask\[6\] a_2869_10927# 0.00335f
C9044 a_8657_2229# net11 3.59e-19
C9045 cal_count\[3\] a_12723_4943# 2.44e-19
C9046 _027_ _116_ 1.29e-20
C9047 a_12691_2527# a_13091_1141# 1.95e-20
C9048 _002_ clk 5.38e-20
C9049 a_9084_4515# a_9207_3311# 4.89e-21
C9050 cal_count\[1\] a_14063_7093# 1.12e-20
C9051 a_3431_10933# a_2787_9845# 1.3e-21
C9052 a_5363_7369# a_6007_7119# 0.0129f
C9053 a_4995_7119# _003_ 1.15e-19
C9054 _114_ a_13091_1141# 8.99e-20
C9055 net3 a_5087_3855# 1.92e-20
C9056 net34 net38 0.481f
C9057 a_9166_4515# VPWR 0.00152f
C9058 a_5915_10927# a_6743_10933# 1.46e-20
C9059 cal_itt\[1\] a_9823_6941# 9.57e-19
C9060 _050_ clk 0.0344f
C9061 en_co_clk _050_ 0.112f
C9062 net34 _061_ 6.04e-19
C9063 net46 a_12424_3689# 0.262f
C9064 net13 a_4621_11305# 1.36e-19
C9065 a_11895_7669# cal_count\[3\] 1.3e-20
C9066 _037_ a_12056_6031# 2.26e-19
C9067 VPWR ctln[1] 0.176f
C9068 a_1095_11305# a_1357_11293# 0.00171f
C9069 a_1313_10901# a_1769_11305# 4.2e-19
C9070 _074_ a_1007_7119# 0.00194f
C9071 net43 a_4259_6031# 5.87e-20
C9072 a_395_7119# a_455_5747# 3.05e-21
C9073 net44 a_3615_8207# 0.296f
C9074 clknet_2_1__leaf_clk a_6515_8534# 3.1e-19
C9075 clknet_2_2__leaf_clk a_13975_3689# 4.83e-20
C9076 a_8298_5487# _107_ 0.0141f
C9077 _101_ a_6007_7119# 0.01f
C9078 a_7689_2589# VPWR 1.22e-19
C9079 _051_ a_5731_4943# 7.24e-19
C9080 clknet_2_2__leaf_clk state\[2\] 2.67e-22
C9081 net15 a_3530_4438# 1.97e-19
C9082 _065_ a_5691_7637# 6.42e-19
C9083 mask\[6\] net53 0.0795f
C9084 net4 _104_ 0.166f
C9085 _053_ a_7460_5807# 1.22e-19
C9086 _133_ a_10864_7387# 0.0012f
C9087 _052_ clk 0.0283f
C9088 net55 net41 9.56e-19
C9089 a_14335_7895# comp 1.17e-19
C9090 net45 a_1585_4777# 6.03e-19
C9091 _110_ ctln[3] 1.44e-20
C9092 net47 _068_ 3.15e-19
C9093 net46 a_12502_4765# 0.00407f
C9094 a_10688_9295# _041_ 3.12e-19
C9095 clknet_0_clk _034_ 0.127f
C9096 _042_ a_1045_9545# 4.64e-22
C9097 a_12231_6005# a_12056_6031# 0.234f
C9098 a_11491_6031# cal_count\[3\] 0.0299f
C9099 a_3053_8457# a_2857_7637# 2.46e-19
C9100 _098_ clk 3.92e-19
C9101 _078_ net30 0.0868f
C9102 _015_ a_3399_2527# 9.37e-19
C9103 _006_ a_1019_7485# 1.65e-21
C9104 a_745_10933# a_2787_10927# 5.49e-20
C9105 a_8455_10383# a_8360_10383# 0.0498f
C9106 a_9602_6614# en_co_clk 0.0029f
C9107 trim_mask\[0\] trim_mask\[2\] 2.63e-20
C9108 clknet_2_1__leaf_clk a_7824_11305# 0.00114f
C9109 _074_ net41 2.02e-19
C9110 _053_ a_6927_3311# 0.00772f
C9111 net46 a_9103_2601# 1.79e-19
C9112 net46 a_11321_3855# 5.19e-20
C9113 _108_ a_13519_4007# 1.9e-19
C9114 a_9007_2601# VPWR 0.21f
C9115 state\[0\] _013_ 7.07e-20
C9116 a_4055_10927# VPWR 0.144f
C9117 net19 cal_itt\[2\] 9.46e-19
C9118 net43 a_4043_7093# 0.313f
C9119 a_13512_4943# _112_ 1.93e-19
C9120 _068_ a_8820_6005# 4.85e-19
C9121 net14 result[5] 8.01e-20
C9122 a_13880_3677# a_14071_3689# 4.61e-19
C9123 a_12231_6005# _058_ 1.27e-20
C9124 net40 _136_ 0.0317f
C9125 a_8495_6895# a_8298_5487# 3.87e-20
C9126 a_3057_4719# VPWR 0.00555f
C9127 _123_ a_12992_8751# 0.0695f
C9128 net18 a_9664_3689# 1.3e-20
C9129 _002_ a_8091_7967# 0.00336f
C9130 a_1467_7923# net45 0.275f
C9131 a_9043_6031# _092_ 0.00324f
C9132 _122_ a_11545_9049# 0.039f
C9133 a_1497_8725# a_2006_8751# 2.6e-19
C9134 _065_ a_4775_6031# 1.69e-19
C9135 a_1129_6273# a_1638_6397# 2.6e-19
C9136 a_911_6031# a_1019_6397# 0.0572f
C9137 trim_mask\[4\] a_7617_2589# 1.36e-19
C9138 a_13607_1513# a_14172_1513# 7.99e-20
C9139 _117_ _116_ 0.224f
C9140 a_9595_5193# _110_ 4.33e-20
C9141 a_11343_3317# a_12424_3689# 0.102f
C9142 trim_mask\[1\] a_11067_3017# 2.65e-19
C9143 a_10975_4105# trim_mask\[3\] 3.89e-20
C9144 _025_ a_12599_3615# 6.78e-21
C9145 _000_ VPWR 0.473f
C9146 _048_ a_3273_4943# 0.017f
C9147 net26 a_5829_9839# 1.97e-19
C9148 a_1313_11989# mask\[7\] 2.25e-19
C9149 net43 a_1660_12393# 0.242f
C9150 clknet_2_1__leaf_clk a_4512_12393# 0.0614f
C9151 net18 a_10689_2223# 5.32e-19
C9152 _075_ _090_ 6.42e-21
C9153 net51 _062_ 7.83e-21
C9154 _026_ a_11413_2767# 2.43e-19
C9155 mask\[4\] _019_ 0.00537f
C9156 a_10005_6031# _038_ 1.62e-19
C9157 _091_ a_11141_6031# 2.12e-20
C9158 a_763_8757# a_1375_9129# 0.00188f
C9159 net46 a_11435_2229# 0.308f
C9160 a_13697_4373# _058_ 0.0124f
C9161 net16 net49 0.433f
C9162 _120_ net3 2.04e-19
C9163 net18 a_11425_5487# 6.37e-19
C9164 _095_ a_3123_3615# 4.44e-20
C9165 cal_itt\[2\] cal_itt\[1\] 0.0472f
C9166 _108_ a_14604_3017# 0.0102f
C9167 net43 a_3565_10205# 0.00401f
C9168 mask\[5\] a_7939_10383# 9.28e-19
C9169 net48 VPWR 0.412f
C9170 net16 a_14733_9545# 7.79e-19
C9171 _063_ a_7571_4943# 1.25e-20
C9172 a_395_6031# _004_ 0.17f
C9173 _050_ _059_ 0.239f
C9174 net15 a_3781_8207# 1.55e-19
C9175 a_15159_9269# trimb[1] 0.00504f
C9176 a_8072_11721# _044_ 0.109f
C9177 _103_ a_7758_4759# 1.66e-19
C9178 a_6763_5193# _104_ 1.47e-22
C9179 a_4167_6575# a_2857_5461# 3.13e-21
C9180 net45 _094_ 1.73e-20
C9181 _041_ cal_count\[1\] 0.0426f
C9182 a_4815_3031# a_4973_2773# 0.0026f
C9183 net4 _110_ 0.326f
C9184 a_1651_7093# a_1651_6005# 5.14e-19
C9185 mask\[5\] a_5997_11247# 0.00214f
C9186 a_7263_7093# _073_ 0.00125f
C9187 _055_ a_14604_2339# 3.39e-19
C9188 mask\[4\] a_6467_9845# 0.228f
C9189 _003_ _062_ 1.18e-20
C9190 net9 a_12047_2601# 7.53e-19
C9191 net5 a_15023_6031# 0.11f
C9192 a_15023_12559# ctlp[2] 0.0101f
C9193 net37 _131_ 0.00604f
C9194 net4 clknet_0_clk 0.12f
C9195 _076_ a_6835_7669# 0.0104f
C9196 _104_ a_11509_3317# 2.53e-20
C9197 cal_count\[3\] _061_ 5.28e-20
C9198 net54 a_4815_3031# 6.47e-20
C9199 _093_ net41 1.4e-19
C9200 net17 net16 0.00167f
C9201 net13 a_2787_9845# 4.31e-21
C9202 _059_ _098_ 1.04e-19
C9203 _074_ a_1137_5487# 0.00107f
C9204 a_7197_7119# _050_ 3.14e-20
C9205 mask\[0\] a_1476_4777# 6.28e-21
C9206 a_13091_1141# VPWR 0.51f
C9207 _102_ result[4] 2.99e-20
C9208 a_2092_8457# clknet_2_0__leaf_clk 5.04e-20
C9209 _009_ _101_ 5.33e-21
C9210 mask\[4\] VPWR 0.488f
C9211 a_1476_4777# valid 5.38e-19
C9212 cal_itt\[2\] _001_ 2.07e-20
C9213 clknet_0_clk a_3303_7119# 8.27e-19
C9214 a_995_3530# a_1867_3317# 4.41e-21
C9215 a_2857_7637# a_4043_7093# 0.00615f
C9216 VPWR trimb[4] 0.577f
C9217 net7 a_1276_565# 1.39e-19
C9218 _092_ _060_ 0.0391f
C9219 calibrate trim_mask\[4\] 0.0447f
C9220 a_10329_1921# a_10207_1679# 3.16e-19
C9221 net19 net55 1.79e-20
C9222 _064_ VPWR 0.74f
C9223 result[7] ctlp[1] 8.79e-20
C9224 clknet_2_1__leaf_clk _046_ 0.0278f
C9225 a_6785_7119# cal_itt\[3\] 1.57e-19
C9226 _136_ _024_ 7.49e-19
C9227 a_14172_1513# a_14334_1135# 0.00645f
C9228 _096_ a_4576_3427# 0.00131f
C9229 a_14193_3285# _055_ 2.51e-21
C9230 _123_ a_14422_7093# 5.11e-22
C9231 a_13975_3689# a_14540_3689# 7.99e-20
C9232 mask\[6\] a_6007_9839# 2.62e-20
C9233 mask\[2\] a_5423_9011# 3.88e-19
C9234 mask\[4\] a_5699_9269# 0.0114f
C9235 a_12612_8725# _041_ 0.0173f
C9236 a_13142_8725# a_12992_8751# 0.344f
C9237 net45 a_2787_7119# 3.7e-19
C9238 a_11343_3317# a_11435_2229# 2.08e-20
C9239 _015_ a_5699_1653# 4.1e-20
C9240 net16 a_12061_7669# 1.08e-20
C9241 _019_ a_2815_9447# 9.77e-21
C9242 cal_itt\[1\] a_11297_7119# 8.64e-20
C9243 a_6703_2197# a_6906_2355# 0.234f
C9244 trim_val\[0\] trim[4] 1.61e-19
C9245 _026_ a_10543_2455# 3.79e-20
C9246 a_4043_10143# a_3868_10217# 0.234f
C9247 a_7447_8041# VPWR 3.35e-19
C9248 _092_ a_10781_5807# 0.00216f
C9249 net9 _131_ 7.01e-21
C9250 clknet_2_2__leaf_clk trim_val\[1\] 2.5e-20
C9251 net46 a_14347_1439# 0.278f
C9252 _076_ a_5515_6005# 0.00101f
C9253 a_10851_1653# VPWR 0.362f
C9254 net32 trim[0] 0.00352f
C9255 net20 VPWR 0.582f
C9256 net34 net40 0.002f
C9257 clknet_2_0__leaf_clk net51 0.0639f
C9258 _012_ _013_ 1.91e-19
C9259 _123_ _132_ 9.06e-21
C9260 trim_mask\[1\] a_9317_3285# 4.87e-20
C9261 a_9802_4007# a_9839_3615# 0.00531f
C9262 _020_ a_8105_10383# 0.227f
C9263 net12 a_5998_11471# 2.76e-19
C9264 net47 a_10774_9661# 1.12e-19
C9265 net35 a_14347_4917# 0.019f
C9266 a_13825_5185# _058_ 0.00357f
C9267 a_13607_4943# a_13697_4373# 0.00114f
C9268 _004_ net30 0.125f
C9269 net33 _123_ 4.06e-22
C9270 net44 a_4227_8207# 1.79e-19
C9271 _016_ a_3411_7485# 6.95e-19
C9272 trim_mask\[4\] a_11292_1251# 2.49e-20
C9273 _051_ a_3339_2767# 3.53e-19
C9274 _108_ a_9839_3615# 0.00369f
C9275 _053_ VPWR 2.55f
C9276 _068_ _072_ 0.015f
C9277 _097_ a_2601_3285# 1.11e-19
C9278 _065_ a_10990_7485# 0.00475f
C9279 net18 _057_ 0.026f
C9280 net31 _055_ 0.131f
C9281 _118_ clknet_2_2__leaf_clk 2.09e-19
C9282 a_6927_12559# a_6375_12021# 4.41e-19
C9283 trim_val\[2\] a_14604_2339# 0.202f
C9284 a_6467_9845# a_7091_9839# 9.73e-19
C9285 trim_mask\[0\] net50 0.00851f
C9286 net54 a_5087_3855# 0.179f
C9287 cal_itt\[2\] a_7916_8041# 0.00769f
C9288 _074_ a_4512_11305# 7.48e-19
C9289 _104_ a_9007_2601# 3.39e-20
C9290 net16 a_14172_1513# 2.65e-19
C9291 a_7001_7669# net30 1.22e-19
C9292 mask\[0\] _120_ 0.00193f
C9293 a_15083_4659# a_14981_4020# 4.49e-19
C9294 a_8749_3317# a_9317_3285# 0.175f
C9295 state\[1\] a_3933_2767# 0.285f
C9296 a_3597_12021# a_4674_12015# 1.46e-19
C9297 _122_ a_12056_6031# 9.16e-20
C9298 a_2815_9447# VPWR 0.26f
C9299 a_14281_1513# VPWR 1.01e-19
C9300 net13 net51 4.16e-20
C9301 clknet_2_0__leaf_clk _003_ 0.00196f
C9302 a_9664_3689# a_10055_2767# 0.00191f
C9303 trim_mask\[2\] a_8298_2767# 1.07e-19
C9304 _110_ a_11509_3317# 4.66e-20
C9305 net43 a_5997_11247# 1.33e-20
C9306 a_13111_6031# a_13441_6281# 0.00899f
C9307 a_10781_5487# _108_ 9.02e-19
C9308 _078_ a_1585_6031# 5.09e-19
C9309 _110_ a_14099_3017# 4.72e-19
C9310 clknet_0_clk a_10586_7371# 1.9e-19
C9311 a_7091_9839# VPWR 0.133f
C9312 a_448_11445# net26 5.05e-21
C9313 net27 mask\[4\] 9.99e-19
C9314 net14 a_395_4405# 0.0117f
C9315 calibrate a_3123_3615# 5.86e-20
C9316 net18 a_10245_5193# 1.3e-20
C9317 a_9195_10357# a_8215_9295# 2.93e-20
C9318 a_8455_10383# _000_ 1.96e-19
C9319 a_1313_10901# VPWR 0.217f
C9320 trim_mask\[1\] a_9773_3689# 2.91e-21
C9321 VPWR trim[0] 0.554f
C9322 trim_mask\[4\] a_10111_1679# 4.33e-20
C9323 a_2961_9545# a_4609_9295# 1.26e-20
C9324 net12 net30 0.011f
C9325 a_12077_3285# a_12533_3689# 4.2e-19
C9326 a_11859_3689# a_12121_3677# 0.00171f
C9327 trim_mask\[3\] a_12047_2601# 1.18e-19
C9328 _092_ a_4498_4373# 0.113f
C9329 a_10239_9295# a_11814_9295# 2.39e-19
C9330 _035_ a_11244_9661# 4.03e-20
C9331 _028_ a_8657_2229# 2e-19
C9332 a_13975_3689# a_14335_2442# 3.33e-19
C9333 _122_ a_13279_8207# 0.107f
C9334 a_14807_8359# trimb[4] 2.54e-20
C9335 a_12900_7663# a_13279_7119# 1.11e-19
C9336 a_14335_7895# a_14199_7369# 5.42e-19
C9337 net22 a_1129_6273# 0.0371f
C9338 _027_ a_11601_2229# 0.00194f
C9339 a_13975_3689# net8 9.56e-21
C9340 a_579_10933# a_911_10217# 6.4e-21
C9341 clknet_2_1__leaf_clk a_3053_8207# 0.0012f
C9342 a_11141_6031# a_11599_6397# 0.0276f
C9343 _110_ a_9166_4515# 4.96e-19
C9344 _108_ a_9207_3311# 3.38e-20
C9345 a_6375_12021# _009_ 0.345f
C9346 a_8301_8207# a_8022_7119# 6.77e-20
C9347 _084_ a_6541_12021# 2.63e-19
C9348 _067_ a_10137_4943# 6.89e-19
C9349 net18 ctlp[4] 0.00798f
C9350 net52 a_4443_9295# 1.87e-19
C9351 net3 a_1867_3317# 1.24e-19
C9352 _036_ _001_ 0.00281f
C9353 a_2787_7119# a_2953_7119# 0.582f
C9354 _136_ _029_ 0.0046f
C9355 a_14564_6397# a_14172_4943# 4.77e-20
C9356 cal_itt\[0\] net2 0.00936f
C9357 net32 a_15023_2767# 0.00155f
C9358 net47 _065_ 0.453f
C9359 net13 _003_ 1.12e-20
C9360 a_763_8757# a_929_8757# 0.887f
C9361 mask\[6\] _101_ 0.509f
C9362 _069_ a_9621_8029# 2.15e-19
C9363 _062_ a_10055_5487# 4.43e-19
C9364 net20 net27 0.0479f
C9365 _081_ VPWR 0.676f
C9366 a_9317_3285# a_9361_3677# 3.69e-19
C9367 a_8749_3317# a_9773_3689# 2.36e-20
C9368 a_1129_7361# a_1173_7119# 3.69e-19
C9369 net2 a_15259_7637# 0.178f
C9370 a_9099_3689# a_9195_3689# 0.0138f
C9371 trim_val\[4\] a_10188_4105# 0.187f
C9372 a_911_7119# a_1007_7119# 0.0138f
C9373 _094_ a_2857_5461# 0.00233f
C9374 a_7891_3617# clk 0.00939f
C9375 net19 a_8636_9295# 0.0028f
C9376 _130_ VPWR 0.543f
C9377 a_10138_5807# a_10055_5487# 2.42e-19
C9378 _078_ a_911_6031# 3.81e-19
C9379 trim_mask\[2\] a_11951_2601# 2.01e-19
C9380 net4 net41 1.15e-19
C9381 a_10864_9269# _124_ 0.00466f
C9382 _035_ _123_ 1.21e-19
C9383 a_10688_9295# a_10747_8970# 3.15e-19
C9384 a_14335_4020# VPWR 0.28f
C9385 _048_ net42 0.454f
C9386 a_13562_8751# a_13470_7663# 1.04e-20
C9387 a_11583_4777# a_11845_4765# 0.00171f
C9388 _041_ a_12900_7663# 9.24e-22
C9389 a_11801_4373# a_12257_4777# 4.2e-19
C9390 a_15023_12559# net34 4.68e-19
C9391 clknet_2_1__leaf_clk a_7456_12393# 1.32e-19
C9392 a_8298_2767# a_9719_1473# 2.09e-21
C9393 a_11204_7485# _136_ 3.08e-19
C9394 net18 _124_ 0.022f
C9395 a_395_2767# clk 0.00131f
C9396 _049_ a_7184_2339# 1.54e-19
C9397 _107_ a_9839_3615# 3.14e-19
C9398 _113_ a_13880_3677# 1.68e-20
C9399 net33 trim_mask\[1\] 2.41e-19
C9400 a_3431_10933# net26 9.87e-21
C9401 a_455_3571# clk 1.65e-19
C9402 a_13825_5185# a_13607_4943# 0.21f
C9403 a_13257_4943# a_14347_4917# 0.0418f
C9404 a_13091_4943# a_14172_4943# 0.102f
C9405 a_12169_2197# a_12625_2601# 4.2e-19
C9406 a_11951_2601# a_12213_2589# 0.00171f
C9407 a_11435_2229# a_12059_2223# 9.73e-19
C9408 net45 a_7181_2589# 6.03e-19
C9409 net45 _096_ 1.24e-19
C9410 a_8215_9295# a_8949_9537# 0.0535f
C9411 _000_ a_8381_9295# 0.214f
C9412 a_5547_5603# _060_ 0.00643f
C9413 _048_ a_4091_5309# 0.0772f
C9414 a_455_5747# VPWR 0.403f
C9415 mask\[4\] a_8455_10383# 8.93e-19
C9416 a_4471_4007# a_5087_3855# 0.0806f
C9417 cal_itt\[3\] a_8935_6895# 3.11e-19
C9418 _078_ a_5691_7637# 5.39e-19
C9419 _062_ _088_ 1.38e-19
C9420 net3 a_3302_3677# 9.82e-20
C9421 a_9003_3829# a_8749_3317# 0.0116f
C9422 net28 a_5578_12131# 8.39e-21
C9423 _136_ a_13349_6031# 0.00637f
C9424 _076_ a_6428_7119# 2.94e-20
C9425 a_6793_8970# a_6631_7485# 6.28e-21
C9426 _123_ _136_ 5.71e-19
C9427 net40 cal_count\[3\] 0.412f
C9428 _062_ a_7262_5461# 0.4f
C9429 _051_ net3 0.0124f
C9430 _064_ _104_ 0.671f
C9431 net44 a_8839_9661# 3.05e-19
C9432 net15 a_2283_4020# 4.65e-20
C9433 _047_ a_14715_3615# 0.0012f
C9434 a_15023_2767# VPWR 0.358f
C9435 a_561_9845# net25 0.0081f
C9436 _050_ a_4725_5487# 0.00217f
C9437 net3 _014_ 0.0126f
C9438 _060_ a_5536_4399# 0.0144f
C9439 net27 a_1313_10901# 4.37e-19
C9440 a_14540_3689# trim_val\[1\] 0.0209f
C9441 a_8298_2767# a_9595_1679# 9.57e-20
C9442 a_2787_7119# a_2857_5461# 4.99e-19
C9443 _062_ trim_val\[4\] 8.95e-19
C9444 a_10005_6031# en_co_clk 0.00148f
C9445 a_395_9845# a_911_10217# 0.115f
C9446 cal_count\[0\] a_12341_8751# 0.0167f
C9447 net31 a_15259_7637# 0.00901f
C9448 calibrate a_1173_4765# 3.62e-20
C9449 mask\[1\] a_4036_8207# 0.0111f
C9450 net14 a_561_9845# 0.0102f
C9451 mask\[6\] _102_ 0.00305f
C9452 _010_ a_3947_12393# 0.00139f
C9453 a_3208_10205# a_3399_10217# 4.61e-19
C9454 a_3891_4943# VPWR 0.234f
C9455 mask\[7\] ctlp[1] 5.33e-20
C9456 net53 _021_ 0.0551f
C9457 _107_ a_9207_3311# 5.99e-19
C9458 _104_ a_10851_1653# 8.76e-20
C9459 net32 a_15299_3311# 0.129f
C9460 trim_mask\[0\] _106_ 0.152f
C9461 net26 a_6198_8534# 6.87e-20
C9462 a_1095_12393# ctlp[0] 0.00126f
C9463 _050_ a_9004_3677# 8.9e-21
C9464 a_10903_7261# a_10975_6031# 4.05e-20
C9465 a_10864_7387# _038_ 7.11e-21
C9466 net46 a_11343_3317# 0.301f
C9467 _010_ a_3425_11721# 0.00151f
C9468 net2 trim_mask\[0\] 1.07e-20
C9469 _101_ a_1763_9295# 1.55e-20
C9470 a_579_10933# a_1000_11293# 0.0931f
C9471 _110_ net48 0.00265f
C9472 cal_itt\[2\] a_8949_6031# 3.56e-19
C9473 net12 state\[2\] 0.261f
C9474 _062_ a_9823_6941# 0.00422f
C9475 a_9460_6807# a_9602_6614# 0.00557f
C9476 clknet_2_2__leaf_clk a_12424_3689# 0.0568f
C9477 a_3840_8867# _040_ 6.46e-21
C9478 _050_ _107_ 0.0466f
C9479 net43 a_3748_6281# 6.96e-20
C9480 _053_ _104_ 0.802f
C9481 _078_ a_6633_9845# 5.67e-20
C9482 mask\[4\] a_8381_9295# 2.28e-19
C9483 a_13821_7119# VPWR 4.85e-19
C9484 _111_ a_12323_4703# 0.0362f
C9485 trim_mask\[1\] trim_val\[3\] 1.05e-21
C9486 net12 state\[0\] 1.7e-20
C9487 a_2971_8457# _040_ 0.0849f
C9488 _052_ a_9004_3677# 1.24e-20
C9489 mask\[6\] _022_ 0.0576f
C9490 en_co_clk _099_ 0.00304f
C9491 cal_count\[0\] a_10864_7387# 7.48e-20
C9492 mask\[6\] a_6375_12021# 5.53e-20
C9493 a_14807_8359# _130_ 8.84e-22
C9494 a_4512_12393# _009_ 4.04e-20
C9495 net47 _067_ 0.0716f
C9496 a_14335_7895# a_14422_7093# 3.62e-19
C9497 _031_ a_13607_1513# 7.35e-20
C9498 a_7999_11231# net26 1.34e-21
C9499 net33 _115_ 1.51e-21
C9500 VPWR result[5] 0.317f
C9501 _052_ _107_ 0.0314f
C9502 _049_ _050_ 0.4f
C9503 trim_mask\[0\] a_14000_4719# 0.0102f
C9504 _074_ a_1375_9129# 2.64e-19
C9505 a_7939_3855# a_9003_3829# 2.25e-20
C9506 trim_mask\[0\] _033_ 0.00407f
C9507 clknet_2_1__leaf_clk a_6743_10933# 0.248f
C9508 _078_ a_1129_9813# 1.96e-19
C9509 _053_ a_7200_3631# 8.87e-19
C9510 _098_ _107_ 0.0442f
C9511 a_15299_3311# VPWR 0.221f
C9512 net2 a_13933_6281# 7.35e-19
C9513 _110_ a_13091_1141# 0.00314f
C9514 a_1651_7093# a_1549_6794# 5.15e-19
C9515 a_7379_2197# VPWR 0.216f
C9516 clknet_2_2__leaf_clk a_11321_3855# 0.00102f
C9517 a_14335_7895# _132_ 0.372f
C9518 clknet_2_2__leaf_clk a_9103_2601# 0.00497f
C9519 net15 result[7] 1.8e-20
C9520 net19 net4 0.346f
C9521 net31 trim_mask\[0\] 3.14e-19
C9522 a_745_12021# a_1660_11305# 5.19e-20
C9523 net43 a_1095_11305# 0.157f
C9524 trim_val\[1\] a_14335_2442# 8.86e-20
C9525 _064_ _110_ 0.00401f
C9526 _124_ a_12153_8757# 1.29e-20
C9527 _123_ a_11987_8757# 0.522f
C9528 _049_ _052_ 0.59f
C9529 a_11116_8983# _036_ 8.26e-20
C9530 _074_ a_4209_12381# 1.15e-20
C9531 net18 a_8583_3317# 7.34e-22
C9532 net32 trim[4] 0.00269f
C9533 a_4995_7119# net55 4.46e-19
C9534 net33 a_14335_7895# 0.0046f
C9535 a_4959_1679# a_5221_1679# 0.00171f
C9536 a_5524_1679# a_5686_2045# 0.00645f
C9537 clknet_0_clk _064_ 1.04e-19
C9538 net44 a_4259_6031# 0.298f
C9539 a_1279_9129# a_1375_9129# 0.0138f
C9540 a_1497_8725# a_1541_9117# 3.69e-19
C9541 a_7088_7119# a_8022_7119# 2.75e-19
C9542 _092_ _066_ 0.0852f
C9543 _049_ _098_ 0.0909f
C9544 net53 a_4655_10071# 0.221f
C9545 _069_ _063_ 0.0696f
C9546 _096_ a_4905_3855# 0.00145f
C9547 a_6891_12393# a_6796_12381# 0.0498f
C9548 a_10699_3311# _025_ 0.116f
C9549 net9 _036_ 0.18f
C9550 net19 a_8360_10383# 0.00137f
C9551 a_11343_3317# a_11149_3017# 3.66e-19
C9552 a_9664_3689# VPWR 0.323f
C9553 a_579_12021# a_1095_12393# 0.115f
C9554 net18 a_11803_10383# 0.00164f
C9555 a_395_6031# a_1651_6005# 0.0435f
C9556 _004_ a_911_6031# 0.00161f
C9557 _127_ _128_ 0.0211f
C9558 clknet_2_1__leaf_clk net45 0.266f
C9559 _063_ a_8022_7119# 0.013f
C9560 net13 net26 0.0114f
C9561 _110_ a_10851_1653# 3.09e-19
C9562 trim_val\[0\] a_13625_3317# 1.49e-20
C9563 _065_ _072_ 0.128f
C9564 net14 a_2283_4020# 2.88e-21
C9565 net40 a_14347_4917# 1.44e-20
C9566 a_14788_7369# a_14870_7369# 0.00477f
C9567 _064_ a_10699_5487# 3.11e-19
C9568 net13 a_5050_8207# 5.11e-19
C9569 en_co_clk a_5537_4943# 1.05e-19
C9570 net4 cal_itt\[1\] 0.407f
C9571 net12 _100_ 0.0959f
C9572 clknet_2_2__leaf_clk a_11435_2229# 0.266f
C9573 a_10689_2223# VPWR 0.197f
C9574 cal_itt\[2\] _062_ 0.00126f
C9575 net15 _017_ 6.48e-20
C9576 _065_ _068_ 0.00939f
C9577 _004_ _012_ 0.00219f
C9578 mask\[7\] a_3852_11293# 5.89e-20
C9579 a_2857_7637# a_3748_6281# 1.45e-21
C9580 _059_ _087_ 6.38e-19
C9581 a_9125_4943# _107_ 1.17e-19
C9582 a_11425_5487# VPWR 0.00563f
C9583 a_4993_6273# a_4871_6031# 3.16e-19
C9584 a_4259_6031# en_co_clk 0.00754f
C9585 net25 _006_ 1.92e-19
C9586 a_2857_5461# _096_ 0.0044f
C9587 _007_ net24 3.43e-21
C9588 _040_ a_4131_8207# 0.0382f
C9589 trim_mask\[4\] a_7184_2339# 5.49e-19
C9590 _053_ _110_ 4.68e-19
C9591 a_4609_9295# a_5423_9011# 0.0108f
C9592 a_14983_9269# net2 1.2e-19
C9593 a_3530_4438# VPWR 0.00203f
C9594 _059_ a_6519_3829# 2.24e-19
C9595 net43 a_4674_12015# 8.2e-20
C9596 _136_ a_10781_5807# 0.00158f
C9597 clknet_0_clk _053_ 0.0952f
C9598 net27 result[5] 0.00579f
C9599 net14 _006_ 0.0111f
C9600 net44 a_4043_7093# 1.61e-19
C9601 a_6007_7119# a_6515_6794# 0.00414f
C9602 net15 net7 0.109f
C9603 net44 a_8563_10749# 5.32e-19
C9604 VPWR trim[4] 0.585f
C9605 a_12631_12559# ctlp[3] 0.157f
C9606 _059_ _099_ 0.0305f
C9607 _092_ a_7571_4943# 0.00229f
C9608 a_2143_2229# a_2564_2589# 0.0931f
C9609 a_12056_6031# a_13111_6031# 3.89e-19
C9610 net13 a_5686_2045# 5.91e-20
C9611 net52 _065_ 0.00701f
C9612 trim_mask\[0\] _054_ 5.81e-20
C9613 net46 a_12059_2223# 0.0122f
C9614 clknet_2_1__leaf_clk a_3868_10217# 0.00232f
C9615 a_10781_3631# VPWR 7.06e-20
C9616 _065_ net46 0.00145f
C9617 _091_ net30 1.3e-19
C9618 _101_ a_1497_8725# 1.29e-19
C9619 trim_mask\[4\] a_9839_3615# 0.052f
C9620 a_14184_1679# VPWR 3.03e-19
C9621 _019_ a_3781_8207# 1.24e-19
C9622 net52 net23 0.00459f
C9623 net23 a_816_7119# 5e-20
C9624 mask\[7\] a_3947_11305# 2.6e-20
C9625 _053_ a_10699_5487# 0.0625f
C9626 _092_ a_4576_3427# 5.9e-22
C9627 a_4512_12393# mask\[6\] 2.19e-20
C9628 a_8307_4943# _106_ 0.0964f
C9629 a_14471_12559# VPWR 0.299f
C9630 clknet_2_3__leaf_clk a_9443_6059# 0.00118f
C9631 calibrate a_1201_3855# 0.00153f
C9632 net4 _001_ 0.0163f
C9633 _006_ a_395_7119# 1.37e-20
C9634 a_763_8757# a_561_7119# 1.51e-19
C9635 _074_ a_448_11445# 2.17e-20
C9636 a_13783_6183# a_13697_4373# 1.43e-20
C9637 a_13459_3317# a_13975_3689# 0.107f
C9638 _037_ a_13142_7271# 0.106f
C9639 _030_ a_14193_3285# 7.67e-19
C9640 a_4043_7093# en_co_clk 2.97e-21
C9641 net12 a_5691_7637# 0.00721f
C9642 net19 a_10586_7371# 1.83e-21
C9643 _036_ a_12436_9129# 9.17e-19
C9644 a_11987_8757# a_13142_8725# 0.0608f
C9645 a_816_6031# a_1007_6031# 4.61e-19
C9646 net15 a_4425_6031# 1.08e-20
C9647 a_10781_5487# trim_mask\[4\] 2.67e-20
C9648 net46 a_9826_3311# 9.87e-20
C9649 _026_ _027_ 1.14e-19
C9650 _018_ a_3303_10217# 2.86e-19
C9651 a_2787_9845# a_4043_10143# 0.0435f
C9652 _051_ a_4973_2773# 0.00165f
C9653 net16 _031_ 2.98e-19
C9654 net31 a_14983_9269# 7.34e-19
C9655 a_4863_4917# a_5081_4943# 0.0326f
C9656 _106_ a_8298_2767# 5.96e-21
C9657 _074_ a_1203_10927# 0.0022f
C9658 a_1651_6005# net30 6.9e-19
C9659 a_15023_2223# trim[2] 0.337f
C9660 _066_ a_11045_5807# 6.81e-19
C9661 clknet_2_1__leaf_clk a_2953_7119# 8.29e-19
C9662 _129_ a_14282_7119# 5.63e-19
C9663 a_5221_1679# VPWR 5.1e-19
C9664 net34 trim_mask\[1\] 5.19e-20
C9665 net14 result[7] 0.0254f
C9666 net46 a_11233_4405# 0.0321f
C9667 a_14467_8751# trimb[4] 1.92e-19
C9668 clknet_2_2__leaf_clk a_14347_1439# 1.24e-20
C9669 _051_ net54 0.00909f
C9670 net55 a_4863_4917# 0.0138f
C9671 a_1493_11721# a_1579_11471# 2.42e-19
C9672 a_8307_6575# a_8473_5193# 8.1e-21
C9673 a_6099_10633# a_6181_10633# 0.171f
C9674 clknet_2_3__leaf_clk a_12061_7669# 0.0106f
C9675 _110_ a_14335_4020# 9.17e-19
C9676 net19 a_9166_4515# 2.11e-19
C9677 a_2033_3317# a_2479_3689# 2.28e-19
C9678 _077_ a_6885_8372# 2.14e-20
C9679 net52 a_2225_7663# 0.00625f
C9680 _059_ a_5537_4943# 8.6e-21
C9681 a_9919_6614# VPWR 8.98e-19
C9682 _108_ a_13233_4737# 1.73e-19
C9683 net2 a_7723_6807# 7.02e-22
C9684 cal_itt\[2\] a_8745_6895# 0.012f
C9685 cal_itt\[1\] a_10586_7371# 0.00177f
C9686 a_3781_8207# VPWR 0.358f
C9687 _062_ net55 0.00671f
C9688 state\[2\] a_5691_2741# 0.26f
C9689 _040_ net30 1.71e-20
C9690 net52 _016_ 0.0278f
C9691 _072_ _067_ 0.0964f
C9692 net49 a_14715_3615# 1.09e-19
C9693 net31 _030_ 1.25e-20
C9694 cal_itt\[3\] a_6515_6794# 5.57e-19
C9695 a_11479_9117# _001_ 4.44e-20
C9696 a_395_4405# VPWR 0.537f
C9697 _083_ a_5829_9839# 3.99e-21
C9698 a_6633_9845# a_6888_10205# 0.0594f
C9699 cal_count\[3\] a_13349_6031# 0.0353f
C9700 a_4259_6031# _059_ 2.77e-19
C9701 a_14604_3017# _056_ 3.39e-19
C9702 a_12056_6031# a_13825_6031# 3.78e-20
C9703 net4 a_3063_591# 0.0341f
C9704 _050_ trim_mask\[4\] 0.228f
C9705 _109_ a_13915_4399# 0.00133f
C9706 clknet_2_1__leaf_clk a_3399_10217# 0.00108f
C9707 _074_ a_3431_10933# 1.71e-20
C9708 _123_ cal_count\[3\] 1.48e-19
C9709 state\[0\] a_5691_2741# 2.4e-19
C9710 _104_ a_7379_2197# 1.29e-21
C9711 a_15023_9839# a_15159_9269# 0.011f
C9712 a_4443_9295# a_4696_8207# 3.32e-20
C9713 _128_ _041_ 0.012f
C9714 net15 a_3868_7119# 9.63e-19
C9715 a_4609_9295# a_4871_8181# 1.65e-20
C9716 net4 a_7916_8041# 2.22e-21
C9717 _068_ _067_ 0.0116f
C9718 net14 a_911_4777# 0.00521f
C9719 mask\[0\] a_1638_6397# 4.86e-21
C9720 _074_ a_929_8757# 0.0142f
C9721 net12 a_6633_9845# 1.11e-19
C9722 net16 a_13356_8457# 1.54e-20
C9723 _057_ VPWR 1.86f
C9724 _131_ a_14788_7369# 0.0477f
C9725 mask\[6\] _046_ 0.075f
C9726 _075_ a_5731_4943# 0.00549f
C9727 _092_ a_3557_5193# 0.00575f
C9728 _033_ a_8298_2767# 0.065f
C9729 _135_ _061_ 5.21e-19
C9730 net9 ctln[3] 0.0104f
C9731 _101_ _021_ 1.28e-19
C9732 net52 a_4696_8207# 2.33e-20
C9733 a_10373_1679# trim_val\[3\] 2.13e-20
C9734 a_9405_9295# _070_ 6.83e-20
C9735 _103_ a_7800_4631# 0.0392f
C9736 a_8389_5193# _107_ 0.00217f
C9737 _052_ trim_mask\[4\] 0.144f
C9738 a_1579_11471# VPWR 3.34e-19
C9739 a_4775_6031# a_5340_6031# 7.99e-20
C9740 a_13825_6031# _058_ 1.75e-19
C9741 _104_ a_9664_3689# 0.0578f
C9742 net15 mask\[7\] 0.0158f
C9743 a_10699_3311# a_10781_3311# 0.171f
C9744 _025_ a_11955_3689# 2.82e-19
C9745 net43 _070_ 6.25e-20
C9746 a_10864_7387# en_co_clk 2.08e-20
C9747 net54 a_5445_4399# 5.19e-19
C9748 a_10239_9295# _035_ 0.114f
C9749 net45 a_6007_7119# 1.56e-20
C9750 _028_ a_7223_2465# 0.458f
C9751 net14 net7 3.57e-21
C9752 a_13880_3677# a_13881_2741# 8.84e-19
C9753 _042_ net24 1.88e-19
C9754 a_929_8757# a_1279_9129# 0.217f
C9755 a_448_9269# _082_ 3.65e-19
C9756 calibrate a_6737_3855# 6.83e-19
C9757 a_10245_5193# VPWR 0.00384f
C9758 _098_ trim_mask\[4\] 1.66e-20
C9759 net19 a_9007_2601# 0.0116f
C9760 a_2787_9845# a_3208_10205# 0.0859f
C9761 a_6633_9845# a_6983_10217# 0.217f
C9762 clknet_0_clk a_3891_4943# 0.0117f
C9763 a_2787_9845# a_2689_8751# 8.73e-21
C9764 _084_ _042_ 6.34e-21
C9765 _001_ a_10586_7371# 6.56e-21
C9766 a_10005_6031# _108_ 2.1e-19
C9767 net30 _048_ 0.468f
C9768 a_11233_4405# a_11343_3317# 2.53e-20
C9769 _014_ a_2645_3677# 3.89e-19
C9770 a_11067_4405# a_11509_3317# 2.52e-20
C9771 _104_ a_10689_2223# 0.0106f
C9772 a_13783_6183# a_13825_5185# 2.67e-19
C9773 state\[0\] a_3110_3311# 8.89e-21
C9774 _093_ a_3224_2601# 8.22e-22
C9775 _058_ a_11067_3017# 7.2e-19
C9776 net44 a_7939_10383# 0.00995f
C9777 a_395_2767# en 0.193f
C9778 a_14347_1439# ctln[2] 8.69e-19
C9779 _051_ a_7019_4407# 5.88e-20
C9780 a_455_8181# mask\[1\] 2.25e-19
C9781 _092_ a_12056_6031# 8.65e-22
C9782 a_455_3571# en 0.00805f
C9783 _023_ net52 6.2e-21
C9784 _045_ a_7153_12381# 5.01e-20
C9785 VPWR ctlp[4] 0.346f
C9786 _053_ net41 8.1e-20
C9787 net2 a_12344_8041# 2.46e-19
C9788 a_9099_3689# _028_ 4.82e-20
C9789 net19 _000_ 0.0338f
C9790 a_10975_6031# a_11141_6031# 0.64f
C9791 _051_ a_4471_4007# 2.4e-20
C9792 net55 a_3817_4697# 3.76e-21
C9793 a_7256_8029# a_7263_7093# 3.74e-19
C9794 net46 clknet_2_2__leaf_clk 0.838f
C9795 state\[2\] _089_ 3.47e-21
C9796 a_9084_4515# a_9503_4399# 7.02e-20
C9797 net45 _092_ 0.00188f
C9798 _107_ a_7891_3617# 0.00152f
C9799 _029_ a_14347_4917# 1.04e-20
C9800 a_7942_2223# clk 0.00869f
C9801 _104_ a_10781_3631# 5.15e-20
C9802 net26 a_9020_10383# 7.59e-19
C9803 trim_mask\[0\] a_13715_5309# 1.2e-19
C9804 _092_ _058_ 9.34e-19
C9805 state\[2\] a_4609_1679# 0.00416f
C9806 net49 a_14099_1929# 9.52e-20
C9807 a_15023_2223# a_15023_1135# 0.00243f
C9808 a_3615_8207# a_4036_8207# 0.0864f
C9809 clknet_2_0__leaf_clk net55 3.53e-19
C9810 _124_ VPWR 0.308f
C9811 a_4863_4917# a_5166_5193# 0.00145f
C9812 a_5686_9661# VPWR 7.93e-19
C9813 net4 a_11116_8983# 7.84e-21
C9814 cal_count\[3\] trim_mask\[1\] 2.64e-20
C9815 a_6885_8372# a_6173_7119# 3.29e-21
C9816 a_561_9845# VPWR 0.277f
C9817 state\[0\] a_4609_1679# 4.22e-20
C9818 a_13441_6281# _136_ 6.58e-19
C9819 _061_ a_14649_6031# 0.001f
C9820 _064_ a_11057_4105# 0.0118f
C9821 a_10676_1679# ctln[4] 2.83e-19
C9822 net37 a_14172_4943# 4.63e-20
C9823 net53 a_8215_9295# 1.37e-21
C9824 _049_ a_7891_3617# 1.45e-19
C9825 clknet_2_3__leaf_clk a_11396_6031# 0.016f
C9826 _101_ a_4655_10071# 0.176f
C9827 trim_mask\[1\] a_12586_3311# 4.1e-19
C9828 _074_ clknet_2_0__leaf_clk 0.167f
C9829 a_4959_9295# a_5055_9295# 0.0138f
C9830 a_5177_9537# a_5221_9295# 3.69e-19
C9831 a_13257_4943# a_13519_4007# 1.72e-20
C9832 net27 a_1579_11471# 6.1e-21
C9833 a_13459_3317# trim_val\[1\] 0.008f
C9834 net47 a_8993_9295# 0.00316f
C9835 a_5455_4943# a_6210_4989# 0.00111f
C9836 net13 a_5081_4943# 0.00116f
C9837 a_4425_6031# a_5449_6031# 2.36e-20
C9838 _081_ a_2775_9071# 0.00151f
C9839 net45 a_6906_2355# 0.255f
C9840 _108_ a_14649_3689# 2.9e-19
C9841 net13 a_4858_8573# 1.5e-19
C9842 a_2659_2601# net7 1.06e-19
C9843 _110_ a_9664_3689# 0.0126f
C9844 net32 a_13625_3317# 1.66e-19
C9845 _074_ a_4687_12319# 3.85e-19
C9846 a_12992_8751# a_13279_8207# 1.16e-19
C9847 net13 net55 0.314f
C9848 a_6375_12021# _021_ 3.92e-20
C9849 net19 mask\[4\] 0.0812f
C9850 _009_ a_6743_10933# 5.42e-21
C9851 en_co_clk _097_ 0.00288f
C9852 a_14249_8725# trimb[4] 9.37e-20
C9853 a_10005_6031# _107_ 4.94e-19
C9854 net43 a_1211_7983# 3.55e-20
C9855 _050_ a_7320_3631# 0.00128f
C9856 net19 _064_ 4.18e-20
C9857 net15 _121_ 0.0264f
C9858 mask\[7\] net25 4.43e-19
C9859 a_3063_591# ctln[1] 0.159f
C9860 cal_count\[2\] a_10864_7387# 1.23e-21
C9861 a_1549_6794# a_395_6031# 0.0025f
C9862 net26 a_8731_9295# 3.75e-20
C9863 net30 a_7021_4105# 8.72e-20
C9864 clknet_2_2__leaf_clk a_11343_3317# 0.862f
C9865 _074_ net13 0.13f
C9866 net14 mask\[7\] 3.5e-19
C9867 trim_mask\[0\] a_12599_3615# 4.74e-19
C9868 clknet_2_2__leaf_clk a_11149_3017# 0.00682f
C9869 _087_ _107_ 0.0797f
C9870 a_13356_7369# VPWR 0.00802f
C9871 _047_ net49 4.23e-21
C9872 _136_ _066_ 0.0391f
C9873 _048_ state\[2\] 0.0104f
C9874 _052_ a_7320_3631# 0.00371f
C9875 net43 a_4349_8449# 2.8e-19
C9876 _100_ _089_ 0.243f
C9877 _107_ a_6519_3829# 0.00492f
C9878 a_3597_12021# _084_ 3.03e-21
C9879 a_14335_2442# a_14686_2339# 1e-19
C9880 _035_ a_11545_9049# 2.02e-20
C9881 a_8473_5193# VPWR 0.18f
C9882 _122_ a_13142_7271# 0.0898f
C9883 a_4512_11305# mask\[4\] 7.84e-19
C9884 a_5915_10927# net26 2.73e-20
C9885 _037_ _131_ 1.12e-19
C9886 _048_ state\[0\] 0.0117f
C9887 net18 a_10903_7261# 0.00548f
C9888 net51 a_7088_7119# 1.37e-21
C9889 _099_ _107_ 0.0643f
C9890 a_3817_4697# _093_ 4.38e-19
C9891 _065_ a_9761_8457# 0.00156f
C9892 a_763_8757# a_1467_7923# 1.41e-19
C9893 cal_itt\[1\] _064_ 0.00142f
C9894 _065_ a_11233_4405# 1.61e-20
C9895 net18 a_11149_2767# 2.46e-19
C9896 net31 a_15083_4659# 0.00233f
C9897 a_4393_8207# VPWR 4.48e-19
C9898 trim_mask\[0\] a_12257_4777# 6.68e-21
C9899 _110_ a_10781_3631# 2.49e-21
C9900 _049_ _087_ 8.72e-19
C9901 mask\[0\] net22 0.297f
C9902 a_11045_5807# _058_ 3.46e-20
C9903 net45 cal 3.14e-19
C9904 a_13625_3317# VPWR 0.623f
C9905 net19 _053_ 0.0347f
C9906 _078_ a_4443_9295# 0.0041f
C9907 _049_ a_6519_3829# 0.025f
C9908 _076_ _051_ 8.68e-19
C9909 _023_ a_1679_10633# 9.1e-19
C9910 _062_ a_9595_5193# 0.125f
C9911 net4 a_3224_2601# 0.0157f
C9912 clknet_2_0__leaf_clk _093_ 0.0107f
C9913 a_561_4405# a_1638_4399# 1.46e-19
C9914 net18 a_11845_4765# 2.75e-19
C9915 a_745_12021# a_579_10933# 3.41e-19
C9916 net40 _135_ 7.13e-19
C9917 a_579_12021# a_745_10933# 7.79e-19
C9918 net43 a_3511_11471# 2.03e-19
C9919 a_15023_2223# trim[1] 7.46e-20
C9920 _049_ _099_ 0.0156f
C9921 net47 a_12924_8029# 0.00215f
C9922 _078_ net52 0.0217f
C9923 a_1129_6273# a_1476_6031# 0.0512f
C9924 _099_ a_3388_4631# 0.0546f
C9925 net23 a_2225_7663# 0.00553f
C9926 cal_itt\[0\] a_11016_6691# 1.11e-19
C9927 a_2283_4020# VPWR 0.24f
C9928 a_14335_2442# a_14347_1439# 6.81e-19
C9929 trim_val\[2\] a_13607_1513# 0.00627f
C9930 _126_ a_14377_7983# 2.58e-20
C9931 _133_ a_13557_7369# 9.81e-19
C9932 a_6007_7119# a_8022_7119# 1.17e-20
C9933 _003_ a_7088_7119# 5.47e-21
C9934 net8 a_14347_1439# 0.0111f
C9935 net23 _016_ 0.0433f
C9936 a_12310_4399# VPWR 7.99e-19
C9937 net9 a_11509_3317# 0.00793f
C9938 _021_ a_7824_11305# 7.95e-20
C9939 a_4512_12393# ctlp[7] 1.83e-19
C9940 a_8583_3317# VPWR 0.513f
C9941 a_8215_9295# _071_ 1.33e-19
C9942 net46 a_14540_3689# 0.236f
C9943 a_1313_10901# a_1822_10927# 2.6e-19
C9944 a_745_10933# a_2869_10927# 1.92e-20
C9945 a_1095_12393# _086_ 9.06e-19
C9946 a_7939_10383# a_8992_9955# 7.54e-19
C9947 a_2143_7663# a_2225_7983# 0.00393f
C9948 cal_itt\[1\] _053_ 0.00161f
C9949 _106_ a_9369_4105# 3.92e-19
C9950 a_1844_9129# VPWR 0.32f
C9951 net18 a_8105_10383# 6.64e-20
C9952 net44 a_6056_8359# 2.12e-20
C9953 net4 trim_mask\[3\] 9.76e-21
C9954 _065_ a_4696_8207# 6.09e-19
C9955 a_5423_9011# a_5535_8181# 0.0152f
C9956 _091_ _118_ 1.49e-21
C9957 _092_ a_6316_5193# 0.0755f
C9958 _064_ a_11067_4405# 4.55e-19
C9959 net2 _133_ 0.00134f
C9960 a_5496_12131# VPWR 0.169f
C9961 net13 _093_ 5.91e-20
C9962 a_11803_10383# VPWR 0.286f
C9963 _006_ VPWR 0.689f
C9964 _092_ a_2857_5461# 0.0808f
C9965 net15 a_3273_4943# 0.0132f
C9966 a_395_4405# a_1007_4777# 0.00188f
C9967 _012_ a_816_4765# 0.16f
C9968 trim_mask\[0\] a_10543_2455# 4.06e-21
C9969 net22 _079_ 0.265f
C9970 a_1549_6794# net30 9.28e-20
C9971 net4 _062_ 0.34f
C9972 _080_ _005_ 0.156f
C9973 _065_ _067_ 0.0259f
C9974 mask\[7\] a_1769_11305# 7.28e-19
C9975 clknet_2_0__leaf_clk _034_ 0.0621f
C9976 _074_ a_561_7119# 0.028f
C9977 trim_val\[2\] a_13881_1653# 0.189f
C9978 _048_ _100_ 0.21f
C9979 _127_ net40 1.19e-19
C9980 net45 a_5067_2045# 0.0122f
C9981 a_8022_7119# _092_ 5e-20
C9982 net4 a_10138_5807# 2.28e-19
C9983 mask\[6\] a_6743_10933# 4.25e-20
C9984 a_15023_1679# net8 2.96e-19
C9985 a_9761_1679# a_10569_1109# 0.00133f
C9986 a_12153_8757# a_12546_9129# 0.00127f
C9987 a_12612_8725# a_12341_8751# 7.79e-20
C9988 a_3781_8207# clknet_0_clk 9.18e-19
C9989 a_3748_6281# en_co_clk 2.2e-21
C9990 net40 a_14063_7093# 0.00375f
C9991 net18 a_9572_2601# 1.78e-36
C9992 net44 a_7710_9839# 3.41e-19
C9993 a_4425_6031# a_5363_4719# 1.46e-20
C9994 net33 _058_ 0.0312f
C9995 net16 _055_ 8.2e-22
C9996 _040_ a_5691_7637# 1.1e-20
C9997 state\[2\] a_7021_4105# 0.00523f
C9998 net52 a_3597_10933# 5.69e-20
C9999 a_13915_4399# trim[1] 7.76e-20
C10000 net43 a_5055_9295# 1.83e-20
C10001 a_12344_8041# a_12249_7663# 0.0356f
C10002 _016_ a_2225_7663# 0.00452f
C10003 _110_ _057_ 0.0685f
C10004 clknet_2_1__leaf_clk a_2787_9845# 0.423f
C10005 net47 a_8551_10383# 9.54e-19
C10006 a_8673_10625# a_8717_10383# 3.69e-19
C10007 net45 a_561_4405# 0.0259f
C10008 a_8105_10383# a_9129_10383# 2.36e-20
C10009 a_4680_6031# VPWR 0.083f
C10010 a_9296_9295# a_10239_9295# 3.5e-19
C10011 a_9471_9269# _035_ 0.00101f
C10012 a_4036_8207# a_4227_8207# 4.61e-19
C10013 a_929_8757# a_911_7119# 8.5e-21
C10014 a_14236_8457# net2 0.183f
C10015 trim_mask\[4\] a_7891_3617# 0.0309f
C10016 a_9478_4105# a_8583_3317# 1.34e-19
C10017 clknet_2_0__leaf_clk a_448_7637# 0.00967f
C10018 _119_ a_8749_3317# 0.00802f
C10019 _065_ clknet_2_2__leaf_clk 0.00202f
C10020 _001_ _053_ 5.28e-19
C10021 net40 a_14649_6031# 7.44e-19
C10022 _053_ a_11067_4405# 7.36e-20
C10023 net13 _034_ 0.00173f
C10024 _049_ a_4259_6031# 0.0504f
C10025 a_9761_1679# a_10329_1921# 0.186f
C10026 net31 _133_ 1.06e-20
C10027 _122_ a_13562_8751# 9.53e-20
C10028 clknet_2_3__leaf_clk _051_ 4.57e-19
C10029 net32 a_14894_3677# 2.91e-19
C10030 VPWR result[7] 0.646f
C10031 _005_ a_816_6031# 2.65e-19
C10032 a_8022_7119# cal_itt\[3\] 0.01f
C10033 a_10569_1109# a_10787_1135# 0.0821f
C10034 a_13091_1141# a_13512_1501# 0.0856f
C10035 a_12424_3689# a_13459_3317# 1.39e-19
C10036 a_5633_9295# VPWR 7.57e-20
C10037 a_12599_3615# _030_ 6.43e-19
C10038 _071_ a_8298_5487# 0.00225f
C10039 a_11545_9049# a_11987_8757# 0.033f
C10040 net47 a_13008_7663# 9.26e-20
C10041 a_7190_3855# VPWR 0.205f
C10042 a_13091_4943# trim[4] 6.64e-20
C10043 _084_ mask\[5\] 0.143f
C10044 a_448_6549# net22 0.171f
C10045 a_2368_9955# a_2787_9845# 8.23e-19
C10046 a_1000_12381# result[6] 9.22e-19
C10047 mask\[4\] a_5829_9839# 4.12e-19
C10048 net47 a_13256_9117# 8.83e-19
C10049 net46 a_14335_2442# 3.52e-20
C10050 a_395_6031# a_1007_6031# 0.00188f
C10051 _108_ a_14686_3017# 5.76e-19
C10052 net46 net8 0.041f
C10053 _040_ a_4775_6031# 8.12e-20
C10054 clknet_2_0__leaf_clk a_3830_6281# 8.17e-21
C10055 _095_ _060_ 3.3e-20
C10056 _129_ a_13557_7369# 1.98e-20
C10057 a_455_12533# result[6] 0.332f
C10058 a_6796_12381# net53 7.79e-20
C10059 a_7571_4943# _105_ 8.03e-20
C10060 a_9503_4399# a_9802_4007# 6.6e-19
C10061 a_6541_12021# a_6197_12015# 8.06e-20
C10062 a_5496_12131# net27 3.65e-20
C10063 _106_ a_8307_4719# 5.59e-19
C10064 clknet_2_2__leaf_clk a_11233_4405# 0.115f
C10065 a_911_4777# VPWR 0.228f
C10066 a_4871_8181# a_5535_8181# 0.0148f
C10067 a_4131_8207# _077_ 2.5e-20
C10068 cal_itt\[0\] a_11709_6273# 1.25e-20
C10069 _108_ a_9503_4399# 0.258f
C10070 _076_ a_5535_8181# 0.00552f
C10071 _078_ a_1679_10633# 0.00324f
C10072 a_4043_7093# _049_ 0.00262f
C10073 _063_ a_9099_3689# 2.94e-21
C10074 _017_ VPWR 0.42f
C10075 net4 a_8745_6895# 1.89e-21
C10076 _129_ net2 0.0365f
C10077 a_9802_4007# a_9369_3855# 2.12e-19
C10078 net4 clknet_2_0__leaf_clk 0.0188f
C10079 _072_ a_7001_7669# 0.134f
C10080 _005_ a_1651_7093# 4.73e-20
C10081 _112_ a_13975_3689# 0.00315f
C10082 state\[0\] a_2033_3317# 5.34e-19
C10083 a_7223_2465# a_7181_2589# 2.56e-19
C10084 net16 trim_val\[2\] 0.111f
C10085 a_12056_6031# _136_ 0.00705f
C10086 net43 net2 3.18e-20
C10087 net37 trimb[4] 0.00207f
C10088 cal_count\[3\] a_13441_6281# 3.69e-19
C10089 _048_ _118_ 3.3e-20
C10090 _100_ a_7021_4105# 8.93e-20
C10091 a_14894_3677# VPWR 8.45e-20
C10092 _068_ a_7001_7669# 2.12e-20
C10093 _108_ a_9369_3855# 0.0194f
C10094 net1 a_1867_3317# 3.65e-20
C10095 clknet_2_1__leaf_clk net51 0.331f
C10096 _014_ a_2564_2589# 0.16f
C10097 net15 a_1835_11231# 9.71e-21
C10098 net7 VPWR 0.521f
C10099 a_816_7119# _004_ 1.79e-20
C10100 clknet_2_0__leaf_clk a_3303_7119# 0.0375f
C10101 a_7939_3855# _119_ 2.72e-19
C10102 a_13111_6031# a_13783_6183# 0.0163f
C10103 a_4775_6031# _048_ 5.1e-21
C10104 a_12520_7637# a_12430_7663# 9.35e-20
C10105 cal_itt\[2\] a_8301_8207# 0.0563f
C10106 net12 _072_ 0.00247f
C10107 state\[1\] a_2755_2601# 1.48e-19
C10108 a_7393_5193# _107_ 6.64e-19
C10109 clknet_2_1__leaf_clk a_4055_12015# 0.00144f
C10110 a_10787_1135# a_11374_1251# 8.01e-20
C10111 _092_ a_6210_4989# 0.0334f
C10112 _136_ _058_ 0.153f
C10113 _104_ a_8583_3317# 0.267f
C10114 clknet_2_0__leaf_clk a_911_7119# 7.75e-19
C10115 a_8298_2767# a_8912_2589# 8.5e-19
C10116 net13 net4 0.00859f
C10117 net27 result[7] 8.81e-19
C10118 net14 _080_ 0.00104f
C10119 _041_ net40 5.18e-22
C10120 clknet_2_3__leaf_clk a_11801_4373# 3e-20
C10121 a_9957_7663# VPWR 0.208f
C10122 a_5625_4943# VPWR 2.43e-19
C10123 _122_ _131_ 0.0065f
C10124 net9 a_13091_1141# 0.00213f
C10125 a_13825_5185# a_14281_4943# 4.2e-19
C10126 _002_ a_7263_7093# 2.36e-19
C10127 net12 a_4443_9295# 6.71e-21
C10128 _108_ a_9747_2527# 4.09e-21
C10129 a_6515_6794# _073_ 0.188f
C10130 net31 _129_ 1.41e-20
C10131 clknet_2_1__leaf_clk _003_ 3.91e-19
C10132 net42 a_7800_4631# 2.25e-19
C10133 a_6541_12021# a_6099_10633# 2.91e-21
C10134 a_8673_10625# _042_ 0.0184f
C10135 net43 net24 0.07f
C10136 net47 a_9871_10383# 6.57e-19
C10137 a_7088_7119# a_7262_5461# 4.15e-22
C10138 a_7263_7093# _050_ 5.67e-21
C10139 en_co_clk a_4308_4917# 0.00756f
C10140 a_7723_10143# a_8083_8181# 5.95e-21
C10141 a_4425_6031# VPWR 0.528f
C10142 net12 net52 4.96e-20
C10143 net47 a_10798_9295# 0.00227f
C10144 cal_count\[3\] _066_ 0.139f
C10145 _095_ a_4498_4373# 4.99e-19
C10146 a_7715_3285# _028_ 0.00369f
C10147 net40 a_9839_3615# 3.24e-21
C10148 _078_ _065_ 0.274f
C10149 _080_ a_395_7119# 1.26e-19
C10150 a_395_4405# net41 1.9e-20
C10151 a_448_7637# a_561_7119# 2.18e-19
C10152 _108_ _111_ 0.0474f
C10153 trim_mask\[3\] a_9007_2601# 5.37e-21
C10154 _014_ net1 1.44e-20
C10155 _107_ a_9503_4399# 0.0841f
C10156 net45 result[0] 3.23e-19
C10157 _036_ _037_ 2.57e-20
C10158 _063_ trim_val\[4\] 6.93e-21
C10159 net53 _041_ 0.106f
C10160 _078_ net23 0.0113f
C10161 calibrate a_6703_2197# 1.23e-19
C10162 mask\[7\] a_1493_11721# 0.0502f
C10163 a_3431_10933# a_4055_10927# 9.73e-19
C10164 net9 a_10851_1653# 1.72e-19
C10165 clknet_0_clk a_8473_5193# 7.06e-19
C10166 a_11116_8983# _053_ 1.01e-19
C10167 _023_ a_816_10205# 4.05e-19
C10168 _074_ a_5915_10927# 3.55e-20
C10169 _107_ a_9369_3855# 5.99e-19
C10170 _070_ a_9459_7895# 0.089f
C10171 a_1644_12533# _085_ 9.81e-20
C10172 net12 a_5931_4105# 0.00101f
C10173 net43 a_4883_6397# 1e-19
C10174 net18 a_11141_6031# 0.00307f
C10175 a_9595_1679# ctln[4] 3.44e-19
C10176 net44 _070_ 0.00138f
C10177 a_13783_6183# a_13825_6031# 0.0175f
C10178 _135_ a_13349_6031# 0.0439f
C10179 a_5087_3855# a_4815_3031# 6.11e-19
C10180 a_6793_8970# a_6173_7119# 3.16e-21
C10181 a_3868_7119# VPWR 0.297f
C10182 a_14983_9269# trimb[1] 7.14e-19
C10183 net9 _053_ 6.64e-20
C10184 a_1125_7663# net22 4.11e-19
C10185 a_1764_10383# VPWR 3.4e-19
C10186 _101_ _018_ 0.0498f
C10187 _060_ calibrate 0.0293f
C10188 net25 a_1677_9545# 0.021f
C10189 _099_ a_3123_3615# 5.48e-21
C10190 _086_ a_1461_10357# 3.17e-21
C10191 cal_count\[3\] a_7571_4943# 2.12e-20
C10192 _029_ a_13519_4007# 7.15e-20
C10193 a_4815_3031# a_4443_1679# 2.83e-20
C10194 cal_itt\[0\] a_10593_9295# 4.41e-19
C10195 a_2288_3677# clk 2.08e-19
C10196 net16 trim_mask\[0\] 0.0753f
C10197 _104_ a_7190_3855# 0.0544f
C10198 a_7310_2223# clk 0.00262f
C10199 _049_ a_9369_3855# 5.81e-20
C10200 a_13512_4943# VPWR 0.0829f
C10201 a_1660_11305# a_1476_10217# 8.34e-21
C10202 a_11435_2229# a_12169_2197# 0.0701f
C10203 a_1835_11231# net25 2.65e-21
C10204 net52 a_1651_10143# 3.73e-19
C10205 a_395_9845# _082_ 1.67e-19
C10206 a_11141_6031# a_12165_6031# 2.36e-20
C10207 _007_ a_448_9269# 0.0163f
C10208 _052_ a_6737_3855# 0.0542f
C10209 _052_ a_6941_2589# 5.97e-20
C10210 a_745_12021# result[6] 0.00342f
C10211 net47 a_12520_7637# 0.159f
C10212 net37 _130_ 0.0221f
C10213 mask\[7\] VPWR 0.736f
C10214 _085_ a_2828_12131# 1.59e-19
C10215 _110_ a_8583_3317# 0.0106f
C10216 net33 _113_ 4.06e-22
C10217 _039_ a_1129_6273# 0.00152f
C10218 _102_ a_1461_10357# 7.47e-19
C10219 _136_ a_13607_4943# 8.86e-19
C10220 _074_ a_1467_7923# 1.42e-19
C10221 _078_ a_2225_7663# 1.34e-20
C10222 _064_ a_10188_4105# 0.00196f
C10223 mask\[7\] a_1769_12393# 6.99e-20
C10224 a_6485_8181# net51 0.144f
C10225 net37 a_14335_4020# 1.32e-20
C10226 clknet_0_clk a_8583_3317# 0.0028f
C10227 a_14377_7983# VPWR 9.42e-19
C10228 clknet_2_0__leaf_clk ctln[1] 4.53e-21
C10229 _070_ en_co_clk 4.53e-21
C10230 a_561_6031# a_1493_5487# 1.15e-19
C10231 _078_ _016_ 3.68e-20
C10232 a_3977_10217# VPWR 4.26e-20
C10233 a_12546_9129# VPWR 5.47e-20
C10234 _094_ a_5081_4943# 0.0481f
C10235 net43 a_1129_6273# 3.38e-19
C10236 net24 a_2857_7637# 0.00181f
C10237 a_4167_6575# _034_ 0.109f
C10238 _045_ _078_ 7.44e-19
C10239 _070_ a_8386_8457# 0.0149f
C10240 net45 a_7010_3311# 2.59e-20
C10241 a_15023_10927# trimb[0] 0.339f
C10242 _101_ mask\[1\] 0.407f
C10243 trim_mask\[0\] a_10699_3311# 6.95e-19
C10244 net34 _058_ 7.39e-20
C10245 _094_ net55 0.323f
C10246 net46 a_13703_4943# 9.54e-19
C10247 a_13059_4631# a_13233_4737# 0.00658f
C10248 a_12148_4777# a_12310_4399# 0.00645f
C10249 _063_ a_8745_4943# 2.79e-19
C10250 mask\[2\] a_4609_9295# 0.0128f
C10251 a_1497_8725# net45 1.46e-19
C10252 _112_ trim_val\[1\] 0.00578f
C10253 a_13415_2442# net48 1.93e-19
C10254 net6 rstn 0.00668f
C10255 _078_ a_4696_8207# 8.98e-19
C10256 _103_ VPWR 0.255f
C10257 a_3557_5193# a_3365_4943# 0.00137f
C10258 a_395_7119# a_1651_7093# 0.0436f
C10259 a_561_7119# a_911_7119# 0.23f
C10260 a_6909_10933# a_7164_11293# 0.0642f
C10261 a_395_9845# a_1007_10217# 0.00188f
C10262 a_8949_9537# a_8839_9661# 0.0977f
C10263 a_9471_9269# a_9296_9295# 0.234f
C10264 a_8731_9295# a_8636_9295# 0.0498f
C10265 _064_ trim_mask\[3\] 0.394f
C10266 net51 a_6007_7119# 0.00529f
C10267 net37 a_15023_2767# 1.08e-19
C10268 en_co_clk _090_ 0.00578f
C10269 _099_ a_3530_4765# 0.00187f
C10270 a_3388_4631# _097_ 0.0806f
C10271 net14 a_937_4105# 0.00183f
C10272 mask\[5\] a_6181_10383# 9.26e-19
C10273 _053_ a_10188_4105# 5.41e-22
C10274 a_10975_4105# a_11067_3017# 1.26e-20
C10275 _064_ a_10689_2543# 8.77e-19
C10276 a_10903_7261# VPWR 0.501f
C10277 _062_ _064_ 0.516f
C10278 cal_itt\[2\] a_7088_7119# 1.91e-20
C10279 a_11859_3689# VPWR 0.209f
C10280 net2 a_14379_6397# 5.73e-21
C10281 a_6173_7119# net30 2.7e-20
C10282 clknet_0_clk a_4680_6031# 6.06e-21
C10283 clknet_2_1__leaf_clk a_763_8757# 0.264f
C10284 _101_ a_1387_8751# 1.95e-20
C10285 calibrate a_7939_3855# 1.26e-19
C10286 net43 a_4801_10159# 3.33e-19
C10287 a_7824_11305# a_8215_9295# 1.54e-20
C10288 _041_ _071_ 1.8e-20
C10289 _100_ a_6197_4399# 6.37e-19
C10290 trim_mask\[3\] a_10851_1653# 0.0277f
C10291 cal_count\[2\] a_14282_7119# 8.88e-19
C10292 mask\[3\] a_5055_9295# 2.74e-19
C10293 cal_itt\[2\] _063_ 0.36f
C10294 calibrate a_4498_4373# 2.97e-19
C10295 mask\[6\] a_4621_11305# 8.65e-19
C10296 _078_ _023_ 3.55e-19
C10297 _086_ a_745_10933# 0.00579f
C10298 a_13415_2442# a_13091_1141# 6.05e-21
C10299 a_6007_7119# _003_ 0.169f
C10300 a_15023_1679# trim[2] 8.02e-19
C10301 _114_ a_13825_1109# 0.00204f
C10302 mask\[7\] net27 0.0419f
C10303 a_11845_4765# VPWR 2.51e-19
C10304 _070_ a_8091_7967# 0.00139f
C10305 net45 a_3148_4399# 0.00113f
C10306 a_6743_10933# _021_ 0.318f
C10307 _131_ comp 0.00527f
C10308 clknet_2_1__leaf_clk net26 0.105f
C10309 cal_itt\[1\] a_9919_6614# 1.1e-19
C10310 a_10405_9295# a_10593_9295# 0.152f
C10311 a_1129_4373# a_1173_4765# 3.69e-19
C10312 net46 a_13459_3317# 0.665f
C10313 a_911_4777# a_1007_4777# 0.0138f
C10314 mask\[0\] a_3977_7119# 8.79e-19
C10315 net13 a_4055_10927# 5.88e-19
C10316 net4 a_2948_3689# 0.00387f
C10317 a_1313_10901# a_1203_10927# 0.0977f
C10318 a_745_10933# _102_ 0.00182f
C10319 net43 a_4993_6273# 6.51e-20
C10320 _136_ a_11488_4765# 5.57e-19
C10321 net44 a_4349_8449# 0.159f
C10322 clknet_2_2__leaf_clk a_14540_3689# 2.36e-21
C10323 net15 a_2971_8457# 0.0109f
C10324 a_9662_3855# VPWR 0.00298f
C10325 _053_ _062_ 0.162f
C10326 a_7140_2223# VPWR 7.89e-19
C10327 _121_ VPWR 0.396f
C10328 cal_itt\[0\] a_9677_8457# 4.74e-19
C10329 a_15259_7637# clkc 5.42e-19
C10330 cal_count\[0\] net2 1.05e-19
C10331 net55 a_4617_3855# 0.00122f
C10332 _065_ a_7001_7669# 7.67e-20
C10333 a_8105_10383# VPWR 0.274f
C10334 _053_ a_10138_5807# 0.00139f
C10335 a_9595_1679# clk 1.35e-21
C10336 net45 a_1019_4399# 0.0122f
C10337 net46 _109_ 3.12e-20
C10338 trim_mask\[0\] a_7019_4407# 9.29e-20
C10339 a_11244_9661# _041_ 3.51e-19
C10340 _123_ a_13279_7119# 0.0215f
C10341 _003_ _092_ 4.53e-21
C10342 a_12056_6031# cal_count\[3\] 0.055f
C10343 a_5515_6005# _051_ 7.17e-19
C10344 a_13307_1707# _114_ 0.18f
C10345 _042_ a_2961_9545# 0.0466f
C10346 net26 a_2368_9955# 8.47e-20
C10347 a_1679_10633# a_1651_10143# 2.28e-19
C10348 _122_ a_11297_7119# 6.43e-19
C10349 _095_ a_4175_4943# 1.35e-20
C10350 _006_ a_1007_7119# 1.56e-20
C10351 net16 _030_ 0.00367f
C10352 a_10383_7093# a_10621_7119# 0.0074f
C10353 a_11098_6691# en_co_clk 8.78e-19
C10354 a_2857_7637# a_4677_7882# 4.1e-19
C10355 net12 _065_ 0.0165f
C10356 _020_ a_6445_10383# 0.00133f
C10357 _094_ a_5166_5193# 0.0159f
C10358 _108_ a_14981_4020# 0.00185f
C10359 a_2283_4020# net41 1.43e-19
C10360 a_9503_4399# trim_mask\[4\] 5.68e-19
C10361 a_9572_2601# VPWR 0.318f
C10362 a_6261_11247# VPWR 7.67e-19
C10363 a_8215_9295# a_10239_9295# 1.71e-19
C10364 _059_ _090_ 0.0303f
C10365 net4 _028_ 0.0109f
C10366 net43 a_3208_7119# 2.77e-19
C10367 _010_ a_4621_12393# 4.2e-20
C10368 cal_count\[3\] _058_ 0.00167f
C10369 a_8935_6895# a_8298_5487# 2.98e-21
C10370 _123_ _041_ 0.0407f
C10371 net2 a_6741_7361# 3.19e-21
C10372 _060_ _015_ 0.0686f
C10373 _002_ _071_ 3.17e-21
C10374 _122_ _036_ 0.00237f
C10375 trim_mask\[4\] a_7942_2223# 1.05e-19
C10376 a_9478_4105# a_9662_3855# 1.91e-19
C10377 trim_mask\[4\] a_9369_3855# 9.91e-21
C10378 _065_ a_5340_6031# 9.33e-19
C10379 _058_ a_12586_3311# 3.74e-20
C10380 a_1129_6273# a_1173_6031# 3.69e-19
C10381 a_911_6031# a_1007_6031# 0.0138f
C10382 _049_ a_3748_6281# 0.0134f
C10383 _003_ cal_itt\[3\] 2.56e-19
C10384 a_14347_1439# a_15023_1135# 9e-19
C10385 net31 cal_count\[0\] 6.25e-20
C10386 a_448_7637# a_1467_7923# 1.78e-20
C10387 a_11343_3317# a_13459_3317# 1.45e-19
C10388 _129_ a_14733_7983# 2.57e-19
C10389 trim_mask\[1\] a_14604_3017# 0.105f
C10390 _063_ net55 5.98e-19
C10391 a_929_8757# _081_ 0.00817f
C10392 _005_ a_395_6031# 1.8e-20
C10393 _127_ a_14565_9295# 3.98e-19
C10394 a_9471_9269# a_9463_8725# 0.0139f
C10395 a_6541_12021# ctlp[6] 1.31e-19
C10396 net46 a_12169_2197# 0.166f
C10397 a_763_8757# a_1953_9129# 2.56e-19
C10398 mask\[1\] a_6515_8534# 2.87e-20
C10399 _034_ _094_ 0.0183f
C10400 _095_ a_4576_3427# 5.79e-20
C10401 net43 a_4222_10205# 0.00438f
C10402 net13 mask\[4\] 0.0131f
C10403 net43 result[1] 1.33e-19
C10404 a_14471_591# VPWR 0.301f
C10405 clknet_0_clk a_4425_6031# 0.0128f
C10406 _101_ _041_ 0.0098f
C10407 a_6375_12021# a_6796_12381# 0.0931f
C10408 clknet_2_2__leaf_clk net8 0.0058f
C10409 net15 a_4131_8207# 6.38e-19
C10410 net37 trim[4] 0.00207f
C10411 _103_ _104_ 0.0652f
C10412 net27 a_8105_10383# 1.6e-19
C10413 mask\[3\] net24 0.0026f
C10414 trim_mask\[4\] a_9747_2527# 4.53e-19
C10415 a_1867_3317# a_2143_2229# 5.3e-21
C10416 net44 a_5055_9295# 0.00274f
C10417 trim_val\[3\] a_10569_1109# 0.185f
C10418 a_15023_1679# a_15023_1135# 0.00787f
C10419 a_9889_6873# VPWR 0.21f
C10420 a_3273_4943# VPWR 0.455f
C10421 mask\[6\] a_2787_9845# 6.01e-19
C10422 net55 _096_ 0.13f
C10423 net47 a_13142_8359# 0.00916f
C10424 _077_ a_5691_7637# 0.0119f
C10425 _112_ a_12424_3689# 1.1e-20
C10426 mask\[5\] a_7164_11293# 7.84e-20
C10427 net18 a_10195_1354# 8.68e-19
C10428 mask\[0\] a_1476_6031# 8.21e-19
C10429 a_8307_6575# net42 1.25e-19
C10430 a_448_11445# result[5] 0.158f
C10431 a_13142_7271# a_14422_7093# 4.16e-20
C10432 a_4443_9295# _040_ 1.61e-20
C10433 a_7001_7669# _067_ 6.85e-20
C10434 _080_ VPWR 0.292f
C10435 a_13825_1109# VPWR 0.223f
C10436 net51 a_5547_5603# 8.31e-21
C10437 a_13933_6281# clkc 7.52e-20
C10438 clknet_0_clk a_3868_7119# 0.0083f
C10439 a_2857_7637# a_3208_7119# 6.83e-19
C10440 net12 a_4696_8207# 7.6e-22
C10441 net30 a_7800_4631# 0.00138f
C10442 net52 _040_ 0.153f
C10443 a_13919_8751# net2 6.55e-20
C10444 _074_ _011_ 0.1f
C10445 _089_ a_5931_4105# 0.113f
C10446 a_7190_3855# net41 1.75e-22
C10447 a_10329_1921# trim_val\[3\] 4.26e-20
C10448 a_10676_1679# a_10838_2045# 0.00645f
C10449 a_10111_1679# a_10373_1679# 0.00171f
C10450 net13 _053_ 5.12e-19
C10451 _094_ a_3830_6281# 7.8e-19
C10452 a_14715_3615# _055_ 0.0274f
C10453 a_14335_7895# a_14063_7093# 4.73e-20
C10454 net33 a_14347_9480# 0.00618f
C10455 mask\[4\] a_4864_9295# 8.95e-19
C10456 a_12992_8751# a_13562_8751# 0.111f
C10457 a_13142_8725# _041_ 0.0204f
C10458 _015_ a_4864_1679# 0.16f
C10459 net45 a_3521_7361# 7.31e-20
C10460 _025_ a_11601_2229# 9.52e-21
C10461 net18 _032_ 4.23e-19
C10462 a_6927_12559# a_8820_12533# 3.07e-21
C10463 a_15023_12015# trimb[0] 6.66e-20
C10464 clknet_2_1__leaf_clk a_2961_9295# 1.25e-19
C10465 _026_ a_11601_2229# 0.228f
C10466 a_6906_2355# a_7223_2465# 0.102f
C10467 a_6703_2197# a_7184_2339# 0.0424f
C10468 a_3868_10217# a_4655_10071# 7.15e-19
C10469 _095_ a_3557_5193# 0.00135f
C10470 a_2857_5461# a_3365_4943# 2.55e-19
C10471 net4 a_9621_8029# 4.12e-19
C10472 _029_ a_14526_4943# 6.53e-22
C10473 net46 a_15023_1135# 8.6e-19
C10474 _005_ net30 5.05e-20
C10475 clknet_2_3__leaf_clk cal_itt\[0\] 0.042f
C10476 a_9296_9295# _069_ 0.00103f
C10477 a_13307_1707# VPWR 0.226f
C10478 _014_ a_2143_2229# 0.17f
C10479 _076_ _075_ 0.0525f
C10480 a_8105_10383# a_8455_10383# 0.217f
C10481 a_6099_10633# _042_ 0.0295f
C10482 a_7939_10383# a_9195_10357# 0.0436f
C10483 a_5455_4943# a_5081_4943# 0.0143f
C10484 net8 ctln[2] 0.00686f
C10485 net23 result[2] 4.23e-19
C10486 _081_ clknet_2_0__leaf_clk 2.17e-20
C10487 a_8072_11721# a_8360_10383# 1.63e-20
C10488 trim_mask\[1\] a_9839_3615# 3.51e-19
C10489 _078_ a_3597_10933# 7.8e-19
C10490 _020_ net47 0.00472f
C10491 _095_ a_1830_4765# 1.1e-19
C10492 net35 a_14972_5193# 2.12e-19
C10493 a_816_6031# VPWR 0.0834f
C10494 a_10785_1679# ctln[4] 6.4e-20
C10495 net2 a_9459_7895# 3.03e-20
C10496 a_14347_4917# _058_ 0.00241f
C10497 state\[1\] a_2309_2229# 1.92e-19
C10498 net55 a_5455_4943# 5.75e-19
C10499 net15 net30 0.429f
C10500 net19 a_8583_3317# 0.0145f
C10501 net44 net2 0.00953f
C10502 trim_val\[3\] a_11374_1251# 1.12e-19
C10503 _037_ a_10586_7371# 7.95e-20
C10504 a_8298_2767# _027_ 0.0137f
C10505 a_6885_8372# VPWR 0.261f
C10506 _051_ a_4815_3031# 0.0381f
C10507 _108_ trim_mask\[2\] 0.167f
C10508 net22 a_1830_6031# 5.12e-19
C10509 _097_ a_3123_3615# 5.84e-19
C10510 _103_ _110_ 4.07e-20
C10511 _058_ _119_ 4.32e-19
C10512 _010_ _022_ 5.28e-19
C10513 _028_ a_7689_2589# 0.00129f
C10514 clknet_2_0__leaf_clk a_455_5747# 0.0847f
C10515 clknet_0_clk _103_ 0.00673f
C10516 _092_ _088_ 6.57e-20
C10517 net46 a_10219_2045# 0.0168f
C10518 a_10781_5487# trim_mask\[1\] 2.79e-21
C10519 _104_ a_9572_2601# 5.9e-20
C10520 a_7351_8041# net30 8.41e-21
C10521 _092_ a_7262_5461# 0.018f
C10522 _049_ a_4308_4917# 0.00826f
C10523 net14 a_395_6031# 0.0096f
C10524 a_9317_3285# a_9099_3689# 0.21f
C10525 a_8749_3317# a_9839_3615# 0.0424f
C10526 a_3597_12021# a_6197_12015# 6.1e-21
C10527 _106_ clk 1.91e-20
C10528 a_1677_9545# VPWR 0.264f
C10529 a_14422_7093# a_14870_7369# 1.95e-19
C10530 _131_ a_14199_7369# 8.44e-19
C10531 a_13715_1135# VPWR 0.155f
C10532 a_3891_4943# a_3817_4697# 9.76e-19
C10533 a_8298_5487# _066_ 5.74e-19
C10534 net26 result[4] 0.00579f
C10535 _096_ _093_ 0.119f
C10536 trim_mask\[2\] a_10655_2932# 0.0345f
C10537 _135_ a_13441_6281# 0.00232f
C10538 a_13783_6183# _136_ 0.144f
C10539 clknet_0_clk a_10903_7261# 1.69e-20
C10540 net45 _095_ 0.0222f
C10541 a_9074_9955# VPWR 0.00228f
C10542 a_7210_5807# a_7019_4407# 1.76e-20
C10543 net2 clk 2.48e-20
C10544 calibrate a_4576_3427# 5.21e-20
C10545 net2 en_co_clk 0.09f
C10546 a_911_10217# _082_ 9.92e-20
C10547 _043_ a_8215_9295# 0.00115f
C10548 _106_ a_9084_4515# 0.149f
C10549 _048_ a_5931_4105# 0.00561f
C10550 a_1835_11231# VPWR 0.43f
C10551 trim_mask\[4\] a_10676_1679# 4.24e-19
C10552 a_4443_9295# a_5177_9537# 0.0532f
C10553 a_11141_6031# VPWR 0.262f
C10554 a_1651_7093# VPWR 0.42f
C10555 a_6519_3829# a_6737_3855# 0.0326f
C10556 a_1203_12015# a_1313_10901# 1.09e-20
C10557 a_12077_3285# a_11967_3311# 0.0977f
C10558 trim_mask\[3\] a_10689_2223# 0.0193f
C10559 a_8105_10383# a_8381_9295# 7.45e-21
C10560 a_7939_10383# a_8949_9537# 1.76e-20
C10561 _092_ a_6519_4631# 3.06e-20
C10562 net2 a_8386_8457# 7.04e-20
C10563 a_14715_3615# trim_val\[2\] 1.8e-20
C10564 _028_ a_9007_2601# 1.48e-21
C10565 net40 a_10005_6031# 4.22e-19
C10566 net44 net24 2.51e-21
C10567 clknet_2_0__leaf_clk a_3891_4943# 1.98e-21
C10568 _101_ a_3615_8207# 7.48e-21
C10569 _132_ a_14870_7369# 8.78e-19
C10570 a_11141_6031# a_12218_6397# 1.46e-19
C10571 net46 a_11599_6397# 0.0122f
C10572 a_3521_9813# a_3977_10217# 4.2e-19
C10573 a_3303_10217# a_3565_10205# 0.00171f
C10574 net9 _057_ 0.0755f
C10575 _027_ a_11951_2601# 1.42e-20
C10576 a_579_10933# a_1476_10217# 4.22e-22
C10577 net28 net52 0.00395f
C10578 a_395_7119# a_395_6031# 5.57e-19
C10579 _084_ net44 1.46e-19
C10580 a_855_4105# cal 0.00651f
C10581 net52 a_5177_9537# 3.59e-21
C10582 a_10903_7261# a_10699_5487# 2.43e-20
C10583 a_11856_2589# a_12047_2601# 4.61e-19
C10584 _096_ a_2865_4460# 1.46e-19
C10585 net3 a_2601_3285# 2.15e-19
C10586 a_2787_7119# a_3303_7119# 0.106f
C10587 a_2953_7119# a_3521_7361# 0.174f
C10588 a_12323_4703# a_12599_3615# 1.65e-19
C10589 a_579_10933# _007_ 0.00105f
C10590 _061_ a_14972_5193# 2.27e-20
C10591 net33 a_14870_7369# 3.68e-19
C10592 a_1099_12533# a_579_10933# 4.86e-21
C10593 cal_itt\[3\] a_7262_5461# 2.17e-19
C10594 en_co_clk a_3667_3829# 9.44e-19
C10595 state\[2\] a_7800_4631# 8.42e-20
C10596 a_15023_6031# trim[1] 8.91e-21
C10597 clknet_2_3__leaf_clk trim_mask\[0\] 0.324f
C10598 _110_ a_9662_3855# 0.00264f
C10599 _097_ a_3530_4765# 2.88e-19
C10600 a_1644_12533# a_745_12021# 0.00864f
C10601 _074_ clknet_2_1__leaf_clk 0.473f
C10602 a_8749_3317# a_9207_3311# 0.0346f
C10603 _033_ clk 2.05e-20
C10604 net18 net30 5.08e-20
C10605 trim_mask\[2\] a_12516_2601# 0.00264f
C10606 a_937_4105# VPWR 0.179f
C10607 a_12631_12559# VPWR 0.301f
C10608 clknet_0_clk _121_ 0.0132f
C10609 a_7939_3855# a_7184_2339# 1.18e-21
C10610 a_911_10217# a_1007_10217# 0.0138f
C10611 a_1129_9813# a_1173_10205# 3.69e-19
C10612 clknet_2_3__leaf_clk a_10405_9295# 0.352f
C10613 a_11801_4373# a_11691_4399# 0.0977f
C10614 _058_ a_11679_4777# 9.54e-19
C10615 _051_ a_5087_3855# 1.21e-20
C10616 _078_ _004_ 1.57e-20
C10617 _063_ a_9595_5193# 0.045f
C10618 a_10055_2767# a_10195_1354# 3e-19
C10619 a_13142_7271# _136_ 0.00209f
C10620 clknet_2_2__leaf_clk a_13703_4943# 5.75e-19
C10621 a_13825_5185# a_14172_4943# 0.0512f
C10622 a_13091_4943# a_13512_4943# 0.0902f
C10623 net44 a_4883_6397# 0.0129f
C10624 net31 en_co_clk 2.05e-20
C10625 a_5578_12131# VPWR 0.00138f
C10626 _052_ a_6703_2197# 2.16e-19
C10627 a_12169_2197# a_12059_2223# 0.0977f
C10628 a_11601_2229# _031_ 1.39e-19
C10629 net45 a_7617_2589# 0.00316f
C10630 _111_ a_12723_4943# 0.19f
C10631 _051_ a_4443_1679# 9.02e-20
C10632 _050_ a_8749_3317# 9.32e-20
C10633 _050_ _060_ 2.31e-19
C10634 a_8215_9295# a_9471_9269# 0.0436f
C10635 calibrate a_1638_4399# 4.47e-19
C10636 _000_ a_8731_9295# 0.00213f
C10637 mask\[4\] a_9020_10383# 0.02f
C10638 clknet_2_1__leaf_clk a_1279_9129# 5.3e-20
C10639 state\[1\] _089_ 3.47e-20
C10640 a_9003_3829# a_9099_3689# 0.00228f
C10641 _074_ a_2368_9955# 4.36e-21
C10642 _136_ a_14181_6031# 4.21e-19
C10643 a_1476_4777# _014_ 3.11e-19
C10644 a_9463_8725# _069_ 0.0024f
C10645 net2 a_8091_7967# 1.58e-19
C10646 _110_ a_9572_2601# 0.0152f
C10647 a_937_3855# valid 1.39e-19
C10648 _090_ _107_ 0.00633f
C10649 _124_ a_11116_8983# 0.0999f
C10650 net14 net30 0.0107f
C10651 a_10747_8970# _123_ 2.48e-19
C10652 cal_itt\[2\] a_6007_7119# 2.48e-21
C10653 state\[1\] a_4609_1679# 2.44e-21
C10654 net20 a_7631_12319# 9.79e-19
C10655 net44 a_5878_9295# 0.00384f
C10656 net15 state\[0\] 0.0042f
C10657 _081_ a_561_7119# 1.5e-21
C10658 net42 VPWR 0.687f
C10659 _052_ a_8749_3317# 1.27e-20
C10660 _047_ _055_ 3.3e-20
C10661 a_9463_8725# a_8022_7119# 2.1e-19
C10662 a_4901_2773# VPWR 1.46e-20
C10663 cal_count\[2\] a_13557_7369# 1.79e-19
C10664 _078_ a_6888_10205# 1.55e-20
C10665 a_10655_2932# a_9595_1679# 2.42e-20
C10666 a_4883_6397# en_co_clk 1.93e-19
C10667 a_395_9845# a_1476_10217# 0.102f
C10668 net4 _063_ 0.0356f
C10669 mask\[1\] a_3053_8207# 7.12e-19
C10670 _010_ a_4512_12393# 3.47e-19
C10671 _078_ net12 0.111f
C10672 a_448_10357# net26 0.18f
C10673 _060_ _098_ 3.68e-19
C10674 a_4091_5309# VPWR 0.31f
C10675 trim_val\[2\] a_14099_1929# 0.0171f
C10676 a_14335_2442# net8 4.41e-20
C10677 a_395_9845# _007_ 0.169f
C10678 _115_ a_13393_1707# 5.76e-19
C10679 net16 _133_ 0.0261f
C10680 a_561_4405# a_855_4105# 9.55e-19
C10681 _049_ _090_ 0.385f
C10682 _090_ a_3388_4631# 0.192f
C10683 a_15023_9839# a_14983_9269# 0.00114f
C10684 net2 cal_count\[2\] 0.244f
C10685 a_561_7119# a_455_5747# 1.86e-20
C10686 a_11059_7356# _038_ 2.52e-20
C10687 a_10990_7485# a_10975_6031# 9.3e-20
C10688 a_14422_7093# _131_ 0.253f
C10689 _130_ a_14788_7369# 0.175f
C10690 _101_ a_3249_9295# 0.00172f
C10691 a_3388_4631# a_3847_4438# 6.64e-19
C10692 cal_itt\[2\] _092_ 0.0943f
C10693 _065_ _040_ 2.39e-19
C10694 clknet_2_2__leaf_clk a_13459_3317# 0.235f
C10695 _054_ clk 0.00996f
C10696 trim_mask\[0\] a_14715_3615# 2.4e-20
C10697 _078_ a_6983_10217# 4.13e-20
C10698 mask\[4\] a_8731_9295# 0.0017f
C10699 a_15289_7119# VPWR 4.45e-20
C10700 _111_ a_13059_4631# 0.109f
C10701 a_10688_9295# net2 2.54e-20
C10702 trim_mask\[3\] _057_ 0.00172f
C10703 _108_ net50 0.13f
C10704 net23 _040_ 0.0546f
C10705 net4 _096_ 3.61e-21
C10706 net43 a_8083_8181# 0.00122f
C10707 net45 calibrate 0.158f
C10708 _122_ a_11479_9117# 0.00369f
C10709 _048_ a_7527_4631# 0.0748f
C10710 a_10239_9295# _041_ 4.85e-19
C10711 _132_ _131_ 0.119f
C10712 net16 a_14236_8457# 5.02e-19
C10713 a_8827_9295# cal_itt\[0\] 1.44e-19
C10714 _050_ a_7939_3855# 0.0108f
C10715 a_745_12021# a_1000_12381# 0.0642f
C10716 a_6316_5193# a_6566_5193# 0.149f
C10717 a_6519_4631# a_6737_4719# 0.0326f
C10718 clknet_2_2__leaf_clk _109_ 0.00148f
C10719 a_5915_10927# mask\[4\] 2.19e-19
C10720 net33 _131_ 0.00541f
C10721 _048_ state\[1\] 6.16e-19
C10722 _095_ a_6316_5193# 2.97e-20
C10723 a_2857_5461# _095_ 0.122f
C10724 _050_ a_4498_4373# 6.01e-21
C10725 a_9003_3829# trim_val\[4\] 0.00958f
C10726 net50 a_10655_2932# 6.72e-19
C10727 _078_ a_1651_10143# 0.00703f
C10728 _053_ _028_ 2.45e-19
C10729 net46 _112_ 0.00936f
C10730 cal_itt\[1\] a_9957_7663# 0.00924f
C10731 a_1476_7119# _039_ 0.00137f
C10732 a_2479_3689# VPWR 1.96e-19
C10733 _110_ a_13825_1109# 6.43e-21
C10734 cal_itt\[2\] cal_itt\[3\] 0.00647f
C10735 a_8491_2229# VPWR 0.429f
C10736 mask\[0\] _039_ 0.0319f
C10737 net47 a_12916_8751# 4.53e-19
C10738 net47 a_10975_6031# 3.98e-21
C10739 _052_ a_7939_3855# 4.28e-20
C10740 _010_ _046_ 9.53e-19
C10741 _067_ _091_ 0.00473f
C10742 _062_ a_10245_5193# 2.94e-21
C10743 _134_ trim_val\[0\] 1.07e-20
C10744 net43 a_1660_11305# 0.237f
C10745 _065_ _048_ 0.0175f
C10746 net30 a_11023_5108# 2.94e-19
C10747 net43 a_1476_7119# 0.264f
C10748 _015_ a_4576_3427# 0.00565f
C10749 mask\[6\] net26 1.39e-19
C10750 net43 mask\[0\] 0.601f
C10751 a_4864_1679# a_5055_1679# 4.61e-19
C10752 net44 a_4993_6273# 0.167f
C10753 net24 a_1184_9117# 0.0164f
C10754 a_8022_7119# a_10383_7093# 1.75e-20
C10755 a_15083_4659# clkc 4.89e-21
C10756 a_1203_10927# a_561_9845# 2.21e-20
C10757 a_3891_4943# a_4091_4943# 8e-19
C10758 clknet_2_3__leaf_clk a_8307_4943# 1.87e-19
C10759 _098_ a_4498_4373# 6.57e-21
C10760 _011_ a_1835_12319# 4.1e-20
C10761 _025_ _026_ 0.00206f
C10762 a_579_12021# a_1660_12393# 0.102f
C10763 a_395_6031# a_2313_6183# 3.94e-21
C10764 net51 _073_ 2.67e-20
C10765 _063_ a_10586_7371# 0.00103f
C10766 _053_ _037_ 0.00216f
C10767 _110_ a_13307_1707# 0.084f
C10768 mask\[5\] a_6099_10633# 0.112f
C10769 net16 _129_ 0.791f
C10770 _092_ a_5081_4943# 0.00256f
C10771 clknet_2_2__leaf_clk a_12169_2197# 4.82e-20
C10772 a_12625_2601# VPWR 6.3e-20
C10773 a_3840_8867# VPWR 0.168f
C10774 a_8307_6575# net30 0.00291f
C10775 cal_count\[1\] net2 0.914f
C10776 mask\[7\] a_1822_10927# 1.46e-19
C10777 _078_ result[2] 4.7e-20
C10778 _092_ net55 0.222f
C10779 net50 _107_ 4.2e-20
C10780 _065_ a_11599_6397# 9.16e-19
C10781 a_4775_6031# a_5037_6031# 0.00171f
C10782 a_2971_8457# VPWR 0.217f
C10783 a_4993_6273# en_co_clk 0.00551f
C10784 a_5340_6031# a_5502_6397# 0.00645f
C10785 _045_ a_3431_12021# 9.7e-21
C10786 clknet_2_0__leaf_clk a_3781_8207# 0.00308f
C10787 _040_ a_4696_8207# 0.0347f
C10788 trim_mask\[4\] a_7310_2223# 5.6e-19
C10789 _119_ a_8657_2229# 2.15e-19
C10790 _042_ clknet_2_3__leaf_clk 1.61e-20
C10791 a_4959_9295# a_5423_9011# 0.00358f
C10792 a_4886_4399# VPWR 0.00452f
C10793 net39 trimb[2] 0.00735f
C10794 a_561_9845# a_929_8757# 8.2e-21
C10795 trim_val\[0\] a_13915_4399# 0.00926f
C10796 clknet_2_0__leaf_clk a_395_4405# 0.271f
C10797 net43 _079_ 2.56e-19
C10798 _003_ _073_ 0.00241f
C10799 net18 a_11030_1679# 3.94e-19
C10800 _112_ a_11343_3317# 2.47e-21
C10801 _042_ a_395_9845# 1.81e-20
C10802 a_11803_10383# net9 6.92e-19
C10803 net46 net10 3.81e-20
C10804 net13 a_5221_1679# 5.87e-19
C10805 a_2309_2229# a_2755_2601# 2.28e-19
C10806 cal_count\[3\] a_13783_6183# 3.02e-19
C10807 a_12056_6031# _135_ 2.01e-19
C10808 net42 _104_ 1.36e-20
C10809 a_11488_4765# a_11679_4777# 4.61e-19
C10810 clknet_2_1__leaf_clk _083_ 0.0112f
C10811 net20 a_8072_11721# 1.58e-20
C10812 a_11764_3677# VPWR 0.0795f
C10813 net29 _023_ 1.43e-21
C10814 a_6835_7669# a_7569_7637# 0.0535f
C10815 _106_ a_9802_4007# 0.00751f
C10816 _108_ a_14604_2339# 0.0279f
C10817 _101_ a_2019_9055# 8.96e-19
C10818 trim_mask\[4\] trim_mask\[2\] 0.014f
C10819 a_10195_1354# VPWR 0.261f
C10820 net7 a_3063_591# 0.173f
C10821 net13 a_3781_8207# 0.00871f
C10822 _074_ result[4] 2.42e-19
C10823 a_11016_6691# _038_ 0.00282f
C10824 _108_ _106_ 0.174f
C10825 net52 a_2143_7663# 0.192f
C10826 a_4165_10901# mask\[2\] 1.27e-19
C10827 net14 a_1585_6031# 2.97e-20
C10828 _135_ _058_ 1.25e-19
C10829 mask\[0\] a_2857_7637# 3.73e-19
C10830 _072_ a_8025_8041# 5.94e-21
C10831 net2 _108_ 4.09e-20
C10832 a_13459_3317# a_14540_3689# 0.102f
C10833 _030_ a_14715_3615# 4.61e-20
C10834 a_11545_9049# _041_ 0.0215f
C10835 net12 a_7001_7669# 3.97e-19
C10836 a_11987_8757# a_13562_8751# 2.39e-19
C10837 _036_ a_12992_8751# 2.02e-20
C10838 mask\[1\] net45 0.124f
C10839 net12 ctln[7] 0.00247f
C10840 a_3748_6281# a_3529_6281# 6.46e-21
C10841 net46 a_12121_3677# 0.00371f
C10842 _018_ a_3868_10217# 2.29e-21
C10843 a_2787_9845# a_4655_10071# 1.74e-20
C10844 a_7916_8041# a_9957_7663# 8.6e-23
C10845 _108_ a_14193_3285# 0.00569f
C10846 a_2225_7983# VPWR 6.05e-19
C10847 trim_mask\[0\] _047_ 2.97e-19
C10848 a_2313_6183# net30 0.00208f
C10849 _066_ a_10781_5487# 0.0697f
C10850 clknet_2_1__leaf_clk a_3303_7119# 6.88e-19
C10851 _032_ VPWR 0.398f
C10852 clknet_2_1__leaf_clk a_8360_10383# 1.99e-19
C10853 a_11141_6031# a_10699_5487# 4.26e-20
C10854 calibrate a_6316_5193# 0.0297f
C10855 net46 a_11583_4777# 0.156f
C10856 a_3667_3829# a_3399_2527# 7.1e-20
C10857 _125_ a_14552_9071# 0.0015f
C10858 a_2857_5461# calibrate 7e-21
C10859 _095_ a_6210_4989# 1.94e-20
C10860 net4 a_9761_1679# 0.00102f
C10861 a_3425_11721# a_3511_11471# 2.42e-19
C10862 a_1099_12533# result[6] 6.17e-19
C10863 net40 a_9503_4399# 1.87e-19
C10864 net43 a_448_6549# 1.91e-19
C10865 clknet_2_3__leaf_clk a_12344_8041# 6.56e-19
C10866 a_2383_3689# a_2479_3689# 0.0138f
C10867 a_2601_3285# a_2645_3677# 3.69e-19
C10868 a_2033_3317# a_3057_3689# 2.36e-20
C10869 trim_mask\[4\] a_11045_3631# 1.57e-19
C10870 cal_count\[3\] a_10975_4105# 3.52e-20
C10871 a_7010_3311# a_7223_2465# 4.97e-21
C10872 trim_val\[3\] a_9805_1473# 1.39e-20
C10873 _108_ a_14000_4719# 1.18e-19
C10874 a_395_6031# VPWR 0.483f
C10875 net28 _045_ 1.65e-19
C10876 cal_itt\[1\] a_10903_7261# 1.28e-19
C10877 a_4131_8207# VPWR 0.197f
C10878 _108_ _033_ 6.2e-21
C10879 clknet_2_1__leaf_clk a_1835_12319# 2.14e-20
C10880 a_2953_9845# a_2961_9545# 1.21e-19
C10881 net45 _015_ 0.0237f
C10882 a_6793_8970# VPWR 0.261f
C10883 net14 a_911_6031# 0.00307f
C10884 _014_ a_1867_3317# 0.0202f
C10885 net49 _055_ 1.29e-20
C10886 a_12249_7663# cal_count\[2\] 1.81e-20
C10887 a_7201_9813# a_7079_10217# 3.16e-19
C10888 a_6983_10217# a_6888_10205# 0.0498f
C10889 _026_ _031_ 1.79e-20
C10890 _083_ a_7245_10205# 1.62e-20
C10891 _048_ clknet_2_2__leaf_clk 2.04e-20
C10892 _092_ _093_ 1.08e-19
C10893 net12 a_5340_6031# 2.05e-19
C10894 _104_ a_8491_2229# 3.03e-20
C10895 clknet_2_1__leaf_clk a_2450_9955# 0.00154f
C10896 net15 a_3411_7485# 0.00187f
C10897 cal_count\[0\] trimb[1] 4.96e-19
C10898 a_4959_9295# a_4871_8181# 1.58e-20
C10899 net31 _108_ 0.0162f
C10900 _074_ _009_ 0.0558f
C10901 net19 a_8105_10383# 0.0188f
C10902 net35 a_14981_4020# 6.06e-22
C10903 _058_ a_13519_4007# 0.00281f
C10904 net50 a_10838_2045# 1.41e-19
C10905 _092_ a_5166_5193# 0.00169f
C10906 _096_ a_3057_4719# 7.33e-19
C10907 a_7527_4631# a_7758_4759# 0.0049f
C10908 net14 _012_ 0.0159f
C10909 _033_ a_10655_2932# 0.109f
C10910 _078_ a_5997_10927# 7.17e-19
C10911 a_395_591# a_1276_565# 1.74e-20
C10912 net52 _077_ 5.79e-19
C10913 net18 _118_ 1.71e-19
C10914 clknet_0_clk net42 0.104f
C10915 _106_ _107_ 0.186f
C10916 trim_mask\[4\] a_9595_1679# 1.83e-22
C10917 a_5998_11471# VPWR 9e-19
C10918 a_395_7119# a_911_6031# 1.1e-20
C10919 _074_ cal 0.00431f
C10920 a_5515_6005# _075_ 0.0308f
C10921 a_14649_6031# _058_ 1.5e-19
C10922 _025_ a_10781_3311# 0.00186f
C10923 a_11059_7356# en_co_clk 2.76e-20
C10924 net54 a_6822_4399# 1.17e-20
C10925 _092_ a_2865_4460# 9.7e-21
C10926 _028_ a_7379_2197# 0.0336f
C10927 a_13459_3317# a_14335_2442# 6.92e-21
C10928 _101_ a_3053_8457# 0.0301f
C10929 net55 a_6737_4719# 2.28e-19
C10930 a_929_8757# a_1844_9129# 0.119f
C10931 state\[2\] a_6927_3311# 0.00858f
C10932 _090_ a_3123_3615# 9.09e-20
C10933 cal_itt\[2\] a_8485_4943# 3.12e-20
C10934 net19 a_9572_2601# 9.02e-20
C10935 a_8657_2229# a_9225_2197# 0.176f
C10936 clknet_0_clk a_4091_5309# 0.013f
C10937 a_2368_9955# a_2450_9955# 0.00477f
C10938 a_448_11445# result[7] 0.00234f
C10939 a_6633_9845# a_7548_10217# 0.119f
C10940 trim_val\[0\] a_15054_5193# 7.82e-19
C10941 net28 _023_ 2.04e-20
C10942 _001_ a_10903_7261# 0.323f
C10943 net15 a_3411_9839# 1.36e-20
C10944 net22 a_1476_4777# 8.95e-21
C10945 net55 a_5547_5603# 1.27e-19
C10946 a_763_8757# a_1497_8725# 0.0701f
C10947 _006_ a_929_8757# 0.252f
C10948 _074_ a_448_10357# 1.55e-19
C10949 net53 a_7939_10383# 0.00178f
C10950 _058_ a_14604_3017# 1.31e-19
C10951 _123_ a_10877_7983# 0.0096f
C10952 net44 a_8673_10625# 0.00124f
C10953 _049_ _106_ 2e-20
C10954 _034_ _092_ 0.00377f
C10955 a_8022_7119# a_8298_5487# 0.00246f
C10956 state\[2\] a_5363_4719# 1.72e-20
C10957 a_1476_7119# a_1638_7485# 0.00645f
C10958 _078_ a_1651_6005# 0.0109f
C10959 net40 _111_ 0.0034f
C10960 net2 a_12900_7663# 1.06e-19
C10961 a_8583_3317# a_9195_3689# 3.82e-19
C10962 _033_ a_9004_3677# 0.158f
C10963 _063_ _064_ 0.219f
C10964 net5 a_15023_5487# 0.00159f
C10965 a_10975_6031# net46 0.296f
C10966 _038_ a_11709_6273# 0.00104f
C10967 _050_ a_7571_4943# 3.15e-19
C10968 net29 _078_ 0.109f
C10969 a_3339_2767# clk 0.00263f
C10970 net55 a_5536_4399# 0.0508f
C10971 net34 _131_ 0.0115f
C10972 a_995_3530# clk 5.57e-20
C10973 _024_ a_9503_4399# 2.56e-20
C10974 clk rstn 0.0354f
C10975 _108_ _054_ 1.4e-20
C10976 a_2815_9447# a_2689_8751# 5.11e-20
C10977 _107_ _033_ 0.00183f
C10978 net21 _045_ 0.00973f
C10979 _088_ a_7010_3311# 2.44e-19
C10980 a_4165_10901# a_4674_10927# 2.6e-19
C10981 a_5363_7369# a_4259_6031# 4.58e-20
C10982 a_4995_7119# a_4425_6031# 4.94e-20
C10983 a_3597_10933# a_5997_10927# 6.47e-20
C10984 a_8912_2589# clk 7.28e-19
C10985 net30 VPWR 4.34f
C10986 net16 a_14379_6397# 0.0078f
C10987 net44 a_7164_11293# 0.00198f
C10988 _078_ _040_ 0.00186f
C10989 state\[2\] a_4959_1679# 7.62e-19
C10990 a_3781_8207# a_4239_8573# 0.0276f
C10991 clknet_2_0__leaf_clk a_4393_8207# 1.55e-19
C10992 _104_ a_10195_1354# 3.86e-19
C10993 net12 a_6197_6281# 4.37e-19
C10994 _060_ _087_ 0.00815f
C10995 net8 trim[2] 2.25e-19
C10996 a_5221_9295# VPWR 2.57e-19
C10997 a_6885_8372# a_6523_7119# 1.06e-19
C10998 a_7939_3855# a_7891_3617# 0.00107f
C10999 net50 trim_mask\[4\] 0.0786f
C11000 _122_ _053_ 0.203f
C11001 a_3388_4631# a_3667_3829# 5.85e-19
C11002 _072_ a_6173_7119# 3.02e-19
C11003 state\[0\] a_4959_1679# 4.69e-20
C11004 _094_ a_3891_4943# 5.63e-20
C11005 _098_ a_7571_4943# 0.191f
C11006 a_3116_12533# _085_ 0.0257f
C11007 _110_ a_8491_2229# 0.00698f
C11008 a_3431_12021# _078_ 0.00921f
C11009 a_1129_9813# net25 0.00128f
C11010 a_911_10217# a_1476_10217# 7.99e-20
C11011 clknet_0_clk a_8491_2229# 5.66e-19
C11012 trim_mask\[2\] _056_ 6.23e-19
C11013 _007_ a_911_10217# 5.1e-19
C11014 _060_ _099_ 0.00621f
C11015 _074_ a_561_4405# 0.0166f
C11016 _063_ _053_ 0.696f
C11017 a_7019_4407# a_6822_4399# 2.88e-19
C11018 net14 a_1129_9813# 0.0115f
C11019 net27 a_5998_11471# 0.00142f
C11020 mask\[3\] a_2961_9545# 0.0583f
C11021 _062_ a_7190_3855# 6.81e-21
C11022 a_6210_4989# calibrate 9.72e-20
C11023 clknet_2_0__leaf_clk a_2283_4020# 0.00103f
C11024 _041_ net45 1.44e-20
C11025 net22 _120_ 0.00171f
C11026 _081_ a_2689_8751# 0.0913f
C11027 net45 a_7184_2339# 0.0314f
C11028 net15 a_3933_2767# 1.04e-19
C11029 net43 a_1125_7663# 0.011f
C11030 _074_ mask\[6\] 0.491f
C11031 a_15083_4659# a_14715_3615# 9.15e-19
C11032 net32 a_13975_3689# 1.22e-19
C11033 net16 cal_count\[0\] 0.081f
C11034 a_1660_11305# mask\[3\] 1.09e-21
C11035 _104_ _032_ 3.44e-21
C11036 a_3868_7119# a_4995_7119# 7.24e-20
C11037 mask\[3\] mask\[0\] 1.07e-20
C11038 net12 a_6631_7485# 0.00178f
C11039 cal_itt\[1\] a_9889_6873# 0.0052f
C11040 clknet_2_1__leaf_clk a_4055_10927# 5.87e-19
C11041 net30 a_9478_4105# 1.45e-19
C11042 net55 a_8485_4943# 3.16e-19
C11043 cal_itt\[0\] a_9443_6059# 0.0479f
C11044 net44 net3 1.09e-20
C11045 net9 a_13512_4943# 7.31e-20
C11046 net4 _092_ 0.0098f
C11047 a_3781_8207# a_4167_6575# 5.64e-21
C11048 _053_ a_7104_3855# 1.26e-19
C11049 clknet_2_3__leaf_clk _133_ 0.00197f
C11050 _101_ a_4043_7093# 8.24e-20
C11051 a_15023_2223# VPWR 0.384f
C11052 _134_ VPWR 0.618f
C11053 _111_ _024_ 7.76e-21
C11054 _123_ a_12341_8751# 0.0146f
C11055 a_2857_5461# _015_ 3.35e-20
C11056 cal_count\[3\] a_10055_5487# 1.5e-19
C11057 _049_ a_4883_6397# 0.00244f
C11058 a_8298_2767# _116_ 3.83e-19
C11059 _105_ a_8745_4943# 0.00164f
C11060 a_11023_5108# _118_ 1.4e-20
C11061 a_13059_4631# trim_mask\[2\] 3.93e-21
C11062 a_6835_7669# a_7723_6807# 1.32e-21
C11063 a_3431_12021# a_3597_10933# 7.04e-19
C11064 net43 a_4871_8181# 3.85e-19
C11065 _050_ a_3557_5193# 3.07e-19
C11066 net23 a_2143_7663# 0.0304f
C11067 a_4687_12319# a_5496_12131# 7.54e-19
C11068 _107_ _054_ 0.00434f
C11069 a_15023_6031# a_15023_5487# 0.00787f
C11070 net43 _076_ 0.00837f
C11071 a_11297_7119# _136_ 1.62e-19
C11072 rstn ctln[0] 2.27e-19
C11073 _035_ _036_ 4.23e-21
C11074 _070_ a_8761_7983# 3.03e-20
C11075 net9 a_12546_9129# 2.06e-19
C11076 net18 a_10990_7485# 0.01f
C11077 a_10990_7485# a_10820_7485# 2.6e-19
C11078 a_10864_7387# a_11204_7485# 0.0346f
C11079 net12 a_5691_2741# 0.00737f
C11080 trim_mask\[0\] a_11691_4399# 2.51e-19
C11081 net3 clk 0.00563f
C11082 en_co_clk net3 0.0269f
C11083 a_11016_6691# en_co_clk 0.0135f
C11084 _060_ a_5537_4943# 8.38e-19
C11085 clknet_2_0__leaf_clk a_4680_6031# 0.00471f
C11086 a_10781_5487# _058_ 0.00122f
C11087 net28 _078_ 0.0029f
C11088 a_13975_3689# VPWR 0.216f
C11089 _110_ a_10195_1354# 0.0273f
C11090 _078_ a_5177_9537# 3.39e-21
C11091 a_4091_5309# net41 2.35e-21
C11092 net54 a_4617_4105# 4.43e-19
C11093 _049_ _054_ 0.243f
C11094 net4 cal_itt\[3\] 7.46e-21
C11095 _131_ a_15299_6575# 0.00106f
C11096 mask\[0\] a_1579_5807# 0.0106f
C11097 net12 a_5726_5807# 1.84e-20
C11098 clknet_2_2__leaf_clk _112_ 0.00632f
C11099 state\[2\] VPWR 1.13f
C11100 _062_ a_5625_4943# 0.00623f
C11101 a_4425_6031# a_4863_4917# 4.82e-19
C11102 a_561_4405# _093_ 1.05e-19
C11103 trim_mask\[0\] net49 5.76e-20
C11104 _123_ a_10864_7387# 0.00196f
C11105 net18 a_12502_4765# 5.71e-20
C11106 cal_itt\[2\] _105_ 9.08e-20
C11107 net43 a_579_10933# 0.307f
C11108 a_579_12021# a_1095_11305# 8.69e-21
C11109 net31 trimb[2] 3.03e-20
C11110 net47 a_13164_8029# 0.00232f
C11111 _013_ a_2033_3317# 0.223f
C11112 _099_ a_4498_4373# 0.0651f
C11113 state\[0\] VPWR 1.13f
C11114 trim_val\[2\] a_14172_1513# 0.00214f
C11115 _004_ a_1651_6005# 1.29e-20
C11116 net8 a_15023_1135# 0.00119f
C11117 a_10569_1109# a_11292_1251# 0.00128f
C11118 net9 a_10903_7261# 0.00441f
C11119 a_13915_4399# VPWR 0.292f
C11120 net9 a_11859_3689# 0.00272f
C11121 net19 a_9074_9955# 4.36e-19
C11122 cal_count\[3\] trim_val\[4\] 1.44e-20
C11123 a_2143_7663# a_2225_7663# 0.171f
C11124 a_11509_3317# a_11067_3017# 8.11e-20
C11125 net47 a_10864_9269# 0.174f
C11126 result[3] result[1] 0.00269f
C11127 net13 a_4680_6031# 0.00342f
C11128 trimb[4] comp 0.0482f
C11129 mask\[7\] a_448_11445# 1.11e-19
C11130 net45 _050_ 4.41e-19
C11131 net12 a_5997_10927# 0.00775f
C11132 net52 a_3852_11293# 1.96e-20
C11133 net4 a_9317_3285# 0.0085f
C11134 a_11233_4405# a_11583_4777# 0.23f
C11135 _106_ trim_mask\[4\] 1.48e-20
C11136 a_13519_4007# _113_ 0.11f
C11137 a_2143_7663# _016_ 0.11f
C11138 net18 net47 0.283f
C11139 clknet_2_1__leaf_clk mask\[4\] 0.0601f
C11140 _110_ _032_ 0.111f
C11141 net44 a_8083_8181# 0.00333f
C11142 net47 a_10820_7485# 4.46e-19
C11143 _065_ _077_ 0.173f
C11144 _092_ a_6763_5193# 0.0722f
C11145 a_4677_7882# _049_ 4.22e-19
C11146 a_395_4405# a_1585_4777# 2.56e-19
C11147 a_11023_5108# a_10137_4943# 2.1e-20
C11148 _108_ a_13715_5309# 0.00129f
C11149 net30 _104_ 0.677f
C11150 _078_ a_4167_11471# 0.0319f
C11151 clknet_2_0__leaf_clk a_911_4777# 0.00107f
C11152 a_4609_1679# ctln[7] 3.63e-20
C11153 net45 _052_ 1.21e-19
C11154 _042_ a_911_10217# 5.03e-21
C11155 _079_ a_1579_5807# 0.0016f
C11156 net45 a_5055_1679# 9.54e-19
C11157 _017_ clknet_2_0__leaf_clk 0.123f
C11158 a_10111_1679# a_10569_1109# 0.0059f
C11159 a_12436_9129# a_12546_9129# 0.00807f
C11160 _041_ a_3922_8867# 4.96e-19
C11161 a_12612_8725# a_12756_9117# 0.00196f
C11162 net12 _089_ 0.0146f
C11163 a_4131_8207# clknet_0_clk 0.00449f
C11164 net41 a_2479_3689# 0.0043f
C11165 net53 a_7710_9839# 4.26e-20
C11166 clknet_2_1__leaf_clk a_7447_8041# 1.98e-20
C11167 clknet_2_3__leaf_clk _129_ 3e-21
C11168 _111_ _029_ 0.00664f
C11169 _122_ a_13821_7119# 1.45e-19
C11170 net45 a_561_6031# 0.0264f
C11171 net52 a_3947_11305# 5.95e-20
C11172 _074_ result[0] 0.0228f
C11173 net16 a_13919_8751# 0.118f
C11174 _042_ a_9182_10749# 3.5e-19
C11175 a_8083_8181# clk 1.37e-19
C11176 a_10752_12533# net17 1.18e-20
C11177 _064_ a_9761_1679# 5e-19
C11178 net20 clknet_2_1__leaf_clk 0.0971f
C11179 net12 a_4609_1679# 8.6e-19
C11180 a_15023_10927# _126_ 2.66e-19
C11181 a_12344_8041# a_12664_8029# 0.00184f
C11182 a_3615_8207# net45 1.04e-20
C11183 a_12520_7637# a_12924_8029# 3.94e-19
C11184 _065_ a_10975_6031# 0.0135f
C11185 net44 mask\[0\] 2.97e-19
C11186 net47 a_9129_10383# 6.03e-19
C11187 _049_ a_5731_4943# 1.13e-19
C11188 a_1585_6031# VPWR 5.67e-20
C11189 clknet_2_0__leaf_clk net7 2.04e-20
C11190 net23 a_1019_7485# 9.76e-19
C11191 net21 _078_ 0.427f
C11192 trim_mask\[4\] _033_ 0.0193f
C11193 a_8083_8181# a_8386_8457# 0.00145f
C11194 net43 a_395_9845# 0.311f
C11195 a_11030_1679# VPWR 7.25e-20
C11196 a_4471_4007# a_4617_4105# 0.171f
C11197 a_14379_6397# clkc 3.36e-19
C11198 net1 a_937_3855# 0.00521f
C11199 mask\[7\] a_3431_10933# 6.45e-19
C11200 _059_ net3 0.0264f
C11201 _096_ a_3891_4943# 3.38e-20
C11202 a_763_8757# a_1129_7361# 3.48e-21
C11203 _100_ VPWR 0.397f
C11204 _006_ a_561_7119# 4.59e-21
C11205 _049_ a_4993_6273# 0.00926f
C11206 net13 _017_ 9.55e-19
C11207 net12 _040_ 1.15e-20
C11208 _047_ a_15083_4659# 0.0241f
C11209 _041_ _069_ 1.36e-19
C11210 a_9761_1679# a_10851_1653# 0.0424f
C11211 a_4259_6031# a_4498_4373# 5.83e-20
C11212 a_10329_1921# a_10111_1679# 0.21f
C11213 net32 trim_val\[1\] 0.00288f
C11214 net39 net38 0.067f
C11215 trim_mask\[1\] a_12077_3285# 0.0188f
C11216 a_2601_3285# a_2564_2589# 1.99e-20
C11217 a_11292_1251# a_11374_1251# 0.00477f
C11218 a_13257_1141# a_13703_1513# 2.28e-19
C11219 a_13183_3311# _030_ 0.109f
C11220 _041_ a_8022_7119# 6.5e-21
C11221 trim_mask\[1\] a_14686_3017# 5.26e-20
C11222 a_9458_9661# VPWR 7.9e-19
C11223 _042_ mask\[2\] 0.0316f
C11224 net55 _105_ 0.112f
C11225 a_11987_8757# _036_ 0.145f
C11226 a_4167_11471# a_3597_10933# 2.65e-20
C11227 a_13091_1141# trim[3] 4.94e-20
C11228 net19 net42 5.45e-21
C11229 a_13825_5185# trim[4] 1.68e-19
C11230 a_2143_2229# a_2877_2197# 0.0701f
C11231 clknet_2_1__leaf_clk a_2815_9447# 0.0724f
C11232 a_2787_9845# _018_ 0.285f
C11233 mask\[4\] a_7245_10205# 0.00207f
C11234 _108_ a_12599_3615# 5.16e-21
C11235 cal_itt\[0\] a_11396_6031# 7.48e-21
C11236 _064_ a_10787_1135# 1.87e-19
C11237 _067_ a_8025_8041# 2.25e-21
C11238 net4 a_9003_3829# 0.0117f
C11239 clk valid 5.35e-20
C11240 clknet_2_2__leaf_clk a_12121_3677# 2.34e-19
C11241 clknet_2_0__leaf_clk a_4425_6031# 0.11f
C11242 _001_ a_11141_6031# 2.94e-19
C11243 a_2953_7119# _050_ 5.42e-21
C11244 a_911_6031# VPWR 0.207f
C11245 net55 a_7010_3311# 3.94e-21
C11246 a_4043_10143# a_3781_8207# 1.97e-19
C11247 _126_ a_14377_9545# 0.00108f
C11248 a_3868_10217# a_3615_8207# 3.64e-21
C11249 a_6541_12021# a_7565_12393# 2.36e-20
C11250 clknet_2_1__leaf_clk a_1313_10901# 4.07e-20
C11251 a_7109_11989# a_7153_12381# 3.69e-19
C11252 _101_ a_5997_11247# 0.00328f
C11253 net29 a_3852_12381# 1.76e-20
C11254 _109_ a_13459_3317# 1.75e-20
C11255 _044_ a_8154_11721# 4.96e-19
C11256 _062_ _103_ 2.33e-19
C11257 clknet_2_2__leaf_clk a_11583_4777# 0.00175f
C11258 a_4696_8207# _077_ 2.9e-19
C11259 _078_ a_1549_6794# 0.0117f
C11260 net29 a_1651_10143# 1.08e-21
C11261 a_13307_1707# a_13512_1501# 2.34e-19
C11262 a_10851_1653# a_10787_1135# 7.21e-20
C11263 _108_ a_12257_4777# 3.22e-20
C11264 _078_ _020_ 3.53e-21
C11265 mask\[6\] _083_ 6.36e-20
C11266 trim_mask\[3\] a_11149_2767# 0.00216f
C11267 a_3339_2767# a_3399_2527# 0.00344f
C11268 mask\[3\] a_5423_9011# 5.26e-20
C11269 net30 _110_ 0.214f
C11270 en_co_clk a_5537_4105# 9.86e-20
C11271 net12 _048_ 0.489f
C11272 _012_ VPWR 0.981f
C11273 net4 a_9602_6941# 7.62e-19
C11274 a_10005_6031# _066_ 0.00683f
C11275 _128_ net2 0.0683f
C11276 a_8083_8181# a_8091_7967# 0.0114f
C11277 _065_ a_6173_7119# 1.17e-20
C11278 a_1313_11989# _078_ 0.00156f
C11279 net49 _030_ 4.69e-20
C11280 _072_ a_7351_8041# 0.00622f
C11281 a_1099_12533# a_1644_12533# 0.00355f
C11282 _005_ a_816_7119# 0.168f
C11283 _011_ result[5] 5.91e-19
C11284 net15 a_4443_9295# 6.81e-20
C11285 clknet_0_clk net30 0.237f
C11286 net14 a_1651_4703# 1.52e-19
C11287 a_15054_5193# VPWR 0.00225f
C11288 net16 en_co_clk 0.045f
C11289 _130_ comp 9.2e-19
C11290 state\[0\] a_2383_3689# 1.56e-19
C11291 net40 a_14282_7119# 2.78e-19
C11292 net36 net31 0.152f
C11293 _092_ a_3057_4719# 0.0603f
C11294 a_5691_7637# VPWR 0.595f
C11295 a_2787_9845# mask\[1\] 3.14e-21
C11296 net13 a_4425_6031# 0.0177f
C11297 trim_val\[1\] VPWR 0.815f
C11298 net47 a_12153_8757# 0.207f
C11299 clknet_2_1__leaf_clk _081_ 1e-19
C11300 net22 _014_ 5.06e-20
C11301 _108_ a_11057_3855# 1.46e-20
C11302 state\[2\] _104_ 0.0326f
C11303 a_9503_4399# a_8749_3317# 1.49e-21
C11304 a_7010_3311# a_7715_3285# 0.016f
C11305 net15 net52 0.228f
C11306 _014_ a_2921_2589# 3.81e-19
C11307 a_3431_12021# a_3852_12381# 0.0867f
C11308 net44 net54 1.35e-20
C11309 trim_val\[4\] _119_ 5.48e-20
C11310 net33 a_14172_4943# 1.36e-19
C11311 clknet_2_0__leaf_clk a_3868_7119# 0.061f
C11312 _054_ trim_mask\[4\] 1.48e-20
C11313 a_13783_6183# _135_ 0.398f
C11314 a_5340_6031# _048_ 2.81e-21
C11315 a_5699_9269# a_5691_7637# 1.06e-20
C11316 _084_ a_6891_12393# 1.05e-19
C11317 a_5089_10159# VPWR 4.34e-19
C11318 state\[1\] a_3333_2601# 1.2e-19
C11319 a_1497_8725# a_1279_9129# 0.21f
C11320 net51 a_7256_8029# 0.00158f
C11321 a_12424_3689# a_12691_2527# 5.34e-20
C11322 a_12599_3615# a_12516_2601# 1.18e-19
C11323 _067_ a_10975_6031# 1.77e-19
C11324 a_2857_5461# _050_ 0.0678f
C11325 a_12454_8041# VPWR 2.04e-19
C11326 _118_ VPWR 0.292f
C11327 net19 a_8491_2229# 0.0187f
C11328 cal_itt\[2\] a_8078_7663# 9.87e-20
C11329 _037_ a_13356_7369# 0.00106f
C11330 a_7184_2339# a_8657_2229# 0.00469f
C11331 a_6467_9845# a_6633_9845# 0.855f
C11332 a_2368_9955# _081_ 1.07e-20
C11333 net9 a_13825_1109# 3.21e-19
C11334 _002_ a_8022_7119# 0.00165f
C11335 a_14604_2339# _056_ 0.105f
C11336 a_2092_8457# mask\[1\] 0.132f
C11337 net44 a_6099_10633# 2.04e-19
C11338 a_4775_6031# VPWR 0.211f
C11339 en_co_clk net54 0.012f
C11340 net13 a_3868_7119# 3.56e-36
C11341 a_7548_10217# _072_ 2.67e-20
C11342 a_2476_6281# net30 1.66e-19
C11343 a_6316_5193# _052_ 1.88e-19
C11344 _064_ a_11067_3017# 0.0867f
C11345 a_6633_9845# VPWR 0.287f
C11346 _074_ ctlp[7] 0.0518f
C11347 net47 a_11268_9295# 0.00264f
C11348 _035_ net4 3.57e-20
C11349 a_8583_3317# _028_ 1.05e-19
C11350 net2 a_11895_7669# 1.21e-19
C11351 _096_ a_3530_4438# 0.00688f
C11352 mask\[3\] a_2489_7983# 7.06e-20
C11353 _098_ a_6316_5193# 0.126f
C11354 trim_mask\[3\] a_9572_2601# 0.00165f
C11355 a_10655_2932# a_10543_2455# 6.15e-20
C11356 a_10975_6031# clknet_2_2__leaf_clk 1.33e-19
C11357 calibrate a_7223_2465# 6.64e-20
C11358 a_448_7637# result[0] 1.11e-20
C11359 a_8657_2229# a_9734_2223# 1.46e-19
C11360 a_395_9845# a_2953_9845# 1.77e-21
C11361 _078_ a_2143_7663# 6.43e-20
C11362 _074_ a_1019_4399# 0.00346f
C11363 _125_ a_13256_9117# 7.89e-21
C11364 mask\[1\] net51 5.71e-20
C11365 mask\[5\] a_6090_10159# 1.96e-20
C11366 a_1129_9813# VPWR 0.22f
C11367 net17 _042_ 0.029f
C11368 cal_count\[3\] net55 6.92e-20
C11369 mask\[3\] a_4871_8181# 4.04e-19
C11370 _092_ _064_ 0.00523f
C11371 _059_ a_5537_4105# 3.87e-19
C11372 net4 _136_ 3e-20
C11373 mask\[3\] _076_ 7.04e-19
C11374 _118_ a_9478_4105# 0.0147f
C11375 net18 net46 0.0539f
C11376 net28 a_3852_12381# 0.0249f
C11377 mask\[5\] a_5915_11721# 0.0821f
C11378 _135_ a_14181_6031# 0.00236f
C11379 a_14983_9269# a_15159_9269# 0.185f
C11380 calibrate a_855_4105# 0.129f
C11381 a_6793_8970# a_6523_7119# 4.26e-21
C11382 _076_ a_6741_7361# 3.26e-20
C11383 net3 a_3399_2527# 4.42e-20
C11384 a_3411_7485# VPWR 0.143f
C11385 clknet_2_3__leaf_clk a_14379_6397# 0.2f
C11386 a_6445_10383# VPWR 3.07e-19
C11387 a_11016_6691# _108_ 1.4e-20
C11388 _099_ a_4576_3427# 7.19e-21
C11389 clknet_0_clk state\[2\] 5.82e-21
C11390 net16 cal_count\[2\] 0.0127f
C11391 a_13625_3317# a_13880_3677# 0.0642f
C11392 a_3388_4631# a_3339_2767# 2.12e-21
C11393 a_4815_3031# a_5177_1921# 0.00109f
C11394 a_14347_9480# _127_ 0.37f
C11395 a_455_12533# a_1099_12533# 0.00151f
C11396 net2 a_6419_8207# 0.00537f
C11397 net2 net35 1.98e-20
C11398 trim_mask\[1\] a_13257_1141# 1.13e-20
C11399 clknet_2_1__leaf_clk result[5] 0.0773f
C11400 _027_ clk 0.00154f
C11401 _101_ a_6056_8359# 0.00106f
C11402 _035_ a_11479_9117# 3.12e-20
C11403 a_10137_4943# VPWR 0.00812f
C11404 a_11435_2229# a_12691_2527# 0.0423f
C11405 net22 a_1638_6397# 2.15e-19
C11406 net52 net25 3.65e-19
C11407 a_11601_2229# a_11951_2601# 0.23f
C11408 net9 a_13715_1135# 4.52e-19
C11409 net46 a_12165_6031# 4.13e-19
C11410 _110_ a_13915_4399# 0.00182f
C11411 net43 result[6] 7.22e-20
C11412 net44 a_5423_9011# 0.00463f
C11413 net19 a_10195_1354# 2.95e-21
C11414 net31 _056_ 9.97e-20
C11415 net47 a_13050_7637# 0.119f
C11416 _085_ a_3597_12021# 0.0013f
C11417 a_13697_4373# a_13625_3317# 2.14e-21
C11418 clknet_2_3__leaf_clk _038_ 0.0816f
C11419 a_15023_6031# trim_val\[0\] 1.76e-19
C11420 a_12992_8751# trimb[4] 2.64e-22
C11421 net21 net12 2.37e-20
C11422 a_1660_12393# _046_ 3.69e-20
C11423 net14 net52 2.19e-20
C11424 a_12430_7663# VPWR 0.00334f
C11425 net52 a_3399_7119# 6.3e-20
C11426 a_7824_11305# a_7939_10383# 2.06e-19
C11427 a_7999_11231# a_8105_10383# 0.00889f
C11428 net9 a_11141_6031# 0.00198f
C11429 mask\[0\] a_3565_7119# 0.00218f
C11430 a_13016_9117# VPWR 1.63e-19
C11431 _053_ _092_ 0.0183f
C11432 a_3411_9839# VPWR 0.143f
C11433 en_co_clk a_4471_4007# 0.00177f
C11434 a_7527_4631# a_7800_4631# 0.168f
C11435 _062_ a_9889_6873# 0.0383f
C11436 net26 a_8215_9295# 6.75e-20
C11437 clknet_2_0__leaf_clk _121_ 0.0275f
C11438 trim_mask\[0\] _025_ 0.00129f
C11439 net46 trim_val\[0\] 0.00414f
C11440 clknet_2_3__leaf_clk cal_count\[0\] 0.36f
C11441 _059_ net54 0.318f
C11442 a_12148_4777# a_13915_4399# 1.68e-20
C11443 a_14655_4399# _109_ 1.08e-19
C11444 _058_ a_13233_4737# 2.95e-19
C11445 trim_mask\[0\] _026_ 1.75e-20
C11446 net3 en 0.0045f
C11447 trim_mask\[1\] a_10676_1679# 3.39e-21
C11448 mask\[2\] a_4959_9295# 7.1e-19
C11449 a_2019_9055# net45 1.36e-20
C11450 _024_ trim_mask\[2\] 3e-21
C11451 _035_ a_10586_7371# 3.54e-20
C11452 _134_ a_14564_6397# 6.6e-19
C11453 trim_val\[2\] _031_ 1.29e-19
C11454 net19 _032_ 1.11e-19
C11455 _078_ _077_ 0.015f
C11456 a_395_7119# a_816_7119# 0.0894f
C11457 net20 a_6927_12559# 0.238f
C11458 a_7259_11305# a_7164_11293# 0.0498f
C11459 a_7477_10901# a_7355_11305# 3.16e-19
C11460 a_395_9845# a_1585_10217# 2.56e-19
C11461 a_8381_9295# a_9458_9661# 1.46e-19
C11462 calibrate _088_ 0.218f
C11463 net18 a_11343_3317# 2.45e-21
C11464 a_15023_1135# trim[2] 0.00212f
C11465 net43 a_6835_7669# 0.921f
C11466 a_4498_4373# _097_ 3.18e-20
C11467 a_1019_4399# _093_ 8.82e-19
C11468 net18 a_11149_3017# 0.00283f
C11469 net31 net35 1.68e-19
C11470 _074_ a_4655_10071# 0.00126f
C11471 en_co_clk a_4970_4399# 2.85e-19
C11472 a_448_9269# result[3] 0.159f
C11473 a_10990_7485# VPWR 0.207f
C11474 net13 _121_ 3.21e-20
C11475 _048_ a_5691_2741# 7.08e-20
C11476 net21 a_3852_12381# 5.49e-20
C11477 a_12424_3689# VPWR 0.294f
C11478 net2 _061_ 1.78e-19
C11479 a_1129_4373# a_1638_4399# 2.6e-19
C11480 a_14184_2767# VPWR 1.86e-19
C11481 a_15023_10927# VPWR 0.497f
C11482 a_9664_3689# a_9761_1679# 3.03e-19
C11483 net12 _020_ 5.58e-20
C11484 a_8298_5487# a_10055_5487# 5.57e-19
C11485 _124_ _122_ 0.00765f
C11486 a_12061_7669# a_12344_8041# 0.215f
C11487 a_10586_7371# _136_ 5.64e-19
C11488 _134_ a_13091_4943# 2.04e-20
C11489 _078_ a_1019_7485# 8.7e-19
C11490 comp trim[4] 6.05e-20
C11491 _118_ _104_ 0.00748f
C11492 en_co_clk clkc 0.00312f
C11493 net15 state\[1\] 1.16e-19
C11494 calibrate a_6519_4631# 0.00314f
C11495 trim_mask\[0\] a_7677_4759# 0.00514f
C11496 net4 _105_ 0.00345f
C11497 _086_ a_1095_11305# 0.00197f
C11498 a_1830_4765# _099_ 5.67e-20
C11499 net28 a_1191_11305# 1.7e-19
C11500 _115_ a_13257_1141# 0.00186f
C11501 a_10689_2223# a_9761_1679# 4.56e-19
C11502 a_4443_1679# a_5177_1921# 0.0701f
C11503 net20 _009_ 0.0217f
C11504 _045_ a_7109_11989# 6.66e-20
C11505 net33 net48 1.38e-20
C11506 net26 a_1461_10357# 0.0495f
C11507 a_6210_4989# _098_ 0.127f
C11508 _070_ _071_ 1.97e-19
C11509 net23 _005_ 0.0439f
C11510 a_12502_4765# VPWR 2.34e-19
C11511 net16 cal_count\[1\] 0.0384f
C11512 net2 a_13257_4943# 2.47e-19
C11513 net15 _065_ 0.00704f
C11514 a_10864_9269# a_10774_9661# 9.35e-20
C11515 a_10688_9295# a_10593_9295# 0.0356f
C11516 _049_ net3 0.0661f
C11517 a_3933_2767# VPWR 0.611f
C11518 a_13142_7271# a_13279_7119# 0.0907f
C11519 a_1095_11305# _102_ 1.05e-19
C11520 net4 a_7010_3311# 7.28e-20
C11521 _130_ a_14199_7369# 0.0553f
C11522 a_13881_2741# a_14604_3017# 0.00128f
C11523 net3 a_3388_4631# 9.98e-19
C11524 net18 a_10774_9661# 5.82e-19
C11525 net44 a_4871_8181# 0.345f
C11526 _072_ a_8307_6575# 3.88e-19
C11527 net44 _076_ 0.148f
C11528 net40 net50 0.0315f
C11529 net15 net23 0.00814f
C11530 net46 a_11023_5108# 8.12e-20
C11531 net39 a_15023_12559# 0.203f
C11532 a_11321_3855# VPWR 1.35e-19
C11533 a_9103_2601# VPWR 4.33e-19
C11534 net38 net31 2.61e-20
C11535 _051_ trim_mask\[0\] 0.0111f
C11536 _074_ a_1129_7361# 0.00835f
C11537 a_7262_5461# a_8298_5487# 0.01f
C11538 net30 a_1137_5487# 5.38e-19
C11539 _065_ a_7351_8041# 3.64e-20
C11540 net47 VPWR 2.15f
C11541 _068_ a_8307_6575# 0.00106f
C11542 a_14377_9545# VPWR 0.26f
C11543 _053_ a_11045_5807# 0.00193f
C11544 net31 _061_ 1.31e-19
C11545 _094_ a_4680_6031# 0.025f
C11546 net45 _099_ 0.0026f
C11547 a_13415_2442# a_13307_1707# 0.00216f
C11548 clknet_2_0__leaf_clk a_3273_4943# 1.79e-19
C11549 trim_mask\[4\] a_11413_2767# 1.19e-19
C11550 _074_ a_1095_12393# 0.00163f
C11551 net29 a_3431_12021# 0.00312f
C11552 _075_ _051_ 0.15f
C11553 a_15023_1679# _114_ 1.25e-20
C11554 _042_ a_4609_9295# 7.52e-20
C11555 a_1677_9545# a_929_8757# 4.52e-20
C11556 net34 a_14172_4943# 4.6e-20
C11557 a_1679_10633# net25 5.91e-19
C11558 net46 a_10055_2767# 0.347f
C11559 _041_ net51 4.43e-20
C11560 _122_ a_13356_7369# 4.73e-19
C11561 net24 a_455_8181# 0.221f
C11562 state\[2\] net41 2.15e-19
C11563 net45 a_6927_591# 5.09e-20
C11564 _110_ trim_val\[1\] 8.48e-19
C11565 net45 a_1129_4373# 0.166f
C11566 a_1660_11305# a_2787_10927# 2.95e-19
C11567 _109_ trim[1] 6.11e-20
C11568 net43 a_911_10217# 0.156f
C11569 a_10586_7371# a_10861_7119# 0.00742f
C11570 a_3868_7119# a_4167_6575# 0.00442f
C11571 net33 trimb[4] 3.24e-19
C11572 a_763_8757# mask\[1\] 5.17e-20
C11573 _048_ _089_ 0.164f
C11574 net46 a_9926_2589# 0.00331f
C11575 a_929_8757# a_1651_7093# 5.28e-20
C11576 a_11895_7669# a_12249_7663# 0.069f
C11577 _076_ en_co_clk 0.129f
C11578 _005_ a_2225_7663# 5e-20
C11579 a_8820_6005# VPWR 0.17f
C11580 _092_ a_3891_4943# 5.22e-19
C11581 _095_ net55 0.0478f
C11582 net16 _108_ 0.253f
C11583 a_7355_11305# VPWR 8.07e-19
C11584 a_11435_2229# VPWR 0.518f
C11585 a_1099_12533# a_745_12021# 0.00632f
C11586 state\[0\] net41 0.272f
C11587 net43 a_1585_7119# 0.00157f
C11588 a_6056_8359# a_6515_8534# 6.64e-19
C11589 net19 net30 0.00891f
C11590 a_9443_6059# a_9529_6059# 0.00658f
C11591 clknet_2_1__leaf_clk a_3781_8207# 1.11e-20
C11592 a_2828_12131# a_3597_12021# 2.04e-19
C11593 _063_ a_8473_5193# 0.0324f
C11594 a_7571_4943# a_7393_5193# 6.01e-20
C11595 net15 a_2225_7663# 4.09e-19
C11596 valid en 0.00147f
C11597 trim[1] trim[2] 3.16e-20
C11598 a_4443_1679# a_5633_1679# 2.56e-19
C11599 net24 a_2006_8751# 4.39e-19
C11600 a_1844_9129# a_2689_8751# 6.28e-19
C11601 mask\[6\] mask\[4\] 5.62e-20
C11602 trim_mask\[4\] a_11057_3855# 2.05e-19
C11603 _058_ a_14649_3689# 1.11e-19
C11604 a_10864_9269# _065_ 7.36e-20
C11605 net15 _016_ 0.0382f
C11606 a_10569_1109# a_10872_1455# 0.00138f
C11607 _118_ _110_ 0.0398f
C11608 cal_count\[3\] a_9595_5193# 0.0689f
C11609 net18 _065_ 0.661f
C11610 clknet_0_clk _118_ 2.72e-21
C11611 _004_ a_1007_6031# 2.31e-19
C11612 a_9296_9295# net4 1.61e-19
C11613 _053_ a_9003_3829# 0.00233f
C11614 a_745_10933# net26 1.15e-20
C11615 net44 ctlp[6] 2.53e-19
C11616 _108_ a_10699_3311# 1.61e-21
C11617 a_763_8757# a_1387_8751# 9.73e-19
C11618 net46 a_12691_2527# 0.35f
C11619 a_7569_7637# a_7613_8029# 3.69e-19
C11620 a_7001_7669# a_8025_8041# 2.36e-20
C11621 net46 _114_ 0.0171f
C11622 cal_itt\[1\] net30 0.00168f
C11623 net43 mask\[2\] 0.00361f
C11624 clknet_0_clk a_4775_6031# 1.84e-19
C11625 a_14686_2339# VPWR 0.00208f
C11626 clknet_2_0__leaf_clk a_816_6031# 0.00107f
C11627 a_1651_4703# VPWR 0.404f
C11628 net50 _024_ 2.32e-20
C11629 _072_ a_7897_6913# 6.42e-19
C11630 trim_mask\[0\] a_11801_4373# 7.95e-19
C11631 net20 mask\[6\] 1.84e-19
C11632 net45 a_4259_6031# 2.29e-20
C11633 a_10699_3311# a_10655_2932# 1.85e-19
C11634 a_2601_3285# a_2143_2229# 0.00112f
C11635 a_2033_3317# a_2309_2229# 9.38e-21
C11636 trim_mask\[4\] a_10543_2455# 0.0667f
C11637 net44 clknet_2_3__leaf_clk 0.00416f
C11638 trim_val\[3\] a_13091_1141# 9.05e-23
C11639 net5 VPWR 0.48f
C11640 net28 net29 0.0207f
C11641 _060_ a_4709_2773# 0.00124f
C11642 _063_ a_8583_3317# 9.79e-21
C11643 net25 net23 2.15e-22
C11644 result[5] result[4] 0.049f
C11645 net4 cal_count\[3\] 0.0122f
C11646 _112_ a_13459_3317# 0.0184f
C11647 net9 a_12625_2601# 4.37e-19
C11648 mask\[0\] _049_ 0.0782f
C11649 _064_ trim_val\[3\] 4.87e-20
C11650 net16 a_12516_2601# 6.01e-21
C11651 _062_ net42 7.43e-19
C11652 a_4308_4917# _060_ 1.36e-20
C11653 net18 a_11233_4405# 0.00863f
C11654 net51 _002_ 0.0071f
C11655 _100_ net41 0.0383f
C11656 a_14063_7093# _131_ 0.0586f
C11657 net14 net23 0.00709f
C11658 _130_ a_14422_7093# 0.0431f
C11659 net33 trim[0] 0.00267f
C11660 net43 a_6428_7119# 5.43e-21
C11661 a_14347_1439# VPWR 0.379f
C11662 net51 _050_ 4.53e-21
C11663 a_4801_9839# a_4871_8181# 1.26e-21
C11664 a_3123_3615# a_3339_2767# 0.0122f
C11665 net43 a_1000_11293# 2.56e-19
C11666 clknet_0_clk a_3411_7485# 3.18e-19
C11667 net30 a_11067_4405# 9.27e-21
C11668 net12 _077_ 0.00266f
C11669 _109_ _112_ 0.00155f
C11670 net40 net2 0.0254f
C11671 net28 a_3431_12021# 0.209f
C11672 clknet_2_0__leaf_clk a_1651_7093# 1.65e-19
C11673 _085_ net43 0.00429f
C11674 clknet_2_3__leaf_clk en_co_clk 0.0129f
C11675 a_10851_1653# trim_val\[3\] 0.0618f
C11676 mask\[6\] a_2815_9447# 1.11e-20
C11677 cal_itt\[2\] a_8298_5487# 0.00843f
C11678 _094_ a_4425_6031# 0.0221f
C11679 _095_ _093_ 1.33e-19
C11680 _057_ a_10787_1135# 2.45e-19
C11681 _132_ _130_ 0.345f
C11682 net9 a_11764_3677# 5.07e-19
C11683 a_13562_8751# _041_ 0.0475f
C11684 _065_ a_5449_6031# 9.91e-20
C11685 a_2491_3311# a_2309_2229# 5.3e-20
C11686 net45 a_4043_7093# 6.73e-19
C11687 clknet_2_3__leaf_clk a_9084_4515# 3.57e-20
C11688 _053_ a_8485_4943# 1.72e-19
C11689 _136_ _064_ 2.37e-19
C11690 net16 a_12900_7663# 8.39e-19
C11691 _019_ a_4443_9295# 0.167f
C11692 _057_ trim[3] 3.31e-19
C11693 net23 a_395_7119# 2.87e-19
C11694 mask\[6\] a_1313_10901# 2.18e-21
C11695 a_6906_2355# a_7379_2197# 7.99e-20
C11696 _026_ a_11951_2601# 0.00195f
C11697 a_7223_2465# a_7184_2339# 0.725f
C11698 _095_ a_5166_5193# 1.16e-19
C11699 net33 _130_ 0.00557f
C11700 clknet_2_1__leaf_clk a_561_9845# 0.596f
C11701 _108_ _027_ 8.23e-22
C11702 _104_ a_11321_3855# 0.00411f
C11703 net33 a_14335_4020# 1.19e-19
C11704 _121_ a_4167_6575# 0.189f
C11705 a_15023_1679# VPWR 0.28f
C11706 _014_ a_2877_2197# 6.4e-19
C11707 _003_ _050_ 3.51e-20
C11708 a_8105_10383# a_9020_10383# 0.119f
C11709 a_6181_10633# _042_ 0.0425f
C11710 net47 a_8455_10383# 0.153f
C11711 net52 _019_ 9.79e-21
C11712 a_7939_10383# _043_ 3.7e-19
C11713 net46 net32 2.32e-19
C11714 _092_ a_3530_4438# 5.89e-19
C11715 mask\[2\] a_2857_7637# 0.014f
C11716 _012_ net41 9.64e-19
C11717 _078_ a_3947_11305# 0.00122f
C11718 trim_mask\[1\] trim_mask\[2\] 0.0266f
C11719 _080_ a_561_7119# 6.57e-20
C11720 a_2857_5461# _099_ 0.00122f
C11721 _095_ a_2865_4460# 0.217f
C11722 net47 a_9650_9295# 0.00392f
C11723 a_2033_3317# a_3110_3311# 1.46e-19
C11724 state\[1\] a_2659_2601# 1.69e-19
C11725 net55 calibrate 0.404f
C11726 net54 _107_ 9.96e-19
C11727 a_14655_4399# trim[1] 0.00212f
C11728 net14 _016_ 1.04e-20
C11729 net18 _067_ 0.0225f
C11730 _037_ a_10903_7261# 0.00269f
C11731 _067_ a_10820_7485# 8.41e-20
C11732 trim_mask\[3\] a_8491_2229# 7.85e-20
C11733 _072_ VPWR 1.06f
C11734 _051_ a_8298_2767# 6.84e-19
C11735 _018_ a_2961_9295# 2.47e-19
C11736 net14 a_1019_6397# 9.07e-20
C11737 _065_ a_4222_7119# 1.27e-19
C11738 a_3431_12021# a_4167_11471# 3.54e-20
C11739 _030_ _031_ 2.09e-19
C11740 _034_ _095_ 4.95e-20
C11741 a_3597_10933# a_3852_11293# 0.0642f
C11742 a_561_9845# a_2368_9955# 2.8e-20
C11743 a_2564_2589# clk 0.00205f
C11744 net31 net40 2.27e-19
C11745 a_4498_4373# a_4709_2773# 1.51e-20
C11746 a_15023_12015# VPWR 0.445f
C11747 _027_ a_9115_2223# 8.49e-19
C11748 _068_ VPWR 0.958f
C11749 _074_ calibrate 0.299f
C11750 _104_ a_11435_2229# 1.59e-19
C11751 a_7916_8041# net30 8.45e-20
C11752 _053_ _136_ 0.0545f
C11753 a_7723_6807# _051_ 7.77e-20
C11754 net33 a_15023_2767# 0.0052f
C11755 a_15023_6031# VPWR 0.259f
C11756 a_9463_8725# net4 0.229f
C11757 _065_ a_11023_5108# 9.5e-22
C11758 _049_ net54 0.392f
C11759 a_395_591# VPWR 0.275f
C11760 a_9317_3285# a_9664_3689# 0.0512f
C11761 a_8749_3317# trim_mask\[2\] 6.73e-20
C11762 a_4443_9295# VPWR 0.48f
C11763 _131_ a_13279_7119# 0.00144f
C11764 a_4512_12393# a_4674_12015# 0.00645f
C11765 a_4308_4917# a_4498_4373# 8.26e-19
C11766 _051_ a_7210_5807# 5.25e-20
C11767 net43 a_4674_10927# 2.88e-19
C11768 _110_ a_12424_3689# 3.3e-20
C11769 net28 a_1191_12393# 0.00177f
C11770 _110_ a_14184_2767# 1.12e-19
C11771 _016_ a_395_7119# 2.75e-21
C11772 a_448_10357# result[5] 0.00311f
C11773 net18 clknet_2_2__leaf_clk 0.123f
C11774 _106_ _024_ 7.33e-22
C11775 a_6835_7669# a_6741_7361# 1.38e-19
C11776 net52 VPWR 1.43f
C11777 a_7001_7669# a_6173_7119# 3.79e-20
C11778 trim_mask\[1\] a_11045_3631# 0.00366f
C11779 net46 VPWR 4.73f
C11780 a_4609_9295# a_4959_9295# 0.212f
C11781 a_4443_9295# a_5699_9269# 0.0436f
C11782 a_816_7119# VPWR 0.0854f
C11783 a_7190_3855# a_7104_3855# 0.00138f
C11784 _054_ a_6737_3855# 7.75e-20
C11785 a_11509_3317# a_12586_3311# 1.46e-19
C11786 net21 a_3431_12021# 7.59e-19
C11787 _007_ _082_ 0.113f
C11788 net47 a_8381_9295# 0.032f
C11789 a_8673_10625# a_8949_9537# 7e-20
C11790 a_8105_10383# a_8731_9295# 3.24e-19
C11791 clknet_2_0__leaf_clk a_4091_5309# 8.64e-21
C11792 _055_ trim_val\[2\] 5.25e-19
C11793 a_3597_10933# a_3947_11305# 0.23f
C11794 _011_ result[7] 0.00565f
C11795 net16 trimb[2] 3.94e-19
C11796 net26 _041_ 5.16e-20
C11797 _084_ net53 6.92e-21
C11798 a_2953_9845# mask\[2\] 0.00833f
C11799 a_3521_9813# a_3411_9839# 0.0977f
C11800 _023_ net25 1.3e-20
C11801 a_11709_6273# a_11587_6031# 3.16e-19
C11802 net46 a_12218_6397# 1.7e-19
C11803 a_1549_6794# a_1651_6005# 0.00116f
C11804 _090_ _060_ 0.00512f
C11805 _129_ a_12061_7669# 0.00163f
C11806 a_10990_7485# a_10699_5487# 4.37e-21
C11807 net55 a_8298_5487# 1.03e-19
C11808 a_13059_4631# a_12599_3615# 3.41e-19
C11809 net3 a_3123_3615# 0.00391f
C11810 _058_ a_12077_3285# 0.0021f
C11811 a_2787_7119# a_3868_7119# 0.102f
C11812 a_3521_7361# a_3303_7119# 0.21f
C11813 a_2953_7119# a_4043_7093# 0.0424f
C11814 _058_ a_14686_3017# 5.6e-20
C11815 net14 _023_ 0.0179f
C11816 net12 a_6173_7119# 0.0173f
C11817 clknet_2_3__leaf_clk cal_count\[2\] 3.1e-20
C11818 net15 a_2755_2601# 0.00103f
C11819 _074_ a_1461_10357# 0.206f
C11820 a_6743_10933# a_7939_10383# 8.63e-20
C11821 _078_ _005_ 2.11e-19
C11822 _050_ a_7223_2465# 7.37e-19
C11823 net13 a_4901_2773# 2.46e-19
C11824 net4 _119_ 0.648f
C11825 net1 clk 2.9e-20
C11826 net29 a_1313_11989# 0.00218f
C11827 a_1644_12533# net43 4.29e-20
C11828 a_7019_4407# _107_ 0.00977f
C11829 a_3057_4719# a_3148_4399# 0.0023f
C11830 a_5931_4105# VPWR 0.362f
C11831 a_9099_3689# a_9207_3311# 0.0572f
C11832 a_9839_3615# a_10018_3677# 0.0074f
C11833 a_9664_3689# a_9773_3689# 0.00742f
C11834 net34 a_13091_1141# 2.68e-20
C11835 net19 a_9458_9661# 9.48e-20
C11836 _064_ _105_ 3.99e-19
C11837 trim_mask\[2\] _115_ 0.0818f
C11838 net25 a_816_10205# 4.37e-20
C11839 net34 trimb[4] 0.0785f
C11840 clknet_2_3__leaf_clk a_10688_9295# 0.0467f
C11841 _058_ a_9503_4399# 0.0014f
C11842 net15 _078_ 0.00631f
C11843 _063_ a_9957_7663# 0.0474f
C11844 trim_mask\[3\] a_10195_1354# 3.63e-19
C11845 net47 clknet_0_clk 5.33e-19
C11846 a_8992_9955# clknet_2_3__leaf_clk 6.28e-21
C11847 a_561_7119# a_1651_7093# 0.0424f
C11848 a_1129_7361# a_911_7119# 0.21f
C11849 clknet_2_2__leaf_clk trim_val\[0\] 2.4e-19
C11850 a_13257_4943# a_13715_5309# 0.0276f
C11851 a_14347_4917# a_14172_4943# 0.234f
C11852 net28 a_4167_11471# 1.04e-20
C11853 a_11951_2601# _031_ 1.22e-19
C11854 net45 a_7942_2223# 2.56e-19
C11855 _051_ a_5177_1921# 4.03e-21
C11856 net14 _013_ 3.23e-20
C11857 _046_ a_4674_12015# 7.93e-21
C11858 a_5915_10927# a_6261_11247# 0.0134f
C11859 calibrate _093_ 1.41f
C11860 _049_ a_7019_4407# 0.0108f
C11861 a_8215_9295# a_8636_9295# 0.0902f
C11862 _000_ a_9296_9295# 5.47e-21
C11863 mask\[0\] sample 1.96e-19
C11864 clknet_2_1__leaf_clk a_1844_9129# 3.88e-21
C11865 sample valid 0.0379f
C11866 _074_ a_6191_12559# 2.4e-19
C11867 a_455_8181# result[1] 0.00235f
C11868 net43 a_2828_12131# 3.83e-20
C11869 _085_ a_2953_9845# 3.94e-21
C11870 clknet_2_1__leaf_clk a_5496_12131# 0.0393f
C11871 trim_val\[4\] a_9839_3615# 0.063f
C11872 clknet_2_1__leaf_clk _006_ 0.00374f
C11873 _049_ a_4471_4007# 6.11e-19
C11874 a_6210_4989# _087_ 0.0132f
C11875 net2 _071_ 1.4e-19
C11876 net47 a_10699_5487# 4.88e-20
C11877 _110_ a_11435_2229# 1.2e-19
C11878 _126_ a_14552_9071# 2.2e-20
C11879 a_11343_3317# VPWR 0.411f
C11880 clknet_0_clk a_8820_6005# 4.96e-19
C11881 clknet_2_3__leaf_clk a_12410_6031# 0.00219f
C11882 a_4995_7119# net30 1.5e-19
C11883 _052_ a_9099_3689# 1.55e-20
C11884 a_11149_3017# VPWR 0.191f
C11885 _044_ a_7939_10383# 4.75e-20
C11886 a_8072_11721# a_8105_10383# 1.58e-20
C11887 _128_ trimb[1] 1.84e-19
C11888 _118_ a_11057_4105# 5.6e-20
C11889 net27 net52 3.96e-19
C11890 _053_ _105_ 0.154f
C11891 a_4043_7093# a_2857_5461# 0.00124f
C11892 trim_mask\[3\] _032_ 0.00318f
C11893 net28 net21 0.0199f
C11894 a_6210_4989# _099_ 1.37e-20
C11895 calibrate a_2865_4460# 9.55e-20
C11896 _048_ a_7758_4759# 1.17e-19
C11897 mask\[1\] a_4858_8573# 4.37e-19
C11898 _056_ a_14931_591# 6.48e-19
C11899 a_3273_4943# a_3461_5193# 0.0101f
C11900 a_8491_2229# net11 1.44e-20
C11901 _121_ _094_ 0.0342f
C11902 a_4425_6031# _096_ 6.48e-19
C11903 net26 _002_ 4.53e-21
C11904 net23 a_2313_6183# 2.59e-19
C11905 net45 _097_ 0.235f
C11906 net37 a_15023_2223# 6.98e-21
C11907 _090_ a_4498_4373# 0.164f
C11908 _053_ a_7010_3311# 0.00615f
C11909 net37 _134_ 1.79e-20
C11910 _049_ a_4970_4399# 0.00703f
C11911 _074_ mask\[1\] 0.0263f
C11912 a_6099_10633# _008_ 1.5e-20
C11913 net43 _120_ 5.67e-20
C11914 net50 trim_mask\[1\] 0.191f
C11915 _079_ sample 0.00111f
C11916 trimb[3] trimb[2] 0.0408f
C11917 _074_ a_745_10933# 0.0206f
C11918 _050_ _088_ 0.121f
C11919 net19 _118_ 3.87e-20
C11920 a_455_5747# result[0] 0.00176f
C11921 _111_ _058_ 0.0177f
C11922 a_7262_5461# _050_ 0.216f
C11923 net33 trim[4] 3.24e-19
C11924 clknet_2_1__leaf_clk result[7] 0.00252f
C11925 a_11023_5108# clknet_2_2__leaf_clk 9.57e-19
C11926 net44 a_6835_7669# 0.0191f
C11927 a_8455_10383# _068_ 6.22e-19
C11928 a_2971_8457# clknet_2_0__leaf_clk 0.0312f
C11929 a_1679_10633# VPWR 0.286f
C11930 a_10774_9661# VPWR 0.00414f
C11931 mask\[3\] mask\[2\] 0.0187f
C11932 net34 trim[0] 0.105f
C11933 net55 _015_ 0.00176f
C11934 trim_mask\[4\] a_10699_3311# 0.0106f
C11935 _051_ a_5633_1679# 5.08e-20
C11936 _042_ _082_ 0.00156f
C11937 a_2019_9055# a_2092_8457# 0.00109f
C11938 _040_ a_2143_7663# 1.86e-19
C11939 net21 a_4167_11471# 0.111f
C11940 a_1313_11989# a_1191_12393# 3.16e-19
C11941 net43 a_1000_12381# 2.56e-19
C11942 net53 a_4801_10159# 0.00406f
C11943 a_6566_5193# a_6763_5193# 0.145f
C11944 _052_ _088_ 0.133f
C11945 a_395_4405# cal 0.00255f
C11946 net50 a_8749_3317# 1.03e-20
C11947 a_579_10933# a_2787_10927# 5.41e-21
C11948 _074_ a_1387_8751# 1.23e-20
C11949 net20 ctlp[7] 4.56e-19
C11950 net28 a_1313_11989# 0.00719f
C11951 net9 _134_ 8.17e-20
C11952 clknet_2_2__leaf_clk a_10055_2767# 0.105f
C11953 net16 net36 2.74e-19
C11954 _078_ net25 0.407f
C11955 net13 a_3840_8867# 9.7e-19
C11956 a_561_9845# result[4] 9.51e-19
C11957 a_395_9845# result[3] 0.00348f
C11958 _098_ _088_ 2.83e-19
C11959 a_3057_3689# VPWR 3.62e-20
C11960 net2 a_13349_6031# 0.0685f
C11961 a_5455_4943# a_5625_4943# 0.00167f
C11962 net46 _104_ 0.688f
C11963 _041_ cal_itt\[2\] 5.23e-20
C11964 _123_ net2 0.0507f
C11965 a_7262_5461# _098_ 1.09e-19
C11966 net47 a_14467_8751# 2.46e-20
C11967 a_3781_8207# a_4805_8207# 2.36e-20
C11968 net50 a_10977_2543# 9.28e-19
C11969 a_6835_7669# clk 0.00415f
C11970 clknet_2_2__leaf_clk a_9926_2589# 4.64e-19
C11971 a_6835_7669# en_co_clk 3.78e-21
C11972 net14 _078_ 0.304f
C11973 net4 a_9225_2197# 0.00111f
C11974 net13 a_2971_8457# 1.03e-19
C11975 net34 _130_ 0.0128f
C11976 _076_ _107_ 2.89e-19
C11977 _112_ trim[1] 4.99e-21
C11978 clknet_2_1__leaf_clk _017_ 6.06e-19
C11979 a_7527_4631# VPWR 0.2f
C11980 net13 a_4886_4399# 9e-19
C11981 _074_ a_6796_12381# 2.76e-20
C11982 a_1476_6031# a_1638_6397# 0.00645f
C11983 cal_count\[3\] _064_ 0.297f
C11984 _080_ a_1467_7923# 8.51e-19
C11985 a_6519_4631# _052_ 0.154f
C11986 _122_ a_10903_7261# 0.0101f
C11987 net41 a_3933_2767# 1.11e-19
C11988 _056_ a_13881_1653# 2.92e-20
C11989 a_10689_2223# trim_val\[3\] 1.23e-20
C11990 a_1279_9129# a_1387_8751# 0.0572f
C11991 a_1844_9129# a_1953_9129# 0.00742f
C11992 a_2019_9055# a_2198_9117# 0.0074f
C11993 a_1497_8725# _081_ 1.59e-19
C11994 net44 a_5515_6005# 0.289f
C11995 a_448_6549# sample 4.4e-21
C11996 _005_ _004_ 0.00243f
C11997 a_10383_7093# a_10586_7371# 0.234f
C11998 a_8022_7119# a_10864_7387# 1.02e-19
C11999 a_6173_7119# a_6631_7485# 0.0346f
C12000 a_10195_1354# net11 4.84e-20
C12001 a_3891_4943# a_4266_4943# 9.37e-20
C12002 a_4091_5309# a_4091_4943# 2.58e-19
C12003 state\[1\] VPWR 0.552f
C12004 net20 _021_ 1.25e-19
C12005 clknet_2_3__leaf_clk _108_ 1.78e-19
C12006 net44 a_7201_9813# 0.165f
C12007 _048_ a_6197_4399# 3.92e-19
C12008 _098_ a_6519_4631# 0.0614f
C12009 _011_ mask\[7\] 2.81e-19
C12010 a_8381_9295# _068_ 0.00885f
C12011 cal_count\[0\] a_14733_9545# 0.00146f
C12012 _000_ a_9463_8725# 1.13e-19
C12013 _091_ a_10975_6031# 0.00191f
C12014 _101_ net2 3.53e-21
C12015 _076_ _049_ 0.143f
C12016 a_13519_4007# a_13693_3883# 0.00658f
C12017 _125_ a_13557_8457# 2.04e-21
C12018 _078_ a_395_7119# 0.00772f
C12019 trim_val\[0\] a_14540_3689# 2.64e-21
C12020 clknet_2_2__leaf_clk a_6927_3311# 1.54e-21
C12021 net40 a_13715_5309# 6.24e-19
C12022 mask\[5\] a_6181_10633# 0.0146f
C12023 _092_ a_8473_5193# 9.77e-20
C12024 clknet_2_2__leaf_clk a_12691_2527# 0.0163f
C12025 a_12059_2223# VPWR 0.145f
C12026 a_2857_7637# _120_ 4.98e-20
C12027 net4 calibrate 2.6e-19
C12028 _065_ VPWR 3.3f
C12029 net16 _128_ 0.0758f
C12030 _062_ net30 0.148f
C12031 net45 a_845_7663# 5.77e-21
C12032 net34 a_15023_2767# 0.0251f
C12033 a_8360_10383# a_8215_9295# 1.6e-20
C12034 _118_ a_11067_4405# 1.7e-20
C12035 net40 a_14733_7983# 0.00189f
C12036 clknet_2_0__leaf_clk a_395_6031# 0.259f
C12037 net23 VPWR 0.72f
C12038 a_5515_6005# en_co_clk 0.125f
C12039 clknet_2_0__leaf_clk a_4131_8207# 0.0014f
C12040 _040_ _077_ 8.91e-20
C12041 a_4576_3427# a_4709_2773# 0.00167f
C12042 trim_mask\[4\] _027_ 3.06e-19
C12043 _032_ net11 1.11e-19
C12044 a_8298_5487# a_9595_5193# 0.00122f
C12045 a_5699_9269# _065_ 0.00339f
C12046 a_5524_9295# a_5423_9011# 0.00157f
C12047 a_5054_4399# VPWR 0.0058f
C12048 _072_ clknet_0_clk 0.00187f
C12049 _053_ cal_count\[3\] 0.0162f
C12050 net33 _057_ 4.43e-21
C12051 _136_ a_11425_5487# 4.88e-19
C12052 trim_mask\[1\] a_14604_2339# 1.33e-19
C12053 net17 cal_count\[0\] 9.79e-21
C12054 clknet_2_3__leaf_clk a_11436_9295# 1.82e-19
C12055 a_395_4405# a_561_4405# 0.888f
C12056 a_7019_4407# trim_mask\[4\] 9.23e-21
C12057 cal_itt\[0\] trim_mask\[0\] 7.46e-19
C12058 a_14471_12559# ctlp[2] 0.158f
C12059 net5 a_14564_6397# 6.96e-19
C12060 mask\[4\] a_4655_10071# 0.0892f
C12061 net54 a_3123_3615# 6.52e-20
C12062 _068_ clknet_0_clk 0.0251f
C12063 _104_ a_11343_3317# 0.0099f
C12064 a_2659_2601# a_2755_2601# 0.0138f
C12065 a_2309_2229# a_3333_2601# 2.36e-20
C12066 a_2877_2197# a_2921_2589# 3.69e-19
C12067 _104_ a_11149_3017# 0.0601f
C12068 net46 a_12678_2223# 3.67e-19
C12069 a_9826_3311# VPWR 0.00122f
C12070 _093_ _015_ 0.0433f
C12071 a_7001_7669# a_7351_8041# 0.219f
C12072 a_6835_7669# a_8091_7967# 0.0435f
C12073 _136_ trim[4] 7.1e-20
C12074 _101_ net24 0.00937f
C12075 cal_itt\[0\] a_10405_9295# 6.21e-19
C12076 a_4443_9295# clknet_0_clk 1.13e-19
C12077 a_1867_3317# a_2601_3285# 0.0701f
C12078 _019_ a_4696_8207# 5.18e-20
C12079 _084_ _101_ 1.37e-19
C12080 a_9761_8457# VPWR 0.00241f
C12081 a_11233_4405# VPWR 0.555f
C12082 cal_itt\[2\] _002_ 0.0339f
C12083 _078_ a_1769_11305# 2.97e-20
C12084 net13 a_4131_8207# 0.00303f
C12085 net46 _110_ 0.393f
C12086 cal_count\[0\] a_12061_7669# 4.99e-21
C12087 a_13142_8725# net2 3.73e-21
C12088 net16 a_12723_4943# 1.21e-20
C12089 a_11141_6031# a_12231_6005# 0.0424f
C12090 _032_ a_10207_1679# 3.71e-19
C12091 a_11709_6273# a_11491_6031# 0.21f
C12092 a_7140_2223# ctln[6] 1.07e-21
C12093 net52 clknet_0_clk 0.119f
C12094 trim_mask\[1\] a_14193_3285# 7.01e-19
C12095 net53 a_4222_10205# 2.16e-19
C12096 a_448_10357# a_561_9845# 2.68e-19
C12097 _095_ a_3057_4719# 0.00346f
C12098 a_2857_5461# _097_ 2.21e-19
C12099 _072_ a_7459_7663# 0.00299f
C12100 net4 a_8298_5487# 0.0209f
C12101 _030_ _055_ 1.99e-20
C12102 net44 mask\[2\] 0.00622f
C12103 net40 a_12599_3615# 1.77e-21
C12104 _036_ _041_ 0.00246f
C12105 net12 a_7351_8041# 3.3e-19
C12106 clknet_2_3__leaf_clk _107_ 0.00643f
C12107 a_2225_7663# VPWR 0.194f
C12108 net46 a_12778_3677# 0.00426f
C12109 a_1467_7923# a_1651_7093# 0.00444f
C12110 _108_ a_14715_3615# 0.0051f
C12111 _106_ a_8749_3317# 7.03e-20
C12112 net16 _056_ 0.00292f
C12113 _016_ VPWR 0.714f
C12114 _074_ _041_ 0.0864f
C12115 _074_ _010_ 0.0801f
C12116 net29 ctlp[1] 5.91e-19
C12117 net46 a_10699_5487# 4.03e-20
C12118 net46 a_12148_4777# 0.252f
C12119 a_1019_6397# VPWR 0.143f
C12120 calibrate a_6763_5193# 0.113f
C12121 _045_ VPWR 0.513f
C12122 state\[0\] a_3224_2601# 1.75e-19
C12123 net34 a_15299_3311# 0.0121f
C12124 net4 a_10111_1679# 3.88e-20
C12125 net13 a_5998_11471# 2.21e-20
C12126 clknet_2_3__leaf_clk a_12900_7663# 9.51e-21
C12127 a_2033_3317# a_2491_3311# 0.0346f
C12128 net37 a_15054_5193# 3.96e-19
C12129 a_7891_3617# a_7223_2465# 6.84e-19
C12130 a_7715_3285# a_7184_2339# 2.79e-21
C12131 a_7010_3311# a_7379_2197# 7.88e-19
C12132 trim_val\[3\] _057_ 0.0206f
C12133 net37 trim_val\[1\] 8.1e-20
C12134 _090_ a_4175_4943# 6.74e-20
C12135 cal_itt\[1\] a_10990_7485# 1.88e-19
C12136 a_4680_6031# _092_ 0.00126f
C12137 a_4696_8207# VPWR 0.294f
C12138 a_745_12021# net43 0.0393f
C12139 clknet_2_1__leaf_clk mask\[7\] 0.00293f
C12140 clknet_2_0__leaf_clk net30 1.38f
C12141 net31 trim_mask\[1\] 4.83e-19
C12142 net44 a_6428_7119# 6.13e-19
C12143 _014_ a_2601_3285# 0.00576f
C12144 net19 a_9103_2601# 8.45e-19
C12145 a_5515_6005# _059_ 4.91e-20
C12146 _067_ VPWR 0.829f
C12147 cal_count\[0\] a_15159_9269# 7.71e-19
C12148 net14 _004_ 0.00343f
C12149 _064_ _119_ 0.0152f
C12150 _111_ a_11488_4765# 9.03e-20
C12151 clknet_2_1__leaf_clk a_3977_10217# 8.36e-20
C12152 a_2953_7119# a_3748_6281# 4.88e-19
C12153 _062_ state\[2\] 2.69e-21
C12154 net47 a_14249_8725# 1.83e-20
C12155 _051_ a_8307_4719# 6.49e-19
C12156 mask\[0\] a_3529_6281# 4.5e-19
C12157 net19 net47 0.152f
C12158 net16 net35 0.0519f
C12159 _033_ a_8749_3317# 0.259f
C12160 a_8583_3317# a_9317_3285# 0.0532f
C12161 net50 a_10373_1679# 2.13e-19
C12162 a_7527_4631# _104_ 1.02e-19
C12163 cal_itt\[0\] a_8949_6281# 0.066f
C12164 _110_ a_11343_3317# 5.55e-20
C12165 a_14564_6397# a_15023_6031# 0.00133f
C12166 _092_ a_7190_3855# 6.21e-19
C12167 _063_ a_9889_6873# 1.54e-19
C12168 _023_ VPWR 0.916f
C12169 mask\[7\] a_2368_9955# 2.69e-19
C12170 net13 net30 0.0102f
C12171 a_6428_7119# clk 7.3e-22
C12172 _025_ a_12533_3689# 2.82e-21
C12173 net22 a_1476_6031# 0.0601f
C12174 a_13142_8359# a_13557_8457# 3.15e-19
C12175 _005_ result[2] 4.79e-21
C12176 _028_ a_8491_2229# 5.1e-19
C12177 a_395_7119# _004_ 2.88e-20
C12178 a_561_7119# a_395_6031# 6.5e-21
C12179 a_2143_2229# clk 0.00834f
C12180 _090_ a_4576_3427# 1.5e-21
C12181 clknet_2_2__leaf_clk VPWR 4.34f
C12182 net19 a_8820_6005# 0.00424f
C12183 a_8657_2229# a_9747_2527# 0.0424f
C12184 a_9225_2197# a_9007_2601# 0.21f
C12185 _038_ a_11396_6031# 0.186f
C12186 a_6983_10217# a_7548_10217# 7.99e-20
C12187 a_10975_6031# a_11599_6397# 9.73e-19
C12188 net45 a_4709_2773# 4.09e-21
C12189 a_5496_12131# _009_ 2.08e-21
C12190 _084_ a_6375_12021# 0.0128f
C12191 _001_ a_10990_7485# 6.85e-20
C12192 net55 _050_ 0.128f
C12193 net13 a_5221_9295# 5.18e-19
C12194 a_763_8757# a_2019_9055# 0.0436f
C12195 net47 cal_itt\[1\] 0.00158f
C12196 net34 trim[4] 0.0953f
C12197 _123_ a_12249_7663# 0.0144f
C12198 _053_ _119_ 0.00168f
C12199 a_1651_7093# a_2787_7119# 2.4e-19
C12200 a_816_7119# a_1007_7119# 4.61e-19
C12201 _045_ net27 6.13e-19
C12202 a_816_10205# VPWR 0.08f
C12203 net2 a_14335_7895# 0.00997f
C12204 mask\[1\] a_911_7119# 1.21e-19
C12205 _013_ VPWR 0.491f
C12206 a_8583_3317# a_9773_3689# 2.56e-19
C12207 _096_ a_3273_4943# 2.67e-20
C12208 net9 a_12454_8041# 7.81e-19
C12209 net4 _015_ 0.0171f
C12210 _101_ a_4801_10159# 2.72e-19
C12211 a_4815_3031# clk 2.62e-20
C12212 net55 _052_ 0.0806f
C12213 _035_ _124_ 0.00385f
C12214 net46 a_13091_4943# 0.331f
C12215 a_3748_6281# a_2857_5461# 0.0126f
C12216 net16 net38 0.0476f
C12217 cal_itt\[1\] a_8820_6005# 0.0396f
C12218 a_4995_7119# a_4775_6031# 0.00143f
C12219 net53 a_7164_11293# 7.43e-19
C12220 a_1095_12393# a_1313_10901# 3.66e-20
C12221 net55 _098_ 0.0966f
C12222 net16 _061_ 2.82e-19
C12223 a_9471_9269# _070_ 2.2e-20
C12224 a_4863_4917# _100_ 3.23e-20
C12225 _104_ a_9826_3311# 3.05e-19
C12226 net33 a_13625_3317# 1.54e-19
C12227 trim_mask\[0\] a_13869_4943# 8.96e-19
C12228 _050_ a_7715_3285# 0.0617f
C12229 state\[2\] a_5524_1679# 0.00311f
C12230 a_8215_9295# _000_ 0.162f
C12231 a_4131_8207# a_4239_8573# 0.0572f
C12232 net28 ctlp[1] 3.32e-19
C12233 net52 a_1830_10205# 5.5e-20
C12234 a_10005_6031# a_10055_5487# 3.63e-19
C12235 cal_count\[2\] a_12824_7663# 1.2e-20
C12236 net15 a_2309_2229# 0.0174f
C12237 a_1201_3855# valid 1.33e-19
C12238 a_9003_3829# a_8583_3317# 0.00922f
C12239 net40 a_11016_6691# 2.83e-21
C12240 clknet_2_2__leaf_clk a_9478_4105# 5.17e-20
C12241 _072_ a_6523_7119# 1.35e-19
C12242 a_11233_4405# _104_ 1.35e-19
C12243 _094_ a_4091_5309# 4.06e-19
C12244 net47 _001_ 0.0228f
C12245 _074_ a_561_6031# 0.0168f
C12246 _081_ a_1129_7361# 9.1e-22
C12247 a_4165_11989# _078_ 6.56e-20
C12248 a_1651_10143# net25 0.129f
C12249 _051_ a_6822_4399# 1.34e-21
C12250 clknet_2_3__leaf_clk a_11587_6031# 0.00133f
C12251 clknet_2_1__leaf_clk a_8105_10383# 0.00196f
C12252 _042_ cal_itt\[0\] 1.18e-20
C12253 a_8381_9295# _065_ 1.73e-20
C12254 trim_mask\[1\] a_14083_3311# 0.00123f
C12255 _052_ a_7715_3285# 0.0801f
C12256 _007_ a_1476_10217# 9.3e-21
C12257 net16 a_13257_4943# 0.0169f
C12258 net27 _023_ 2.27e-19
C12259 _078_ _019_ 5.23e-20
C12260 a_7843_3677# clk 7.46e-19
C12261 mask\[3\] a_4609_9295# 0.627f
C12262 VPWR ctln[2] 0.182f
C12263 a_5340_6031# a_5449_6031# 0.00742f
C12264 net45 a_2288_3677# 7.54e-19
C12265 a_9443_6059# en_co_clk 0.0101f
C12266 a_5515_6005# a_5694_6031# 0.0074f
C12267 a_4425_6031# _092_ 5.56e-19
C12268 clknet_2_0__leaf_clk state\[0\] 2.17e-20
C12269 a_1129_4373# a_855_4105# 3.84e-19
C12270 _108_ _047_ 0.00591f
C12271 _078_ a_1493_11721# 0.05f
C12272 net45 a_7310_2223# 0.169f
C12273 net43 a_7613_8029# 0.0019f
C12274 net32 a_14540_3689# 5.89e-19
C12275 a_15083_4659# _055_ 6.66e-22
C12276 a_6541_12021# a_6909_10933# 7.32e-21
C12277 _039_ a_1638_6397# 3.69e-19
C12278 _114_ net8 3.77e-19
C12279 _122_ a_11141_6031# 5.13e-19
C12280 clknet_2_1__leaf_clk a_6261_11247# 2.72e-19
C12281 _064_ a_9225_2197# 1.87e-21
C12282 _118_ a_10188_4105# 0.0224f
C12283 net13 state\[2\] 0.127f
C12284 net34 _057_ 0.00351f
C12285 net26 a_8839_9661# 1.01e-19
C12286 _029_ a_12599_3615# 5.83e-21
C12287 _063_ a_11141_6031# 1.35e-20
C12288 _050_ _093_ 2.32e-20
C12289 _065_ clknet_0_clk 0.288f
C12290 en_co_clk a_5087_3855# 0.00156f
C12291 a_2755_2601# VPWR 1.75e-20
C12292 clknet_2_3__leaf_clk trim_mask\[4\] 1.03e-21
C12293 _078_ a_6467_9845# 2.01e-19
C12294 _101_ a_6181_10383# 0.00599f
C12295 mask\[4\] a_8215_9295# 9.47e-20
C12296 _087_ _088_ 4.44e-20
C12297 net13 state\[0\] 0.143f
C12298 _058_ trim_mask\[2\] 0.00127f
C12299 a_3431_12021# a_3947_11305# 8.17e-21
C12300 a_911_4777# cal 0.00152f
C12301 a_7569_7637# a_7723_6807# 1.9e-20
C12302 a_4443_1679# clk 0.0539f
C12303 trim_mask\[0\] a_8307_4943# 0.00833f
C12304 net43 a_5535_8181# 3.21e-20
C12305 net9 a_12430_7663# 6.51e-19
C12306 a_4512_12393# _084_ 1.37e-20
C12307 mask\[6\] a_5496_12131# 0.193f
C12308 _088_ a_6519_3829# 0.0908f
C12309 a_9572_2601# a_9761_1679# 1.74e-20
C12310 a_13356_7369# _136_ 6.7e-20
C12311 cal_itt\[2\] a_8389_5193# 7.66e-20
C12312 net9 a_13016_9117# 2.24e-19
C12313 _083_ _041_ 3.53e-21
C12314 a_15299_6575# trim[4] 0.00118f
C12315 _078_ VPWR 4.55f
C12316 a_10864_7387# a_13142_7271# 4.02e-20
C12317 net14 result[2] 6.6e-20
C12318 a_11059_7356# a_11204_7485# 0.0572f
C12319 a_10903_7261# a_11622_7485# 0.0826f
C12320 _065_ a_6198_8207# 0.00117f
C12321 net45 _090_ 1.49e-20
C12322 _065_ a_10699_5487# 0.0274f
C12323 _110_ a_9826_3311# 1.39e-19
C12324 _060_ a_5731_4943# 0.00137f
C12325 _054_ a_7939_3855# 0.23f
C12326 net43 _082_ 0.00876f
C12327 net19 _072_ 7.43e-19
C12328 net46 a_11057_4105# 2.51e-20
C12329 _087_ a_6519_4631# 5.14e-20
C12330 a_455_8181# a_448_6549# 9.71e-21
C12331 trim_mask\[0\] a_8298_2767# 4.42e-20
C12332 a_14540_3689# VPWR 0.293f
C12333 _078_ a_5699_9269# 0.0128f
C12334 net2 a_13441_6281# 0.00683f
C12335 a_2869_11247# VPWR 4.28e-19
C12336 mask\[0\] a_1493_5487# 0.0502f
C12337 a_1764_10383# result[4] 1.3e-20
C12338 a_11233_4405# _110_ 6.59e-21
C12339 net4 _041_ 0.0577f
C12340 a_6519_4631# a_6519_3829# 0.0132f
C12341 net19 _068_ 0.276f
C12342 _062_ _118_ 0.0742f
C12343 a_4775_6031# a_4863_4917# 1.39e-19
C12344 net4 a_7184_2339# 1.66e-19
C12345 clknet_2_2__leaf_clk _104_ 0.0678f
C12346 a_579_12021# a_1660_11305# 2.25e-20
C12347 a_11116_8983# a_10990_7485# 9.16e-22
C12348 _034_ _050_ 2.82e-20
C12349 a_6891_12393# ctlp[6] 9.17e-19
C12350 _124_ a_11987_8757# 2.96e-21
C12351 _013_ a_2383_3689# 9.07e-19
C12352 a_15023_5487# trim[1] 9.24e-19
C12353 a_10138_5807# _118_ 9.57e-20
C12354 _099_ a_6519_4631# 5.38e-19
C12355 a_395_7119# result[2] 9.42e-19
C12356 net14 a_2309_2229# 5.64e-19
C12357 net14 a_1191_11305# 0.00129f
C12358 net9 a_12424_3689# 0.0101f
C12359 mask\[7\] result[4] 5.8e-20
C12360 _095_ a_3891_4943# 0.0579f
C12361 a_2857_5461# a_4308_4917# 4.09e-20
C12362 _042_ a_7723_10143# 7.31e-20
C12363 a_4043_10143# a_3840_8867# 0.00127f
C12364 net15 a_4609_1679# 7.1e-21
C12365 net18 a_9871_10383# 0.111f
C12366 net47 a_11394_9509# 0.143f
C12367 clknet_2_1__leaf_clk _080_ 5.41e-19
C12368 _075_ a_7210_5807# 1.97e-19
C12369 a_8381_9295# _067_ 9.32e-21
C12370 net29 net15 0.0176f
C12371 _072_ cal_itt\[1\] 2.1e-20
C12372 a_14604_3017# a_14099_3017# 0.00615f
C12373 a_11067_3017# a_11149_2767# 0.00393f
C12374 a_1660_11305# a_2869_10927# 1.24e-19
C12375 net52 a_1822_10927# 5.26e-21
C12376 net4 a_9839_3615# 5.48e-19
C12377 a_11233_4405# a_12148_4777# 0.125f
C12378 a_10699_5487# a_11233_4405# 5.93e-20
C12379 net19 net46 0.00497f
C12380 clknet_0_clk _016_ 7.76e-21
C12381 _053_ calibrate 0.145f
C12382 _063_ net42 0.00633f
C12383 a_3597_10933# VPWR 0.591f
C12384 clknet_2_0__leaf_clk a_911_6031# 6.3e-19
C12385 trim_val\[0\] a_13459_3317# 2.17e-20
C12386 net43 a_1007_10217# 0.00168f
C12387 _092_ _103_ 0.0584f
C12388 _068_ cal_itt\[1\] 0.171f
C12389 net13 _100_ 0.00763f
C12390 a_6835_7669# _049_ 5.51e-20
C12391 a_395_4405# a_1019_4399# 9.73e-19
C12392 a_4167_6575# net30 0.0273f
C12393 net15 _040_ 0.0131f
C12394 a_8298_5487# _064_ 0.0533f
C12395 a_1467_7923# a_2225_7983# 5.73e-20
C12396 a_4959_1679# ctln[7] 1.28e-19
C12397 a_561_4405# a_911_4777# 0.229f
C12398 _042_ a_1476_10217# 1.99e-19
C12399 a_4687_11231# a_4609_9295# 1.15e-20
C12400 _120_ en_co_clk 0.129f
C12401 net33 a_14894_3677# 7.82e-19
C12402 _079_ a_1493_5487# 0.0909f
C12403 _048_ a_7800_4631# 0.0208f
C12404 net44 a_4609_9295# 0.0319f
C12405 clknet_2_0__leaf_clk _012_ 0.00553f
C12406 a_9195_10357# clknet_2_3__leaf_clk 7.04e-22
C12407 _059_ a_5087_3855# 0.00398f
C12408 _041_ a_11479_9117# 0.00175f
C12409 a_12612_8725# a_13184_9117# 1.57e-19
C12410 net41 a_3057_3689# 8.27e-19
C12411 _042_ _007_ 0.00131f
C12412 net47 a_11116_8983# 2.22e-19
C12413 trim_val\[0\] _109_ 0.00388f
C12414 a_14471_591# trim[3] 6.33e-19
C12415 net15 a_3431_12021# 0.00107f
C12416 net27 _078_ 0.445f
C12417 a_5515_6005# _107_ 2.03e-19
C12418 clknet_2_3__leaf_clk _128_ 1.4e-20
C12419 clknet_2_0__leaf_clk a_5691_7637# 0.005f
C12420 net16 net40 0.129f
C12421 net52 a_4512_11305# 2.36e-21
C12422 clknet_0_clk _067_ 0.00189f
C12423 net12 a_4959_1679# 7.82e-19
C12424 net55 a_8389_5193# 0.0133f
C12425 ctlp[6] ctlp[5] 1.96e-20
C12426 a_12061_7669# cal_count\[2\] 1.45e-19
C12427 net47 net9 0.131f
C12428 a_5502_6397# VPWR 7.85e-19
C12429 net30 _028_ 6.27e-21
C12430 a_14335_2442# VPWR 0.231f
C12431 net4 a_9207_3311# 0.00382f
C12432 _072_ _001_ 1.65e-20
C12433 _119_ a_9664_3689# 3.82e-20
C12434 a_7256_8029# a_7447_8041# 4.61e-19
C12435 net8 VPWR 0.557f
C12436 _062_ a_10137_4943# 0.0522f
C12437 _076_ a_6419_8207# 6.37e-19
C12438 _061_ clkc 4.9e-19
C12439 state\[1\] net41 0.00658f
C12440 clknet_2_1__leaf_clk a_6885_8372# 0.012f
C12441 _096_ a_4091_5309# 2.5e-20
C12442 _049_ a_5515_6005# 0.0176f
C12443 _068_ _001_ 1.8e-20
C12444 net4 _002_ 7.04e-21
C12445 _105_ a_8473_5193# 0.00869f
C12446 a_7571_4943# _106_ 1.27e-20
C12447 _067_ a_10699_5487# 0.00366f
C12448 _053_ a_8298_5487# 0.133f
C12449 a_10329_1921# a_10676_1679# 0.0512f
C12450 net15 _048_ 0.0177f
C12451 trim_mask\[1\] a_12599_3615# 0.0871f
C12452 _119_ a_10689_2223# 1.16e-20
C12453 a_13607_1513# a_13703_1513# 0.0138f
C12454 clknet_2_2__leaf_clk _110_ 1.01f
C12455 a_6191_12559# net20 0.111f
C12456 net4 _050_ 0.773f
C12457 a_8993_9295# VPWR 2.3e-19
C12458 net40 a_10699_3311# 5.9e-22
C12459 cal_count\[3\] a_10245_5193# 9.2e-19
C12460 clknet_0_clk clknet_2_2__leaf_clk 0.0836f
C12461 a_4167_11471# a_3947_11305# 1.05e-19
C12462 _121_ _092_ 1.03e-21
C12463 net9 a_11435_2229# 0.0128f
C12464 a_6909_10933# a_7723_10143# 4.08e-19
C12465 a_13825_1109# trim[3] 9.11e-20
C12466 a_6541_12021# mask\[5\] 1.47e-20
C12467 a_2143_2229# a_3399_2527# 0.0435f
C12468 a_2309_2229# a_2659_2601# 0.217f
C12469 a_14347_4917# trim[4] 4.74e-19
C12470 net22 _039_ 0.412f
C12471 mask\[4\] a_7902_10205# 0.00185f
C12472 _070_ _069_ 0.13f
C12473 clknet_2_2__leaf_clk a_12778_3677# 2.16e-19
C12474 clknet_2_0__leaf_clk a_4775_6031# 0.00278f
C12475 a_1313_10901# a_1461_10357# 1.8e-19
C12476 clknet_2_3__leaf_clk a_8949_9537# 0.0429f
C12477 net37 net5 0.00267f
C12478 _070_ a_8022_7119# 0.00201f
C12479 net27 a_3597_10933# 9.9e-20
C12480 net13 a_5089_10159# 6.47e-19
C12481 net46 a_11067_4405# 0.3f
C12482 net43 net22 2.63e-19
C12483 a_4043_10143# a_4131_8207# 1.26e-21
C12484 net55 a_7891_3617# 2.98e-20
C12485 a_6541_12021# a_6999_12015# 0.0346f
C12486 net44 a_7565_12393# 6.03e-19
C12487 net34 a_13625_3317# 2.12e-20
C12488 clknet_2_1__leaf_clk a_1835_11231# 4.23e-20
C12489 a_11204_7485# a_11016_6691# 3e-20
C12490 _101_ a_7164_11293# 4.94e-21
C12491 net4 _052_ 8.16e-20
C12492 net29 a_1822_12015# 1.14e-19
C12493 _004_ VPWR 0.353f
C12494 a_10699_5487# clknet_2_2__leaf_clk 2.3e-20
C12495 clknet_2_2__leaf_clk a_12148_4777# 3.11e-19
C12496 clknet_2_3__leaf_clk a_11895_7669# 0.24f
C12497 net50 _058_ 0.0378f
C12498 trim_mask\[0\] a_15083_4659# 7.18e-21
C12499 net29 net25 7.99e-20
C12500 net21 a_3947_11305# 0.00162f
C12501 a_8820_6005# a_8949_6031# 0.0101f
C12502 a_2857_5461# _090_ 0.00855f
C12503 net4 a_9602_6614# 7.36e-19
C12504 trim_mask\[1\] a_11057_3855# 0.00217f
C12505 a_14377_7983# a_14422_7093# 4.23e-20
C12506 _018_ a_2815_9447# 0.116f
C12507 a_5455_4943# net42 4.92e-20
C12508 net14 net29 0.0335f
C12509 net28 net15 0.0994f
C12510 _072_ a_7916_8041# 0.059f
C12511 _065_ a_6523_7119# 2.85e-21
C12512 state\[0\] a_2948_3689# 0.00316f
C12513 a_6906_2355# a_7140_2223# 0.00645f
C12514 a_7379_2197# a_7617_2589# 0.00171f
C12515 net12 a_5878_1679# 3.18e-19
C12516 a_7223_2465# a_7942_2223# 0.0902f
C12517 a_7184_2339# a_7689_2589# 2.28e-19
C12518 a_6467_9845# a_6888_10205# 0.0897f
C12519 a_7001_7669# VPWR 0.524f
C12520 net13 a_4775_6031# 0.014f
C12521 _085_ a_2787_10927# 1.1e-19
C12522 VPWR ctln[7] 0.391f
C12523 net47 a_12436_9129# 0.206f
C12524 _125_ a_15023_8751# 0.0129f
C12525 _108_ net49 0.119f
C12526 _068_ a_7916_8041# 1.61e-21
C12527 clknet_2_3__leaf_clk a_11491_6031# 0.0431f
C12528 a_9503_4399# a_9099_3689# 8.17e-20
C12529 net12 a_6467_9845# 7.12e-21
C12530 a_7715_3285# a_7891_3617# 0.185f
C12531 a_2828_12131# a_2910_12131# 0.00477f
C12532 a_3597_12021# a_4043_12393# 2.28e-19
C12533 a_10752_565# ctln[4] 0.159f
C12534 clknet_2_0__leaf_clk a_3411_7485# 0.00604f
C12535 net43 a_3133_11247# 6.22e-20
C12536 net16 a_15023_12559# 0.00133f
C12537 a_14335_7895# a_14733_7983# 0.00369f
C12538 a_12900_7663# a_12824_7663# 0.00212f
C12539 _084_ a_7456_12393# 1.83e-20
C12540 a_15259_7637# _133_ 1.69e-19
C12541 _132_ a_14377_7983# 0.067f
C12542 a_561_7119# a_911_6031# 1.91e-19
C12543 a_6888_10205# VPWR 0.0796f
C12544 net12 VPWR 1.57f
C12545 _113_ trim_mask\[2\] 2.11e-19
C12546 clknet_2_1__leaf_clk a_5578_12131# 0.00148f
C12547 a_1497_8725# a_1844_9129# 0.0512f
C12548 trim_mask\[1\] a_10543_2455# 6.42e-20
C12549 _050_ a_6763_5193# 0.148f
C12550 a_12924_8029# VPWR 4.86e-19
C12551 a_4801_9839# a_4609_9295# 3.84e-19
C12552 a_13715_1135# trim[3] 5.61e-20
C12553 a_2815_9447# mask\[1\] 4.05e-20
C12554 _006_ a_1497_8725# 6.55e-19
C12555 state\[2\] _028_ 0.00598f
C12556 a_6467_9845# a_6983_10217# 0.111f
C12557 _008_ a_7201_9813# 6.55e-19
C12558 a_11141_6031# a_13111_6031# 2.39e-19
C12559 net12 a_5699_9269# 0.00904f
C12560 net4 a_9125_4943# 1.27e-19
C12561 net46 a_13512_1501# 0.0181f
C12562 net53 a_6099_10633# 0.242f
C12563 net55 _087_ 0.0879f
C12564 a_11067_4405# a_11149_3017# 6.37e-21
C12565 net44 a_6181_10633# 2.66e-20
C12566 a_5340_6031# VPWR 0.288f
C12567 _092_ a_3273_4943# 0.0974f
C12568 a_3411_9839# clknet_2_0__leaf_clk 4.04e-20
C12569 net43 a_4165_10901# 0.17f
C12570 _094_ net30 2.27e-19
C12571 net55 a_6519_3829# 3.8e-20
C12572 a_6885_8372# a_6485_8181# 0.00391f
C12573 a_6056_8359# net51 0.00203f
C12574 a_6763_5193# _052_ 2.78e-19
C12575 mask\[7\] mask\[6\] 0.224f
C12576 net20 a_6796_12381# 0.0146f
C12577 a_6983_10217# VPWR 0.211f
C12578 a_745_10933# a_1313_10901# 0.186f
C12579 net47 a_11508_9295# 0.0028f
C12580 _000_ _041_ 0.2f
C12581 trim_val\[0\] a_14655_4399# 0.0344f
C12582 a_14552_9071# a_14467_8751# 1.48e-19
C12583 a_1867_3317# clk 2.74e-19
C12584 _096_ a_4886_4399# 3.87e-19
C12585 _098_ a_6763_5193# 0.00811f
C12586 net55 _099_ 0.103f
C12587 net37 a_15023_6031# 0.0139f
C12588 trim_mask\[3\] a_11435_2229# 0.00556f
C12589 _097_ a_855_4105# 7.99e-20
C12590 a_14715_3615# _056_ 1.36e-20
C12591 cal_count\[3\] a_8473_5193# 5.67e-19
C12592 clknet_2_2__leaf_clk a_13091_4943# 0.262f
C12593 a_3852_12381# VPWR 0.0836f
C12594 a_10543_2455# a_10977_2543# 0.00393f
C12595 _062_ a_8820_6005# 0.125f
C12596 a_9460_6807# a_9443_6059# 1.86e-19
C12597 net19 _065_ 0.00893f
C12598 net44 _051_ 0.00365f
C12599 _081_ mask\[1\] 0.274f
C12600 net15 net21 1.66e-20
C12601 _078_ clknet_0_clk 3.17e-20
C12602 _017_ a_3317_8207# 1.97e-19
C12603 net2 a_12056_6031# 2.97e-19
C12604 a_1651_10143# VPWR 0.392f
C12605 net26 a_7939_10383# 4.04e-19
C12606 _114_ trim[2] 9.22e-20
C12607 _095_ a_395_4405# 5.58e-22
C12608 a_9503_4399# trim_val\[4\] 3.83e-19
C12609 net37 net46 1.7e-19
C12610 a_5496_12131# ctlp[7] 0.00111f
C12611 net4 a_10747_8970# 1.58e-19
C12612 a_9463_8725# _124_ 2.13e-19
C12613 a_7800_4631# a_7758_4759# 1.84e-19
C12614 a_6885_8372# a_6007_7119# 7.75e-22
C12615 a_7190_3855# a_7010_3311# 4.36e-19
C12616 a_6056_8359# _003_ 4.11e-20
C12617 _126_ _125_ 0.272f
C12618 trim_mask\[0\] a_9369_4105# 0.0472f
C12619 a_1830_7119# VPWR 4.04e-19
C12620 _074_ a_1129_4373# 0.00545f
C12621 a_8551_10383# VPWR 7.45e-19
C12622 clknet_2_3__leaf_clk _061_ 0.00543f
C12623 a_2787_7119# net30 1.48e-19
C12624 _106_ _058_ 5.05e-19
C12625 _049_ a_4815_3031# 6.23e-21
C12626 net16 _029_ 4.6e-19
C12627 net27 net12 0.331f
C12628 a_14193_3285# a_14071_3689# 3.16e-19
C12629 a_13975_3689# a_13880_3677# 0.0498f
C12630 a_9003_3829# a_9662_3855# 0.00414f
C12631 mask\[3\] _082_ 0.0846f
C12632 cal_itt\[0\] a_9405_9295# 1.13e-19
C12633 net40 clkc 1.65e-19
C12634 net2 a_13279_8207# 0.0383f
C12635 net28 net14 0.398f
C12636 trim_mask\[1\] a_13607_1513# 8.39e-22
C12637 _065_ cal_itt\[1\] 0.00318f
C12638 a_13703_4943# VPWR 0.00379f
C12639 _051_ clk 0.357f
C12640 net15 a_2033_3317# 2.68e-19
C12641 a_11601_2229# a_12516_2601# 0.125f
C12642 a_11435_2229# a_13415_2442# 8.25e-21
C12643 net22 a_1173_6031# 7.15e-19
C12644 net53 a_5423_9011# 3.34e-19
C12645 en_co_clk _051_ 0.00346f
C12646 a_1387_8751# _081_ 8.91e-20
C12647 _129_ a_15259_7637# 3.05e-19
C12648 a_15023_12559# trimb[3] 0.34f
C12649 mask\[4\] _041_ 1.8e-20
C12650 net47 a_13470_7663# 0.00218f
C12651 net35 a_14715_3615# 1.16e-19
C12652 _107_ a_7843_3677# 2.5e-19
C12653 _085_ a_3947_12393# 1.84e-19
C12654 _058_ a_14193_3285# 6.41e-19
C12655 net32 a_13459_3317# 7.72e-20
C12656 _013_ net41 0.107f
C12657 mask\[5\] a_7723_10143# 5.66e-20
C12658 a_6909_10933# _042_ 8.79e-20
C12659 _014_ clk 0.0041f
C12660 _136_ a_13512_4943# 0.00156f
C12661 net3 _060_ 0.0282f
C12662 a_9443_6059# _107_ 2.31e-19
C12663 a_14063_7093# _130_ 0.135f
C12664 clknet_2_0__leaf_clk a_3933_2767# 1.92e-20
C12665 net52 a_4995_7119# 4.86e-20
C12666 _051_ a_9084_4515# 4.76e-20
C12667 a_13008_7663# VPWR 0.00306f
C12668 net45 a_3667_3829# 6.11e-19
C12669 net9 net46 1.8f
C12670 _101_ a_2961_9545# 0.0133f
C12671 a_13256_9117# VPWR 1.86e-19
C12672 a_6197_6281# VPWR 0.00439f
C12673 a_14604_3017# trim[0] 5.41e-20
C12674 a_13519_4007# a_14335_4020# 3.49e-20
C12675 _085_ a_3425_11721# 0.0972f
C12676 VPWR result[2] 0.514f
C12677 trim_mask\[2\] a_10569_1109# 2.87e-21
C12678 a_4259_6031# net55 2.11e-19
C12679 a_13697_4373# a_13915_4399# 0.0821f
C12680 _124_ a_11258_9117# 2.88e-19
C12681 _058_ a_14000_4719# 1.18e-19
C12682 _049_ a_7843_3677# 7.02e-19
C12683 a_1660_11305# _101_ 6.61e-20
C12684 mask\[2\] a_5524_9295# 8.23e-21
C12685 net24 net45 2.76e-20
C12686 a_561_9845# a_1638_9839# 1.46e-19
C12687 _101_ mask\[0\] 0.115f
C12688 net16 a_13349_6031# 2.73e-19
C12689 net16 _123_ 0.036f
C12690 a_8657_2229# a_9595_1679# 0.00461f
C12691 _064_ a_9839_3615# 2.96e-19
C12692 a_6796_12381# a_6987_12393# 4.61e-19
C12693 a_395_9845# a_1019_9839# 9.73e-19
C12694 _056_ a_14099_1929# 9.9e-20
C12695 trim_val\[0\] trim[1] 0.00234f
C12696 a_8949_9537# a_8827_9295# 3.16e-19
C12697 net13 a_3933_2767# 1.79e-19
C12698 net43 a_7569_7637# 0.203f
C12699 _065_ _001_ 0.437f
C12700 _099_ _093_ 0.0555f
C12701 net31 _058_ 5.96e-20
C12702 _065_ a_11067_4405# 2.04e-20
C12703 _092_ a_11141_6031# 7.25e-19
C12704 net32 trim[2] 6.26e-20
C12705 clknet_2_1__leaf_clk a_3840_8867# 4.36e-21
C12706 en_co_clk a_5445_4399# 1.73e-19
C12707 _110_ a_14335_2442# 9.81e-20
C12708 a_6631_7485# VPWR 0.143f
C12709 _041_ _053_ 2.62e-20
C12710 _110_ net8 5.18e-21
C12711 a_13459_3317# VPWR 0.436f
C12712 net12 _104_ 0.034f
C12713 a_7088_7119# net30 6.43e-20
C12714 _053_ a_7184_2339# 1.48e-22
C12715 a_1129_4373# _093_ 1.4e-19
C12716 _133_ a_14485_7663# 0.00272f
C12717 a_2309_2229# VPWR 0.273f
C12718 a_1191_11305# VPWR 0.00132f
C12719 clknet_2_1__leaf_clk a_2971_8457# 0.00409f
C12720 _064_ a_10781_5487# 0.00114f
C12721 net44 a_7613_8029# 4.25e-19
C12722 clknet_2_2__leaf_clk a_11057_4105# 0.00629f
C12723 a_12061_7669# a_12900_7663# 0.0573f
C12724 a_10903_7261# _136_ 0.00313f
C12725 a_1651_6005# a_2313_6183# 0.0135f
C12726 a_10055_2767# a_10219_2045# 1.44e-19
C12727 net19 _067_ 0.0106f
C12728 _134_ a_13825_5185# 2.32e-19
C12729 a_579_12021# a_579_10933# 0.002f
C12730 _063_ net30 0.0247f
C12731 trim_mask\[0\] a_8307_4719# 0.0762f
C12732 net45 a_4883_6397# 6.88e-20
C12733 mask\[6\] a_6261_11247# 0.00163f
C12734 a_745_10933# result[5] 7.03e-19
C12735 a_2865_4460# _099_ 0.0595f
C12736 a_4609_1679# a_4959_1679# 0.217f
C12737 a_4443_1679# a_5699_1653# 0.0436f
C12738 _048_ a_7460_5807# 0.0814f
C12739 _109_ VPWR 0.355f
C12740 a_1476_4777# a_3388_4631# 7.92e-21
C12741 net9 a_11343_3317# 0.00722f
C12742 net46 a_10188_4105# 2.99e-19
C12743 net2 a_13607_4943# 1.14e-19
C12744 net9 a_11149_3017# 7.53e-20
C12745 a_911_4777# a_1019_4399# 0.0572f
C12746 a_14249_8725# a_14552_9071# 0.00138f
C12747 _001_ a_9761_8457# 0.0158f
C12748 a_5691_2741# VPWR 0.629f
C12749 _020_ a_7548_10217# 1.4e-20
C12750 a_14604_3017# a_15023_2767# 0.001f
C12751 net4 a_7891_3617# 3.44e-21
C12752 a_1660_11305# _102_ 0.00202f
C12753 net52 a_1203_10927# 1.99e-20
C12754 net3 a_4498_4373# 0.00234f
C12755 _136_ a_11845_4765# 1.89e-19
C12756 _051_ _059_ 0.0305f
C12757 _034_ _099_ 1.39e-21
C12758 net53 a_4871_8181# 4.06e-21
C12759 a_11067_4405# a_11233_4405# 0.863f
C12760 a_2143_7663# _005_ 7.7e-20
C12761 net18 a_11352_9661# 3.91e-19
C12762 net53 _076_ 0.0282f
C12763 net44 a_5535_8181# 0.00315f
C12764 a_14347_4917# a_13625_3317# 5.72e-21
C12765 _072_ _062_ 5.18e-20
C12766 calibrate a_395_4405# 0.00333f
C12767 net19 clknet_2_2__leaf_clk 0.125f
C12768 a_9871_10383# VPWR 0.246f
C12769 a_7524_2223# VPWR 0.144f
C12770 _067_ cal_itt\[1\] 0.258f
C12771 clknet_2_0__leaf_clk a_1651_4703# 0.00635f
C12772 _078_ a_1830_10205# 2.33e-19
C12773 _078_ a_2775_9071# 2.65e-19
C12774 VPWR trim[2] 0.606f
C12775 net30 _096_ 1.8e-20
C12776 mask\[2\] a_4036_8207# 1.38e-19
C12777 _068_ _062_ 0.0311f
C12778 net14 a_2033_3317# 3.78e-20
C12779 net15 a_2143_7663# 6.52e-19
C12780 a_5726_5807# VPWR 1.43e-19
C12781 _115_ a_13881_1653# 0.00215f
C12782 _048_ a_5363_4719# 0.00665f
C12783 net45 a_1129_6273# 0.166f
C12784 _002_ a_7447_8041# 0.00467f
C12785 a_9595_1679# a_10569_1109# 3.69e-19
C12786 _042_ a_4959_9295# 3.29e-20
C12787 a_9761_1679# a_10195_1354# 0.00452f
C12788 a_15023_9839# net40 2.1e-20
C12789 _036_ a_12341_8751# 0.148f
C12790 a_1313_11989# a_1822_12015# 2.6e-19
C12791 net43 a_4043_12393# 2.48e-19
C12792 _092_ net42 0.0793f
C12793 net46 trim_mask\[3\] 0.0635f
C12794 net16 trim_mask\[1\] 0.0189f
C12795 _122_ _134_ 0.084f
C12796 net14 a_1549_6794# 0.113f
C12797 net43 a_1476_10217# 0.257f
C12798 a_10903_7261# a_10861_7119# 2.56e-19
C12799 net52 a_3431_10933# 0.00612f
C12800 a_1660_11305# _022_ 4.8e-20
C12801 a_8455_10383# a_8551_10383# 0.0138f
C12802 net16 a_13142_8725# 8.18e-19
C12803 state\[0\] a_4617_3855# 6.15e-20
C12804 net26 a_6056_8359# 1.14e-21
C12805 net46 a_10689_2543# 1.02e-19
C12806 a_3110_3311# VPWR 7.19e-19
C12807 net29 a_1493_11721# 0.00958f
C12808 net43 _007_ 7.35e-19
C12809 _092_ a_4091_5309# 0.00143f
C12810 _091_ VPWR 0.348f
C12811 net1 a_1201_3855# 0.00105f
C12812 net14 a_1313_11989# 0.00489f
C12813 a_5997_10927# VPWR 0.204f
C12814 a_1099_12533# net43 0.0031f
C12815 a_12169_2197# VPWR 0.224f
C12816 _069_ net2 0.0612f
C12817 _070_ net51 1.36e-20
C12818 a_13880_3677# trim_val\[1\] 9.97e-20
C12819 net4 a_10005_6031# 0.005f
C12820 _119_ a_8583_3317# 0.0126f
C12821 _019_ _040_ 8.42e-20
C12822 net45 a_4677_7882# 0.0379f
C12823 a_9369_4105# a_8298_2767# 1.04e-20
C12824 _059_ a_5445_4399# 0.016f
C12825 a_3431_12021# a_4165_11989# 0.0535f
C12826 net2 a_8022_7119# 3.61e-20
C12827 clknet_2_1__leaf_clk a_6793_8970# 0.0024f
C12828 _049_ _120_ 0.0916f
C12829 net35 _047_ 2.85e-19
C12830 clknet_2_3__leaf_clk net40 0.00271f
C12831 _001_ _067_ 9.01e-19
C12832 _060_ a_5537_4105# 0.00175f
C12833 a_9595_1679# a_10329_1921# 0.0701f
C12834 _032_ a_9761_1679# 0.224f
C12835 _053_ _050_ 0.183f
C12836 a_5177_1921# a_5633_1679# 4.2e-19
C12837 a_5997_10927# a_5699_9269# 1.33e-21
C12838 _101_ a_6099_10633# 0.103f
C12839 net12 clknet_0_clk 0.0103f
C12840 a_395_7119# a_1549_6794# 0.0116f
C12841 _058_ a_14083_3311# 6.29e-19
C12842 a_10975_4105# trim_mask\[2\] 5.93e-21
C12843 trim_mask\[1\] a_10699_3311# 0.18f
C12844 a_11292_1251# _057_ 0.106f
C12845 _129_ a_14485_7663# 0.00335f
C12846 a_11987_8757# a_10903_7261# 2.67e-20
C12847 net18 net10 0.228f
C12848 net26 a_7710_9839# 4.38e-19
C12849 cal_itt\[3\] net42 2.24e-19
C12850 a_2857_5461# a_3667_3829# 5.09e-19
C12851 net4 _087_ 2.67e-20
C12852 net46 a_9195_3689# 1.79e-19
C12853 _089_ VPWR 0.255f
C12854 a_1095_11305# net26 2.32e-20
C12855 mask\[5\] _042_ 0.00943f
C12856 net22 a_1579_5807# 1.55e-19
C12857 _128_ a_13184_9117# 1.82e-19
C12858 a_14655_4399# net32 1.88e-19
C12859 net46 a_13415_2442# 0.0272f
C12860 _103_ a_7010_3311# 1.08e-20
C12861 a_7001_7669# a_7459_7663# 0.0346f
C12862 _064_ a_10872_1455# 8.95e-20
C12863 _034_ a_4259_6031# 0.139f
C12864 a_12520_7637# VPWR 0.25f
C12865 a_1651_6005# VPWR 0.389f
C12866 _053_ _052_ 0.0087f
C12867 net12 a_6198_8207# 1.76e-19
C12868 clknet_0_clk a_5340_6031# 8.64e-21
C12869 a_4609_1679# VPWR 0.291f
C12870 net16 a_14565_9295# 5.96e-19
C12871 net29 VPWR 1.12f
C12872 a_6375_12021# a_6197_12015# 5.89e-20
C12873 clknet_2_1__leaf_clk a_5998_11471# 2.53e-20
C12874 net50 a_10569_1109# 0.00491f
C12875 a_816_4765# VPWR 0.0865f
C12876 net29 a_1769_12393# 1.37e-19
C12877 _053_ _098_ 4.65e-21
C12878 clknet_2_2__leaf_clk a_11067_4405# 0.3f
C12879 a_8749_3317# a_10699_3311# 1.28e-19
C12880 trim_mask\[4\] a_7843_3677# 3.87e-19
C12881 a_937_4105# cal 0.00146f
C12882 net53 clknet_2_3__leaf_clk 1.23e-20
C12883 trim_mask\[0\] a_12323_4703# 0.129f
C12884 net45 a_4993_6273# 4.08e-19
C12885 trim_mask\[2\] a_13881_2741# 1.32e-20
C12886 trim_mask\[4\] a_11601_2229# 1.26e-19
C12887 a_3123_3615# a_2143_2229# 4.57e-20
C12888 a_2383_3689# a_2309_2229# 2.29e-20
C12889 cal_itt\[0\] _038_ 6.38e-20
C12890 net12 a_7459_7663# 3.15e-19
C12891 trim_mask\[3\] a_11149_3017# 0.00299f
C12892 _005_ a_1019_7485# 1.23e-20
C12893 _040_ VPWR 0.343f
C12894 _068_ a_8745_6895# 0.00437f
C12895 a_5694_6031# _051_ 3.32e-20
C12896 _065_ a_4995_7119# 0.024f
C12897 _113_ a_14193_3285# 7.33e-21
C12898 mask\[5\] a_7521_11293# 9.25e-20
C12899 net9 a_12059_2223# 0.00203f
C12900 a_1095_12393# result[7] 3.7e-20
C12901 net9 _065_ 3.57e-20
C12902 net16 _115_ 0.013f
C12903 net54 _060_ 0.214f
C12904 state\[2\] a_7104_3855# 8.2e-20
C12905 _107_ a_6822_4105# 2.25e-19
C12906 net18 a_11583_4777# 0.00215f
C12907 a_7916_8041# _067_ 7.47e-19
C12908 a_3431_12021# VPWR 0.441f
C12909 cal_itt\[0\] cal_count\[0\] 4.18e-21
C12910 net43 a_3977_7119# 4.13e-19
C12911 a_4043_7093# _034_ 1.22e-20
C12912 net50 a_10329_1921# 0.00471f
C12913 a_15023_1135# VPWR 0.421f
C12914 net27 a_5997_10927# 6.97e-20
C12915 a_7190_3855# _119_ 5.69e-21
C12916 mask\[1\] a_3781_8207# 0.402f
C12917 net43 a_1357_11293# 0.00316f
C12918 _101_ a_5423_9011# 0.0103f
C12919 a_6007_9839# _076_ 5.93e-20
C12920 _096_ state\[0\] 2.01e-19
C12921 a_14655_4399# VPWR 0.242f
C12922 a_11895_7669# a_12824_7663# 0.00159f
C12923 _037_ a_12430_7663# 1.08e-19
C12924 net52 clknet_2_0__leaf_clk 0.139f
C12925 net28 a_4165_11989# 0.022f
C12926 clknet_2_0__leaf_clk a_816_7119# 0.00154f
C12927 _125_ VPWR 0.441f
C12928 clknet_2_1__leaf_clk net30 2.02e-20
C12929 a_8767_11471# VPWR 0.293f
C12930 _094_ a_4775_6031# 0.038f
C12931 _049_ a_6822_4105# 2.38e-19
C12932 VPWR trimb[0] 0.581f
C12933 a_1461_10357# a_561_9845# 0.00844f
C12934 net55 _097_ 1.31e-20
C12935 net16 a_14335_7895# 1.68e-20
C12936 mask\[6\] a_1835_11231# 2.47e-19
C12937 a_7184_2339# a_7379_2197# 0.223f
C12938 a_7223_2465# a_7310_2223# 0.0623f
C12939 _026_ a_12516_2601# 3.46e-19
C12940 _048_ VPWR 2.55f
C12941 result[6] ctlp[0] 4.71e-19
C12942 net28 a_1493_11721# 0.0628f
C12943 mask\[5\] a_6909_10933# 5.97e-19
C12944 net31 _113_ 2.53e-20
C12945 net13 a_4443_9295# 0.0193f
C12946 net9 a_11233_4405# 9.64e-20
C12947 _051_ _108_ 1.4e-20
C12948 a_10219_2045# VPWR 0.145f
C12949 _014_ a_3399_2527# 1.29e-20
C12950 a_6375_12021# a_6099_10633# 3.88e-21
C12951 a_14379_6397# trim_mask\[0\] 5.9e-21
C12952 a_8673_10625# _043_ 2.03e-21
C12953 net47 a_9020_10383# 0.24f
C12954 clknet_2_2__leaf_clk a_13512_1501# 5.24e-19
C12955 net29 net27 0.284f
C12956 net43 _042_ 0.377f
C12957 net13 net52 0.0204f
C12958 net15 ctlp[1] 0.037f
C12959 net35 a_14334_5309# 8.41e-20
C12960 _128_ a_14733_9545# 2.33e-19
C12961 net43 a_7723_6807# 1.14e-20
C12962 a_13142_8359# a_13050_7637# 0.00813f
C12963 a_13715_5309# _058_ 9.61e-19
C12964 state\[1\] a_3224_2601# 0.00189f
C12965 _033_ a_8657_2229# 4.32e-20
C12966 net32 trim[1] 0.16f
C12967 _037_ a_10990_7485# 1.29e-19
C12968 a_561_6031# a_455_5747# 6.7e-19
C12969 a_1476_10217# a_2953_9845# 2.49e-20
C12970 _050_ a_3891_4943# 0.115f
C12971 net45 result[1] 3.22e-20
C12972 _038_ trim_mask\[0\] 3.83e-20
C12973 _082_ a_1184_9117# 1.16e-19
C12974 net3 a_4175_4943# 0.00123f
C12975 a_4165_11989# a_4167_11471# 0.00138f
C12976 a_3947_11305# a_3852_11293# 0.0498f
C12977 a_4165_10901# a_4043_11305# 3.16e-19
C12978 a_2921_2589# clk 2.74e-19
C12979 a_1191_12393# VPWR 4.68e-19
C12980 net46 a_10207_1679# 0.00482f
C12981 a_11599_6397# VPWR 0.133f
C12982 _134_ comp 1.07e-19
C12983 calibrate a_2283_4020# 0.0273f
C12984 _101_ a_2489_7983# 8.5e-19
C12985 _060_ a_4471_4007# 0.233f
C12986 a_4863_4917# state\[1\] 1.16e-21
C12987 net28 VPWR 2.08f
C12988 _131_ a_14282_7119# 0.00298f
C12989 net12 net41 5.07e-20
C12990 a_9839_3615# a_9664_3689# 0.234f
C12991 a_9099_3689# trim_mask\[2\] 1.15e-20
C12992 a_3431_12021# net27 3.51e-20
C12993 a_5177_9537# VPWR 0.214f
C12994 mask\[6\] a_5578_12131# 2.29e-19
C12995 net54 a_4498_4373# 0.172f
C12996 _096_ _100_ 0.0909f
C12997 net18 a_10975_6031# 0.017f
C12998 _062_ a_7527_4631# 1.75e-20
C12999 _110_ a_13459_3317# 6.35e-19
C13000 _107_ a_7677_4759# 2.25e-19
C13001 net28 a_1769_12393# 2.55e-20
C13002 a_11396_6031# a_11587_6031# 4.61e-19
C13003 net34 a_14471_591# 8.93e-19
C13004 a_10903_7261# cal_count\[3\] 8.79e-21
C13005 clknet_2_3__leaf_clk _071_ 7.99e-20
C13006 a_6793_8970# a_6007_7119# 2.16e-21
C13007 _076_ a_5363_7369# 2.71e-19
C13008 a_7001_7669# a_6523_7119# 0.00115f
C13009 trim_mask\[2\] a_12047_2601# 1.57e-19
C13010 trim_mask\[1\] a_11955_3689# 6.86e-21
C13011 a_6835_7669# a_7263_7093# 9.58e-19
C13012 net14 a_1276_565# 0.0251f
C13013 a_1677_9545# a_1763_9295# 2.42e-19
C13014 a_4609_9295# a_5524_9295# 0.125f
C13015 a_2815_9447# a_3249_9295# 0.00393f
C13016 a_4443_9295# a_4864_9295# 0.0931f
C13017 net50 a_10975_4105# 0.00768f
C13018 net21 a_4165_11989# 9.46e-19
C13019 net27 a_8767_11471# 0.00138f
C13020 a_12424_3689# a_13880_3677# 6.86e-21
C13021 net47 a_8731_9295# 0.155f
C13022 trim_mask\[3\] a_12059_2223# 6.01e-19
C13023 a_8298_5487# a_8473_5193# 0.00178f
C13024 a_10405_9295# cal_count\[0\] 1.45e-19
C13025 _104_ _089_ 0.00112f
C13026 a_3597_10933# a_4512_11305# 0.125f
C13027 _101_ a_4871_8181# 5.34e-21
C13028 _051_ a_9004_3677# 8.21e-21
C13029 _132_ a_15289_7119# 0.00948f
C13030 a_3303_10217# mask\[2\] 6.01e-19
C13031 net46 a_11753_6031# 0.00322f
C13032 _101_ _076_ 0.036f
C13033 a_10975_6031# a_12165_6031# 2.56e-19
C13034 _039_ a_1476_6031# 0.0336f
C13035 a_11141_6031# _136_ 0.0113f
C13036 _049_ a_7677_4759# 2.88e-19
C13037 _125_ a_14807_8359# 0.122f
C13038 _129_ a_12344_8041# 6.87e-21
C13039 _110_ _109_ 0.126f
C13040 a_6541_12021# net44 0.0322f
C13041 a_816_6031# result[0] 6.73e-19
C13042 a_579_12021# result[6] 0.00742f
C13043 VPWR trim[1] 0.488f
C13044 net14 a_1019_7485# 0.00291f
C13045 net47 _037_ 0.00229f
C13046 _058_ a_12599_3615# 0.0034f
C13047 _065_ _062_ 1.86e-19
C13048 net3 a_4576_3427# 7.88e-22
C13049 a_2787_7119# a_3411_7485# 9.73e-19
C13050 a_2953_7119# a_3208_7119# 0.0612f
C13051 a_3521_7361# a_3868_7119# 0.0512f
C13052 a_745_10933# a_561_9845# 3.85e-21
C13053 net43 a_1476_6031# 1.76e-19
C13054 _051_ _107_ 0.156f
C13055 net12 a_6523_7119# 0.00752f
C13056 net15 a_3333_2601# 2.97e-20
C13057 _004_ a_1137_5487# 0.0113f
C13058 _108_ a_11801_4373# 2.33e-19
C13059 a_929_8757# net23 6.13e-20
C13060 _050_ a_7379_2197# 0.00129f
C13061 a_7021_4105# VPWR 0.238f
C13062 _097_ _093_ 0.507f
C13063 net34 a_13825_1109# 5.32e-21
C13064 a_4425_6031# _095_ 0.00207f
C13065 net19 a_8993_9295# 6.71e-19
C13066 net9 clknet_2_2__leaf_clk 0.185f
C13067 a_4167_11471# VPWR 0.243f
C13068 _053_ a_11369_7119# 8.12e-19
C13069 a_911_10217# a_1019_9839# 0.0572f
C13070 a_1651_10143# a_1830_10205# 0.0074f
C13071 a_1476_10217# a_1585_10217# 0.00742f
C13072 net45 a_3339_2767# 0.181f
C13073 clknet_2_3__leaf_clk a_11244_9661# 0.0853f
C13074 a_12148_4777# _109_ 2.67e-20
C13075 _058_ a_12257_4777# 1.84e-19
C13076 _063_ _118_ 0.00299f
C13077 clknet_0_clk a_5726_5807# 4.75e-19
C13078 a_395_7119# a_1019_7485# 9.73e-19
C13079 a_561_7119# a_816_7119# 0.0604f
C13080 _049_ _051_ 0.0328f
C13081 a_13607_4943# a_13715_5309# 0.0572f
C13082 a_13257_4943# a_14334_5309# 1.46e-19
C13083 a_13091_4943# a_13703_4943# 0.00188f
C13084 net44 a_4871_6031# 1.79e-19
C13085 a_14172_4943# a_14972_5193# 5.3e-19
C13086 _052_ a_7379_2197# 2.78e-21
C13087 clknet_2_3__leaf_clk a_11204_7485# 6.03e-20
C13088 net14 a_1173_10205# 5.85e-19
C13089 _053_ a_8389_5193# 0.00481f
C13090 _074_ a_845_7663# 0.0012f
C13091 _134_ a_13111_6031# 7.21e-19
C13092 a_12516_2601# _031_ 8.91e-19
C13093 a_12169_2197# a_12678_2223# 2.6e-19
C13094 a_6743_10933# a_7164_11293# 0.0931f
C13095 _021_ a_6261_11247# 0.00133f
C13096 a_5455_4943# _100_ 1.35e-20
C13097 _049_ _014_ 1.21e-21
C13098 a_2865_4460# _097_ 8.1e-19
C13099 _082_ result[3] 5.94e-19
C13100 _099_ a_3057_4719# 0.114f
C13101 a_3388_4631# _014_ 7.24e-19
C13102 _065_ a_6198_8534# 0.00203f
C13103 a_3116_12533# a_3513_12809# 5.98e-20
C13104 a_13142_8359# VPWR 0.278f
C13105 a_15023_2223# trim[3] 6.66e-20
C13106 a_1835_12319# a_1660_12393# 0.234f
C13107 trim_val\[4\] trim_mask\[2\] 0.00455f
C13108 a_1095_12393# mask\[7\] 0.00299f
C13109 net28 net27 0.41f
C13110 net43 a_3597_12021# 0.0394f
C13111 _085_ a_3303_10217# 3.19e-20
C13112 cal_itt\[0\] a_9459_7895# 0.0715f
C13113 net21 VPWR 0.803f
C13114 _041_ a_3781_8207# 0.00174f
C13115 _110_ a_12169_2197# 7.05e-19
C13116 _090_ _088_ 1.46e-20
C13117 clknet_2_3__leaf_clk a_13349_6031# 0.0447f
C13118 a_4498_4373# a_4471_4007# 0.0115f
C13119 a_3817_4697# state\[1\] 3.95e-20
C13120 net2 a_13783_6183# 0.00226f
C13121 a_6007_7119# net30 6.46e-21
C13122 _067_ a_10188_4105# 3.4e-20
C13123 calibrate a_7190_3855# 0.0066f
C13124 clknet_2_3__leaf_clk _123_ 0.156f
C13125 net4 a_10864_7387# 8.89e-21
C13126 a_8657_2229# ctln[5] 1.07e-20
C13127 a_1476_10217# mask\[3\] 0.00101f
C13128 a_11895_7669# a_12061_7669# 0.779f
C13129 net19 a_7001_7669# 1.43e-20
C13130 _078_ a_5829_9839# 0.00526f
C13131 trim_mask\[0\] a_10270_4105# 9.24e-19
C13132 a_4871_6031# en_co_clk 4.18e-19
C13133 _007_ mask\[3\] 1.14e-19
C13134 cal_count\[0\] a_11258_8790# 0.00688f
C13135 _048_ _104_ 0.0872f
C13136 _086_ a_579_10933# 2.59e-20
C13137 a_3273_4943# a_3365_4943# 0.0606f
C13138 clknet_2_0__leaf_clk state\[1\] 0.027f
C13139 a_2787_9845# net24 1.24e-20
C13140 net52 a_4239_8573# 1.67e-19
C13141 _104_ a_10219_2045# 1.87e-19
C13142 a_4775_6031# _096_ 4.24e-19
C13143 cal_count\[0\] a_14983_9269# 0.00352f
C13144 a_816_4765# a_1007_4777# 4.61e-19
C13145 _074_ a_1045_9545# 0.00223f
C13146 _058_ a_10543_2455# 1.34e-20
C13147 _042_ a_2953_9845# 0.00809f
C13148 _053_ a_7891_3617# 1.27e-19
C13149 calibrate a_911_4777# 0.00737f
C13150 _090_ a_6519_4631# 1.33e-20
C13151 a_2033_3317# VPWR 0.613f
C13152 a_10005_6031# _064_ 7e-19
C13153 net4 a_9503_4399# 0.00976f
C13154 clknet_0_clk _089_ 2.95e-21
C13155 a_10239_9295# a_10593_9295# 0.0685f
C13156 _049_ a_5445_4399# 2.17e-20
C13157 a_12612_8725# a_12522_8751# 9.35e-20
C13158 a_13142_7271# a_13557_7369# 3.15e-19
C13159 a_579_10933# _102_ 7.75e-20
C13160 a_12631_591# ctln[3] 0.159f
C13161 cal_itt\[0\] clk 7.41e-21
C13162 cal_itt\[0\] en_co_clk 0.426f
C13163 a_4498_4373# a_4970_4399# 0.00132f
C13164 _092_ net30 0.0074f
C13165 _065_ clknet_2_0__leaf_clk 0.113f
C13166 a_13091_4943# a_13459_3317# 5.12e-19
C13167 trim_val\[4\] a_11045_3631# 2.41e-20
C13168 _074_ a_1095_11305# 0.0147f
C13169 a_10975_6031# a_11023_5108# 2.11e-19
C13170 _112_ VPWR 0.709f
C13171 _101_ a_395_9845# 5.73e-22
C13172 net27 a_4167_11471# 0.0334f
C13173 mask\[4\] a_8839_9661# 4.61e-20
C13174 _078_ a_1375_9129# 9.62e-19
C13175 a_14347_9480# net2 5.01e-19
C13176 a_1549_6794# VPWR 0.257f
C13177 a_7758_4759# VPWR 4.83e-20
C13178 _122_ a_12430_7663# 7.19e-20
C13179 net4 a_9369_3855# 0.00201f
C13180 net44 a_7569_7637# 0.0065f
C13181 _063_ a_10137_4943# 3.44e-19
C13182 net23 clknet_2_0__leaf_clk 7.41e-19
C13183 a_11352_9661# VPWR 0.00336f
C13184 _067_ _062_ 0.302f
C13185 _020_ VPWR 0.452f
C13186 trim_mask\[4\] _025_ 0.016f
C13187 net2 net51 0.0602f
C13188 net13 state\[1\] 0.144f
C13189 _134_ a_13825_6031# 0.0353f
C13190 a_1313_11989# VPWR 0.212f
C13191 _067_ a_10138_5807# 0.00191f
C13192 trim_mask\[4\] _026_ 1.16e-19
C13193 a_10329_1921# a_10785_1679# 4.2e-19
C13194 net24 a_2092_8457# 1.86e-19
C13195 a_1844_9129# mask\[1\] 1.15e-19
C13196 _040_ clknet_0_clk 0.0218f
C13197 net43 a_1357_12381# 0.00316f
C13198 a_1313_11989# a_1769_12393# 4.2e-19
C13199 net53 a_6090_10159# 4.92e-21
C13200 a_13091_4943# _109_ 4.37e-19
C13201 net44 a_7079_10217# 5.93e-19
C13202 net41 a_2309_2229# 6.96e-21
C13203 _006_ mask\[1\] 3.35e-19
C13204 a_579_10933# _022_ 6.41e-22
C13205 net12 a_4512_11305# 7.56e-21
C13206 clknet_2_2__leaf_clk trim_mask\[3\] 0.0111f
C13207 net45 net3 0.264f
C13208 net43 a_4959_9295# 2.97e-20
C13209 net13 _065_ 0.058f
C13210 net21 net27 0.448f
C13211 a_2491_3311# VPWR 0.142f
C13212 VPWR ctlp[3] 0.283f
C13213 _053_ a_10005_6031# 8.17e-19
C13214 a_7939_10383# a_8360_10383# 0.0931f
C13215 cal_itt\[3\] net30 0.176f
C13216 a_13257_4943# net49 1.04e-19
C13217 clknet_2_2__leaf_clk a_10689_2543# 3.54e-21
C13218 a_7569_7637# clk 3.45e-19
C13219 _040_ a_6198_8207# 3.98e-20
C13220 net4 a_9747_2527# 4.47e-19
C13221 a_15023_5487# trim_val\[0\] 6.59e-20
C13222 _076_ a_6515_8534# 0.00551f
C13223 _078_ a_4995_7119# 5.71e-21
C13224 _086_ a_395_9845# 3.93e-22
C13225 _124_ _041_ 0.112f
C13226 net13 a_5054_4399# 0.00141f
C13227 net2 _003_ 4.96e-20
C13228 _122_ a_10990_7485# 0.00631f
C13229 net4 _097_ 0.00243f
C13230 a_2019_9055# _081_ 0.00119f
C13231 net44 _075_ 0.0155f
C13232 _070_ cal_itt\[2\] 0.166f
C13233 net55 a_4709_2773# 1.7e-20
C13234 a_6523_7119# a_6631_7485# 0.0572f
C13235 a_10383_7093# a_10903_7261# 0.0436f
C13236 a_10586_7371# a_10864_7387# 0.125f
C13237 a_9719_1473# a_9805_1473# 0.00658f
C13238 net53 a_7201_9813# 0.00351f
C13239 clknet_2_1__leaf_clk a_5691_7637# 0.011f
C13240 _053_ _087_ 3.09e-20
C13241 net8 a_13512_1501# 0.00107f
C13242 a_4091_5309# a_4266_4943# 0.00228f
C13243 _129_ _133_ 0.108f
C13244 a_11509_3317# a_12077_3285# 0.171f
C13245 net44 a_7723_10143# 0.284f
C13246 _048_ _110_ 0.017f
C13247 a_13625_3317# a_14604_3017# 3.32e-19
C13248 net19 a_8551_10383# 8.84e-19
C13249 cal_count\[0\] a_11008_9295# 2.06e-20
C13250 a_8731_9295# _068_ 0.0027f
C13251 net30 a_9317_3285# 2.25e-21
C13252 cal_itt\[0\] a_8091_7967# 1.59e-20
C13253 clknet_2_0__leaf_clk _016_ 0.0814f
C13254 _104_ a_7021_4105# 0.021f
C13255 clknet_0_clk _048_ 0.0719f
C13256 a_14099_3017# a_14686_3017# 8.01e-20
C13257 a_6375_12021# ctlp[6] 6.16e-19
C13258 _110_ a_10219_2045# 7.89e-21
C13259 net42 _105_ 0.00141f
C13260 net10 VPWR 0.359f
C13261 _134_ a_14199_7369# 4.26e-21
C13262 clknet_2_2__leaf_clk a_13415_2442# 3.4e-20
C13263 _034_ a_3748_6281# 1.49e-19
C13264 trim_mask\[0\] clk 0.00535f
C13265 en_co_clk trim_mask\[0\] 4.6e-20
C13266 net43 mask\[5\] 2.36e-21
C13267 a_1638_4399# valid 2.99e-20
C13268 net27 _020_ 2.32e-20
C13269 _075_ en_co_clk 0.17f
C13270 _121_ _095_ 7.97e-19
C13271 trim_mask\[0\] a_9084_4515# 9.75e-19
C13272 a_3615_8207# a_3781_8207# 0.85f
C13273 clknet_2_0__leaf_clk a_4696_8207# 1.96e-19
C13274 a_448_7637# a_845_7663# 5.98e-20
C13275 net42 a_7010_3311# 5.04e-19
C13276 _119_ a_9572_2601# 7.31e-20
C13277 trim_val\[3\] a_10195_1354# 4.8e-19
C13278 _051_ trim_mask\[4\] 0.266f
C13279 a_6197_4399# VPWR 0.00584f
C13280 a_1313_11989# net27 3.66e-19
C13281 _042_ mask\[3\] 0.768f
C13282 _129_ a_14236_8457# 0.00941f
C13283 a_2143_7663# VPWR 0.213f
C13284 _092_ state\[2\] 2.44e-20
C13285 net44 a_4030_7485# 1.27e-20
C13286 clknet_2_3__leaf_clk a_10781_5807# 0.00176f
C13287 _113_ a_12599_3615# 0.0215f
C13288 net44 a_8717_10383# 1.74e-19
C13289 _037_ net46 1.3e-20
C13290 net47 _122_ 0.1f
C13291 net50 trim_val\[4\] 7.69e-20
C13292 net54 a_4576_3427# 0.167f
C13293 a_2309_2229# a_2767_2223# 0.0276f
C13294 a_11491_6031# a_11396_6031# 0.0498f
C13295 a_15259_7637# cal_count\[2\] 9.26e-21
C13296 a_12121_3677# VPWR 2.71e-19
C13297 clknet_2_1__leaf_clk a_6633_9845# 0.00421f
C13298 a_7001_7669# a_7916_8041# 0.119f
C13299 cal_itt\[0\] a_10688_9295# 3.8e-19
C13300 a_1867_3317# a_3123_3615# 0.0436f
C13301 _072_ a_8301_8207# 0.00672f
C13302 a_2033_3317# a_2383_3689# 0.23f
C13303 net47 _063_ 0.0107f
C13304 mask\[1\] _017_ 0.00371f
C13305 en_co_clk a_13933_6281# 5.5e-20
C13306 a_13557_8457# VPWR 0.00253f
C13307 a_11583_4777# VPWR 0.22f
C13308 _078_ a_1203_10927# 9.07e-20
C13309 net13 a_4696_8207# 0.014f
C13310 a_13562_8751# net2 3.98e-20
C13311 net34 a_15289_7119# 1.59e-19
C13312 cal_count\[0\] a_12344_8041# 7.26e-21
C13313 _068_ a_8301_8207# 2.69e-19
C13314 _085_ a_579_12021# 1.58e-21
C13315 _089_ net41 4.47e-19
C13316 a_11141_6031# cal_count\[3\] 0.547f
C13317 _032_ trim_val\[3\] 2.72e-19
C13318 a_11709_6273# a_12056_6031# 0.0512f
C13319 net46 a_12231_6005# 0.293f
C13320 net53 mask\[2\] 0.0021f
C13321 net23 a_561_7119# 4.14e-19
C13322 _096_ a_3933_2767# 4.21e-21
C13323 clknet_2_1__leaf_clk a_1129_9813# 0.0198f
C13324 _110_ trim[1] 5.23e-20
C13325 a_8025_8041# VPWR 9.49e-21
C13326 a_3748_6281# a_3830_6281# 0.00477f
C13327 net46 a_13880_3677# 0.0181f
C13328 net52 a_1467_7923# 6.06e-19
C13329 net9 net8 0.00149f
C13330 net30 a_9003_3829# 0.00106f
C13331 a_816_4765# net41 5.39e-20
C13332 _106_ a_9099_3689# 7.17e-19
C13333 _108_ _055_ 0.00609f
C13334 net45 a_1476_7119# 0.012f
C13335 state\[2\] a_6906_2355# 6.44e-20
C13336 _063_ a_8820_6005# 0.0782f
C13337 a_7689_2589# a_7942_2223# 4.61e-19
C13338 a_6090_10159# a_6007_9839# 2.42e-19
C13339 a_1461_10357# a_1764_10383# 0.00138f
C13340 net3 a_4905_3855# 8.21e-21
C13341 net45 mask\[0\] 0.203f
C13342 net45 valid 3.94e-19
C13343 _080_ a_1129_7361# 4.22e-19
C13344 _020_ a_8455_10383# 2.71e-19
C13345 net12 a_5829_9839# 4.53e-19
C13346 clknet_2_1__leaf_clk a_6445_10383# 0.00105f
C13347 calibrate _103_ 0.00146f
C13348 net46 a_13697_4373# 0.00127f
C13349 a_1007_6031# VPWR 4.04e-19
C13350 clknet_2_2__leaf_clk net11 3.85e-20
C13351 net50 a_9805_1473# 1.8e-20
C13352 clknet_2_0__leaf_clk _013_ 0.0347f
C13353 _125_ a_14467_8751# 0.00884f
C13354 a_1644_12533# ctlp[0] 6.9e-19
C13355 _078_ a_3431_10933# 0.0104f
C13356 net43 _039_ 0.0278f
C13357 a_2948_3689# a_3057_3689# 0.00742f
C13358 a_3123_3615# a_3302_3677# 0.0074f
C13359 a_2383_3689# a_2491_3311# 0.0572f
C13360 trim_mask\[4\] a_10781_3311# 0.0018f
C13361 a_6541_12021# a_7618_12015# 1.46e-19
C13362 _078_ a_929_8757# 0.0278f
C13363 a_4308_4917# _093_ 1.76e-20
C13364 mask\[7\] a_1461_10357# 0.0581f
C13365 net14 _005_ 8.37e-20
C13366 net51 a_4677_7882# 3.52e-20
C13367 en_co_clk a_8949_6281# 0.0454f
C13368 _077_ VPWR 0.279f
C13369 a_7824_11305# clknet_2_3__leaf_clk 2.62e-19
C13370 net15 net25 4.23e-21
C13371 a_4043_10143# a_4443_9295# 1.92e-19
C13372 net30 a_561_4405# 1.98e-21
C13373 net16 a_14071_3689# 0.0015f
C13374 _014_ a_3123_3615# 3.34e-20
C13375 a_2787_10927# a_3133_11247# 0.0134f
C13376 _095_ a_3273_4943# 0.152f
C13377 net55 _090_ 0.339f
C13378 a_2857_5461# net3 0.0132f
C13379 a_2971_8457# a_3317_8207# 0.0134f
C13380 net19 a_9871_10383# 8.67e-19
C13381 a_4043_11305# _042_ 1.01e-19
C13382 a_8657_2229# a_8912_2589# 0.0612f
C13383 _075_ _059_ 2.71e-19
C13384 _092_ _100_ 9.61e-20
C13385 net14 net15 6.76e-20
C13386 clknet_2_1__leaf_clk a_3411_9839# 0.0045f
C13387 a_1276_565# VPWR 0.267f
C13388 net15 a_3399_7119# 7.77e-19
C13389 a_5699_9269# _077_ 4.15e-20
C13390 a_5067_9661# a_4871_8181# 2.66e-20
C13391 a_5524_9295# a_5535_8181# 1.04e-19
C13392 a_4471_4007# a_4576_3427# 8.18e-19
C13393 net16 a_13279_8207# 0.00111f
C13394 _033_ a_9099_3689# 4.76e-19
C13395 net16 _058_ 0.0446f
C13396 a_8583_3317# a_9839_3615# 0.0436f
C13397 a_14422_7093# _134_ 4.24e-20
C13398 net12 a_7442_7119# 1.18e-19
C13399 _005_ a_395_7119# 0.213f
C13400 net45 _079_ 0.004f
C13401 a_1019_7485# VPWR 0.144f
C13402 cal_count\[3\] net42 9.22e-20
C13403 _106_ _088_ 3.91e-20
C13404 _048_ net41 2.36e-19
C13405 a_5691_7637# a_6007_7119# 0.0041f
C13406 a_12916_8751# VPWR 0.00405f
C13407 _078_ a_6198_8534# 4.08e-19
C13408 a_10975_6031# VPWR 0.456f
C13409 a_5087_3855# a_6737_3855# 3.22e-20
C13410 net22 _049_ 2.83e-19
C13411 a_11343_3317# a_13880_3677# 1.96e-21
C13412 a_7939_10383# _000_ 4.43e-20
C13413 _034_ a_4308_4917# 3.76e-21
C13414 a_8105_10383# a_8215_9295# 4.37e-21
C13415 a_10405_9295# a_10688_9295# 0.196f
C13416 a_14236_8457# a_14318_8457# 0.00477f
C13417 net2 _131_ 0.157f
C13418 a_3431_10933# a_3597_10933# 0.852f
C13419 trim_mask\[1\] a_14099_1929# 1.52e-20
C13420 a_2877_2197# clk 0.00393f
C13421 calibrate a_7140_2223# 2.39e-20
C13422 a_9225_2197# a_9572_2601# 0.0512f
C13423 net18 a_10864_9269# 0.0113f
C13424 net30 a_8485_4943# 1.49e-19
C13425 a_14099_3017# a_13257_1141# 2.19e-21
C13426 net44 _042_ 0.0115f
C13427 _106_ trim_val\[4\] 0.0101f
C13428 net44 a_7723_6807# 1.65e-19
C13429 a_763_8757# net24 0.0466f
C13430 _065_ a_4167_6575# 0.0287f
C13431 a_7527_4631# _028_ 6.9e-20
C13432 _058_ a_10699_3311# 3.18e-19
C13433 mask\[1\] a_3868_7119# 2.41e-19
C13434 _108_ trim_val\[2\] 0.0396f
C13435 net33 a_15023_2223# 0.251f
C13436 a_13783_6183# a_13715_5309# 5.55e-20
C13437 net33 _134_ 3.12e-20
C13438 a_395_6031# result[0] 0.0108f
C13439 net52 a_2787_7119# 5.23e-20
C13440 _096_ a_1651_4703# 8.71e-21
C13441 net44 a_7210_5807# 1.14e-20
C13442 state\[2\] a_6737_4719# 0.00228f
C13443 a_1476_7119# a_2953_7119# 9.39e-20
C13444 net45 net54 0.00148f
C13445 mask\[0\] a_2953_7119# 0.0252f
C13446 a_1173_10205# VPWR 4.15e-19
C13447 a_3057_4719# _097_ 0.0499f
C13448 a_8583_3317# a_9207_3311# 9.73e-19
C13449 a_1644_12533# a_579_12021# 0.0106f
C13450 _110_ _112_ 0.251f
C13451 net9 a_12924_8029# 3.98e-19
C13452 a_8298_2767# clk 0.00318f
C13453 net46 a_13825_5185# 0.181f
C13454 clknet_2_3__leaf_clk a_10239_9295# 0.781f
C13455 _024_ a_11691_4399# 0.00219f
C13456 a_11067_4405# _109_ 2.68e-21
C13457 VPWR ctlp[1] 0.348f
C13458 a_5915_11721# _101_ 1.76e-20
C13459 cal_itt\[1\] _091_ 0.00111f
C13460 net26 net24 6.35e-21
C13461 mask\[7\] a_745_10933# 0.0143f
C13462 a_4512_11305# a_5997_10927# 7.36e-20
C13463 _064_ a_9503_4399# 3.08e-19
C13464 a_9084_4515# a_8298_2767# 1.71e-19
C13465 a_7723_6807# clk 0.0113f
C13466 net44 a_7521_11293# 0.00374f
C13467 _074_ a_1211_7983# 4.22e-19
C13468 net43 a_2857_7637# 0.00886f
C13469 _078_ clknet_2_0__leaf_clk 0.006f
C13470 a_5536_4399# state\[2\] 7.14e-20
C13471 _050_ a_8583_3317# 2.14e-19
C13472 state\[2\] a_5067_2045# 9.5e-19
C13473 net15 a_4222_7119# 6.83e-20
C13474 a_1000_12381# ctlp[0] 5.04e-19
C13475 a_3781_8207# a_4227_8207# 2.28e-19
C13476 a_4349_8449# a_4858_8573# 2.6e-19
C13477 net52 a_3208_10205# 6.06e-21
C13478 a_7210_5807# clk 0.00194f
C13479 net31 _131_ 0.0059f
C13480 cal_count\[2\] a_14485_7663# 5.95e-20
C13481 net15 a_2659_2601# 0.00815f
C13482 _129_ a_14318_8457# 3.83e-19
C13483 a_15023_5487# net32 0.00105f
C13484 trim_val\[4\] _033_ 5.22e-21
C13485 a_579_12021# a_2828_12131# 2.64e-21
C13486 _072_ a_7088_7119# 4.11e-19
C13487 a_455_12533# ctlp[0] 0.0347f
C13488 mask\[4\] a_7939_10383# 0.00766f
C13489 _128_ a_13356_8457# 0.00566f
C13490 _101_ a_5515_6005# 4.33e-21
C13491 a_4687_12319# _078_ 3.27e-20
C13492 _053_ a_10864_7387# 0.00902f
C13493 _092_ _118_ 9.2e-20
C13494 a_6173_7119# VPWR 0.602f
C13495 a_10747_8970# _124_ 0.242f
C13496 _090_ _093_ 0.0849f
C13497 clknet_2_3__leaf_clk a_13441_6281# 2.43e-21
C13498 clknet_2_1__leaf_clk net47 6.21e-20
C13499 cal_itt\[0\] a_9460_6807# 0.379f
C13500 _068_ a_7088_7119# 9.75e-21
C13501 _072_ _063_ 0.00253f
C13502 _052_ a_8583_3317# 3.51e-20
C13503 _093_ a_3847_4438# 7.79e-20
C13504 _127_ a_14377_7983# 7.44e-21
C13505 net16 a_13607_4943# 0.00336f
C13506 a_13512_4943# a_13519_4007# 4.39e-20
C13507 net14 net25 0.00744f
C13508 net4 a_4709_2773# 0.0196f
C13509 mask\[3\] a_4959_9295# 0.0512f
C13510 a_4775_6031# _092_ 3.51e-19
C13511 _075_ a_5694_6031# 6.2e-19
C13512 net45 a_2645_3677# 0.00215f
C13513 _068_ _063_ 0.647f
C13514 _065_ _037_ 1.04e-20
C13515 a_13415_2442# a_14335_2442# 1.32e-20
C13516 _078_ net13 0.0381f
C13517 mask\[0\] a_2857_5461# 0.00815f
C13518 _115_ a_14099_1929# 5.06e-19
C13519 net43 a_8270_8029# 0.00288f
C13520 _106_ a_8745_4943# 5.46e-19
C13521 net44 a_6909_10933# 0.0485f
C13522 _122_ net46 1.07e-20
C13523 a_3116_12533# a_2787_10927# 7.82e-21
C13524 a_15159_9269# net40 1.87e-20
C13525 _126_ a_15023_8751# 0.0463f
C13526 _125_ a_14249_8725# 0.206f
C13527 _090_ a_2865_4460# 1.71e-19
C13528 net12 a_6619_7119# 0.00108f
C13529 clknet_2_1__leaf_clk a_7355_11305# 3.14e-19
C13530 _064_ a_9747_2527# 1.96e-19
C13531 net19 a_8767_11471# 0.118f
C13532 _110_ net10 1.95e-20
C13533 _099_ a_3530_4438# 2.1e-19
C13534 trim_mask\[0\] a_9802_4007# 0.028f
C13535 _123_ a_12824_7663# 0.00237f
C13536 _063_ net46 1.01e-21
C13537 net43 a_2953_9845# 0.0461f
C13538 a_3333_2601# VPWR 2.84e-20
C13539 _076_ a_6515_6794# 7.8e-20
C13540 cal_count\[0\] a_14236_8457# 4.41e-19
C13541 a_15023_5487# VPWR 0.494f
C13542 net19 _048_ 0.0218f
C13543 a_395_4405# a_455_3571# 3.29e-20
C13544 cal_itt\[0\] _107_ 3.22e-19
C13545 _049_ a_4871_6031# 7.11e-19
C13546 net14 a_395_7119# 0.00787f
C13547 a_4165_11989# a_3947_11305# 3.29e-20
C13548 a_3947_12393# a_4165_10901# 4.07e-20
C13549 trim_mask\[0\] _108_ 0.295f
C13550 a_5177_1921# clk 0.0185f
C13551 net9 a_13008_7663# 1.65e-19
C13552 _088_ _054_ 0.0123f
C13553 clknet_2_3__leaf_clk _066_ 0.29f
C13554 _134_ _136_ 0.00622f
C13555 a_10543_2455# a_10329_1921# 2.67e-19
C13556 _070_ a_10043_7983# 3.51e-21
C13557 mask\[5\] mask\[3\] 7.12e-22
C13558 cal_itt\[2\] _106_ 1.12e-20
C13559 _012_ cal 0.00363f
C13560 net48 a_13257_1141# 6.36e-19
C13561 _050_ a_7190_3855# 0.0186f
C13562 net47 a_13111_6031# 1.31e-20
C13563 a_7262_5461# _054_ 3.69e-21
C13564 a_579_12021# a_1000_12381# 0.0931f
C13565 a_5536_4399# _100_ 2.66e-19
C13566 _065_ a_8301_8207# 2.28e-19
C13567 _007_ result[3] 0.00262f
C13568 a_1129_9813# result[4] 2.56e-19
C13569 _042_ a_4801_9839# 3.94e-19
C13570 net23 a_1467_7923# 0.0294f
C13571 cal_itt\[2\] net2 0.0512f
C13572 _118_ a_9317_3285# 3.01e-19
C13573 net13 a_3597_10933# 0.00405f
C13574 a_1638_7485# _039_ 1.6e-20
C13575 _079_ a_2857_5461# 8.04e-21
C13576 net18 a_11023_5108# 0.0112f
C13577 net54 a_4905_3855# 1.14e-19
C13578 a_455_12533# a_579_12021# 0.0132f
C13579 _086_ a_911_10217# 2.06e-21
C13580 net12 _062_ 0.00931f
C13581 net5 comp 6.19e-20
C13582 _101_ mask\[2\] 0.269f
C13583 _094_ state\[1\] 3.09e-22
C13584 a_3852_11293# VPWR 0.0857f
C13585 net43 a_1638_7485# 2.06e-19
C13586 a_13091_4943# _112_ 6.36e-19
C13587 a_11583_4777# _110_ 1.92e-20
C13588 _052_ a_7190_3855# 0.00659f
C13589 net37 _109_ 7.01e-21
C13590 net42 a_6566_5193# 2.29e-19
C13591 a_5515_6005# _060_ 3.9e-20
C13592 net30 _105_ 0.0135f
C13593 _013_ a_2948_3689# 4.03e-21
C13594 net22 sample 2.63e-19
C13595 net41 a_2033_3317# 0.0258f
C13596 net6 clk 0.00704f
C13597 clknet_2_3__leaf_clk a_11545_9049# 0.0797f
C13598 _098_ a_7190_3855# 1.2e-21
C13599 cal_itt\[0\] a_8495_6895# 1.53e-19
C13600 _065_ _094_ 0.191f
C13601 _058_ a_11955_3689# 5.31e-19
C13602 _062_ a_5340_6031# 9.67e-20
C13603 a_13091_1141# a_13257_1141# 0.902f
C13604 net4 _070_ 0.138f
C13605 net14 a_2659_2601# 1.93e-19
C13606 net9 a_13459_3317# 2.54e-21
C13607 _095_ a_4091_5309# 0.0496f
C13608 cal_count\[0\] _129_ 0.0507f
C13609 a_6822_4105# a_6737_3855# 8.13e-19
C13610 a_10688_9295# a_11008_9295# 0.00184f
C13611 a_3830_6281# _090_ 2.4e-20
C13612 _078_ a_561_7119# 0.00934f
C13613 a_10864_9269# a_11268_9295# 3.94e-19
C13614 net47 a_11814_9295# 0.0549f
C13615 net13 a_5502_6397# 6.96e-20
C13616 net4 trim_mask\[2\] 9.27e-20
C13617 a_11583_4777# a_12148_4777# 7.99e-20
C13618 a_10975_4105# a_11057_3855# 0.00393f
C13619 net16 _113_ 0.00136f
C13620 net18 a_11268_9295# 4e-19
C13621 net47 a_11622_7485# 1.1e-20
C13622 a_3947_11305# VPWR 0.202f
C13623 clknet_2_2__leaf_clk _028_ 0.00261f
C13624 net43 a_1585_10217# 0.00157f
C13625 net12 a_6198_8534# 6.82e-19
C13626 _101_ a_6428_7119# 8.21e-21
C13627 net45 a_1125_7663# 0.00109f
C13628 a_7109_11989# VPWR 0.203f
C13629 a_395_4405# _099_ 1.82e-20
C13630 clknet_2_0__leaf_clk _004_ 0.107f
C13631 _073_ net30 0.348f
C13632 _108_ a_13869_4943# 6.71e-19
C13633 net33 a_15054_5193# 3.83e-19
C13634 _010_ mask\[7\] 0.00329f
C13635 a_1467_7923# _016_ 2.63e-19
C13636 net53 a_4609_9295# 2.02e-19
C13637 net33 trim_val\[1\] 0.127f
C13638 a_1651_10143# a_929_8757# 5.38e-20
C13639 _017_ a_3615_8207# 0.383f
C13640 trim_mask\[0\] _107_ 0.0667f
C13641 net4 _090_ 3.3e-20
C13642 _119_ a_8491_2229# 8.06e-19
C13643 net44 a_4959_9295# 0.159f
C13644 _012_ a_561_4405# 0.263f
C13645 a_395_4405# a_1129_4373# 0.0701f
C13646 a_12992_8751# a_13016_9117# 0.0016f
C13647 _041_ a_12546_9129# 0.0018f
C13648 a_745_12021# ctlp[0] 0.00268f
C13649 a_8389_5193# a_8473_5193# 0.0927f
C13650 _075_ _107_ 5.06e-19
C13651 _065_ a_2787_7119# 2.03e-19
C13652 net5 a_13111_6031# 7.07e-21
C13653 _118_ a_9003_3829# 0.052f
C13654 _064_ a_10676_1679# 0.00192f
C13655 net12 a_5524_1679# 0.00278f
C13656 a_4425_6031# _050_ 1.33e-19
C13657 net55 _106_ 0.00408f
C13658 a_4871_8181# net45 4.09e-19
C13659 a_12344_8041# cal_count\[2\] 2.99e-20
C13660 a_13050_7637# a_13164_8029# 1.84e-19
C13661 a_12900_7663# a_13092_8029# 0.00536f
C13662 net43 mask\[3\] 0.0301f
C13663 net15 _019_ -1.01e-36
C13664 a_5037_6031# VPWR 1.5e-19
C13665 _076_ net45 1.28e-20
C13666 a_4471_4007# a_4905_3855# 0.00393f
C13667 net23 a_2787_7119# 6.85e-20
C13668 net43 a_6741_7361# 1.24e-20
C13669 _049_ trim_mask\[0\] 0.00997f
C13670 _077_ a_6198_8207# 2.88e-19
C13671 net19 a_7810_12381# 9.63e-20
C13672 net4 a_9719_1473# 7.64e-22
C13673 en_co_clk a_9529_6059# 1.15e-19
C13674 clknet_2_1__leaf_clk _072_ 1.55e-20
C13675 a_7800_4631# VPWR 0.165f
C13676 net34 a_15023_2223# 0.0216f
C13677 _049_ _075_ 0.178f
C13678 net34 _134_ 1.5e-20
C13679 net30 a_3148_4399# 3.79e-19
C13680 net12 clknet_2_0__leaf_clk 1.37e-19
C13681 _036_ net2 0.152f
C13682 a_10851_1653# a_10676_1679# 0.234f
C13683 trim_mask\[1\] a_13183_3311# 0.118f
C13684 net6 ctln[0] 0.0657f
C13685 a_13257_1141# a_14281_1513# 2.36e-20
C13686 a_13825_1109# a_13869_1501# 3.69e-19
C13687 a_4266_4943# state\[0\] 3.57e-20
C13688 a_5455_4943# a_5931_4105# 1.02e-19
C13689 mask\[1\] _080_ 0.0845f
C13690 net9 a_12169_2197# 0.00805f
C13691 a_7259_11305# a_7723_10143# 0.00122f
C13692 net26 a_6181_10383# 0.00123f
C13693 a_14347_1439# trim[3] 2.13e-19
C13694 net13 ctln[7] 0.101f
C13695 calibrate a_937_4105# 0.0387f
C13696 net44 mask\[5\] 0.0328f
C13697 a_2309_2229# a_3224_2601# 0.119f
C13698 a_14972_5193# trim[4] 0.00111f
C13699 clknet_2_1__leaf_clk a_4443_9295# 0.243f
C13700 a_11067_3017# a_11435_2229# 0.0111f
C13701 a_1000_11293# _102_ 3.52e-20
C13702 net47 _092_ 0.0024f
C13703 _108_ _030_ 1.99e-20
C13704 net55 a_3667_3829# 8.54e-19
C13705 _067_ a_9621_8029# 0.00258f
C13706 net12 net11 0.00123f
C13707 _005_ VPWR 0.428f
C13708 clknet_2_2__leaf_clk a_13880_3677# 1.96e-20
C13709 clknet_2_0__leaf_clk a_5340_6031# 7.25e-20
C13710 clknet_2_3__leaf_clk a_9471_9269# 0.0739f
C13711 a_3868_7119# _050_ 3.91e-20
C13712 net27 a_3947_11305# 1.05e-19
C13713 a_10975_6031# a_10699_5487# 4.17e-19
C13714 net44 a_6999_12015# 0.0135f
C13715 a_7109_11989# net27 3.47e-19
C13716 clknet_2_1__leaf_clk net52 0.743f
C13717 _101_ a_4674_10927# 1.05e-20
C13718 net4 a_9595_1679# 2.87e-19
C13719 _123_ a_12061_7669# 0.0182f
C13720 net13 net12 0.0452f
C13721 clknet_2_2__leaf_clk a_13697_4373# 0.00101f
C13722 net15 VPWR 2.08f
C13723 a_9802_4007# a_8298_2767# 8.19e-20
C13724 state\[2\] a_7010_3311# 0.00652f
C13725 net21 a_4512_11305# 0.00558f
C13726 _016_ a_2787_7119# 0.156f
C13727 a_4030_7485# _049_ 3.27e-20
C13728 a_8820_6005# _092_ 0.0621f
C13729 net9 a_12520_7637# 0.00712f
C13730 _065_ _122_ 0.0791f
C13731 a_579_12021# a_745_12021# 0.883f
C13732 trim_mask\[1\] net49 0.17f
C13733 a_14193_3285# a_14702_3311# 2.6e-19
C13734 calibrate net42 3.11e-19
C13735 cal_count\[3\] net30 0.00416f
C13736 a_2787_9845# a_2961_9545# 3.77e-20
C13737 _108_ a_8298_2767# 7.12e-19
C13738 a_7379_2197# a_7942_2223# 0.0498f
C13739 a_7310_2223# a_7689_2589# 3.16e-19
C13740 a_7184_2339# a_7140_2223# 1.46e-19
C13741 a_7223_2465# a_8912_2589# 3.88e-21
C13742 _074_ net24 0.05f
C13743 a_7351_8041# VPWR 0.214f
C13744 a_8949_6281# _107_ 4.95e-20
C13745 net46 a_9761_1679# 0.051f
C13746 a_13919_8751# _129_ 0.00317f
C13747 net13 a_5340_6031# 0.00163f
C13748 _085_ _022_ 0.00128f
C13749 a_10903_7261# a_10781_5487# 4.56e-21
C13750 net37 _125_ 0.00738f
C13751 net47 a_12992_8751# 0.216f
C13752 a_14347_9480# trimb[1] 6.6e-19
C13753 _065_ _063_ 4.66e-19
C13754 clknet_2_3__leaf_clk a_12056_6031# 0.0465f
C13755 net19 _020_ 0.0017f
C13756 a_9503_4399# a_9664_3689# 1.59e-20
C13757 _074_ _084_ 0.0777f
C13758 net52 a_2368_9955# 0.00178f
C13759 a_4091_5309# calibrate 4.35e-21
C13760 a_7891_3617# a_8583_3317# 4.62e-21
C13761 a_3597_12021# a_2910_12131# 9.72e-20
C13762 a_3947_12393# a_4043_12393# 0.0138f
C13763 mask\[3\] a_2857_7637# 8.09e-21
C13764 mask\[1\] a_6885_8372# 2.18e-20
C13765 a_855_4105# a_995_3530# 3.78e-19
C13766 net43 a_4043_11305# 0.00118f
C13767 a_3781_8207# a_4043_7093# 8.37e-21
C13768 _060_ a_4815_3031# 5.66e-19
C13769 a_6541_12021# a_6891_12393# 0.23f
C13770 clknet_0_clk a_6173_7119# 8.12e-20
C13771 a_4030_9839# VPWR 7.5e-19
C13772 a_4883_6397# net55 4.2e-19
C13773 _096_ state\[1\] 2.16e-19
C13774 a_561_7119# _004_ 1.44e-20
C13775 _119_ _032_ 2.87e-21
C13776 a_1279_9129# net24 0.0302f
C13777 a_2019_9055# a_1844_9129# 0.234f
C13778 a_8298_2767# a_9115_2223# 2.2e-19
C13779 _050_ _103_ 0.0737f
C13780 _069_ a_9677_8457# 0.0097f
C13781 a_911_6031# result[0] 0.00117f
C13782 clknet_2_3__leaf_clk _058_ 6.52e-19
C13783 _006_ a_2019_9055# 4.1e-20
C13784 a_13164_8029# VPWR 5.16e-19
C13785 net46 a_13111_6031# 6.86e-20
C13786 a_6467_9845# a_7548_10217# 0.102f
C13787 _008_ a_7723_10143# 3.61e-20
C13788 a_8491_2229# a_9225_2197# 0.0535f
C13789 _027_ a_8657_2229# 0.74f
C13790 a_11141_6031# _135_ 0.00145f
C13791 a_13881_2741# a_13607_1513# 1.89e-20
C13792 a_745_10933# a_1677_9545# 7.22e-21
C13793 net31 a_13693_3883# 2.11e-20
C13794 _024_ _025_ 6.82e-20
C13795 net46 a_10787_1135# 6.39e-20
C13796 _065_ _096_ 2.11e-19
C13797 net53 a_6181_10633# 0.0573f
C13798 net14 a_1493_11721# 5.51e-19
C13799 net43 a_9459_7895# 7.84e-20
C13800 net43 a_4687_11231# 0.273f
C13801 mask\[1\] a_1651_7093# 0.00118f
C13802 net46 trim[3] 1.66e-19
C13803 a_10864_9269# VPWR 0.242f
C13804 a_8298_5487# net42 0.00341f
C13805 net55 _054_ 4.54e-20
C13806 _103_ _052_ 9.12e-20
C13807 a_2092_8457# mask\[0\] 0.00105f
C13808 a_8307_4943# _107_ 0.00775f
C13809 net43 net44 0.0814f
C13810 a_7548_10217# VPWR 0.285f
C13811 a_1313_10901# a_1095_11305# 0.21f
C13812 a_745_10933# a_1835_11231# 0.0424f
C13813 a_15023_8751# VPWR 0.499f
C13814 trim_val\[0\] net32 1.68e-19
C13815 clknet_2_0__leaf_clk result[2] 0.00281f
C13816 net18 VPWR 1.45f
C13817 _078_ a_1585_4777# 6.12e-20
C13818 a_2601_3285# clk 2.77e-19
C13819 a_10820_7485# VPWR 7.67e-19
C13820 _093_ a_3667_3829# 0.0694f
C13821 a_9664_3689# a_9747_2527# 1.45e-19
C13822 _078_ a_5915_10927# 0.00401f
C13823 a_9839_3615# a_9572_2601# 8.54e-21
C13824 a_9004_3677# a_8298_2767# 9.38e-19
C13825 net15 net27 0.008f
C13826 net29 a_448_11445# 5.41e-20
C13827 _134_ cal_count\[3\] 0.0058f
C13828 _098_ _103_ 0.0872f
C13829 trim_mask\[3\] a_12169_2197# 8.85e-19
C13830 a_3977_7119# _049_ 5.28e-20
C13831 a_12153_8757# a_13050_7637# 1.55e-19
C13832 a_12612_8725# a_12344_8041# 4.26e-20
C13833 a_12436_9129# a_12520_7637# 4.14e-22
C13834 a_1019_9839# _082_ 9.17e-19
C13835 mask\[3\] a_2953_9845# 2.82e-19
C13836 clknet_2_2__leaf_clk a_13825_5185# 2.34e-19
C13837 net16 a_13783_6183# 0.0132f
C13838 _000_ _070_ 6.75e-20
C13839 _107_ a_8298_2767# 0.00242f
C13840 a_1822_12015# VPWR 7.89e-19
C13841 _062_ _091_ 0.00153f
C13842 a_9572_2601# a_9734_2223# 0.00645f
C13843 a_11435_2229# a_11856_2589# 0.0931f
C13844 net45 a_2564_2589# 2.47e-19
C13845 _049_ a_8307_4943# 0.00201f
C13846 net29 a_1203_10927# 1.1e-19
C13847 _129_ en_co_clk 4.52e-19
C13848 net33 a_15023_10927# 0.0323f
C13849 a_12165_6031# VPWR 3.07e-20
C13850 cal_count\[0\] a_13100_8751# 1.36e-19
C13851 net25 VPWR 0.637f
C13852 net26 a_8673_10625# 3.76e-20
C13853 _074_ a_1129_6273# 0.00439f
C13854 cal_count\[2\] _133_ 0.308f
C13855 net43 clk 0.00926f
C13856 net43 en_co_clk 1.22e-20
C13857 a_7800_4631# _104_ 0.00139f
C13858 a_2198_9117# mask\[0\] 2.34e-20
C13859 _054_ a_7715_3285# 3.69e-20
C13860 net28 a_4209_12381# 0.0021f
C13861 _072_ a_6007_7119# 2.88e-19
C13862 trim_mask\[0\] trim_mask\[4\] 0.115f
C13863 net51 mask\[0\] 6.26e-20
C13864 net14 VPWR 1.38f
C13865 _060_ a_5087_3855# 0.078f
C13866 _121_ _050_ 4.53e-21
C13867 a_3399_7119# VPWR 2.37e-19
C13868 _078_ a_1467_7923# 0.053f
C13869 a_7210_5807# _107_ 0.00102f
C13870 clknet_2_0__leaf_clk a_2309_2229# 0.584f
C13871 _122_ _067_ 1.5e-19
C13872 net14 a_1769_12393# 1.84e-19
C13873 a_9129_10383# VPWR 1.75e-19
C13874 net37 trim[1] 0.0301f
C13875 trim_mask\[2\] net48 0.139f
C13876 _097_ a_3530_4438# 9.3e-19
C13877 a_4498_4373# a_4815_3031# 1.86e-20
C13878 a_13625_3317# a_14649_3689# 2.36e-20
C13879 a_14193_3285# a_14237_3677# 3.69e-19
C13880 _062_ _089_ 5.29e-21
C13881 net9 a_11599_6397# 3.15e-19
C13882 trim_mask\[1\] a_14172_1513# 9.68e-21
C13883 trim_val\[0\] VPWR 0.354f
C13884 _067_ _063_ 0.54f
C13885 a_11601_2229# _115_ 7.12e-20
C13886 a_11951_2601# a_12516_2601# 7.99e-20
C13887 a_7723_6807# _049_ 7.54e-22
C13888 a_3597_10933# a_5915_10927# 5.85e-20
C13889 _106_ a_9595_5193# 5e-19
C13890 net47 _132_ 4.97e-20
C13891 a_7259_11305# _042_ 8.95e-20
C13892 _049_ a_7210_5807# 9.24e-19
C13893 net16 a_14347_9480# 0.00571f
C13894 net52 a_6007_7119# 2.88e-20
C13895 a_395_7119# VPWR 0.509f
C13896 _072_ _092_ 4.89e-20
C13897 net34 trim_val\[1\] 0.00267f
C13898 net33 a_14377_9545# 0.00361f
C13899 net16 a_13142_7271# 1.26e-20
C13900 net30 _119_ 6.18e-19
C13901 _101_ a_4609_9295# 0.0138f
C13902 a_11575_8790# VPWR 1e-19
C13903 a_5449_6031# VPWR 1.14e-19
C13904 a_14335_4020# a_14981_4020# 3.09e-20
C13905 net45 net1 1.51e-20
C13906 a_3615_8207# _121_ 2.11e-20
C13907 net44 a_2857_7637# 0.00139f
C13908 _126_ VPWR 0.852f
C13909 _078_ a_4043_10143# 1.24e-21
C13910 a_4993_6273# net55 0.00343f
C13911 trim_mask\[2\] a_13091_1141# 0.00247f
C13912 _049_ a_4658_3427# 3.24e-20
C13913 _105_ _118_ 0.00226f
C13914 a_3431_12021# a_3431_10933# 7.57e-19
C13915 net16 a_14181_6031# 0.00162f
C13916 trim_val\[2\] _056_ 0.228f
C13917 _027_ a_10329_1921# 1.21e-19
C13918 _064_ trim_mask\[2\] 0.525f
C13919 a_7259_11305# a_7521_11293# 0.00171f
C13920 a_7477_10901# a_7933_11305# 4.2e-19
C13921 a_8731_9295# a_8993_9295# 0.00171f
C13922 a_8949_9537# cal_itt\[0\] 1.93e-19
C13923 a_9296_9295# a_9458_9661# 0.00645f
C13924 net4 _106_ 0.0182f
C13925 net13 a_5691_2741# 1.58e-19
C13926 net43 a_8091_7967# 0.285f
C13927 net30 _095_ 1.44e-19
C13928 _015_ a_4901_2773# 2.51e-20
C13929 _092_ net46 9.46e-20
C13930 a_10975_4105# a_10699_3311# 8.33e-19
C13931 _072_ cal_itt\[3\] 0.352f
C13932 _034_ a_4883_6397# 7.15e-19
C13933 clknet_2_1__leaf_clk _065_ 0.0218f
C13934 net4 net2 0.00902f
C13935 a_14981_4020# a_15023_2767# 8.1e-20
C13936 net16 a_13881_2741# 0.00875f
C13937 a_4222_7119# VPWR 1.14e-19
C13938 _048_ a_4863_4917# 0.0273f
C13939 net14 net27 0.00986f
C13940 net21 a_4209_12381# 7.65e-20
C13941 a_12153_8757# VPWR 0.294f
C13942 _068_ cal_itt\[3\] 3.49e-19
C13943 a_4091_5309# _015_ 1.97e-19
C13944 a_2659_2601# VPWR 0.205f
C13945 a_1769_11305# VPWR 1.17e-19
C13946 trim_mask\[2\] a_10851_1653# 2.02e-20
C13947 clknet_2_1__leaf_clk net23 0.00695f
C13948 clknet_2_3__leaf_clk _069_ 4.01e-20
C13949 a_7800_4631# _110_ 4.49e-21
C13950 a_12344_8041# a_12900_7663# 0.00329f
C13951 clknet_2_2__leaf_clk a_7181_2589# 2.72e-20
C13952 a_10990_7485# _136_ 0.00121f
C13953 _078_ a_2787_7119# 1.06e-21
C13954 _124_ a_10864_7387# 5.74e-22
C13955 net43 _059_ 1.7e-19
C13956 cal_count\[1\] _133_ 0.00162f
C13957 a_11023_5108# VPWR 0.242f
C13958 _129_ cal_count\[2\] 0.127f
C13959 _011_ _023_ 0.00513f
C13960 clknet_0_clk a_7800_4631# 2.5e-19
C13961 _062_ _048_ 0.118f
C13962 _050_ a_3273_4943# 0.018f
C13963 clknet_2_3__leaf_clk a_8022_7119# 5.7e-20
C13964 _085_ _046_ 0.0687f
C13965 net45 a_1830_6031# 0.00342f
C13966 a_1095_11305# result[5] 2.17e-19
C13967 _070_ _053_ 1.58e-19
C13968 net28 a_1203_10927# 7.39e-20
C13969 a_4609_1679# a_5524_1679# 0.119f
C13970 a_4443_1679# a_4864_1679# 0.0931f
C13971 a_6173_7119# a_6523_7119# 0.23f
C13972 cal_itt\[0\] a_11491_6031# 5.19e-21
C13973 net4 a_3667_3829# 3.57e-20
C13974 _117_ a_10569_1109# 0.014f
C13975 a_6909_10933# a_7259_11305# 0.23f
C13976 _042_ _008_ 6.43e-21
C13977 _064_ a_11045_3631# 1.56e-20
C13978 a_11343_3317# a_11067_3017# 1.75e-19
C13979 _132_ net5 0.00278f
C13980 net12 _028_ 0.00295f
C13981 net47 _035_ 0.144f
C13982 a_11244_9661# a_11168_9661# 0.00212f
C13983 net18 _104_ 0.0279f
C13984 clknet_2_0__leaf_clk a_1651_6005# 3.93e-19
C13985 a_10055_2767# VPWR 0.418f
C13986 a_11067_3017# a_11149_3017# 0.171f
C13987 net4 _033_ 0.0333f
C13988 _136_ a_12502_4765# 1.06e-19
C13989 _024_ a_11801_4373# 0.00253f
C13990 a_11067_4405# a_11583_4777# 0.115f
C13991 clknet_2_0__leaf_clk a_4609_1679# 0.00447f
C13992 net33 net5 3.09e-19
C13993 _012_ a_1019_4399# 1.08e-20
C13994 net43 a_1184_9117# 2.79e-19
C13995 a_9926_2589# VPWR 0.00178f
C13996 clknet_2_0__leaf_clk a_816_4765# 0.00154f
C13997 _078_ a_2689_8751# 0.129f
C13998 a_8307_6575# VPWR 0.31f
C13999 a_561_4405# a_1651_4703# 0.0424f
C14000 a_1129_4373# a_911_4777# 0.21f
C14001 _105_ a_10137_4943# 8.14e-20
C14002 cal_count\[1\] a_14236_8457# 0.145f
C14003 a_9802_4007# a_9369_4105# 7.66e-19
C14004 _053_ _090_ 2.67e-20
C14005 net15 clknet_0_clk 0.0846f
C14006 a_7460_5807# VPWR 0.00252f
C14007 net28 a_3431_10933# 9.8e-20
C14008 a_4259_6031# a_4680_6031# 0.0897f
C14009 a_11435_2229# trim_val\[3\] 8.78e-20
C14010 _057_ a_12631_591# 0.0557f
C14011 cal_count\[0\] a_13919_8751# 0.0451f
C14012 a_3053_8457# _017_ 0.00387f
C14013 _040_ clknet_2_0__leaf_clk 0.0704f
C14014 a_13307_1707# a_13393_1707# 0.00658f
C14015 a_10329_1921# _117_ 0.00241f
C14016 a_10111_1679# a_10195_1354# 6.3e-19
C14017 net46 a_9317_3285# 0.159f
C14018 a_3891_4943# a_4308_4917# 0.103f
C14019 a_11987_8757# a_13016_9117# 0.00248f
C14020 _126_ a_14807_8359# 0.0258f
C14021 net47 _136_ 0.00242f
C14022 a_855_4105# valid 0.00378f
C14023 _103_ a_8389_5193# 1.2e-19
C14024 _087_ a_5625_4943# 3.03e-20
C14025 clknet_2_1__leaf_clk _016_ 0.0775f
C14026 _108_ a_9369_4105# 0.0131f
C14027 a_3840_8867# mask\[1\] 0.00832f
C14028 trim_mask\[0\] a_12723_4943# 6.85e-19
C14029 net9 _112_ 1.19e-20
C14030 a_10864_7387# a_13356_7369# 8.14e-21
C14031 a_10903_7261# a_11369_7119# 0.00188f
C14032 a_11059_7356# a_11297_7119# 0.00171f
C14033 a_10990_7485# a_10861_7119# 4.2e-19
C14034 net16 a_13562_8751# 0.00389f
C14035 _074_ result[1] 0.00166f
C14036 _045_ clknet_2_1__leaf_clk 0.0454f
C14037 _064_ a_9595_1679# 4.61e-20
C14038 net13 a_4609_1679# 0.0212f
C14039 net46 a_11856_2589# 2.48e-19
C14040 net24 a_911_7119# 7.21e-21
C14041 net12 a_5915_10927# 0.0117f
C14042 a_6927_3311# VPWR 0.332f
C14043 a_11895_7669# a_13092_8029# 1.63e-19
C14044 net9 a_11352_9661# 1.04e-19
C14045 mask\[1\] a_2971_8457# 0.06f
C14046 a_12691_2527# VPWR 0.375f
C14047 a_7933_11305# VPWR 1.16e-19
C14048 net43 a_3565_7119# 0.00206f
C14049 a_6885_8372# _002_ 1.05e-19
C14050 a_763_8757# a_1476_7119# 4.8e-19
C14051 _114_ VPWR 0.274f
C14052 _048_ a_3817_4697# 0.0416f
C14053 trim_mask\[4\] a_8298_2767# 2.14e-19
C14054 a_13783_6183# clkc 7.43e-20
C14055 en_co_clk a_14379_6397# 0.0927f
C14056 clknet_2_1__leaf_clk a_4696_8207# 6.67e-22
C14057 a_5363_4719# VPWR 0.00535f
C14058 a_3597_12021# a_3947_12393# 0.22f
C14059 a_3431_12021# a_4687_12319# 0.0436f
C14060 net13 _040_ 0.171f
C14061 _047_ _058_ 2.25e-19
C14062 _101_ a_6181_10633# 0.0106f
C14063 a_9595_1679# a_10851_1653# 0.0436f
C14064 _032_ a_10111_1679# 0.00164f
C14065 a_4425_6031# _099_ 7.41e-21
C14066 a_14335_4020# trim_mask\[2\] 6.01e-22
C14067 trim_mask\[1\] _025_ 0.12f
C14068 a_13257_1141# _057_ 5.45e-20
C14069 net33 a_15023_1679# 0.11f
C14070 a_9529_6059# _107_ 8.43e-20
C14071 trim_mask\[1\] _026_ 1.47e-19
C14072 net26 a_448_9269# 6.71e-20
C14073 cal_count\[3\] _118_ 0.0221f
C14074 a_14193_3285# a_14099_3017# 2.18e-19
C14075 clknet_2_0__leaf_clk _048_ 7.83e-20
C14076 a_4167_11471# a_3431_10933# 4.34e-20
C14077 a_5423_9011# net51 9.02e-20
C14078 _065_ a_6485_8181# 0.0772f
C14079 cal_count\[1\] _129_ 0.0153f
C14080 net46 a_9773_3689# 2.95e-19
C14081 en_co_clk _038_ 2.04e-19
C14082 net22 a_1493_5487# 0.00758f
C14083 _103_ a_7891_3617# 3.34e-21
C14084 a_7351_8041# a_7459_7663# 0.0572f
C14085 a_8091_7967# a_8270_8029# 0.0074f
C14086 a_7916_8041# a_8025_8041# 0.00742f
C14087 a_13050_7637# VPWR 0.234f
C14088 a_561_6031# a_816_6031# 0.0642f
C14089 _034_ a_4993_6273# 3.46e-19
C14090 a_2313_6183# VPWR 0.186f
C14091 net30 calibrate 0.00261f
C14092 a_4959_1679# VPWR 0.205f
C14093 _001_ a_10975_6031# 5.83e-20
C14094 a_10975_6031# a_11067_4405# 4.43e-21
C14095 a_14983_9269# _128_ 3.1e-21
C14096 net47 a_10861_7119# 8.02e-19
C14097 net18 _110_ 0.0157f
C14098 clknet_2_1__leaf_clk _023_ 0.184f
C14099 a_6375_12021# a_7565_12393# 2.56e-19
C14100 a_7477_10901# VPWR 0.22f
C14101 _132_ a_15023_6031# 4.11e-22
C14102 net34 a_15023_10927# 0.0153f
C14103 net29 a_1203_12015# 9.55e-19
C14104 a_8072_11721# net12 4.73e-20
C14105 a_8749_3317# _025_ 1.26e-20
C14106 net43 result[3] 6.6e-20
C14107 trim_mask\[0\] a_13059_4631# 0.0743f
C14108 trim_mask\[0\] net35 0.012f
C14109 net33 a_15023_6031# 0.00552f
C14110 a_2948_3689# a_2309_2229# 9.92e-21
C14111 a_2383_3689# a_2659_2601# 9.85e-20
C14112 _053_ a_11098_6691# 3.68e-19
C14113 a_7897_6913# VPWR 1.48e-19
C14114 _064_ net50 0.465f
C14115 mask\[1\] a_2225_7983# 0.00256f
C14116 net44 mask\[3\] 0.295f
C14117 en_co_clk a_4617_4105# 7.06e-19
C14118 net46 a_9003_3829# 7.7e-19
C14119 _068_ a_9602_6941# 2.88e-19
C14120 net14 a_1007_4777# 7.18e-19
C14121 net13 _048_ 0.00631f
C14122 net9 net10 2.17e-19
C14123 net44 a_6741_7361# 0.168f
C14124 _065_ a_6007_7119# 9.37e-21
C14125 _107_ a_9369_4105# 0.00207f
C14126 a_745_12021# _086_ 8.56e-20
C14127 mask\[5\] a_8178_11293# 6.42e-19
C14128 _113_ a_14715_3615# 3.12e-21
C14129 net5 _136_ 5.3e-20
C14130 _074_ a_995_3530# 0.00827f
C14131 a_3521_9813# a_4030_9839# 2.6e-19
C14132 a_4655_10071# a_5089_10159# 0.00393f
C14133 a_2953_9845# a_4801_9839# 2.5e-19
C14134 net12 _094_ 1.21e-20
C14135 net18 a_10699_5487# 0.0108f
C14136 _088_ a_5537_4105# 9.11e-21
C14137 net18 a_12148_4777# 5.62e-19
C14138 clknet_2_1__leaf_clk a_816_10205# 0.0289f
C14139 a_4864_9295# _040_ 2.36e-19
C14140 net47 a_11987_8757# 0.0527f
C14141 net33 net46 0.0155f
C14142 a_4165_11989# VPWR 0.225f
C14143 a_9503_4399# a_8583_3317# 1.96e-20
C14144 net16 _131_ 0.0107f
C14145 a_11023_5108# _104_ 2.43e-21
C14146 a_1129_7361# a_911_6031# 7.82e-20
C14147 a_911_7119# a_1129_6273# 2.14e-20
C14148 net50 a_10851_1653# 0.00823f
C14149 a_2828_12131# _046_ 0.106f
C14150 clknet_2_2__leaf_clk a_9761_1679# 0.00249f
C14151 _092_ state\[1\] 0.00946f
C14152 mask\[1\] a_4131_8207# 0.0346f
C14153 net43 a_2014_11293# 0.00288f
C14154 a_4576_3427# a_4815_3031# 3.85e-19
C14155 net32 VPWR 0.552f
C14156 _019_ VPWR 0.476f
C14157 a_12900_7663# _133_ 0.0121f
C14158 net28 a_4687_12319# 0.15f
C14159 _090_ a_3891_4943# 0.00181f
C14160 a_1493_11721# VPWR 0.24f
C14161 _094_ a_5340_6031# 0.004f
C14162 net30 a_8298_5487# 0.00182f
C14163 a_4259_6031# a_4425_6031# 0.855f
C14164 _123_ a_13356_8457# 0.00337f
C14165 a_6741_7361# clk 6.33e-21
C14166 trim_val\[0\] _110_ 0.00507f
C14167 cal_count\[3\] a_10137_4943# 1.1e-19
C14168 _065_ _092_ 0.0108f
C14169 _104_ a_10055_2767# 0.0101f
C14170 net45 a_1585_7119# 6.07e-20
C14171 a_7223_2465# _027_ 4.98e-19
C14172 a_7184_2339# a_8491_2229# 0.00133f
C14173 a_7379_2197# a_7310_2223# 0.21f
C14174 mask\[6\] net52 0.201f
C14175 mask\[5\] a_7259_11305# 2.57e-19
C14176 net28 net13 3.54e-20
C14177 a_9020_10383# a_9871_10383# 2.94e-19
C14178 a_9195_10357# _042_ 0.0354f
C14179 net13 a_5177_9537# 9.37e-19
C14180 net15 net41 0.00739f
C14181 _000_ net2 9.24e-22
C14182 a_11233_4405# a_11067_3017# 7.13e-19
C14183 a_5878_1679# VPWR 0.00178f
C14184 _061_ trim_mask\[0\] 5.78e-19
C14185 net43 a_2787_10927# 1.31e-19
C14186 _050_ net42 0.00488f
C14187 a_4871_8181# net51 2e-20
C14188 a_4696_8207# a_6485_8181# 5.98e-21
C14189 a_6467_9845# VPWR 0.423f
C14190 trim_val\[0\] a_12148_4777# 1.75e-21
C14191 a_14334_5309# _058_ 3.02e-20
C14192 _076_ net51 0.092f
C14193 a_2948_3689# a_3110_3311# 0.00645f
C14194 net54 _088_ 6.12e-21
C14195 trim_val\[4\] a_10699_3311# 0.00148f
C14196 _097_ a_2283_4020# 0.183f
C14197 _051_ a_8749_3317# 0.00327f
C14198 a_8993_9295# _063_ 6.23e-21
C14199 net25 a_3521_9813# 4.62e-21
C14200 _051_ _060_ 0.26f
C14201 mask\[2\] net45 6.57e-20
C14202 _050_ a_4091_5309# 0.00179f
C14203 net16 a_14281_4943# 1.59e-19
C14204 a_8083_8181# cal_itt\[2\] 0.00349f
C14205 trim_mask\[1\] _031_ 2.04e-20
C14206 net3 a_5081_4943# 0.0409f
C14207 a_14193_3285# net48 6.02e-21
C14208 a_4043_7093# a_4425_6031# 3.92e-20
C14209 _028_ a_7524_2223# 0.00136f
C14210 a_3868_7119# a_4259_6031# 3.29e-20
C14211 a_3578_2589# clk 2.24e-19
C14212 net42 _052_ 5.72e-21
C14213 a_3840_8867# _041_ 0.109f
C14214 calibrate state\[2\] 0.62f
C14215 _104_ a_6927_3311# 0.0126f
C14216 a_1769_12393# VPWR 1.22e-19
C14217 a_448_7637# result[1] 0.157f
C14218 _093_ a_3339_2767# 2.06e-20
C14219 cal_count\[1\] a_14318_8457# 0.00101f
C14220 _112_ a_13415_2442# 4.98e-19
C14221 trim_mask\[0\] a_13257_4943# 0.00645f
C14222 net46 trim_val\[3\] 0.075f
C14223 a_395_9845# a_2787_9845# 5.48e-21
C14224 net55 net3 0.134f
C14225 a_12218_6397# VPWR 4.89e-19
C14226 net26 a_6099_10633# 8.35e-19
C14227 calibrate state\[0\] 0.00673f
C14228 net42 _098_ 0.174f
C14229 a_4165_11989# net27 2.51e-21
C14230 a_9664_3689# trim_mask\[2\] 1.12e-19
C14231 a_5699_9269# VPWR 0.404f
C14232 net54 a_6519_4631# 1.39e-19
C14233 _107_ a_8307_4719# 0.00512f
C14234 _118_ _119_ 3.49e-19
C14235 net28 a_1203_12015# 0.00362f
C14236 a_5535_8181# a_5363_7369# 7.42e-20
C14237 a_4167_11471# net13 2.62e-19
C14238 a_15023_6031# _136_ 3.66e-21
C14239 a_10990_7485# cal_count\[3\] 9.6e-21
C14240 _125_ a_14788_7369# 6.58e-20
C14241 _076_ _003_ 0.149f
C14242 net34 a_14686_2339# 2.58e-19
C14243 clknet_2_3__leaf_clk a_13783_6183# 0.117f
C14244 net27 _019_ 4.53e-21
C14245 _074_ net3 3.09e-20
C14246 a_7001_7669# a_7088_7119# 2.86e-19
C14247 a_6835_7669# a_8022_7119# 7.19e-20
C14248 trim_mask\[1\] a_10781_3311# 0.0163f
C14249 a_7569_7637# a_7263_7093# 0.00118f
C14250 trim_mask\[2\] a_10689_2223# 8.17e-20
C14251 a_4609_9295# a_5067_9661# 0.0306f
C14252 a_4959_9295# a_5524_9295# 7.99e-20
C14253 trim_mask\[3\] net10 0.00217f
C14254 net21 a_4687_12319# 0.00744f
C14255 a_12424_3689# a_12586_3311# 0.00645f
C14256 a_13459_3317# a_13880_3677# 0.0864f
C14257 net27 a_1493_11721# 0.0472f
C14258 net47 a_9296_9295# 0.251f
C14259 a_10688_9295# cal_count\[0\] 0.00994f
C14260 _064_ _106_ 0.00126f
C14261 net45 a_6428_7119# 4.42e-22
C14262 clknet_2_1__leaf_clk _078_ 0.0378f
C14263 a_3947_11305# a_4512_11305# 7.99e-20
C14264 _101_ a_5535_8181# 0.0126f
C14265 net34 net5 0.217f
C14266 net2 trimb[4] 1.08e-19
C14267 a_7001_7669# _063_ 7.72e-20
C14268 _039_ _049_ 1.46e-19
C14269 a_6541_12021# net53 5.31e-20
C14270 mask\[3\] a_4801_9839# 0.0051f
C14271 _038_ a_12410_6031# 3.39e-20
C14272 a_3868_10217# mask\[2\] 0.00219f
C14273 net46 _136_ 0.0557f
C14274 _123_ a_12522_8751# 0.00224f
C14275 net45 a_2143_2229# 0.299f
C14276 _129_ a_12900_7663# 4.17e-19
C14277 net14 a_1007_7119# 7.18e-19
C14278 _107_ a_7010_3631# 7.02e-20
C14279 a_13697_4373# a_13459_3317# 8.6e-21
C14280 _058_ a_13183_3311# 0.00186f
C14281 a_3521_7361# a_3411_7485# 0.0977f
C14282 mask\[5\] _008_ 1.37e-19
C14283 a_4043_7093# a_3868_7119# 0.234f
C14284 a_3303_7119# a_3208_7119# 0.0498f
C14285 a_1095_11305# a_561_9845# 5.84e-21
C14286 clknet_2_0__leaf_clk a_2033_3317# 0.00439f
C14287 _007_ a_455_8181# 4.85e-19
C14288 _048_ a_4091_4943# 0.00353f
C14289 _060_ a_5445_4399# 2.06e-19
C14290 a_14564_6397# trim_val\[0\] 1.02e-19
C14291 net19 a_7800_4631# 5.86e-21
C14292 _110_ a_10055_2767# 0.00447f
C14293 net21 net13 0.13f
C14294 net43 _049_ 0.006f
C14295 net12 a_7088_7119# 0.00227f
C14296 a_9478_4105# VPWR 0.237f
C14297 a_7999_11231# _020_ 8.91e-19
C14298 net15 a_2767_2223# 0.00245f
C14299 net9 a_12916_8751# 2.92e-19
C14300 _108_ a_12323_4703# 1.58e-19
C14301 a_10699_5487# a_11023_5108# 1.03e-19
C14302 net9 a_10975_6031# 0.00101f
C14303 _101_ _082_ 8.79e-21
C14304 trim[3] ctln[2] 2.75e-19
C14305 ctln[7] ctln[6] 0.00465f
C14306 cal_itt\[0\] net40 5.38e-21
C14307 a_7019_4407# _088_ 0.00314f
C14308 trim_mask\[2\] a_10781_3631# 4.58e-19
C14309 net34 a_14347_1439# 0.0166f
C14310 net27 a_6467_9845# 1.98e-21
C14311 _110_ a_9926_2589# 4.63e-19
C14312 a_8749_3317# a_10781_3311# 1.7e-19
C14313 a_9317_3285# a_9826_3311# 2.6e-19
C14314 a_4775_6031# _095_ 3.65e-19
C14315 _067_ _092_ 0.0862f
C14316 a_7262_5461# a_7019_4407# 4.91e-19
C14317 clknet_2_2__leaf_clk a_11067_3017# 0.0569f
C14318 _078_ a_2368_9955# 5.82e-19
C14319 trim_mask\[2\] a_14184_1679# 0.0101f
C14320 clknet_0_clk a_8307_6575# 0.0106f
C14321 a_1129_9813# a_1638_9839# 2.6e-19
C14322 net45 a_4815_3031# 2.97e-19
C14323 _051_ a_7939_3855# 0.0094f
C14324 _090_ a_3530_4438# 1.53e-19
C14325 _058_ a_11691_4399# 0.00331f
C14326 a_13697_4373# _109_ 0.125f
C14327 net47 cal_count\[3\] 9.79e-21
C14328 net40 a_15259_7637# 2.19e-20
C14329 a_9459_7895# en_co_clk 1.18e-19
C14330 net38 a_14983_9269# 4.06e-21
C14331 clknet_0_clk a_7460_5807# 0.0521f
C14332 a_395_7119# a_1007_7119# 0.00188f
C14333 a_11343_3317# trim_val\[3\] 8.55e-21
C14334 net44 clk 0.00764f
C14335 a_13091_4943# trim_val\[0\] 1.33e-19
C14336 net44 en_co_clk 0.165f
C14337 a_13825_5185# a_13703_4943# 3.16e-19
C14338 net27 VPWR 1.22f
C14339 clknet_2_3__leaf_clk a_13142_7271# 1.63e-19
C14340 a_11149_3017# trim_val\[3\] 3.19e-20
C14341 net12 ctln[6] 0.02f
C14342 _053_ _106_ 0.00112f
C14343 _115_ _031_ 0.00257f
C14344 _134_ _135_ 0.259f
C14345 _051_ a_4498_4373# 1.22e-21
C14346 _064_ _033_ 0.00276f
C14347 net14 net41 0.0116f
C14348 _045_ a_6927_12559# 6.23e-19
C14349 _021_ a_7355_11305# 1.9e-19
C14350 a_5915_10927# a_5997_10927# 0.171f
C14351 calibrate _100_ 0.631f
C14352 _084_ mask\[4\] 3.07e-20
C14353 a_6741_7361# a_7197_7119# 4.2e-19
C14354 net44 a_8386_8457# 2.86e-19
C14355 a_4498_4373# _014_ 1.2e-20
C14356 a_6519_4631# a_7019_4407# 7.45e-19
C14357 _058_ net49 0.00402f
C14358 net2 _053_ 8.1e-20
C14359 clknet_2_1__leaf_clk a_3597_10933# 0.00758f
C14360 a_14807_8359# VPWR 0.212f
C14361 net31 trimb[4] 0.109f
C14362 net43 a_3947_12393# 0.161f
C14363 a_1660_12393# mask\[7\] 8.56e-19
C14364 a_9889_6873# a_10005_6031# 0.0015f
C14365 a_1476_4777# a_1638_4399# 0.00645f
C14366 a_911_7119# result[1] 2.56e-19
C14367 net34 a_15023_1679# 0.0156f
C14368 _110_ a_12691_2527# 2.51e-19
C14369 a_6793_8970# _041_ 0.0359f
C14370 _126_ a_14467_8751# 0.0549f
C14371 clknet_2_3__leaf_clk a_14181_6031# 0.0029f
C14372 _110_ _114_ 0.103f
C14373 a_1099_12533# ctlp[0] 0.338f
C14374 a_9664_3689# a_9595_1679# 1.46e-19
C14375 net3 _093_ 0.0565f
C14376 a_11895_7669# a_12344_8041# 0.211f
C14377 a_9369_4105# trim_mask\[4\] 1.27e-19
C14378 _037_ a_12520_7637# 7.99e-19
C14379 _107_ a_6822_4399# 3.55e-19
C14380 _023_ result[4] 5.22e-19
C14381 en_co_clk clk 0.00988f
C14382 net43 a_3425_11721# 1.63e-19
C14383 a_4167_6575# _048_ 8.48e-21
C14384 cal_count\[0\] cal_count\[1\] 0.112f
C14385 a_763_8757# a_1125_7663# 1.24e-20
C14386 net3 a_5166_5193# 2.21e-19
C14387 a_12341_8751# a_12546_9129# 3.7e-19
C14388 mask\[2\] a_3922_8867# 3.43e-19
C14389 net52 a_3317_8207# 0.00141f
C14390 a_10689_2223# a_9595_1679# 8.28e-19
C14391 _045_ _009_ 0.00719f
C14392 net20 _084_ 0.00131f
C14393 _121_ a_4259_6031# 0.051f
C14394 net34 a_15023_12015# 0.0944f
C14395 _042_ a_3303_10217# 0.0026f
C14396 net18 a_11057_4105# 0.00587f
C14397 a_2383_3689# VPWR 0.209f
C14398 net37 a_15023_5487# 0.0127f
C14399 a_10239_9295# a_11168_9661# 0.00294f
C14400 net34 a_15023_6031# 0.00426f
C14401 _035_ a_10774_9661# 3.7e-19
C14402 _049_ a_6822_4399# 3.21e-19
C14403 a_14063_7093# _134_ 0.082f
C14404 _074_ a_448_9269# 4.25e-19
C14405 calibrate _012_ 0.189f
C14406 a_3273_4943# _099_ 7.1e-21
C14407 _064_ a_10785_1679# 3.56e-20
C14408 a_2857_7637# _049_ 0.00147f
C14409 net4 a_3339_2767# 0.213f
C14410 a_3840_8867# a_3615_8207# 8.61e-19
C14411 a_816_10205# result[4] 6.75e-19
C14412 _072_ _073_ 0.00309f
C14413 a_13257_4943# _030_ 6.47e-22
C14414 _038_ _108_ 1.47e-19
C14415 _048_ _028_ 8.13e-20
C14416 clknet_2_2__leaf_clk a_6906_2355# 1.1e-19
C14417 a_14471_12559# net39 0.01f
C14418 net40 trim_mask\[0\] 0.00625f
C14419 a_8455_10383# VPWR 0.197f
C14420 trim_mask\[2\] _057_ 2.32e-20
C14421 _074_ mask\[0\] 1.13e-20
C14422 net45 a_5087_3855# 1.48e-20
C14423 _078_ a_1953_9129# 0.0011f
C14424 net4 rstn 0.00313f
C14425 _122_ a_13008_7663# 2.73e-19
C14426 _104_ VPWR 1.95f
C14427 _074_ valid 0.0171f
C14428 a_2971_8457# a_3615_8207# 2.32e-20
C14429 net5 a_15299_6575# 0.197f
C14430 a_14083_3311# net48 6.72e-21
C14431 a_1467_7923# a_1651_6005# 3.85e-22
C14432 a_9650_9295# VPWR 2.56e-19
C14433 _034_ net3 2.54e-21
C14434 a_2815_9447# net24 5.06e-20
C14435 net55 a_5537_4105# 2.48e-19
C14436 net34 net46 0.00589f
C14437 _122_ a_13256_9117# 9.69e-20
C14438 net2 _130_ 0.137f
C14439 net47 a_9463_8725# 0.19f
C14440 net45 a_4443_1679# 0.297f
C14441 _048_ a_3751_4765# 0.00406f
C14442 cal_count\[0\] a_12612_8725# 0.0264f
C14443 net43 a_2014_12381# 0.00288f
C14444 a_1313_11989# a_1203_12015# 0.0977f
C14445 net19 a_7548_10217# 5.66e-19
C14446 net53 a_7079_10217# 6.89e-19
C14447 net45 a_1476_4777# 0.245f
C14448 a_7393_5193# _103_ 0.0123f
C14449 net19 net18 3.97e-19
C14450 net14 a_2767_2223# 2.17e-19
C14451 mask\[3\] result[3] 1.45e-19
C14452 net14 a_1137_5487# 9.08e-19
C14453 a_14335_4020# a_14193_3285# 7.71e-20
C14454 a_2019_9055# a_1651_7093# 4.89e-20
C14455 net12 a_5455_4943# 2.37e-20
C14456 clknet_2_2__leaf_clk a_9317_3285# 0.00214f
C14457 state\[2\] _015_ 8.91e-20
C14458 a_929_8757# a_1019_7485# 4.01e-21
C14459 net50 a_9664_3689# 1.67e-20
C14460 a_4043_7093# _121_ 0.00141f
C14461 net44 _059_ 0.00165f
C14462 net31 trim[0] 0.0191f
C14463 a_7200_3631# VPWR 1.94e-19
C14464 _120_ a_3557_5193# 6.75e-19
C14465 a_8105_10383# a_8563_10749# 0.0276f
C14466 net26 _076_ 0.00189f
C14467 state\[0\] _015_ 0.268f
C14468 a_1099_12533# a_579_12021# 0.0023f
C14469 _077_ a_6198_8534# 1.1e-19
C14470 a_8091_7967# clk 0.00454f
C14471 net50 a_10689_2223# 0.00887f
C14472 clknet_2_2__leaf_clk a_11856_2589# 1.12e-19
C14473 a_4871_8181# a_5050_8207# 0.0074f
C14474 net32 _110_ 4.19e-20
C14475 a_4696_8207# a_4805_8207# 0.00742f
C14476 net42 a_8389_5193# 0.0131f
C14477 a_2313_6183# a_2476_6281# 0.00477f
C14478 a_1651_6005# _094_ 8.61e-21
C14479 a_561_7119# a_1549_6794# 7.99e-20
C14480 a_5340_6031# a_5455_4943# 9.99e-20
C14481 clk ctln[0] 0.0136f
C14482 trim_val\[2\] a_13703_1513# 1.48e-19
C14483 net24 _081_ 0.277f
C14484 _074_ _079_ 0.0789f
C14485 a_6173_7119# a_6619_7119# 2.28e-19
C14486 a_6741_7361# a_7250_7485# 2.6e-19
C14487 a_10864_7387# a_10903_7261# 0.827f
C14488 a_10586_7371# a_11059_7356# 7.99e-20
C14489 net53 a_7723_10143# 2.38e-20
C14490 clknet_2_1__leaf_clk a_7001_7669# 9.3e-19
C14491 a_10569_1109# _116_ 0.115f
C14492 net18 cal_itt\[1\] 2.96e-20
C14493 _117_ a_9805_1473# 5.76e-19
C14494 _035_ _065_ 5.27e-20
C14495 net54 a_5081_4943# 0.00733f
C14496 _104_ a_9478_4105# 5.82e-19
C14497 a_12077_3285# a_11859_3689# 0.21f
C14498 a_11509_3317# a_12599_3615# 0.0424f
C14499 a_7456_12393# a_7565_12393# 0.00742f
C14500 a_6891_12393# a_6999_12015# 0.0572f
C14501 a_8381_9295# VPWR 0.581f
C14502 a_7631_12319# a_7810_12381# 0.0074f
C14503 net44 a_8992_9955# 1.91e-19
C14504 _042_ a_1019_9839# 1.29e-20
C14505 _128_ _133_ 5.69e-19
C14506 net19 a_9129_10383# 2.55e-19
C14507 _053_ _054_ 0.339f
C14508 en_co_clk _059_ 0.091f
C14509 net8 trim[3] 2.86e-19
C14510 net44 a_7197_7119# 6.03e-19
C14511 cal_itt\[0\] _071_ 9.45e-19
C14512 net31 _130_ 0.00142f
C14513 a_579_10933# net26 0.00144f
C14514 _023_ a_448_10357# 0.00178f
C14515 mask\[4\] a_4801_10159# 5.55e-19
C14516 net55 net54 0.395f
C14517 a_10005_6031# a_11141_6031# 3.72e-19
C14518 net35 a_15083_4659# 0.00348f
C14519 net16 a_13693_3883# 4.09e-19
C14520 net31 a_14335_4020# 6.95e-19
C14521 clknet_2_1__leaf_clk a_6888_10205# 1.68e-20
C14522 cal_count\[2\] en_co_clk 1.66e-19
C14523 _134_ a_13279_7119# 0.00196f
C14524 a_1007_4777# VPWR 8.62e-19
C14525 a_395_6031# a_561_6031# 0.806f
C14526 a_12678_2223# VPWR 8.28e-19
C14527 clknet_2_1__leaf_clk net12 1.46f
C14528 _101_ a_3133_11247# 3.04e-19
C14529 _013_ cal 4.03e-19
C14530 _093_ valid 9.09e-19
C14531 trim_mask\[4\] a_7010_3631# 1.83e-20
C14532 _065_ _136_ 0.0334f
C14533 net15 a_3063_591# 0.00137f
C14534 a_3615_8207# a_4131_8207# 0.11f
C14535 trim_mask\[0\] _024_ 0.123f
C14536 a_3781_8207# a_4349_8449# 0.181f
C14537 net42 a_7891_3617# 3.84e-21
C14538 _045_ mask\[6\] 0.0215f
C14539 net45 _120_ 4.53e-21
C14540 a_8298_5487# _118_ 2.47e-19
C14541 a_10329_1921# _116_ 1.75e-20
C14542 _032_ a_10872_1455# 7.95e-20
C14543 a_13919_8751# cal_count\[1\] 0.0563f
C14544 a_3891_4943# a_3667_3829# 1.86e-20
C14545 net2 a_13821_7119# 1.11e-19
C14546 _110_ VPWR 3.18f
C14547 a_9802_4007# a_10270_4105# 1.25e-19
C14548 _067_ a_9602_6941# 1.53e-20
C14549 net4 net3 0.416f
C14550 clknet_0_clk VPWR 3.19f
C14551 _078_ result[4] 5.53e-20
C14552 _128_ a_14236_8457# 2.16e-20
C14553 clknet_2_3__leaf_clk a_10055_5487# 0.0227f
C14554 _113_ a_13183_3311# 0.201f
C14555 a_7263_7093# a_7723_6807# 0.00131f
C14556 a_14983_9269# net40 1.78e-19
C14557 clknet_2_2__leaf_clk a_9003_3829# 5.22e-19
C14558 _126_ a_14249_8725# 8.39e-19
C14559 a_3224_2601# a_3333_2601# 0.00742f
C14560 net31 a_15023_2767# 0.235f
C14561 a_2659_2601# a_2767_2223# 0.0572f
C14562 a_3399_2527# a_3578_2589# 0.0074f
C14563 net18 _001_ 0.00937f
C14564 net47 a_10383_7093# 0.286f
C14565 _100_ _015_ 3.26e-20
C14566 net18 a_11067_4405# 0.0237f
C14567 a_12778_3677# VPWR 1.46e-19
C14568 clknet_2_1__leaf_clk a_6983_10217# 3.51e-20
C14569 a_395_9845# a_763_8757# 2.63e-19
C14570 _108_ a_10270_4105# 5.77e-19
C14571 a_7351_8041# a_7916_8041# 7.99e-20
C14572 _074_ a_448_6549# 0.00596f
C14573 a_2033_3317# a_2948_3689# 0.125f
C14574 a_1867_3317# a_4576_3427# 6.01e-22
C14575 _101_ a_4165_10901# 1.37e-19
C14576 a_5087_3855# a_4905_3855# 1.5e-19
C14577 _074_ a_6099_10633# 4.66e-19
C14578 a_6198_8207# VPWR 2.26e-19
C14579 _094_ _048_ 0.00253f
C14580 a_10699_5487# VPWR 0.216f
C14581 a_12148_4777# VPWR 0.309f
C14582 a_11895_7669# _133_ 2.33e-22
C14583 _002_ net30 0.00184f
C14584 net13 _077_ 2.18e-20
C14585 cal_count\[0\] a_12900_7663# 2.03e-20
C14586 mask\[0\] _034_ 8.13e-22
C14587 net26 clknet_2_3__leaf_clk 8.28e-19
C14588 net46 cal_count\[3\] 0.0794f
C14589 a_4609_9295# net45 5.96e-21
C14590 clknet_2_1__leaf_clk a_3852_12381# 0.0149f
C14591 trim_mask\[1\] _055_ 0.00218f
C14592 net30 _050_ 4.74e-19
C14593 _049_ a_4617_4105# 0.00162f
C14594 _136_ a_11233_4405# 0.0014f
C14595 _072_ a_8078_7663# 5.67e-19
C14596 a_8022_7119# a_9443_6059# 8.11e-20
C14597 net44 a_5694_6031# 0.00312f
C14598 _053_ a_12249_7663# 8.64e-20
C14599 net26 a_395_9845# 1.7e-19
C14600 a_3748_6281# a_4425_6031# 2.71e-19
C14601 clknet_2_1__leaf_clk a_1651_10143# 0.0376f
C14602 a_7459_7663# VPWR 0.144f
C14603 net55 a_7019_4407# 0.181f
C14604 _113_ net49 0.0029f
C14605 state\[2\] a_7184_2339# 1.43e-20
C14606 _106_ a_9664_3689# 3.75e-20
C14607 mask\[4\] a_6181_10383# 0.00134f
C14608 _063_ _091_ 0.0171f
C14609 cal_itt\[0\] _123_ 0.00309f
C14610 _065_ a_10861_7119# 2.55e-19
C14611 _110_ a_9478_4105# 0.00536f
C14612 _051_ a_7571_4943# 2.15e-20
C14613 net55 a_4471_4007# 0.149f
C14614 a_2283_4020# a_2288_3677# 5.77e-19
C14615 net30 _052_ 1.34e-20
C14616 a_2476_6281# VPWR 0.00231f
C14617 net50 _057_ 8.88e-20
C14618 a_1129_4373# a_937_4105# 3.22e-19
C14619 _128_ _129_ 4.32e-20
C14620 _065_ a_4266_4943# 7.4e-21
C14621 a_7939_10383# a_8105_10383# 0.9f
C14622 a_3521_9813# VPWR 0.218f
C14623 net42 _087_ 2.68e-20
C14624 net44 a_7618_12015# 3.47e-19
C14625 trim_mask\[2\] a_13625_3317# 2.63e-20
C14626 net30 _098_ 8.93e-20
C14627 a_561_6031# net30 1.28e-19
C14628 net54 _093_ 0.0386f
C14629 _122_ a_12520_7637# 0.00191f
C14630 a_13697_4373# trim[1] 4.51e-20
C14631 _095_ a_1651_4703# 8.55e-19
C14632 _051_ a_4576_3427# 1.82e-20
C14633 net51 a_6835_7669# 0.0281f
C14634 a_6741_7361# _049_ 4.88e-20
C14635 a_1651_10143# a_2368_9955# 9.04e-19
C14636 a_9602_6614# net30 8.83e-21
C14637 en_co_clk a_5694_6031# 5.11e-19
C14638 a_4655_10071# a_4443_9295# 2.75e-19
C14639 net44 a_7250_7485# 2.98e-19
C14640 a_7527_4631# a_7010_3311# 4.03e-19
C14641 a_14335_4020# a_14083_3311# 1.13e-19
C14642 net16 a_14237_3677# 0.00127f
C14643 _022_ a_3133_11247# 1.97e-19
C14644 net31 a_15299_3311# 0.00232f
C14645 a_3431_10933# a_3852_11293# 0.0897f
C14646 a_2953_7119# _120_ 1.44e-20
C14647 _104_ a_7200_3631# 5.22e-19
C14648 a_9225_2197# a_9103_2601# 3.16e-19
C14649 a_9007_2601# a_8912_2589# 0.0498f
C14650 trim_mask\[0\] _029_ 0.00237f
C14651 a_6983_10217# a_7245_10205# 0.00171f
C14652 a_7201_9813# a_7657_10217# 4.2e-19
C14653 _111_ a_11845_4765# 1.11e-19
C14654 net1 a_855_4105# 0.0853f
C14655 a_3868_7119# a_3748_6281# 4.85e-20
C14656 net55 a_4970_4399# 7.38e-19
C14657 _068_ a_9463_8725# 3.24e-19
C14658 a_14564_6397# VPWR 0.209f
C14659 mask\[0\] a_3830_6281# 6.75e-20
C14660 _074_ a_5423_9011# 0.334f
C14661 a_4036_8207# a_2857_7637# 9.72e-19
C14662 a_8583_3317# trim_mask\[2\] 2.46e-19
C14663 _033_ a_9664_3689# 1.94e-21
C14664 clknet_2_2__leaf_clk trim_val\[3\] 0.00266f
C14665 clknet_2_1__leaf_clk result[2] 2.89e-20
C14666 _067_ _136_ 8.31e-19
C14667 a_4091_5309# _099_ 4.16e-20
C14668 cal_itt\[0\] a_9043_6031# 3.38e-19
C14669 clknet_2_0__leaf_clk a_6173_7119# 0.00196f
C14670 _074_ a_1229_8457# 0.00107f
C14671 a_1007_7119# VPWR 7.36e-19
C14672 a_8455_10383# a_8381_9295# 2.56e-20
C14673 a_7001_7669# a_6007_7119# 1.34e-19
C14674 calibrate a_3933_2767# 1.95e-20
C14675 a_14467_8751# VPWR 0.282f
C14676 net47 a_8215_9295# 0.304f
C14677 a_10405_9295# a_11244_9661# 0.0573f
C14678 a_8949_9537# a_9405_9295# 4.2e-19
C14679 a_1137_11721# ctlp[0] 4.39e-19
C14680 a_1019_6397# result[0] 5.48e-19
C14681 _022_ a_4165_10901# 7.67e-19
C14682 trim_val\[1\] a_14604_3017# 0.239f
C14683 a_3431_10933# a_3947_11305# 0.111f
C14684 a_3399_2527# clk 0.00588f
C14685 a_13091_4943# VPWR 0.484f
C14686 cal_itt\[1\] a_8307_6575# 7.64e-19
C14687 net51 a_5515_6005# 9.5e-20
C14688 a_9747_2527# a_9572_2601# 0.234f
C14689 net53 _042_ 0.369f
C14690 net18 a_11394_9509# 0.00254f
C14691 net37 a_15023_8751# 0.00597f
C14692 _038_ a_11587_6031# 0.00196f
C14693 a_2787_9845# mask\[2\] 9e-19
C14694 a_6375_12021# a_6541_12021# 0.897f
C14695 _129_ a_11895_7669# 1.16e-20
C14696 _108_ clk 2.39e-21
C14697 en_co_clk _108_ 7.36e-21
C14698 _125_ _122_ 8.39e-20
C14699 _058_ _025_ 0.00193f
C14700 _065_ _073_ 3.23e-20
C14701 clknet_2_1__leaf_clk a_6631_7485# 7.92e-19
C14702 _136_ clknet_2_2__leaf_clk 0.00225f
C14703 _058_ _026_ 4.85e-19
C14704 net12 a_6007_7119# 0.0176f
C14705 a_11023_5108# a_11067_4405# 3.91e-19
C14706 _108_ a_9084_4515# 0.00179f
C14707 _064_ a_11413_2767# 6.38e-21
C14708 mask\[0\] a_3303_7119# 0.036f
C14709 a_1830_10205# VPWR 2.01e-19
C14710 _050_ state\[2\] 0.711f
C14711 net41 VPWR 0.501f
C14712 net29 _011_ 0.00552f
C14713 _120_ a_2857_5461# 0.0439f
C14714 _104_ _110_ 0.0117f
C14715 _071_ a_8949_6281# 4.88e-19
C14716 a_7001_7669# _092_ 1.07e-20
C14717 net45 a_1867_3317# 0.305f
C14718 a_10864_9269# a_11116_8983# 1.79e-19
C14719 a_10405_9295# _123_ 0.00678f
C14720 a_561_7119# a_1019_7485# 0.0346f
C14721 a_911_7119# a_1476_7119# 7.99e-20
C14722 _054_ a_7379_2197# 1.12e-20
C14723 net46 a_14347_4917# 0.282f
C14724 clknet_0_clk _104_ 0.0857f
C14725 net31 trim[4] 0.109f
C14726 _050_ state\[0\] 5.44e-19
C14727 _093_ a_4471_4007# 0.0328f
C14728 net18 a_11116_8983# 0.0103f
C14729 _074_ a_1125_7663# 0.0208f
C14730 _067_ a_10861_7119# 1.37e-19
C14731 mask\[7\] a_1095_11305# 0.00755f
C14732 _112_ a_13880_3677# 0.00367f
C14733 _063_ _048_ 0.268f
C14734 _029_ a_13869_4943# 9.23e-20
C14735 net44 a_8178_11293# 0.00323f
C14736 a_9460_6807# en_co_clk 0.0344f
C14737 net14 a_1375_9129# 0.00144f
C14738 net33 a_14540_3689# 0.00671f
C14739 net9 a_10864_9269# 5.31e-20
C14740 _052_ state\[2\] 0.346f
C14741 _078_ a_561_4405# 1.25e-19
C14742 net19 a_7477_10901# 2.59e-19
C14743 state\[2\] a_5055_1679# 2.38e-19
C14744 a_4349_8449# a_4393_8207# 3.69e-19
C14745 net46 _119_ 0.0655f
C14746 a_4131_8207# a_4227_8207# 0.0138f
C14747 _038_ trim_mask\[4\] 1.02e-19
C14748 net18 net9 0.0456f
C14749 en_co_clk a_4725_5487# 2.11e-19
C14750 net12 _092_ 0.00962f
C14751 clk en 0.0348f
C14752 a_448_7637# a_448_6549# 5.69e-19
C14753 net15 a_3224_2601# 0.0035f
C14754 _074_ a_5363_12559# 0.0341f
C14755 _062_ a_7800_4631# 6.61e-21
C14756 _098_ state\[2\] 0.0595f
C14757 clknet_2_3__leaf_clk cal_itt\[2\] 2.4e-19
C14758 a_10699_5487# _104_ 4.46e-22
C14759 mask\[4\] a_8673_10625# 0.00101f
C14760 a_4259_6031# a_4091_5309# 1.43e-21
C14761 _064_ a_11057_3855# 0.00344f
C14762 net37 trim_val\[0\] 0.0153f
C14763 _053_ a_11059_7356# 0.0172f
C14764 mask\[6\] _078_ 0.307f
C14765 cal_count\[1\] cal_count\[2\] 4.34e-19
C14766 a_6523_7119# VPWR 0.221f
C14767 a_5455_4943# _089_ 2.73e-19
C14768 a_7001_7669# cal_itt\[3\] 6.76e-21
C14769 a_8072_11721# _020_ 0.00129f
C14770 a_3273_4943# _097_ 3.28e-19
C14771 net16 a_14172_4943# 0.0106f
C14772 _041_ a_5691_7637# 4.56e-21
C14773 mask\[3\] a_5524_9295# 0.058f
C14774 a_5340_6031# _092_ 2.64e-19
C14775 net45 a_3302_3677# 0.00196f
C14776 _048_ _096_ 0.0551f
C14777 net44 _049_ 0.0558f
C14778 mask\[6\] a_2869_11247# 0.00286f
C14779 _115_ trim_val\[2\] 0.0012f
C14780 net45 _051_ 0.00193f
C14781 net53 a_6909_10933# 0.00258f
C14782 net43 a_8761_7983# 3.14e-20
C14783 calibrate a_1651_4703# 0.0914f
C14784 net44 a_7259_11305# 0.164f
C14785 net4 net54 1.14e-19
C14786 _107_ clk 0.0308f
C14787 net15 a_3431_10933# 8.47e-19
C14788 net45 _014_ 0.346f
C14789 net37 _126_ 0.458f
C14790 net12 cal_itt\[3\] 0.012f
C14791 clknet_2_1__leaf_clk a_5997_10927# 9.25e-19
C14792 _101_ a_1476_10217# 1.33e-21
C14793 _121_ a_3748_6281# 0.106f
C14794 a_10864_7387# a_11141_6031# 1.89e-21
C14795 a_8820_6005# a_8298_5487# 0.00682f
C14796 net24 a_3781_8207# 9.63e-20
C14797 _064_ a_10543_2455# 0.0954f
C14798 net12 a_6906_2355# 0.00143f
C14799 _107_ a_9084_4515# 0.00884f
C14800 trim_mask\[0\] trim_mask\[1\] 0.0496f
C14801 _029_ _030_ 3.04e-21
C14802 _074_ a_579_10933# 0.0207f
C14803 _065_ cal_count\[3\] 0.0151f
C14804 net43 a_3303_10217# 0.188f
C14805 _050_ _100_ 8.69e-21
C14806 a_2767_2223# VPWR 0.133f
C14807 a_11057_4105# VPWR 0.184f
C14808 a_1137_5487# VPWR 0.00632f
C14809 _123_ a_11258_8790# 0.00109f
C14810 a_12723_4943# a_12323_4703# 0.01f
C14811 a_11116_8983# a_11575_8790# 6.64e-19
C14812 _049_ clk 0.483f
C14813 _049_ en_co_clk 0.459f
C14814 _105_ clknet_2_2__leaf_clk 4.87e-20
C14815 a_2971_8457# a_3053_8457# 0.171f
C14816 mask\[6\] a_3597_10933# 0.0254f
C14817 a_7916_8041# a_8307_6575# 4.06e-20
C14818 en_co_clk a_3388_4631# 4.52e-20
C14819 a_5699_1653# clk 0.031f
C14820 a_4512_12393# a_6541_12021# 9.89e-22
C14821 a_10543_2455# a_10851_1653# 3.08e-19
C14822 net46 a_11679_4777# 0.00142f
C14823 net33 a_14335_2442# 5.32e-20
C14824 net30 a_8389_5193# 1.47e-19
C14825 clknet_0_clk _110_ 1.84e-21
C14826 net51 a_6428_7119# 6.51e-21
C14827 a_4512_11305# _019_ 2.67e-19
C14828 net19 a_6467_9845# 7.96e-22
C14829 net33 net8 1.21e-19
C14830 a_561_6031# a_1585_6031# 2.36e-20
C14831 _052_ _100_ 0.00194f
C14832 a_1651_10143# result[4] 3.24e-19
C14833 net50 a_8583_3317# 2.82e-21
C14834 clknet_2_2__leaf_clk a_7010_3311# 1.05e-20
C14835 _118_ a_9839_3615# 1.64e-20
C14836 net13 a_3947_11305# 0.00146f
C14837 _045_ ctlp[7] 0.0227f
C14838 trim[2] trim[3] 0.0486f
C14839 net28 _011_ 0.0751f
C14840 net16 a_14099_3017# 0.00983f
C14841 _009_ net12 8.32e-19
C14842 net29 clknet_2_1__leaf_clk 0.00238f
C14843 _098_ _100_ 0.048f
C14844 a_14249_8725# VPWR 0.211f
C14845 _078_ a_1763_9295# 0.00136f
C14846 a_1822_10927# VPWR 8.42e-19
C14847 net19 VPWR 1.54f
C14848 a_1467_7923# a_2143_7663# 0.0216f
C14849 net43 a_1173_7119# 0.00368f
C14850 _048_ a_5455_4943# 0.0335f
C14851 _059_ a_4725_5487# 4.7e-21
C14852 a_12148_4777# _110_ 0.00254f
C14853 a_1099_12533# _086_ 0.00109f
C14854 a_14335_7895# a_15259_7637# 1.11e-19
C14855 _046_ a_3133_11247# 2.01e-19
C14856 net42 a_7393_5193# 5.63e-19
C14857 net4 _027_ 2.02e-19
C14858 _075_ _060_ 0.245f
C14859 _122_ a_13142_8359# 0.0843f
C14860 clknet_2_1__leaf_clk _040_ 0.00956f
C14861 a_11116_8983# a_12153_8757# 4.61e-20
C14862 net41 a_2383_3689# 0.0356f
C14863 _102_ a_1476_10217# 0.00168f
C14864 clknet_2_3__leaf_clk _036_ 0.0321f
C14865 _002_ a_5691_7637# 2.85e-20
C14866 cal_itt\[0\] a_8935_6895# 0.102f
C14867 net18 trim_mask\[3\] 0.692f
C14868 _015_ a_3933_2767# 0.0131f
C14869 net48 a_13881_1653# 0.00566f
C14870 a_8949_6281# a_9043_6031# 1.26e-19
C14871 _003_ a_6428_7119# 0.158f
C14872 _058_ a_10781_3311# 2.86e-19
C14873 a_6007_7119# a_6631_7485# 9.73e-19
C14874 _114_ a_13512_1501# 2.07e-19
C14875 a_13257_1141# a_13825_1109# 0.186f
C14876 a_13091_1141# a_13607_1513# 0.107f
C14877 net14 a_1203_10927# 0.00477f
C14878 net26 a_6090_10159# 1.86e-19
C14879 net44 _008_ 0.00112f
C14880 net9 a_12153_8757# 0.0164f
C14881 clknet_2_1__leaf_clk a_3431_12021# 0.851f
C14882 a_7021_4105# a_7104_3855# 1.48e-19
C14883 net29 a_2368_9955# 1.71e-20
C14884 net4 a_4471_4007# 3.76e-21
C14885 a_561_6031# a_911_6031# 0.227f
C14886 a_14347_9480# a_14733_9545# 0.00641f
C14887 _127_ a_14377_9545# 0.0557f
C14888 a_8215_9295# _068_ 0.00323f
C14889 cal_count\[0\] _128_ 0.0184f
C14890 a_4425_6031# _090_ 2.84e-21
C14891 net47 _127_ 1.52e-20
C14892 net18 _062_ 2.2e-19
C14893 net13 a_5037_6031# 4.26e-19
C14894 clknet_2_0__leaf_clk _005_ 0.00317f
C14895 a_9296_9295# _067_ 5.17e-21
C14896 net30 a_7891_3617# 0.00119f
C14897 _104_ net41 1.28e-20
C14898 a_12323_4703# a_13059_4631# 0.0141f
C14899 a_11801_4373# _058_ 0.0126f
C14900 net46 a_9225_2197# 0.159f
C14901 _074_ a_395_9845# 0.0175f
C14902 net18 a_11508_9295# 2.78e-19
C14903 cal_itt\[1\] VPWR 0.95f
C14904 a_4512_11305# VPWR 0.309f
C14905 net43 a_2006_8751# 1.7e-19
C14906 net43 a_1019_9839# 0.0122f
C14907 _059_ _107_ 9.45e-19
C14908 _046_ a_4165_10901# 0.00305f
C14909 net12 a_6737_4719# 4.52e-19
C14910 _078_ result[0] 4.11e-20
C14911 a_2368_9955# _040_ 1.18e-21
C14912 trimb[1] trimb[4] 0.0486f
C14913 net15 clknet_2_0__leaf_clk 0.154f
C14914 net12 a_5547_5603# 1.95e-19
C14915 _065_ a_9463_8725# 1e-19
C14916 _080_ a_845_7663# 0.00379f
C14917 a_5067_2045# ctln[7] 3.69e-20
C14918 net40 _133_ 0.00147f
C14919 a_561_9845# net24 2.6e-21
C14920 net25 a_929_8757# 3.78e-20
C14921 _017_ a_4349_8449# 7.03e-19
C14922 _053_ a_11016_6691# 0.171f
C14923 net19 a_9478_4105# 3.29e-19
C14924 _076_ _034_ 1.79e-20
C14925 net34 ctln[2] 0.00136f
C14926 _053_ net3 1.05e-20
C14927 net44 a_5524_9295# 0.255f
C14928 a_13881_1653# a_13091_1141# 4.16e-20
C14929 a_12992_8751# a_13256_9117# 0.00384f
C14930 _041_ a_13016_9117# 0.00208f
C14931 net26 a_7201_9813# 0.0191f
C14932 a_395_9845# a_1279_9129# 1.16e-20
C14933 a_8473_5193# _106_ 0.00367f
C14934 a_911_10217# a_763_8757# 1.17e-20
C14935 _049_ _059_ 0.00658f
C14936 net14 a_929_8757# 0.0121f
C14937 a_3781_8207# a_4677_7882# 0.00913f
C14938 a_10137_4943# a_9839_3615# 2.4e-21
C14939 _067_ cal_count\[3\] 0.0363f
C14940 net5 _135_ 1.05e-19
C14941 a_13625_3317# a_14604_2339# 8.23e-20
C14942 a_5363_591# ctln[7] 0.362f
C14943 net49 a_13881_2741# 8.25e-19
C14944 a_4775_6031# _050_ 5.57e-20
C14945 a_5340_6031# a_5547_5603# 0.00254f
C14946 trim_mask\[0\] a_7939_3855# 3.71e-19
C14947 a_12900_7663# cal_count\[2\] 0.0129f
C14948 a_10005_6031# net30 7.08e-21
C14949 net43 a_7263_7093# 0.00135f
C14950 cal_itt\[0\] a_10239_9295# 0.00494f
C14951 net19 net27 0.0249f
C14952 net15 net13 0.00271f
C14953 a_2092_8457# a_2174_8457# 0.00477f
C14954 _001_ VPWR 1.83f
C14955 _101_ _042_ 0.0277f
C14956 _051_ a_6316_5193# 0.00417f
C14957 a_11067_4405# VPWR 0.493f
C14958 net12 a_5363_591# 0.00349f
C14959 net26 a_911_10217# 2.08e-19
C14960 cal_count\[0\] a_11895_7669# 3.14e-19
C14961 net4 a_9677_8457# 7.7e-19
C14962 net40 a_14236_8457# 0.00492f
C14963 net23 a_1129_7361# 2.72e-19
C14964 _038_ a_11491_6031# 0.00788f
C14965 a_10975_6031# a_12231_6005# 0.0436f
C14966 a_9761_1679# a_10219_2045# 0.0346f
C14967 a_5340_6031# a_5536_4399# 3.12e-19
C14968 a_6763_5193# a_7019_4407# 7.83e-20
C14969 a_929_8757# a_395_7119# 4.17e-21
C14970 a_2383_3689# a_2767_2223# 3.6e-21
C14971 trim_mask\[1\] _030_ 0.104f
C14972 a_13257_1141# a_13715_1135# 0.0346f
C14973 calibrate a_5931_4105# 0.0647f
C14974 a_13091_4943# _110_ 0.00426f
C14975 a_13625_3317# a_14193_3285# 0.186f
C14976 _068_ a_8298_5487# 2.29e-19
C14977 a_12153_8757# a_12436_9129# 0.198f
C14978 mask\[5\] net53 0.188f
C14979 a_7824_11305# a_7723_10143# 1.27e-20
C14980 net9 a_12691_2527# 3.47e-19
C14981 a_8022_7119# _051_ 4.12e-20
C14982 a_15023_1135# trim[3] 0.337f
C14983 _072_ a_7256_8029# 2.59e-19
C14984 _108_ a_9802_4007# 0.235f
C14985 net28 clknet_2_1__leaf_clk 0.242f
C14986 mask\[6\] net12 0.00824f
C14987 a_2953_9845# a_3303_10217# 0.22f
C14988 a_13715_5309# trim[4] 1.32e-19
C14989 a_2659_2601# a_3224_2601# 7.99e-20
C14990 mask\[2\] a_763_8757# 7.45e-21
C14991 _106_ a_8583_3317# 0.0015f
C14992 net16 net48 0.22f
C14993 clknet_2_2__leaf_clk a_12586_3311# 2.74e-19
C14994 _104_ a_11057_4105# 0.00732f
C14995 _039_ a_1493_5487# 6.7e-20
C14996 net52 a_1461_10357# 1.82e-19
C14997 clknet_2_3__leaf_clk a_8636_9295# 0.0138f
C14998 net30 _099_ 7.54e-20
C14999 _078_ a_1497_8725# 0.0257f
C15000 a_2689_8751# a_2143_7663# 2.2e-20
C15001 _123_ a_12344_8041# 0.0324f
C15002 net43 a_1493_5487# 1.58e-19
C15003 _065_ _095_ 0.178f
C15004 a_10188_4105# a_10055_2767# 0.00121f
C15005 trim_mask\[4\] clk 0.00945f
C15006 a_6056_8359# a_6885_8372# 5.21e-19
C15007 a_3116_12533# _046_ 0.00266f
C15008 net44 a_4036_8207# 5.91e-20
C15009 _074_ net1 0.113f
C15010 _016_ a_3521_7361# 3.37e-19
C15011 net26 mask\[2\] 7.52e-20
C15012 a_3565_7119# _049_ 2.4e-20
C15013 _091_ _092_ 0.115f
C15014 net9 a_13050_7637# 9.58e-19
C15015 a_579_12021# net43 0.311f
C15016 _011_ a_1313_11989# 7.65e-19
C15017 _065_ a_10383_7093# 0.00232f
C15018 a_9084_4515# trim_mask\[4\] 1.75e-20
C15019 a_1125_7663# a_911_7119# 4.65e-19
C15020 a_3063_591# VPWR 0.292f
C15021 net31 a_13625_3317# 9.64e-20
C15022 _118_ a_9125_4943# 1.73e-20
C15023 net19 a_8455_10383# 0.00603f
C15024 net37 net32 0.129f
C15025 a_8491_2229# a_7942_2223# 3.88e-21
C15026 _102_ _042_ 1.59e-20
C15027 a_7310_2223# a_7140_2223# 2.6e-19
C15028 a_7916_8041# VPWR 0.28f
C15029 cal_itt\[2\] a_6835_7669# 0.00131f
C15030 net19 _104_ 0.122f
C15031 net46 a_10111_1679# 0.187f
C15032 net40 _129_ 0.083f
C15033 net47 _041_ 0.611f
C15034 _128_ a_13919_8751# 0.00276f
C15035 a_9463_8725# _067_ 5.48e-19
C15036 net52 _018_ 0.19f
C15037 _062_ a_11023_5108# 9.39e-20
C15038 a_8583_3317# _033_ 0.168f
C15039 a_4165_11989# a_4209_12381# 3.69e-19
C15040 _005_ a_561_7119# 0.308f
C15041 a_3597_12021# a_4621_12393# 2.36e-20
C15042 a_13512_1501# VPWR 0.0857f
C15043 clknet_2_1__leaf_clk a_4167_11471# 8.29e-20
C15044 net14 clknet_2_0__leaf_clk 0.527f
C15045 net16 trimb[4] 3e-20
C15046 a_8749_3317# a_8298_2767# 0.0151f
C15047 a_14379_6397# _061_ 0.00275f
C15048 _135_ a_15023_6031# 1.17e-19
C15049 a_5829_9839# VPWR 0.00866f
C15050 net44 a_6891_12393# 0.155f
C15051 a_10055_2767# trim_mask\[3\] 0.0016f
C15052 a_14335_7895# a_14485_7663# 0.00899f
C15053 a_6541_12021# a_7456_12393# 0.125f
C15054 _101_ a_6909_10933# 5.02e-20
C15055 _092_ _089_ 1.2e-20
C15056 _049_ a_5694_6031# 4.02e-19
C15057 a_1844_9129# net24 0.0587f
C15058 a_2815_9447# a_2961_9545# 0.171f
C15059 a_11509_3317# a_11955_3689# 2.28e-19
C15060 _078_ ctlp[7] 5.41e-19
C15061 trim_mask\[3\] a_9926_2589# 4.97e-19
C15062 net3 a_3891_4943# 0.0657f
C15063 a_10239_9295# a_10405_9295# 0.55f
C15064 a_4443_9295# mask\[1\] 2.06e-20
C15065 _006_ net24 0.0752f
C15066 _122_ a_13557_8457# 0.0107f
C15067 _027_ a_9007_2601# 0.0336f
C15068 a_8491_2229# a_9747_2527# 0.0436f
C15069 net46 _135_ 6e-20
C15070 _107_ a_9802_4007# 0.0022f
C15071 _113_ _031_ 0.00248f
C15072 a_5496_12131# _084_ 8.19e-19
C15073 _004_ result[0] 0.00119f
C15074 net46 a_13869_1501# 0.0036f
C15075 clknet_2_0__leaf_clk a_395_7119# 0.266f
C15076 net21 clknet_2_1__leaf_clk 0.00953f
C15077 _085_ net26 1.3e-20
C15078 a_8307_6575# _062_ 2.48e-19
C15079 net52 mask\[1\] 0.114f
C15080 _064_ a_10699_3311# 0.109f
C15081 net43 net53 0.0135f
C15082 a_11394_9509# VPWR 0.231f
C15083 a_4259_6031# net30 2.09e-19
C15084 _108_ _107_ 0.412f
C15085 a_1313_10901# a_1660_11305# 0.0512f
C15086 a_745_10933# net52 0.00214f
C15087 net37 VPWR 0.557f
C15088 net34 a_14335_2442# 4.93e-19
C15089 a_1375_9129# VPWR 4.66e-19
C15090 net34 net8 0.0332f
C15091 net19 a_8381_9295# 0.0168f
C15092 a_3123_3615# clk 5.68e-19
C15093 en_co_clk a_3123_3615# 3.25e-21
C15094 _087_ state\[2\] 0.00261f
C15095 a_7442_7119# VPWR 1.48e-19
C15096 _060_ a_4658_3427# 4.96e-19
C15097 _078_ _021_ 5.51e-21
C15098 a_11233_4405# a_11679_4777# 2.28e-19
C15099 _093_ net1 0.00112f
C15100 state\[2\] a_6519_3829# 2.59e-20
C15101 net45 net22 0.156f
C15102 mask\[7\] a_3511_11471# 5.21e-21
C15103 mask\[3\] a_3303_10217# 2.36e-20
C15104 a_10699_3311# a_10851_1653# 1.03e-20
C15105 clknet_2_2__leaf_clk a_14347_4917# 2.36e-21
C15106 _051_ a_6210_4989# 0.116f
C15107 net33 a_13459_3317# 2.82e-20
C15108 a_4209_12381# VPWR 3.71e-20
C15109 a_10543_2455# a_10689_2223# 0.171f
C15110 a_11601_2229# a_12047_2601# 2.28e-19
C15111 _049_ _108_ 2.47e-20
C15112 net45 a_2921_2589# 0.00316f
C15113 _099_ state\[2\] 1.26e-19
C15114 net16 a_14281_1513# 6.83e-21
C15115 a_13193_6031# VPWR 3.57e-19
C15116 calibrate a_7527_4631# 2.51e-19
C15117 _050_ a_3933_2767# 1.97e-20
C15118 a_11116_8983# VPWR 0.105f
C15119 mask\[5\] a_6007_9839# 9e-21
C15120 _081_ a_1476_7119# 3.75e-21
C15121 a_10699_5487# a_11057_4105# 4.61e-21
C15122 a_11067_4405# _104_ 7.3e-20
C15123 clknet_2_2__leaf_clk _119_ 0.358f
C15124 _081_ mask\[0\] 1.69e-19
C15125 _099_ state\[0\] 3.09e-20
C15126 net28 a_4866_12381# 0.002f
C15127 mask\[4\] a_6099_10633# 0.0611f
C15128 a_1461_10357# a_1679_10633# 0.0821f
C15129 clknet_2_3__leaf_clk net4 0.0256f
C15130 net19 _110_ 0.0477f
C15131 calibrate state\[1\] 0.00217f
C15132 net16 trim[0] 3.49e-20
C15133 net46 a_13519_4007# 1.89e-20
C15134 clknet_2_0__leaf_clk a_2659_2601# 0.0306f
C15135 a_4995_7119# VPWR 0.305f
C15136 net9 VPWR 1.25f
C15137 clknet_2_1__leaf_clk _020_ 0.349f
C15138 net14 a_1203_12015# 0.00311f
C15139 a_4043_7093# net30 1.19e-19
C15140 trim_mask\[2\] a_14471_591# 3e-19
C15141 _092_ _048_ 0.273f
C15142 net19 clknet_0_clk 0.0411f
C15143 net44 a_8949_9537# 2.45e-19
C15144 net33 _109_ 9.17e-21
C15145 _067_ a_10383_7093# 0.013f
C15146 a_5547_5603# a_5726_5807# 0.00698f
C15147 trim_mask\[0\] _066_ 0.0715f
C15148 a_13625_3317# a_14083_3311# 0.0346f
C15149 clknet_2_1__leaf_clk a_1313_11989# 4.07e-20
C15150 net9 a_12218_6397# 9.87e-20
C15151 net15 a_2948_3689# 0.00642f
C15152 _086_ a_1137_11721# 0.00114f
C15153 _065_ calibrate 3.98e-20
C15154 _053_ net54 1.84e-19
C15155 a_12691_2527# a_13415_2442# 0.0112f
C15156 mask\[0\] a_455_5747# 2.42e-21
C15157 a_13415_2442# _114_ 0.00163f
C15158 a_9747_2527# a_10195_1354# 1.37e-19
C15159 net40 a_14318_8457# 2.58e-19
C15160 _107_ a_9004_3677# 5.02e-19
C15161 a_6541_12021# a_6743_10933# 2.78e-21
C15162 a_6375_12021# a_6909_10933# 1.15e-19
C15163 a_7824_11305# _042_ 1.03e-19
C15164 _049_ a_4725_5487# 7.62e-20
C15165 net40 a_12323_4703# 5.37e-20
C15166 _122_ a_10975_6031# 5.3e-19
C15167 net33 trim[2] 0.11f
C15168 _125_ a_12992_8751# 1.43e-20
C15169 clknet_2_3__leaf_clk a_14172_4943# 1.88e-21
C15170 net16 _130_ 0.0061f
C15171 net15 a_4167_6575# 5.67e-19
C15172 net24 _017_ 0.00128f
C15173 _064_ _027_ 0.00142f
C15174 _101_ a_4959_9295# 0.00139f
C15175 a_8949_6031# VPWR 2.27e-19
C15176 net16 a_14335_4020# 0.00604f
C15177 net46 a_14604_3017# 0.00178f
C15178 clknet_0_clk cal_itt\[1\] 0.0151f
C15179 _062_ a_7897_6913# 6.54e-20
C15180 _123_ _133_ 0.143f
C15181 _012_ a_455_3571# 9.78e-19
C15182 a_395_4405# a_995_3530# 1.03e-21
C15183 _074_ a_5915_11721# 3.15e-19
C15184 _063_ a_10975_6031# 2.69e-20
C15185 cal_itt\[3\] _048_ 2.38e-19
C15186 net14 a_561_7119# 0.0121f
C15187 trim_mask\[2\] a_13825_1109# 1.47e-20
C15188 _078_ a_4655_10071# 4.2e-21
C15189 a_816_4765# cal 0.00123f
C15190 _090_ a_3273_4943# 0.139f
C15191 _087_ _100_ 0.0124f
C15192 a_14281_4943# net49 3.38e-20
C15193 net37 a_14807_8359# 0.00414f
C15194 clknet_2_3__leaf_clk a_11479_9117# 3.34e-19
C15195 a_4165_11989# a_3431_10933# 4.52e-22
C15196 trim_mask\[0\] a_7571_4943# 4.51e-19
C15197 _100_ a_6519_3829# 0.0112f
C15198 _088_ a_5087_3855# 6.68e-21
C15199 a_3431_12021# _009_ 1.71e-21
C15200 a_9747_2527# _032_ 4.72e-19
C15201 a_10569_1109# a_10752_565# 8.07e-20
C15202 a_9572_2601# a_9595_1679# 8.91e-19
C15203 a_6909_10933# a_7986_10927# 1.46e-19
C15204 a_7477_10901# a_7367_10927# 0.0977f
C15205 _049_ _107_ 0.0962f
C15206 a_9471_9269# cal_itt\[0\] 0.102f
C15207 a_8636_9295# a_8827_9295# 4.61e-19
C15208 a_448_11445# VPWR 0.329f
C15209 net43 _071_ 0.00629f
C15210 mask\[4\] a_5423_9011# 1.07e-21
C15211 _099_ _100_ 0.0406f
C15212 a_10975_4105# _025_ 2.61e-20
C15213 a_455_5747# _079_ 0.00107f
C15214 _041_ _072_ 5.23e-20
C15215 a_10188_4105# VPWR 0.16f
C15216 a_7190_3855# _054_ 0.119f
C15217 a_395_7119# a_561_7119# 0.864f
C15218 net12 _073_ 0.00478f
C15219 net21 a_4866_12381# 1.36e-19
C15220 a_12436_9129# VPWR 0.285f
C15221 _125_ a_15111_9295# 0.00172f
C15222 _123_ a_14236_8457# 6.19e-21
C15223 a_1203_10927# VPWR 0.145f
C15224 a_745_10933# a_1679_10633# 3.25e-19
C15225 a_3224_2601# VPWR 0.277f
C15226 trim_mask\[2\] a_13307_1707# 0.0537f
C15227 _068_ _041_ 0.0507f
C15228 a_11067_4405# _110_ 1.76e-20
C15229 clknet_2_2__leaf_clk a_7617_2589# 8.94e-20
C15230 _040_ a_4805_8207# 0.00103f
C15231 mask\[5\] _101_ 0.382f
C15232 a_13050_7637# a_13470_7663# 0.144f
C15233 _124_ a_11059_7356# 8.48e-20
C15234 net15 a_3461_5193# 9.27e-19
C15235 net40 a_14379_6397# 0.00448f
C15236 _053_ a_7019_4407# 0.0101f
C15237 _049_ a_3388_4631# 2.74e-19
C15238 clknet_2_3__leaf_clk a_10586_7371# 1.68e-19
C15239 _128_ cal_count\[2\] 0.00309f
C15240 a_6885_8372# _070_ 5.08e-20
C15241 net45 a_4871_6031# 3.56e-20
C15242 mask\[6\] a_5997_10927# 0.0116f
C15243 a_1660_11305# result[5] 1.11e-19
C15244 clknet_2_1__leaf_clk a_2143_7663# 0.00291f
C15245 a_4443_9295# _041_ 7.15e-20
C15246 a_4609_1679# a_5067_2045# 0.0276f
C15247 a_4959_1679# a_5524_1679# 7.99e-20
C15248 a_6173_7119# a_7088_7119# 0.125f
C15249 _074_ a_911_10217# 0.0136f
C15250 net53 a_2953_9845# 7.04e-20
C15251 _000_ _076_ 1.78e-20
C15252 _078_ a_1129_7361# 3.77e-19
C15253 a_6909_10933# a_7824_11305# 0.125f
C15254 a_9195_10357# a_8992_9955# 0.00781f
C15255 net30 a_9503_4399# 0.0977f
C15256 net18 a_9020_10383# 2.68e-19
C15257 net2 a_13512_4943# 1.91e-19
C15258 net52 _041_ 0.00218f
C15259 _035_ a_10798_9295# 3.33e-19
C15260 a_4863_4917# VPWR 0.254f
C15261 a_8215_9295# _067_ 1.31e-22
C15262 a_14249_8725# a_14467_8751# 0.0821f
C15263 a_1095_12393# _078_ 6.41e-19
C15264 net40 _038_ 2.03e-19
C15265 trim_mask\[3\] VPWR 0.53f
C15266 a_4709_2773# a_4901_2773# 1.81e-19
C15267 a_10699_5487# a_11067_4405# 8.93e-19
C15268 a_1129_6273# a_911_4777# 5.13e-21
C15269 a_911_6031# a_1129_4373# 5.13e-21
C15270 _136_ _109_ 0.00114f
C15271 _024_ a_12323_4703# 2.09e-19
C15272 a_11067_4405# a_12148_4777# 0.102f
C15273 _125_ a_14422_7093# 1.04e-19
C15274 a_3431_10933# VPWR 0.43f
C15275 net43 a_1541_9117# 0.00378f
C15276 a_10005_6031# _118_ 3.89e-19
C15277 net2 a_14377_7983# 0.00117f
C15278 clknet_2_2__leaf_clk a_9225_2197# 0.0325f
C15279 net50 a_9572_2601# 1.17e-20
C15280 a_10689_2543# VPWR 2.07e-19
C15281 _078_ a_1638_9839# 1.98e-19
C15282 a_929_8757# VPWR 0.291f
C15283 _062_ VPWR 3.68f
C15284 a_561_4405# a_816_4765# 0.0642f
C15285 net30 a_7942_2223# 5.29e-20
C15286 net22 a_2857_5461# 1.84e-20
C15287 a_1651_10143# a_1497_8725# 3.87e-22
C15288 mask\[2\] a_4858_8573# 1.03e-21
C15289 a_9802_4007# trim_mask\[4\] 0.0227f
C15290 _080_ a_1211_7983# 0.00151f
C15291 a_1467_7923# _005_ 4.32e-19
C15292 _012_ a_1129_4373# 8.16e-19
C15293 a_10138_5807# VPWR 2.07e-19
C15294 a_10787_1135# net10 4.27e-19
C15295 a_4425_6031# a_4883_6397# 0.0346f
C15296 a_448_6549# a_455_5747# 7.06e-19
C15297 _057_ a_14931_591# 0.206f
C15298 _094_ a_5037_6031# 0.00271f
C15299 cal_count\[0\] net40 0.0315f
C15300 _048_ a_6737_4719# 0.0482f
C15301 net29 mask\[6\] 6.37e-19
C15302 net28 _009_ 8.18e-21
C15303 a_13881_1653# a_14184_1679# 0.00138f
C15304 _042_ a_5067_9661# 2.18e-20
C15305 net46 a_9839_3615# 0.319f
C15306 _123_ _129_ 8.37e-20
C15307 a_4308_4917# a_4091_5309# 0.267f
C15308 net43 a_4621_12393# 2.95e-19
C15309 a_5547_5603# _048_ 2.7e-20
C15310 net47 a_10747_8970# 0.0126f
C15311 net33 a_15023_1135# 0.00131f
C15312 _103_ _106_ 0.00163f
C15313 _108_ trim_mask\[4\] 0.183f
C15314 _125_ _132_ 0.00249f
C15315 net27 a_448_11445# 0.18f
C15316 _065_ mask\[1\] 0.00925f
C15317 net33 a_14655_4399# 0.00559f
C15318 _074_ mask\[2\] 0.00154f
C15319 net51 _051_ 3.7e-20
C15320 a_10990_7485# a_11369_7119# 3.16e-19
C15321 a_9195_10357# a_9374_10383# 0.0074f
C15322 a_9020_10383# a_9129_10383# 0.00742f
C15323 clknet_0_clk a_7916_8041# 1.24e-19
C15324 net13 a_4959_1679# 0.0122f
C15325 net9 _104_ 3.84e-19
C15326 net33 _125_ 0.401f
C15327 _048_ a_9003_3829# 0.00276f
C15328 a_9195_3689# VPWR 5.1e-19
C15329 net46 a_9734_2223# 8.41e-20
C15330 a_11895_7669# cal_count\[2\] 0.00358f
C15331 net12 _021_ 7.98e-19
C15332 _110_ a_13512_1501# 1.14e-20
C15333 mask\[1\] net23 0.958f
C15334 a_13415_2442# VPWR 0.281f
C15335 a_7367_10927# VPWR 0.144f
C15336 mask\[4\] a_4871_8181# 7.02e-20
C15337 net43 a_5363_7369# 0.00135f
C15338 a_9471_9269# a_10405_9295# 1.98e-19
C15339 _072_ _002_ 0.0998f
C15340 net33 trimb[0] 0.00141f
C15341 a_8992_9955# a_8949_9537# 5.23e-19
C15342 _048_ a_5536_4399# 0.154f
C15343 state\[1\] _015_ 0.0493f
C15344 trim_mask\[4\] a_10655_2932# 2.45e-20
C15345 a_6198_8534# VPWR 0.00215f
C15346 clknet_2_1__leaf_clk _077_ 2.07e-20
C15347 en_co_clk _061_ 0.0379f
C15348 a_3597_12021# a_4512_12393# 0.125f
C15349 a_3431_12021# mask\[6\] 4.14e-19
C15350 net30 _097_ 4.53e-21
C15351 _068_ _002_ 6.92e-19
C15352 a_12992_8751# a_13142_8359# 0.00155f
C15353 net26 a_4609_9295# 2.09e-20
C15354 _032_ a_10676_1679# 1.92e-19
C15355 a_4775_6031# _099_ 1.53e-21
C15356 net18 _037_ 1.21e-20
C15357 a_13607_1513# _057_ 1.22e-19
C15358 calibrate _013_ 0.0224f
C15359 net21 a_6927_12559# 4.43e-21
C15360 a_5363_12559# net20 6.94e-19
C15361 _045_ a_6191_12559# 0.197f
C15362 _067_ a_8298_5487# 0.00377f
C15363 net43 _101_ 0.139f
C15364 _037_ a_10820_7485# 8.96e-21
C15365 a_6743_10933# a_7723_10143# 2.45e-20
C15366 _065_ _015_ 2.22e-19
C15367 net46 a_9207_3311# 0.0122f
C15368 net15 _094_ 0.00573f
C15369 a_6375_12021# mask\[5\] 1.04e-19
C15370 _128_ cal_count\[1\] 0.18f
C15371 a_7001_7669# a_8078_7663# 1.46e-19
C15372 a_13470_7663# VPWR 0.181f
C15373 _034_ a_5515_6005# 7.08e-20
C15374 _081_ a_1229_8457# 7.96e-20
C15375 net46 a_13393_1707# 3.61e-19
C15376 _074_ a_1000_11293# 0.00612f
C15377 _023_ a_1461_10357# 0.114f
C15378 a_1579_5807# a_1493_5487# 2.42e-19
C15379 a_10005_6031# a_10137_4943# 3.92e-20
C15380 net52 _002_ 2.55e-20
C15381 clknet_2_3__leaf_clk _000_ 0.0294f
C15382 a_3817_4697# VPWR 0.224f
C15383 net27 a_3431_10933# 1.97e-20
C15384 net37 _110_ 5.19e-20
C15385 a_5524_1679# VPWR 0.309f
C15386 net13 _019_ 0.105f
C15387 a_7571_4943# a_8307_4943# 3.51e-19
C15388 net47 a_11369_7119# 9.54e-19
C15389 _038_ _024_ 0.00259f
C15390 _085_ _074_ 0.0914f
C15391 a_6375_12021# a_6999_12015# 9.73e-19
C15392 a_7999_11231# VPWR 0.371f
C15393 clknet_2_2__leaf_clk a_11292_1251# 3.17e-20
C15394 net55 a_4815_3031# 1.35e-20
C15395 mask\[1\] a_2225_7663# 0.0105f
C15396 trim_mask\[4\] a_9004_3677# 0.025f
C15397 a_9664_3689# a_10699_3311# 3.7e-19
C15398 trim_mask\[0\] _058_ 0.142f
C15399 a_3123_3615# a_3399_2527# 1.13e-19
C15400 net53 mask\[3\] 0.00181f
C15401 a_8745_6895# VPWR 0.00182f
C15402 mask\[1\] _016_ 0.00155f
C15403 net16 trim[4] 4.7e-20
C15404 clknet_2_0__leaf_clk VPWR 7.25f
C15405 net21 _009_ 5.24e-21
C15406 net14 a_1585_4777# 2.37e-19
C15407 net44 a_7263_7093# 0.341f
C15408 _104_ a_10188_4105# 2.89e-19
C15409 _107_ trim_mask\[4\] 0.0049f
C15410 net43 _086_ 0.011f
C15411 net9 a_12678_2223# 1.44e-19
C15412 _026_ a_12047_2601# 7.96e-19
C15413 net13 a_5878_1679# 1.57e-19
C15414 _083_ a_6090_10159# 0.003f
C15415 _048_ a_8485_4943# 3.16e-19
C15416 a_15023_9839# trimb[4] 2.97e-20
C15417 _088_ a_6822_4105# 0.0156f
C15418 net15 a_2787_7119# 0.0217f
C15419 net4 a_6835_7669# 3.13e-22
C15420 a_4687_12319# VPWR 0.374f
C15421 clknet_2_2__leaf_clk a_10111_1679# 1.7e-19
C15422 net11 VPWR 0.572f
C15423 a_3597_12021# _046_ 9.45e-19
C15424 net16 a_14471_12559# 0.174f
C15425 mask\[1\] a_4696_8207# 0.0542f
C15426 net9 _110_ 0.138f
C15427 net43 _102_ 0.00624f
C15428 clknet_0_clk a_4995_7119# 1.96e-21
C15429 _081_ a_1125_7663# 1.76e-20
C15430 a_14335_7895# _133_ 0.148f
C15431 net33 trim[1] 0.00648f
C15432 net52 a_3615_8207# 0.00489f
C15433 _049_ trim_mask\[4\] 0.161f
C15434 net28 mask\[6\] 0.365f
C15435 net51 a_7613_8029# 1.55e-19
C15436 net34 trim[2] 0.0157f
C15437 _090_ a_4091_5309# 4.94e-20
C15438 net13 VPWR 1.38f
C15439 a_1651_6005# result[0] 1.48e-19
C15440 a_7010_3311# a_7524_2223# 9.66e-21
C15441 a_4259_6031# a_4775_6031# 0.111f
C15442 a_4425_6031# a_4993_6273# 0.186f
C15443 a_7263_7093# clk 0.0142f
C15444 a_2288_3677# a_2479_3689# 4.61e-19
C15445 net9 a_12778_3677# 2.57e-19
C15446 a_10699_3311# a_10781_3631# 0.00393f
C15447 net14 a_1467_7923# 0.00189f
C15448 mask\[4\] clknet_2_3__leaf_clk 1.27e-19
C15449 net46 a_14526_4943# 0.00196f
C15450 a_13919_8751# net40 2.09e-19
C15451 _104_ trim_mask\[3\] 0.257f
C15452 _052_ a_5931_4105# 3.29e-20
C15453 mask\[0\] a_395_4405# 1.54e-19
C15454 _019_ a_4864_9295# 0.159f
C15455 a_395_4405# valid 0.0101f
C15456 net49 a_14702_3311# 1.1e-19
C15457 a_10975_6031# a_13111_6031# 1.01e-20
C15458 a_14604_2339# a_14471_591# 8.9e-21
C15459 _083_ a_7201_9813# 1.99e-20
C15460 _101_ a_2857_7637# 0.0272f
C15461 a_14972_5193# a_15054_5193# 0.00477f
C15462 a_14172_4943# _047_ 1.66e-19
C15463 clknet_2_3__leaf_clk _064_ 0.211f
C15464 _051_ a_7223_2465# 0.0011f
C15465 net49 a_13693_3883# 2.9e-19
C15466 mask\[5\] a_7824_11305# 0.00427f
C15467 net15 a_3208_10205# 0.00623f
C15468 net17 _036_ 0.00164f
C15469 net15 a_2689_8751# 1.13e-20
C15470 net20 ctlp[6] 0.0904f
C15471 _043_ _042_ 0.019f
C15472 a_5081_4943# a_5087_3855# 8.79e-20
C15473 _103_ _054_ 5.3e-21
C15474 _098_ a_5931_4105# 4.93e-19
C15475 trim_val\[0\] a_13880_3677# 5.91e-20
C15476 net9 a_12148_4777# 0.00184f
C15477 _104_ a_10689_2543# 0.00178f
C15478 a_2033_3317# cal 2.27e-19
C15479 clknet_2_1__leaf_clk a_6173_7119# 1.45e-19
C15480 cal_itt\[0\] _069_ 0.257f
C15481 _062_ _104_ 4.39e-20
C15482 a_11583_4777# a_11067_3017# 1.14e-20
C15483 _093_ a_2143_2229# 6.21e-22
C15484 a_10207_1679# VPWR 7.26e-19
C15485 _009_ _020_ 1.89e-20
C15486 net43 _022_ 0.00451f
C15487 net55 a_5087_3855# 0.0294f
C15488 _078_ calibrate 2.42e-20
C15489 cal_itt\[0\] a_8022_7119# 0.0265f
C15490 _077_ a_6485_8181# 4.91e-20
C15491 a_5535_8181# net51 0.00296f
C15492 _045_ a_6796_12381# 2.21e-19
C15493 net27 a_7999_11231# 0.00397f
C15494 _023_ a_745_10933# 0.259f
C15495 a_579_10933# a_1313_10901# 0.0701f
C15496 a_13869_4943# _058_ 4.09e-19
C15497 trim_val\[0\] a_13697_4373# 0.189f
C15498 a_14236_8457# a_14335_7895# 4.35e-19
C15499 a_4576_3427# a_4658_3427# 0.00477f
C15500 a_7715_3285# a_7843_3677# 0.00476f
C15501 a_3748_6281# net30 1.63e-19
C15502 _097_ state\[0\] 4.23e-21
C15503 trim_val\[4\] _025_ 1.11e-20
C15504 a_1467_7923# a_395_7119# 0.00358f
C15505 a_9664_3689# _027_ 1.01e-21
C15506 _033_ a_9572_2601# 5.66e-20
C15507 _051_ a_9099_3689# 4.44e-21
C15508 _108_ a_12723_4943# 0.0365f
C15509 _036_ a_12061_7669# 1.63e-19
C15510 a_12153_8757# _037_ 2.07e-20
C15511 net19 cal_itt\[1\] 0.215f
C15512 _008_ a_5524_9295# 0.00155f
C15513 mask\[6\] a_4167_11471# 2.6e-19
C15514 a_4165_10901# a_4621_11305# 4.2e-19
C15515 a_3947_11305# a_4209_11293# 0.00171f
C15516 _065_ _041_ 0.204f
C15517 _104_ a_9195_3689# 0.00118f
C15518 a_1203_12015# VPWR 0.143f
C15519 _027_ a_10689_2223# 0.00475f
C15520 trim_mask\[0\] a_13607_4943# 0.00719f
C15521 net16 _057_ 1.4e-20
C15522 _108_ _056_ 0.00425f
C15523 _040_ a_3317_8207# 0.00356f
C15524 a_15023_5487# comp 3.98e-20
C15525 net26 a_6181_10633# 6.35e-20
C15526 _079_ a_395_4405# 1.26e-20
C15527 clknet_2_3__leaf_clk _053_ 1.13f
C15528 _110_ a_10188_4105# 3.09e-19
C15529 a_11067_4405# a_11057_4105# 3.33e-19
C15530 a_4687_12319# net27 1.17e-20
C15531 a_4864_9295# VPWR 0.0794f
C15532 _088_ a_7677_4759# 5.81e-20
C15533 a_11204_7485# _038_ 2.17e-20
C15534 a_11599_6397# _136_ 0.00138f
C15535 a_7631_12319# a_7477_10901# 9.96e-21
C15536 _101_ a_2953_9845# 0.493f
C15537 a_7456_12393# a_6909_10933# 1.89e-19
C15538 a_7351_8041# a_7088_7119# 5.01e-19
C15539 a_3388_4631# a_3123_3615# 1.98e-19
C15540 _078_ a_1461_10357# 0.011f
C15541 trim_mask\[2\] a_12625_2601# 1.33e-19
C15542 a_4959_9295# a_5067_9661# 0.0572f
C15543 clknet_2_2__leaf_clk a_13519_4007# 0.0016f
C15544 net21 mask\[6\] 0.00186f
C15545 _099_ a_3933_2767# 4.06e-21
C15546 _028_ a_6927_3311# 9.92e-19
C15547 net27 net13 0.074f
C15548 net47 a_8839_9661# 0.0129f
C15549 a_11244_9661# cal_count\[0\] 0.00966f
C15550 net12 a_6566_5193# 0.00306f
C15551 net40 en_co_clk 0.084f
C15552 trim_val\[1\] a_14686_3017# 0.00172f
C15553 _094_ a_5449_6031# 3.29e-19
C15554 net12 _095_ 6.2e-21
C15555 a_7351_8041# _063_ 1.33e-20
C15556 net44 net53 0.123f
C15557 a_561_9845# a_448_9269# 2.18e-19
C15558 _123_ a_13100_8751# 0.00177f
C15559 net45 a_2877_2197# 0.166f
C15560 _129_ a_14335_7895# 0.0732f
C15561 a_12323_4703# trim_mask\[1\] 5.11e-23
C15562 a_561_7119# VPWR 0.605f
C15563 net52 a_3249_9295# 0.00475f
C15564 a_14471_12559# trimb[3] 6.54e-19
C15565 _128_ a_12900_7663# 0.0117f
C15566 _107_ a_7320_3631# 2.35e-19
C15567 _058_ _030_ 0.00101f
C15568 a_6743_10933# _042_ 7.87e-20
C15569 a_7999_11231# a_8455_10383# 3.32e-19
C15570 a_2787_7119# a_3399_7119# 3.82e-19
C15571 a_2953_7119# a_4030_7485# 1.46e-19
C15572 clknet_2_0__leaf_clk a_2383_3689# 2.38e-19
C15573 net19 _001_ 2.07e-19
C15574 _048_ a_4266_4943# 0.00275f
C15575 _110_ trim_mask\[3\] 0.121f
C15576 a_911_4777# a_995_3530# 2.16e-20
C15577 _125_ a_11987_8757# 2.29e-20
C15578 _051_ _088_ 2.97e-19
C15579 _065_ a_10781_5487# 3.33e-21
C15580 clknet_0_clk a_4863_4917# 8.61e-20
C15581 clknet_2_1__leaf_clk a_3852_11293# 0.00239f
C15582 a_1313_10901# a_395_9845# 3.13e-20
C15583 net35 _108_ 0.00122f
C15584 _108_ a_13059_4631# 9.5e-19
C15585 net15 _096_ 0.00182f
C15586 _122_ a_13164_8029# 6.42e-19
C15587 _051_ a_7262_5461# 0.114f
C15588 net34 a_15023_1135# 0.22f
C15589 _062_ _110_ 3.13e-19
C15590 net9 a_13091_4943# 4.94e-19
C15591 _050_ a_7527_4631# 0.00104f
C15592 cal_count\[0\] _123_ 0.293f
C15593 net34 a_14655_4399# 3.82e-22
C15594 clknet_0_clk _062_ 0.142f
C15595 _078_ _018_ 0.00646f
C15596 _120_ net55 2.09e-21
C15597 net25 a_3208_10205# 8.78e-21
C15598 a_14788_7369# VPWR 0.156f
C15599 _090_ a_4886_4399# 0.00148f
C15600 _049_ a_7320_3631# 0.00435f
C15601 net34 _125_ 0.0132f
C15602 net24 _080_ 0.0117f
C15603 a_395_7119# a_2787_7119# 1.75e-19
C15604 net49 a_14237_3677# 6.71e-19
C15605 _048_ _105_ 0.237f
C15606 a_13607_4943# a_13869_4943# 0.00171f
C15607 a_13825_5185# trim_val\[0\] 0.00308f
C15608 _050_ state\[1\] 4.82e-20
C15609 a_14172_4943# a_14334_5309# 0.00645f
C15610 _093_ a_5087_3855# 3.26e-20
C15611 a_8491_2229# a_9595_1679# 9.7e-19
C15612 net18 _122_ 0.155f
C15613 _051_ a_6519_4631# 2.03e-20
C15614 a_4091_4943# VPWR 6.94e-20
C15615 _001_ cal_itt\[1\] 0.00103f
C15616 _021_ a_5997_10927# 0.0018f
C15617 net48 a_14099_1929# 0.0911f
C15618 _000_ a_8827_9295# 9.32e-19
C15619 net34 trimb[0] 0.0659f
C15620 a_6885_8372# net2 0.0326f
C15621 _052_ a_7527_4631# 2.19e-20
C15622 _065_ _002_ 0.0293f
C15623 _118_ a_9503_4399# 0.0112f
C15624 a_3388_4631# a_3530_4765# 0.00783f
C15625 clknet_2_1__leaf_clk a_3947_11305# 0.00214f
C15626 _092_ a_10975_6031# 0.00324f
C15627 a_4239_8573# VPWR 0.134f
C15628 trim_mask\[0\] a_11488_4765# 7.47e-20
C15629 clknet_2_1__leaf_clk a_7109_11989# 4.98e-19
C15630 net43 a_4512_12393# 0.216f
C15631 net18 _063_ 2.7e-19
C15632 _059_ a_6737_3855# 8.65e-21
C15633 _048_ a_7010_3311# 4.7e-21
C15634 _065_ _050_ 0.0226f
C15635 _110_ a_13415_2442# 0.0044f
C15636 _091_ cal_count\[3\] 2.04e-19
C15637 _098_ a_7527_4631# 7.16e-19
C15638 clkc trim[4] 0.0371f
C15639 a_455_8181# result[3] 0.00182f
C15640 _041_ _067_ 2.26e-20
C15641 a_11895_7669# a_12900_7663# 0.178f
C15642 _037_ a_13050_7637# 0.00151f
C15643 net4 a_2143_2229# 0.0101f
C15644 _078_ mask\[1\] 0.975f
C15645 trim_mask\[0\] _113_ 3.43e-19
C15646 _012_ _097_ 7.01e-20
C15647 _073_ _048_ 7.12e-19
C15648 net47 a_10877_7983# 3.32e-19
C15649 _074_ a_1000_12381# 1.14e-19
C15650 _078_ a_745_10933# 0.0225f
C15651 a_579_10933# result[5] 0.00691f
C15652 a_7631_12319# VPWR 0.392f
C15653 net2 a_11141_6031# 9.68e-20
C15654 _022_ a_2953_9845# 7.1e-19
C15655 a_6007_7119# a_6173_7119# 0.906f
C15656 a_2953_7119# a_3977_7119# 2.36e-20
C15657 _104_ a_10207_1679# 7.42e-20
C15658 a_14099_1929# a_13091_1141# 2.64e-20
C15659 _004_ calibrate 2.09e-19
C15660 a_9719_1473# a_10195_1354# 0.0157f
C15661 a_1651_4703# _099_ 3e-19
C15662 a_1476_4777# a_2865_4460# 5.06e-20
C15663 a_6743_10933# a_6909_10933# 0.901f
C15664 _074_ a_4609_9295# 0.0117f
C15665 _042_ a_3868_10217# 0.016f
C15666 a_2948_3689# VPWR 0.314f
C15667 a_12992_8751# a_12916_8751# 0.00212f
C15668 a_12520_7637# cal_count\[3\] 8.19e-20
C15669 _101_ mask\[3\] 0.341f
C15670 clknet_2_0__leaf_clk a_1007_4777# 1.44e-19
C15671 a_14981_4020# a_15023_2223# 2.14e-20
C15672 a_1173_10205# result[4] 1.99e-19
C15673 net4 a_4815_3031# 0.0534f
C15674 _065_ a_3615_8207# 1.76e-20
C15675 net40 cal_count\[2\] 0.00976f
C15676 _101_ a_6741_7361# 1.05e-20
C15677 _118_ a_9747_2527# 3.87e-22
C15678 a_7916_8041# cal_itt\[1\] 3.79e-21
C15679 clknet_2_2__leaf_clk a_7184_2339# 0.00247f
C15680 _071_ a_9459_7895# 1.22e-20
C15681 a_9020_10383# VPWR 0.28f
C15682 _078_ a_1387_8751# 0.00281f
C15683 a_4167_6575# VPWR 0.224f
C15684 net44 _071_ 2.38e-20
C15685 net23 a_3615_8207# 1.89e-20
C15686 _108_ a_13257_4943# 0.397f
C15687 net45 a_1476_6031# 0.237f
C15688 ctlp[3] ctlp[2] 0.00303f
C15689 _122_ a_11575_8790# 2.48e-19
C15690 net45 a_5177_1921# 0.166f
C15691 cal_count\[0\] a_13142_8725# 0.065f
C15692 a_8022_7119# a_8949_6281# 6.87e-20
C15693 _067_ a_10781_5487# 0.00139f
C15694 _032_ a_9719_1473# 0.0323f
C15695 a_9595_1679# a_10195_1354# 2.48e-20
C15696 clknet_2_0__leaf_clk clknet_0_clk 0.825f
C15697 a_14807_8359# a_14788_7369# 1.56e-20
C15698 net43 _046_ 0.0132f
C15699 net53 a_4801_9839# 0.00625f
C15700 clknet_2_1__leaf_clk _005_ 1.3e-21
C15701 _126_ _122_ 1.19e-19
C15702 net41 a_3224_2601# 3.16e-21
C15703 _082_ a_763_8757# 5.57e-20
C15704 _048_ a_3365_4943# 0.00302f
C15705 net34 trim[1] 0.0403f
C15706 net16 a_13625_3317# 0.0161f
C15707 clknet_2_2__leaf_clk a_9839_3615# 0.00137f
C15708 a_1844_9129# a_1476_7119# 2.99e-21
C15709 net12 calibrate 0.0079f
C15710 a_1844_9129# mask\[0\] 3.55e-19
C15711 _028_ VPWR 0.442f
C15712 _110_ net11 2.59e-19
C15713 net47 a_8563_10749# 0.0122f
C15714 net15 clknet_2_1__leaf_clk 1.21f
C15715 net14 _011_ 0.00251f
C15716 a_14172_4943# net49 2.02e-19
C15717 _071_ clk 6.42e-20
C15718 net4 a_9443_6059# 0.012f
C15719 _071_ en_co_clk 0.125f
C15720 net42 _106_ 2.06e-19
C15721 a_7456_12393# mask\[5\] 2.34e-20
C15722 a_3751_4765# VPWR 1.95e-19
C15723 a_2313_6183# _094_ 5.3e-20
C15724 trim_val\[1\] a_13257_1141# 5.84e-22
C15725 trim_val\[3\] net10 5.28e-22
C15726 _060_ a_4617_4105# 0.0101f
C15727 a_10781_5487# clknet_2_2__leaf_clk 5.41e-20
C15728 _002_ _067_ 1.66e-21
C15729 net13 clknet_0_clk 0.0596f
C15730 a_9595_1679# _032_ 0.169f
C15731 _122_ a_12153_8757# 6.01e-21
C15732 net32 a_13880_3677# 6.05e-20
C15733 a_6173_7119# cal_itt\[3\] 4.34e-19
C15734 a_10864_7387# a_10990_7485# 0.186f
C15735 a_6741_7361# a_6785_7119# 3.69e-19
C15736 a_10903_7261# a_11059_7356# 0.113f
C15737 a_6523_7119# a_6619_7119# 0.0138f
C15738 _102_ mask\[3\] 1.05e-19
C15739 _117_ _057_ 7.58e-20
C15740 clknet_2_1__leaf_clk a_7351_8041# 6.69e-20
C15741 net8 a_13869_1501# 4.44e-19
C15742 a_3461_5193# VPWR 0.00302f
C15743 a_11509_3317# a_13183_3311# 1.96e-19
C15744 a_12077_3285# a_12424_3689# 0.0512f
C15745 a_7631_12319# net27 0.0716f
C15746 a_8731_9295# VPWR 0.222f
C15747 _042_ a_3399_10217# 3.04e-19
C15748 a_561_6031# a_1019_6397# 0.0346f
C15749 a_14715_3615# a_15023_2767# 0.00807f
C15750 net28 ctlp[7] 0.00152f
C15751 a_14540_3689# a_14604_3017# 1.43e-19
C15752 a_5915_10927# a_6467_9845# 1.96e-20
C15753 cal_count\[3\] _048_ 0.0554f
C15754 cal_count\[0\] a_14565_9295# 0.00164f
C15755 a_8839_9661# _068_ 2.26e-19
C15756 mask\[4\] a_6090_10159# 0.0106f
C15757 net47 a_12341_8751# 1.31e-20
C15758 _058_ a_15083_4659# 0.0029f
C15759 state\[2\] a_4709_2773# 0.0798f
C15760 net4 a_5087_3855# 2.18e-20
C15761 a_4425_6031# net3 6.11e-19
C15762 _037_ VPWR 1.06f
C15763 _125_ a_14981_8235# 5.76e-19
C15764 _134_ a_14282_7119# 5.12e-19
C15765 clknet_2_1__leaf_clk a_4030_9839# 6.85e-20
C15766 a_5915_11721# mask\[4\] 1.03e-20
C15767 a_1585_4777# VPWR 2.13e-19
C15768 a_6835_7669# a_7447_8041# 3.82e-19
C15769 a_7001_7669# a_7256_8029# 0.0612f
C15770 _063_ a_11023_5108# 6.07e-20
C15771 a_3521_9813# clknet_2_0__leaf_clk 1.49e-20
C15772 a_5915_10927# VPWR 0.313f
C15773 state\[0\] a_4709_2773# 0.034f
C15774 net50 a_10195_1354# 0.00108f
C15775 _037_ a_12218_6397# 8.1e-21
C15776 net4 a_4443_1679# 5.02e-19
C15777 a_8583_3317# a_10699_3311# 6.17e-21
C15778 trim_mask\[4\] a_7320_3631# 4.14e-20
C15779 net30 _090_ 9.79e-21
C15780 a_3781_8207# a_4871_8181# 0.0424f
C15781 a_3615_8207# a_4696_8207# 0.102f
C15782 a_4349_8449# a_4131_8207# 0.21f
C15783 net45 a_5633_1679# 6.03e-19
C15784 _050_ clknet_2_2__leaf_clk 0.00221f
C15785 net40 cal_count\[1\] 0.0105f
C15786 a_4308_4917# state\[0\] 1.55e-21
C15787 a_4091_5309# a_3667_3829# 1.47e-20
C15788 a_5915_10927# a_5699_9269# 9.71e-22
C15789 a_2143_2229# ctln[1] 1.75e-20
C15790 a_12231_6005# VPWR 0.36f
C15791 net19 a_8949_6031# 6.7e-19
C15792 net44 a_5363_7369# 0.0642f
C15793 net12 a_7256_8029# 2.34e-19
C15794 a_11394_9509# _001_ 5.8e-20
C15795 a_6056_8359# a_5691_7637# 0.00349f
C15796 _113_ _030_ 0.0189f
C15797 mask\[4\] a_7201_9813# 0.0219f
C15798 net49 a_14099_3017# 0.0484f
C15799 a_2877_2197# a_3386_2223# 2.6e-19
C15800 a_11491_6031# a_11587_6031# 0.0138f
C15801 cal_count\[3\] a_11599_6397# 0.0265f
C15802 a_4043_10143# _019_ 0.002f
C15803 net47 a_10864_7387# 0.0345f
C15804 a_6191_12559# net12 2.04e-19
C15805 a_13880_3677# VPWR 0.1f
C15806 clknet_2_1__leaf_clk a_7548_10217# 0.00435f
C15807 _063_ a_8307_6575# 0.0985f
C15808 a_8091_7967# _071_ 0.0266f
C15809 a_1467_7923# VPWR 0.456f
C15810 clknet_2_2__leaf_clk _052_ 2.54e-20
C15811 net50 _032_ 0.0063f
C15812 a_2383_3689# a_2948_3689# 7.99e-20
C15813 _101_ a_4687_11231# 0.00102f
C15814 _087_ a_5931_4105# 0.0965f
C15815 clknet_2_0__leaf_clk a_1007_7119# 1.44e-19
C15816 _074_ a_6181_10633# 3.35e-20
C15817 net44 _101_ 0.158f
C15818 _051_ a_5081_4943# 1.85e-20
C15819 _078_ _041_ 0.409f
C15820 a_8301_8207# VPWR 0.00785f
C15821 a_13697_4373# VPWR 0.245f
C15822 _123_ en_co_clk 5.23e-20
C15823 _010_ _078_ 8.71e-19
C15824 net52 a_3053_8457# 0.0143f
C15825 cal_count\[0\] a_14335_7895# 4.49e-21
C15826 _074_ a_745_12021# 0.00484f
C15827 a_6519_3829# a_5931_4105# 5.4e-20
C15828 net29 a_1095_12393# 0.00118f
C15829 a_1644_12533# a_1835_12319# 5.15e-19
C15830 a_911_4777# valid 0.00124f
C15831 a_4959_9295# net45 4.28e-20
C15832 a_8072_11721# VPWR 0.175f
C15833 a_1461_10357# a_1651_10143# 6.89e-19
C15834 net55 _051_ 0.121f
C15835 _136_ a_11583_4777# 0.00139f
C15836 a_11116_8983# _001_ 1.8e-19
C15837 a_11057_4105# trim_mask\[3\] 1.18e-20
C15838 a_14715_3615# a_15299_3311# 4.74e-19
C15839 a_5363_7369# en_co_clk 3.94e-20
C15840 _047_ trim[0] 5.54e-19
C15841 a_4498_4373# a_4617_4105# 8.58e-19
C15842 clknet_2_1__leaf_clk net25 0.367f
C15843 net18 a_9761_1679# 1.54e-19
C15844 a_9621_8029# VPWR 2.14e-19
C15845 net46 a_14649_3689# 6.24e-19
C15846 net40 _108_ 1.01f
C15847 mask\[4\] a_9182_10749# 2.86e-20
C15848 net21 ctlp[7] 0.0401f
C15849 a_8455_10383# a_9020_10383# 7.99e-20
C15850 mask\[5\] a_6743_10933# 2.68e-19
C15851 net31 a_15289_7119# 1.37e-19
C15852 net9 _001_ 0.00129f
C15853 net9 a_11067_4405# 5.13e-22
C15854 net14 clknet_2_1__leaf_clk 0.0168f
C15855 _065_ a_11369_7119# 1.91e-19
C15856 net38 trimb[2] 0.0166f
C15857 state\[0\] a_2288_3677# 1.44e-20
C15858 net12 mask\[1\] 1.8e-20
C15859 a_13783_6183# trim_mask\[0\] 3.95e-20
C15860 a_4680_6031# net54 5.27e-21
C15861 _094_ VPWR 0.382f
C15862 _101_ en_co_clk 0.00249f
C15863 clknet_2_0__leaf_clk net41 0.123f
C15864 _074_ _014_ 1.05e-21
C15865 net27 a_5915_10927# 8.68e-19
C15866 a_8105_10383# a_8673_10625# 0.181f
C15867 a_4043_10143# VPWR 0.39f
C15868 a_7939_10383# net47 0.296f
C15869 a_14347_4917# a_14655_4399# 0.0125f
C15870 trim_mask\[2\] a_13975_3689# 2.97e-20
C15871 _122_ a_13050_7637# 0.00579f
C15872 _033_ a_8491_2229# 6.44e-20
C15873 _051_ a_7715_3285# 0.21f
C15874 _065_ a_4227_8207# 2.56e-20
C15875 net42 _054_ 1.86e-19
C15876 net51 a_7569_7637# 4.95e-19
C15877 a_1651_10143# _018_ 3.75e-19
C15878 a_1476_10217# a_2787_9845# 3.19e-20
C15879 a_8298_2767# a_8657_2229# 0.0169f
C15880 net25 a_2368_9955# 0.12f
C15881 _080_ result[1] 8.38e-19
C15882 a_13279_8207# _133_ 1.3e-20
C15883 net44 a_6785_7119# 0.00316f
C15884 _079_ a_911_4777# 8.18e-20
C15885 a_4655_10071# a_5177_9537# 0.00173f
C15886 _093_ a_1867_3317# 2.78e-20
C15887 a_7527_4631# a_7891_3617# 6.04e-21
C15888 a_14981_4020# trim_val\[1\] 3.66e-20
C15889 _010_ a_3597_10933# 3.98e-19
C15890 calibrate a_2309_2229# 4.8e-21
C15891 a_2787_10927# a_2869_10927# 0.171f
C15892 net18 a_10787_1135# 0.00664f
C15893 a_3303_7119# _120_ 1.27e-19
C15894 a_6927_12559# a_7109_11989# 0.0034f
C15895 _104_ _028_ 4.91e-20
C15896 a_8657_2229# a_9681_2601# 2.36e-20
C15897 a_9007_2601# a_9269_2589# 0.00171f
C15898 a_6633_9845# a_7710_9839# 1.46e-19
C15899 net19 _062_ 0.248f
C15900 a_7201_9813# a_7091_9839# 0.0977f
C15901 _092_ a_7800_4631# 4.21e-21
C15902 _111_ a_12502_4765# 7.11e-19
C15903 net55 a_5445_4399# 0.00139f
C15904 mask\[0\] a_4425_6031# 5.23e-20
C15905 a_4239_8573# clknet_0_clk 4.43e-19
C15906 net13 net41 0.00634f
C15907 _107_ a_6737_3855# 7.76e-19
C15908 a_10903_7261# a_11016_6691# 1.21e-20
C15909 _090_ state\[2\] 3.14e-19
C15910 _096_ a_5363_4719# 1.97e-20
C15911 clknet_2_0__leaf_clk a_6523_7119# 1.49e-19
C15912 mask\[5\] _044_ 0.162f
C15913 a_13783_6183# a_13933_6281# 0.00899f
C15914 _048_ _119_ 6.77e-19
C15915 a_2787_7119# VPWR 0.479f
C15916 a_8455_10383# a_8731_9295# 1.15e-19
C15917 a_9195_10357# a_8949_9537# 2.87e-20
C15918 a_9020_10383# a_8381_9295# 0.00107f
C15919 _090_ state\[0\] 1.04e-19
C15920 a_8563_10749# _068_ 1.1e-21
C15921 net27 a_8072_11721# 0.107f
C15922 _047_ a_15023_2767# 2.51e-19
C15923 a_10239_9295# cal_count\[0\] 1.14e-19
C15924 a_10688_9295# a_11244_9661# 0.00329f
C15925 trim_mask\[0\] a_10975_4105# 0.177f
C15926 net19 a_9195_3689# 7.16e-19
C15927 a_3431_10933# a_4512_11305# 0.102f
C15928 _022_ a_4687_11231# 4.61e-20
C15929 _049_ a_6737_3855# 0.0486f
C15930 a_6703_2197# clk 5.3e-21
C15931 a_13825_5185# VPWR 0.221f
C15932 net24 a_3840_8867# 0.105f
C15933 cal_itt\[1\] _062_ 0.363f
C15934 _132_ a_15023_5487# 4.05e-20
C15935 a_1313_10901# a_911_10217# 0.00116f
C15936 a_745_10933# a_1651_10143# 3.39e-19
C15937 net18 a_11814_9295# 7.99e-19
C15938 a_9572_2601# a_10543_2455# 3.98e-19
C15939 net9 a_13512_1501# 3.67e-19
C15940 a_10975_6031# _136_ 0.0151f
C15941 net30 net50 3.8e-20
C15942 _024_ a_9802_4007# 1.08e-20
C15943 a_6375_12021# net44 0.299f
C15944 net49 net48 0.00261f
C15945 _036_ a_13356_8457# 0.00106f
C15946 net15 _092_ 0.167f
C15947 a_579_10933# a_561_9845# 2.81e-21
C15948 cal_count\[2\] a_13349_6031# 1.85e-20
C15949 _048_ a_6566_5193# 0.0172f
C15950 a_15023_6031# a_14972_5193# 1.06e-20
C15951 result[6] result[5] 0.035f
C15952 _123_ cal_count\[2\] 0.277f
C15953 a_2019_9055# net23 0.00142f
C15954 net33 a_15023_5487# 0.0075f
C15955 a_1095_12393# a_1191_12393# 0.0138f
C15956 _095_ _048_ 0.0407f
C15957 _051_ _093_ 1.44e-20
C15958 a_4617_3855# VPWR 2.85e-19
C15959 _006_ a_1229_8457# 0.0155f
C15960 _108_ _024_ 0.0014f
C15961 mask\[0\] a_3868_7119# 0.0388f
C15962 a_3208_10205# VPWR 0.0842f
C15963 a_2689_8751# VPWR 0.235f
C15964 _014_ _093_ 0.0073f
C15965 net28 a_1095_12393# 0.0102f
C15966 _121_ net3 1.77e-21
C15967 clknet_2_0__leaf_clk a_2767_2223# 0.0267f
C15968 _060_ clk 1.07e-20
C15969 clknet_2_0__leaf_clk a_1137_5487# 0.00371f
C15970 _101_ a_4801_9839# 0.0373f
C15971 en_co_clk _060_ 0.00965f
C15972 a_11394_9509# a_11116_8983# 7.41e-21
C15973 net45 a_2601_3285# 0.165f
C15974 a_10688_9295# _123_ 9.46e-22
C15975 clknet_0_clk a_4167_6575# 0.00409f
C15976 a_561_7119# a_1007_7119# 2.28e-19
C15977 net46 a_14972_5193# 0.00116f
C15978 _078_ a_561_6031# 0.0115f
C15979 net40 a_12900_7663# 8.48e-21
C15980 trim_mask\[0\] a_13881_2741# 3.76e-20
C15981 mask\[2\] a_2815_9447# 0.0574f
C15982 mask\[7\] a_1660_11305# 0.0223f
C15983 a_9084_4515# a_8749_3317# 2.02e-21
C15984 a_7019_4407# a_7190_3855# 8.07e-20
C15985 a_11067_4405# trim_mask\[3\] 1.68e-20
C15986 net44 a_7986_10927# 3.33e-19
C15987 net21 a_4655_10071# 8.05e-21
C15988 net9 a_11394_9509# 0.0012f
C15989 _078_ a_3615_8207# 3.44e-19
C15990 net19 a_7999_11231# 0.00291f
C15991 net45 _039_ 0.214f
C15992 a_8381_9295# a_8731_9295# 0.22f
C15993 a_2865_4460# _014_ 0.171f
C15994 a_6793_8970# net2 4.99e-20
C15995 a_1651_7093# result[1] 1.68e-19
C15996 mask\[1\] result[2] 0.00154f
C15997 net18 a_11067_3017# 0.00591f
C15998 _122_ VPWR 1.1f
C15999 a_4425_6031# net54 3.54e-19
C16000 net43 net45 0.392f
C16001 _038_ _066_ 0.257f
C16002 net19 a_8745_6895# 0.00242f
C16003 a_11508_9295# _001_ 1.29e-19
C16004 a_1651_4703# _097_ 7.8e-21
C16005 a_1476_4777# a_3057_4719# 2e-20
C16006 a_7088_7119# VPWR 0.306f
C16007 clknet_0_clk _028_ 8.37e-20
C16008 a_2019_9055# a_2225_7663# 7.64e-22
C16009 _099_ state\[1\] 6.04e-22
C16010 _090_ _100_ 0.179f
C16011 clknet_2_3__leaf_clk _124_ 2.19e-19
C16012 calibrate _089_ 0.0219f
C16013 a_7351_8041# cal_itt\[3\] 6.56e-19
C16014 _033_ _032_ 5.83e-21
C16015 _074_ a_5535_8181# 0.00126f
C16016 net16 a_13512_4943# 4.27e-19
C16017 _041_ a_7001_7669# 7.19e-21
C16018 net38 net36 0.0522f
C16019 a_10055_2767# a_9761_1679# 1.22e-19
C16020 _063_ VPWR 2.18f
C16021 mask\[3\] a_5067_9661# 0.0228f
C16022 net9 a_13193_6031# 4.46e-19
C16023 cal_itt\[0\] a_10055_5487# 3.46e-19
C16024 a_14471_591# a_14931_591# 1.48e-19
C16025 mask\[6\] a_3852_11293# 0.0248f
C16026 mask\[2\] _081_ 0.0816f
C16027 net19 net11 0.0983f
C16028 net53 a_7259_11305# 8.7e-19
C16029 _065_ _099_ 3.14e-19
C16030 a_395_9845# a_561_9845# 0.887f
C16031 calibrate a_816_4765# 8.06e-19
C16032 net18 _092_ 4.21e-19
C16033 a_5363_12559# a_5496_12131# 0.005f
C16034 net44 a_7824_11305# 0.248f
C16035 a_14099_1929# a_14184_1679# 1.48e-19
C16036 net8 a_13393_1707# 1.62e-20
C16037 a_14347_9480# a_14983_9269# 0.0019f
C16038 VPWR ctln[6] 0.364f
C16039 _042_ a_2787_9845# 0.106f
C16040 _074_ _082_ 0.102f
C16041 a_395_4405# net1 4.25e-19
C16042 cal_itt\[1\] a_8745_6895# 0.0111f
C16043 a_11059_7356# a_11141_6031# 9.04e-20
C16044 a_9443_6059# _064_ 0.00158f
C16045 net12 _041_ 0.00956f
C16046 _091_ a_8298_5487# 0.00418f
C16047 _053_ a_4815_3031# 0.128f
C16048 a_11987_8757# a_12916_8751# 0.00159f
C16049 net46 a_12077_3285# 0.169f
C16050 _064_ a_11601_2229# 5.56e-20
C16051 a_745_10933# a_1191_11305# 2.28e-19
C16052 net12 a_7184_2339# 1.35e-19
C16053 _107_ _024_ 6.14e-21
C16054 trim_mask\[2\] trim_val\[1\] 1.73e-20
C16055 net43 a_3868_10217# 0.254f
C16056 a_7939_3855# clk 0.0124f
C16057 a_7104_3855# VPWR 5.39e-20
C16058 a_7181_2589# VPWR 6.18e-20
C16059 _096_ VPWR 0.938f
C16060 _123_ cal_count\[1\] 0.0248f
C16061 a_14335_7895# en_co_clk 2.85e-20
C16062 _108_ _029_ 0.104f
C16063 net23 a_3053_8457# 7.55e-20
C16064 a_4512_12393# a_4687_11231# 8.78e-21
C16065 mask\[6\] a_3947_11305# 0.0357f
C16066 en_co_clk a_4498_4373# 0.00613f
C16067 a_3273_4943# net3 1.3e-20
C16068 _082_ a_1279_9129# 9.95e-19
C16069 a_4864_1679# clk 0.0164f
C16070 cal_count\[0\] a_11545_9049# 0.258f
C16071 _136_ a_15023_5487# 4.5e-19
C16072 a_7939_10383# _068_ 1.08e-20
C16073 net46 a_9503_4399# 4.18e-20
C16074 a_15259_7637# _131_ 0.0115f
C16075 _011_ VPWR 0.714f
C16076 a_3399_7119# _092_ 1.66e-20
C16077 net48 a_14172_1513# 4.81e-19
C16078 _032_ a_10785_1679# 1.04e-20
C16079 net30 _106_ 0.084f
C16080 _059_ _060_ 0.654f
C16081 a_12992_8751# a_15023_8751# 1.1e-20
C16082 clknet_2_2__leaf_clk a_13233_4737# 3.94e-19
C16083 _015_ a_2309_2229# 5.56e-20
C16084 net29 a_1461_10357# 8.48e-19
C16085 net25 result[4] 1.25e-20
C16086 clknet_2_2__leaf_clk a_7891_3617# 6.96e-20
C16087 a_13519_4007# a_13459_3317# 0.00308f
C16088 net13 a_4512_11305# 0.0152f
C16089 _074_ a_1007_10217# 0.00204f
C16090 trim_mask\[0\] a_9099_3689# 4.83e-20
C16091 clknet_2_1__leaf_clk a_7477_10901# 4.73e-19
C16092 _084_ a_5998_11471# 0.00151f
C16093 net49 trim[0] 1.66e-19
C16094 _047_ trim[4] 0.0025f
C16095 _053_ a_9443_6059# 0.0834f
C16096 _076_ a_4680_6031# 3.97e-20
C16097 net14 result[4] 8.01e-20
C16098 net45 a_2857_7637# 0.158f
C16099 a_4209_11293# VPWR 3.44e-19
C16100 mask\[0\] _121_ 0.00291f
C16101 net4 a_3302_3677# 4.88e-20
C16102 _048_ calibrate 0.262f
C16103 net43 a_2953_7119# 0.0243f
C16104 _065_ a_10877_7983# 8.6e-21
C16105 a_13697_4373# _110_ 0.00533f
C16106 _010_ a_3852_12381# 0.159f
C16107 _067_ a_10005_6031# 0.0161f
C16108 _122_ a_14807_8359# 5.33e-20
C16109 net4 _051_ 0.333f
C16110 _123_ a_12612_8725# 0.0317f
C16111 net41 a_2948_3689# 0.0403f
C16112 a_4617_4105# a_4576_3427# 7.35e-20
C16113 cal_itt\[0\] a_9823_6941# 7.96e-19
C16114 _109_ a_13519_4007# 1.23e-19
C16115 _002_ a_7001_7669# 0.23f
C16116 _071_ _107_ 2.52e-19
C16117 net4 _014_ 5.39e-20
C16118 trim_mask\[0\] a_10055_5487# 0.0872f
C16119 a_1493_5487# sample 3.8e-19
C16120 _058_ a_12533_3689# 1e-20
C16121 trim_mask\[4\] a_6737_3855# 1.96e-19
C16122 _065_ a_4259_6031# 0.0302f
C16123 trim_mask\[4\] a_6941_2589# 0.00102f
C16124 a_13091_1141# a_14172_1513# 0.102f
C16125 net53 _008_ 0.028f
C16126 a_13257_1141# a_14347_1439# 0.0424f
C16127 a_13825_1109# a_13607_1513# 0.21f
C16128 _025_ a_11509_3317# 0.219f
C16129 a_11343_3317# a_12077_3285# 0.0535f
C16130 a_929_8757# a_1375_9129# 2.28e-19
C16131 net9 a_12436_9129# 0.0108f
C16132 a_937_4105# a_995_3530# 7.12e-21
C16133 _013_ a_455_3571# 2.01e-20
C16134 a_13459_3317# a_14604_3017# 3.35e-19
C16135 _030_ a_13881_2741# 0.00419f
C16136 a_11509_3317# _026_ 1.18e-19
C16137 a_1313_11989# a_1095_12393# 0.21f
C16138 a_745_12021# a_1835_12319# 0.0424f
C16139 clknet_2_1__leaf_clk a_4165_11989# 0.0433f
C16140 a_11394_9509# a_11508_9295# 1.84e-19
C16141 a_11244_9661# a_11436_9295# 0.00536f
C16142 a_4775_6031# _090_ 8.11e-22
C16143 _053_ a_5087_3855# 8.25e-20
C16144 net30 _033_ 2.25e-21
C16145 a_12148_4777# a_13697_4373# 4.92e-20
C16146 a_12323_4703# _058_ 0.0143f
C16147 net46 a_9747_2527# 0.336f
C16148 a_14335_4020# net49 0.111f
C16149 _053_ a_12061_7669# 1.6e-19
C16150 a_14604_2339# a_15023_2223# 0.001f
C16151 _004_ a_561_6031# 0.223f
C16152 a_395_6031# a_1129_6273# 0.0626f
C16153 a_5455_4943# VPWR 0.422f
C16154 _095_ a_2033_3317# 1.18e-19
C16155 net18 a_11045_5807# 5.13e-19
C16156 a_13557_7369# _134_ 8.56e-20
C16157 clknet_2_1__leaf_clk _019_ 0.00835f
C16158 net43 a_3399_10217# 0.00449f
C16159 net12 _002_ 4.08e-19
C16160 a_15159_9269# trimb[4] 9.58e-19
C16161 clknet_0_clk _094_ 0.0166f
C16162 net50 a_11030_1679# 1.92e-19
C16163 net12 _050_ 0.0242f
C16164 a_5055_1679# ctln[7] 6.41e-20
C16165 net53 a_5524_9295# 9.34e-20
C16166 net40 trim_mask\[4\] 0.00108f
C16167 trim_mask\[0\] _088_ 0.0317f
C16168 net46 _111_ 0.00637f
C16169 _017_ a_4871_8181# 3.61e-20
C16170 net45 a_1173_6031# 0.00316f
C16171 a_13307_1707# a_13607_1513# 2.63e-20
C16172 a_13881_1653# a_13825_1109# 6.84e-20
C16173 net44 a_5067_9661# 0.0122f
C16174 net9 trim_mask\[3\] 0.0183f
C16175 a_13142_8725# cal_count\[1\] 0.00358f
C16176 _041_ a_13256_9117# 0.00205f
C16177 _011_ net27 0.0592f
C16178 a_10055_2767# a_11067_3017# 2.53e-20
C16179 a_3933_2767# a_4709_2773# 3.05e-19
C16180 net2 _134_ 0.501f
C16181 a_15023_12559# trimb[2] 0.00275f
C16182 net26 a_7723_10143# 0.11f
C16183 a_7262_5461# trim_mask\[0\] 3.41e-19
C16184 _048_ a_8298_5487# 0.00413f
C16185 a_1476_10217# a_763_8757# 3.96e-19
C16186 _071_ a_8495_6895# 0.00714f
C16187 net15 mask\[6\] 0.0927f
C16188 _065_ a_4043_7093# 8.51e-19
C16189 net43 a_2857_5461# 4.53e-20
C16190 a_6173_7119# _073_ 0.00579f
C16191 _003_ a_7723_6807# 4.94e-20
C16192 a_395_9845# _006_ 1.34e-21
C16193 _126_ a_12992_8751# 1.28e-21
C16194 _059_ a_4498_4373# 4.28e-19
C16195 _007_ a_763_8757# 1.26e-19
C16196 net46 a_12631_591# 1.71e-19
C16197 net12 _052_ 0.00248f
C16198 a_5340_6031# _050_ 3.29e-20
C16199 net12 a_5055_1679# 2.31e-19
C16200 _075_ a_7262_5461# 4.85e-20
C16201 net43 _069_ 7.84e-21
C16202 _074_ net22 0.191f
C16203 trim_mask\[0\] trim_val\[4\] 0.0422f
C16204 net29 a_745_10933# 1.03e-19
C16205 clknet_2_1__leaf_clk a_6467_9845# 0.266f
C16206 a_14335_7895# cal_count\[2\] 8.68e-19
C16207 _063_ _104_ 4.99e-20
C16208 net43 a_8022_7119# 4.46e-19
C16209 net12 _098_ 0.0253f
C16210 _101_ a_2787_10927# 0.118f
C16211 VPWR comp 0.245f
C16212 net14 cal 0.0197f
C16213 trim_mask\[0\] a_6519_4631# 2.03e-20
C16214 mask\[1\] _040_ 0.41f
C16215 en_co_clk a_13441_6281# 3.47e-21
C16216 _051_ a_6763_5193# 4.51e-19
C16217 a_2857_7637# a_2953_7119# 0.0204f
C16218 clknet_0_clk a_2787_7119# 0.00149f
C16219 net26 a_1476_10217# 1.19e-19
C16220 a_448_10357# net25 3.74e-20
C16221 a_11016_6691# a_11141_6031# 2.51e-20
C16222 net12 a_3615_8207# 1.15e-21
C16223 a_1000_11293# result[5] 2.53e-19
C16224 clknet_2_1__leaf_clk VPWR 6.38f
C16225 net34 a_15023_5487# 0.018f
C16226 a_10111_1679# a_10219_2045# 0.0572f
C16227 a_13307_1707# a_13881_1653# 0.00979f
C16228 a_10975_6031# cal_count\[3\] 0.0348f
C16229 _038_ a_12056_6031# 3.1e-19
C16230 _103_ a_7019_4407# 0.00696f
C16231 a_15023_8751# _132_ 7.25e-21
C16232 a_14172_1513# a_14281_1513# 0.00742f
C16233 a_14347_1439# a_14526_1501# 0.0074f
C16234 a_13825_1109# a_14334_1135# 2.6e-19
C16235 a_13607_1513# a_13715_1135# 0.0572f
C16236 _116_ _057_ 6.5e-20
C16237 net26 _007_ 0.00175f
C16238 _061_ net35 0.0122f
C16239 a_14379_6397# _058_ 1.98e-20
C16240 a_13825_5185# _110_ 7.59e-20
C16241 calibrate a_7021_4105# 0.0408f
C16242 a_13625_3317# a_14715_3615# 0.0424f
C16243 a_14193_3285# a_13975_3689# 0.21f
C16244 mask\[4\] a_4609_9295# 0.0011f
C16245 cal_itt\[0\] cal_itt\[2\] 0.136f
C16246 a_12153_8757# a_12992_8751# 0.0573f
C16247 net45 a_1638_7485# 1.41e-19
C16248 _015_ a_4609_1679# 0.255f
C16249 a_8307_6575# _092_ 3.77e-20
C16250 net33 a_15023_8751# 0.00169f
C16251 _108_ trim_mask\[1\] 0.0105f
C16252 a_14334_5309# trim[4] 9.46e-21
C16253 clknet_2_1__leaf_clk a_5699_9269# 5.83e-20
C16254 a_2953_9845# a_3868_10217# 0.125f
C16255 net16 a_14471_591# 2.4e-20
C16256 net30 _054_ 0.0194f
C16257 _067_ a_10877_7983# 1.96e-20
C16258 _092_ a_7460_5807# 0.00259f
C16259 net31 a_15023_2223# 0.00225f
C16260 trim_mask\[0\] a_14281_4943# 0.00108f
C16261 net31 _134_ 4.59e-22
C16262 net46 a_13257_1141# 0.042f
C16263 _104_ a_7104_3855# 3.55e-19
C16264 _076_ a_4425_6031# 3.9e-20
C16265 a_9761_1679# VPWR 0.627f
C16266 _126_ a_15111_9295# 1.43e-19
C16267 _083_ a_5535_8181# 1.29e-20
C16268 _038_ _058_ 0.00111f
C16269 _081_ a_2174_8457# 0.00117f
C16270 a_1129_6273# net30 4.59e-21
C16271 _078_ a_2019_9055# 0.0767f
C16272 _123_ a_12900_7663# 0.0867f
C16273 net19 a_7631_12319# 0.00166f
C16274 a_2368_9955# VPWR 0.159f
C16275 a_9802_4007# a_8749_3317# 0.0013f
C16276 a_6099_10633# a_8105_10383# 1.81e-20
C16277 net35 a_13257_4943# 8.54e-19
C16278 a_13091_4943# a_13697_4373# 3.01e-20
C16279 trim_mask\[2\] a_12424_3689# 7.08e-20
C16280 a_13881_1653# a_13715_1135# 5.04e-20
C16281 a_8381_9295# _063_ 8.5e-21
C16282 a_3667_3829# state\[0\] 0.234f
C16283 _092_ a_6927_3311# 4.55e-21
C16284 a_8298_2767# a_7223_2465# 3.93e-19
C16285 _016_ a_4043_7093# 6.74e-20
C16286 a_5363_7369# _049_ 7.59e-19
C16287 _108_ a_8749_3317# 3.78e-19
C16288 en_co_clk _066_ 2.69e-21
C16289 _062_ a_10188_4105# 3.02e-20
C16290 _024_ trim_mask\[4\] 4.44e-19
C16291 _065_ a_10864_7387# 0.0205f
C16292 net1 a_2283_4020# 1.02e-19
C16293 cal_itt\[3\] a_8307_6575# 0.169f
C16294 a_2787_10927# _102_ 0.00446f
C16295 _118_ net50 0.00284f
C16296 net19 a_9020_10383# 0.0132f
C16297 a_7184_2339# a_7524_2223# 0.0346f
C16298 _008_ a_6007_9839# 0.15f
C16299 a_8491_2229# a_8912_2589# 0.0867f
C16300 trim_mask\[0\] a_8745_4943# 4.46e-19
C16301 _092_ a_5363_4719# 0.0243f
C16302 a_9043_6031# _107_ 8.43e-20
C16303 _127_ _125_ 0.0731f
C16304 _051_ a_7689_2589# 2.63e-19
C16305 net46 a_10676_1679# 0.268f
C16306 cal_itt\[2\] a_7569_7637# 6.11e-19
C16307 a_14000_4719# a_13915_4399# 1.48e-19
C16308 _053_ a_11396_6031# 2.94e-20
C16309 cal_itt\[3\] a_7460_5807# 1.94e-19
C16310 _128_ net40 2.4e-21
C16311 a_13111_6031# VPWR 0.389f
C16312 _074_ a_6541_12021# 2.25e-19
C16313 _101_ _049_ 0.00159f
C16314 _126_ a_14422_7093# 4.82e-20
C16315 a_10787_1135# VPWR 0.236f
C16316 a_3597_12021# a_4055_12015# 0.0346f
C16317 en_co_clk a_4175_4943# 9.46e-20
C16318 net33 trim_val\[0\] 0.0273f
C16319 clknet_2_0__leaf_clk a_4995_7119# 0.0446f
C16320 net14 a_561_4405# 0.0145f
C16321 net43 a_4621_11305# 3.93e-19
C16322 a_9099_3689# a_8298_2767# 0.00882f
C16323 clknet_0_clk a_7088_7119# 3.47e-19
C16324 a_7245_10205# VPWR 1.18e-19
C16325 net44 a_7456_12393# 0.247f
C16326 VPWR trim[3] 0.564f
C16327 net52 a_6056_8359# 0.00104f
C16328 calibrate a_2033_3317# 4.87e-20
C16329 _063_ _110_ 6.44e-20
C16330 net47 _070_ 0.00159f
C16331 _048_ _015_ 2.39e-20
C16332 cal_count\[1\] a_14335_7895# 5.21e-20
C16333 clknet_2_1__leaf_clk net27 0.0557f
C16334 a_2815_9447# a_4609_9295# 1.58e-20
C16335 mask\[3\] net45 4.53e-21
C16336 net14 mask\[6\] 4.06e-22
C16337 clknet_0_clk _063_ 0.0459f
C16338 a_11859_3689# a_11955_3689# 0.0138f
C16339 trim_mask\[1\] a_12516_2601# 2.78e-20
C16340 _020_ a_8215_9295# 0.00106f
C16341 trim_mask\[3\] a_10689_2543# 0.00366f
C16342 _035_ a_10864_9269# 1.2e-19
C16343 a_10239_9295# a_10688_9295# 0.209f
C16344 net3 a_4091_5309# 0.0689f
C16345 net19 _028_ 0.00127f
C16346 net18 trim_val\[3\] 0.00706f
C16347 a_2787_10927# _022_ 0.11f
C16348 a_5177_9537# mask\[1\] 2.24e-20
C16349 _126_ _132_ 9.98e-21
C16350 a_2953_9845# a_3399_10217# 2.28e-19
C16351 net18 _035_ 0.0212f
C16352 _027_ a_9572_2601# 0.0566f
C16353 a_8491_2229# a_10543_2455# 1.16e-20
C16354 _090_ a_3933_2767# 8.23e-21
C16355 _035_ a_10820_7485# 1.07e-21
C16356 net16 a_13307_1707# 3.67e-19
C16357 net44 _043_ 1.13e-20
C16358 cal_itt\[2\] trim_mask\[0\] 1.07e-20
C16359 a_7571_4943# clk 0.00295f
C16360 net28 a_745_10933# 4.64e-20
C16361 net44 a_6515_6794# 1.06e-20
C16362 net46 a_14526_1501# 0.00288f
C16363 _108_ _115_ 0.00253f
C16364 net33 _126_ 0.46f
C16365 cal_count\[2\] a_13441_6281# 2.46e-19
C16366 net13 a_4995_7119# 0.00419f
C16367 mask\[2\] a_3781_8207# 5.9e-19
C16368 _064_ _025_ 1.51e-19
C16369 a_11814_9295# VPWR 0.184f
C16370 _064_ _026_ 9.32e-20
C16371 net40 a_12723_4943# 0.0221f
C16372 a_1095_11305# net52 1.38e-19
C16373 net20 a_7565_12393# 8.49e-20
C16374 a_1835_11231# a_1660_11305# 0.234f
C16375 a_1953_9129# VPWR 5.34e-19
C16376 _014_ a_3057_4719# 0.0476f
C16377 a_1129_7361# a_1019_7485# 0.0977f
C16378 a_1651_7093# a_1476_7119# 0.234f
C16379 a_8749_3317# a_9004_3677# 0.0642f
C16380 a_7459_7663# a_7088_7119# 1.35e-19
C16381 a_11141_6031# a_11709_6273# 0.169f
C16382 a_6485_8181# VPWR 0.166f
C16383 a_15299_6575# a_15023_5487# 3.56e-20
C16384 net19 a_8731_9295# 0.0109f
C16385 a_11622_7485# VPWR 0.0846f
C16386 mask\[0\] a_1651_7093# 0.0103f
C16387 trim_mask\[2\] a_11435_2229# 2.31e-19
C16388 clknet_0_clk _096_ 0.0288f
C16389 net18 _136_ 0.0321f
C16390 a_12992_8751# a_13050_7637# 5.58e-20
C16391 state\[2\] _054_ 1.37e-20
C16392 a_13142_8725# a_12900_7663# 7.12e-20
C16393 a_11583_4777# a_11679_4777# 0.0138f
C16394 a_10820_7485# _136_ 1.97e-21
C16395 net21 a_6191_12559# 1.65e-19
C16396 _108_ a_7939_3855# 1.1e-19
C16397 _107_ a_8749_3317# 0.00241f
C16398 mask\[7\] a_579_10933# 0.0132f
C16399 trim_val\[1\] a_14604_2339# 5.65e-19
C16400 mask\[3\] a_3868_10217# 1.86e-21
C16401 net15 a_3317_8207# 4.75e-19
C16402 a_13091_4943# a_13825_5185# 0.0623f
C16403 net50 a_10137_4943# 1.62e-19
C16404 _060_ _107_ 0.00674f
C16405 a_4866_12381# VPWR 8.13e-20
C16406 a_6515_6794# clk 4.17e-19
C16407 a_11601_2229# a_10689_2223# 3.97e-19
C16408 net26 _042_ 0.0409f
C16409 a_11951_2601# a_12047_2601# 0.0138f
C16410 net45 a_3578_2589# 0.00342f
C16411 net29 _010_ 8.13e-20
C16412 _046_ a_2910_12131# 4.96e-19
C16413 a_448_7637# net22 6.71e-20
C16414 net45 a_1579_5807# 1.19e-19
C16415 a_13825_6031# VPWR 0.0118f
C16416 _050_ a_5691_2741# 0.327f
C16417 _058_ a_10270_4105# 9.62e-19
C16418 cal_itt\[3\] a_7897_6913# 0.00121f
C16419 clknet_2_1__leaf_clk a_8455_10383# 1.49e-19
C16420 _136_ a_12165_6031# 1.18e-19
C16421 mask\[4\] a_6181_10633# 0.0015f
C16422 _120_ a_3891_4943# 0.183f
C16423 net2 a_5691_7637# 5.89e-19
C16424 _041_ _040_ 4.32e-20
C16425 a_3116_12533# _074_ 3.47e-20
C16426 trim_val\[4\] a_8298_2767# 1.41e-19
C16427 clknet_2_0__leaf_clk a_3224_2601# 0.0701f
C16428 a_6007_7119# VPWR 0.502f
C16429 a_7210_5807# _088_ 6.59e-20
C16430 a_1313_11989# a_1461_10357# 1.88e-22
C16431 net25 a_1763_9295# 5.39e-20
C16432 _101_ _008_ 0.00877f
C16433 _049_ _060_ 0.00176f
C16434 a_3208_7119# net30 5.56e-19
C16435 _067_ a_10864_7387# 2.16e-19
C16436 a_11067_3017# VPWR 0.205f
C16437 a_937_4105# valid 0.00145f
C16438 a_561_9845# a_911_10217# 0.217f
C16439 a_7262_5461# a_7210_5807# 0.0212f
C16440 a_14193_3285# trim_val\[1\] 9.6e-19
C16441 a_14540_3689# a_14649_3689# 0.00742f
C16442 a_14715_3615# a_14894_3677# 0.0074f
C16443 a_13975_3689# a_14083_3311# 0.0572f
C16444 a_13519_4007# trim[1] 2.55e-20
C16445 a_911_4777# net1 0.00105f
C16446 _010_ a_3431_12021# 0.168f
C16447 _133_ a_13142_7271# 0.243f
C16448 a_12516_2601# _115_ 5.13e-21
C16449 a_2775_9071# a_2689_8751# 2.42e-19
C16450 a_4512_11305# a_5915_10927# 8.86e-20
C16451 _031_ net48 0.00259f
C16452 _106_ _118_ 0.00544f
C16453 _107_ a_9361_3677# 1.48e-19
C16454 net44 a_6743_10933# 0.319f
C16455 net40 net35 0.175f
C16456 _104_ a_9761_1679# 0.0025f
C16457 net40 a_13059_4631# 2.5e-20
C16458 _125_ _041_ 0.0167f
C16459 net37 a_14788_7369# 8.7e-20
C16460 calibrate a_6197_4399# 1.7e-21
C16461 net19 a_8072_11721# 0.00139f
C16462 net13 a_3224_2601# 2.3e-20
C16463 en_co_clk a_3557_5193# 0.00324f
C16464 _051_ _064_ 0.00148f
C16465 _101_ a_5524_9295# 0.0104f
C16466 net55 trim_mask\[0\] 0.0775f
C16467 _092_ VPWR 3.61f
C16468 a_12631_12559# net16 5.69e-19
C16469 cal_itt\[2\] a_8949_6281# 0.0327f
C16470 _062_ a_8745_6895# 0.00215f
C16471 clknet_0_clk a_5455_4943# 5.47e-20
C16472 a_9460_6807# a_8935_6895# 6.49e-20
C16473 clknet_2_2__leaf_clk a_12077_3285# 0.0443f
C16474 net43 a_2787_9845# 0.446f
C16475 trim_mask\[2\] a_14347_1439# 4.78e-20
C16476 _075_ net55 2.15e-19
C16477 a_14199_7369# VPWR 0.195f
C16478 a_14347_9480# a_14236_8457# 3.32e-19
C16479 _111_ a_11233_4405# 1.95e-19
C16480 net31 a_15054_5193# 2.19e-20
C16481 a_8307_4943# a_8745_4943# 0.013f
C16482 net31 trim_val\[1\] 0.0297f
C16483 a_7351_8041# _073_ 4.8e-21
C16484 _107_ a_7939_3855# 0.00468f
C16485 net44 net45 0.00514f
C16486 net14 result[0] 0.00258f
C16487 a_1129_6273# a_1585_6031# 4.2e-19
C16488 VPWR result[4] 0.264f
C16489 _035_ a_12153_8757# 7.63e-21
C16490 _038_ a_11488_4765# 2.76e-19
C16491 _001_ _037_ 7.89e-19
C16492 a_6909_10933# net26 2.1e-21
C16493 _129_ a_13783_6183# 6.02e-20
C16494 _031_ a_13091_1141# 0.167f
C16495 a_8636_9295# cal_itt\[0\] 7.63e-20
C16496 result[6] result[7] 0.0507f
C16497 _050_ _089_ 5.45e-21
C16498 net13 a_4863_4917# 0.0118f
C16499 clknet_2_2__leaf_clk a_9503_4399# 7.38e-19
C16500 a_4498_4373# _107_ 6.74e-19
C16501 a_5536_4399# a_5363_4719# 0.0326f
C16502 net13 a_3431_10933# 0.00283f
C16503 net44 _044_ 9.19e-19
C16504 en_co_clk a_12056_6031# 1.08e-19
C16505 cal_itt\[3\] VPWR 0.557f
C16506 a_9459_7895# a_9693_8029# 0.00517f
C16507 net15 a_3148_4399# 0.00192f
C16508 a_911_7119# net22 5.67e-19
C16509 a_12992_8751# VPWR 0.459f
C16510 a_455_12533# result[5] 6.68e-19
C16511 _049_ a_7939_3855# 0.00707f
C16512 a_6927_12559# VPWR 0.41f
C16513 a_6906_2355# VPWR 0.31f
C16514 a_9664_3689# a_10016_1679# 3.67e-21
C16515 _053_ _051_ 0.0391f
C16516 net34 a_15023_8751# 0.0147f
C16517 net43 a_2092_8457# 3.96e-19
C16518 a_12900_7663# a_14335_7895# 6.74e-20
C16519 _052_ _089_ 0.00686f
C16520 a_13050_7637# _132_ 5.78e-20
C16521 clknet_2_2__leaf_clk a_7942_2223# 6.21e-19
C16522 net15 a_3365_4943# 0.00261f
C16523 a_395_7119# result[0] 0.00211f
C16524 a_1313_11989# a_745_10933# 5.38e-22
C16525 cal_itt\[2\] a_8307_4943# 1.31e-19
C16526 a_745_12021# a_1313_10901# 5.17e-21
C16527 net40 _061_ 0.0224f
C16528 _049_ a_4498_4373# 0.0563f
C16529 net45 clk 0.323f
C16530 clknet_2_3__leaf_clk a_10903_7261# 0.469f
C16531 _015_ a_2033_3317# 7.75e-21
C16532 _072_ _070_ 0.0703f
C16533 _074_ a_4043_12393# 1.35e-20
C16534 net45 en_co_clk 2.3e-20
C16535 a_1007_6031# calibrate 2.23e-20
C16536 a_10851_1653# a_10752_565# 1.15e-19
C16537 clknet_2_1__leaf_clk clknet_0_clk 0.00737f
C16538 a_5177_9537# _041_ 5.07e-21
C16539 net28 _010_ 0.0643f
C16540 a_5177_1921# a_5686_2045# 2.6e-19
C16541 a_11601_2229# _057_ 3.06e-19
C16542 a_4959_1679# a_5067_2045# 0.0572f
C16543 a_4609_1679# a_5055_1679# 2.28e-19
C16544 _136_ a_11023_5108# 0.0027f
C16545 _074_ a_1476_10217# 5.17e-19
C16546 a_6523_7119# a_7088_7119# 7.99e-20
C16547 a_1129_6273# a_911_6031# 0.21f
C16548 a_561_6031# a_1651_6005# 0.0424f
C16549 _068_ _070_ 0.0108f
C16550 en_co_clk _058_ 9.63e-19
C16551 a_7259_11305# a_7824_11305# 7.99e-20
C16552 _043_ a_8992_9955# 0.105f
C16553 a_14347_9480# _129_ 7.54e-21
C16554 net41 a_7104_3855# 4.96e-22
C16555 a_9317_3285# VPWR 0.211f
C16556 _064_ a_10781_3311# 0.0165f
C16557 _065_ a_3748_6281# 0.181f
C16558 _074_ _007_ 0.117f
C16559 _096_ net41 1.83e-20
C16560 a_11244_9661# _128_ 2.37e-20
C16561 a_10239_9295# a_11436_9295# 1.63e-19
C16562 a_1099_12533# _074_ 1.54e-19
C16563 a_1660_12393# _078_ 7.59e-21
C16564 a_9084_4515# _058_ 3.24e-19
C16565 _129_ a_13142_7271# 1.27e-19
C16566 a_13519_4007# _112_ 0.171f
C16567 a_11067_4405# a_13697_4373# 1.9e-21
C16568 _110_ a_9761_1679# 0.0115f
C16569 clknet_2_0__leaf_clk a_3817_4697# 7.15e-20
C16570 a_4959_1679# a_5363_591# 1.95e-19
C16571 _065_ a_6056_8359# 0.158f
C16572 net40 a_13257_4943# 0.0137f
C16573 net43 a_2198_9117# 0.00196f
C16574 _009_ VPWR 0.35f
C16575 clknet_2_2__leaf_clk a_9747_2527# 0.00182f
C16576 _080_ a_1125_7663# 0.0993f
C16577 a_11856_2589# VPWR 0.0853f
C16578 _046_ a_2787_10927# 5.07e-19
C16579 net43 net51 0.382f
C16580 a_1476_10217# a_1279_9129# 2.66e-20
C16581 net25 a_1497_8725# 1.47e-19
C16582 trim_mask\[1\] trim_mask\[4\] 0.0742f
C16583 a_8495_6895# a_8935_6895# 0.0234f
C16584 a_10781_3311# a_10851_1653# 8.88e-21
C16585 a_395_4405# a_1476_4777# 0.102f
C16586 net12 _087_ 0.00185f
C16587 a_13562_8751# _133_ 6.44e-21
C16588 a_4775_6031# a_4883_6397# 0.0572f
C16589 a_911_10217# _006_ 2.82e-20
C16590 _040_ a_3615_8207# 0.359f
C16591 trim_mask\[4\] a_6703_2197# 0.0893f
C16592 net14 a_1497_8725# 6.88e-19
C16593 a_11987_8757# a_11575_8790# 7e-20
C16594 a_4091_5309# net54 0.0437f
C16595 net46 trim_mask\[2\] 0.25f
C16596 net34 trim_val\[0\] 8.77e-19
C16597 net12 a_6519_3829# 0.00707f
C16598 net43 a_4055_12015# 0.0173f
C16599 _050_ _048_ 0.175f
C16600 a_579_12021# ctlp[0] 0.00196f
C16601 VPWR cal 0.226f
C16602 a_12723_4943# _029_ 0.116f
C16603 _111_ clknet_2_2__leaf_clk 0.0731f
C16604 a_6927_591# ctln[7] 4.45e-20
C16605 _128_ _123_ 0.281f
C16606 cal_itt\[0\] a_10043_7983# 0.0109f
C16607 net44 a_2953_7119# 4.35e-20
C16608 net33 net32 1.61e-19
C16609 _126_ a_11987_8757# 1.75e-20
C16610 _118_ _054_ 8.99e-21
C16611 net12 _099_ 0.00188f
C16612 net13 a_5524_1679# 0.00312f
C16613 _066_ _108_ 0.0118f
C16614 a_9773_3689# VPWR 5.34e-19
C16615 _097_ _013_ 0.00171f
C16616 _104_ a_11067_3017# 0.233f
C16617 net46 a_12213_2589# 0.00316f
C16618 clknet_2_1__leaf_clk a_3521_9813# 0.00609f
C16619 _110_ a_10787_1135# 0.0517f
C16620 a_448_10357# VPWR 0.322f
C16621 net43 _003_ 0.00181f
C16622 trim_mask\[4\] a_8749_3317# 0.0256f
C16623 a_9369_4105# a_9099_3689# 5.26e-20
C16624 a_14083_3311# trim_val\[1\] 4.79e-19
C16625 net12 a_6927_591# 0.24f
C16626 _048_ _052_ 0.119f
C16627 a_855_4105# a_937_3855# 0.00393f
C16628 net18 a_9296_9295# 2.39e-19
C16629 a_14422_7093# VPWR 0.245f
C16630 a_4805_8207# VPWR 2.71e-20
C16631 mask\[1\] a_2143_7663# 0.0982f
C16632 a_6737_4719# VPWR 0.00429f
C16633 a_4165_11989# mask\[6\] 1.34e-21
C16634 a_929_8757# a_561_7119# 1.43e-21
C16635 a_3947_12393# a_4512_12393# 7.99e-20
C16636 net13 clknet_2_0__leaf_clk 0.164f
C16637 net34 _126_ 0.00327f
C16638 a_8301_8207# a_7916_8041# 3.77e-19
C16639 a_5340_6031# _099_ 2.94e-21
C16640 _048_ _098_ 0.24f
C16641 a_5547_5603# VPWR 0.137f
C16642 mask\[2\] a_1844_9129# 6.47e-20
C16643 a_15023_12559# net38 4.96e-20
C16644 net39 a_15023_12015# 0.0374f
C16645 trim_mask\[4\] a_10977_2543# 5.34e-19
C16646 a_14172_1513# _057_ 2.11e-20
C16647 mask\[6\] _019_ 1.18e-20
C16648 net55 a_8307_4943# 0.133f
C16649 net19 a_7088_7119# 2.19e-21
C16650 a_11987_8757# a_12153_8757# 0.549f
C16651 _092_ _104_ 1.49e-20
C16652 cal_itt\[0\] net4 0.122f
C16653 a_9003_3829# VPWR 0.277f
C16654 a_4687_12319# net13 4.31e-19
C16655 a_7456_12393# a_7618_12015# 0.00645f
C16656 net45 _059_ 1.18e-20
C16657 a_2787_9845# a_2953_9845# 0.586f
C16658 _132_ VPWR 0.778f
C16659 net19 _063_ 0.824f
C16660 _090_ a_5931_4105# 0.159f
C16661 net46 a_9719_1473# 3.42e-21
C16662 _074_ a_1357_11293# 5.87e-19
C16663 a_5536_4399# VPWR 0.252f
C16664 _129_ a_14870_7369# 1.39e-19
C16665 a_5067_2045# VPWR 0.136f
C16666 clknet_2_2__leaf_clk a_13257_1141# 0.00461f
C16667 _009_ net27 3.17e-19
C16668 net33 VPWR 1.02f
C16669 net18 cal_count\[3\] 0.423f
C16670 _123_ a_11895_7669# 0.519f
C16671 net55 a_8298_2767# 3.7e-19
C16672 a_13279_8207# cal_count\[2\] 4.49e-19
C16673 _029_ a_13059_4631# 1.07e-19
C16674 a_9664_3689# _025_ 6.48e-20
C16675 trim_mask\[4\] a_9361_3677# 0.00213f
C16676 trim_mask\[2\] a_11343_3317# 3.93e-19
C16677 state\[1\] a_4709_2773# 0.134f
C16678 _069_ a_9459_7895# 0.044f
C16679 en_co_clk a_4905_3855# 4.69e-20
C16680 a_4696_8207# a_6056_8359# 6.13e-20
C16681 _122_ cal_itt\[1\] 1.33e-20
C16682 trim_mask\[2\] a_11149_3017# 0.0116f
C16683 a_9602_6941# VPWR 8.79e-20
C16684 _076_ a_6885_8372# 0.246f
C16685 a_9459_7895# a_8022_7119# 0.0095f
C16686 a_5363_591# VPWR 0.472f
C16687 a_561_4405# VPWR 0.452f
C16688 net9 _037_ 0.11f
C16689 state\[2\] a_3339_2767# 2.77e-20
C16690 net14 a_1019_4399# 0.00176f
C16691 _133_ _131_ 0.00247f
C16692 a_4091_5309# a_4471_4007# 4.67e-19
C16693 net44 a_8022_7119# 0.00349f
C16694 net47 net2 0.0188f
C16695 a_12249_7663# a_12454_8041# 3.7e-19
C16696 net49 a_13625_3317# 0.0129f
C16697 mask\[5\] net26 0.00797f
C16698 mask\[0\] a_2225_7983# 0.0011f
C16699 cal_itt\[1\] _063_ 0.39f
C16700 a_15023_10927# net31 0.00817f
C16701 _026_ a_10689_2223# 1.11e-19
C16702 _083_ a_7079_10217# 2.45e-20
C16703 a_3868_10217# a_4801_9839# 2.52e-19
C16704 net12 a_4259_6031# 1.79e-21
C16705 _005_ a_1129_7361# 9.52e-19
C16706 state\[0\] a_3339_2767# 4.75e-21
C16707 net46 a_9595_1679# 0.345f
C16708 net15 a_3521_7361# 0.00236f
C16709 _128_ a_13142_8725# 0.0153f
C16710 mask\[6\] VPWR 0.717f
C16711 _074_ _042_ 0.448f
C16712 a_8307_6575# _105_ 9.22e-20
C16713 _050_ a_7021_4105# 0.00539f
C16714 clknet_2_2__leaf_clk a_10676_1679# 8.02e-20
C16715 a_3947_12393# _046_ 2.94e-19
C16716 net27 a_448_10357# 7.85e-21
C16717 a_8820_6005# _106_ 1.09e-20
C16718 mask\[2\] a_5633_9295# 3.77e-21
C16719 mask\[1\] _077_ 4.87e-19
C16720 _060_ a_3123_3615# 6.36e-21
C16721 a_9003_3829# a_9478_4105# 0.0127f
C16722 a_7939_3855# trim_mask\[4\] 7.91e-20
C16723 trim_val\[4\] a_9369_4105# 0.0263f
C16724 _065_ a_4308_4917# 0.131f
C16725 a_13783_6183# a_14379_6397# 0.0264f
C16726 en_co_clk a_2857_5461# 0.0217f
C16727 a_6375_12021# a_6891_12393# 0.115f
C16728 net9 a_12231_6005# 0.0146f
C16729 clknet_0_clk a_6007_7119# 1.07e-20
C16730 _078_ a_5997_11247# 1.96e-19
C16731 a_1476_7119# a_395_6031# 3.02e-20
C16732 net52 a_4349_8449# 7.52e-19
C16733 mask\[0\] a_395_6031# 0.0111f
C16734 a_4131_8207# mask\[0\] 1.57e-20
C16735 _082_ a_2815_9447# 1.82e-20
C16736 a_4259_6031# a_5340_6031# 0.102f
C16737 a_4993_6273# a_4775_6031# 0.21f
C16738 a_4425_6031# a_5515_6005# 0.0418f
C16739 a_8022_7119# clk 0.315f
C16740 _104_ a_9317_3285# 0.0473f
C16741 _046_ a_3425_11721# 0.0555f
C16742 a_8022_7119# en_co_clk 3.63e-19
C16743 net54 a_4886_4399# 0.00231f
C16744 _052_ a_7021_4105# 0.0718f
C16745 _007_ a_448_7637# 4.13e-20
C16746 _122_ _001_ 0.589f
C16747 a_8485_4943# VPWR 1.16e-19
C16748 clknet_2_0__leaf_clk a_561_7119# 0.00336f
C16749 a_8491_2229# _027_ 0.617f
C16750 a_10975_6031# _135_ 1.04e-20
C16751 _083_ a_7723_10143# 7.61e-22
C16752 _051_ a_7379_2197# 0.00194f
C16753 a_14604_2339# a_14686_2339# 0.00477f
C16754 a_579_10933# a_1677_9545# 5.86e-22
C16755 net13 a_4864_9295# 0.00788f
C16756 mask\[1\] a_1019_7485# 2.4e-19
C16757 net4 trim_mask\[0\] 0.0222f
C16758 a_2383_3689# cal 5.95e-20
C16759 clknet_2_1__leaf_clk a_6523_7119# 1.07e-19
C16760 trim_val\[3\] VPWR 0.258f
C16761 VPWR ctlp[2] 0.274f
C16762 _049_ a_4175_4943# 4.47e-20
C16763 mask\[2\] _017_ 0.0217f
C16764 _035_ VPWR 0.222f
C16765 a_7571_4943# _107_ 0.00449f
C16766 _023_ a_1095_11305# 0.00115f
C16767 clknet_0_clk _092_ 0.206f
C16768 a_579_10933# a_1835_11231# 0.0436f
C16769 _128_ a_14565_9295# 0.00206f
C16770 a_10569_1109# ctln[4] 8.88e-19
C16771 a_7010_3311# a_6927_3311# 0.188f
C16772 a_14807_8359# _132_ 9.11e-19
C16773 _085_ result[7] 1.61e-21
C16774 net43 a_763_8757# 0.303f
C16775 a_7256_8029# a_6173_7119# 2.4e-19
C16776 net33 a_14807_8359# 0.00892f
C16777 net46 net50 0.0769f
C16778 net15 _095_ 0.0835f
C16779 a_11987_8757# a_13050_7637# 2.07e-19
C16780 _036_ a_12344_8041# 6.1e-19
C16781 a_4165_10901# a_4055_10927# 0.0977f
C16782 a_4995_7119# _094_ 5.81e-20
C16783 mask\[3\] a_2787_9845# 0.00649f
C16784 a_3386_2223# clk 8.78e-20
C16785 a_395_6031# _079_ 2.27e-19
C16786 _029_ a_13257_4943# 0.218f
C16787 cal_count\[1\] a_13279_8207# 0.05f
C16788 _092_ a_10699_5487# 0.0688f
C16789 _049_ a_7571_4943# 0.00225f
C16790 trim_mask\[0\] a_14172_4943# 0.0462f
C16791 net2 net5 9.9e-19
C16792 _136_ VPWR 0.642f
C16793 _040_ a_4227_8207# 0.00527f
C16794 net17 a_11803_10383# 0.112f
C16795 _087_ a_5691_2741# 1.03e-19
C16796 _074_ a_6909_10933# 8.1e-21
C16797 mask\[6\] net27 0.348f
C16798 a_12249_7663# a_12430_7663# 8.75e-19
C16799 a_1763_9295# VPWR 1.28e-19
C16800 _088_ a_8307_4719# 2.94e-20
C16801 _129_ _131_ 0.00886f
C16802 net43 net26 0.0143f
C16803 a_12218_6397# _136_ 8.32e-20
C16804 _061_ a_13349_6031# 2.76e-20
C16805 _065_ _070_ 0.657f
C16806 clknet_0_clk cal_itt\[3\] 0.0237f
C16807 _069_ a_8091_7967# 5.34e-20
C16808 net3 state\[2\] 6.86e-20
C16809 _049_ a_4576_3427# 3.65e-19
C16810 a_7456_12393# a_7259_11305# 4.48e-20
C16811 _101_ a_3303_10217# 0.0338f
C16812 a_7631_12319# a_7999_11231# 9.77e-20
C16813 net43 a_5050_8207# 1.48e-19
C16814 trim_mask\[1\] a_11967_3311# 0.0265f
C16815 a_8091_7967# a_8022_7119# 0.00428f
C16816 a_4443_9295# a_5055_9295# 0.00188f
C16817 a_4609_9295# a_5686_9661# 1.46e-19
C16818 cal_count\[3\] a_11023_5108# 0.012f
C16819 _014_ a_3530_4438# 1.21e-19
C16820 a_13459_3317# a_14649_3689# 2.56e-19
C16821 net3 state\[0\] 0.135f
C16822 a_14347_9480# cal_count\[0\] 0.103f
C16823 _090_ state\[1\] 5.04e-20
C16824 _104_ a_9003_3829# 0.0821f
C16825 mask\[0\] net30 0.228f
C16826 _091_ a_10005_6031# 0.222f
C16827 a_8657_2229# clk 0.00144f
C16828 a_7916_8041# _063_ 2.71e-19
C16829 net18 _119_ 1.51e-19
C16830 net45 a_3399_2527# 0.337f
C16831 a_13059_4631# trim_mask\[1\] 2.13e-21
C16832 _026_ _057_ 0.00227f
C16833 _027_ a_10195_1354# 3.83e-21
C16834 a_2143_2229# net7 1.44e-20
C16835 net13 a_4239_8573# 0.00125f
C16836 net18 a_11258_9117# 3.63e-19
C16837 _128_ a_14335_7895# 1.51e-21
C16838 clknet_2_3__leaf_clk a_11141_6031# 0.526f
C16839 _110_ a_9317_3285# 0.00634f
C16840 _074_ a_3597_12021# 6.67e-19
C16841 net40 _024_ 5.23e-20
C16842 a_2787_7119# a_4995_7119# 6.12e-21
C16843 a_3521_7361# a_3399_7119# 3.16e-19
C16844 _048_ a_8389_5193# 0.0145f
C16845 clknet_2_0__leaf_clk a_2948_3689# 2.11e-21
C16846 net19 clknet_2_1__leaf_clk 5.46e-19
C16847 _065_ _090_ 1.37e-19
C16848 a_1549_6794# a_561_6031# 0.00105f
C16849 a_2019_9055# _040_ 3.64e-19
C16850 _108_ _058_ 0.228f
C16851 _012_ a_995_3530# 5.56e-21
C16852 VPWR result[0] 0.335f
C16853 net14 a_1129_7361# 0.0137f
C16854 net31 net5 0.0416f
C16855 a_9664_3689# a_10781_3311# 1.54e-19
C16856 _073_ a_7897_6913# 5.76e-19
C16857 a_1007_4777# cal 3.17e-19
C16858 a_448_6549# a_395_6031# 0.0112f
C16859 clknet_2_0__leaf_clk a_4167_6575# 0.0101f
C16860 net50 a_11343_3317# 5.21e-21
C16861 net9 a_13825_5185# 8.16e-20
C16862 _074_ a_1137_11721# 0.00107f
C16863 _070_ a_9761_8457# 1.01e-19
C16864 net14 a_1095_12393# 0.00272f
C16865 net34 net32 0.459f
C16866 a_10861_7119# VPWR 7.1e-20
C16867 net25 a_1638_9839# 2.35e-19
C16868 _090_ a_5054_4399# 0.0179f
C16869 a_11394_9509# _122_ 0.00536f
C16870 net37 _122_ 7.04e-21
C16871 a_14347_4917# trim_val\[0\] 0.0699f
C16872 _058_ a_10655_2932# 1.64e-19
C16873 trim_val\[2\] net48 0.0604f
C16874 net19 a_9761_1679# 2.89e-20
C16875 _027_ _032_ 5.79e-20
C16876 _115_ _056_ 4.69e-21
C16877 _078_ a_6056_8359# 9.44e-19
C16878 net8 a_12631_591# 3.66e-19
C16879 mask\[3\] net51 4.53e-21
C16880 a_4266_4943# VPWR 1.11e-19
C16881 a_929_8757# a_1467_7923# 3.37e-20
C16882 _021_ a_7933_11305# 2.14e-20
C16883 _000_ cal_itt\[0\] 1.21e-20
C16884 calibrate a_7800_4631# 3.13e-20
C16885 net51 a_6741_7361# 2.89e-19
C16886 _072_ net2 0.234f
C16887 net30 _079_ 0.0937f
C16888 _087_ _089_ 0.162f
C16889 a_395_7119# a_1129_7361# 0.0701f
C16890 clknet_2_1__leaf_clk a_4512_11305# 5.88e-20
C16891 a_3317_8207# VPWR 5.57e-19
C16892 _110_ a_9773_3689# 1.59e-19
C16893 _049_ a_3557_5193# 3.38e-21
C16894 _041_ _077_ 5.12e-20
C16895 _068_ net2 0.00928f
C16896 _048_ a_7891_3617# 3.58e-20
C16897 _089_ a_6519_3829# 0.111f
C16898 a_10699_5487# a_11045_5807# 0.0134f
C16899 a_11987_8757# VPWR 0.404f
C16900 a_1644_12533# result[7] 0.159f
C16901 net2 a_15023_6031# 0.00103f
C16902 a_11116_8983# _122_ 0.0652f
C16903 net3 _100_ 3.82e-21
C16904 net14 _095_ 1.78e-20
C16905 _099_ _089_ 9.94e-20
C16906 _037_ a_13470_7663# 5.93e-20
C16907 a_11764_3677# a_11955_3689# 4.61e-19
C16908 _094_ a_4863_4917# 0.0948f
C16909 net4 a_2877_2197# 0.00189f
C16910 _105_ VPWR 0.27f
C16911 net18 a_11679_4777# 6.77e-19
C16912 net46 _106_ 9.94e-21
C16913 net47 a_12249_7663# 1.05e-20
C16914 _078_ a_1095_11305# 0.00326f
C16915 a_395_4405# _014_ 1.2e-20
C16916 _066_ trim_mask\[4\] 2.16e-20
C16917 clknet_0_clk a_5547_5603# 0.0422f
C16918 a_14335_2442# a_13257_1141# 1.5e-19
C16919 a_9572_2601# _116_ 1.53e-20
C16920 trim_val\[2\] a_13091_1141# 2.46e-19
C16921 net31 a_15023_1679# 5.31e-19
C16922 net9 _122_ 0.0809f
C16923 _092_ net41 5.14e-20
C16924 net20 a_6541_12021# 0.0347f
C16925 _081_ net22 3.65e-20
C16926 net34 VPWR 1.22f
C16927 _104_ trim_val\[3\] 5.05e-20
C16928 a_6007_7119# a_6523_7119# 0.115f
C16929 _022_ a_3303_10217# 8.25e-19
C16930 _003_ a_6741_7361# 2.33e-20
C16931 net2 net46 1.9e-19
C16932 a_10195_1354# _117_ 0.212f
C16933 net8 a_13257_1141# 0.0163f
C16934 net15 calibrate 0.00828f
C16935 net23 a_1211_7983# 0.0015f
C16936 _110_ a_9003_3829# 0.00346f
C16937 _070_ _067_ 0.0808f
C16938 _021_ a_7477_10901# 1.27e-19
C16939 _074_ a_4959_9295# 0.00617f
C16940 a_6743_10933# a_7259_11305# 0.115f
C16941 _042_ _083_ 8.1e-20
C16942 a_7010_3311# VPWR 0.142f
C16943 clknet_0_clk a_9003_3829# 1.14e-20
C16944 _055_ trim[0] 0.0624f
C16945 net46 a_14193_3285# 0.167f
C16946 a_12992_8751# a_14467_8751# 4.14e-20
C16947 net12 a_5997_11247# 3.88e-20
C16948 a_6519_4631# a_6822_4399# 0.00145f
C16949 _107_ _058_ 4.44e-19
C16950 _065_ a_11098_6691# 0.00156f
C16951 clknet_2_0__leaf_clk a_1585_4777# 2.56e-19
C16952 a_1497_8725# VPWR 0.204f
C16953 net16 a_15023_2223# 7.09e-19
C16954 net4 a_8298_2767# 0.214f
C16955 net16 _134_ 0.335f
C16956 a_1830_10205# result[4] 2.78e-20
C16957 _065_ a_4349_8449# 7.65e-21
C16958 a_561_4405# a_1007_4777# 2.28e-19
C16959 a_911_4777# a_1476_4777# 7.99e-20
C16960 net33 _110_ 1.3e-20
C16961 clknet_0_clk a_5536_4399# 4.48e-22
C16962 net40 _029_ 0.0203f
C16963 a_5423_9011# a_6793_8970# 2.19e-20
C16964 clknet_2_2__leaf_clk a_7310_2223# 1.82e-19
C16965 _073_ VPWR 0.396f
C16966 net22 a_455_5747# 0.00146f
C16967 cal_itt\[2\] a_8307_4719# 8.54e-20
C16968 _108_ a_13607_4943# 0.042f
C16969 _002_ a_8025_8041# 0.00102f
C16970 net45 _049_ 0.00196f
C16971 mask\[7\] a_1000_11293# 8.14e-20
C16972 cal_itt\[0\] _064_ 2.64e-19
C16973 net45 a_3388_4631# 3.57e-21
C16974 _057_ a_10752_565# 4.11e-19
C16975 cal_count\[0\] a_13562_8751# 0.0475f
C16976 _040_ a_3053_8457# 7.16e-19
C16977 net3 _012_ 2.04e-20
C16978 net45 a_5699_1653# 0.33f
C16979 a_13279_8207# a_12900_7663# 8.4e-19
C16980 _085_ mask\[7\] 2e-19
C16981 _032_ _117_ 0.278f
C16982 _031_ _057_ 6.44e-20
C16983 net43 cal_itt\[2\] 0.00853f
C16984 net46 _033_ 0.176f
C16985 a_15259_7637# trimb[4] 0.00219f
C16986 _013_ a_2288_3677# 0.167f
C16987 net26 a_2953_9845# 1.99e-19
C16988 net44 a_7657_10217# 4.56e-19
C16989 _086_ ctlp[0] 1.04e-19
C16990 _048_ _087_ 0.463f
C16991 net52 net24 0.0116f
C16992 clknet_2_2__leaf_clk trim_mask\[2\] 0.59f
C16993 net24 a_816_7119# 9.84e-21
C16994 a_14981_4020# a_14540_3689# 0.00116f
C16995 net16 a_13975_3689# 0.0106f
C16996 _063_ a_8949_6031# 0.00187f
C16997 _042_ a_8360_10383# 0.0161f
C16998 _074_ a_937_3855# 0.00145f
C16999 _048_ a_6519_3829# 0.185f
C17000 net31 net46 9.91e-19
C17001 _074_ mask\[5\] 5.12e-19
C17002 a_8072_11721# a_7999_11231# 0.00189f
C17003 a_7939_10383# a_8551_10383# 0.00188f
C17004 a_8105_10383# a_9182_10749# 1.46e-19
C17005 _010_ ctlp[1] 0.00232f
C17006 a_8381_9295# _035_ 1.09e-21
C17007 a_10975_6031# a_10781_5487# 5.29e-20
C17008 _048_ _099_ 0.0926f
C17009 _119_ a_10055_2767# 0.0686f
C17010 en_co_clk a_13783_6183# 0.00143f
C17011 a_3148_4399# VPWR 0.0139f
C17012 _123_ net40 1.12e-20
C17013 VPWR ctlp[7] 0.639f
C17014 net30 a_7019_4407# 5.12e-21
C17015 net1 a_937_4105# 0.00511f
C17016 net16 a_13915_4399# 0.00719f
C17017 trim_val\[2\] a_14281_1513# 1.34e-19
C17018 a_11059_7356# a_10990_7485# 0.21f
C17019 a_6523_7119# cal_itt\[3\] 3.33e-19
C17020 net8 a_14526_1501# 4.63e-19
C17021 clknet_2_1__leaf_clk a_7916_8041# 9.63e-21
C17022 a_3365_4943# VPWR 0.00365f
C17023 cal_itt\[0\] _053_ 0.037f
C17024 a_12599_3615# a_12424_3689# 0.234f
C17025 cal_itt\[1\] a_11622_7485# 7.03e-20
C17026 a_11509_3317# _030_ 0.0025f
C17027 a_9296_9295# VPWR 0.292f
C17028 _042_ a_2450_9955# 4.96e-19
C17029 net47 a_14733_7983# 2.49e-20
C17030 clknet_0_clk a_8485_4943# 1.91e-20
C17031 _021_ a_6467_9845# 7.16e-21
C17032 _055_ a_15023_2767# 0.224f
C17033 a_561_6031# a_1007_6031# 2.28e-19
C17034 a_6743_10933# _008_ 2.16e-20
C17035 net44 net51 0.158f
C17036 mask\[4\] a_7079_10217# 0.00428f
C17037 net47 a_12756_9117# 7.37e-19
C17038 _110_ trim_val\[3\] 0.211f
C17039 state\[2\] a_4973_2773# 1.35e-19
C17040 a_455_12533# result[7] 0.0564f
C17041 net15 _018_ 0.00157f
C17042 a_4775_6031# net3 1.35e-21
C17043 net46 a_10785_1679# 0.0013f
C17044 _040_ a_4259_6031# 4.82e-21
C17045 clknet_2_0__leaf_clk _094_ 0.0325f
C17046 a_4609_9295# a_5633_9295# 2.36e-20
C17047 a_1019_4399# VPWR 0.138f
C17048 a_7351_8041# a_7256_8029# 0.0498f
C17049 a_7569_7637# a_7447_8041# 3.16e-19
C17050 clknet_2_2__leaf_clk a_9719_1473# 8.39e-22
C17051 _021_ VPWR 0.367f
C17052 state\[0\] a_4973_2773# 0.00443f
C17053 a_6541_12021# a_6987_12393# 2.28e-19
C17054 _101_ a_2869_10927# 0.0603f
C17055 net41 cal 0.0709f
C17056 _132_ a_14564_6397# 8.94e-20
C17057 net54 state\[2\] 0.00408f
C17058 a_8583_3317# _025_ 2.56e-21
C17059 a_3615_8207# _077_ 3.13e-20
C17060 a_3781_8207# a_5535_8181# 2.58e-19
C17061 net33 a_14564_6397# 0.0027f
C17062 a_4349_8449# a_4696_8207# 0.0512f
C17063 _033_ a_11149_3017# 6.44e-20
C17064 a_15299_6575# VPWR 0.283f
C17065 _108_ a_11488_4765# 9.48e-19
C17066 net54 state\[0\] 0.126f
C17067 net14 calibrate 0.0958f
C17068 mask\[1\] _005_ 2.2e-19
C17069 _069_ a_9460_6807# 5.64e-21
C17070 a_2953_7119# _049_ 0.00111f
C17071 a_2877_2197# ctln[1] 2.4e-20
C17072 _064_ trim_mask\[0\] 0.46f
C17073 cal_count\[3\] VPWR 2.99f
C17074 a_6793_8970# _076_ 0.212f
C17075 net19 _092_ 0.00741f
C17076 net55 a_8307_4719# 0.00894f
C17077 net51 en_co_clk 1.77e-19
C17078 net37 comp 8.58e-19
C17079 net44 _003_ 0.00554f
C17080 a_6885_8372# a_6835_7669# 8.38e-19
C17081 a_579_12021# _086_ 0.00916f
C17082 _011_ a_448_11445# 0.00178f
C17083 a_6891_12393# a_7456_12393# 7.99e-20
C17084 net18 a_11292_1251# 0.00254f
C17085 mask\[4\] a_7723_10143# 0.0672f
C17086 a_8022_7119# a_9460_6807# 0.011f
C17087 mask\[3\] a_763_8757# 1.75e-19
C17088 _136_ _110_ 5.58e-19
C17089 a_2283_4020# a_1867_3317# 9.84e-19
C17090 a_14249_8725# a_14199_7369# 2.3e-21
C17091 a_6703_2197# a_6941_2589# 0.0074f
C17092 a_4655_10071# _019_ 0.117f
C17093 cal_count\[3\] a_12218_6397# 4.21e-19
C17094 _048_ a_5537_4943# 0.00218f
C17095 net47 a_11059_7356# 0.153f
C17096 net13 _094_ 0.0763f
C17097 net43 net55 0.00162f
C17098 _100_ a_5537_4105# 0.00279f
C17099 _001_ a_11622_7485# 0.177f
C17100 a_12586_3311# VPWR 4.98e-19
C17101 net15 mask\[1\] 0.00484f
C17102 _108_ _113_ 9.94e-20
C17103 _063_ _062_ 0.322f
C17104 mask\[0\] a_911_6031# 2.09e-20
C17105 net13 a_4043_10143# 0.0043f
C17106 _074_ _039_ 4.18e-20
C17107 _105_ _104_ 8.7e-20
C17108 clknet_2_2__leaf_clk a_9595_1679# 0.247f
C17109 _101_ net53 0.0933f
C17110 net33 a_13091_4943# 7.1e-21
C17111 clknet_2_0__leaf_clk a_2787_7119# 0.854f
C17112 a_14981_8235# VPWR 4.87e-19
C17113 net4 net6 0.0663f
C17114 a_4259_6031# _048_ 1.76e-20
C17115 a_3339_2767# a_3933_2767# 1.28e-19
C17116 net12 a_6056_8359# 0.0113f
C17117 _074_ net43 0.0394f
C17118 a_1644_12533# mask\[7\] 1.67e-19
C17119 net29 a_1660_12393# 0.0124f
C17120 net27 ctlp[7] 1.3e-20
C17121 a_6316_5193# _107_ 0.00144f
C17122 _106_ a_7527_4631# 5.89e-20
C17123 a_455_3571# a_2033_3317# 9.62e-20
C17124 net26 mask\[3\] 0.00358f
C17125 _120_ a_4425_6031# 9.35e-20
C17126 a_1461_10357# net25 8.35e-19
C17127 cal_itt\[1\] _092_ 0.00235f
C17128 net40 trim_mask\[1\] 8.96e-22
C17129 _136_ a_10699_5487# 0.0986f
C17130 _136_ a_12148_4777# 0.00119f
C17131 _003_ clk 2.86e-19
C17132 _055_ a_15299_3311# 0.197f
C17133 a_15259_7637# _130_ 0.0114f
C17134 _104_ a_7010_3311# 0.0789f
C17135 _003_ en_co_clk 9.3e-20
C17136 _012_ valid 0.0086f
C17137 net52 a_4677_7882# 0.0406f
C17138 _096_ a_4863_4917# 0.00268f
C17139 net19 cal_itt\[3\] 4.96e-20
C17140 a_13562_8751# a_13919_8751# 2.69e-19
C17141 a_12992_8751# a_14249_8725# 1.08e-19
C17142 a_13142_8725# net40 4.04e-20
C17143 a_8078_7663# VPWR 5.12e-19
C17144 net46 a_14083_3311# 0.0122f
C17145 net14 a_1461_10357# 0.00317f
C17146 cal_itt\[2\] a_8270_8029# 8.36e-19
C17147 _053_ trim_mask\[0\] 0.396f
C17148 a_3868_10217# _008_ 1.37e-20
C17149 _102_ a_2869_10927# 6.74e-19
C17150 _002_ a_6173_7119# 0.00792f
C17151 a_8912_2589# a_9103_2601# 4.61e-19
C17152 a_9195_10357# _043_ 0.0167f
C17153 mask\[4\] a_8717_10383# 2.83e-19
C17154 _097_ a_2309_2229# 4.42e-21
C17155 a_11067_4405# a_11067_3017# 2.01e-21
C17156 net43 a_1279_9129# 0.157f
C17157 a_7939_10383# a_9871_10383# 1.06e-20
C17158 a_6173_7119# _050_ 1.23e-21
C17159 _049_ a_6316_5193# 0.00562f
C17160 net13 a_2787_7119# 1.88e-21
C17161 a_2689_8751# clknet_2_0__leaf_clk 1.88e-20
C17162 a_10405_9295# _053_ 1.27e-21
C17163 state\[2\] a_7019_4407# 0.166f
C17164 _049_ a_2857_5461# 0.0271f
C17165 a_561_4405# net41 2.66e-21
C17166 mask\[7\] a_2828_12131# 0.188f
C17167 a_1660_12393# a_3431_12021# 1.43e-20
C17168 net1 a_2479_3689# 7.19e-21
C17169 a_1467_7923# a_561_7119# 0.00553f
C17170 a_4655_10071# VPWR 0.288f
C17171 a_8673_10625# net47 0.166f
C17172 a_2857_5461# a_3388_4631# 8.03e-19
C17173 a_7010_3311# a_7200_3631# 0.0119f
C17174 a_911_6031# _079_ 4.49e-19
C17175 net54 _100_ 0.0442f
C17176 state\[2\] a_4471_4007# 5.29e-21
C17177 _122_ a_13470_7663# 0.00134f
C17178 _014_ a_2283_4020# 0.00786f
C17179 net45 sample 4.04e-20
C17180 net19 a_9317_3285# 6.83e-19
C17181 net45 trim_mask\[4\] 0.103f
C17182 _051_ a_8583_3317# 5.67e-19
C17183 _065_ net2 1.15f
C17184 cal_itt\[1\] cal_itt\[3\] 0.00338f
C17185 net25 _018_ 0.00104f
C17186 a_8298_2767# a_9007_2601# 0.00978f
C17187 a_4871_8181# net30 4.43e-21
C17188 _058_ trim_mask\[4\] 0.134f
C17189 _093_ a_2601_3285# 8.41e-20
C17190 a_3667_3829# state\[1\] 2.13e-19
C17191 state\[0\] a_4471_4007# 0.0209f
C17192 _076_ net30 0.0106f
C17193 net16 trim_val\[1\] 0.0116f
C17194 a_1095_12393# a_1493_11721# 9.8e-19
C17195 _022_ a_2869_10927# 0.00252f
C17196 net50 clknet_2_2__leaf_clk 0.0136f
C17197 net14 _018_ 9.06e-21
C17198 _134_ clkc 2.48e-19
C17199 a_8657_2229# a_9115_2223# 0.0346f
C17200 a_9463_8725# VPWR 0.339f
C17201 a_4055_10927# _042_ 4.99e-19
C17202 _111_ _109_ 9.95e-19
C17203 net13 a_4617_3855# 1.99e-19
C17204 net55 a_6822_4399# 0.00129f
C17205 net4 a_9529_6059# 7.2e-19
C17206 a_10990_7485# a_11016_6691# 1.96e-20
C17207 a_8022_7119# a_8495_6895# 0.00413f
C17208 clknet_2_0__leaf_clk a_7088_7119# 6.95e-20
C17209 a_14564_6397# _136_ 1.66e-19
C17210 a_13111_6031# a_13193_6031# 0.00369f
C17211 a_3521_7361# VPWR 0.225f
C17212 cal_count\[2\] a_13142_7271# 0.0138f
C17213 _063_ a_8745_6895# 0.0185f
C17214 _042_ _000_ 1.3e-20
C17215 a_9020_10383# a_8731_9295# 3.42e-20
C17216 trim_val\[4\] a_10270_4105# 8.47e-19
C17217 clknet_0_clk _105_ 0.0125f
C17218 a_11394_9509# a_11814_9295# 0.144f
C17219 a_561_9845# _082_ 0.00178f
C17220 trim_mask\[0\] a_14335_4020# 2.87e-20
C17221 net9 a_13111_6031# 0.00155f
C17222 a_14807_8359# a_14981_8235# 0.00658f
C17223 net2 a_9761_8457# 3.07e-19
C17224 clknet_2_1__leaf_clk a_448_11445# 0.0124f
C17225 a_745_12021# result[7] 0.0012f
C17226 a_7223_2465# clk 0.0236f
C17227 a_1129_7361# VPWR 0.227f
C17228 net24 _065_ 3.63e-21
C17229 a_14347_4917# VPWR 0.37f
C17230 a_6375_12021# net53 1.2e-19
C17231 _062_ a_5455_4943# 0.14f
C17232 a_7164_11293# a_7355_11305# 4.61e-19
C17233 a_745_10933# net25 1.29e-19
C17234 a_10543_2455# a_11435_2229# 7.3e-21
C17235 a_9572_2601# a_11601_2229# 1.79e-21
C17236 _024_ trim_mask\[1\] 1.13e-19
C17237 net14 mask\[1\] 0.00984f
C17238 _096_ a_3817_4697# 0.247f
C17239 a_14249_8725# a_14422_7093# 9.18e-21
C17240 a_1095_12393# VPWR 0.209f
C17241 mask\[5\] _083_ 0.00101f
C17242 _048_ a_7393_5193# 0.0011f
C17243 _136_ a_13091_4943# 0.00475f
C17244 net3 a_3933_2767# 0.0394f
C17245 net24 net23 3.22e-19
C17246 net14 a_745_10933# 0.00884f
C17247 a_1099_12533# a_1313_10901# 2.73e-21
C17248 _119_ VPWR 0.494f
C17249 _053_ a_8949_6281# 2.12e-19
C17250 a_1638_9839# VPWR 5.57e-19
C17251 a_11258_9117# VPWR 9.7e-20
C17252 net4 a_9369_4105# 0.00558f
C17253 a_15023_10927# trimb[1] 6.66e-20
C17254 a_2019_9055# a_2143_7663# 1.68e-20
C17255 net28 a_1660_12393# 1.46e-19
C17256 trim_mask\[2\] a_14335_2442# 0.053f
C17257 clknet_2_0__leaf_clk _096_ 0.00191f
C17258 _071_ a_9043_6031# 6.01e-19
C17259 _101_ a_6007_9839# 2.38e-19
C17260 net22 a_395_4405# 2.45e-20
C17261 a_11244_9661# _123_ 6.77e-19
C17262 net11 ctln[6] 6.71e-19
C17263 cal_count\[3\] _104_ 1.88e-20
C17264 net45 a_3123_3615# 0.275f
C17265 net47 a_11016_6691# 0.00446f
C17266 clknet_0_clk _073_ 5.34e-22
C17267 a_561_7119# a_2787_7119# 8.25e-20
C17268 net19 a_9003_3829# 0.0147f
C17269 trim_mask\[2\] net8 0.0279f
C17270 net25 a_1387_8751# 1.1e-19
C17271 net46 a_13715_5309# 0.0388f
C17272 net40 a_14335_7895# 0.015f
C17273 a_11801_4373# a_12310_4399# 2.6e-19
C17274 calibrate a_6927_3311# 0.0157f
C17275 _100_ a_4471_4007# 0.0743f
C17276 net43 _034_ 0.021f
C17277 a_9084_4515# a_9099_3689# 1.1e-20
C17278 mask\[1\] a_395_7119# 3.15e-20
C17279 a_7631_12319# a_8072_11721# 3.24e-19
C17280 a_561_9845# a_1007_10217# 2.28e-19
C17281 a_7527_4631# _054_ 5.12e-20
C17282 net44 net26 0.0747f
C17283 net14 a_1387_8751# 0.00184f
C17284 net9 a_11814_9295# 0.00333f
C17285 _078_ a_4349_8449# 1.24e-19
C17286 a_6566_5193# VPWR 0.183f
C17287 a_14972_5193# trim[1] 2.18e-19
C17288 a_6210_4989# _107_ 0.00576f
C17289 a_8381_9295# a_9296_9295# 0.125f
C17290 _095_ VPWR 0.976f
C17291 _064_ a_8298_2767# 2.53e-20
C17292 mask\[4\] _042_ 0.0476f
C17293 _074_ a_1173_6031# 6.43e-19
C17294 net44 a_5050_8207# 0.00331f
C17295 a_816_7119# result[1] 6.45e-20
C17296 net15 _010_ 0.00749f
C17297 clknet_2_1__leaf_clk a_3431_10933# 0.253f
C17298 _048_ a_9503_4399# 0.00146f
C17299 clknet_2_3__leaf_clk net30 3.13e-21
C17300 _074_ a_2953_9845# 1.2e-19
C17301 clknet_2_1__leaf_clk a_929_8757# 0.00269f
C17302 a_4775_6031# net54 1.26e-21
C17303 _128_ a_13279_8207# 0.00844f
C17304 net44 a_7262_5461# 3.35e-21
C17305 net2 _067_ 3.42e-19
C17306 _123_ a_13349_6031# 1.36e-19
C17307 a_8307_6575# a_8298_5487# 0.00108f
C17308 a_10383_7093# VPWR 0.389f
C17309 net13 _096_ 0.649f
C17310 a_911_4777# _014_ 4.82e-21
C17311 a_7916_8041# cal_itt\[3\] 4.63e-19
C17312 a_14377_9545# trimb[1] 5.07e-19
C17313 trim_val\[0\] a_13519_4007# 1.89e-21
C17314 _119_ a_9478_4105# 3.48e-19
C17315 _049_ a_6210_4989# 0.00157f
C17316 _053_ a_8307_4943# 0.111f
C17317 trim_mask\[3\] a_9761_1679# 0.00315f
C17318 a_10055_2767# a_10111_1679# 1.78e-19
C17319 a_10655_2932# a_10329_1921# 1.36e-21
C17320 mask\[3\] a_2961_9295# 0.00178f
C17321 net9 a_13825_6031# 9.99e-20
C17322 a_14347_9480# cal_count\[1\] 4.78e-21
C17323 _087_ a_6197_4399# 0.00257f
C17324 net53 a_7824_11305# 1.86e-21
C17325 trim_val\[2\] a_14184_1679# 3.41e-19
C17326 a_13783_6183# _108_ 1.67e-20
C17327 _106_ clknet_2_2__leaf_clk 1.18e-19
C17328 _045_ _084_ 0.0144f
C17329 net20 _042_ 1.83e-22
C17330 a_4995_7119# a_6007_7119# 3.47e-21
C17331 _088_ clk 8.97e-20
C17332 _121_ _120_ 0.00179f
C17333 _131_ en_co_clk 0.00178f
C17334 en_co_clk _088_ 9.79e-21
C17335 _127_ _126_ 0.0402f
C17336 _070_ a_7001_7669# 2.92e-20
C17337 a_11679_4777# VPWR 5.1e-19
C17338 a_1095_12393# net27 9.2e-20
C17339 a_7262_5461# clk 0.0122f
C17340 cal_itt\[1\] a_9602_6941# 1.04e-19
C17341 net9 a_11067_3017# 6.46e-19
C17342 en_co_clk a_7262_5461# 4.84e-21
C17343 _053_ a_8298_2767# 4.79e-19
C17344 net46 a_12599_3615# 0.347f
C17345 a_11987_8757# a_14467_8751# 3.38e-20
C17346 _037_ a_12231_6005# 9.46e-20
C17347 net12 a_7310_2223# 7.17e-20
C17348 a_1313_10901# a_1357_11293# 3.69e-19
C17349 net13 a_4209_11293# 1.81e-19
C17350 a_1095_11305# a_1191_11305# 0.0138f
C17351 a_6099_10633# a_6633_9845# 3.43e-19
C17352 a_745_10933# a_1769_11305# 2.36e-20
C17353 _099_ a_6197_4399# 0.0113f
C17354 _029_ trim_mask\[1\] 5.78e-21
C17355 a_13562_8751# cal_count\[2\] 8.14e-20
C17356 clknet_2_2__leaf_clk a_14193_3285# 1.54e-20
C17357 _101_ a_5363_7369# 0.17f
C17358 _050_ a_7800_4631# 1.83e-20
C17359 a_7617_2589# VPWR 5.66e-20
C17360 _051_ a_5625_4943# 2.74e-19
C17361 a_12723_4943# _058_ 0.00368f
C17362 trim_mask\[3\] a_10787_1135# 0.059f
C17363 a_5423_9011# a_5691_7637# 1.96e-19
C17364 mask\[6\] a_4512_11305# 0.0417f
C17365 _053_ a_7210_5807# 1.94e-19
C17366 a_5686_2045# clk 3.55e-19
C17367 net55 a_4617_4105# 0.0477f
C17368 net19 trim_val\[3\] 5.82e-23
C17369 net45 a_1173_4765# 0.00316f
C17370 a_9572_2601# a_10016_1679# 2.39e-19
C17371 _048_ _097_ 0.0686f
C17372 cal_count\[3\] _110_ 4.11e-20
C17373 a_14172_1513# a_14471_591# 0.00177f
C17374 a_8673_10625# _068_ 1.5e-21
C17375 a_10864_9269# _041_ 1.13e-19
C17376 a_395_591# rstn 0.195f
C17377 net46 a_12257_4777# 8.19e-19
C17378 cal_count\[0\] _036_ 0.083f
C17379 _042_ a_2815_9447# 0.0322f
C17380 a_11491_6031# a_12056_6031# 7.99e-20
C17381 net37 a_12992_8751# 4.63e-21
C17382 _082_ _006_ 0.00503f
C17383 clknet_2_3__leaf_clk _134_ 0.0566f
C17384 net34 a_13091_4943# 2.82e-21
C17385 a_579_12021# _046_ 6.7e-21
C17386 cal_itt\[3\] a_7442_7119# 6.42e-19
C17387 clknet_0_clk cal_count\[3\] 1.76e-20
C17388 _011_ a_1203_12015# 0.00105f
C17389 net43 net4 2.72e-21
C17390 net18 _041_ 0.00946f
C17391 a_6909_10933# mask\[4\] 1.34e-20
C17392 clknet_2_2__leaf_clk _033_ 0.759f
C17393 trim_mask\[0\] a_9664_3689# 5.1e-20
C17394 net16 a_14184_2767# 4.9e-19
C17395 net16 a_15023_10927# 3.37e-19
C17396 clknet_2_1__leaf_clk a_7999_11231# 9.42e-19
C17397 net46 a_8912_2589# 2.46e-19
C17398 a_6099_10633# a_6445_10383# 0.0134f
C17399 _108_ a_10975_4105# 1.48e-19
C17400 a_9225_2197# VPWR 0.209f
C17401 a_4866_11293# VPWR 1.68e-19
C17402 net43 a_3303_7119# 0.153f
C17403 net15 _050_ 3.54e-20
C17404 net12 _090_ 0.0052f
C17405 _046_ a_2869_10927# 1.51e-19
C17406 cal_count\[3\] a_10699_5487# 0.0968f
C17407 clknet_2_1__leaf_clk clknet_2_0__leaf_clk 0.028f
C17408 _123_ a_13142_8725# 0.0138f
C17409 a_15023_1679# a_14931_591# 1.77e-20
C17410 cal_itt\[0\] a_9919_6614# 0.00591f
C17411 _002_ a_7351_8041# 0.0364f
C17412 trim_val\[2\] _057_ 5.23e-20
C17413 a_8949_6031# _092_ 0.00314f
C17414 a_816_10205# net24 2.92e-21
C17415 net43 a_911_7119# 0.156f
C17416 a_6007_7119# a_6619_7119# 0.00188f
C17417 _058_ a_11967_3311# 5.41e-19
C17418 _005_ a_561_6031# 4.58e-20
C17419 _065_ a_4993_6273# 8.96e-21
C17420 a_1129_6273# a_1019_6397# 0.0977f
C17421 a_10195_1354# _116_ 0.0372f
C17422 a_13825_1109# a_14172_1513# 0.0512f
C17423 a_13257_1141# a_15023_1135# 2.12e-19
C17424 _104_ _119_ 0.103f
C17425 a_8215_9295# VPWR 0.49f
C17426 net20 a_6909_10933# 5.31e-21
C17427 _025_ a_11859_3689# 6.4e-19
C17428 a_11343_3317# a_12599_3615# 0.0435f
C17429 net9 a_12992_8751# 7.41e-19
C17430 a_929_8757# a_1953_9129# 2.36e-20
C17431 a_745_12021# mask\[7\] 5.51e-19
C17432 clknet_2_1__leaf_clk a_4687_12319# 0.0609f
C17433 a_1313_11989# a_1660_12393# 0.0512f
C17434 _074_ mask\[3\] 0.116f
C17435 net43 a_1835_12319# 0.281f
C17436 a_8381_9295# a_9463_8725# 2.48e-19
C17437 a_10005_6031# a_10975_6031# 4.77e-19
C17438 a_9443_6059# a_11141_6031# 6.55e-21
C17439 a_763_8757# a_1184_9117# 0.0931f
C17440 net35 _058_ 0.00401f
C17441 net37 a_15111_9295# 0.00147f
C17442 a_13059_4631# _058_ 0.00906f
C17443 net46 a_10543_2455# 0.00358f
C17444 _053_ a_12344_8041# 5.85e-20
C17445 _120_ a_3273_4943# 0.0845f
C17446 calibrate VPWR 4.54f
C17447 _095_ a_2383_3689# 4.5e-19
C17448 net18 a_10781_5487# 0.0044f
C17449 net43 a_2450_9955# 3.43e-19
C17450 a_1493_11721# a_1461_10357# 1.29e-21
C17451 _053_ a_5177_1921# 8.36e-20
C17452 _059_ _088_ 7.29e-21
C17453 net16 net47 7.59e-20
C17454 net16 a_14377_9545# 0.00445f
C17455 net44 cal_itt\[2\] 4.51e-19
C17456 a_13470_7663# a_13111_6031# 6.18e-20
C17457 _101_ _102_ 0.00317f
C17458 clknet_2_1__leaf_clk net13 7.95e-20
C17459 net15 a_3615_8207# 4.44e-21
C17460 cal_count\[2\] _131_ 0.643f
C17461 _103_ a_7677_4759# 2.7e-19
C17462 mask\[3\] a_1279_9129# 0.00691f
C17463 _040_ a_6056_8359# 1.12e-19
C17464 _017_ a_5535_8181# 7.14e-22
C17465 _032_ _116_ 0.0668f
C17466 a_13562_8751# cal_count\[1\] 0.0975f
C17467 _041_ a_11575_8790# 3.12e-19
C17468 a_4815_3031# a_4901_2773# 0.0049f
C17469 trim_mask\[3\] a_11067_3017# 0.0609f
C17470 net26 a_8992_9955# 0.104f
C17471 _071_ a_8935_6895# 6.61e-21
C17472 net40 _066_ 4.32e-20
C17473 a_448_11445# result[4] 1.02e-19
C17474 _035_ _001_ 1.09e-19
C17475 a_4696_8207# a_4677_7882# 2e-19
C17476 a_6523_7119# _073_ 9.17e-19
C17477 a_14715_3615# a_15023_2223# 9.71e-21
C17478 net9 a_11856_2589# 0.00125f
C17479 _076_ a_5691_7637# 0.0222f
C17480 a_9463_8725# clknet_0_clk 3.52e-21
C17481 a_6793_8970# a_6835_7669# 6.02e-20
C17482 _093_ a_4617_4105# 0.00354f
C17483 net29 a_1095_11305# 1.9e-19
C17484 _078_ net2 6.06e-20
C17485 cal_itt\[2\] clk 0.0131f
C17486 net17 a_12631_12559# 0.174f
C17487 cal_itt\[2\] en_co_clk 0.253f
C17488 a_11292_1251# VPWR 0.171f
C17489 _101_ _022_ 0.0144f
C17490 a_1461_10357# VPWR 0.226f
C17491 a_1651_4703# valid 1.44e-19
C17492 _051_ _103_ 0.0432f
C17493 cal_itt\[2\] a_8386_8457# 2.25e-19
C17494 a_2857_7637# a_3303_7119# 0.0132f
C17495 clknet_0_clk a_3521_7361# 0.00127f
C17496 mask\[5\] _000_ 1.37e-19
C17497 _092_ a_4863_4917# 0.0527f
C17498 a_9761_1679# a_10207_1679# 2.28e-19
C17499 a_10329_1921# a_10838_2045# 2.6e-19
C17500 net37 _132_ 0.00591f
C17501 a_8298_5487# VPWR 1.25f
C17502 _001_ _136_ 0.00119f
C17503 a_6619_7119# cal_itt\[3\] 2.69e-19
C17504 _136_ a_11067_4405# 0.00263f
C17505 net51 _049_ 0.00338f
C17506 a_12900_7663# a_13142_7271# 0.00129f
C17507 _030_ a_15299_3311# 1.16e-20
C17508 a_14193_3285# a_14540_3689# 0.0512f
C17509 a_13625_3317# _055_ 1.23e-19
C17510 a_12153_8757# _041_ 0.275f
C17511 a_12436_9129# a_12992_8751# 0.00329f
C17512 mask\[2\] a_3840_8867# 0.201f
C17513 a_11987_8757# a_14249_8725# 5.65e-20
C17514 _036_ a_13919_8751# 6.61e-21
C17515 _015_ a_4959_1679# 9.18e-19
C17516 net33 net37 0.841f
C17517 _062_ _092_ 0.0592f
C17518 _006_ net22 7.26e-21
C17519 cal_itt\[1\] a_10861_7119# 1.09e-19
C17520 a_3303_10217# a_3868_10217# 7.99e-20
C17521 net16 a_14686_2339# 3.12e-19
C17522 a_7256_8029# VPWR 0.0851f
C17523 mask\[2\] a_2971_8457# 0.112f
C17524 _019_ mask\[1\] 2.67e-20
C17525 cal_itt\[0\] _124_ 7.19e-19
C17526 net46 a_13607_1513# 0.177f
C17527 net19 _105_ 0.0167f
C17528 _110_ _119_ 0.00786f
C17529 net23 result[1] 0.00612f
C17530 clknet_2_3__leaf_clk a_9458_9661# 3.05e-19
C17531 a_10111_1679# VPWR 0.212f
C17532 _076_ a_4775_6031# 1.22e-19
C17533 clknet_0_clk _119_ 0.0394f
C17534 a_15083_4659# trim[0] 1.44e-19
C17535 a_6191_12559# VPWR 0.277f
C17536 _078_ net24 0.506f
C17537 trim_mask\[1\] a_8749_3317# 0.00141f
C17538 a_5915_11721# a_5998_11471# 2.42e-19
C17539 a_1493_11721# a_745_10933# 4.52e-20
C17540 _018_ VPWR 0.477f
C17541 _020_ a_7939_10383# 0.288f
C17542 net47 a_10593_9295# 0.0215f
C17543 net16 net5 3.66e-20
C17544 a_13257_4943# _058_ 0.00777f
C17545 a_13825_5185# a_13697_4373# 3.19e-19
C17546 _084_ _078_ 0.00638f
C17547 a_8083_8181# _072_ 0.171f
C17548 _122_ _037_ 0.00898f
C17549 net44 a_4858_8573# 1.7e-19
C17550 net44 net55 0.00485f
C17551 _003_ _049_ 1.6e-19
C17552 _016_ a_3208_7119# 0.157f
C17553 _108_ a_9099_3689# 4.04e-19
C17554 _068_ a_8083_8181# 0.00218f
C17555 _097_ a_2033_3317# 0.00178f
C17556 _065_ a_11059_7356# 0.00211f
C17557 _022_ _102_ 1.9e-20
C17558 cal_itt\[3\] _062_ 2.91e-19
C17559 a_2787_7119# _094_ 3.12e-21
C17560 net15 a_3249_9295# 9.36e-19
C17561 net31 a_14540_3689# 0.00298f
C17562 _028_ a_7181_2589# 1.84e-19
C17563 cal_count\[1\] _131_ 1.02e-20
C17564 a_14335_2442# a_14604_2339# 0.0215f
C17565 cal_itt\[1\] _105_ 4.25e-19
C17566 a_7310_2223# a_7524_2223# 0.0977f
C17567 a_8298_5487# a_9478_4105# 2.91e-21
C17568 net14 a_561_6031# 0.0105f
C17569 net46 a_13881_1653# 0.00853f
C17570 cal_itt\[2\] a_8091_7967# 0.0914f
C17571 _074_ a_4687_11231# 0.00417f
C17572 mask\[5\] mask\[4\] 0.071f
C17573 a_6835_7669# net30 4.23e-20
C17574 _053_ a_9529_6059# 4.01e-19
C17575 net16 a_14347_1439# 0.00492f
C17576 _104_ a_9225_2197# 3.01e-20
C17577 clknet_0_clk _095_ 0.166f
C17578 _135_ VPWR 0.394f
C17579 _074_ net44 0.137f
C17580 a_14788_7369# comp 1.28e-19
C17581 a_3947_12393# a_4055_12015# 0.0572f
C17582 a_4471_4007# a_3933_2767# 0.0011f
C17583 a_4687_12319# a_4866_12381# 0.0074f
C17584 a_4512_12393# a_4621_12393# 0.00742f
C17585 state\[1\] a_3339_2767# 0.0119f
C17586 a_13869_1501# VPWR 0.0022f
C17587 en_co_clk a_5081_4943# 0.00145f
C17588 clknet_2_0__leaf_clk a_6007_7119# 0.248f
C17589 net43 a_4055_10927# 0.0173f
C17590 a_9664_3689# a_8298_2767# 0.00155f
C17591 a_9839_3615# a_10055_2767# 0.0114f
C17592 a_10781_5487# a_11023_5108# 1.6e-19
C17593 a_10055_5487# _108_ 5.02e-19
C17594 a_448_11445# a_448_10357# 0.00269f
C17595 a_7902_10205# VPWR 7.21e-20
C17596 mask\[1\] VPWR 2.43f
C17597 net55 clk 0.00591f
C17598 en_co_clk net55 0.0459f
C17599 a_8455_10383# a_8215_9295# 1.92e-20
C17600 a_745_10933# VPWR 0.589f
C17601 trim_mask\[1\] _115_ 1.95e-19
C17602 a_12077_3285# a_12121_3677# 3.69e-19
C17603 a_11509_3317# a_12533_3689# 2.36e-20
C17604 trim_mask\[3\] a_11856_2589# 8.81e-19
C17605 a_4866_12381# net13 3.89e-20
C17606 trim_mask\[2\] trim[2] 1.25e-19
C17607 a_10239_9295# a_11244_9661# 0.183f
C17608 _092_ a_3817_4697# 3.2e-21
C17609 _035_ a_11394_9509# 1.83e-21
C17610 a_14193_3285# a_14335_2442# 2.09e-20
C17611 a_395_7119# a_561_6031# 1.21e-19
C17612 net55 a_9084_4515# 5.3e-21
C17613 a_14236_8457# trimb[4] 1.71e-19
C17614 _027_ a_11435_2229# 2.54e-19
C17615 cal_itt\[1\] _073_ 4.66e-20
C17616 a_3303_10217# a_3399_10217# 0.0138f
C17617 a_11141_6031# a_11396_6031# 0.0564f
C17618 calibrate _104_ 0.145f
C17619 trim_val\[0\] a_14526_4943# 1.25e-19
C17620 _090_ a_5691_2741# 1.39e-20
C17621 net28 a_1095_11305# 7.67e-20
C17622 a_5496_12131# a_6541_12021# 1.03e-20
C17623 net20 mask\[5\] 0.0649f
C17624 net52 a_2961_9545# 0.0105f
C17625 a_10752_12533# ctlp[4] 0.168f
C17626 _078_ a_5878_9295# 5.11e-19
C17627 net46 a_14334_1135# 2.06e-19
C17628 a_14379_6397# a_14172_4943# 0.00112f
C17629 a_14564_6397# a_14347_4917# 4.47e-19
C17630 a_15083_4659# a_15023_2767# 1.88e-19
C17631 _053_ a_9369_4105# 1.27e-20
C17632 net22 a_911_4777# 8.02e-19
C17633 mask\[2\] a_4131_8207# 3.55e-19
C17634 _127_ VPWR 0.264f
C17635 clknet_2_3__leaf_clk _118_ 5.75e-20
C17636 clknet_2_0__leaf_clk _092_ 0.144f
C17637 net20 a_6999_12015# 0.00219f
C17638 a_1660_11305# net52 9.47e-19
C17639 a_6191_12559# net27 3.71e-20
C17640 a_1387_8751# VPWR 0.134f
C17641 cal_count\[0\] net4 2.07e-19
C17642 _015_ VPWR 0.564f
C17643 trim_val\[4\] a_9802_4007# 0.085f
C17644 a_1129_7361# a_1007_7119# 3.16e-19
C17645 a_9099_3689# a_9004_3677# 0.0498f
C17646 a_9317_3285# a_9195_3689# 3.16e-19
C17647 net19 a_9296_9295# 0.00455f
C17648 a_11709_6273# net46 0.162f
C17649 a_7715_3285# clk 0.0154f
C17650 net52 mask\[0\] 6.74e-19
C17651 _078_ a_1129_6273# 0.00235f
C17652 a_14063_7093# VPWR 0.207f
C17653 trim_mask\[2\] a_12169_2197# 2.59e-19
C17654 _035_ a_11116_8983# 1.97e-19
C17655 a_10239_9295# _123_ 0.0015f
C17656 a_10405_9295# _124_ 1.13e-19
C17657 a_10864_9269# a_10747_8970# 7.07e-19
C17658 net37 _136_ 2.66e-20
C17659 a_13519_4007# VPWR 0.25f
C17660 _047_ a_15023_2223# 4.2e-22
C17661 clknet_2_1__leaf_clk a_7631_12319# 3.11e-20
C17662 _041_ a_13050_7637# 4.68e-21
C17663 a_11801_4373# a_11845_4765# 3.69e-19
C17664 calibrate a_7200_3631# 0.00602f
C17665 _063_ a_9621_8029# 1.28e-19
C17666 a_12992_8751# a_13470_7663# 1.29e-19
C17667 a_11233_4405# a_12257_4777# 2.36e-20
C17668 net16 a_15023_12015# 0.00105f
C17669 net18 a_10747_8970# 2.08e-19
C17670 _049_ a_7223_2465# 2.8e-20
C17671 _108_ trim_val\[4\] 0.299f
C17672 a_7800_4631# a_7891_3617# 1.68e-19
C17673 _107_ a_9099_3689# 0.00213f
C17674 net9 trim_val\[3\] 4.6e-19
C17675 mask\[3\] _083_ 6.93e-20
C17676 a_13091_4943# a_14347_4917# 0.0427f
C17677 a_13257_4943# a_13607_4943# 0.21f
C17678 a_5524_9295# net51 3.81e-20
C17679 a_6796_12381# VPWR 0.0824f
C17680 a_11601_2229# a_12625_2601# 2.36e-20
C17681 a_12169_2197# a_12213_2589# 3.69e-19
C17682 net45 a_6941_2589# 0.00288f
C17683 net45 a_1493_5487# 0.00159f
C17684 a_8215_9295# a_8381_9295# 0.584f
C17685 _048_ a_4308_4917# 0.0203f
C17686 net13 _092_ 0.0585f
C17687 a_13059_4631# _113_ 6.11e-20
C17688 cal_itt\[3\] a_8745_6895# 8.18e-20
C17689 clknet_2_1__leaf_clk a_9020_10383# 6.95e-20
C17690 _136_ a_13193_6031# 0.00104f
C17691 a_9296_9295# cal_itt\[1\] 1.16e-20
C17692 _129_ trimb[4] 0.00203f
C17693 net2 a_7001_7669# 1.92e-19
C17694 _110_ a_9225_2197# 2.26e-19
C17695 _062_ a_5547_5603# 0.00558f
C17696 net16 net46 0.0561f
C17697 a_10055_5487# _107_ 5.69e-20
C17698 a_8298_5487# _104_ 1.77e-19
C17699 net19 cal_count\[3\] 0.00666f
C17700 net43 mask\[4\] 2.88e-19
C17701 net44 a_8636_9295# 4.4e-19
C17702 a_14604_3017# VPWR 0.156f
C17703 a_561_9845# a_1476_10217# 0.117f
C17704 _050_ a_7460_5807# 0.0867f
C17705 _060_ a_4498_4373# 0.0107f
C17706 _060_ a_4864_1679# 3.19e-20
C17707 net27 a_745_10933# 3.19e-20
C17708 a_14715_3615# trim_val\[1\] 0.103f
C17709 _059_ a_5081_4943# 1.17e-19
C17710 _062_ a_9003_3829# 1.82e-19
C17711 net9 _136_ 0.0501f
C17712 a_395_9845# a_1129_9813# 0.0701f
C17713 net10 a_12631_591# 3.69e-20
C17714 a_4680_6031# a_4871_6031# 4.61e-19
C17715 _007_ a_561_9845# 0.252f
C17716 a_14981_4020# trim[1] 6.46e-19
C17717 calibrate a_1007_4777# 2.29e-19
C17718 _010_ a_4165_11989# 4.31e-19
C17719 _133_ _130_ 3.75e-19
C17720 net3 state\[1\] 0.00998f
C17721 _090_ _089_ 0.205f
C17722 net53 a_6743_10933# 0.0107f
C17723 a_4512_11305# _021_ 1.91e-20
C17724 _062_ a_5536_4399# 3.44e-19
C17725 net55 _059_ 0.186f
C17726 net12 net2 0.00487f
C17727 _012_ net1 0.0346f
C17728 a_10975_4105# trim_mask\[4\] 0.0098f
C17729 a_15083_4659# a_15299_3311# 5.36e-21
C17730 _104_ a_10111_1679# 1.71e-19
C17731 _046_ _101_ 0.00309f
C17732 net40 _058_ 0.00678f
C17733 _094_ _096_ 2.17e-19
C17734 trim_mask\[0\] a_8473_5193# 3.38e-19
C17735 _019_ _041_ 8.1e-20
C17736 en_co_clk _093_ 0.00338f
C17737 net43 a_7447_8041# 1.79e-19
C17738 _050_ a_6927_3311# 0.00209f
C17739 a_10864_7387# a_10975_6031# 3.33e-21
C17740 net46 a_10699_3311# 1.93e-20
C17741 cal_itt\[1\] cal_count\[3\] 7.38e-21
C17742 en_co_clk a_5166_5193# 3.21e-19
C17743 net44 _034_ 7.88e-19
C17744 _065_ a_11016_6691# 0.164f
C17745 _107_ _088_ 0.0421f
C17746 _062_ a_9602_6941# 0.00222f
C17747 _065_ net3 0.0566f
C17748 clknet_0_clk calibrate 1.42e-19
C17749 a_7460_5807# _098_ 9.31e-21
C17750 clknet_2_2__leaf_clk a_12599_3615# 0.0763f
C17751 _050_ a_5363_4719# 2.23e-20
C17752 a_7262_5461# _107_ 0.00319f
C17753 trim_mask\[0\] a_13625_3317# 1.91e-19
C17754 clknet_2_2__leaf_clk a_11413_2767# 0.00199f
C17755 _053_ a_8307_4719# 0.00554f
C17756 _111_ a_11583_4777# 2.05e-19
C17757 a_9296_9295# _001_ 2.64e-20
C17758 _095_ net41 4.84e-20
C17759 _124_ a_11258_8790# 2.88e-19
C17760 a_13279_7119# VPWR 0.0103f
C17761 mask\[2\] a_5221_9295# 1.81e-19
C17762 _052_ a_6927_3311# 0.00804f
C17763 mask\[6\] a_3431_10933# 0.224f
C17764 mask\[3\] a_2450_9955# 2.27e-19
C17765 _107_ trim_val\[4\] 9.3e-19
C17766 a_4512_12393# a_6375_12021# 1.26e-20
C17767 a_14236_8457# _130_ 3.28e-21
C17768 a_11244_9661# a_11545_9049# 0.00227f
C17769 clknet_2_0__leaf_clk cal 0.00552f
C17770 _035_ a_12436_9129# 1.11e-21
C17771 a_6796_12381# net27 5.98e-20
C17772 net33 a_13415_2442# 7.24e-21
C17773 a_7824_11305# a_7986_10927# 0.00645f
C17774 _049_ _088_ 0.0514f
C17775 a_15023_10927# a_15023_9839# 0.00254f
C17776 a_6519_4631# _107_ 0.0112f
C17777 _049_ a_7262_5461# 4.05e-19
C17778 trim_mask\[0\] a_12310_4399# 7.89e-20
C17779 net5 clkc 0.0669f
C17780 _074_ a_1184_9117# 0.0102f
C17781 _034_ en_co_clk 5.03e-19
C17782 trim_mask\[0\] a_8583_3317# 8.59e-20
C17783 clknet_2_1__leaf_clk a_5915_10927# 0.045f
C17784 net43 a_2815_9447# 4.34e-21
C17785 _084_ net12 0.00227f
C17786 a_15023_12015# trimb[3] 9.86e-19
C17787 _098_ a_5363_4719# 1.51e-19
C17788 net21 a_4674_12015# 5.17e-20
C17789 _110_ a_11292_1251# 0.0586f
C17790 _041_ VPWR 1.69f
C17791 _010_ VPWR 0.372f
C17792 net34 net37 2.05f
C17793 a_7184_2339# VPWR 0.602f
C17794 a_13257_4943# _113_ 1.3e-20
C17795 clknet_2_0__leaf_clk a_4805_8207# 1.2e-21
C17796 clknet_2_2__leaf_clk a_8912_2589# 0.0254f
C17797 a_13470_7663# _132_ 6.93e-20
C17798 a_3116_12533# result[7] 4.15e-20
C17799 trim_mask\[3\] trim_val\[3\] 0.57f
C17800 _001_ cal_count\[3\] 3.63e-20
C17801 net19 a_9463_8725# 0.00323f
C17802 a_15023_5487# a_14972_5193# 0.00583f
C17803 a_14083_3311# a_14335_2442# 4.98e-20
C17804 net43 a_1313_10901# 0.175f
C17805 a_1313_11989# a_1095_11305# 3.17e-20
C17806 _049_ a_6519_4631# 0.0147f
C17807 a_11116_8983# a_11987_8757# 5.71e-21
C17808 a_10747_8970# a_12153_8757# 4.91e-21
C17809 _123_ a_11545_9049# 0.136f
C17810 a_8298_5487# _110_ 1.11e-20
C17811 clknet_2_3__leaf_clk a_10990_7485# 0.00101f
C17812 a_15083_4659# trim[4] 0.00125f
C17813 clknet_2_0__leaf_clk a_5547_5603# 5.13e-20
C17814 a_5699_9269# _041_ 7.76e-20
C17815 clknet_0_clk a_8298_5487# 0.327f
C17816 a_4959_1679# a_5055_1679# 0.0138f
C17817 _048_ _090_ 0.549f
C17818 a_5177_1921# a_5221_1679# 3.69e-19
C17819 _031_ a_13307_1707# 0.00952f
C17820 a_1497_8725# a_1375_9129# 3.16e-19
C17821 a_1279_9129# a_1184_9117# 0.0498f
C17822 ctln[2] VGND 0.737f
C17823 ctln[3] VGND 0.623f
C17824 ctln[4] VGND 0.632f
C17825 ctln[5] VGND 0.606f
C17826 ctln[6] VGND 0.818f
C17827 ctln[7] VGND 1.01f
C17828 ctln[1] VGND 0.617f
C17829 ctln[0] VGND 0.57f
C17830 rstn VGND 0.377f
C17831 trim[3] VGND 0.508f
C17832 trim[2] VGND 0.452f
C17833 trim[0] VGND 0.443f
C17834 en VGND 0.464f
C17835 valid VGND 0.69f
C17836 cal VGND 0.56f
C17837 trim[1] VGND 0.403f
C17838 trim[4] VGND 0.429f
C17839 sample VGND 0.392f
C17840 clkc VGND 0.269f
C17841 result[0] VGND 0.248f
C17842 clk VGND 5.72f
C17843 result[1] VGND 0.28f
C17844 comp VGND 0.325f
C17845 result[2] VGND 0.441f
C17846 trimb[4] VGND 0.441f
C17847 result[3] VGND 0.355f
C17848 trimb[1] VGND 0.418f
C17849 result[4] VGND 0.345f
C17850 trimb[0] VGND 0.459f
C17851 result[5] VGND 0.385f
C17852 trimb[2] VGND 0.496f
C17853 trimb[3] VGND 0.5f
C17854 ctlp[2] VGND 0.631f
C17855 ctlp[3] VGND 0.684f
C17856 ctlp[4] VGND 0.661f
C17857 ctlp[5] VGND 0.635f
C17858 ctlp[6] VGND 0.803f
C17859 ctlp[7] VGND 0.795f
C17860 ctlp[1] VGND 0.627f
C17861 result[7] VGND 0.506f
C17862 ctlp[0] VGND 0.707f
C17863 result[6] VGND 0.597f
C17864 VPWR VGND 0.798p
C17865 a_14931_591# VGND 0.268f
C17866 a_14471_591# VGND 0.39f
C17867 a_12631_591# VGND 0.367f
C17868 net10 VGND 0.439f
C17869 a_10752_565# VGND 0.368f
C17870 a_8767_591# VGND 0.382f
C17871 a_6927_591# VGND 0.695f
C17872 a_5363_591# VGND 0.675f
C17873 a_3063_591# VGND 0.384f
C17874 a_1276_565# VGND 0.366f
C17875 a_395_591# VGND 0.291f
C17876 a_14334_1135# VGND 2.69e-19
C17877 a_13715_1135# VGND 0.00733f
C17878 a_14526_1501# VGND 0.00405f
C17879 a_14281_1513# VGND 0.00103f
C17880 a_13869_1501# VGND 0.00579f
C17881 a_11374_1251# VGND 1.44e-19
C17882 a_10787_1135# VGND 0.00742f
C17883 a_13703_1513# VGND 0.00863f
C17884 a_13512_1501# VGND 0.08f
C17885 _057_ VGND 1.19f
C17886 a_10872_1455# VGND 0.00344f
C17887 a_9805_1473# VGND 0.00466f
C17888 _116_ VGND 0.293f
C17889 net11 VGND 0.492f
C17890 net7 VGND 0.479f
C17891 net6 VGND 0.513f
C17892 a_15023_1135# VGND 0.605f
C17893 a_14172_1513# VGND 0.305f
C17894 a_14347_1439# VGND 0.537f
C17895 a_13607_1513# VGND 0.276f
C17896 a_13825_1109# VGND 0.203f
C17897 a_13257_1141# VGND 0.34f
C17898 a_13091_1141# VGND 0.638f
C17899 a_11292_1251# VGND 0.242f
C17900 a_10569_1109# VGND 0.322f
C17901 _117_ VGND 0.302f
C17902 a_10195_1354# VGND 0.259f
C17903 a_9719_1473# VGND 0.261f
C17904 a_14184_1679# VGND 0.00343f
C17905 a_13393_1707# VGND 0.00339f
C17906 net8 VGND 0.838f
C17907 a_14099_1929# VGND 0.00736f
C17908 a_11030_1679# VGND 0.00135f
C17909 a_10785_1679# VGND 5.42e-19
C17910 _114_ VGND 0.185f
C17911 trim_val\[3\] VGND 0.737f
C17912 a_10373_1679# VGND 0.0052f
C17913 a_10207_1679# VGND 0.00754f
C17914 a_10838_2045# VGND 6.88e-20
C17915 a_5878_1679# VGND 0.00221f
C17916 a_5633_1679# VGND 9.68e-19
C17917 a_10219_2045# VGND 0.0101f
C17918 a_10016_1679# VGND 0.0801f
C17919 a_15023_1679# VGND 0.277f
C17920 a_13881_1653# VGND 0.29f
C17921 a_13307_1707# VGND 0.238f
C17922 a_10676_1679# VGND 0.27f
C17923 a_10851_1653# VGND 0.507f
C17924 a_10111_1679# VGND 0.274f
C17925 a_10329_1921# VGND 0.203f
C17926 a_9761_1679# VGND 0.333f
C17927 _032_ VGND 0.545f
C17928 a_9595_1679# VGND 0.687f
C17929 a_5221_1679# VGND 0.00579f
C17930 a_5055_1679# VGND 0.00863f
C17931 a_5067_2045# VGND 0.00472f
C17932 a_4864_1679# VGND 0.0818f
C17933 a_5524_1679# VGND 0.284f
C17934 a_5699_1653# VGND 0.525f
C17935 a_4959_1679# VGND 0.28f
C17936 a_5177_1921# VGND 0.189f
C17937 a_4609_1679# VGND 0.335f
C17938 a_4443_1679# VGND 0.715f
C17939 a_14686_2339# VGND 5.84e-19
C17940 _056_ VGND 0.351f
C17941 a_12678_2223# VGND 4.28e-20
C17942 net48 VGND 0.274f
C17943 _031_ VGND 0.364f
C17944 a_12059_2223# VGND 0.00862f
C17945 a_12870_2589# VGND 0.00257f
C17946 a_12625_2601# VGND 0.00104f
C17947 a_12213_2589# VGND 0.00639f
C17948 a_10689_2223# VGND 0.0119f
C17949 a_9734_2223# VGND 2.57e-20
C17950 a_12047_2601# VGND 0.00988f
C17951 a_11856_2589# VGND 0.0853f
C17952 a_10977_2543# VGND 0.00717f
C17953 a_10689_2543# VGND 0.00363f
C17954 a_9115_2223# VGND 0.00807f
C17955 a_9926_2589# VGND 0.00221f
C17956 a_9681_2601# VGND 0.00104f
C17957 a_7524_2223# VGND 0.00785f
C17958 a_9269_2589# VGND 0.0053f
C17959 a_9103_2601# VGND 0.00754f
C17960 a_8912_2589# VGND 0.0763f
C17961 a_7140_2223# VGND 1.07e-19
C17962 a_7942_2223# VGND 0.0836f
C17963 a_7689_2589# VGND 0.01f
C17964 a_7617_2589# VGND 0.00648f
C17965 a_3386_2223# VGND 1.01e-19
C17966 a_7181_2589# VGND 0.00122f
C17967 a_6941_2589# VGND 0.00282f
C17968 a_2767_2223# VGND 0.0114f
C17969 a_3578_2589# VGND 0.00276f
C17970 a_3333_2601# VGND 0.00109f
C17971 a_2921_2589# VGND 0.00658f
C17972 a_2755_2601# VGND 0.0123f
C17973 a_2564_2589# VGND 0.0904f
C17974 a_15023_2223# VGND 0.571f
C17975 a_14604_2339# VGND 0.242f
C17976 trim_val\[2\] VGND 0.858f
C17977 a_14335_2442# VGND 0.269f
C17978 _115_ VGND 0.329f
C17979 a_13415_2442# VGND 0.259f
C17980 a_12516_2601# VGND 0.28f
C17981 a_12691_2527# VGND 0.515f
C17982 a_11951_2601# VGND 0.273f
C17983 a_12169_2197# VGND 0.198f
C17984 a_11601_2229# VGND 0.334f
C17985 a_11435_2229# VGND 0.713f
C17986 a_10543_2455# VGND 0.399f
C17987 a_9572_2601# VGND 0.269f
C17988 a_9747_2527# VGND 0.499f
C17989 a_9007_2601# VGND 0.269f
C17990 a_9225_2197# VGND 0.195f
C17991 a_8657_2229# VGND 0.299f
C17992 _027_ VGND 0.35f
C17993 a_8491_2229# VGND 0.534f
C17994 a_7310_2223# VGND 0.187f
C17995 a_7379_2197# VGND 0.277f
C17996 a_7184_2339# VGND 0.331f
C17997 a_7223_2465# VGND 0.684f
C17998 a_6906_2355# VGND 0.294f
C17999 a_6703_2197# VGND 0.529f
C18000 a_3224_2601# VGND 0.299f
C18001 a_3399_2527# VGND 0.533f
C18002 a_2659_2601# VGND 0.299f
C18003 a_2877_2197# VGND 0.203f
C18004 a_2309_2229# VGND 0.358f
C18005 a_2143_2229# VGND 0.733f
C18006 a_14184_2767# VGND 0.00375f
C18007 a_11413_2767# VGND 0.00224f
C18008 a_11149_2767# VGND 0.00652f
C18009 a_14686_3017# VGND 3.32e-19
C18010 a_14099_3017# VGND 0.0101f
C18011 _026_ VGND 0.523f
C18012 a_11149_3017# VGND 0.00582f
C18013 a_4973_2773# VGND 0.00247f
C18014 a_4901_2773# VGND 4.78e-19
C18015 a_4709_2773# VGND 0.192f
C18016 a_15023_2767# VGND 0.553f
C18017 a_14604_3017# VGND 0.234f
C18018 a_13881_2741# VGND 0.271f
C18019 a_11067_3017# VGND 0.384f
C18020 trim_mask\[3\] VGND 1.66f
C18021 a_10655_2932# VGND 0.245f
C18022 a_10055_2767# VGND 0.569f
C18023 a_8298_2767# VGND 1.97f
C18024 a_5691_2741# VGND 0.77f
C18025 a_4815_3031# VGND 0.347f
C18026 a_3933_2767# VGND 0.755f
C18027 a_3339_2767# VGND 0.361f
C18028 a_395_2767# VGND 0.275f
C18029 a_14702_3311# VGND 1.2e-19
C18030 trim_val\[1\] VGND 0.476f
C18031 a_14083_3311# VGND 0.00798f
C18032 a_14894_3677# VGND 0.0025f
C18033 a_14649_3689# VGND 0.0014f
C18034 a_14237_3677# VGND 0.00631f
C18035 a_12586_3311# VGND 5.15e-20
C18036 a_14071_3689# VGND 0.0096f
C18037 a_13880_3677# VGND 0.0787f
C18038 a_11967_3311# VGND 0.00863f
C18039 a_12778_3677# VGND 0.00135f
C18040 a_12533_3689# VGND 4.73e-19
C18041 a_12121_3677# VGND 0.00613f
C18042 a_10781_3311# VGND 0.00581f
C18043 a_11955_3689# VGND 0.00936f
C18044 a_11764_3677# VGND 0.0839f
C18045 a_11045_3631# VGND 0.00244f
C18046 a_10781_3631# VGND 0.00755f
C18047 a_9207_3311# VGND 0.00587f
C18048 a_10018_3677# VGND 0.00127f
C18049 a_9773_3689# VGND 4.65e-19
C18050 a_9361_3677# VGND 0.00513f
C18051 a_9195_3689# VGND 0.00719f
C18052 a_9004_3677# VGND 0.0747f
C18053 a_6927_3311# VGND 0.0221f
C18054 a_4658_3427# VGND 1.36e-19
C18055 a_3110_3311# VGND 1.17e-19
C18056 a_7843_3677# VGND 0.00547f
C18057 _028_ VGND 0.391f
C18058 a_7320_3631# VGND 0.00262f
C18059 a_7200_3631# VGND 0.00368f
C18060 a_7010_3631# VGND 0.00556f
C18061 a_2491_3311# VGND 0.0147f
C18062 a_3302_3677# VGND 0.00146f
C18063 a_3057_3689# VGND 5.91e-19
C18064 a_2645_3677# VGND 0.00649f
C18065 a_2479_3689# VGND 0.00909f
C18066 a_2288_3677# VGND 0.0785f
C18067 a_15299_3311# VGND 0.223f
C18068 _055_ VGND 0.351f
C18069 a_14540_3689# VGND 0.291f
C18070 a_14715_3615# VGND 0.498f
C18071 a_13975_3689# VGND 0.279f
C18072 a_14193_3285# VGND 0.21f
C18073 a_13625_3317# VGND 0.33f
C18074 _030_ VGND 0.268f
C18075 a_13459_3317# VGND 0.553f
C18076 a_13183_3311# VGND 0.219f
C18077 a_12424_3689# VGND 0.262f
C18078 a_12599_3615# VGND 0.495f
C18079 a_11859_3689# VGND 0.283f
C18080 a_12077_3285# VGND 0.198f
C18081 a_11509_3317# VGND 0.33f
C18082 _025_ VGND 0.42f
C18083 a_11343_3317# VGND 0.622f
C18084 a_10699_3311# VGND 0.374f
C18085 trim_mask\[2\] VGND 3.02f
C18086 a_9664_3689# VGND 0.263f
C18087 a_9839_3615# VGND 0.489f
C18088 a_9099_3689# VGND 0.255f
C18089 a_9317_3285# VGND 0.177f
C18090 a_8749_3317# VGND 0.288f
C18091 _033_ VGND 0.328f
C18092 a_8583_3317# VGND 0.548f
C18093 a_7891_3617# VGND 0.248f
C18094 a_7715_3285# VGND 0.225f
C18095 a_7010_3311# VGND 0.358f
C18096 a_4576_3427# VGND 0.233f
C18097 a_2948_3689# VGND 0.267f
C18098 a_3123_3615# VGND 0.508f
C18099 a_2383_3689# VGND 0.289f
C18100 a_2601_3285# VGND 0.206f
C18101 a_2033_3317# VGND 0.343f
C18102 a_1867_3317# VGND 0.57f
C18103 a_995_3530# VGND 0.271f
C18104 a_455_3571# VGND 0.553f
C18105 a_13693_3883# VGND 0.0047f
C18106 net49 VGND 0.526f
C18107 a_11321_3855# VGND 0.00282f
C18108 a_11057_3855# VGND 0.00645f
C18109 a_9662_3855# VGND 0.0126f
C18110 a_9369_3855# VGND 0.00768f
C18111 _112_ VGND 0.343f
C18112 _113_ VGND 0.465f
C18113 a_7104_3855# VGND 0.0034f
C18114 a_6737_3855# VGND 0.17f
C18115 a_11057_4105# VGND 0.00531f
C18116 a_10270_4105# VGND 2.7e-19
C18117 trim_mask\[4\] VGND 2.77f
C18118 a_9478_4105# VGND 0.00643f
C18119 a_9369_4105# VGND 0.00636f
C18120 _119_ VGND 0.541f
C18121 a_4905_3855# VGND 0.00627f
C18122 a_4617_3855# VGND 0.00263f
C18123 a_1201_3855# VGND 0.00366f
C18124 a_937_3855# VGND 0.00604f
C18125 a_7021_4105# VGND 0.00686f
C18126 a_6822_4105# VGND 2.68e-19
C18127 a_5931_4105# VGND 0.00823f
C18128 a_5537_4105# VGND 9.13e-20
C18129 net41 VGND 3.33f
C18130 a_4617_4105# VGND 0.00357f
C18131 _015_ VGND 0.563f
C18132 _013_ VGND 0.443f
C18133 a_937_4105# VGND 0.00409f
C18134 a_14981_4020# VGND 0.252f
C18135 a_14335_4020# VGND 0.303f
C18136 a_13519_4007# VGND 0.269f
C18137 a_10975_4105# VGND 0.387f
C18138 trim_mask\[1\] VGND 1.73f
C18139 a_10188_4105# VGND 0.241f
C18140 a_9802_4007# VGND 0.174f
C18141 trim_val\[4\] VGND 0.538f
C18142 a_9003_3829# VGND 0.604f
C18143 a_7939_3855# VGND 0.375f
C18144 _054_ VGND 0.452f
C18145 a_7190_3855# VGND 0.288f
C18146 a_6519_3829# VGND 0.278f
C18147 _089_ VGND 0.343f
C18148 a_5087_3855# VGND 0.352f
C18149 state\[1\] VGND 1.15f
C18150 a_4471_4007# VGND 0.369f
C18151 state\[0\] VGND 1.03f
C18152 a_3667_3829# VGND 0.712f
C18153 a_2283_4020# VGND 0.264f
C18154 a_855_4105# VGND 0.39f
C18155 net1 VGND 0.448f
C18156 a_13915_4399# VGND 0.0106f
C18157 a_14000_4719# VGND 0.00327f
C18158 a_12310_4399# VGND 4.68e-20
C18159 a_13233_4737# VGND 0.00339f
C18160 _109_ VGND 0.232f
C18161 a_11691_4399# VGND 0.00866f
C18162 a_12502_4765# VGND 0.00221f
C18163 a_12257_4777# VGND 0.00102f
C18164 a_11845_4765# VGND 0.00596f
C18165 a_9503_4399# VGND 0.0149f
C18166 a_9166_4515# VGND 9.13e-22
C18167 a_11679_4777# VGND 0.00901f
C18168 a_11488_4765# VGND 0.0816f
C18169 _110_ VGND 2.32f
C18170 a_6822_4399# VGND 2.91e-19
C18171 a_6197_4399# VGND 2.42e-19
C18172 a_5445_4399# VGND 6.69e-20
C18173 a_5054_4399# VGND 2.21e-19
C18174 a_4970_4399# VGND 1.4e-19
C18175 a_4886_4399# VGND 4.88e-20
C18176 a_3847_4438# VGND 4.27e-19
C18177 a_3530_4438# VGND 4.4e-19
C18178 _104_ VGND 1.72f
C18179 a_8307_4719# VGND 0.295f
C18180 a_7758_4759# VGND 4.85e-19
C18181 a_7677_4759# VGND 0.00252f
C18182 net32 VGND 0.741f
C18183 a_15083_4659# VGND 0.612f
C18184 a_14655_4399# VGND 0.26f
C18185 _058_ VGND 1.68f
C18186 a_13697_4373# VGND 0.275f
C18187 a_13059_4631# VGND 0.231f
C18188 a_12148_4777# VGND 0.285f
C18189 a_12323_4703# VGND 0.629f
C18190 a_11583_4777# VGND 0.28f
C18191 a_11801_4373# VGND 0.197f
C18192 a_11233_4405# VGND 0.315f
C18193 _024_ VGND 0.361f
C18194 a_11067_4405# VGND 0.714f
C18195 a_9084_4515# VGND 0.23f
C18196 a_7800_4631# VGND 0.208f
C18197 _088_ VGND 0.271f
C18198 a_6737_4719# VGND 0.136f
C18199 _100_ VGND 0.344f
C18200 _107_ VGND 1.69f
C18201 a_5363_4719# VGND 0.167f
C18202 _093_ VGND 0.885f
C18203 a_3148_4399# VGND 0.00113f
C18204 a_1638_4399# VGND 2.91e-20
C18205 a_3751_4765# VGND 0.00301f
C18206 a_3530_4765# VGND 0.00264f
C18207 _097_ VGND 0.476f
C18208 a_3057_4719# VGND 0.161f
C18209 _014_ VGND 0.678f
C18210 a_7527_4631# VGND 0.236f
C18211 a_7019_4407# VGND 0.313f
C18212 state\[2\] VGND 1.11f
C18213 _052_ VGND 1.11f
C18214 a_6519_4631# VGND 0.27f
C18215 a_5536_4399# VGND 0.241f
C18216 a_4498_4373# VGND 0.605f
C18217 a_3817_4697# VGND 0.344f
C18218 a_3388_4631# VGND 0.263f
C18219 _099_ VGND 2.14f
C18220 a_2865_4460# VGND 0.212f
C18221 a_1019_4399# VGND 0.00515f
C18222 a_1830_4765# VGND 0.00221f
C18223 a_1585_4777# VGND 9.68e-19
C18224 a_1173_4765# VGND 0.00579f
C18225 a_1007_4777# VGND 0.00863f
C18226 a_816_4765# VGND 0.0803f
C18227 a_1476_4777# VGND 0.283f
C18228 a_1651_4703# VGND 0.527f
C18229 a_911_4777# VGND 0.26f
C18230 a_1129_4373# VGND 0.18f
C18231 a_561_4405# VGND 0.318f
C18232 _012_ VGND 0.461f
C18233 a_395_4405# VGND 0.699f
C18234 a_14526_4943# VGND 0.00219f
C18235 a_14281_4943# VGND 5.42e-19
C18236 _047_ VGND 0.443f
C18237 a_15054_5193# VGND 1.71e-19
C18238 trim_val\[0\] VGND 1.06f
C18239 a_13869_4943# VGND 0.00579f
C18240 a_13703_4943# VGND 0.00863f
C18241 a_14334_5309# VGND 2.69e-19
C18242 a_10137_4943# VGND 0.193f
C18243 a_13715_5309# VGND 0.00605f
C18244 a_13512_4943# VGND 0.0818f
C18245 a_14972_5193# VGND 0.222f
C18246 a_14172_4943# VGND 0.288f
C18247 a_14347_4917# VGND 0.508f
C18248 a_13607_4943# VGND 0.283f
C18249 a_13825_5185# VGND 0.187f
C18250 a_13257_4943# VGND 0.339f
C18251 a_13091_4943# VGND 0.678f
C18252 clknet_2_2__leaf_clk VGND 4.96f
C18253 _029_ VGND 0.548f
C18254 net50 VGND 0.543f
C18255 a_10245_5193# VGND 1.45e-19
C18256 a_9125_4943# VGND 0.0019f
C18257 a_8745_4943# VGND 0.00239f
C18258 a_8485_4943# VGND 0.00156f
C18259 _118_ VGND 0.331f
C18260 a_5731_4943# VGND 0.00334f
C18261 a_5625_4943# VGND 0.00333f
C18262 a_5537_4943# VGND 0.00162f
C18263 a_9595_5193# VGND 0.00889f
C18264 _106_ VGND 0.96f
C18265 a_8473_5193# VGND 0.00115f
C18266 a_8389_5193# VGND 8.69e-19
C18267 a_5081_4943# VGND 0.127f
C18268 a_4266_4943# VGND 0.00184f
C18269 a_4175_4943# VGND 0.00342f
C18270 a_4091_4943# VGND 0.00355f
C18271 _103_ VGND 0.596f
C18272 a_7393_5193# VGND 5.03e-19
C18273 a_6763_5193# VGND 0.0159f
C18274 a_6566_5193# VGND 0.0226f
C18275 a_6316_5193# VGND 0.0377f
C18276 _087_ VGND 0.642f
C18277 a_3365_4943# VGND 0.211f
C18278 a_3557_5193# VGND 2.75e-19
C18279 a_3461_5193# VGND 4e-19
C18280 a_12723_4943# VGND 0.27f
C18281 _111_ VGND 0.577f
C18282 _108_ VGND 3.92f
C18283 a_11023_5108# VGND 0.277f
C18284 a_8307_4943# VGND 0.539f
C18285 _105_ VGND 0.42f
C18286 a_7571_4943# VGND 0.262f
C18287 _098_ VGND 1.52f
C18288 net42 VGND 0.405f
C18289 calibrate VGND 0.991f
C18290 a_6210_4989# VGND 0.4f
C18291 a_5455_4943# VGND 0.245f
C18292 _060_ VGND 1.09f
C18293 a_4863_4917# VGND 0.234f
C18294 net54 VGND 0.961f
C18295 a_4091_5309# VGND 0.311f
C18296 a_4308_4917# VGND 0.221f
C18297 a_3891_4943# VGND 0.183f
C18298 net3 VGND 2.35f
C18299 a_3273_4943# VGND 0.236f
C18300 _090_ VGND 0.899f
C18301 a_11425_5487# VGND 5.61e-19
C18302 a_10781_5487# VGND 0.00732f
C18303 a_10055_5487# VGND 0.0101f
C18304 a_11045_5807# VGND 0.00231f
C18305 a_10781_5807# VGND 0.00653f
C18306 a_10138_5807# VGND 0.00434f
C18307 a_4725_5487# VGND 5.53e-20
C18308 a_7460_5807# VGND 0.182f
C18309 a_7210_5807# VGND 0.274f
C18310 a_5726_5807# VGND 0.00474f
C18311 _059_ VGND 0.587f
C18312 _096_ VGND 0.657f
C18313 a_1493_5487# VGND 0.0114f
C18314 a_1137_5487# VGND 4.14e-19
C18315 a_1579_5807# VGND 0.00411f
C18316 a_15023_5487# VGND 0.615f
C18317 net35 VGND 0.707f
C18318 a_10699_5487# VGND 0.378f
C18319 _066_ VGND 0.49f
C18320 trim_mask\[0\] VGND 3.21f
C18321 _064_ VGND 1.72f
C18322 a_8298_5487# VGND 2.02f
C18323 _048_ VGND 4.17f
C18324 _050_ VGND 2.06f
C18325 a_7262_5461# VGND 0.315f
C18326 a_5547_5603# VGND 0.23f
C18327 _051_ VGND 4.08f
C18328 net55 VGND 1.09f
C18329 _095_ VGND 1.08f
C18330 a_2857_5461# VGND 2.02f
C18331 _079_ VGND 0.473f
C18332 net30 VGND 3.33f
C18333 a_455_5747# VGND 0.636f
C18334 a_14649_6031# VGND 0.00703f
C18335 a_14181_6031# VGND 0.00565f
C18336 a_13825_6031# VGND 0.223f
C18337 a_13349_6031# VGND 0.223f
C18338 a_13193_6031# VGND 0.0057f
C18339 a_12410_6031# VGND 0.00143f
C18340 a_12165_6031# VGND 5.76e-19
C18341 _136_ VGND 1.24f
C18342 a_13441_6281# VGND 4.18e-19
C18343 a_11753_6031# VGND 0.00631f
C18344 a_11587_6031# VGND 0.00976f
C18345 a_12218_6397# VGND 8.12e-20
C18346 a_9529_6059# VGND 0.00355f
C18347 a_11599_6397# VGND 0.00878f
C18348 a_11396_6031# VGND 0.0749f
C18349 a_15023_6031# VGND 0.286f
C18350 _061_ VGND 0.376f
C18351 a_14564_6397# VGND 0.372f
C18352 a_14379_6397# VGND 0.29f
C18353 _135_ VGND 0.282f
C18354 a_13783_6183# VGND 0.253f
C18355 a_13111_6031# VGND 0.259f
C18356 cal_count\[3\] VGND 0.86f
C18357 a_12056_6031# VGND 0.266f
C18358 a_12231_6005# VGND 0.51f
C18359 a_11491_6031# VGND 0.285f
C18360 net46 VGND 7.59f
C18361 a_11709_6273# VGND 0.195f
C18362 a_11141_6031# VGND 0.333f
C18363 _038_ VGND 0.556f
C18364 a_10975_6031# VGND 0.674f
C18365 _092_ VGND 4.12f
C18366 a_9043_6031# VGND 0.00528f
C18367 a_8949_6031# VGND 0.00583f
C18368 a_5694_6031# VGND 0.00248f
C18369 a_5449_6031# VGND 0.00108f
C18370 a_8949_6281# VGND 0.00718f
C18371 a_6197_6281# VGND 3.87e-19
C18372 en_co_clk VGND 1.64f
C18373 a_5037_6031# VGND 0.00525f
C18374 a_4871_6031# VGND 0.0074f
C18375 a_5502_6397# VGND 5.36e-20
C18376 a_1830_6031# VGND 0.00248f
C18377 a_1585_6031# VGND 0.00103f
C18378 a_4883_6397# VGND 0.00719f
C18379 a_4680_6031# VGND 0.0771f
C18380 a_10005_6031# VGND 0.767f
C18381 _091_ VGND 0.362f
C18382 a_9443_6059# VGND 0.227f
C18383 a_8820_6005# VGND 0.322f
C18384 _075_ VGND 0.892f
C18385 a_5340_6031# VGND 0.293f
C18386 a_5515_6005# VGND 0.528f
C18387 a_4775_6031# VGND 0.269f
C18388 a_4993_6273# VGND 0.202f
C18389 a_4425_6031# VGND 0.336f
C18390 a_4259_6031# VGND 0.54f
C18391 a_3830_6281# VGND 2.64e-19
C18392 _120_ VGND 0.397f
C18393 _094_ VGND 1.31f
C18394 a_3529_6281# VGND 9.65e-19
C18395 a_2476_6281# VGND 3.36e-19
C18396 a_1173_6031# VGND 0.00613f
C18397 a_1007_6031# VGND 0.00927f
C18398 a_1638_6397# VGND 3.88e-20
C18399 a_1019_6397# VGND 0.00839f
C18400 a_816_6031# VGND 0.0836f
C18401 a_3748_6281# VGND 0.223f
C18402 _049_ VGND 3.35f
C18403 a_2313_6183# VGND 0.245f
C18404 a_1476_6031# VGND 0.283f
C18405 a_1651_6005# VGND 0.51f
C18406 a_911_6031# VGND 0.28f
C18407 a_1129_6273# VGND 0.203f
C18408 a_561_6031# VGND 0.331f
C18409 _004_ VGND 0.791f
C18410 a_395_6031# VGND 0.71f
C18411 a_11098_6691# VGND 2.82e-19
C18412 a_9919_6614# VGND 2.7e-19
C18413 a_9602_6614# VGND 5.37e-20
C18414 a_9823_6941# VGND 0.00331f
C18415 a_9602_6941# VGND 0.00263f
C18416 a_8935_6895# VGND 0.183f
C18417 a_8745_6895# VGND 0.193f
C18418 a_8495_6895# VGND 0.176f
C18419 a_7897_6913# VGND 0.00502f
C18420 _034_ VGND 0.383f
C18421 a_15299_6575# VGND 0.284f
C18422 net5 VGND 0.393f
C18423 a_11016_6691# VGND 0.244f
C18424 a_9889_6873# VGND 0.3f
C18425 _062_ VGND 1.91f
C18426 a_9460_6807# VGND 0.247f
C18427 a_8307_6575# VGND 0.34f
C18428 a_7723_6807# VGND 0.252f
C18429 _073_ VGND 0.777f
C18430 a_6515_6794# VGND 0.315f
C18431 a_4167_6575# VGND 0.255f
C18432 _121_ VGND 0.329f
C18433 _039_ VGND 0.325f
C18434 a_1549_6794# VGND 0.257f
C18435 net22 VGND 1.22f
C18436 a_448_6549# VGND 0.354f
C18437 a_15289_7119# VGND 0.00178f
C18438 a_14282_7119# VGND 0.00446f
C18439 a_13821_7119# VGND 0.0019f
C18440 a_13279_7119# VGND 0.322f
C18441 a_14870_7369# VGND 2.53e-19
C18442 a_14199_7369# VGND 0.0125f
C18443 _134_ VGND 0.531f
C18444 a_13557_7369# VGND 3.11e-20
C18445 a_13356_7369# VGND 1.01e-19
C18446 a_11369_7119# VGND 0.0094f
C18447 a_11297_7119# VGND 0.00622f
C18448 a_10861_7119# VGND 0.00116f
C18449 a_10621_7119# VGND 0.00405f
C18450 a_14788_7369# VGND 0.222f
C18451 _131_ VGND 1.47f
C18452 a_14422_7093# VGND 0.233f
C18453 _130_ VGND 0.376f
C18454 a_14063_7093# VGND 0.393f
C18455 a_13142_7271# VGND 0.193f
C18456 a_11622_7485# VGND 0.0817f
C18457 a_11204_7485# VGND 0.00897f
C18458 a_7442_7119# VGND 0.00255f
C18459 a_7197_7119# VGND 0.00115f
C18460 a_10820_7485# VGND 1e-19
C18461 cal_itt\[3\] VGND 0.684f
C18462 a_6785_7119# VGND 0.00723f
C18463 a_6619_7119# VGND 0.0132f
C18464 a_7250_7485# VGND 9.17e-20
C18465 a_4222_7119# VGND 0.00139f
C18466 a_3977_7119# VGND 5.49e-19
C18467 a_6631_7485# VGND 0.0132f
C18468 a_6428_7119# VGND 0.0838f
C18469 a_10990_7485# VGND 0.203f
C18470 a_11059_7356# VGND 0.276f
C18471 a_10903_7261# VGND 0.644f
C18472 a_10864_7387# VGND 0.321f
C18473 a_10586_7371# VGND 0.3f
C18474 a_10383_7093# VGND 0.548f
C18475 a_8022_7119# VGND 2.03f
C18476 a_7088_7119# VGND 0.279f
C18477 a_7263_7093# VGND 0.497f
C18478 a_6523_7119# VGND 0.292f
C18479 a_6741_7361# VGND 0.203f
C18480 a_6173_7119# VGND 0.34f
C18481 _003_ VGND 0.583f
C18482 a_6007_7119# VGND 0.693f
C18483 a_5363_7369# VGND 0.0091f
C18484 a_4995_7119# VGND 0.363f
C18485 a_3565_7119# VGND 0.00527f
C18486 a_3399_7119# VGND 0.0075f
C18487 a_4030_7485# VGND 6.7e-20
C18488 a_1830_7119# VGND 0.00236f
C18489 a_1585_7119# VGND 4.86e-19
C18490 a_3411_7485# VGND 0.00642f
C18491 a_3208_7119# VGND 0.0761f
C18492 a_3868_7119# VGND 0.264f
C18493 a_4043_7093# VGND 0.494f
C18494 a_3303_7119# VGND 0.254f
C18495 a_3521_7361# VGND 0.177f
C18496 a_2953_7119# VGND 0.29f
C18497 a_2787_7119# VGND 0.569f
C18498 a_1173_7119# VGND 0.00596f
C18499 a_1007_7119# VGND 0.00895f
C18500 a_1638_7485# VGND 3.11e-20
C18501 a_1019_7485# VGND 0.00526f
C18502 a_816_7119# VGND 0.0809f
C18503 a_1476_7119# VGND 0.261f
C18504 a_1651_7093# VGND 0.505f
C18505 a_911_7119# VGND 0.263f
C18506 a_1129_7361# VGND 0.183f
C18507 a_561_7119# VGND 0.304f
C18508 a_395_7119# VGND 0.687f
C18509 a_14485_7663# VGND 0.00413f
C18510 a_12824_7663# VGND 3.4e-19
C18511 a_14733_7983# VGND 0.00585f
C18512 a_14377_7983# VGND 0.247f
C18513 _133_ VGND 0.303f
C18514 cal_count\[2\] VGND 0.788f
C18515 a_13164_8029# VGND 0.00523f
C18516 a_13092_8029# VGND 0.00169f
C18517 a_12924_8029# VGND 0.00386f
C18518 a_12664_8029# VGND 0.00583f
C18519 a_12454_8041# VGND 0.00172f
C18520 a_12249_7663# VGND 0.101f
C18521 a_9957_7663# VGND 0.0116f
C18522 a_10877_7983# VGND 0.00209f
C18523 a_10043_7983# VGND 0.00387f
C18524 a_8078_7663# VGND 3.27e-20
C18525 a_9693_8029# VGND 8.26e-19
C18526 a_9621_8029# VGND 0.00221f
C18527 a_8761_7983# VGND 0.002f
C18528 a_7459_7663# VGND 0.00576f
C18529 a_8270_8029# VGND 0.00232f
C18530 a_8025_8041# VGND 4.71e-19
C18531 a_7613_8029# VGND 0.00514f
C18532 a_2225_7663# VGND 0.00637f
C18533 a_1125_7663# VGND 0.00463f
C18534 a_7447_8041# VGND 0.00725f
C18535 a_7256_8029# VGND 0.0756f
C18536 _016_ VGND 0.349f
C18537 a_2489_7983# VGND 0.00382f
C18538 a_2225_7983# VGND 0.00649f
C18539 a_1211_7983# VGND 0.00379f
C18540 _005_ VGND 0.388f
C18541 a_15259_7637# VGND 0.356f
C18542 _132_ VGND 0.444f
C18543 a_14335_7895# VGND 0.325f
C18544 a_13470_7663# VGND 0.205f
C18545 a_12900_7663# VGND 0.42f
C18546 a_13050_7637# VGND 0.176f
C18547 a_12344_8041# VGND 0.453f
C18548 a_12520_7637# VGND 0.197f
C18549 a_12061_7669# VGND 0.518f
C18550 _037_ VGND 0.386f
C18551 a_11895_7669# VGND 0.539f
C18552 _053_ VGND 3.56f
C18553 _063_ VGND 1.71f
C18554 cal_itt\[1\] VGND 1.27f
C18555 a_9459_7895# VGND 0.247f
C18556 _067_ VGND 2.03f
C18557 _071_ VGND 0.312f
C18558 a_7916_8041# VGND 0.268f
C18559 a_8091_7967# VGND 0.491f
C18560 a_7351_8041# VGND 0.267f
C18561 a_7569_7637# VGND 0.177f
C18562 a_7001_7669# VGND 0.301f
C18563 a_6835_7669# VGND 0.6f
C18564 a_5691_7637# VGND 0.737f
C18565 a_4677_7882# VGND 0.262f
C18566 clknet_0_clk VGND 5.41f
C18567 a_2857_7637# VGND 1.97f
C18568 a_2143_7663# VGND 0.393f
C18569 mask\[0\] VGND 3.75f
C18570 net45 VGND 6.51f
C18571 a_1467_7923# VGND 0.529f
C18572 _080_ VGND 0.21f
C18573 a_448_7637# VGND 0.346f
C18574 a_14981_8235# VGND 0.00495f
C18575 a_13279_8207# VGND 0.305f
C18576 a_8301_8207# VGND 0.185f
C18577 a_6419_8207# VGND 0.00381f
C18578 a_6198_8207# VGND 0.00336f
C18579 a_14318_8457# VGND 2.64e-19
C18580 a_13557_8457# VGND 3.14e-20
C18581 a_13356_8457# VGND 1.8e-19
C18582 a_9761_8457# VGND 1.59e-20
C18583 a_9677_8457# VGND 2.46e-19
C18584 _001_ VGND 0.769f
C18585 a_8386_8457# VGND 2.39e-19
C18586 _002_ VGND 0.933f
C18587 a_5050_8207# VGND 0.00221f
C18588 a_4805_8207# VGND 4.65e-19
C18589 a_6515_8534# VGND 0.00133f
C18590 a_6198_8534# VGND 5.68e-19
C18591 net51 VGND 0.914f
C18592 a_6485_8181# VGND 0.308f
C18593 net2 VGND 6.73f
C18594 a_4393_8207# VGND 0.00507f
C18595 a_4227_8207# VGND 0.00711f
C18596 a_4858_8573# VGND 5.39e-20
C18597 a_3317_8207# VGND 0.00257f
C18598 a_3053_8207# VGND 0.00679f
C18599 a_4239_8573# VGND 0.00834f
C18600 a_4036_8207# VGND 0.0797f
C18601 a_14807_8359# VGND 0.277f
C18602 a_14236_8457# VGND 0.246f
C18603 a_13142_8359# VGND 0.18f
C18604 _069_ VGND 0.224f
C18605 cal_itt\[2\] VGND 0.881f
C18606 _070_ VGND 0.54f
C18607 _072_ VGND 0.607f
C18608 a_8083_8181# VGND 0.26f
C18609 a_6885_8372# VGND 0.256f
C18610 a_6056_8359# VGND 0.281f
C18611 _077_ VGND 0.189f
C18612 a_5535_8181# VGND 0.482f
C18613 a_4696_8207# VGND 0.275f
C18614 a_4871_8181# VGND 0.507f
C18615 a_4131_8207# VGND 0.279f
C18616 a_4349_8449# VGND 0.196f
C18617 a_3781_8207# VGND 0.319f
C18618 a_3615_8207# VGND 0.53f
C18619 clknet_2_0__leaf_clk VGND 5.23f
C18620 _017_ VGND 0.267f
C18621 a_3053_8457# VGND 0.0103f
C18622 _040_ VGND 1.4f
C18623 a_2174_8457# VGND 9.13e-22
C18624 net23 VGND 1.7f
C18625 a_1229_8457# VGND 0.00114f
C18626 a_2971_8457# VGND 0.378f
C18627 mask\[1\] VGND 1.52f
C18628 a_2092_8457# VGND 0.229f
C18629 a_455_8181# VGND 0.617f
C18630 a_14467_8751# VGND 0.0243f
C18631 a_13100_8751# VGND 6.77e-20
C18632 a_12916_8751# VGND 5.26e-19
C18633 a_12522_8751# VGND 1.7e-19
C18634 a_14552_9071# VGND 0.00472f
C18635 _129_ VGND 0.727f
C18636 cal_count\[1\] VGND 0.637f
C18637 a_11575_8790# VGND 4.71e-19
C18638 a_11258_8790# VGND 6.4e-19
C18639 a_13256_9117# VGND 0.00474f
C18640 a_13184_9117# VGND 0.00119f
C18641 a_13016_9117# VGND 0.00337f
C18642 a_12756_9117# VGND 0.00535f
C18643 a_12546_9129# VGND 8.52e-19
C18644 a_12341_8751# VGND 0.0985f
C18645 a_11479_9117# VGND 0.00328f
C18646 a_11258_9117# VGND 0.00302f
C18647 a_3922_8867# VGND 2.45e-19
C18648 a_2689_8751# VGND 0.0166f
C18649 a_2775_9071# VGND 0.00523f
C18650 _081_ VGND 0.625f
C18651 a_1387_8751# VGND 0.008f
C18652 a_2198_9117# VGND 0.00145f
C18653 a_1953_9129# VGND 4.65e-19
C18654 a_1541_9117# VGND 0.00628f
C18655 a_1375_9129# VGND 0.00941f
C18656 a_1184_9117# VGND 0.083f
C18657 a_15023_8751# VGND 0.653f
C18658 net40 VGND 2.02f
C18659 a_14249_8725# VGND 0.305f
C18660 a_13919_8751# VGND 0.222f
C18661 _041_ VGND 4.88f
C18662 a_13562_8751# VGND 0.184f
C18663 a_12992_8751# VGND 0.41f
C18664 a_13142_8725# VGND 0.168f
C18665 a_12436_9129# VGND 0.451f
C18666 a_12612_8725# VGND 0.196f
C18667 a_12153_8757# VGND 0.37f
C18668 _036_ VGND 0.269f
C18669 a_11987_8757# VGND 0.521f
C18670 a_11545_9049# VGND 0.3f
C18671 _122_ VGND 2.02f
C18672 _123_ VGND 1.17f
C18673 a_11116_8983# VGND 0.279f
C18674 _124_ VGND 0.254f
C18675 a_10747_8970# VGND 0.249f
C18676 net4 VGND 3.56f
C18677 a_9463_8725# VGND 0.411f
C18678 _068_ VGND 0.547f
C18679 _076_ VGND 1.08f
C18680 a_6793_8970# VGND 0.275f
C18681 _065_ VGND 3.18f
C18682 a_5423_9011# VGND 0.642f
C18683 a_3840_8867# VGND 0.244f
C18684 net24 VGND 0.959f
C18685 a_1844_9129# VGND 0.261f
C18686 a_2019_9055# VGND 0.477f
C18687 a_1279_9129# VGND 0.288f
C18688 a_1497_8725# VGND 0.202f
C18689 a_929_8757# VGND 0.317f
C18690 _006_ VGND 0.439f
C18691 a_763_8757# VGND 0.729f
C18692 a_15111_9295# VGND 0.00528f
C18693 a_14565_9295# VGND 0.00886f
C18694 a_11508_9295# VGND 0.00475f
C18695 a_11436_9295# VGND 0.00121f
C18696 a_11268_9295# VGND 0.00341f
C18697 a_11008_9295# VGND 0.00541f
C18698 a_10798_9295# VGND 8.36e-19
C18699 a_14733_9545# VGND 0.00143f
C18700 a_14377_9545# VGND 0.0334f
C18701 _128_ VGND 0.71f
C18702 a_9650_9295# VGND 0.00242f
C18703 a_9405_9295# VGND 0.00107f
C18704 a_11352_9661# VGND 3.5e-19
C18705 a_11168_9661# VGND 9.02e-19
C18706 a_10774_9661# VGND 5.72e-19
C18707 a_10593_9295# VGND 0.112f
C18708 _125_ VGND 1.1f
C18709 a_15159_9269# VGND 0.235f
C18710 _126_ VGND 0.724f
C18711 a_14983_9269# VGND 0.222f
C18712 cal_count\[0\] VGND 1.39f
C18713 _127_ VGND 0.349f
C18714 a_14347_9480# VGND 0.366f
C18715 a_11814_9295# VGND 0.22f
C18716 a_11244_9661# VGND 0.465f
C18717 a_11394_9509# VGND 0.193f
C18718 a_10688_9295# VGND 0.469f
C18719 a_10864_9269# VGND 0.201f
C18720 a_10405_9295# VGND 0.402f
C18721 _035_ VGND 0.496f
C18722 a_10239_9295# VGND 0.568f
C18723 cal_itt\[0\] VGND 1.61f
C18724 a_8993_9295# VGND 0.00604f
C18725 a_8827_9295# VGND 0.00915f
C18726 a_9458_9661# VGND 5.06e-20
C18727 a_5878_9295# VGND 0.00221f
C18728 a_5633_9295# VGND 5.27e-19
C18729 a_8839_9661# VGND 0.00584f
C18730 a_8636_9295# VGND 0.0836f
C18731 a_9296_9295# VGND 0.288f
C18732 a_9471_9269# VGND 0.615f
C18733 a_8731_9295# VGND 0.262f
C18734 a_8949_9537# VGND 0.193f
C18735 a_8381_9295# VGND 0.328f
C18736 _000_ VGND 0.753f
C18737 a_8215_9295# VGND 0.709f
C18738 clknet_2_3__leaf_clk VGND 3.83f
C18739 a_5221_9295# VGND 0.00604f
C18740 a_5055_9295# VGND 0.00915f
C18741 a_5686_9661# VGND 5.06e-20
C18742 a_3249_9295# VGND 0.00675f
C18743 a_2961_9295# VGND 0.00218f
C18744 a_1763_9295# VGND 0.00429f
C18745 a_5067_9661# VGND 0.00562f
C18746 a_4864_9295# VGND 0.0814f
C18747 a_5524_9295# VGND 0.268f
C18748 a_5699_9269# VGND 0.498f
C18749 a_4959_9295# VGND 0.284f
C18750 a_5177_9537# VGND 0.186f
C18751 a_4609_9295# VGND 0.312f
C18752 a_4443_9295# VGND 0.695f
C18753 a_2961_9545# VGND 0.00485f
C18754 a_1677_9545# VGND 0.00848f
C18755 a_1045_9545# VGND 3.87e-19
C18756 a_2815_9447# VGND 0.388f
C18757 _082_ VGND 0.319f
C18758 a_448_9269# VGND 0.333f
C18759 a_9074_9955# VGND 1.18e-19
C18760 a_7710_9839# VGND 8.96e-20
C18761 a_7091_9839# VGND 0.00796f
C18762 a_7902_10205# VGND 0.00141f
C18763 a_7657_10217# VGND 5.6e-19
C18764 a_7245_10205# VGND 0.0053f
C18765 a_6007_9839# VGND 0.0058f
C18766 a_5829_9839# VGND 1.66e-20
C18767 a_4801_9839# VGND 0.00455f
C18768 a_4030_9839# VGND 8.16e-20
C18769 a_7079_10217# VGND 0.00756f
C18770 a_6888_10205# VGND 0.0779f
C18771 a_6090_10159# VGND 0.00382f
C18772 a_5089_10159# VGND 0.00646f
C18773 a_4801_10159# VGND 0.00263f
C18774 _019_ VGND 0.277f
C18775 mask\[2\] VGND 2.7f
C18776 a_3411_9839# VGND 0.00904f
C18777 a_4222_10205# VGND 0.00247f
C18778 a_3977_10217# VGND 5.51e-19
C18779 a_3565_10205# VGND 0.00527f
C18780 a_2450_9955# VGND 1.78e-19
C18781 a_1638_9839# VGND 4.62e-20
C18782 a_3399_10217# VGND 0.00744f
C18783 a_3208_10205# VGND 0.0755f
C18784 a_1019_9839# VGND 0.00625f
C18785 a_1830_10205# VGND 0.00134f
C18786 a_1585_10217# VGND 4.86e-19
C18787 a_1173_10205# VGND 0.00597f
C18788 a_1007_10217# VGND 0.00897f
C18789 a_816_10205# VGND 0.0809f
C18790 a_15023_9839# VGND 0.595f
C18791 net37 VGND 1.61f
C18792 a_8992_9955# VGND 0.231f
C18793 a_7548_10217# VGND 0.267f
C18794 a_7723_10143# VGND 0.501f
C18795 a_6983_10217# VGND 0.275f
C18796 a_7201_9813# VGND 0.194f
C18797 a_6633_9845# VGND 0.327f
C18798 _008_ VGND 0.387f
C18799 a_6467_9845# VGND 0.586f
C18800 _083_ VGND 0.424f
C18801 a_4655_10071# VGND 0.365f
C18802 a_3868_10217# VGND 0.279f
C18803 a_4043_10143# VGND 0.487f
C18804 a_3303_10217# VGND 0.274f
C18805 a_3521_9813# VGND 0.193f
C18806 a_2953_9845# VGND 0.313f
C18807 _018_ VGND 0.501f
C18808 a_2787_9845# VGND 0.525f
C18809 a_2368_9955# VGND 0.234f
C18810 mask\[3\] VGND 1.48f
C18811 net25 VGND 1.13f
C18812 a_1476_10217# VGND 0.26f
C18813 a_1651_10143# VGND 0.484f
C18814 a_911_10217# VGND 0.285f
C18815 a_1129_9813# VGND 0.183f
C18816 a_561_9845# VGND 0.302f
C18817 _007_ VGND 0.442f
C18818 a_395_9845# VGND 0.699f
C18819 net9 VGND 1.43f
C18820 a_9374_10383# VGND 0.00133f
C18821 a_9129_10383# VGND 0.00103f
C18822 a_8717_10383# VGND 0.00595f
C18823 a_8551_10383# VGND 0.00896f
C18824 a_9182_10749# VGND 2.27e-20
C18825 a_6445_10383# VGND 0.00485f
C18826 a_6181_10383# VGND 0.0068f
C18827 a_1764_10383# VGND 0.0037f
C18828 a_8563_10749# VGND 0.00734f
C18829 a_8360_10383# VGND 0.0814f
C18830 net31 VGND 2.51f
C18831 a_11803_10383# VGND 0.287f
C18832 _042_ VGND 3.6f
C18833 a_9871_10383# VGND 0.249f
C18834 _043_ VGND 0.988f
C18835 a_9020_10383# VGND 0.288f
C18836 a_9195_10357# VGND 0.492f
C18837 a_8455_10383# VGND 0.285f
C18838 net47 VGND 5.48f
C18839 a_8673_10625# VGND 0.197f
C18840 a_8105_10383# VGND 0.322f
C18841 a_7939_10383# VGND 0.658f
C18842 _020_ VGND 1.08f
C18843 a_6181_10633# VGND 0.0048f
C18844 a_1679_10633# VGND 0.00703f
C18845 a_6099_10633# VGND 0.42f
C18846 mask\[4\] VGND 3.02f
C18847 a_1461_10357# VGND 0.286f
C18848 net26 VGND 3.39f
C18849 a_448_10357# VGND 0.353f
C18850 a_7986_10927# VGND 3.52e-20
C18851 a_7367_10927# VGND 0.0084f
C18852 a_8178_11293# VGND 0.00233f
C18853 a_7933_11305# VGND 0.00103f
C18854 a_7521_11293# VGND 0.00602f
C18855 a_5997_10927# VGND 0.00428f
C18856 a_7355_11305# VGND 0.00915f
C18857 a_7164_11293# VGND 0.084f
C18858 a_6261_11247# VGND 0.00372f
C18859 a_5997_11247# VGND 0.00623f
C18860 a_4055_10927# VGND 0.00788f
C18861 a_4866_11293# VGND 0.00127f
C18862 a_4621_11305# VGND 4.65e-19
C18863 a_4209_11293# VGND 0.00509f
C18864 a_2869_10927# VGND 0.00886f
C18865 a_4043_11305# VGND 0.00713f
C18866 a_3852_11293# VGND 0.075f
C18867 a_3133_11247# VGND 0.00239f
C18868 a_2869_11247# VGND 0.00847f
C18869 _102_ VGND 0.548f
C18870 a_1203_10927# VGND 0.00471f
C18871 a_2014_11293# VGND 0.00221f
C18872 a_1769_11305# VGND 9.68e-19
C18873 a_1357_11293# VGND 0.00579f
C18874 a_1191_11305# VGND 0.00863f
C18875 a_1000_11293# VGND 0.0818f
C18876 a_15023_10927# VGND 0.62f
C18877 net36 VGND 0.36f
C18878 net33 VGND 1.29f
C18879 a_7824_11305# VGND 0.277f
C18880 a_7999_11231# VGND 0.516f
C18881 a_7259_11305# VGND 0.28f
C18882 a_7477_10901# VGND 0.196f
C18883 a_6909_10933# VGND 0.327f
C18884 _021_ VGND 0.541f
C18885 a_6743_10933# VGND 0.653f
C18886 a_5915_10927# VGND 0.376f
C18887 net53 VGND 1.83f
C18888 a_4512_11305# VGND 0.265f
C18889 a_4687_11231# VGND 0.513f
C18890 a_3947_11305# VGND 0.282f
C18891 a_4165_10901# VGND 0.195f
C18892 a_3597_10933# VGND 0.322f
C18893 _022_ VGND 0.261f
C18894 a_3431_10933# VGND 0.539f
C18895 a_2787_10927# VGND 0.383f
C18896 _101_ VGND 2.46f
C18897 net52 VGND 2.89f
C18898 a_1660_11305# VGND 0.28f
C18899 a_1835_11231# VGND 0.507f
C18900 a_1095_11305# VGND 0.264f
C18901 a_1313_10901# VGND 0.186f
C18902 a_745_10933# VGND 0.315f
C18903 _023_ VGND 0.344f
C18904 a_579_10933# VGND 0.657f
C18905 a_5998_11471# VGND 0.00418f
C18906 a_3511_11471# VGND 0.00399f
C18907 a_1579_11471# VGND 0.00384f
C18908 a_8154_11721# VGND 2.29e-19
C18909 net12 VGND 2.33f
C18910 a_5915_11721# VGND 0.00526f
C18911 net13 VGND 1.36f
C18912 a_3425_11721# VGND 0.0103f
C18913 a_1493_11721# VGND 0.00787f
C18914 a_1137_11721# VGND 4.16e-19
C18915 a_8767_11471# VGND 0.285f
C18916 _044_ VGND 0.489f
C18917 a_8072_11721# VGND 0.253f
C18918 mask\[5\] VGND 1.26f
C18919 a_4167_11471# VGND 0.253f
C18920 _078_ VGND 3.19f
C18921 _086_ VGND 0.232f
C18922 a_448_11445# VGND 0.363f
C18923 a_7618_12015# VGND 1.66e-19
C18924 net27 VGND 4.33f
C18925 a_6999_12015# VGND 0.0118f
C18926 a_7810_12381# VGND 0.00257f
C18927 a_7565_12393# VGND 0.00115f
C18928 a_7153_12381# VGND 0.00634f
C18929 a_6197_12015# VGND 4.76e-19
C18930 a_5578_12131# VGND 1.76e-19
C18931 a_4674_12015# VGND 1.18e-19
C18932 a_6987_12393# VGND 0.00977f
C18933 a_6796_12381# VGND 0.0868f
C18934 a_4055_12015# VGND 0.00836f
C18935 a_4866_12381# VGND 0.00137f
C18936 a_4621_12393# VGND 5.28e-19
C18937 a_4209_12381# VGND 0.00526f
C18938 a_2910_12131# VGND 5.09e-19
C18939 a_1822_12015# VGND 1.18e-19
C18940 a_4043_12393# VGND 0.00748f
C18941 a_3852_12381# VGND 0.0799f
C18942 _046_ VGND 0.346f
C18943 a_1203_12015# VGND 0.00755f
C18944 a_2014_12381# VGND 0.00221f
C18945 a_1769_12393# VGND 0.00107f
C18946 a_1357_12381# VGND 0.00605f
C18947 a_1191_12393# VGND 0.00911f
C18948 a_1000_12381# VGND 0.0837f
C18949 a_15023_12015# VGND 0.635f
C18950 net38 VGND 0.701f
C18951 net34 VGND 1.93f
C18952 a_7456_12393# VGND 0.294f
C18953 a_7631_12319# VGND 0.515f
C18954 a_6891_12393# VGND 0.293f
C18955 net44 VGND 5.07f
C18956 a_7109_11989# VGND 0.211f
C18957 a_6541_12021# VGND 0.37f
C18958 _009_ VGND 0.582f
C18959 a_6375_12021# VGND 0.715f
C18960 _084_ VGND 0.262f
C18961 a_5496_12131# VGND 0.228f
C18962 mask\[6\] VGND 2.95f
C18963 a_4512_12393# VGND 0.265f
C18964 a_4687_12319# VGND 0.505f
C18965 a_3947_12393# VGND 0.262f
C18966 a_4165_11989# VGND 0.181f
C18967 a_3597_12021# VGND 0.334f
C18968 a_3431_12021# VGND 0.543f
C18969 a_2828_12131# VGND 0.258f
C18970 mask\[7\] VGND 2.23f
C18971 a_1660_12393# VGND 0.288f
C18972 a_1835_12319# VGND 0.543f
C18973 a_1095_12393# VGND 0.277f
C18974 net43 VGND 11.2f
C18975 a_1313_11989# VGND 0.191f
C18976 a_745_12021# VGND 0.323f
C18977 _011_ VGND 0.41f
C18978 a_579_12021# VGND 0.66f
C18979 clknet_2_1__leaf_clk VGND 5.95f
C18980 a_15023_12559# VGND 0.611f
C18981 net39 VGND 0.73f
C18982 a_14471_12559# VGND 0.406f
C18983 net16 VGND 2.48f
C18984 a_12631_12559# VGND 0.359f
C18985 net17 VGND 1.36f
C18986 net18 VGND 2.76f
C18987 a_10752_12533# VGND 0.381f
C18988 net19 VGND 2.07f
C18989 a_3513_12809# VGND 9.28e-19
C18990 _010_ VGND 0.55f
C18991 a_8820_12533# VGND 0.372f
C18992 a_6927_12559# VGND 0.637f
C18993 net20 VGND 1.21f
C18994 a_6191_12559# VGND 0.292f
C18995 _045_ VGND 0.614f
C18996 a_5363_12559# VGND 0.641f
C18997 net21 VGND 0.868f
C18998 _074_ VGND 4.98f
C18999 _085_ VGND 0.39f
C19000 net15 VGND 1.58f
C19001 a_3116_12533# VGND 0.372f
C19002 net29 VGND 1.51f
C19003 a_1644_12533# VGND 0.365f
C19004 net14 VGND 1.56f
C19005 a_1099_12533# VGND 0.629f
C19006 net28 VGND 2.38f
C19007 a_455_12533# VGND 0.599f
C19008 net3.t2 VGND 0.0332f
C19009 net3.t4 VGND 0.0225f
C19010 net3.n0 VGND 0.0941f
C19011 net3.t3 VGND 0.0318f
C19012 net3.t5 VGND 0.0253f
C19013 net3.n1 VGND 0.0758f
C19014 net3.n2 VGND 0.0852f
C19015 net3.n3 VGND 0.922f
C19016 net3.t1 VGND 0.0409f
C19017 net3.n4 VGND 0.0617f
C19018 net3.n5 VGND 0.0267f
C19019 net3.t0 VGND 0.0388f
C19020 net3.n6 VGND 0.176f
C19021 net4.n0 VGND 1.08f
C19022 net4.n1 VGND 0.423f
C19023 net4.t5 VGND 0.0302f
C19024 net4.t2 VGND 0.0165f
C19025 net4.n2 VGND 0.0466f
C19026 net4.n3 VGND 0.00408f
C19027 net4.t6 VGND 0.0151f
C19028 net4.n4 VGND 0.0108f
C19029 net4.n5 VGND 0.0244f
C19030 net4.n6 VGND 0.00363f
C19031 net4.t3 VGND 0.0297f
C19032 net4.n7 VGND 0.0281f
C19033 net4.n8 VGND 0.0042f
C19034 net4.t1 VGND 0.0293f
C19035 net4.n9 VGND 0.0453f
C19036 net4.n10 VGND 0.0192f
C19037 net4.t0 VGND 0.0278f
C19038 net4.n11 VGND 0.531f
C19039 net4.t4 VGND 0.0163f
C19040 net4.t7 VGND 0.0252f
C19041 net4.n12 VGND 0.0598f
C19042 net4.n13 VGND 0.0193f
C19043 net4.n14 VGND 0.00419f
C19044 net4.n15 VGND 0.00419f
C19045 net4.n16 VGND 0.808f
C19046 net4.n17 VGND 0.0427f
C19047 _042_.n0 VGND 2.63f
C19048 _042_.t1 VGND 0.195f
C19049 _042_.n1 VGND 0.376f
C19050 _042_.t0 VGND 0.186f
C19051 _042_.t3 VGND 0.0424f
C19052 _042_.t2 VGND 0.0672f
C19053 _042_.n2 VGND 0.143f
C19054 _042_.n3 VGND 0.236f
C19055 clk.t0 VGND 0.0277f
C19056 clk.t3 VGND 0.013f
C19057 clk.t1 VGND 0.0277f
C19058 clk.t5 VGND 0.013f
C19059 clk.t2 VGND 0.0277f
C19060 clk.t6 VGND 0.013f
C19061 clk.t4 VGND 0.0277f
C19062 clk.t7 VGND 0.013f
C19063 clk.n0 VGND 0.0632f
C19064 clk.n1 VGND 0.0833f
C19065 clk.n2 VGND 0.0833f
C19066 clk.n3 VGND 0.0983f
C19067 clk.n4 VGND 1.05f
C19068 _110_.t1 VGND 0.0776f
C19069 _110_.n0 VGND 0.149f
C19070 _110_.t0 VGND 0.0738f
C19071 _110_.t5 VGND 0.0189f
C19072 _110_.t7 VGND 0.013f
C19073 _110_.n1 VGND 0.055f
C19074 _110_.n2 VGND 0.00767f
C19075 _110_.n3 VGND 0.0221f
C19076 _110_.t8 VGND 0.0133f
C19077 _110_.t4 VGND 0.0191f
C19078 _110_.n4 VGND 0.0469f
C19079 _110_.n5 VGND 0.0667f
C19080 _110_.t6 VGND 0.0189f
C19081 _110_.t3 VGND 0.013f
C19082 _110_.n6 VGND 0.055f
C19083 _110_.n7 VGND 0.0131f
C19084 _110_.n8 VGND 0.0553f
C19085 _110_.n9 VGND 0.464f
C19086 _110_.n10 VGND 0.247f
C19087 _110_.t9 VGND 0.013f
C19088 _110_.t2 VGND 0.0189f
C19089 _110_.n11 VGND 0.055f
C19090 _110_.n12 VGND 0.0138f
C19091 _110_.n13 VGND 0.916f
C19092 _110_.n14 VGND 0.296f
C19093 net20.n0 VGND -0.175f
C19094 net20.t0 VGND -0.0403f
C19095 net20.n1 VGND -0.0187f
C19096 net20.t5 VGND -0.0295f
C19097 net20.t2 VGND -0.0161f
C19098 net20.n2 VGND -0.0455f
C19099 net20.n3 VGND -0.0206f
C19100 net20.t4 VGND -0.0273f
C19101 net20.t7 VGND -0.0161f
C19102 net20.t3 VGND -0.0273f
C19103 net20.t6 VGND -0.0161f
C19104 net20.n4 VGND -0.0459f
C19105 net20.n5 VGND -0.0543f
C19106 net20.n6 VGND -0.185f
C19107 net20.n7 VGND -0.017f
C19108 net20.t1 VGND -0.0143f
C19109 net20.n8 VGND -0.0561f
C19110 _062_.n0 VGND 0.00872f
C19111 _062_.n1 VGND 0.132f
C19112 _062_.n2 VGND 0.0143f
C19113 _062_.n3 VGND 0.0114f
C19114 _062_.t4 VGND 0.0136f
C19115 _062_.t5 VGND 0.0136f
C19116 _062_.n4 VGND 0.0465f
C19117 _062_.t7 VGND 0.0209f
C19118 _062_.t6 VGND 0.0209f
C19119 _062_.n5 VGND 0.0445f
C19120 _062_.t1 VGND 0.0209f
C19121 _062_.t0 VGND 0.0209f
C19122 _062_.n6 VGND 0.0581f
C19123 _062_.n7 VGND 0.182f
C19124 _062_.t2 VGND 0.0209f
C19125 _062_.t3 VGND 0.0209f
C19126 _062_.n8 VGND 0.0442f
C19127 _062_.n9 VGND 0.091f
C19128 _062_.t10 VGND 0.0325f
C19129 _062_.t14 VGND 0.0192f
C19130 _062_.n10 VGND 0.0467f
C19131 _062_.t18 VGND 0.0325f
C19132 _062_.t8 VGND 0.0192f
C19133 _062_.n11 VGND 0.041f
C19134 _062_.n12 VGND 0.0275f
C19135 _062_.n13 VGND 0.0325f
C19136 _062_.t9 VGND 0.0346f
C19137 _062_.t11 VGND 0.0215f
C19138 _062_.n14 VGND 0.0236f
C19139 _062_.n15 VGND 0.0339f
C19140 _062_.n16 VGND 0.0208f
C19141 _062_.n17 VGND 0.197f
C19142 _062_.n18 VGND 0.00265f
C19143 _062_.t17 VGND 0.035f
C19144 _062_.t19 VGND 0.0207f
C19145 _062_.n19 VGND 0.0195f
C19146 _062_.n20 VGND 0.00356f
C19147 _062_.n21 VGND 0.0261f
C19148 _062_.n22 VGND 0.00327f
C19149 _062_.n23 VGND 0.00944f
C19150 _062_.t13 VGND 0.0154f
C19151 _062_.t15 VGND 0.0423f
C19152 _062_.n24 VGND 0.0654f
C19153 _062_.n25 VGND 0.0946f
C19154 _062_.n26 VGND 0.315f
C19155 _062_.n27 VGND 0.39f
C19156 _062_.t12 VGND 0.0283f
C19157 _062_.t16 VGND 0.0193f
C19158 _062_.n28 VGND 0.0571f
C19159 _062_.n29 VGND 0.198f
C19160 _062_.n30 VGND 0.596f
C19161 _062_.n31 VGND 0.0269f
C19162 net37.t5 VGND 0.0192f
C19163 net37.t4 VGND 0.0351f
C19164 net37.n0 VGND 0.0536f
C19165 net37.n1 VGND 0.0138f
C19166 net37.n2 VGND 0.698f
C19167 net37.t3 VGND 0.0136f
C19168 net37.t2 VGND 0.0136f
C19169 net37.n3 VGND 0.0314f
C19170 net37.n4 VGND 0.0295f
C19171 net37.n5 VGND 0.0193f
C19172 net37.t0 VGND 0.0209f
C19173 net37.t1 VGND 0.0209f
C19174 net37.n6 VGND 0.0535f
C19175 net37.n7 VGND 0.0923f
C19176 _051_.t10 VGND 0.00601f
C19177 _051_.t6 VGND 0.00601f
C19178 _051_.n0 VGND 0.0171f
C19179 _051_.t2 VGND 0.00924f
C19180 _051_.t4 VGND 0.00924f
C19181 _051_.n1 VGND 0.0248f
C19182 _051_.t11 VGND 0.00601f
C19183 _051_.t7 VGND 0.00601f
C19184 _051_.n2 VGND 0.0132f
C19185 _051_.t1 VGND 0.00924f
C19186 _051_.t0 VGND 0.00924f
C19187 _051_.n3 VGND 0.0208f
C19188 _051_.t9 VGND 0.00601f
C19189 _051_.t8 VGND 0.00601f
C19190 _051_.n4 VGND 0.0132f
C19191 _051_.n5 VGND 0.0384f
C19192 _051_.t20 VGND 0.014f
C19193 _051_.t13 VGND 0.00665f
C19194 _051_.n6 VGND 0.0505f
C19195 _051_.n7 VGND 0.00978f
C19196 _051_.t12 VGND 0.0123f
C19197 _051_.t16 VGND 0.00846f
C19198 _051_.n8 VGND 0.0303f
C19199 _051_.n9 VGND 0.0691f
C19200 _051_.t17 VGND 0.00617f
C19201 _051_.n10 VGND 0.0232f
C19202 _051_.t14 VGND 0.00857f
C19203 _051_.n11 VGND 0.0258f
C19204 _051_.n12 VGND 0.00791f
C19205 _051_.n13 VGND 0.0194f
C19206 _051_.n14 VGND 0.211f
C19207 _051_.n15 VGND 0.0859f
C19208 _051_.n16 VGND 0.00509f
C19209 _051_.n17 VGND 0.0014f
C19210 _051_.t19 VGND 0.00937f
C19211 _051_.n18 VGND 0.01f
C19212 _051_.t15 VGND 0.0153f
C19213 _051_.n19 VGND 0.0143f
C19214 _051_.n20 VGND 0.0767f
C19215 _051_.t21 VGND 0.0125f
C19216 _051_.t18 VGND 0.00633f
C19217 _051_.n21 VGND 0.0244f
C19218 _051_.n22 VGND 0.0273f
C19219 _051_.n23 VGND 0.239f
C19220 _051_.n24 VGND 0.379f
C19221 _051_.n25 VGND 0.0873f
C19222 _051_.t3 VGND 0.00924f
C19223 _051_.t5 VGND 0.00924f
C19224 _051_.n26 VGND 0.0208f
C19225 _051_.n27 VGND 0.102f
C19226 _123_.t1 VGND 0.0471f
C19227 _123_.n0 VGND 0.0384f
C19228 _123_.n1 VGND 0.0459f
C19229 _123_.n2 VGND 0.0174f
C19230 _123_.t0 VGND 0.0245f
C19231 _123_.n3 VGND 0.014f
C19232 _123_.t2 VGND 0.0264f
C19233 _123_.n4 VGND 0.0274f
C19234 _123_.n5 VGND 0.0304f
C19235 _123_.t6 VGND 0.0461f
C19236 _123_.t8 VGND 0.029f
C19237 _123_.n6 VGND 0.0656f
C19238 _123_.n7 VGND 0.0467f
C19239 _123_.t3 VGND 0.0219f
C19240 _123_.t5 VGND 0.0791f
C19241 _123_.n8 VGND 0.171f
C19242 _123_.n9 VGND 0.414f
C19243 _123_.n10 VGND 0.47f
C19244 _123_.t4 VGND 0.0461f
C19245 _123_.t7 VGND 0.029f
C19246 _123_.n11 VGND 0.0656f
C19247 _123_.n12 VGND 0.0703f
C19248 _123_.n13 VGND 0.495f
C19249 _123_.n14 VGND 0.465f
C19250 _123_.n15 VGND 0.0593f
C19251 _065_.n0 VGND 0.124f
C19252 _065_.t0 VGND 0.013f
C19253 _065_.t1 VGND 0.013f
C19254 _065_.n1 VGND 0.0262f
C19255 _065_.t13 VGND 0.0119f
C19256 _065_.t9 VGND 0.0218f
C19257 _065_.n2 VGND 0.0333f
C19258 _065_.n3 VGND 0.0086f
C19259 _065_.n4 VGND 0.0546f
C19260 _065_.t18 VGND 0.0214f
C19261 _065_.t5 VGND 0.0135f
C19262 _065_.n5 VGND 0.0424f
C19263 _065_.t8 VGND 0.0116f
C19264 _065_.t15 VGND 0.00922f
C19265 _065_.n6 VGND 0.0432f
C19266 _065_.n7 VGND 0.0327f
C19267 _065_.n8 VGND 0.197f
C19268 _065_.t6 VGND 0.0215f
C19269 _065_.t12 VGND 0.0134f
C19270 _065_.n9 VGND 0.0485f
C19271 _065_.n10 VGND 0.0401f
C19272 _065_.n11 VGND 0.492f
C19273 _065_.t10 VGND 0.0263f
C19274 _065_.t19 VGND 0.00957f
C19275 _065_.n12 VGND 0.0436f
C19276 _065_.n13 VGND 0.414f
C19277 _065_.n14 VGND 0.21f
C19278 _065_.n15 VGND 0.0706f
C19279 _065_.n16 VGND 0.00953f
C19280 _065_.n17 VGND 0.00164f
C19281 _065_.t17 VGND 0.0202f
C19282 _065_.t4 VGND 0.0119f
C19283 _065_.n18 VGND 0.0284f
C19284 _065_.t7 VGND 0.0202f
C19285 _065_.t14 VGND 0.0119f
C19286 _065_.n19 VGND 0.0234f
C19287 _065_.n20 VGND 0.00493f
C19288 _065_.n21 VGND 0.0027f
C19289 _065_.n22 VGND 0.00842f
C19290 _065_.n23 VGND 0.0105f
C19291 _065_.n24 VGND 0.0169f
C19292 _065_.n25 VGND 0.182f
C19293 _065_.t11 VGND 0.00957f
C19294 _065_.t16 VGND 0.012f
C19295 _065_.n26 VGND 0.0271f
C19296 _065_.n27 VGND 0.401f
C19297 _065_.n28 VGND 0.0645f
C19298 _065_.t3 VGND 0.00845f
C19299 _065_.t2 VGND 0.00845f
C19300 _065_.n29 VGND 0.0195f
C19301 net43.n0 VGND 0.111f
C19302 net43.n1 VGND 0.00322f
C19303 net43.n2 VGND 0.0245f
C19304 net43.n3 VGND 0.144f
C19305 net43.n4 VGND 0.00322f
C19306 net43.n5 VGND 0.0245f
C19307 net43.n6 VGND 0.021f
C19308 net43.n7 VGND 0.0918f
C19309 net43.n8 VGND 0.0245f
C19310 net43.n9 VGND 0.0156f
C19311 net43.n10 VGND 0.0156f
C19312 net43.n11 VGND 0.0156f
C19313 net43.n12 VGND 0.0254f
C19314 net43.n13 VGND 0.00493f
C19315 net43.n14 VGND 0.0254f
C19316 net43.n15 VGND 0.00493f
C19317 net43.n16 VGND 0.0254f
C19318 net43.n17 VGND 0.00493f
C19319 net43.n18 VGND 0.0254f
C19320 net43.n19 VGND 0.00493f
C19321 net43.n20 VGND 0.0254f
C19322 net43.n21 VGND 0.00493f
C19323 net43.n22 VGND 0.0254f
C19324 net43.n23 VGND 0.00493f
C19325 net43.n24 VGND 0.00583f
C19326 net43.n25 VGND 0.00824f
C19327 net43.n26 VGND 0.0178f
C19328 net43.n27 VGND 0.00824f
C19329 net43.n28 VGND 0.0178f
C19330 net43.n29 VGND 0.00824f
C19331 net43.n30 VGND 0.0178f
C19332 net43.n31 VGND 0.00335f
C19333 net43.n32 VGND 0.00335f
C19334 net43.n33 VGND 0.00335f
C19335 net43.n34 VGND 4.67e-19
C19336 net43.t6 VGND 0.00795f
C19337 net43.t7 VGND 0.00795f
C19338 net43.n35 VGND 0.0357f
C19339 net43.t4 VGND 0.00795f
C19340 net43.t5 VGND 0.00795f
C19341 net43.n36 VGND 0.0191f
C19342 net43.n37 VGND 0.0969f
C19343 net43.n38 VGND 0.00756f
C19344 net43.n39 VGND 0.00425f
C19345 net43.t8 VGND 0.0156f
C19346 net43.n40 VGND 0.0197f
C19347 net43.t17 VGND 0.0252f
C19348 net43.n41 VGND 0.00675f
C19349 net43.n42 VGND 0.031f
C19350 net43.n43 VGND 0.00508f
C19351 net43.n44 VGND 0.0681f
C19352 net43.t34 VGND 0.0298f
C19353 net43.t41 VGND 0.0118f
C19354 net43.n45 VGND 0.0605f
C19355 net43.n46 VGND 0.0492f
C19356 net43.n47 VGND 0.0244f
C19357 net43.n48 VGND 0.0434f
C19358 net43.n49 VGND 0.0351f
C19359 net43.n50 VGND 0.00425f
C19360 net43.t36 VGND 0.0156f
C19361 net43.n51 VGND 0.0197f
C19362 net43.t47 VGND 0.0252f
C19363 net43.n52 VGND 0.00675f
C19364 net43.n53 VGND 0.031f
C19365 net43.n54 VGND 0.00508f
C19366 net43.n55 VGND 0.0681f
C19367 net43.t19 VGND 0.0298f
C19368 net43.t28 VGND 0.0118f
C19369 net43.n56 VGND 0.0605f
C19370 net43.n57 VGND 0.0492f
C19371 net43.n58 VGND 0.0244f
C19372 net43.n59 VGND 0.0434f
C19373 net43.n60 VGND 0.0113f
C19374 net43.n61 VGND 0.16f
C19375 net43.n62 VGND 0.00425f
C19376 net43.t23 VGND 0.0156f
C19377 net43.n63 VGND 0.0197f
C19378 net43.t24 VGND 0.0252f
C19379 net43.n64 VGND 0.00675f
C19380 net43.n65 VGND 0.031f
C19381 net43.n66 VGND 0.004f
C19382 net43.n67 VGND 0.00516f
C19383 net43.t37 VGND 0.0298f
C19384 net43.t15 VGND 0.0118f
C19385 net43.n68 VGND 0.0605f
C19386 net43.n69 VGND 0.0492f
C19387 net43.n70 VGND 0.0693f
C19388 net43.n71 VGND 0.00756f
C19389 net43.t46 VGND 0.0298f
C19390 net43.t12 VGND 0.0118f
C19391 net43.n72 VGND 0.051f
C19392 net43.n73 VGND 0.00425f
C19393 net43.t33 VGND 0.0156f
C19394 net43.n74 VGND 0.0197f
C19395 net43.t45 VGND 0.0252f
C19396 net43.n75 VGND 0.00675f
C19397 net43.n76 VGND 0.031f
C19398 net43.n77 VGND 0.00508f
C19399 net43.n78 VGND 0.0651f
C19400 net43.n79 VGND 0.00451f
C19401 net43.n80 VGND 0.0205f
C19402 net43.n81 VGND 0.134f
C19403 net43.t31 VGND 0.0298f
C19404 net43.t43 VGND 0.0118f
C19405 net43.n82 VGND 0.051f
C19406 net43.n83 VGND 0.00425f
C19407 net43.t20 VGND 0.0156f
C19408 net43.n84 VGND 0.0197f
C19409 net43.t30 VGND 0.0252f
C19410 net43.n85 VGND 0.00675f
C19411 net43.n86 VGND 0.031f
C19412 net43.n87 VGND 0.00508f
C19413 net43.n88 VGND 0.0651f
C19414 net43.n89 VGND 0.00451f
C19415 net43.n90 VGND 0.0205f
C19416 net43.n91 VGND 0.0196f
C19417 net43.t21 VGND 0.0298f
C19418 net43.t27 VGND 0.0118f
C19419 net43.n92 VGND 0.0605f
C19420 net43.n93 VGND 0.0492f
C19421 net43.n94 VGND 0.0693f
C19422 net43.t13 VGND 0.0156f
C19423 net43.n95 VGND 0.0197f
C19424 net43.t35 VGND 0.0252f
C19425 net43.n96 VGND 0.00404f
C19426 net43.n97 VGND 0.00675f
C19427 net43.n98 VGND 0.031f
C19428 net43.n99 VGND 0.0049f
C19429 net43.n100 VGND 0.294f
C19430 net43.n101 VGND 0.224f
C19431 net43.n102 VGND 0.112f
C19432 net43.t26 VGND 0.0298f
C19433 net43.t16 VGND 0.0118f
C19434 net43.n103 VGND 0.051f
C19435 net43.n104 VGND 0.00425f
C19436 net43.t25 VGND 0.0156f
C19437 net43.n105 VGND 0.0197f
C19438 net43.t14 VGND 0.0252f
C19439 net43.n106 VGND 0.00675f
C19440 net43.n107 VGND 0.031f
C19441 net43.n108 VGND 0.00508f
C19442 net43.n109 VGND 0.0651f
C19443 net43.n110 VGND 0.00451f
C19444 net43.n111 VGND 0.0205f
C19445 net43.n112 VGND 0.0196f
C19446 net43.n113 VGND 0.00425f
C19447 net43.t42 VGND 0.0252f
C19448 net43.n114 VGND 0.0161f
C19449 net43.n115 VGND 0.00675f
C19450 net43.t22 VGND 0.0155f
C19451 net43.n116 VGND 0.0193f
C19452 net43.n117 VGND 0.0314f
C19453 net43.n118 VGND 0.004f
C19454 net43.n119 VGND 0.00516f
C19455 net43.t18 VGND 0.0118f
C19456 net43.t11 VGND 0.0298f
C19457 net43.n120 VGND 0.0605f
C19458 net43.n121 VGND 0.0492f
C19459 net43.n122 VGND 0.0693f
C19460 net43.n123 VGND 0.00425f
C19461 net43.t9 VGND 0.0156f
C19462 net43.n124 VGND 0.0197f
C19463 net43.t39 VGND 0.0252f
C19464 net43.n125 VGND 0.00675f
C19465 net43.n126 VGND 0.031f
C19466 net43.n127 VGND 0.004f
C19467 net43.n128 VGND 0.00516f
C19468 net43.t38 VGND 0.0298f
C19469 net43.t29 VGND 0.0118f
C19470 net43.n129 VGND 0.0605f
C19471 net43.n130 VGND 0.0492f
C19472 net43.n131 VGND 0.0693f
C19473 net43.n132 VGND 0.00425f
C19474 net43.t10 VGND 0.0252f
C19475 net43.t32 VGND 0.0155f
C19476 net43.n133 VGND 0.0193f
C19477 net43.t44 VGND 0.0118f
C19478 net43.t40 VGND 0.0298f
C19479 net43.n134 VGND 0.0605f
C19480 net43.n135 VGND 0.0492f
C19481 net43.n136 VGND 0.0693f
C19482 net43.n137 VGND 0.00508f
C19483 net43.n138 VGND 0.0314f
C19484 net43.n139 VGND 0.00675f
C19485 net43.n140 VGND 0.0159f
C19486 net43.n141 VGND 0.0185f
C19487 net43.n142 VGND 0.731f
C19488 net43.n143 VGND 0.497f
C19489 net43.n144 VGND 0.214f
C19490 net43.n145 VGND 0.0414f
C19491 net43.t1 VGND 0.0189f
C19492 net43.t2 VGND 0.0189f
C19493 net43.n146 VGND 0.0396f
C19494 net43.t3 VGND 0.0189f
C19495 net43.t0 VGND 0.0189f
C19496 net43.n147 VGND 0.0479f
C19497 net43.n148 VGND 0.109f
C19498 net30.t1 VGND 0.0206f
C19499 net30.t0 VGND 0.0206f
C19500 net30.n0 VGND 0.0441f
C19501 net30.t11 VGND 0.0189f
C19502 net30.t8 VGND 0.032f
C19503 net30.n1 VGND 0.0432f
C19504 net30.t7 VGND 0.0189f
C19505 net30.t5 VGND 0.032f
C19506 net30.n2 VGND 0.0432f
C19507 net30.n3 VGND 0.0212f
C19508 net30.n4 VGND 0.0233f
C19509 net30.t9 VGND 0.0235f
C19510 net30.t4 VGND 0.0282f
C19511 net30.n5 VGND 0.0702f
C19512 net30.n6 VGND 0.295f
C19513 net30.n7 VGND 0.495f
C19514 net30.t6 VGND 0.0189f
C19515 net30.t10 VGND 0.0346f
C19516 net30.n8 VGND 0.0528f
C19517 net30.n9 VGND 0.0136f
C19518 net30.n10 VGND 0.00652f
C19519 net30.n11 VGND 1.31f
C19520 net30.n12 VGND 0.0584f
C19521 net30.t3 VGND 0.00865f
C19522 net30.t2 VGND 0.00865f
C19523 net30.n13 VGND 0.0243f
C19524 net34.t7 VGND 0.011f
C19525 net34.t4 VGND 0.0201f
C19526 net34.n0 VGND 0.0307f
C19527 net34.n1 VGND 0.0106f
C19528 net34.t5 VGND 0.011f
C19529 net34.t2 VGND 0.0187f
C19530 net34.t6 VGND 0.011f
C19531 net34.t3 VGND 0.0187f
C19532 net34.n2 VGND 0.0313f
C19533 net34.n3 VGND 0.0366f
C19534 net34.n4 VGND 0.703f
C19535 net34.n5 VGND 0.845f
C19536 net34.n6 VGND 0.0253f
C19537 net34.t1 VGND 0.0195f
C19538 net34.n7 VGND 0.0302f
C19539 net34.t0 VGND 0.0183f
C19540 net34.n8 VGND 0.0128f
C19541 net34.n9 VGND 0.00291f
C19542 net34.n10 VGND 0.0148f
C19543 net34.n11 VGND 0.0265f
C19544 _048_.t1 VGND 0.00867f
C19545 _048_.t4 VGND 0.00867f
C19546 _048_.n0 VGND 0.0232f
C19547 _048_.t10 VGND 0.00564f
C19548 _048_.t7 VGND 0.00564f
C19549 _048_.n1 VGND 0.0161f
C19550 _048_.n2 VGND 0.0504f
C19551 _048_.t3 VGND 0.00867f
C19552 _048_.t0 VGND 0.00867f
C19553 _048_.n3 VGND 0.0195f
C19554 _048_.t6 VGND 0.00564f
C19555 _048_.t9 VGND 0.00564f
C19556 _048_.n4 VGND 0.0123f
C19557 _048_.t12 VGND 0.00638f
C19558 _048_.t14 VGND 0.0175f
C19559 _048_.n5 VGND 0.0305f
C19560 _048_.n6 VGND 0.0337f
C19561 _048_.t21 VGND 0.0135f
C19562 _048_.t28 VGND 0.00795f
C19563 _048_.n7 VGND 0.0196f
C19564 _048_.t29 VGND 0.0135f
C19565 _048_.t36 VGND 0.00795f
C19566 _048_.n8 VGND 0.0168f
C19567 _048_.n9 VGND 0.00931f
C19568 _048_.t37 VGND 0.0146f
C19569 _048_.t33 VGND 0.00915f
C19570 _048_.n10 VGND 0.0215f
C19571 _048_.n11 VGND 0.0115f
C19572 _048_.t30 VGND 0.00824f
C19573 _048_.t23 VGND 0.0138f
C19574 _048_.n12 VGND 0.0174f
C19575 _048_.t20 VGND 0.00824f
C19576 _048_.t32 VGND 0.0138f
C19577 _048_.n13 VGND 0.0174f
C19578 _048_.n14 VGND 0.00734f
C19579 _048_.t18 VGND 0.0143f
C19580 _048_.t22 VGND 0.00903f
C19581 _048_.n15 VGND 0.0286f
C19582 _048_.n16 VGND 0.0412f
C19583 _048_.t34 VGND 0.0135f
C19584 _048_.t16 VGND 0.00795f
C19585 _048_.t27 VGND 0.0135f
C19586 _048_.t31 VGND 0.00795f
C19587 _048_.n17 VGND 0.0226f
C19588 _048_.n18 VGND 0.0225f
C19589 _048_.n19 VGND 0.00803f
C19590 _048_.n20 VGND 0.00873f
C19591 _048_.n21 VGND 0.11f
C19592 _048_.n22 VGND 0.122f
C19593 _048_.t24 VGND 0.00807f
C19594 _048_.t26 VGND 0.00629f
C19595 _048_.n23 VGND 0.02f
C19596 _048_.n24 VGND 0.116f
C19597 _048_.n25 VGND 0.135f
C19598 _048_.t25 VGND 0.00918f
C19599 _048_.t35 VGND 0.0146f
C19600 _048_.n26 VGND 0.0203f
C19601 _048_.n27 VGND 0.116f
C19602 _048_.n28 VGND 0.134f
C19603 _048_.n29 VGND 0.133f
C19604 _048_.t17 VGND 0.00915f
C19605 _048_.t19 VGND 0.0146f
C19606 _048_.n30 VGND 0.021f
C19607 _048_.n31 VGND 0.142f
C19608 _048_.t13 VGND 0.0138f
C19609 _048_.t15 VGND 0.00603f
C19610 _048_.n32 VGND 0.0236f
C19611 _048_.n33 VGND 0.00578f
C19612 _048_.n34 VGND 0.00567f
C19613 _048_.n35 VGND 0.116f
C19614 _048_.n36 VGND 0.0686f
C19615 _048_.t11 VGND 0.00564f
C19616 _048_.t8 VGND 0.00564f
C19617 _048_.n37 VGND 0.0123f
C19618 _048_.t2 VGND 0.00867f
C19619 _048_.t5 VGND 0.00867f
C19620 _048_.n38 VGND 0.0195f
C19621 _048_.n39 VGND 0.036f
C19622 _048_.n40 VGND 0.0554f
C19623 _048_.n41 VGND 0.0863f
C19624 _063_.n0 VGND 0.0121f
C19625 _063_.n1 VGND 0.019f
C19626 _063_.t4 VGND 0.00872f
C19627 _063_.t5 VGND 0.00869f
C19628 _063_.n2 VGND 0.0184f
C19629 _063_.t16 VGND 0.0138f
C19630 _063_.t11 VGND 0.0219f
C19631 _063_.n3 VGND 0.0451f
C19632 _063_.t10 VGND 0.0207f
C19633 _063_.t12 VGND 0.0122f
C19634 _063_.n4 VGND 0.0279f
C19635 _063_.t14 VGND 0.0207f
C19636 _063_.t17 VGND 0.0122f
C19637 _063_.n5 VGND 0.0279f
C19638 _063_.n6 VGND 0.0176f
C19639 _063_.n7 VGND 0.12f
C19640 _063_.t18 VGND 0.0142f
C19641 _063_.t15 VGND 0.0223f
C19642 _063_.n8 VGND 0.0332f
C19643 _063_.n9 VGND 0.214f
C19644 _063_.t13 VGND 0.0103f
C19645 _063_.t19 VGND 0.0147f
C19646 _063_.n10 VGND 0.0367f
C19647 _063_.n11 VGND 0.0882f
C19648 _063_.n12 VGND 0.177f
C19649 _063_.n13 VGND 0.276f
C19650 _063_.n14 VGND 0.0579f
C19651 _063_.t9 VGND 0.0133f
C19652 _063_.t8 VGND 0.0133f
C19653 _063_.n15 VGND 0.0327f
C19654 _063_.t6 VGND 0.0133f
C19655 _063_.t7 VGND 0.0133f
C19656 _063_.n16 VGND 0.0449f
C19657 _063_.t1 VGND 0.0133f
C19658 _063_.t0 VGND 0.0133f
C19659 _063_.n17 VGND 0.0327f
C19660 _063_.n18 VGND 0.156f
C19661 _063_.n19 VGND 0.0927f
C19662 _063_.n20 VGND 0.0218f
C19663 _063_.t2 VGND 0.0133f
C19664 _063_.t3 VGND 0.0133f
C19665 _063_.n21 VGND 0.0316f
C19666 clknet_2_1__leaf_clk.n0 VGND 0.00948f
C19667 clknet_2_1__leaf_clk.t30 VGND 0.00536f
C19668 clknet_2_1__leaf_clk.t27 VGND 0.00536f
C19669 clknet_2_1__leaf_clk.n1 VGND 0.024f
C19670 clknet_2_1__leaf_clk.t16 VGND 0.00536f
C19671 clknet_2_1__leaf_clk.t18 VGND 0.00536f
C19672 clknet_2_1__leaf_clk.n2 VGND 0.0135f
C19673 clknet_2_1__leaf_clk.n3 VGND 0.0711f
C19674 clknet_2_1__leaf_clk.t20 VGND 0.00536f
C19675 clknet_2_1__leaf_clk.t21 VGND 0.00536f
C19676 clknet_2_1__leaf_clk.n4 VGND 0.0135f
C19677 clknet_2_1__leaf_clk.n5 VGND 0.0452f
C19678 clknet_2_1__leaf_clk.t17 VGND 0.00536f
C19679 clknet_2_1__leaf_clk.t19 VGND 0.00536f
C19680 clknet_2_1__leaf_clk.n6 VGND 0.0135f
C19681 clknet_2_1__leaf_clk.n7 VGND 0.0466f
C19682 clknet_2_1__leaf_clk.t25 VGND 0.00536f
C19683 clknet_2_1__leaf_clk.t22 VGND 0.00536f
C19684 clknet_2_1__leaf_clk.n8 VGND 0.0135f
C19685 clknet_2_1__leaf_clk.n9 VGND 0.0452f
C19686 clknet_2_1__leaf_clk.t23 VGND 0.00536f
C19687 clknet_2_1__leaf_clk.t24 VGND 0.00536f
C19688 clknet_2_1__leaf_clk.n10 VGND 0.0135f
C19689 clknet_2_1__leaf_clk.n11 VGND 0.0454f
C19690 clknet_2_1__leaf_clk.t28 VGND 0.00504f
C19691 clknet_2_1__leaf_clk.t26 VGND 0.00565f
C19692 clknet_2_1__leaf_clk.n12 VGND 0.011f
C19693 clknet_2_1__leaf_clk.n13 VGND 0.0108f
C19694 clknet_2_1__leaf_clk.n14 VGND 0.00936f
C19695 clknet_2_1__leaf_clk.t44 VGND 0.0134f
C19696 clknet_2_1__leaf_clk.t34 VGND 0.0199f
C19697 clknet_2_1__leaf_clk.n15 VGND 0.0382f
C19698 clknet_2_1__leaf_clk.n16 VGND 0.0888f
C19699 clknet_2_1__leaf_clk.t35 VGND 0.0134f
C19700 clknet_2_1__leaf_clk.t52 VGND 0.0199f
C19701 clknet_2_1__leaf_clk.n17 VGND 0.0382f
C19702 clknet_2_1__leaf_clk.n18 VGND 0.0505f
C19703 clknet_2_1__leaf_clk.n19 VGND 0.239f
C19704 clknet_2_1__leaf_clk.n20 VGND 0.00568f
C19705 clknet_2_1__leaf_clk.t46 VGND 0.0134f
C19706 clknet_2_1__leaf_clk.t40 VGND 0.0199f
C19707 clknet_2_1__leaf_clk.n21 VGND 0.0368f
C19708 clknet_2_1__leaf_clk.n22 VGND 0.0148f
C19709 clknet_2_1__leaf_clk.n23 VGND 0.00178f
C19710 clknet_2_1__leaf_clk.n24 VGND 0.0101f
C19711 clknet_2_1__leaf_clk.n25 VGND 0.0578f
C19712 clknet_2_1__leaf_clk.n26 VGND 0.15f
C19713 clknet_2_1__leaf_clk.t53 VGND 0.0134f
C19714 clknet_2_1__leaf_clk.t36 VGND 0.02f
C19715 clknet_2_1__leaf_clk.n27 VGND 0.0373f
C19716 clknet_2_1__leaf_clk.n28 VGND 0.0237f
C19717 clknet_2_1__leaf_clk.n29 VGND 0.204f
C19718 clknet_2_1__leaf_clk.t32 VGND 0.0134f
C19719 clknet_2_1__leaf_clk.t43 VGND 0.02f
C19720 clknet_2_1__leaf_clk.n30 VGND 0.0373f
C19721 clknet_2_1__leaf_clk.n31 VGND 0.0108f
C19722 clknet_2_1__leaf_clk.n32 VGND 0.197f
C19723 clknet_2_1__leaf_clk.t49 VGND 0.02f
C19724 clknet_2_1__leaf_clk.t57 VGND 0.0134f
C19725 clknet_2_1__leaf_clk.n33 VGND 0.0365f
C19726 clknet_2_1__leaf_clk.n34 VGND 0.0108f
C19727 clknet_2_1__leaf_clk.t41 VGND 0.0134f
C19728 clknet_2_1__leaf_clk.t33 VGND 0.02f
C19729 clknet_2_1__leaf_clk.n35 VGND 0.0373f
C19730 clknet_2_1__leaf_clk.n36 VGND 0.0146f
C19731 clknet_2_1__leaf_clk.t55 VGND 0.0134f
C19732 clknet_2_1__leaf_clk.t45 VGND 0.02f
C19733 clknet_2_1__leaf_clk.n37 VGND 0.0373f
C19734 clknet_2_1__leaf_clk.n38 VGND 0.0109f
C19735 clknet_2_1__leaf_clk.t37 VGND 0.0134f
C19736 clknet_2_1__leaf_clk.t54 VGND 0.02f
C19737 clknet_2_1__leaf_clk.n39 VGND 0.0373f
C19738 clknet_2_1__leaf_clk.n40 VGND 0.0434f
C19739 clknet_2_1__leaf_clk.t56 VGND 0.02f
C19740 clknet_2_1__leaf_clk.t38 VGND 0.0134f
C19741 clknet_2_1__leaf_clk.n41 VGND 0.0365f
C19742 clknet_2_1__leaf_clk.n42 VGND 0.0108f
C19743 clknet_2_1__leaf_clk.t48 VGND 0.0134f
C19744 clknet_2_1__leaf_clk.t42 VGND 0.0199f
C19745 clknet_2_1__leaf_clk.n43 VGND 0.0382f
C19746 clknet_2_1__leaf_clk.n44 VGND 0.0366f
C19747 clknet_2_1__leaf_clk.t51 VGND 0.0134f
C19748 clknet_2_1__leaf_clk.t47 VGND 0.0199f
C19749 clknet_2_1__leaf_clk.n45 VGND 0.0382f
C19750 clknet_2_1__leaf_clk.n46 VGND 0.165f
C19751 clknet_2_1__leaf_clk.n47 VGND 0.268f
C19752 clknet_2_1__leaf_clk.n48 VGND 0.202f
C19753 clknet_2_1__leaf_clk.n49 VGND 0.16f
C19754 clknet_2_1__leaf_clk.n50 VGND 0.282f
C19755 clknet_2_1__leaf_clk.t50 VGND 0.0134f
C19756 clknet_2_1__leaf_clk.t39 VGND 0.02f
C19757 clknet_2_1__leaf_clk.n51 VGND 0.0373f
C19758 clknet_2_1__leaf_clk.n52 VGND 0.0109f
C19759 clknet_2_1__leaf_clk.n53 VGND 0.279f
C19760 clknet_2_1__leaf_clk.n54 VGND 0.251f
C19761 clknet_2_1__leaf_clk.n55 VGND 0.145f
C19762 clknet_2_1__leaf_clk.n56 VGND 0.176f
C19763 clknet_2_1__leaf_clk.n57 VGND 0.0101f
C19764 clknet_2_1__leaf_clk.n58 VGND 0.0966f
C19765 clknet_2_1__leaf_clk.n59 VGND 0.0058f
C19766 clknet_2_1__leaf_clk.n60 VGND 0.00783f
C19767 clknet_2_1__leaf_clk.n61 VGND 0.0227f
C19768 clknet_2_1__leaf_clk.t29 VGND 0.00536f
C19769 clknet_2_1__leaf_clk.t31 VGND 0.00536f
C19770 clknet_2_1__leaf_clk.n62 VGND 0.0129f
C19771 clknet_2_1__leaf_clk.n63 VGND 0.0523f
C19772 clknet_2_1__leaf_clk.t0 VGND 0.0128f
C19773 clknet_2_1__leaf_clk.t2 VGND 0.0128f
C19774 clknet_2_1__leaf_clk.n64 VGND 0.0275f
C19775 clknet_2_1__leaf_clk.t1 VGND 0.0128f
C19776 clknet_2_1__leaf_clk.t14 VGND 0.0128f
C19777 clknet_2_1__leaf_clk.n65 VGND 0.0378f
C19778 clknet_2_1__leaf_clk.t3 VGND 0.0128f
C19779 clknet_2_1__leaf_clk.t5 VGND 0.0128f
C19780 clknet_2_1__leaf_clk.n66 VGND 0.0282f
C19781 clknet_2_1__leaf_clk.n67 VGND 0.116f
C19782 clknet_2_1__leaf_clk.t7 VGND 0.0128f
C19783 clknet_2_1__leaf_clk.t8 VGND 0.0128f
C19784 clknet_2_1__leaf_clk.n68 VGND 0.0282f
C19785 clknet_2_1__leaf_clk.n69 VGND 0.0693f
C19786 clknet_2_1__leaf_clk.t4 VGND 0.0128f
C19787 clknet_2_1__leaf_clk.t6 VGND 0.0128f
C19788 clknet_2_1__leaf_clk.n70 VGND 0.0282f
C19789 clknet_2_1__leaf_clk.n71 VGND 0.069f
C19790 clknet_2_1__leaf_clk.t12 VGND 0.0128f
C19791 clknet_2_1__leaf_clk.t9 VGND 0.0128f
C19792 clknet_2_1__leaf_clk.n72 VGND 0.0282f
C19793 clknet_2_1__leaf_clk.n73 VGND 0.069f
C19794 clknet_2_1__leaf_clk.t10 VGND 0.0128f
C19795 clknet_2_1__leaf_clk.t11 VGND 0.0128f
C19796 clknet_2_1__leaf_clk.n74 VGND 0.0282f
C19797 clknet_2_1__leaf_clk.n75 VGND 0.0693f
C19798 clknet_2_1__leaf_clk.t13 VGND 0.0128f
C19799 clknet_2_1__leaf_clk.t15 VGND 0.0128f
C19800 clknet_2_1__leaf_clk.n76 VGND 0.0282f
C19801 clknet_2_1__leaf_clk.n77 VGND 0.0596f
C19802 clknet_2_1__leaf_clk.n78 VGND 0.0399f
C19803 VPWR.n0 VGND 6.83e-19
C19804 VPWR.n1 VGND 5.12e-19
C19805 VPWR.n2 VGND 5.05e-19
C19806 VPWR.n3 VGND 0.00138f
C19807 VPWR.n4 VGND 5.48e-19
C19808 VPWR.n5 VGND 9.06e-19
C19809 VPWR.n6 VGND 6.54e-19
C19810 VPWR.n7 VGND 8.67e-19
C19811 VPWR.n8 VGND 4.11e-19
C19812 VPWR.n9 VGND 4.11e-19
C19813 VPWR.n10 VGND 7.39e-19
C19814 VPWR.n11 VGND 5.19e-19
C19815 VPWR.n12 VGND 7.39e-19
C19816 VPWR.n13 VGND 4.11e-19
C19817 VPWR.n14 VGND 4.11e-19
C19818 VPWR.n15 VGND 8.67e-19
C19819 VPWR.n16 VGND 6.54e-19
C19820 VPWR.n17 VGND 9.06e-19
C19821 VPWR.n18 VGND 0.00626f
C19822 VPWR.n20 VGND 0.0057f
C19823 VPWR.n21 VGND 6.54e-19
C19824 VPWR.n22 VGND 9.06e-19
C19825 VPWR.n23 VGND 0.00139f
C19826 VPWR.n24 VGND 5.48e-19
C19827 VPWR.t878 VGND 0.00654f
C19828 VPWR.n26 VGND 0.0109f
C19829 VPWR.n27 VGND 8.11e-19
C19830 VPWR.n28 VGND 3.95e-19
C19831 VPWR.n29 VGND 6.26e-19
C19832 VPWR.t1347 VGND 0.00102f
C19833 VPWR.t1609 VGND 0.00154f
C19834 VPWR.n30 VGND 0.00486f
C19835 VPWR.n31 VGND 0.00622f
C19836 VPWR.n32 VGND 0.0218f
C19837 VPWR.n33 VGND 0.0031f
C19838 VPWR.t242 VGND 0.00387f
C19839 VPWR.t1556 VGND 0.00676f
C19840 VPWR.t2294 VGND 0.00631f
C19841 VPWR.t3019 VGND 0.00239f
C19842 VPWR.n34 VGND 0.00417f
C19843 VPWR.n35 VGND 0.00589f
C19844 VPWR.t2296 VGND 0.00632f
C19845 VPWR.n36 VGND 0.007f
C19846 VPWR.t1378 VGND 6.73e-19
C19847 VPWR.t1558 VGND 0.00127f
C19848 VPWR.n37 VGND 0.00203f
C19849 VPWR.t618 VGND 0.00387f
C19850 VPWR.t3569 VGND 0.0179f
C19851 VPWR.n38 VGND 0.0133f
C19852 VPWR.n39 VGND 0.0103f
C19853 VPWR.n40 VGND 0.0173f
C19854 VPWR.n41 VGND 0.00493f
C19855 VPWR.t619 VGND 0.00387f
C19856 VPWR.n42 VGND 0.00837f
C19857 VPWR.t256 VGND 0.00387f
C19858 VPWR.n43 VGND 0.00493f
C19859 VPWR.t2870 VGND 0.00234f
C19860 VPWR.t3439 VGND 0.0179f
C19861 VPWR.n44 VGND 0.0173f
C19862 VPWR.n45 VGND 0.0103f
C19863 VPWR.n46 VGND 0.00829f
C19864 VPWR.n47 VGND 0.00941f
C19865 VPWR.t257 VGND 0.00387f
C19866 VPWR.n48 VGND 0.00695f
C19867 VPWR.t1172 VGND 0.00102f
C19868 VPWR.t1828 VGND 0.00102f
C19869 VPWR.n49 VGND 0.00221f
C19870 VPWR.t3110 VGND 0.00184f
C19871 VPWR.t1349 VGND 0.00166f
C19872 VPWR.n50 VGND 0.0036f
C19873 VPWR.n51 VGND 0.0082f
C19874 VPWR.n52 VGND 0.00525f
C19875 VPWR.t3027 VGND 0.00102f
C19876 VPWR.t2247 VGND 0.00154f
C19877 VPWR.n53 VGND 0.00483f
C19878 VPWR.n54 VGND 0.0127f
C19879 VPWR.n55 VGND 0.00927f
C19880 VPWR.n56 VGND 0.0133f
C19881 VPWR.t565 VGND 0.00387f
C19882 VPWR.n57 VGND 0.00837f
C19883 VPWR.t228 VGND 0.0462f
C19884 VPWR.t3245 VGND 0.0253f
C19885 VPWR.t3247 VGND 0.0198f
C19886 VPWR.t1882 VGND 0.0109f
C19887 VPWR.t2104 VGND 0.0052f
C19888 VPWR.t1309 VGND 0.0154f
C19889 VPWR.t421 VGND 0.0389f
C19890 VPWR.t935 VGND 0.0361f
C19891 VPWR.t3220 VGND 0.021f
C19892 VPWR.t883 VGND 0.0166f
C19893 VPWR.t1308 VGND 0.0121f
C19894 VPWR.t1030 VGND 0.00604f
C19895 VPWR.t2739 VGND 0.0151f
C19896 VPWR.t1363 VGND 0.0116f
C19897 VPWR.t2899 VGND 0.0233f
C19898 VPWR.t3024 VGND 0.0242f
C19899 VPWR.t2668 VGND 0.0149f
C19900 VPWR.t3099 VGND 0.0166f
C19901 VPWR.t1307 VGND 0.0208f
C19902 VPWR.t3219 VGND 0.0191f
C19903 VPWR.t2650 VGND 0.0322f
C19904 VPWR.t2747 VGND 0.0322f
C19905 VPWR.t1630 VGND 0.0196f
C19906 VPWR.t451 VGND 0.0361f
C19907 VPWR.t2648 VGND 0.0512f
C19908 VPWR.t671 VGND 0.0339f
C19909 VPWR.n58 VGND 0.0392f
C19910 VPWR.t672 VGND 0.00387f
C19911 VPWR.n59 VGND 0.00493f
C19912 VPWR.t3557 VGND 0.0179f
C19913 VPWR.n60 VGND 0.0173f
C19914 VPWR.n61 VGND 0.0103f
C19915 VPWR.t453 VGND 0.00387f
C19916 VPWR.n62 VGND 0.00837f
C19917 VPWR.n63 VGND 0.00186f
C19918 VPWR.t884 VGND 0.00654f
C19919 VPWR.n64 VGND 0.0108f
C19920 VPWR.t936 VGND 0.00235f
C19921 VPWR.t3495 VGND 0.00911f
C19922 VPWR.t422 VGND 0.00391f
C19923 VPWR.n65 VGND 0.0253f
C19924 VPWR.t423 VGND 0.00391f
C19925 VPWR.n67 VGND 0.0138f
C19926 VPWR.n68 VGND 0.0115f
C19927 VPWR.t1310 VGND 0.00102f
C19928 VPWR.t2105 VGND 0.00102f
C19929 VPWR.n69 VGND 0.00221f
C19930 VPWR.n70 VGND 0.00572f
C19931 VPWR.t1883 VGND 0.00137f
C19932 VPWR.t3248 VGND -2.18e-20
C19933 VPWR.n71 VGND 0.00629f
C19934 VPWR.n72 VGND 0.00755f
C19935 VPWR.t3246 VGND 0.00663f
C19936 VPWR.n73 VGND 0.00884f
C19937 VPWR.t3399 VGND 0.00911f
C19938 VPWR.t230 VGND 0.00391f
C19939 VPWR.n74 VGND 0.0253f
C19940 VPWR.t229 VGND 0.00391f
C19941 VPWR.n76 VGND 0.0138f
C19942 VPWR.t3339 VGND 0.00911f
C19943 VPWR.t699 VGND 0.00391f
C19944 VPWR.n77 VGND 0.0253f
C19945 VPWR.t700 VGND 0.00391f
C19946 VPWR.n79 VGND 0.0138f
C19947 VPWR.n80 VGND 0.0109f
C19948 VPWR.n81 VGND 0.00444f
C19949 VPWR.n82 VGND 0.00333f
C19950 VPWR.n83 VGND 0.00121f
C19951 VPWR.n84 VGND 0.00393f
C19952 VPWR.n85 VGND 0.00262f
C19953 VPWR.n86 VGND 0.00179f
C19954 VPWR.n87 VGND 0.00444f
C19955 VPWR.n88 VGND 0.00393f
C19956 VPWR.n89 VGND 0.00146f
C19957 VPWR.n90 VGND 0.00473f
C19958 VPWR.n91 VGND 0.00182f
C19959 VPWR.n92 VGND 0.00199f
C19960 VPWR.n93 VGND 0.00109f
C19961 VPWR.t1364 VGND 6.73e-19
C19962 VPWR.t2740 VGND 9.96e-19
C19963 VPWR.n94 VGND 0.0018f
C19964 VPWR.n95 VGND 0.00483f
C19965 VPWR.n96 VGND 0.00103f
C19966 VPWR.n97 VGND 0.0031f
C19967 VPWR.n98 VGND 0.00155f
C19968 VPWR.n99 VGND 0.00524f
C19969 VPWR.t3100 VGND 0.00184f
C19970 VPWR.t3025 VGND 0.00166f
C19971 VPWR.n100 VGND 0.00358f
C19972 VPWR.t2669 VGND 0.00453f
C19973 VPWR.n101 VGND 0.00559f
C19974 VPWR.n102 VGND 0.00226f
C19975 VPWR.n103 VGND 9.58e-19
C19976 VPWR.n104 VGND 0.00524f
C19977 VPWR.n105 VGND 0.00393f
C19978 VPWR.n106 VGND 0.00173f
C19979 VPWR.n107 VGND 0.00525f
C19980 VPWR.n108 VGND 0.0031f
C19981 VPWR.t2748 VGND 6.73e-19
C19982 VPWR.t2651 VGND 0.00127f
C19983 VPWR.n109 VGND 0.00203f
C19984 VPWR.n110 VGND 0.00368f
C19985 VPWR.n111 VGND 0.0059f
C19986 VPWR.n112 VGND 0.0123f
C19987 VPWR.n113 VGND 0.00387f
C19988 VPWR.n114 VGND 0.00203f
C19989 VPWR.n115 VGND 0.00156f
C19990 VPWR.n116 VGND 4.27e-19
C19991 VPWR.n117 VGND 8.54e-20
C19992 VPWR.n118 VGND 0.0012f
C19993 VPWR.n119 VGND 0.00673f
C19994 VPWR.n120 VGND 4.27e-19
C19995 VPWR.n121 VGND 6.83e-19
C19996 VPWR.n122 VGND 3.7e-19
C19997 VPWR.n123 VGND 9.68e-19
C19998 VPWR.n124 VGND 9.96e-19
C19999 VPWR.n125 VGND 5.41e-19
C20000 VPWR.n126 VGND 7.4e-19
C20001 VPWR.n127 VGND 0.00127f
C20002 VPWR.n128 VGND 0.00665f
C20003 VPWR.n129 VGND 3.42e-19
C20004 VPWR.n130 VGND 2.56e-19
C20005 VPWR.n131 VGND 4.27e-19
C20006 VPWR.n132 VGND 9.68e-19
C20007 VPWR.n133 VGND 9.96e-19
C20008 VPWR.n134 VGND 3.13e-19
C20009 VPWR.n135 VGND 4.84e-19
C20010 VPWR.n136 VGND 6.83e-19
C20011 VPWR.n137 VGND 7.73e-19
C20012 VPWR.n138 VGND 2.84e-19
C20013 VPWR.n139 VGND 0.00123f
C20014 VPWR.n140 VGND 3.95e-19
C20015 VPWR.n141 VGND 5.05e-19
C20016 VPWR.n142 VGND 5.05e-19
C20017 VPWR.n143 VGND 9.06e-19
C20018 VPWR.n144 VGND 9e-19
C20019 VPWR.n145 VGND 0.00138f
C20020 VPWR.n146 VGND 6.14e-19
C20021 VPWR.n147 VGND 5.48e-19
C20022 VPWR.n148 VGND 0.00138f
C20023 VPWR.n149 VGND 6.54e-19
C20024 VPWR.n150 VGND 8.67e-19
C20025 VPWR.n151 VGND 7.39e-19
C20026 VPWR.n152 VGND 4.11e-19
C20027 VPWR.n153 VGND 5.27e-19
C20028 VPWR.n154 VGND 3.73e-19
C20029 VPWR.n155 VGND 2.41e-19
C20030 VPWR.n156 VGND 4.83e-19
C20031 VPWR.n157 VGND 4.17e-19
C20032 VPWR.n158 VGND 4.83e-19
C20033 VPWR.n159 VGND 4.61e-19
C20034 VPWR.n160 VGND 4.61e-19
C20035 VPWR.n161 VGND 4.11e-19
C20036 VPWR.n163 VGND 0.0581f
C20037 VPWR.n164 VGND 1.01f
C20038 VPWR.n165 VGND 0.0452f
C20039 VPWR.n166 VGND 0.0057f
C20040 VPWR.n167 VGND 6.54e-19
C20041 VPWR.n168 VGND 8.67e-19
C20042 VPWR.n169 VGND 6.14e-19
C20043 VPWR.n170 VGND 4.39e-19
C20044 VPWR.n171 VGND 1.76e-19
C20045 VPWR.n172 VGND 4.83e-19
C20046 VPWR.n173 VGND 2.41e-19
C20047 VPWR.n174 VGND 3.73e-19
C20048 VPWR.n175 VGND 3.07e-19
C20049 VPWR.n176 VGND 4.11e-19
C20050 VPWR.n177 VGND 4.11e-19
C20051 VPWR.n178 VGND 7.39e-19
C20052 VPWR.n179 VGND 5.19e-19
C20053 VPWR.n180 VGND 7.39e-19
C20054 VPWR.n181 VGND 4.11e-19
C20055 VPWR.n182 VGND 5.71e-19
C20056 VPWR.n183 VGND 3.29e-19
C20057 VPWR.n184 VGND 3.95e-19
C20058 VPWR.n185 VGND 4.17e-19
C20059 VPWR.n186 VGND 2.85e-19
C20060 VPWR.n187 VGND 4.17e-19
C20061 VPWR.n188 VGND 6.26e-19
C20062 VPWR.n189 VGND 3.95e-19
C20063 VPWR.n190 VGND 8.11e-19
C20064 VPWR.n191 VGND 3.95e-19
C20065 VPWR.n192 VGND 6.26e-19
C20066 VPWR.t576 VGND 0.00387f
C20067 VPWR.n193 VGND 0.0107f
C20068 VPWR.n194 VGND 0.00199f
C20069 VPWR.t2491 VGND 0.00676f
C20070 VPWR.n195 VGND 0.0119f
C20071 VPWR.n196 VGND 0.00646f
C20072 VPWR.t2425 VGND 0.00634f
C20073 VPWR.n197 VGND 0.0117f
C20074 VPWR.n198 VGND 0.0169f
C20075 VPWR.t2423 VGND 0.00647f
C20076 VPWR.n199 VGND 0.00688f
C20077 VPWR.n200 VGND 9.25e-19
C20078 VPWR.n201 VGND 3.95e-19
C20079 VPWR.n202 VGND 5.05e-19
C20080 VPWR.n203 VGND 5.05e-19
C20081 VPWR.n204 VGND 9.06e-19
C20082 VPWR.n205 VGND 9e-19
C20083 VPWR.t850 VGND 0.00166f
C20084 VPWR.t3023 VGND 0.00166f
C20085 VPWR.n206 VGND 0.00381f
C20086 VPWR.n207 VGND 0.00759f
C20087 VPWR.t206 VGND 0.00387f
C20088 VPWR.t3423 VGND 0.0231f
C20089 VPWR.n208 VGND 0.0138f
C20090 VPWR.n209 VGND 0.0384f
C20091 VPWR.n210 VGND 0.00837f
C20092 VPWR.n211 VGND 0.00525f
C20093 VPWR.t207 VGND 0.00387f
C20094 VPWR.n212 VGND 0.00837f
C20095 VPWR.t898 VGND 0.00137f
C20096 VPWR.t2701 VGND -2.18e-20
C20097 VPWR.n213 VGND 0.00629f
C20098 VPWR.n214 VGND 0.00755f
C20099 VPWR.t1336 VGND 0.00102f
C20100 VPWR.t2088 VGND 0.00102f
C20101 VPWR.n215 VGND 0.00221f
C20102 VPWR.t2699 VGND 0.00663f
C20103 VPWR.n216 VGND 0.00884f
C20104 VPWR.t3585 VGND 0.00911f
C20105 VPWR.t722 VGND 0.00391f
C20106 VPWR.n217 VGND 0.0253f
C20107 VPWR.t721 VGND 0.00391f
C20108 VPWR.n219 VGND 0.0138f
C20109 VPWR.t3520 VGND 0.00911f
C20110 VPWR.t478 VGND 0.00391f
C20111 VPWR.n220 VGND 0.0253f
C20112 VPWR.t479 VGND 0.00391f
C20113 VPWR.n222 VGND 0.0138f
C20114 VPWR.n223 VGND 0.0109f
C20115 VPWR.n224 VGND 0.00444f
C20116 VPWR.n225 VGND 0.00333f
C20117 VPWR.n226 VGND 0.00121f
C20118 VPWR.n227 VGND 0.00393f
C20119 VPWR.n228 VGND 0.00262f
C20120 VPWR.n229 VGND 0.00179f
C20121 VPWR.n230 VGND 0.00599f
C20122 VPWR.n231 VGND 0.00483f
C20123 VPWR.n232 VGND 0.0031f
C20124 VPWR.n233 VGND 0.0119f
C20125 VPWR.n234 VGND 0.00524f
C20126 VPWR.t2188 VGND 0.00234f
C20127 VPWR.n235 VGND 0.00986f
C20128 VPWR.n236 VGND 0.00829f
C20129 VPWR.n237 VGND 0.00524f
C20130 VPWR.n238 VGND 0.00524f
C20131 VPWR.n239 VGND 0.00524f
C20132 VPWR.n240 VGND 0.00393f
C20133 VPWR.n241 VGND 0.00199f
C20134 VPWR.n242 VGND 9.6e-19
C20135 VPWR.t2750 VGND 6.73e-19
C20136 VPWR.t1182 VGND 9.96e-19
C20137 VPWR.n243 VGND 0.0018f
C20138 VPWR.n244 VGND 0.00483f
C20139 VPWR.n245 VGND 0.00103f
C20140 VPWR.n246 VGND 0.0031f
C20141 VPWR.t1210 VGND 0.00587f
C20142 VPWR.n247 VGND 0.00681f
C20143 VPWR.n248 VGND 9.38e-19
C20144 VPWR.n249 VGND 0.00524f
C20145 VPWR.t2878 VGND 0.00453f
C20146 VPWR.n250 VGND 0.00561f
C20147 VPWR.n251 VGND 0.00123f
C20148 VPWR.n252 VGND 0.00524f
C20149 VPWR.n253 VGND 0.0015f
C20150 VPWR.n254 VGND 0.00524f
C20151 VPWR.n255 VGND 0.00524f
C20152 VPWR.n256 VGND 0.00116f
C20153 VPWR.n257 VGND 0.00367f
C20154 VPWR.n258 VGND 9.06e-19
C20155 VPWR.n259 VGND 0.00112f
C20156 VPWR.n260 VGND 4.27e-19
C20157 VPWR.n261 VGND 0.0012f
C20158 VPWR.n262 VGND 4.55e-19
C20159 VPWR.t1965 VGND 0.00239f
C20160 VPWR.n263 VGND 0.00784f
C20161 VPWR.n264 VGND 0.00202f
C20162 VPWR.n265 VGND 4.84e-19
C20163 VPWR.n266 VGND 6.83e-19
C20164 VPWR.n267 VGND 4.84e-19
C20165 VPWR.n268 VGND 3.13e-19
C20166 VPWR.n269 VGND 9.96e-19
C20167 VPWR.n270 VGND 0.00426f
C20168 VPWR.n271 VGND 9.68e-19
C20169 VPWR.n272 VGND 4.27e-19
C20170 VPWR.n273 VGND 2.56e-19
C20171 VPWR.n274 VGND 0.00127f
C20172 VPWR.n275 VGND 0.00643f
C20173 VPWR.n276 VGND 3.42e-19
C20174 VPWR.n277 VGND 7.4e-19
C20175 VPWR.n278 VGND 5.41e-19
C20176 VPWR.n279 VGND 9.96e-19
C20177 VPWR.n280 VGND 9.68e-19
C20178 VPWR.n281 VGND 3.7e-19
C20179 VPWR.n282 VGND 6.83e-19
C20180 VPWR.t65 VGND 0.00387f
C20181 VPWR.n283 VGND 0.008f
C20182 VPWR.n284 VGND 8.97e-19
C20183 VPWR.n285 VGND 4.48e-19
C20184 VPWR.n286 VGND 4.27e-19
C20185 VPWR.n287 VGND 8.54e-20
C20186 VPWR.n288 VGND 4.27e-19
C20187 VPWR.t3118 VGND 6.73e-19
C20188 VPWR.t2111 VGND 0.00127f
C20189 VPWR.n289 VGND 0.00196f
C20190 VPWR.n290 VGND 0.00208f
C20191 VPWR.n291 VGND 0.00161f
C20192 VPWR.n292 VGND 0.00192f
C20193 VPWR.n293 VGND 0.00149f
C20194 VPWR.n294 VGND 4.84e-19
C20195 VPWR.n295 VGND 8.26e-19
C20196 VPWR.n296 VGND 0.00138f
C20197 VPWR.n297 VGND 6.14e-19
C20198 VPWR.n298 VGND 5.48e-19
C20199 VPWR.n299 VGND 0.00138f
C20200 VPWR.n300 VGND 6.54e-19
C20201 VPWR.n301 VGND 8.67e-19
C20202 VPWR.n302 VGND 5.27e-19
C20203 VPWR.n303 VGND 3.73e-19
C20204 VPWR.n304 VGND 2.41e-19
C20205 VPWR.n305 VGND 4.83e-19
C20206 VPWR.n306 VGND 5.71e-19
C20207 VPWR.n307 VGND 4.17e-19
C20208 VPWR.n308 VGND 4.83e-19
C20209 VPWR.n309 VGND 4.61e-19
C20210 VPWR.n310 VGND 4.61e-19
C20211 VPWR.n311 VGND 5.19e-19
C20212 VPWR.n312 VGND 7.39e-19
C20213 VPWR.n313 VGND 4.11e-19
C20214 VPWR.n314 VGND 4.11e-19
C20215 VPWR.n316 VGND 0.0057f
C20216 VPWR.n317 VGND 6.54e-19
C20217 VPWR.n318 VGND 8.67e-19
C20218 VPWR.n319 VGND 3.51e-19
C20219 VPWR.n320 VGND 4.61e-19
C20220 VPWR.n321 VGND 5.27e-19
C20221 VPWR.n322 VGND 2.85e-19
C20222 VPWR.n323 VGND 2.85e-19
C20223 VPWR.n324 VGND 4.17e-19
C20224 VPWR.n325 VGND 4.11e-19
C20225 VPWR.n326 VGND 4.11e-19
C20226 VPWR.n327 VGND 7.39e-19
C20227 VPWR.n328 VGND 5.19e-19
C20228 VPWR.n329 VGND 7.39e-19
C20229 VPWR.n330 VGND 4.11e-19
C20230 VPWR.n331 VGND 5.27e-19
C20231 VPWR.n332 VGND 3.73e-19
C20232 VPWR.n333 VGND 2.41e-19
C20233 VPWR.n334 VGND 4.83e-19
C20234 VPWR.n335 VGND 4.17e-19
C20235 VPWR.n336 VGND 4.84e-19
C20236 VPWR.t3474 VGND 0.0289f
C20237 VPWR.t561 VGND 0.00387f
C20238 VPWR.n337 VGND 0.0604f
C20239 VPWR.n338 VGND 0.0146f
C20240 VPWR.n339 VGND 3.42e-19
C20241 VPWR.n340 VGND 6.26e-19
C20242 VPWR.n341 VGND 3.95e-19
C20243 VPWR.n342 VGND 5.05e-19
C20244 VPWR.n343 VGND 5.05e-19
C20245 VPWR.n344 VGND 0.00139f
C20246 VPWR.n345 VGND 0.0057f
C20247 VPWR.n346 VGND 6.54e-19
C20248 VPWR.n347 VGND 8.67e-19
C20249 VPWR.n348 VGND 4.61e-19
C20250 VPWR.n349 VGND 5.27e-19
C20251 VPWR.t2746 VGND 6.73e-19
C20252 VPWR.t2007 VGND 0.00127f
C20253 VPWR.n350 VGND 0.00207f
C20254 VPWR.n351 VGND 0.0048f
C20255 VPWR.t2005 VGND 0.00692f
C20256 VPWR.n352 VGND 0.00156f
C20257 VPWR.t3108 VGND 0.00184f
C20258 VPWR.t3189 VGND 0.00166f
C20259 VPWR.n353 VGND 0.00362f
C20260 VPWR.n354 VGND 0.00387f
C20261 VPWR.t1733 VGND 0.025f
C20262 VPWR.t1734 VGND 0.00676f
C20263 VPWR.n355 VGND 0.00938f
C20264 VPWR.n356 VGND 6.26e-19
C20265 VPWR.n357 VGND 5.05e-19
C20266 VPWR.n358 VGND 8.67e-19
C20267 VPWR.n359 VGND 6.54e-19
C20268 VPWR.n360 VGND 9.06e-19
C20269 VPWR.n362 VGND 0.071f
C20270 VPWR.n363 VGND 1.01f
C20271 VPWR.n364 VGND 0.0057f
C20272 VPWR.n365 VGND 6.54e-19
C20273 VPWR.n366 VGND 8.67e-19
C20274 VPWR.n367 VGND 3.51e-19
C20275 VPWR.n368 VGND 4.61e-19
C20276 VPWR.n369 VGND 5.27e-19
C20277 VPWR.n370 VGND 2.85e-19
C20278 VPWR.n371 VGND 2.85e-19
C20279 VPWR.n372 VGND 4.17e-19
C20280 VPWR.n373 VGND 4.11e-19
C20281 VPWR.n374 VGND 4.11e-19
C20282 VPWR.n375 VGND 7.39e-19
C20283 VPWR.n376 VGND 5.19e-19
C20284 VPWR.n377 VGND 7.39e-19
C20285 VPWR.n378 VGND 4.11e-19
C20286 VPWR.n379 VGND 4.83e-19
C20287 VPWR.n380 VGND 4.17e-19
C20288 VPWR.n381 VGND 4.84e-19
C20289 VPWR.t1796 VGND 0.00524f
C20290 VPWR.t3491 VGND 0.0179f
C20291 VPWR.n382 VGND 0.0173f
C20292 VPWR.n383 VGND 0.00351f
C20293 VPWR.n384 VGND 0.0108f
C20294 VPWR.n385 VGND 0.0132f
C20295 VPWR.t38 VGND 0.00387f
C20296 VPWR.n386 VGND 0.00837f
C20297 VPWR.n387 VGND 0.00524f
C20298 VPWR.n388 VGND 3.42e-19
C20299 VPWR.n389 VGND 6.26e-19
C20300 VPWR.n390 VGND 3.95e-19
C20301 VPWR.n391 VGND 5.05e-19
C20302 VPWR.n392 VGND 5.05e-19
C20303 VPWR.n393 VGND 0.00139f
C20304 VPWR.n395 VGND 8.67e-19
C20305 VPWR.n396 VGND 6.54e-19
C20306 VPWR.n397 VGND 9.06e-19
C20307 VPWR.n398 VGND 3.29e-19
C20308 VPWR.n399 VGND 4.39e-19
C20309 VPWR.n400 VGND 9e-19
C20310 VPWR.t396 VGND 0.0046f
C20311 VPWR.n401 VGND 0.00407f
C20312 VPWR.t3218 VGND 0.00136f
C20313 VPWR.t1812 VGND 0.00136f
C20314 VPWR.n402 VGND 0.00328f
C20315 VPWR.n403 VGND 0.0079f
C20316 VPWR.t3468 VGND 0.0289f
C20317 VPWR.t607 VGND 0.00387f
C20318 VPWR.n404 VGND 0.0604f
C20319 VPWR.n405 VGND 0.0146f
C20320 VPWR.n406 VGND 0.0117f
C20321 VPWR.t608 VGND 0.00387f
C20322 VPWR.n407 VGND 0.00837f
C20323 VPWR.t1300 VGND 0.00102f
C20324 VPWR.t1768 VGND 0.00102f
C20325 VPWR.n408 VGND 0.00221f
C20326 VPWR.n409 VGND 0.00563f
C20327 VPWR.t3166 VGND 0.00137f
C20328 VPWR.t2770 VGND -2.18e-20
C20329 VPWR.n410 VGND 0.00629f
C20330 VPWR.n411 VGND 0.00759f
C20331 VPWR.t2772 VGND 0.00663f
C20332 VPWR.n412 VGND 0.00848f
C20333 VPWR.t3446 VGND 0.00911f
C20334 VPWR.t538 VGND 0.00391f
C20335 VPWR.n413 VGND 0.0253f
C20336 VPWR.t537 VGND 0.00391f
C20337 VPWR.n415 VGND 0.0138f
C20338 VPWR.t3394 VGND 0.00911f
C20339 VPWR.t137 VGND 0.00391f
C20340 VPWR.n416 VGND 0.0253f
C20341 VPWR.t138 VGND 0.00391f
C20342 VPWR.n418 VGND 0.0138f
C20343 VPWR.n419 VGND 0.0109f
C20344 VPWR.n420 VGND 0.00444f
C20345 VPWR.n421 VGND 0.0031f
C20346 VPWR.n422 VGND 0.00524f
C20347 VPWR.n423 VGND 0.00475f
C20348 VPWR.n424 VGND 0.00179f
C20349 VPWR.n425 VGND 0.00123f
C20350 VPWR.t1629 VGND 0.00235f
C20351 VPWR.n426 VGND 0.00646f
C20352 VPWR.n427 VGND 0.00201f
C20353 VPWR.n428 VGND 0.0031f
C20354 VPWR.n429 VGND 0.0133f
C20355 VPWR.n430 VGND 0.00524f
C20356 VPWR.n431 VGND 0.0138f
C20357 VPWR.n432 VGND 0.00524f
C20358 VPWR.n433 VGND 0.0113f
C20359 VPWR.n434 VGND 0.0104f
C20360 VPWR.n435 VGND 0.00903f
C20361 VPWR.t2504 VGND 6.73e-19
C20362 VPWR.t3202 VGND 9.96e-19
C20363 VPWR.n436 VGND 0.00176f
C20364 VPWR.t1617 VGND 0.00453f
C20365 VPWR.n437 VGND 0.00968f
C20366 VPWR.n438 VGND 0.00996f
C20367 VPWR.n439 VGND 0.00123f
C20368 VPWR.n440 VGND 0.00393f
C20369 VPWR.n441 VGND 0.00475f
C20370 VPWR.n442 VGND 0.00262f
C20371 VPWR.n443 VGND 0.00126f
C20372 VPWR.t2516 VGND 6.73e-19
C20373 VPWR.t2890 VGND 0.00127f
C20374 VPWR.n444 VGND 0.00204f
C20375 VPWR.n445 VGND 0.00462f
C20376 VPWR.n446 VGND 9.08e-19
C20377 VPWR.n447 VGND 0.0031f
C20378 VPWR.t2811 VGND 0.00239f
C20379 VPWR.n448 VGND 0.00608f
C20380 VPWR.n449 VGND 0.00513f
C20381 VPWR.n450 VGND 0.00387f
C20382 VPWR.n451 VGND 0.0136f
C20383 VPWR.t395 VGND 0.00463f
C20384 VPWR.n452 VGND 0.00578f
C20385 VPWR.n453 VGND 0.0185f
C20386 VPWR.n454 VGND 0.0179f
C20387 VPWR.t323 VGND 0.0046f
C20388 VPWR.n455 VGND 0.01f
C20389 VPWR.t3049 VGND 0.00633f
C20390 VPWR.n456 VGND 0.0121f
C20391 VPWR.n457 VGND 0.00352f
C20392 VPWR.t3370 VGND 0.0592f
C20393 VPWR.n458 VGND 0.0066f
C20394 VPWR.t3314 VGND 0.00102f
C20395 VPWR.t2793 VGND 0.00154f
C20396 VPWR.n459 VGND 0.00488f
C20397 VPWR.t3264 VGND 0.00136f
C20398 VPWR.t2334 VGND 0.00136f
C20399 VPWR.n460 VGND 0.00328f
C20400 VPWR.n461 VGND 0.0031f
C20401 VPWR.n462 VGND 0.00393f
C20402 VPWR.t1047 VGND 0.00102f
C20403 VPWR.t1770 VGND 0.00102f
C20404 VPWR.n463 VGND 0.00221f
C20405 VPWR.t465 VGND 0.00387f
C20406 VPWR.n464 VGND 0.00837f
C20407 VPWR.t3426 VGND 0.0289f
C20408 VPWR.t464 VGND 0.00387f
C20409 VPWR.n465 VGND 0.0604f
C20410 VPWR.n466 VGND 0.0146f
C20411 VPWR.n467 VGND 0.0117f
C20412 VPWR.t2839 VGND 6.73e-19
C20413 VPWR.t3287 VGND 9.96e-19
C20414 VPWR.n468 VGND 0.00177f
C20415 VPWR.n469 VGND 0.0149f
C20416 VPWR.t2782 VGND 0.00453f
C20417 VPWR.t136 VGND 0.0463f
C20418 VPWR.t1767 VGND 0.0111f
C20419 VPWR.t2771 VGND 0.0141f
C20420 VPWR.t1299 VGND 0.0141f
C20421 VPWR.t2769 VGND 0.0161f
C20422 VPWR.t3165 VGND 0.0211f
C20423 VPWR.t1628 VGND 0.0235f
C20424 VPWR.t2624 VGND 0.0321f
C20425 VPWR.t1301 VGND 0.0334f
C20426 VPWR.t606 VGND 0.0235f
C20427 VPWR.t3201 VGND 0.023f
C20428 VPWR.t2503 VGND 0.0493f
C20429 VPWR.t1616 VGND 0.0497f
C20430 VPWR.t1298 VGND 0.0215f
C20431 VPWR.t1811 VGND 0.0144f
C20432 VPWR.t2625 VGND 0.0148f
C20433 VPWR.t3217 VGND 0.0104f
C20434 VPWR.t2889 VGND 0.0154f
C20435 VPWR.t2515 VGND 0.0205f
C20436 VPWR.t2810 VGND 0.0502f
C20437 VPWR.t2891 VGND 0.0673f
C20438 VPWR.t394 VGND 0.042f
C20439 VPWR.t1197 VGND 0.027f
C20440 VPWR.t3167 VGND 0.0284f
C20441 VPWR.t3053 VGND 0.0242f
C20442 VPWR.n470 VGND 0.0344f
C20443 VPWR.t45 VGND 0.0775f
C20444 VPWR.t321 VGND 0.0287f
C20445 VPWR.t3048 VGND 0.0305f
C20446 VPWR.t1194 VGND 0.0171f
C20447 VPWR.t2948 VGND 0.0299f
C20448 VPWR.t3313 VGND 0.0284f
C20449 VPWR.t2333 VGND 0.0151f
C20450 VPWR.t3263 VGND 0.0109f
C20451 VPWR.t1769 VGND 0.0148f
C20452 VPWR.t1046 VGND 0.02f
C20453 VPWR.t2468 VGND 0.0544f
C20454 VPWR.t3161 VGND 0.018f
C20455 VPWR.t463 VGND 0.0166f
C20456 VPWR.t1048 VGND 0.0376f
C20457 VPWR.t3286 VGND 0.0398f
C20458 VPWR.t2838 VGND 0.0294f
C20459 VPWR.n471 VGND 0.0235f
C20460 VPWR.t711 VGND 0.0046f
C20461 VPWR.n472 VGND 0.00407f
C20462 VPWR.n473 VGND 0.00274f
C20463 VPWR.n474 VGND 6.26e-19
C20464 VPWR.n475 VGND 5.71e-19
C20465 VPWR.n476 VGND 3.29e-19
C20466 VPWR.n477 VGND 3.95e-19
C20467 VPWR.n478 VGND 4.17e-19
C20468 VPWR.n479 VGND 2.85e-19
C20469 VPWR.n480 VGND 6.54e-19
C20470 VPWR.n481 VGND 8.67e-19
C20471 VPWR.n482 VGND 0.1f
C20472 VPWR.n483 VGND 0.1f
C20473 VPWR.n484 VGND 0.00139f
C20474 VPWR.n485 VGND 9.06e-19
C20475 VPWR.t710 VGND 0.00463f
C20476 VPWR.n486 VGND 0.00578f
C20477 VPWR.t369 VGND 0.00463f
C20478 VPWR.t2549 VGND 0.00136f
C20479 VPWR.t2627 VGND 0.00136f
C20480 VPWR.n487 VGND 0.00317f
C20481 VPWR.n488 VGND 0.0185f
C20482 VPWR.n489 VGND 0.0179f
C20483 VPWR.t547 VGND 0.00387f
C20484 VPWR.n490 VGND 0.0107f
C20485 VPWR.n491 VGND 0.00796f
C20486 VPWR.t3453 VGND 0.0179f
C20487 VPWR.n492 VGND 0.00352f
C20488 VPWR.t2781 VGND 0.0126f
C20489 VPWR.t1045 VGND 0.0205f
C20490 VPWR.t3160 VGND 0.0285f
C20491 VPWR.t3077 VGND 0.0322f
C20492 VPWR.t2828 VGND 0.0322f
C20493 VPWR.t2911 VGND 0.0351f
C20494 VPWR.t709 VGND 0.0361f
C20495 VPWR.t3075 VGND 0.0493f
C20496 VPWR.t1383 VGND 0.0463f
C20497 VPWR.t1190 VGND 0.0171f
C20498 VPWR.t2626 VGND 0.0411f
C20499 VPWR.t2548 VGND 0.02f
C20500 VPWR.t367 VGND 0.0569f
C20501 VPWR.t545 VGND 0.0973f
C20502 VPWR.t294 VGND 0.0492f
C20503 VPWR.t905 VGND 0.0386f
C20504 VPWR.n493 VGND 0.0216f
C20505 VPWR.t459 VGND 0.00387f
C20506 VPWR.n494 VGND 0.00546f
C20507 VPWR.t3514 VGND 0.0289f
C20508 VPWR.t458 VGND 0.00387f
C20509 VPWR.n495 VGND 0.0604f
C20510 VPWR.n496 VGND 0.0146f
C20511 VPWR.t2340 VGND 0.00608f
C20512 VPWR.t2954 VGND 0.00231f
C20513 VPWR.n497 VGND 0.0138f
C20514 VPWR.n498 VGND 0.0117f
C20515 VPWR.n499 VGND 0.0099f
C20516 VPWR.t2538 VGND 0.00874f
C20517 VPWR.t2607 VGND 0.00265f
C20518 VPWR.n500 VGND 0.00606f
C20519 VPWR.n501 VGND 0.00138f
C20520 VPWR.n502 VGND 4.83e-19
C20521 VPWR.n503 VGND 2.85e-19
C20522 VPWR.n504 VGND 3.95e-19
C20523 VPWR.n505 VGND 6.54e-19
C20524 VPWR.n506 VGND 8.67e-19
C20525 VPWR.n507 VGND 3.95e-19
C20526 VPWR.n508 VGND 4.61e-19
C20527 VPWR.n509 VGND 2.41e-19
C20528 VPWR.n510 VGND 3.95e-19
C20529 VPWR.n511 VGND 3.07e-19
C20530 VPWR.n512 VGND 0.1f
C20531 VPWR.n513 VGND 0.0194f
C20532 VPWR.n515 VGND 8.67e-19
C20533 VPWR.n516 VGND 6.54e-19
C20534 VPWR.n517 VGND 9.06e-19
C20535 VPWR.n518 VGND 3.29e-19
C20536 VPWR.n519 VGND 5.71e-19
C20537 VPWR.n520 VGND 5.92e-19
C20538 VPWR.n521 VGND 5.05e-19
C20539 VPWR.t2149 VGND 0.00166f
C20540 VPWR.t2151 VGND 0.00166f
C20541 VPWR.n522 VGND 0.00359f
C20542 VPWR.n523 VGND 0.00606f
C20543 VPWR.n524 VGND 6.78e-19
C20544 VPWR.t2235 VGND 0.0016f
C20545 VPWR.t2241 VGND 0.0016f
C20546 VPWR.n525 VGND 0.00379f
C20547 VPWR.n526 VGND 0.00763f
C20548 VPWR.t2141 VGND 0.00166f
C20549 VPWR.t2147 VGND 0.00166f
C20550 VPWR.n527 VGND 0.00359f
C20551 VPWR.n528 VGND 0.00574f
C20552 VPWR.t2137 VGND 0.00166f
C20553 VPWR.t2139 VGND 0.00166f
C20554 VPWR.n529 VGND 0.00354f
C20555 VPWR.t3391 VGND 0.00911f
C20556 VPWR.t173 VGND 0.00391f
C20557 VPWR.n530 VGND 0.0253f
C20558 VPWR.t174 VGND 0.00391f
C20559 VPWR.n532 VGND 0.0138f
C20560 VPWR.n533 VGND 0.0128f
C20561 VPWR.t2643 VGND 0.00632f
C20562 VPWR.t2145 VGND 0.0016f
C20563 VPWR.t2155 VGND 0.00166f
C20564 VPWR.n534 VGND 0.00347f
C20565 VPWR.n535 VGND 0.00465f
C20566 VPWR.n536 VGND 0.00767f
C20567 VPWR.t2125 VGND 0.00166f
C20568 VPWR.t2153 VGND 0.00166f
C20569 VPWR.n537 VGND 0.00353f
C20570 VPWR.n538 VGND 0.00522f
C20571 VPWR.t2353 VGND 0.00632f
C20572 VPWR.t2133 VGND 0.00166f
C20573 VPWR.t2127 VGND 0.00166f
C20574 VPWR.n539 VGND 0.00353f
C20575 VPWR.n540 VGND 0.00522f
C20576 VPWR.t2600 VGND 0.00531f
C20577 VPWR.n541 VGND 0.00637f
C20578 VPWR.t2135 VGND 0.00166f
C20579 VPWR.t1064 VGND 0.00166f
C20580 VPWR.n542 VGND 0.0039f
C20581 VPWR.n543 VGND 0.00636f
C20582 VPWR.t1056 VGND 0.00166f
C20583 VPWR.t1058 VGND 0.00166f
C20584 VPWR.n544 VGND 0.00391f
C20585 VPWR.n545 VGND 0.00653f
C20586 VPWR.n546 VGND 0.00133f
C20587 VPWR.t1062 VGND 0.00614f
C20588 VPWR.t2325 VGND 0.0065f
C20589 VPWR.n547 VGND 0.00763f
C20590 VPWR.t494 VGND 0.00387f
C20591 VPWR.n548 VGND 0.00837f
C20592 VPWR.t2253 VGND 0.00653f
C20593 VPWR.n549 VGND 0.0108f
C20594 VPWR.n550 VGND 0.00393f
C20595 VPWR.t3511 VGND 0.0231f
C20596 VPWR.n551 VGND 0.0384f
C20597 VPWR.n552 VGND 0.00475f
C20598 VPWR.t493 VGND 0.00387f
C20599 VPWR.n553 VGND 0.00837f
C20600 VPWR.n554 VGND 0.00475f
C20601 VPWR.t2641 VGND 0.00527f
C20602 VPWR.t1533 VGND 0.00136f
C20603 VPWR.t1463 VGND 0.00136f
C20604 VPWR.n555 VGND 0.00328f
C20605 VPWR.t1461 VGND 0.0016f
C20606 VPWR.t2406 VGND 0.00208f
C20607 VPWR.n556 VGND 0.00422f
C20608 VPWR.t497 VGND 0.0046f
C20609 VPWR.n557 VGND 0.00644f
C20610 VPWR.t236 VGND 0.0046f
C20611 VPWR.n558 VGND 0.00407f
C20612 VPWR.t202 VGND 0.053f
C20613 VPWR.t1230 VGND 0.0493f
C20614 VPWR.t1232 VGND 0.02f
C20615 VPWR.t1234 VGND 0.0253f
C20616 VPWR.t3306 VGND 0.0144f
C20617 VPWR.t1228 VGND 0.0163f
C20618 VPWR.t948 VGND 0.0161f
C20619 VPWR.t1319 VGND 0.0121f
C20620 VPWR.t1896 VGND 0.0111f
C20621 VPWR.t1317 VGND 0.0196f
C20622 VPWR.t1315 VGND 0.0151f
C20623 VPWR.t1284 VGND 0.0371f
C20624 VPWR.t1518 VGND 0.0413f
C20625 VPWR.t982 VGND 0.027f
C20626 VPWR.t1286 VGND 0.0322f
C20627 VPWR.t1747 VGND 0.0285f
C20628 VPWR.t1325 VGND 0.0253f
C20629 VPWR.t715 VGND 0.0166f
C20630 VPWR.t2284 VGND 0.0388f
C20631 VPWR.t984 VGND 0.0493f
C20632 VPWR.t1183 VGND 0.0181f
C20633 VPWR.t1328 VGND 0.0383f
C20634 VPWR.t1748 VGND 0.0321f
C20635 VPWR.t747 VGND 0.0592f
C20636 VPWR.t234 VGND 0.0448f
C20637 VPWR.t1326 VGND 0.0151f
C20638 VPWR.t1022 VGND 0.025f
C20639 VPWR.t492 VGND 0.0311f
C20640 VPWR.t2867 VGND 0.025f
C20641 VPWR.t788 VGND 0.0453f
C20642 VPWR.t2640 VGND 0.0322f
C20643 VPWR.t1462 VGND 0.0158f
C20644 VPWR.t1532 VGND 0.02f
C20645 VPWR.t1460 VGND 0.0154f
C20646 VPWR.t3318 VGND 0.0228f
C20647 VPWR.t2601 VGND 0.0354f
C20648 VPWR.t318 VGND 0.0878f
C20649 VPWR.t495 VGND 0.0975f
C20650 VPWR.t42 VGND 0.0618f
C20651 VPWR.t1512 VGND 0.0257f
C20652 VPWR.t1405 VGND 0.0383f
C20653 VPWR.n559 VGND 0.0396f
C20654 VPWR.n560 VGND 0.00653f
C20655 VPWR.n561 VGND 0.00138f
C20656 VPWR.n562 VGND 4.83e-19
C20657 VPWR.n563 VGND 4.61e-19
C20658 VPWR.n564 VGND 6.54e-19
C20659 VPWR.n565 VGND 8.67e-19
C20660 VPWR.n566 VGND 4.39e-19
C20661 VPWR.n567 VGND 3.29e-19
C20662 VPWR.n568 VGND 5.27e-19
C20663 VPWR.n569 VGND 2.85e-19
C20664 VPWR.n570 VGND 2.85e-19
C20665 VPWR.n571 VGND 4.17e-19
C20666 VPWR.n572 VGND 5.71e-19
C20667 VPWR.n573 VGND 4.17e-19
C20668 VPWR.n574 VGND 3.51e-19
C20669 VPWR.n575 VGND 4.61e-19
C20670 VPWR.n576 VGND 4.17e-19
C20671 VPWR.n577 VGND 0.0057f
C20672 VPWR.n578 VGND 8.67e-19
C20673 VPWR.n579 VGND 6.54e-19
C20674 VPWR.n580 VGND 9.06e-19
C20675 VPWR.n581 VGND 0.00139f
C20676 VPWR.n582 VGND 5.27e-19
C20677 VPWR.n583 VGND 3.95e-19
C20678 VPWR.n584 VGND 5.05e-19
C20679 VPWR.n585 VGND 5.05e-19
C20680 VPWR.n586 VGND 2.63e-19
C20681 VPWR.t2216 VGND 0.00652f
C20682 VPWR.n587 VGND 0.00911f
C20683 VPWR.n588 VGND 1.99e-19
C20684 VPWR.n589 VGND 4.83e-19
C20685 VPWR.n590 VGND 4.61e-19
C20686 VPWR.n591 VGND 4.61e-19
C20687 VPWR.t1166 VGND 0.00633f
C20688 VPWR.t2998 VGND 0.0076f
C20689 VPWR.t1564 VGND 0.00166f
C20690 VPWR.t2986 VGND 0.00166f
C20691 VPWR.n592 VGND 0.00347f
C20692 VPWR.n593 VGND 0.0107f
C20693 VPWR.t1560 VGND 0.0016f
C20694 VPWR.n594 VGND 0.00706f
C20695 VPWR.n595 VGND 0.00211f
C20696 VPWR.t3381 VGND 0.00911f
C20697 VPWR.t317 VGND 0.00391f
C20698 VPWR.n596 VGND 0.0253f
C20699 VPWR.t316 VGND 0.00391f
C20700 VPWR.n598 VGND 0.0138f
C20701 VPWR.t2411 VGND 0.00102f
C20702 VPWR.t2308 VGND 0.00154f
C20703 VPWR.n599 VGND 0.00487f
C20704 VPWR.n600 VGND 0.0146f
C20705 VPWR.t2591 VGND 0.00622f
C20706 VPWR.n601 VGND 0.00123f
C20707 VPWR.t2119 VGND 0.00166f
C20708 VPWR.t2655 VGND 0.00219f
C20709 VPWR.n602 VGND 0.00445f
C20710 VPWR.t3488 VGND 0.00911f
C20711 VPWR.t624 VGND 0.00391f
C20712 VPWR.n603 VGND 0.0253f
C20713 VPWR.t623 VGND 0.00391f
C20714 VPWR.n605 VGND 0.0138f
C20715 VPWR.t3348 VGND 0.00911f
C20716 VPWR.t383 VGND 0.00391f
C20717 VPWR.n606 VGND 0.0253f
C20718 VPWR.t384 VGND 0.00391f
C20719 VPWR.n608 VGND 0.0138f
C20720 VPWR.n609 VGND 0.0112f
C20721 VPWR.n610 VGND 0.00345f
C20722 VPWR.n611 VGND 0.00177f
C20723 VPWR.t3083 VGND 0.0065f
C20724 VPWR.n612 VGND 0.0153f
C20725 VPWR.n613 VGND 0.00147f
C20726 VPWR.n614 VGND 0.00478f
C20727 VPWR.t2657 VGND 0.00529f
C20728 VPWR.n615 VGND 0.00518f
C20729 VPWR.t2984 VGND 0.00632f
C20730 VPWR.n616 VGND 0.00751f
C20731 VPWR.n617 VGND 8.07e-20
C20732 VPWR.n618 VGND 0.00393f
C20733 VPWR.n619 VGND 0.00444f
C20734 VPWR.n620 VGND 0.00179f
C20735 VPWR.n621 VGND 0.0067f
C20736 VPWR.n622 VGND 0.00143f
C20737 VPWR.n623 VGND 0.00262f
C20738 VPWR.n624 VGND 0.00179f
C20739 VPWR.n625 VGND 0.00339f
C20740 VPWR.t3085 VGND 0.00227f
C20741 VPWR.n626 VGND 0.00298f
C20742 VPWR.n627 VGND 0.00424f
C20743 VPWR.t1562 VGND 0.0016f
C20744 VPWR.n628 VGND 0.00706f
C20745 VPWR.n629 VGND 4.03e-19
C20746 VPWR.n630 VGND 0.00173f
C20747 VPWR.n631 VGND 6.86e-19
C20748 VPWR.n632 VGND 0.00475f
C20749 VPWR.n633 VGND 0.0015f
C20750 VPWR.n634 VGND 0.00524f
C20751 VPWR.n635 VGND 0.00148f
C20752 VPWR.n636 VGND 0.00524f
C20753 VPWR.n637 VGND 0.00393f
C20754 VPWR.n638 VGND 0.00199f
C20755 VPWR.n639 VGND 0.00139f
C20756 VPWR.n640 VGND 0.0107f
C20757 VPWR.t389 VGND 0.00387f
C20758 VPWR.n641 VGND 0.00493f
C20759 VPWR.n642 VGND 0.00213f
C20760 VPWR.n643 VGND 0.00393f
C20761 VPWR.t3406 VGND 0.0179f
C20762 VPWR.n644 VGND 0.0173f
C20763 VPWR.n645 VGND 0.00934f
C20764 VPWR.n646 VGND 0.0037f
C20765 VPWR.n647 VGND 9e-19
C20766 VPWR.n648 VGND 0.00138f
C20767 VPWR.n649 VGND 9.06e-19
C20768 VPWR.n650 VGND 5.48e-19
C20769 VPWR.n651 VGND 6.14e-19
C20770 VPWR.n652 VGND 0.00138f
C20771 VPWR.n653 VGND 8.88e-19
C20772 VPWR.n654 VGND 9.39e-19
C20773 VPWR.n655 VGND 0.00665f
C20774 VPWR.n656 VGND 0.00125f
C20775 VPWR.n657 VGND 4.27e-19
C20776 VPWR.n658 VGND 1.14e-19
C20777 VPWR.t2415 VGND 0.00632f
C20778 VPWR.n659 VGND 0.00785f
C20779 VPWR.n660 VGND 5.23e-19
C20780 VPWR.n661 VGND 0.00643f
C20781 VPWR.n662 VGND 4.27e-19
C20782 VPWR.n663 VGND 6.83e-19
C20783 VPWR.n664 VGND 3.7e-19
C20784 VPWR.n665 VGND 9.68e-19
C20785 VPWR.n666 VGND 9.96e-19
C20786 VPWR.n667 VGND 5.41e-19
C20787 VPWR.n668 VGND 4.39e-19
C20788 VPWR.n669 VGND 3.29e-19
C20789 VPWR.n670 VGND 5.27e-19
C20790 VPWR.n671 VGND 2.85e-19
C20791 VPWR.n672 VGND 2.85e-19
C20792 VPWR.n673 VGND 6.54e-19
C20793 VPWR.n674 VGND 8.67e-19
C20794 VPWR.n675 VGND 0.59f
C20795 VPWR.n676 VGND 0.071f
C20796 VPWR.n678 VGND 4.11e-19
C20797 VPWR.n679 VGND 4.11e-19
C20798 VPWR.n680 VGND 7.39e-19
C20799 VPWR.n681 VGND 5.19e-19
C20800 VPWR.n682 VGND 7.39e-19
C20801 VPWR.n683 VGND 4.11e-19
C20802 VPWR.n684 VGND 4.11e-19
C20803 VPWR.n685 VGND 4.17e-19
C20804 VPWR.n686 VGND 4.61e-19
C20805 VPWR.n687 VGND 3.51e-19
C20806 VPWR.n688 VGND 4.17e-19
C20807 VPWR.n689 VGND 4.17e-19
C20808 VPWR.n690 VGND 5.71e-19
C20809 VPWR.n691 VGND 7.4e-19
C20810 VPWR.t390 VGND 0.00387f
C20811 VPWR.n692 VGND 0.008f
C20812 VPWR.n693 VGND 0.00127f
C20813 VPWR.n694 VGND 4.48e-19
C20814 VPWR.n695 VGND 3.13e-19
C20815 VPWR.n696 VGND 2.56e-19
C20816 VPWR.n697 VGND 4.55e-19
C20817 VPWR.n698 VGND 0.00344f
C20818 VPWR.n699 VGND 2.56e-19
C20819 VPWR.n700 VGND 8.26e-19
C20820 VPWR.n701 VGND 4.83e-19
C20821 VPWR.n702 VGND 2.41e-19
C20822 VPWR.n703 VGND 3.73e-19
C20823 VPWR.n704 VGND 4.84e-19
C20824 VPWR.n705 VGND 6.83e-19
C20825 VPWR.n706 VGND 7.65e-19
C20826 VPWR.n707 VGND 2.92e-19
C20827 VPWR.n708 VGND 7.94e-19
C20828 VPWR.t2213 VGND 0.00659f
C20829 VPWR.n709 VGND 0.0102f
C20830 VPWR.t930 VGND 8.82e-19
C20831 VPWR.t3226 VGND 0.00144f
C20832 VPWR.n710 VGND 0.00533f
C20833 VPWR.n711 VGND 0.0069f
C20834 VPWR.t3230 VGND 0.00225f
C20835 VPWR.n712 VGND 0.00127f
C20836 VPWR.n713 VGND 0.00199f
C20837 VPWR.t382 VGND 0.046f
C20838 VPWR.t2118 VGND 0.0153f
C20839 VPWR.t2654 VGND 0.0201f
C20840 VPWR.t2656 VGND 0.053f
C20841 VPWR.t315 VGND 0.042f
C20842 VPWR.t2307 VGND 0.0183f
C20843 VPWR.t2410 VGND 0.0131f
C20844 VPWR.t2214 VGND 0.0144f
C20845 VPWR.t2590 VGND 0.0154f
C20846 VPWR.t1559 VGND 0.0154f
C20847 VPWR.t3084 VGND 0.0193f
C20848 VPWR.t1561 VGND 0.0262f
C20849 VPWR.t2592 VGND 0.0176f
C20850 VPWR.t2726 VGND 0.0161f
C20851 VPWR.t2997 VGND 0.0141f
C20852 VPWR.t1563 VGND 0.018f
C20853 VPWR.t2985 VGND 0.0258f
C20854 VPWR.t1165 VGND 0.0361f
C20855 VPWR.t388 VGND 0.0316f
C20856 VPWR.t2414 VGND 0.026f
C20857 VPWR.t2215 VGND 0.0156f
C20858 VPWR.t929 VGND 0.0205f
C20859 VPWR.t2212 VGND 0.0151f
C20860 VPWR.t2095 VGND 0.0129f
C20861 VPWR.t3225 VGND 0.0208f
C20862 VPWR.t1655 VGND 0.0316f
C20863 VPWR.t3227 VGND 0.0129f
C20864 VPWR.t3170 VGND 0.0161f
C20865 VPWR.t1695 VGND 0.03f
C20866 VPWR.t838 VGND 0.0269f
C20867 VPWR.t3229 VGND 0.0126f
C20868 VPWR.n714 VGND 0.00874f
C20869 VPWR.t3157 VGND 0.00614f
C20870 VPWR.n715 VGND 0.00827f
C20871 VPWR.n716 VGND 0.00901f
C20872 VPWR.t761 VGND 0.00661f
C20873 VPWR.n717 VGND 0.0167f
C20874 VPWR.t2920 VGND 0.0016f
C20875 VPWR.t2431 VGND 0.00208f
C20876 VPWR.n718 VGND 0.00422f
C20877 VPWR.n719 VGND 0.00606f
C20878 VPWR.t1086 VGND 0.00561f
C20879 VPWR.t2874 VGND 0.00102f
C20880 VPWR.t1778 VGND 0.00102f
C20881 VPWR.n720 VGND 0.00221f
C20882 VPWR.n721 VGND 0.00569f
C20883 VPWR.n722 VGND 0.0072f
C20884 VPWR.t1539 VGND 0.00692f
C20885 VPWR.t1074 VGND 0.00614f
C20886 VPWR.t2722 VGND 0.00136f
C20887 VPWR.t2033 VGND 0.00136f
C20888 VPWR.n723 VGND 0.00317f
C20889 VPWR.t3390 VGND 0.0179f
C20890 VPWR.n724 VGND 0.0173f
C20891 VPWR.t510 VGND 0.00387f
C20892 VPWR.n725 VGND 0.00493f
C20893 VPWR.t759 VGND -2.18e-20
C20894 VPWR.t2526 VGND 0.00137f
C20895 VPWR.n726 VGND 0.00618f
C20896 VPWR.t3505 VGND 0.0179f
C20897 VPWR.t3336 VGND 0.00911f
C20898 VPWR.t186 VGND 0.00391f
C20899 VPWR.n727 VGND 0.0253f
C20900 VPWR.t185 VGND 0.00391f
C20901 VPWR.n729 VGND 0.0138f
C20902 VPWR.t3317 VGND 0.0016f
C20903 VPWR.t2388 VGND 0.0016f
C20904 VPWR.n730 VGND 0.00371f
C20905 VPWR.n731 VGND 0.0144f
C20906 VPWR.t2639 VGND 0.0016f
C20907 VPWR.t2631 VGND 0.0016f
C20908 VPWR.n732 VGND 0.00379f
C20909 VPWR.n733 VGND 6.55e-19
C20910 VPWR.n734 VGND 4.58e-19
C20911 VPWR.n735 VGND 6.26e-19
C20912 VPWR.n736 VGND 5.12e-19
C20913 VPWR.n737 VGND 0.00108f
C20914 VPWR.n738 VGND 0.00122f
C20915 VPWR.n739 VGND 3.95e-19
C20916 VPWR.n740 VGND 3.95e-19
C20917 VPWR.n741 VGND 7.68e-19
C20918 VPWR.n742 VGND 5.05e-19
C20919 VPWR.n743 VGND 8.67e-19
C20920 VPWR.n744 VGND 6.54e-19
C20921 VPWR.n745 VGND 9.06e-19
C20922 VPWR.n747 VGND 0.1f
C20923 VPWR.n748 VGND 0.00139f
C20924 VPWR.n749 VGND 9.06e-19
C20925 VPWR.t1125 VGND 0.00631f
C20926 VPWR.t2084 VGND 0.00234f
C20927 VPWR.t3496 VGND 0.0179f
C20928 VPWR.n750 VGND 0.0173f
C20929 VPWR.n751 VGND 0.0103f
C20930 VPWR.n752 VGND 0.0133f
C20931 VPWR.t654 VGND 0.00387f
C20932 VPWR.n753 VGND 0.00837f
C20933 VPWR.n754 VGND 0.00525f
C20934 VPWR.t1580 VGND 0.00166f
C20935 VPWR.t1582 VGND 0.00166f
C20936 VPWR.n755 VGND 0.00353f
C20937 VPWR.t3033 VGND 0.00632f
C20938 VPWR.t919 VGND 0.00652f
C20939 VPWR.n756 VGND 0.00108f
C20940 VPWR.t1584 VGND 0.00166f
C20941 VPWR.t1586 VGND 0.00166f
C20942 VPWR.n757 VGND 0.00359f
C20943 VPWR.n758 VGND 0.00546f
C20944 VPWR.t1605 VGND 0.0016f
C20945 VPWR.t1589 VGND 0.00166f
C20946 VPWR.n759 VGND 0.00347f
C20947 VPWR.n760 VGND 0.0105f
C20948 VPWR.t476 VGND 0.00387f
C20949 VPWR.n761 VGND 0.0033f
C20950 VPWR.n762 VGND 0.00202f
C20951 VPWR.t1601 VGND 0.00166f
C20952 VPWR.t1593 VGND 0.00166f
C20953 VPWR.n763 VGND 0.00359f
C20954 VPWR.n764 VGND 0.00643f
C20955 VPWR.t737 VGND 0.00387f
C20956 VPWR.n765 VGND 0.00755f
C20957 VPWR.n766 VGND 5.69e-19
C20958 VPWR.n767 VGND 3.29e-19
C20959 VPWR.n768 VGND 5.71e-19
C20960 VPWR.n769 VGND 5.92e-19
C20961 VPWR.n770 VGND 5.05e-19
C20962 VPWR.n771 VGND 8.67e-19
C20963 VPWR.n772 VGND 6.54e-19
C20964 VPWR.n773 VGND 9.06e-19
C20965 VPWR.n774 VGND 0.1f
C20966 VPWR.n775 VGND 0.00139f
C20967 VPWR.n776 VGND 9.06e-19
C20968 VPWR.n777 VGND 8.11e-19
C20969 VPWR.n778 VGND 3.95e-19
C20970 VPWR.n779 VGND 1.76e-19
C20971 VPWR.n780 VGND 3.95e-19
C20972 VPWR.n781 VGND 7.68e-19
C20973 VPWR.n782 VGND 5.05e-19
C20974 VPWR.n783 VGND 1.76e-19
C20975 VPWR.n784 VGND 5.48e-19
C20976 VPWR.n786 VGND 0.0976f
C20977 VPWR.n787 VGND 0.071f
C20978 VPWR.n788 VGND 6.54e-19
C20979 VPWR.n789 VGND 8.67e-19
C20980 VPWR.n790 VGND 3.95e-19
C20981 VPWR.n791 VGND 4.61e-19
C20982 VPWR.n792 VGND 2.41e-19
C20983 VPWR.n793 VGND 3.95e-19
C20984 VPWR.n794 VGND 3.07e-19
C20985 VPWR.n795 VGND 4.83e-19
C20986 VPWR.n796 VGND 2.85e-19
C20987 VPWR.n797 VGND 3.95e-19
C20988 VPWR.n798 VGND 3.95e-19
C20989 VPWR.t3479 VGND 0.0231f
C20990 VPWR.t3068 VGND 0.00676f
C20991 VPWR.n799 VGND 0.00956f
C20992 VPWR.n800 VGND 0.00168f
C20993 VPWR.t3361 VGND 0.00911f
C20994 VPWR.t251 VGND 0.00391f
C20995 VPWR.n801 VGND 0.0253f
C20996 VPWR.t250 VGND 0.00391f
C20997 VPWR.n803 VGND 0.0138f
C20998 VPWR.t1312 VGND 0.00239f
C20999 VPWR.t3066 VGND 0.00127f
C21000 VPWR.t1694 VGND 6.73e-19
C21001 VPWR.n804 VGND 0.00204f
C21002 VPWR.n805 VGND 0.00705f
C21003 VPWR.n806 VGND 0.00782f
C21004 VPWR.t763 VGND 0.00453f
C21005 VPWR.t1941 VGND 9.96e-19
C21006 VPWR.t1700 VGND 6.73e-19
C21007 VPWR.n807 VGND 0.00176f
C21008 VPWR.n808 VGND 0.0102f
C21009 VPWR.n809 VGND 0.0101f
C21010 VPWR.n810 VGND 0.0115f
C21011 VPWR.n811 VGND 0.0111f
C21012 VPWR.t159 VGND 0.00387f
C21013 VPWR.n812 VGND 0.00374f
C21014 VPWR.t3583 VGND 0.0289f
C21015 VPWR.t158 VGND 0.00387f
C21016 VPWR.n813 VGND 0.0604f
C21017 VPWR.n814 VGND 0.0146f
C21018 VPWR.n815 VGND 0.0117f
C21019 VPWR.t2255 VGND 0.00235f
C21020 VPWR.n816 VGND 0.0148f
C21021 VPWR.t1909 VGND 0.00102f
C21022 VPWR.t1516 VGND 0.00102f
C21023 VPWR.n817 VGND 0.00217f
C21024 VPWR.n818 VGND 0.00284f
C21025 VPWR.t2398 VGND 6.73e-19
C21026 VPWR.t2396 VGND 6.73e-19
C21027 VPWR.n819 VGND 0.00141f
C21028 VPWR.t1698 VGND 9.71e-19
C21029 VPWR.t1170 VGND 9.22e-19
C21030 VPWR.n820 VGND 0.00196f
C21031 VPWR.n821 VGND 0.00797f
C21032 VPWR.t3417 VGND 0.0289f
C21033 VPWR.t595 VGND 0.00387f
C21034 VPWR.n822 VGND 0.0604f
C21035 VPWR.n823 VGND 0.0146f
C21036 VPWR.n824 VGND 0.0117f
C21037 VPWR.n825 VGND 0.00996f
C21038 VPWR.n826 VGND 0.00199f
C21039 VPWR.n827 VGND 0.00903f
C21040 VPWR.n828 VGND 0.0113f
C21041 VPWR.n829 VGND 0.0104f
C21042 VPWR.n830 VGND 0.0138f
C21043 VPWR.n831 VGND 0.00524f
C21044 VPWR.n832 VGND 0.0133f
C21045 VPWR.n833 VGND 0.00524f
C21046 VPWR.t835 VGND 0.00461f
C21047 VPWR.n834 VGND 0.00352f
C21048 VPWR.t596 VGND 0.00387f
C21049 VPWR.n835 VGND 0.00815f
C21050 VPWR.n836 VGND 0.0014f
C21051 VPWR.n837 VGND 0.00239f
C21052 VPWR.n838 VGND 0.0031f
C21053 VPWR.n839 VGND 0.00179f
C21054 VPWR.n840 VGND 0.00152f
C21055 VPWR.n841 VGND 0.00472f
C21056 VPWR.t1939 VGND 0.00102f
C21057 VPWR.t1911 VGND 0.00102f
C21058 VPWR.n842 VGND 0.00217f
C21059 VPWR.n843 VGND 0.00472f
C21060 VPWR.n844 VGND 4.03e-20
C21061 VPWR.n845 VGND 0.00475f
C21062 VPWR.n846 VGND 0.00184f
C21063 VPWR.n847 VGND 0.0031f
C21064 VPWR.n848 VGND 0.00141f
C21065 VPWR.n849 VGND 0.00199f
C21066 VPWR.n850 VGND 0.00901f
C21067 VPWR.n851 VGND 0.00807f
C21068 VPWR.n852 VGND 0.0104f
C21069 VPWR.n853 VGND 0.00524f
C21070 VPWR.n854 VGND 0.00524f
C21071 VPWR.n855 VGND 0.0031f
C21072 VPWR.n856 VGND 0.00487f
C21073 VPWR.t2605 VGND 0.00652f
C21074 VPWR.n857 VGND 0.00903f
C21075 VPWR.n858 VGND 0.00393f
C21076 VPWR.n859 VGND 0.00135f
C21077 VPWR.n860 VGND 0.00524f
C21078 VPWR.t2173 VGND 0.00652f
C21079 VPWR.n861 VGND 0.00925f
C21080 VPWR.n862 VGND 0.00313f
C21081 VPWR.n863 VGND 0.00444f
C21082 VPWR.n864 VGND 0.00199f
C21083 VPWR.n865 VGND 0.00262f
C21084 VPWR.n866 VGND 0.00202f
C21085 VPWR.n867 VGND 0.00525f
C21086 VPWR.t736 VGND 0.00387f
C21087 VPWR.n868 VGND 0.00837f
C21088 VPWR.n869 VGND 0.00688f
C21089 VPWR.n870 VGND 0.0376f
C21090 VPWR.n871 VGND 0.00364f
C21091 VPWR.n872 VGND 0.00259f
C21092 VPWR.n873 VGND 2.85e-19
C21093 VPWR.n874 VGND 2.28e-19
C21094 VPWR.n875 VGND 6.26e-19
C21095 VPWR.n876 VGND 5.12e-19
C21096 VPWR.n877 VGND 3.13e-19
C21097 VPWR.n878 VGND 0.00122f
C21098 VPWR.n879 VGND 0.00108f
C21099 VPWR.n880 VGND 5.12e-19
C21100 VPWR.n881 VGND 5.98e-19
C21101 VPWR.t922 VGND 0.00184f
C21102 VPWR.t2547 VGND 0.00166f
C21103 VPWR.n882 VGND 0.00358f
C21104 VPWR.n883 VGND 9.71e-19
C21105 VPWR.n884 VGND 0.00248f
C21106 VPWR.n885 VGND 0.00665f
C21107 VPWR.n886 VGND 9.71e-19
C21108 VPWR.n887 VGND 8.97e-19
C21109 VPWR.n888 VGND 0.00673f
C21110 VPWR.n889 VGND 0.0123f
C21111 VPWR.n890 VGND 3.13e-19
C21112 VPWR.n891 VGND 5.41e-19
C21113 VPWR.n892 VGND 9.68e-19
C21114 VPWR.n893 VGND 9.96e-19
C21115 VPWR.n894 VGND 5.41e-19
C21116 VPWR.n895 VGND 1.76e-19
C21117 VPWR.n896 VGND 4.39e-19
C21118 VPWR.n897 VGND 6.14e-19
C21119 VPWR.n898 VGND 4.17e-19
C21120 VPWR.n899 VGND 5.05e-19
C21121 VPWR.n900 VGND 6.55e-19
C21122 VPWR.n901 VGND 6.26e-19
C21123 VPWR.n902 VGND 3.7e-19
C21124 VPWR.n903 VGND 3.42e-19
C21125 VPWR.n904 VGND 3.7e-19
C21126 VPWR.n905 VGND 4.84e-19
C21127 VPWR.n906 VGND 0.00128f
C21128 VPWR.n907 VGND 2.56e-19
C21129 VPWR.n908 VGND 4.27e-19
C21130 VPWR.n909 VGND 5.12e-19
C21131 VPWR.n910 VGND 3.7e-19
C21132 VPWR.n911 VGND 4.17e-19
C21133 VPWR.n912 VGND 2.85e-19
C21134 VPWR.n913 VGND 2.85e-19
C21135 VPWR.n914 VGND 4.11e-19
C21136 VPWR.n915 VGND 4.11e-19
C21137 VPWR.n916 VGND 7.39e-19
C21138 VPWR.n917 VGND 5.19e-19
C21139 VPWR.n918 VGND 7.39e-19
C21140 VPWR.n919 VGND 4.11e-19
C21141 VPWR.n920 VGND 4.11e-19
C21142 VPWR.n922 VGND 0.0057f
C21143 VPWR.n923 VGND 0.00138f
C21144 VPWR.n924 VGND 5.48e-19
C21145 VPWR.n925 VGND 4.17e-19
C21146 VPWR.n926 VGND 1.33e-19
C21147 VPWR.n927 VGND 6.58e-20
C21148 VPWR.n928 VGND 0.00118f
C21149 VPWR.n929 VGND 8.05e-19
C21150 VPWR.n930 VGND 4.84e-19
C21151 VPWR.n931 VGND 8.54e-20
C21152 VPWR.n932 VGND 0.00595f
C21153 VPWR.t1633 VGND 6.73e-19
C21154 VPWR.t2540 VGND 6.73e-19
C21155 VPWR.n933 VGND 0.00166f
C21156 VPWR.n934 VGND 0.0104f
C21157 VPWR.t1603 VGND 0.00556f
C21158 VPWR.n935 VGND 0.00642f
C21159 VPWR.n936 VGND 0.00105f
C21160 VPWR.n937 VGND 0.00393f
C21161 VPWR.n938 VGND 0.0015f
C21162 VPWR.n939 VGND 0.00524f
C21163 VPWR.t1576 VGND 0.00166f
C21164 VPWR.t1599 VGND 0.00166f
C21165 VPWR.n940 VGND 0.00359f
C21166 VPWR.n941 VGND 0.00523f
C21167 VPWR.t924 VGND 9.96e-19
C21168 VPWR.t1039 VGND -0.00105f
C21169 VPWR.n942 VGND 0.00655f
C21170 VPWR.n943 VGND 0.00489f
C21171 VPWR.n944 VGND 0.00524f
C21172 VPWR.n945 VGND 0.00393f
C21173 VPWR.n946 VGND 0.00128f
C21174 VPWR.n947 VGND 0.00628f
C21175 VPWR.t475 VGND 0.00387f
C21176 VPWR.t3440 VGND 0.0179f
C21177 VPWR.t1597 VGND 0.00166f
C21178 VPWR.t1578 VGND 0.00166f
C21179 VPWR.n948 VGND 0.00353f
C21180 VPWR.n949 VGND 0.012f
C21181 VPWR.n950 VGND 0.0078f
C21182 VPWR.n951 VGND 0.00746f
C21183 VPWR.n952 VGND 0.0165f
C21184 VPWR.n953 VGND 0.00495f
C21185 VPWR.n954 VGND 0.00496f
C21186 VPWR.n955 VGND 0.00393f
C21187 VPWR.n956 VGND 0.00524f
C21188 VPWR.n957 VGND 0.00524f
C21189 VPWR.n958 VGND 0.0031f
C21190 VPWR.n959 VGND 0.00489f
C21191 VPWR.n960 VGND 0.00121f
C21192 VPWR.n961 VGND 0.00722f
C21193 VPWR.n962 VGND 0.00393f
C21194 VPWR.n963 VGND 0.00524f
C21195 VPWR.n964 VGND 0.00313f
C21196 VPWR.n965 VGND 9.64e-19
C21197 VPWR.n966 VGND 0.00785f
C21198 VPWR.n967 VGND 0.00521f
C21199 VPWR.n968 VGND 0.00143f
C21200 VPWR.n969 VGND 0.00393f
C21201 VPWR.t1855 VGND 0.00676f
C21202 VPWR.n970 VGND 0.00959f
C21203 VPWR.t1595 VGND 0.00166f
C21204 VPWR.t1588 VGND 0.00166f
C21205 VPWR.n971 VGND 0.00353f
C21206 VPWR.n972 VGND 0.00522f
C21207 VPWR.n973 VGND 3.53e-19
C21208 VPWR.n974 VGND 0.00524f
C21209 VPWR.t1794 VGND 0.00242f
C21210 VPWR.n975 VGND 0.0048f
C21211 VPWR.n976 VGND 6.64e-19
C21212 VPWR.n977 VGND 0.00524f
C21213 VPWR.t1591 VGND 0.00166f
C21214 VPWR.t3155 VGND 0.00166f
C21215 VPWR.n978 VGND 0.00389f
C21216 VPWR.n979 VGND 0.00504f
C21217 VPWR.n980 VGND 9.03e-19
C21218 VPWR.n981 VGND 0.00524f
C21219 VPWR.t1372 VGND 6.73e-19
C21220 VPWR.t1853 VGND 0.00127f
C21221 VPWR.n982 VGND 0.00207f
C21222 VPWR.n983 VGND 0.00431f
C21223 VPWR.n984 VGND 0.00524f
C21224 VPWR.t3153 VGND 0.00166f
C21225 VPWR.t3151 VGND 0.00166f
C21226 VPWR.n985 VGND 0.00391f
C21227 VPWR.n986 VGND 0.00641f
C21228 VPWR.n987 VGND 0.00524f
C21229 VPWR.n988 VGND 0.00121f
C21230 VPWR.n989 VGND 0.00524f
C21231 VPWR.n990 VGND 0.0031f
C21232 VPWR.n991 VGND 0.00199f
C21233 VPWR.t1253 VGND 0.00453f
C21234 VPWR.n992 VGND 0.00562f
C21235 VPWR.n993 VGND 0.00151f
C21236 VPWR.n994 VGND 0.00393f
C21237 VPWR.t1969 VGND 0.00676f
C21238 VPWR.n995 VGND 0.00956f
C21239 VPWR.t1370 VGND 6.73e-19
C21240 VPWR.t3283 VGND 9.96e-19
C21241 VPWR.n996 VGND 0.00176f
C21242 VPWR.n997 VGND 0.00421f
C21243 VPWR.n998 VGND 4.74e-19
C21244 VPWR.n999 VGND 0.00524f
C21245 VPWR.t3285 VGND 0.00242f
C21246 VPWR.n1000 VGND 0.00484f
C21247 VPWR.n1001 VGND 5.14e-19
C21248 VPWR.n1002 VGND 0.00524f
C21249 VPWR.n1003 VGND 0.00105f
C21250 VPWR.n1004 VGND 0.00524f
C21251 VPWR.t2837 VGND 6.73e-19
C21252 VPWR.t1967 VGND 0.00127f
C21253 VPWR.n1005 VGND 0.00207f
C21254 VPWR.n1006 VGND 0.00496f
C21255 VPWR.n1007 VGND 0.00524f
C21256 VPWR.n1008 VGND 0.00141f
C21257 VPWR.n1009 VGND 0.00524f
C21258 VPWR.t1727 VGND 0.00238f
C21259 VPWR.n1010 VGND 0.0053f
C21260 VPWR.n1011 VGND 0.00524f
C21261 VPWR.n1012 VGND 0.00141f
C21262 VPWR.n1013 VGND 0.00524f
C21263 VPWR.t2370 VGND 0.00453f
C21264 VPWR.n1014 VGND 0.00562f
C21265 VPWR.n1015 VGND 0.00123f
C21266 VPWR.n1016 VGND 0.00524f
C21267 VPWR.t791 VGND 0.00102f
C21268 VPWR.t1838 VGND 0.00102f
C21269 VPWR.n1017 VGND 0.00217f
C21270 VPWR.n1018 VGND 0.00472f
C21271 VPWR.n1019 VGND 6.45e-19
C21272 VPWR.n1020 VGND 0.00524f
C21273 VPWR.n1021 VGND 0.0031f
C21274 VPWR.n1022 VGND 0.00106f
C21275 VPWR.t2841 VGND 6.73e-19
C21276 VPWR.t2312 VGND 9.96e-19
C21277 VPWR.n1023 VGND 0.00178f
C21278 VPWR.n1024 VGND 0.00661f
C21279 VPWR.t653 VGND 0.00387f
C21280 VPWR.n1025 VGND 0.00493f
C21281 VPWR.n1026 VGND 0.00254f
C21282 VPWR.n1027 VGND 0.00393f
C21283 VPWR.n1028 VGND 0.00524f
C21284 VPWR.n1029 VGND 0.00524f
C21285 VPWR.n1030 VGND 0.0031f
C21286 VPWR.n1031 VGND 0.00182f
C21287 VPWR.n1032 VGND 9.91e-19
C21288 VPWR.n1033 VGND 0.00356f
C21289 VPWR.n1034 VGND 0.00523f
C21290 VPWR.n1035 VGND 0.00127f
C21291 VPWR.n1036 VGND 0.00473f
C21292 VPWR.n1037 VGND 0.00142f
C21293 VPWR.n1038 VGND 0.00504f
C21294 VPWR.t2637 VGND 0.0016f
C21295 VPWR.t2633 VGND 0.0016f
C21296 VPWR.n1039 VGND 0.00379f
C21297 VPWR.n1040 VGND 8.37e-19
C21298 VPWR.n1041 VGND 0.00737f
C21299 VPWR.n1042 VGND 3.13e-19
C21300 VPWR.n1043 VGND 5.71e-19
C21301 VPWR.n1044 VGND 3.29e-19
C21302 VPWR.n1045 VGND 3.95e-19
C21303 VPWR.n1046 VGND 4.17e-19
C21304 VPWR.n1047 VGND 2.85e-19
C21305 VPWR.n1048 VGND 6.54e-19
C21306 VPWR.n1049 VGND 8.67e-19
C21307 VPWR.n1050 VGND 7.97e-19
C21308 VPWR.n1051 VGND 6.14e-19
C21309 VPWR.n1052 VGND 4.39e-19
C21310 VPWR.n1053 VGND 1.76e-19
C21311 VPWR.n1054 VGND 4.83e-19
C21312 VPWR.n1055 VGND 2.41e-19
C21313 VPWR.n1056 VGND 9.68e-19
C21314 VPWR.n1057 VGND 0.00103f
C21315 VPWR.n1058 VGND 3.13e-19
C21316 VPWR.n1059 VGND 5.12e-19
C21317 VPWR.n1060 VGND 3.73e-19
C21318 VPWR.n1061 VGND 3.07e-19
C21319 VPWR.n1062 VGND 4.11e-19
C21320 VPWR.n1063 VGND 4.11e-19
C21321 VPWR.n1064 VGND 7.39e-19
C21322 VPWR.n1065 VGND 5.19e-19
C21323 VPWR.n1066 VGND 7.39e-19
C21324 VPWR.n1067 VGND 4.11e-19
C21325 VPWR.n1068 VGND 4.11e-19
C21326 VPWR.n1069 VGND 2.85e-19
C21327 VPWR.n1070 VGND 3.95e-19
C21328 VPWR.n1071 VGND 2.85e-19
C21329 VPWR.n1072 VGND 4.83e-19
C21330 VPWR.n1073 VGND 4.17e-19
C21331 VPWR.n1074 VGND 5.05e-19
C21332 VPWR.n1075 VGND 6.26e-19
C21333 VPWR.n1076 VGND 1.14e-19
C21334 VPWR.n1077 VGND 4.29e-19
C21335 VPWR.n1078 VGND 4.54e-19
C21336 VPWR.n1079 VGND 7.4e-19
C21337 VPWR.n1080 VGND 5.41e-19
C21338 VPWR.n1081 VGND 5.12e-19
C21339 VPWR.n1082 VGND 4.27e-19
C21340 VPWR.n1083 VGND 9.96e-19
C21341 VPWR.n1084 VGND 0.00131f
C21342 VPWR.n1085 VGND 5.98e-19
C21343 VPWR.t1127 VGND 0.0016f
C21344 VPWR.t2629 VGND 0.0016f
C21345 VPWR.n1086 VGND 0.00365f
C21346 VPWR.n1087 VGND 0.00503f
C21347 VPWR.t1035 VGND 0.00102f
C21348 VPWR.t1780 VGND 0.00102f
C21349 VPWR.n1088 VGND 0.00217f
C21350 VPWR.n1089 VGND 0.00462f
C21351 VPWR.n1090 VGND 4.54e-19
C21352 VPWR.n1091 VGND 6.99e-19
C21353 VPWR.n1092 VGND 0.00218f
C21354 VPWR.n1093 VGND 0.00137f
C21355 VPWR.n1094 VGND 5.92e-19
C21356 VPWR.n1095 VGND 5.05e-19
C21357 VPWR.n1096 VGND 4.17e-19
C21358 VPWR.n1097 VGND 5.48e-19
C21359 VPWR.n1099 VGND 0.0057f
C21360 VPWR.n1100 VGND 0.00138f
C21361 VPWR.n1101 VGND 5.48e-19
C21362 VPWR.n1102 VGND 1.76e-19
C21363 VPWR.n1103 VGND 8.11e-19
C21364 VPWR.n1104 VGND 3.95e-19
C21365 VPWR.n1105 VGND 1.77e-19
C21366 VPWR.n1106 VGND 3.13e-19
C21367 VPWR.n1107 VGND 5.12e-19
C21368 VPWR.n1108 VGND 5.98e-19
C21369 VPWR.n1109 VGND 8.39e-20
C21370 VPWR.n1110 VGND 0.00819f
C21371 VPWR.n1111 VGND 0.00103f
C21372 VPWR.n1112 VGND 0.00393f
C21373 VPWR.t2635 VGND 0.00655f
C21374 VPWR.n1113 VGND 0.0108f
C21375 VPWR.n1114 VGND 0.00393f
C21376 VPWR.n1115 VGND 0.0044f
C21377 VPWR.n1116 VGND 0.00199f
C21378 VPWR.n1117 VGND 0.0031f
C21379 VPWR.n1118 VGND 0.00524f
C21380 VPWR.n1119 VGND 0.00393f
C21381 VPWR.n1120 VGND 0.00487f
C21382 VPWR.t678 VGND 0.00387f
C21383 VPWR.n1121 VGND 0.00493f
C21384 VPWR.n1122 VGND 0.0168f
C21385 VPWR.n1123 VGND 0.00894f
C21386 VPWR.n1124 VGND 0.0074f
C21387 VPWR.n1125 VGND 0.0126f
C21388 VPWR.t679 VGND 0.00399f
C21389 VPWR.n1126 VGND 0.0129f
C21390 VPWR.n1127 VGND 0.00443f
C21391 VPWR.n1128 VGND 0.00179f
C21392 VPWR.n1129 VGND 0.00179f
C21393 VPWR.n1130 VGND 0.0103f
C21394 VPWR.t511 VGND 0.00387f
C21395 VPWR.n1131 VGND 0.0049f
C21396 VPWR.n1132 VGND 0.00837f
C21397 VPWR.n1133 VGND 0.0188f
C21398 VPWR.n1134 VGND 0.00475f
C21399 VPWR.n1135 VGND 0.0031f
C21400 VPWR.n1136 VGND 0.00179f
C21401 VPWR.n1137 VGND 0.00787f
C21402 VPWR.n1138 VGND 0.0106f
C21403 VPWR.n1139 VGND 0.00475f
C21404 VPWR.t1052 VGND 0.00166f
C21405 VPWR.t1054 VGND 0.00166f
C21406 VPWR.n1140 VGND 0.00379f
C21407 VPWR.n1141 VGND 0.0052f
C21408 VPWR.t3262 VGND 0.00239f
C21409 VPWR.n1142 VGND 0.00421f
C21410 VPWR.n1143 VGND 4.13e-19
C21411 VPWR.n1144 VGND 0.00524f
C21412 VPWR.n1145 VGND 0.00132f
C21413 VPWR.n1146 VGND 0.00524f
C21414 VPWR.t1050 VGND 0.00166f
C21415 VPWR.t1084 VGND 0.00166f
C21416 VPWR.n1147 VGND 0.00377f
C21417 VPWR.n1148 VGND 0.0054f
C21418 VPWR.t1380 VGND 6.73e-19
C21419 VPWR.t1541 VGND 0.00127f
C21420 VPWR.n1149 VGND 0.00203f
C21421 VPWR.n1150 VGND 0.00359f
C21422 VPWR.n1151 VGND 3.21e-19
C21423 VPWR.n1152 VGND 0.00524f
C21424 VPWR.n1153 VGND 0.00119f
C21425 VPWR.n1154 VGND 0.00524f
C21426 VPWR.t1110 VGND 0.00166f
C21427 VPWR.t1088 VGND 0.00166f
C21428 VPWR.n1155 VGND 0.00359f
C21429 VPWR.n1156 VGND 0.0057f
C21430 VPWR.n1157 VGND 9.96e-19
C21431 VPWR.n1158 VGND 0.00524f
C21432 VPWR.n1159 VGND 0.0012f
C21433 VPWR.n1160 VGND 0.00524f
C21434 VPWR.t1509 VGND 0.00455f
C21435 VPWR.t1092 VGND 0.00166f
C21436 VPWR.t1096 VGND 0.00166f
C21437 VPWR.n1161 VGND 0.00359f
C21438 VPWR.n1162 VGND 0.00562f
C21439 VPWR.n1163 VGND 0.00655f
C21440 VPWR.n1164 VGND 0.00524f
C21441 VPWR.t1098 VGND 0.00166f
C21442 VPWR.t1090 VGND 0.00166f
C21443 VPWR.n1165 VGND 0.00359f
C21444 VPWR.n1166 VGND 0.0057f
C21445 VPWR.n1167 VGND 3.84e-19
C21446 VPWR.n1168 VGND 0.00524f
C21447 VPWR.t1374 VGND 6.73e-19
C21448 VPWR.t1189 VGND 9.96e-19
C21449 VPWR.n1169 VGND 0.0018f
C21450 VPWR.n1170 VGND 0.00488f
C21451 VPWR.n1171 VGND 3.94e-19
C21452 VPWR.n1172 VGND 0.00524f
C21453 VPWR.t1094 VGND 0.00166f
C21454 VPWR.t1106 VGND 0.0016f
C21455 VPWR.n1173 VGND 0.00353f
C21456 VPWR.n1174 VGND 0.00557f
C21457 VPWR.n1175 VGND 0.00524f
C21458 VPWR.n1176 VGND 0.00128f
C21459 VPWR.n1177 VGND 0.00524f
C21460 VPWR.t1100 VGND 0.00166f
C21461 VPWR.t1102 VGND 0.00166f
C21462 VPWR.n1178 VGND 0.00359f
C21463 VPWR.n1179 VGND 0.00636f
C21464 VPWR.n1180 VGND 0.00524f
C21465 VPWR.n1181 VGND 0.00153f
C21466 VPWR.n1182 VGND 0.00524f
C21467 VPWR.t1104 VGND 0.00166f
C21468 VPWR.t1108 VGND 0.00166f
C21469 VPWR.n1183 VGND 0.00353f
C21470 VPWR.t2363 VGND 0.00234f
C21471 VPWR.n1184 VGND 0.00392f
C21472 VPWR.n1185 VGND 0.0042f
C21473 VPWR.n1186 VGND 9.65e-19
C21474 VPWR.n1187 VGND 0.00524f
C21475 VPWR.n1188 VGND 0.00134f
C21476 VPWR.n1189 VGND 0.00524f
C21477 VPWR.t1112 VGND 0.00166f
C21478 VPWR.t1082 VGND 0.00166f
C21479 VPWR.n1190 VGND 0.00359f
C21480 VPWR.n1191 VGND 0.00622f
C21481 VPWR.n1192 VGND 0.00524f
C21482 VPWR.n1193 VGND 0.00524f
C21483 VPWR.n1194 VGND 0.0031f
C21484 VPWR.n1195 VGND 0.00524f
C21485 VPWR.t37 VGND 0.00387f
C21486 VPWR.n1196 VGND 0.00493f
C21487 VPWR.n1197 VGND 0.00507f
C21488 VPWR.n1198 VGND 0.00393f
C21489 VPWR.n1199 VGND 0.00199f
C21490 VPWR.n1200 VGND 0.00199f
C21491 VPWR.n1201 VGND 0.00977f
C21492 VPWR.t503 VGND 0.0463f
C21493 VPWR.t1765 VGND 0.0111f
C21494 VPWR.t3239 VGND 0.0141f
C21495 VPWR.t1814 VGND 0.0141f
C21496 VPWR.t3237 VGND 0.0161f
C21497 VPWR.t1651 VGND 0.0211f
C21498 VPWR.t2974 VGND 0.0107f
C21499 VPWR.t2965 VGND 0.0149f
C21500 VPWR.t879 VGND 0.0126f
C21501 VPWR.t1002 VGND 0.0171f
C21502 VPWR.t1816 VGND 0.0228f
C21503 VPWR.t1653 VGND 0.0173f
C21504 VPWR.t1272 VGND 0.0144f
C21505 VPWR.t1799 VGND 0.0163f
C21506 VPWR.t1381 VGND 0.0149f
C21507 VPWR.t3105 VGND 0.0331f
C21508 VPWR.t2356 VGND 0.0332f
C21509 VPWR.t1262 VGND 0.0166f
C21510 VPWR.t1813 VGND 0.0144f
C21511 VPWR.t1260 VGND 0.0144f
C21512 VPWR.t1003 VGND 0.0144f
C21513 VPWR.t1258 VGND 0.0141f
C21514 VPWR.t2773 VGND 0.0144f
C21515 VPWR.t1264 VGND 0.0181f
C21516 VPWR.t1375 VGND 0.0161f
C21517 VPWR.t2529 VGND 0.00906f
C21518 VPWR.t1004 VGND 0.0153f
C21519 VPWR.t2775 VGND 0.0311f
C21520 VPWR.t3052 VGND 0.0154f
C21521 VPWR.t1554 VGND 0.026f
C21522 VPWR.t36 VGND 0.0312f
C21523 VPWR.t1795 VGND 0.0305f
C21524 VPWR.t2430 VGND 0.0213f
C21525 VPWR.t2919 VGND 0.018f
C21526 VPWR.n1202 VGND 0.0244f
C21527 VPWR.t1777 VGND 0.0139f
C21528 VPWR.t1085 VGND 0.0141f
C21529 VPWR.t2873 VGND 0.0144f
C21530 VPWR.t1081 VGND 0.0178f
C21531 VPWR.t1111 VGND 0.0289f
C21532 VPWR.t1107 VGND 0.027f
C21533 VPWR.t2362 VGND 0.0144f
C21534 VPWR.t1103 VGND 0.0154f
C21535 VPWR.t2003 VGND 0.0144f
C21536 VPWR.t1101 VGND 0.0153f
C21537 VPWR.t1099 VGND 0.0158f
C21538 VPWR.t2875 VGND 0.0144f
C21539 VPWR.t1105 VGND 0.0235f
C21540 VPWR.t1188 VGND 0.0143f
C21541 VPWR.t1093 VGND 0.0163f
C21542 VPWR.t1373 VGND 0.0144f
C21543 VPWR.t1089 VGND 0.0164f
C21544 VPWR.t1097 VGND 0.0289f
C21545 VPWR.t1095 VGND 0.0166f
C21546 VPWR.t1508 VGND 0.0144f
C21547 VPWR.t1091 VGND 0.0166f
C21548 VPWR.t2876 VGND 0.0144f
C21549 VPWR.t1087 VGND 0.0144f
C21550 VPWR.t2002 VGND 0.0144f
C21551 VPWR.t1109 VGND 0.0141f
C21552 VPWR.t1540 VGND 0.0144f
C21553 VPWR.t1083 VGND 0.0181f
C21554 VPWR.t1379 VGND 0.0144f
C21555 VPWR.t1049 VGND 0.0141f
C21556 VPWR.t3261 VGND 0.0144f
C21557 VPWR.t1053 VGND 0.0215f
C21558 VPWR.t1051 VGND 0.0289f
C21559 VPWR.t1073 VGND 0.0146f
C21560 VPWR.t1538 VGND 0.00537f
C21561 VPWR.t2032 VGND 0.0257f
C21562 VPWR.t2721 VGND 0.0151f
C21563 VPWR.t509 VGND 0.0052f
C21564 VPWR.t677 VGND 0.0109f
C21565 VPWR.t2525 VGND 0.0163f
C21566 VPWR.t758 VGND 0.03f
C21567 VPWR.t760 VGND 0.0223f
C21568 VPWR.n1203 VGND 0.0246f
C21569 VPWR.t2387 VGND 0.0181f
C21570 VPWR.t184 VGND 0.0141f
C21571 VPWR.t3316 VGND 0.0215f
C21572 VPWR.t1128 VGND 0.0282f
C21573 VPWR.t1123 VGND 0.0175f
C21574 VPWR.t2634 VGND 0.0175f
C21575 VPWR.t2630 VGND 0.0198f
C21576 VPWR.t2638 VGND 0.0225f
C21577 VPWR.t2632 VGND 0.0227f
C21578 VPWR.t2636 VGND 0.0109f
C21579 VPWR.t1779 VGND 0.0141f
C21580 VPWR.t2628 VGND 0.0141f
C21581 VPWR.t1034 VGND 0.0141f
C21582 VPWR.t1126 VGND 0.0228f
C21583 VPWR.t1124 VGND 0.0279f
C21584 VPWR.t2083 VGND 0.0156f
C21585 VPWR.t1565 VGND 0.0247f
C21586 VPWR.t1036 VGND 0.018f
C21587 VPWR.t652 VGND 0.0235f
C21588 VPWR.t2311 VGND 0.0358f
C21589 VPWR.t2840 VGND 0.0109f
C21590 VPWR.t1837 VGND 0.0223f
C21591 VPWR.t790 VGND 0.0248f
C21592 VPWR.t2369 VGND 0.0274f
C21593 VPWR.t1037 VGND 0.0311f
C21594 VPWR.t1566 VGND 0.0175f
C21595 VPWR.t1726 VGND 0.0141f
C21596 VPWR.t1966 VGND 0.0154f
C21597 VPWR.t1451 VGND 0.0181f
C21598 VPWR.t2836 VGND 0.0166f
C21599 VPWR.t789 VGND 0.0141f
C21600 VPWR.t3284 VGND 0.0235f
C21601 VPWR.t3282 VGND 0.0285f
C21602 VPWR.t1369 VGND 0.0238f
C21603 VPWR.t1968 VGND 0.0311f
C21604 VPWR.n1204 VGND 0.029f
C21605 VPWR.t1252 VGND 0.0126f
C21606 VPWR.t792 VGND 0.00822f
C21607 VPWR.t3156 VGND 0.0144f
C21608 VPWR.t1452 VGND 0.0144f
C21609 VPWR.t3150 VGND 0.0141f
C21610 VPWR.t1852 VGND 0.0144f
C21611 VPWR.t3152 VGND 0.0181f
C21612 VPWR.t1371 VGND 0.0144f
C21613 VPWR.t3154 VGND 0.0141f
C21614 VPWR.t1793 VGND 0.0144f
C21615 VPWR.t1590 VGND 0.0164f
C21616 VPWR.t1587 VGND 0.0289f
C21617 VPWR.t1594 VGND 0.0196f
C21618 VPWR.t1854 VGND 0.0144f
C21619 VPWR.t1581 VGND 0.0205f
C21620 VPWR.t1579 VGND 0.0117f
C21621 VPWR.t3032 VGND 0.0144f
C21622 VPWR.t1585 VGND 0.0141f
C21623 VPWR.t918 VGND 0.0144f
C21624 VPWR.t1583 VGND 0.0206f
C21625 VPWR.t1604 VGND 0.026f
C21626 VPWR.t474 VGND 0.0144f
C21627 VPWR.t1577 VGND 0.0171f
C21628 VPWR.t1596 VGND 0.0289f
C21629 VPWR.t1592 VGND 0.019f
C21630 VPWR.t1600 VGND 0.0243f
C21631 VPWR.t1598 VGND 0.0161f
C21632 VPWR.t1038 VGND 0.0144f
C21633 VPWR.t1575 VGND 0.0159f
C21634 VPWR.t923 VGND 0.0144f
C21635 VPWR.t1602 VGND 0.0156f
C21636 VPWR.t2539 VGND 0.0185f
C21637 VPWR.t1632 VGND 0.0193f
C21638 VPWR.t1636 VGND 0.026f
C21639 VPWR.t735 VGND 0.0294f
C21640 VPWR.t921 VGND 0.0356f
C21641 VPWR.t3067 VGND 0.0339f
C21642 VPWR.n1205 VGND 0.0235f
C21643 VPWR.t1311 VGND 0.0183f
C21644 VPWR.t249 VGND 0.0141f
C21645 VPWR.t1693 VGND 0.0279f
C21646 VPWR.t3065 VGND 0.0117f
C21647 VPWR.t2172 VGND 0.0141f
C21648 VPWR.t950 VGND 0.0141f
C21649 VPWR.t2604 VGND 0.0144f
C21650 VPWR.t1514 VGND 0.0206f
C21651 VPWR.t762 VGND 0.0339f
C21652 VPWR.t1699 VGND 0.0493f
C21653 VPWR.t1940 VGND 0.023f
C21654 VPWR.t157 VGND 0.0235f
C21655 VPWR.t1517 VGND 0.0334f
C21656 VPWR.t951 VGND 0.0321f
C21657 VPWR.t2254 VGND 0.0336f
C21658 VPWR.t1910 VGND 0.00873f
C21659 VPWR.t1515 VGND 0.0141f
C21660 VPWR.t1938 VGND 0.0141f
C21661 VPWR.t1908 VGND 0.00587f
C21662 VPWR.t834 VGND 0.0265f
C21663 VPWR.t1979 VGND 0.0304f
C21664 VPWR.t1936 VGND 0.0304f
C21665 VPWR.t594 VGND 0.0201f
C21666 VPWR.t1169 VGND 0.0217f
C21667 VPWR.t1697 VGND 0.0319f
C21668 VPWR.t2395 VGND 0.0282f
C21669 VPWR.t2397 VGND 0.0269f
C21670 VPWR.t1937 VGND 0.0171f
C21671 VPWR.t1978 VGND 0.018f
C21672 VPWR.n1206 VGND 0.0158f
C21673 VPWR.n1207 VGND 0.0108f
C21674 VPWR.n1208 VGND 0.00274f
C21675 VPWR.n1209 VGND 0.00247f
C21676 VPWR.n1210 VGND 0.0031f
C21677 VPWR.n1211 VGND 0.00135f
C21678 VPWR.n1212 VGND 0.00524f
C21679 VPWR.t3228 VGND 0.00148f
C21680 VPWR.t1696 VGND 9.71e-19
C21681 VPWR.n1213 VGND 0.00358f
C21682 VPWR.n1214 VGND 0.00613f
C21683 VPWR.t839 VGND 0.00569f
C21684 VPWR.t3171 VGND 0.00557f
C21685 VPWR.n1215 VGND 0.00756f
C21686 VPWR.n1216 VGND 0.0139f
C21687 VPWR.n1217 VGND 5.44e-19
C21688 VPWR.n1218 VGND 0.00524f
C21689 VPWR.n1219 VGND 0.00172f
C21690 VPWR.n1220 VGND 0.00524f
C21691 VPWR.n1221 VGND 0.00179f
C21692 VPWR.n1222 VGND 0.00524f
C21693 VPWR.n1223 VGND 0.00524f
C21694 VPWR.n1224 VGND 0.00387f
C21695 VPWR.n1225 VGND 9.42e-19
C21696 VPWR.n1226 VGND 0.00131f
C21697 VPWR.n1227 VGND 5.98e-19
C21698 VPWR.n1228 VGND 3.42e-19
C21699 VPWR.n1229 VGND 1.99e-19
C21700 VPWR.n1230 VGND 1.76e-19
C21701 VPWR.n1231 VGND 3.07e-19
C21702 VPWR.n1232 VGND 5.48e-19
C21703 VPWR.n1234 VGND 0.1f
C21704 VPWR.n1235 VGND 0.1f
C21705 VPWR.n1236 VGND 6.54e-19
C21706 VPWR.n1237 VGND 8.67e-19
C21707 VPWR.n1238 VGND 4.39e-19
C21708 VPWR.n1239 VGND 3.29e-19
C21709 VPWR.n1240 VGND 5.27e-19
C21710 VPWR.n1241 VGND 2.85e-19
C21711 VPWR.n1242 VGND 2.85e-19
C21712 VPWR.n1243 VGND 4.17e-19
C21713 VPWR.n1244 VGND 5.71e-19
C21714 VPWR.n1245 VGND 4.17e-19
C21715 VPWR.n1246 VGND 3.51e-19
C21716 VPWR.n1247 VGND 4.61e-19
C21717 VPWR.n1248 VGND 4.17e-19
C21718 VPWR.n1249 VGND 4.83e-19
C21719 VPWR.n1250 VGND 4.61e-19
C21720 VPWR.n1251 VGND 3.73e-19
C21721 VPWR.n1252 VGND 2.41e-19
C21722 VPWR.n1253 VGND 4.83e-19
C21723 VPWR.n1254 VGND 4.61e-19
C21724 VPWR.n1255 VGND 4.11e-19
C21725 VPWR.n1256 VGND 4.11e-19
C21726 VPWR.n1257 VGND 7.39e-19
C21727 VPWR.n1258 VGND 5.19e-19
C21728 VPWR.n1259 VGND 7.39e-19
C21729 VPWR.n1260 VGND 4.11e-19
C21730 VPWR.n1261 VGND 4.11e-19
C21731 VPWR.n1263 VGND 0.0057f
C21732 VPWR.n1264 VGND 8.67e-19
C21733 VPWR.n1265 VGND 6.54e-19
C21734 VPWR.n1266 VGND 9.06e-19
C21735 VPWR.n1267 VGND 0.00139f
C21736 VPWR.n1268 VGND 5.27e-19
C21737 VPWR.n1269 VGND 3.95e-19
C21738 VPWR.n1270 VGND 5.05e-19
C21739 VPWR.n1271 VGND 5.05e-19
C21740 VPWR.t2725 VGND 0.00618f
C21741 VPWR.t3560 VGND 0.0592f
C21742 VPWR.n1272 VGND 0.0356f
C21743 VPWR.t3268 VGND 0.00385f
C21744 VPWR.n1273 VGND 0.00351f
C21745 VPWR.t605 VGND 0.00387f
C21746 VPWR.n1274 VGND 0.00837f
C21747 VPWR.n1275 VGND 0.00524f
C21748 VPWR.t3467 VGND 0.0231f
C21749 VPWR.t1392 VGND 0.00136f
C21750 VPWR.t1208 VGND 0.00136f
C21751 VPWR.n1276 VGND 0.00317f
C21752 VPWR.t3401 VGND 0.00911f
C21753 VPWR.t417 VGND 0.00391f
C21754 VPWR.n1277 VGND 0.0253f
C21755 VPWR.t416 VGND 0.00391f
C21756 VPWR.n1279 VGND 0.0138f
C21757 VPWR.t3352 VGND 0.00911f
C21758 VPWR.t730 VGND 0.00391f
C21759 VPWR.n1280 VGND 0.0253f
C21760 VPWR.t731 VGND 0.00391f
C21761 VPWR.n1282 VGND 0.0138f
C21762 VPWR.n1283 VGND 0.0109f
C21763 VPWR.t1660 VGND 0.00136f
C21764 VPWR.t3173 VGND 0.00136f
C21765 VPWR.n1284 VGND 0.0032f
C21766 VPWR.n1285 VGND 0.00393f
C21767 VPWR.n1286 VGND 0.00345f
C21768 VPWR.n1287 VGND 0.00444f
C21769 VPWR.t3445 VGND 0.00911f
C21770 VPWR.t271 VGND 0.00391f
C21771 VPWR.n1288 VGND 0.0253f
C21772 VPWR.t272 VGND 0.00391f
C21773 VPWR.n1290 VGND 0.0138f
C21774 VPWR.n1291 VGND 0.0143f
C21775 VPWR.n1292 VGND 0.00487f
C21776 VPWR.t604 VGND 0.00387f
C21777 VPWR.n1293 VGND 0.00837f
C21778 VPWR.n1294 VGND 0.0439f
C21779 VPWR.t3270 VGND 0.00614f
C21780 VPWR.n1295 VGND 0.0133f
C21781 VPWR.n1296 VGND 0.00702f
C21782 VPWR.n1297 VGND 0.013f
C21783 VPWR.n1298 VGND 0.0136f
C21784 VPWR.n1299 VGND 0.0031f
C21785 VPWR.n1300 VGND 0.00393f
C21786 VPWR.n1301 VGND 0.00524f
C21787 VPWR.n1302 VGND 0.0031f
C21788 VPWR.n1303 VGND 0.00607f
C21789 VPWR.n1304 VGND 0.00347f
C21790 VPWR.t2659 VGND 9.22e-19
C21791 VPWR.n1305 VGND 0.00265f
C21792 VPWR.n1306 VGND 0.00333f
C21793 VPWR.n1307 VGND 0.00128f
C21794 VPWR.n1308 VGND 0.00393f
C21795 VPWR.t111 VGND 0.00463f
C21796 VPWR.n1309 VGND 0.00567f
C21797 VPWR.n1310 VGND 0.00588f
C21798 VPWR.n1311 VGND 0.00524f
C21799 VPWR.n1312 VGND 0.00337f
C21800 VPWR.n1313 VGND 0.00524f
C21801 VPWR.t2788 VGND 0.00115f
C21802 VPWR.t1921 VGND 6.73e-19
C21803 VPWR.n1314 VGND 0.00192f
C21804 VPWR.n1315 VGND 0.00673f
C21805 VPWR.n1316 VGND 0.00499f
C21806 VPWR.n1317 VGND 0.00307f
C21807 VPWR.n1318 VGND 0.00179f
C21808 VPWR.n1319 VGND 0.00158f
C21809 VPWR.n1320 VGND 0.00786f
C21810 VPWR.n1321 VGND 0.00588f
C21811 VPWR.n1322 VGND 0.00651f
C21812 VPWR.n1323 VGND 0.0111f
C21813 VPWR.t1861 VGND 0.00581f
C21814 VPWR.t1863 VGND 0.00581f
C21815 VPWR.n1324 VGND 0.00607f
C21816 VPWR.n1325 VGND 0.0101f
C21817 VPWR.n1326 VGND 0.00536f
C21818 VPWR.n1327 VGND 9e-19
C21819 VPWR.n1328 VGND 0.00138f
C21820 VPWR.n1329 VGND 9.06e-19
C21821 VPWR.n1330 VGND 5.48e-19
C21822 VPWR.n1331 VGND 6.14e-19
C21823 VPWR.n1332 VGND 0.00138f
C21824 VPWR.n1333 VGND 0.00408f
C21825 VPWR.n1334 VGND 0.00276f
C21826 VPWR.n1335 VGND 0.00153f
C21827 VPWR.n1336 VGND 6.1e-19
C21828 VPWR.n1337 VGND 4.27e-19
C21829 VPWR.n1338 VGND 1.14e-19
C21830 VPWR.n1339 VGND 0.00326f
C21831 VPWR.n1340 VGND 4.27e-19
C21832 VPWR.n1341 VGND 6.83e-19
C21833 VPWR.n1342 VGND 3.7e-19
C21834 VPWR.n1343 VGND 9.68e-19
C21835 VPWR.n1344 VGND 9.96e-19
C21836 VPWR.n1345 VGND 5.41e-19
C21837 VPWR.n1346 VGND 7.4e-19
C21838 VPWR.n1347 VGND 6.1e-19
C21839 VPWR.n1348 VGND 0.00316f
C21840 VPWR.n1349 VGND 3.13e-19
C21841 VPWR.n1350 VGND 2.56e-19
C21842 VPWR.n1351 VGND 4.55e-19
C21843 VPWR.n1352 VGND 0.00276f
C21844 VPWR.n1353 VGND 9.68e-19
C21845 VPWR.n1354 VGND 9.96e-19
C21846 VPWR.n1355 VGND 3.13e-19
C21847 VPWR.n1356 VGND 4.84e-19
C21848 VPWR.n1357 VGND 6.83e-19
C21849 VPWR.n1358 VGND 0.00248f
C21850 VPWR.n1359 VGND 4.84e-19
C21851 VPWR.t2720 VGND 0.00757f
C21852 VPWR.n1360 VGND 0.00485f
C21853 VPWR.n1361 VGND 3.59e-19
C21854 VPWR.n1362 VGND 4.27e-19
C21855 VPWR.n1363 VGND 4.66e-19
C21856 VPWR.n1364 VGND 4.27e-19
C21857 VPWR.n1365 VGND 0.00309f
C21858 VPWR.n1366 VGND 6.26e-19
C21859 VPWR.n1367 VGND 4.84e-19
C21860 VPWR.n1368 VGND 3.42e-19
C21861 VPWR.n1369 VGND 5.98e-19
C21862 VPWR.t112 VGND 0.0046f
C21863 VPWR.n1370 VGND 0.00378f
C21864 VPWR.n1371 VGND 0.00123f
C21865 VPWR.t2409 VGND 0.00618f
C21866 VPWR.n1372 VGND 0.00786f
C21867 VPWR.t415 VGND 0.0515f
C21868 VPWR.t1659 VGND 0.0463f
C21869 VPWR.t270 VGND 0.0148f
C21870 VPWR.t3172 VGND 0.0183f
C21871 VPWR.t1391 VGND 0.0354f
C21872 VPWR.t1207 VGND 0.0257f
C21873 VPWR.t603 VGND 0.021f
C21874 VPWR.t3269 VGND 0.0302f
C21875 VPWR.t3267 VGND 0.0253f
C21876 VPWR.t2658 VGND 0.0336f
C21877 VPWR.t2787 VGND 0.0321f
C21878 VPWR.t1920 VGND 0.028f
C21879 VPWR.t2724 VGND 0.0203f
C21880 VPWR.t110 VGND 0.0141f
C21881 VPWR.t1860 VGND 0.0299f
C21882 VPWR.t1862 VGND 0.0416f
C21883 VPWR.t2723 VGND 0.0282f
C21884 VPWR.t2719 VGND 0.0458f
C21885 VPWR.t1542 VGND 0.0247f
C21886 VPWR.t2412 VGND 0.0282f
C21887 VPWR.t2644 VGND 0.0416f
C21888 VPWR.t2646 VGND 0.0436f
C21889 VPWR.t2408 VGND 0.0264f
C21890 VPWR.t376 VGND 0.0126f
C21891 VPWR.n1373 VGND 0.0451f
C21892 VPWR.n1374 VGND 0.0066f
C21893 VPWR.t904 VGND 0.00676f
C21894 VPWR.n1375 VGND 0.0119f
C21895 VPWR.t378 VGND 0.0046f
C21896 VPWR.n1376 VGND 0.00407f
C21897 VPWR.t1271 VGND 0.0024f
C21898 VPWR.t443 VGND 0.0046f
C21899 VPWR.n1377 VGND 0.00407f
C21900 VPWR.t444 VGND 0.0046f
C21901 VPWR.n1378 VGND 0.00407f
C21902 VPWR.t2609 VGND 0.00102f
C21903 VPWR.t864 VGND 0.00154f
C21904 VPWR.n1379 VGND 0.00495f
C21905 VPWR.n1380 VGND 0.00787f
C21906 VPWR.t2210 VGND 0.00102f
C21907 VPWR.t1913 VGND 0.00102f
C21908 VPWR.n1381 VGND 0.00221f
C21909 VPWR.n1382 VGND 0.00626f
C21910 VPWR.t3529 VGND 0.0179f
C21911 VPWR.t19 VGND 0.00395f
C21912 VPWR.n1383 VGND 0.028f
C21913 VPWR.t20 VGND 0.00432f
C21914 VPWR.t807 VGND 0.00634f
C21915 VPWR.n1384 VGND 0.00976f
C21916 VPWR.t803 VGND 0.0016f
C21917 VPWR.t805 VGND 0.0016f
C21918 VPWR.n1385 VGND 0.00367f
C21919 VPWR.t903 VGND 0.0462f
C21920 VPWR.t1270 VGND 0.0245f
C21921 VPWR.t990 VGND 0.0322f
C21922 VPWR.t901 VGND 0.0322f
C21923 VPWR.t2777 VGND 0.0285f
C21924 VPWR.t2208 VGND 0.0311f
C21925 VPWR.t2670 VGND 0.0264f
C21926 VPWR.t442 VGND 0.0331f
C21927 VPWR.t956 VGND 0.0396f
C21928 VPWR.t1841 VGND 0.0398f
C21929 VPWR.t2211 VGND 0.0401f
C21930 VPWR.t2778 VGND 0.0247f
C21931 VPWR.t1657 VGND 0.0311f
C21932 VPWR.t863 VGND 0.0399f
C21933 VPWR.t2608 VGND 0.0211f
C21934 VPWR.t2209 VGND 0.0121f
C21935 VPWR.t3315 VGND 0.0141f
C21936 VPWR.t1912 VGND 0.0178f
C21937 VPWR.t637 VGND 0.0312f
C21938 VPWR.t18 VGND 0.0206f
C21939 VPWR.t806 VGND 0.026f
C21940 VPWR.t802 VGND 0.0126f
C21941 VPWR.t2798 VGND 0.0126f
C21942 VPWR.t2955 VGND 0.0154f
C21943 VPWR.t457 VGND 0.0312f
C21944 VPWR.t2953 VGND 0.0423f
C21945 VPWR.t2339 VGND 0.0457f
C21946 VPWR.t2337 VGND 0.0196f
C21947 VPWR.t3040 VGND 0.0153f
C21948 VPWR.t3046 VGND 0.0109f
C21949 VPWR.t3005 VGND 0.0201f
C21950 VPWR.t3044 VGND 0.0264f
C21951 VPWR.t1637 VGND 0.0158f
C21952 VPWR.t2545 VGND 0.0141f
C21953 VPWR.t1639 VGND 0.0161f
C21954 VPWR.t1634 VGND 0.0171f
C21955 VPWR.t2543 VGND 0.0161f
C21956 VPWR.t2239 VGND 0.0141f
C21957 VPWR.t2537 VGND 0.0324f
C21958 VPWR.t2075 VGND 0.0094f
C21959 VPWR.t2606 VGND 0.0183f
C21960 VPWR.t2541 VGND 0.0141f
C21961 VPWR.t2177 VGND 0.0173f
C21962 VPWR.t2238 VGND 0.0181f
C21963 VPWR.t1522 VGND 0.0309f
C21964 VPWR.t920 VGND 0.0171f
C21965 VPWR.t2897 VGND 0.0144f
C21966 VPWR.t1303 VGND 0.0161f
C21967 VPWR.t2535 VGND 0.0141f
C21968 VPWR.t1305 VGND 0.0144f
C21969 VPWR.t798 VGND 0.0279f
C21970 VPWR.t808 VGND 0.0144f
C21971 VPWR.t800 VGND 0.0282f
C21972 VPWR.t804 VGND 0.0195f
C21973 VPWR.n1386 VGND 0.0176f
C21974 VPWR.n1387 VGND 0.00126f
C21975 VPWR.t801 VGND 0.0016f
C21976 VPWR.t809 VGND 0.0016f
C21977 VPWR.n1388 VGND 0.00379f
C21978 VPWR.n1389 VGND 0.00819f
C21979 VPWR.n1390 VGND 9.28e-19
C21980 VPWR.n1391 VGND 4.55e-19
C21981 VPWR.n1392 VGND 1.31e-19
C21982 VPWR.n1393 VGND 3.7e-19
C21983 VPWR.n1394 VGND 1.21e-19
C21984 VPWR.n1395 VGND 3.42e-19
C21985 VPWR.n1396 VGND 5.65e-19
C21986 VPWR.n1397 VGND 3.7e-19
C21987 VPWR.n1398 VGND 6.26e-19
C21988 VPWR.n1399 VGND 1.76e-19
C21989 VPWR.n1400 VGND 4.39e-19
C21990 VPWR.n1401 VGND 6.14e-19
C21991 VPWR.n1402 VGND 4.17e-19
C21992 VPWR.n1403 VGND 5.05e-19
C21993 VPWR.n1404 VGND 6.55e-19
C21994 VPWR.n1405 VGND 5.41e-19
C21995 VPWR.n1406 VGND 9.96e-19
C21996 VPWR.n1407 VGND 9.68e-19
C21997 VPWR.n1408 VGND 5.41e-19
C21998 VPWR.t2536 VGND 7.22e-19
C21999 VPWR.t2898 VGND 9.22e-19
C22000 VPWR.n1409 VGND 0.00189f
C22001 VPWR.n1410 VGND 0.00367f
C22002 VPWR.t1304 VGND 0.00631f
C22003 VPWR.n1411 VGND 0.0053f
C22004 VPWR.n1412 VGND 8.07e-19
C22005 VPWR.n1413 VGND 3.13e-19
C22006 VPWR.n1414 VGND 5.98e-19
C22007 VPWR.n1415 VGND 5.12e-19
C22008 VPWR.n1416 VGND 0.00108f
C22009 VPWR.n1417 VGND 0.00122f
C22010 VPWR.n1418 VGND 3.13e-19
C22011 VPWR.n1419 VGND 5.12e-19
C22012 VPWR.n1420 VGND 4.64e-19
C22013 VPWR.n1421 VGND 6.26e-19
C22014 VPWR.n1422 VGND 1.71e-19
C22015 VPWR.n1423 VGND 2.28e-19
C22016 VPWR.n1424 VGND 2.85e-19
C22017 VPWR.n1425 VGND 2.52e-19
C22018 VPWR.n1426 VGND 0.00259f
C22019 VPWR.t799 VGND 0.0016f
C22020 VPWR.t1306 VGND 0.0016f
C22021 VPWR.n1427 VGND 0.00377f
C22022 VPWR.n1428 VGND 0.0053f
C22023 VPWR.n1429 VGND 0.00105f
C22024 VPWR.n1430 VGND 0.00364f
C22025 VPWR.n1431 VGND 0.00333f
C22026 VPWR.n1432 VGND 0.00393f
C22027 VPWR.n1433 VGND 0.00199f
C22028 VPWR.n1434 VGND 0.00908f
C22029 VPWR.n1435 VGND 0.00672f
C22030 VPWR.n1436 VGND 0.00169f
C22031 VPWR.n1437 VGND 0.0031f
C22032 VPWR.n1438 VGND 0.00393f
C22033 VPWR.n1439 VGND 5.24e-19
C22034 VPWR.n1440 VGND 0.0295f
C22035 VPWR.n1441 VGND 0.00139f
C22036 VPWR.n1442 VGND 0.0031f
C22037 VPWR.t3572 VGND 0.00911f
C22038 VPWR.t638 VGND 0.00391f
C22039 VPWR.n1443 VGND 0.0253f
C22040 VPWR.t639 VGND 0.00391f
C22041 VPWR.n1445 VGND 0.0126f
C22042 VPWR.n1446 VGND 0.00609f
C22043 VPWR.n1447 VGND 0.00393f
C22044 VPWR.n1448 VGND 0.00199f
C22045 VPWR.n1449 VGND 0.00186f
C22046 VPWR.n1450 VGND 0.0015f
C22047 VPWR.n1451 VGND 0.0031f
C22048 VPWR.n1452 VGND 0.00524f
C22049 VPWR.n1453 VGND 0.00524f
C22050 VPWR.n1454 VGND 7.56e-19
C22051 VPWR.n1455 VGND 0.00524f
C22052 VPWR.n1456 VGND 0.00475f
C22053 VPWR.t1658 VGND 0.00238f
C22054 VPWR.n1457 VGND 0.00521f
C22055 VPWR.n1458 VGND 0.00267f
C22056 VPWR.n1459 VGND 0.0031f
C22057 VPWR.n1460 VGND 0.00639f
C22058 VPWR.n1461 VGND 0.00524f
C22059 VPWR.n1462 VGND 0.0066f
C22060 VPWR.n1463 VGND 0.00524f
C22061 VPWR.n1464 VGND 0.00506f
C22062 VPWR.n1465 VGND 0.00524f
C22063 VPWR.t957 VGND 6.73e-19
C22064 VPWR.t1842 VGND 9.96e-19
C22065 VPWR.n1466 VGND 0.00176f
C22066 VPWR.n1467 VGND 0.00658f
C22067 VPWR.n1468 VGND 0.00484f
C22068 VPWR.n1469 VGND 0.00524f
C22069 VPWR.n1470 VGND 0.00553f
C22070 VPWR.n1471 VGND 0.00524f
C22071 VPWR.t2671 VGND 0.00453f
C22072 VPWR.n1472 VGND 0.00799f
C22073 VPWR.n1473 VGND 0.00438f
C22074 VPWR.n1474 VGND 0.00524f
C22075 VPWR.t3416 VGND 0.0592f
C22076 VPWR.n1475 VGND 0.0356f
C22077 VPWR.n1476 VGND 0.00484f
C22078 VPWR.n1477 VGND 0.00524f
C22079 VPWR.n1478 VGND 0.00506f
C22080 VPWR.n1479 VGND 0.00524f
C22081 VPWR.n1480 VGND 0.00614f
C22082 VPWR.n1481 VGND 0.00524f
C22083 VPWR.t991 VGND 6.73e-19
C22084 VPWR.t902 VGND 0.00127f
C22085 VPWR.n1482 VGND 0.00203f
C22086 VPWR.n1483 VGND 0.00594f
C22087 VPWR.n1484 VGND 0.00355f
C22088 VPWR.n1485 VGND 0.00524f
C22089 VPWR.n1486 VGND 0.00475f
C22090 VPWR.n1487 VGND 0.00166f
C22091 VPWR.n1488 VGND 0.00564f
C22092 VPWR.n1489 VGND 0.00119f
C22093 VPWR.n1490 VGND 0.0031f
C22094 VPWR.n1491 VGND 0.00323f
C22095 VPWR.n1492 VGND 0.00524f
C22096 VPWR.n1493 VGND 0.00393f
C22097 VPWR.n1494 VGND 0.00646f
C22098 VPWR.n1495 VGND 0.0066f
C22099 VPWR.n1496 VGND 0.00333f
C22100 VPWR.n1497 VGND 0.00393f
C22101 VPWR.n1498 VGND 0.00199f
C22102 VPWR.n1499 VGND 0.0147f
C22103 VPWR.n1500 VGND 0.00334f
C22104 VPWR.n1501 VGND 0.0031f
C22105 VPWR.t3385 VGND 0.0592f
C22106 VPWR.n1502 VGND 0.0356f
C22107 VPWR.n1503 VGND 0.00481f
C22108 VPWR.n1504 VGND 0.00524f
C22109 VPWR.t2645 VGND 0.00584f
C22110 VPWR.t2647 VGND 0.00584f
C22111 VPWR.n1505 VGND 0.00573f
C22112 VPWR.n1506 VGND 0.0108f
C22113 VPWR.n1507 VGND 0.00334f
C22114 VPWR.n1508 VGND 0.00524f
C22115 VPWR.n1509 VGND 0.00502f
C22116 VPWR.n1510 VGND 0.00524f
C22117 VPWR.n1511 VGND 0.00639f
C22118 VPWR.n1512 VGND 0.00524f
C22119 VPWR.t1543 VGND 0.00757f
C22120 VPWR.n1513 VGND 0.00609f
C22121 VPWR.t377 VGND 0.0046f
C22122 VPWR.n1514 VGND 0.00407f
C22123 VPWR.n1515 VGND 0.00251f
C22124 VPWR.n1516 VGND 0.00475f
C22125 VPWR.n1517 VGND 0.00174f
C22126 VPWR.n1518 VGND 0.00131f
C22127 VPWR.n1519 VGND 9.42e-19
C22128 VPWR.n1520 VGND 2.63e-19
C22129 VPWR.n1521 VGND 1.76e-19
C22130 VPWR.n1522 VGND 3.07e-19
C22131 VPWR.n1523 VGND 5.48e-19
C22132 VPWR.n1525 VGND 0.1f
C22133 VPWR.n1526 VGND 0.1f
C22134 VPWR.n1527 VGND 0.0194f
C22135 VPWR.n1528 VGND 8.67e-19
C22136 VPWR.n1529 VGND 6.54e-19
C22137 VPWR.n1530 VGND 9.06e-19
C22138 VPWR.n1531 VGND 0.00139f
C22139 VPWR.n1532 VGND 5.27e-19
C22140 VPWR.n1533 VGND 3.95e-19
C22141 VPWR.n1534 VGND 5.05e-19
C22142 VPWR.n1535 VGND 5.05e-19
C22143 VPWR.n1536 VGND 3.07e-19
C22144 VPWR.n1537 VGND 5.48e-19
C22145 VPWR.t3502 VGND 0.0289f
C22146 VPWR.t716 VGND 0.00387f
C22147 VPWR.n1539 VGND 0.0604f
C22148 VPWR.n1540 VGND 0.0146f
C22149 VPWR.n1541 VGND 0.0117f
C22150 VPWR.t983 VGND 6.73e-19
C22151 VPWR.t1287 VGND 0.00127f
C22152 VPWR.n1542 VGND 0.00204f
C22153 VPWR.n1543 VGND 0.0143f
C22154 VPWR.t1316 VGND 0.00644f
C22155 VPWR.t1318 VGND 0.00651f
C22156 VPWR.n1544 VGND 0.00179f
C22157 VPWR.t1233 VGND 0.00166f
C22158 VPWR.t1235 VGND 0.00166f
C22159 VPWR.n1545 VGND 0.00345f
C22160 VPWR.t1231 VGND 0.00695f
C22161 VPWR.t3587 VGND 0.00911f
C22162 VPWR.t204 VGND 0.00391f
C22163 VPWR.n1546 VGND 0.0253f
C22164 VPWR.t203 VGND 0.00391f
C22165 VPWR.n1548 VGND 0.0138f
C22166 VPWR.n1549 VGND 0.00345f
C22167 VPWR.t3523 VGND 0.00911f
C22168 VPWR.t518 VGND 0.00391f
C22169 VPWR.n1550 VGND 0.0253f
C22170 VPWR.t519 VGND 0.00391f
C22171 VPWR.n1552 VGND 0.0138f
C22172 VPWR.n1553 VGND 0.011f
C22173 VPWR.n1554 VGND 0.00819f
C22174 VPWR.n1555 VGND 0.00393f
C22175 VPWR.n1556 VGND 0.00333f
C22176 VPWR.n1557 VGND 0.00122f
C22177 VPWR.n1558 VGND 0.00502f
C22178 VPWR.n1559 VGND 0.00393f
C22179 VPWR.n1560 VGND 0.00126f
C22180 VPWR.n1561 VGND 0.00524f
C22181 VPWR.t1229 VGND 0.00225f
C22182 VPWR.t1320 VGND 0.00166f
C22183 VPWR.n1562 VGND 0.00438f
C22184 VPWR.t949 VGND 0.00102f
C22185 VPWR.t3307 VGND 0.00154f
C22186 VPWR.n1563 VGND 0.00483f
C22187 VPWR.n1564 VGND 0.00665f
C22188 VPWR.n1565 VGND 0.00574f
C22189 VPWR.n1566 VGND 9.88e-19
C22190 VPWR.n1567 VGND 0.00524f
C22191 VPWR.n1568 VGND 0.0031f
C22192 VPWR.n1569 VGND 0.00164f
C22193 VPWR.n1570 VGND 0.0082f
C22194 VPWR.n1571 VGND 0.00125f
C22195 VPWR.n1572 VGND 0.00393f
C22196 VPWR.n1573 VGND 0.00393f
C22197 VPWR.t1285 VGND 0.00692f
C22198 VPWR.n1574 VGND 0.0163f
C22199 VPWR.n1575 VGND 6.86e-19
C22200 VPWR.n1576 VGND 0.00393f
C22201 VPWR.t1519 VGND 0.00242f
C22202 VPWR.n1577 VGND 0.00484f
C22203 VPWR.n1578 VGND 8.77e-19
C22204 VPWR.n1579 VGND 0.00333f
C22205 VPWR.n1580 VGND 0.00899f
C22206 VPWR.t2285 VGND 0.00453f
C22207 VPWR.n1581 VGND 0.0116f
C22208 VPWR.n1582 VGND 0.00665f
C22209 VPWR.n1583 VGND 0.0104f
C22210 VPWR.n1584 VGND 0.00688f
C22211 VPWR.n1585 VGND 0.0105f
C22212 VPWR.n1586 VGND 0.0039f
C22213 VPWR.n1587 VGND 0.00351f
C22214 VPWR.n1588 VGND 2.56e-19
C22215 VPWR.n1589 VGND 4.55e-19
C22216 VPWR.n1590 VGND 2.56e-19
C22217 VPWR.t717 VGND 0.00387f
C22218 VPWR.n1591 VGND 0.00508f
C22219 VPWR.n1592 VGND 0.00127f
C22220 VPWR.n1593 VGND 4.48e-19
C22221 VPWR.n1594 VGND 3.13e-19
C22222 VPWR.n1595 VGND 7.4e-19
C22223 VPWR.n1596 VGND 5.41e-19
C22224 VPWR.n1597 VGND 9.96e-19
C22225 VPWR.n1598 VGND 9.68e-19
C22226 VPWR.n1599 VGND 3.7e-19
C22227 VPWR.n1600 VGND 6.83e-19
C22228 VPWR.n1601 VGND 0.00127f
C22229 VPWR.t985 VGND 6.73e-19
C22230 VPWR.t1184 VGND 9.96e-19
C22231 VPWR.n1602 VGND 0.00176f
C22232 VPWR.n1603 VGND 0.00941f
C22233 VPWR.n1604 VGND 0.00321f
C22234 VPWR.n1605 VGND 4.27e-19
C22235 VPWR.n1606 VGND 1.14e-19
C22236 VPWR.n1607 VGND 4.27e-19
C22237 VPWR.n1608 VGND 0.00153f
C22238 VPWR.n1609 VGND 0.00206f
C22239 VPWR.n1610 VGND 0.00138f
C22240 VPWR.n1611 VGND 9e-19
C22241 VPWR.n1612 VGND 6.14e-19
C22242 VPWR.n1613 VGND 9.06e-19
C22243 VPWR.n1614 VGND 5.48e-19
C22244 VPWR.n1615 VGND 0.00138f
C22245 VPWR.n1616 VGND 0.0057f
C22246 VPWR.n1618 VGND 4.11e-19
C22247 VPWR.n1619 VGND 4.11e-19
C22248 VPWR.n1620 VGND 7.39e-19
C22249 VPWR.n1621 VGND 5.19e-19
C22250 VPWR.n1622 VGND 7.39e-19
C22251 VPWR.n1623 VGND 4.11e-19
C22252 VPWR.n1624 VGND 4.11e-19
C22253 VPWR.n1625 VGND 4.61e-19
C22254 VPWR.n1626 VGND 3.73e-19
C22255 VPWR.n1627 VGND 2.41e-19
C22256 VPWR.n1628 VGND 4.83e-19
C22257 VPWR.n1629 VGND 8.26e-19
C22258 VPWR.n1630 VGND 1.99e-19
C22259 VPWR.n1631 VGND 4.84e-19
C22260 VPWR.n1632 VGND 6.83e-19
C22261 VPWR.n1633 VGND 0.00156f
C22262 VPWR.n1634 VGND 4.84e-19
C22263 VPWR.n1635 VGND 5.38e-19
C22264 VPWR.n1636 VGND 4.27e-19
C22265 VPWR.n1637 VGND 4.66e-19
C22266 VPWR.n1638 VGND 4.27e-19
C22267 VPWR.t235 VGND 0.0046f
C22268 VPWR.n1639 VGND 0.00105f
C22269 VPWR.n1640 VGND 0.00309f
C22270 VPWR.n1641 VGND 9.6e-19
C22271 VPWR.n1642 VGND 0.00217f
C22272 VPWR.n1643 VGND 0.00632f
C22273 VPWR.n1644 VGND 0.00451f
C22274 VPWR.n1645 VGND 0.0066f
C22275 VPWR.n1646 VGND 0.00524f
C22276 VPWR.t748 VGND 0.00234f
C22277 VPWR.n1647 VGND 0.00474f
C22278 VPWR.n1648 VGND 0.00398f
C22279 VPWR.n1649 VGND 0.00524f
C22280 VPWR.t3342 VGND 0.0592f
C22281 VPWR.n1650 VGND 0.0349f
C22282 VPWR.n1651 VGND 0.00484f
C22283 VPWR.n1652 VGND 0.00524f
C22284 VPWR.n1653 VGND 0.0066f
C22285 VPWR.n1654 VGND 0.00524f
C22286 VPWR.t1327 VGND 0.00102f
C22287 VPWR.t1023 VGND 0.00102f
C22288 VPWR.n1655 VGND 0.00217f
C22289 VPWR.n1656 VGND 0.0071f
C22290 VPWR.n1657 VGND 0.00337f
C22291 VPWR.n1658 VGND 0.00524f
C22292 VPWR.n1659 VGND 0.0031f
C22293 VPWR.n1660 VGND 0.00199f
C22294 VPWR.n1661 VGND 0.0147f
C22295 VPWR.n1662 VGND 0.0066f
C22296 VPWR.n1663 VGND 0.00393f
C22297 VPWR.t1406 VGND 0.00136f
C22298 VPWR.t1513 VGND 0.00136f
C22299 VPWR.n1664 VGND 0.00317f
C22300 VPWR.n1665 VGND 0.0119f
C22301 VPWR.n1666 VGND 0.00524f
C22302 VPWR.n1667 VGND 0.0031f
C22303 VPWR.n1668 VGND 0.00237f
C22304 VPWR.n1669 VGND 0.00166f
C22305 VPWR.t496 VGND 0.0046f
C22306 VPWR.n1670 VGND 0.00407f
C22307 VPWR.n1671 VGND 0.00122f
C22308 VPWR.n1672 VGND 0.00393f
C22309 VPWR.n1673 VGND 0.00477f
C22310 VPWR.n1674 VGND 0.00524f
C22311 VPWR.t3359 VGND 0.0176f
C22312 VPWR.n1675 VGND 0.00891f
C22313 VPWR.n1676 VGND 0.00228f
C22314 VPWR.t43 VGND 0.00387f
C22315 VPWR.n1677 VGND 0.00634f
C22316 VPWR.n1678 VGND 0.0109f
C22317 VPWR.t44 VGND 0.00432f
C22318 VPWR.n1679 VGND 0.0318f
C22319 VPWR.n1680 VGND 0.00492f
C22320 VPWR.n1681 VGND 0.00524f
C22321 VPWR.n1682 VGND 0.0031f
C22322 VPWR.n1683 VGND 0.0055f
C22323 VPWR.t3433 VGND 0.0597f
C22324 VPWR.n1684 VGND 0.034f
C22325 VPWR.t319 VGND 0.0046f
C22326 VPWR.n1685 VGND 0.011f
C22327 VPWR.n1686 VGND 0.00644f
C22328 VPWR.n1687 VGND 0.00396f
C22329 VPWR.n1688 VGND 0.00393f
C22330 VPWR.n1689 VGND 0.00524f
C22331 VPWR.n1690 VGND 0.0113f
C22332 VPWR.n1691 VGND 0.00524f
C22333 VPWR.n1692 VGND 0.0087f
C22334 VPWR.n1693 VGND 0.00524f
C22335 VPWR.t3449 VGND 0.0592f
C22336 VPWR.n1694 VGND 0.038f
C22337 VPWR.n1695 VGND 0.00833f
C22338 VPWR.n1696 VGND 0.00524f
C22339 VPWR.n1697 VGND 0.0113f
C22340 VPWR.n1698 VGND 0.00524f
C22341 VPWR.n1699 VGND 0.011f
C22342 VPWR.n1700 VGND 0.00524f
C22343 VPWR.n1701 VGND 0.0031f
C22344 VPWR.n1702 VGND 0.00535f
C22345 VPWR.t2602 VGND 0.00633f
C22346 VPWR.n1703 VGND 0.0121f
C22347 VPWR.n1704 VGND 0.00333f
C22348 VPWR.n1705 VGND 0.00475f
C22349 VPWR.n1706 VGND 0.00639f
C22350 VPWR.n1707 VGND 0.00524f
C22351 VPWR.n1708 VGND 0.00307f
C22352 VPWR.n1709 VGND 0.00639f
C22353 VPWR.t320 VGND 0.0046f
C22354 VPWR.n1710 VGND 0.00407f
C22355 VPWR.n1711 VGND 0.00228f
C22356 VPWR.n1712 VGND 0.00179f
C22357 VPWR.n1713 VGND 0.00262f
C22358 VPWR.n1714 VGND 0.00612f
C22359 VPWR.n1715 VGND 0.0074f
C22360 VPWR.n1716 VGND 0.00619f
C22361 VPWR.n1717 VGND 0.00393f
C22362 VPWR.n1718 VGND 0.00393f
C22363 VPWR.n1719 VGND 0.00524f
C22364 VPWR.n1720 VGND 0.0031f
C22365 VPWR.n1721 VGND 0.0138f
C22366 VPWR.n1722 VGND 0.0138f
C22367 VPWR.n1723 VGND 0.0133f
C22368 VPWR.n1724 VGND 0.00333f
C22369 VPWR.t1895 VGND 0.00166f
C22370 VPWR.t1623 VGND 0.00184f
C22371 VPWR.n1725 VGND 0.00362f
C22372 VPWR.n1726 VGND 0.00393f
C22373 VPWR.t2143 VGND 0.00561f
C22374 VPWR.n1727 VGND 0.00744f
C22375 VPWR.n1728 VGND 5.69e-19
C22376 VPWR.n1729 VGND 0.00131f
C22377 VPWR.n1730 VGND 9.96e-19
C22378 VPWR.n1731 VGND 4.27e-19
C22379 VPWR.n1732 VGND 5.12e-19
C22380 VPWR.n1733 VGND 5.41e-19
C22381 VPWR.n1734 VGND 7.76e-19
C22382 VPWR.n1735 VGND 5.41e-19
C22383 VPWR.n1736 VGND 1.31e-19
C22384 VPWR.n1737 VGND 3.7e-19
C22385 VPWR.n1738 VGND 1.21e-19
C22386 VPWR.n1739 VGND 3.42e-19
C22387 VPWR.n1740 VGND 4.74e-19
C22388 VPWR.n1741 VGND 3.7e-19
C22389 VPWR.n1742 VGND 6.26e-19
C22390 VPWR.n1743 VGND 6.55e-19
C22391 VPWR.n1744 VGND 5.41e-19
C22392 VPWR.n1745 VGND 9.96e-19
C22393 VPWR.n1746 VGND 9.68e-19
C22394 VPWR.n1747 VGND 5.41e-19
C22395 VPWR.n1748 VGND 3.13e-19
C22396 VPWR.n1749 VGND 5.98e-19
C22397 VPWR.n1750 VGND 5.12e-19
C22398 VPWR.n1751 VGND 7.12e-19
C22399 VPWR.n1752 VGND 5.98e-19
C22400 VPWR.n1753 VGND 8.11e-19
C22401 VPWR.n1754 VGND 3.95e-19
C22402 VPWR.n1755 VGND 3.95e-19
C22403 VPWR.n1756 VGND 7.68e-19
C22404 VPWR.n1757 VGND 5.05e-19
C22405 VPWR.n1758 VGND 0.00139f
C22406 VPWR.n1759 VGND 9.06e-19
C22407 VPWR.n1760 VGND 5.48e-19
C22408 VPWR.n1761 VGND 1.76e-19
C22409 VPWR.n1762 VGND 1.76e-19
C22410 VPWR.n1763 VGND 3.13e-19
C22411 VPWR.n1764 VGND 5.12e-19
C22412 VPWR.n1765 VGND 6.26e-19
C22413 VPWR.t769 VGND 0.0042f
C22414 VPWR.n1766 VGND 0.00704f
C22415 VPWR.n1767 VGND 4.61e-20
C22416 VPWR.n1768 VGND 4.67e-19
C22417 VPWR.n1769 VGND 0.00259f
C22418 VPWR.n1770 VGND 0.00495f
C22419 VPWR.n1771 VGND 0.00127f
C22420 VPWR.n1772 VGND 0.00473f
C22421 VPWR.n1773 VGND 0.00179f
C22422 VPWR.n1774 VGND 0.00179f
C22423 VPWR.n1775 VGND 0.0129f
C22424 VPWR.n1776 VGND 0.0188f
C22425 VPWR.t2252 VGND 0.00571f
C22426 VPWR.t2405 VGND 0.0121f
C22427 VPWR.t744 VGND 0.0144f
C22428 VPWR.t1894 VGND 0.018f
C22429 VPWR.t1622 VGND 0.0151f
C22430 VPWR.t768 VGND 0.0344f
C22431 VPWR.t2171 VGND 0.0346f
C22432 VPWR.t2142 VGND 0.0141f
C22433 VPWR.t2174 VGND 0.0144f
C22434 VPWR.t2148 VGND 0.0141f
C22435 VPWR.t2234 VGND 0.0144f
C22436 VPWR.t2150 VGND 0.0141f
C22437 VPWR.t2240 VGND 0.0144f
C22438 VPWR.t2140 VGND 0.0114f
C22439 VPWR.t2146 VGND 0.0188f
C22440 VPWR.t2136 VGND 0.0238f
C22441 VPWR.t172 VGND 0.0144f
C22442 VPWR.t2138 VGND 0.0183f
C22443 VPWR.t2144 VGND 0.0153f
C22444 VPWR.t2154 VGND 0.00604f
C22445 VPWR.t2642 VGND 0.0144f
C22446 VPWR.t2124 VGND 0.0141f
C22447 VPWR.t2352 VGND 0.0144f
C22448 VPWR.t2152 VGND 0.0233f
C22449 VPWR.t2132 VGND 0.0232f
C22450 VPWR.t1236 VGND 0.0144f
C22451 VPWR.t2126 VGND 0.0156f
C22452 VPWR.t2175 VGND 0.0144f
C22453 VPWR.t2128 VGND 0.0161f
C22454 VPWR.t2599 VGND 0.0144f
C22455 VPWR.t2130 VGND 0.0173f
C22456 VPWR.t2134 VGND 0.0287f
C22457 VPWR.t1725 VGND 0.0144f
C22458 VPWR.t1063 VGND 0.0141f
C22459 VPWR.t3017 VGND 0.0144f
C22460 VPWR.t1055 VGND 0.0141f
C22461 VPWR.t772 VGND 0.0144f
C22462 VPWR.t1057 VGND 0.0107f
C22463 VPWR.t1061 VGND 0.0128f
C22464 VPWR.t2329 VGND 0.0196f
C22465 VPWR.t2324 VGND 0.0255f
C22466 VPWR.t2757 VGND 0.0124f
C22467 VPWR.n1777 VGND 0.0218f
C22468 VPWR.t2758 VGND 0.00108f
C22469 VPWR.t2321 VGND 0.0028f
C22470 VPWR.n1778 VGND 0.00485f
C22471 VPWR.n1779 VGND 0.00641f
C22472 VPWR.t2328 VGND 0.0016f
C22473 VPWR.t2619 VGND 0.0016f
C22474 VPWR.n1780 VGND 0.00331f
C22475 VPWR.t2916 VGND 0.00136f
C22476 VPWR.t1032 VGND 0.00136f
C22477 VPWR.n1781 VGND 0.00328f
C22478 VPWR.n1782 VGND 0.00965f
C22479 VPWR.t1611 VGND 0.00532f
C22480 VPWR.n1783 VGND 0.0053f
C22481 VPWR.t2611 VGND 0.00532f
C22482 VPWR.t2861 VGND 0.00654f
C22483 VPWR.n1784 VGND 0.0106f
C22484 VPWR.t1613 VGND 0.00531f
C22485 VPWR.n1785 VGND 0.00619f
C22486 VPWR.t2613 VGND 0.0016f
C22487 VPWR.t2621 VGND 0.0016f
C22488 VPWR.n1786 VGND 0.0037f
C22489 VPWR.t244 VGND 0.0046f
C22490 VPWR.n1787 VGND 0.004f
C22491 VPWR.n1788 VGND 0.0039f
C22492 VPWR.n1789 VGND 0.00137f
C22493 VPWR.n1790 VGND 4.66e-19
C22494 VPWR.n1791 VGND 3.7e-19
C22495 VPWR.n1792 VGND 3.23e-19
C22496 VPWR.n1793 VGND 3.7e-19
C22497 VPWR.t245 VGND 0.0046f
C22498 VPWR.n1794 VGND 0.00113f
C22499 VPWR.n1795 VGND 0.00309f
C22500 VPWR.n1796 VGND 5.12e-19
C22501 VPWR.n1797 VGND 5.71e-19
C22502 VPWR.n1798 VGND 3.29e-19
C22503 VPWR.n1799 VGND 3.95e-19
C22504 VPWR.n1800 VGND 3.95e-19
C22505 VPWR.n1801 VGND 6.54e-19
C22506 VPWR.n1802 VGND 8.67e-19
C22507 VPWR.n1803 VGND 0.1f
C22508 VPWR.n1804 VGND 0.0839f
C22509 VPWR.n1805 VGND 0.59f
C22510 VPWR.n1806 VGND 0.0057f
C22511 VPWR.n1807 VGND 6.54e-19
C22512 VPWR.n1808 VGND 8.67e-19
C22513 VPWR.n1809 VGND 3.95e-19
C22514 VPWR.n1810 VGND 4.61e-19
C22515 VPWR.n1811 VGND 2.41e-19
C22516 VPWR.n1812 VGND 0.00143f
C22517 VPWR.n1813 VGND 3.13e-19
C22518 VPWR.t1529 VGND 0.0016f
C22519 VPWR.t1859 VGND 0.00225f
C22520 VPWR.n1814 VGND 0.00444f
C22521 VPWR.n1815 VGND 0.00764f
C22522 VPWR.t757 VGND 0.0016f
C22523 VPWR.t752 VGND 0.0016f
C22524 VPWR.n1816 VGND 0.00377f
C22525 VPWR.n1817 VGND 0.00627f
C22526 VPWR.n1818 VGND 3.29e-19
C22527 VPWR.n1819 VGND 5.71e-19
C22528 VPWR.n1820 VGND 5.92e-19
C22529 VPWR.n1821 VGND 5.05e-19
C22530 VPWR.n1822 VGND 8.67e-19
C22531 VPWR.n1823 VGND 6.54e-19
C22532 VPWR.n1824 VGND 9.06e-19
C22533 VPWR.n1825 VGND 0.00138f
C22534 VPWR.n1826 VGND 5.48e-19
C22535 VPWR.n1827 VGND 4.17e-19
C22536 VPWR.n1828 VGND 0.00138f
C22537 VPWR.t755 VGND 0.0016f
C22538 VPWR.t750 VGND 0.0016f
C22539 VPWR.n1829 VGND 0.00379f
C22540 VPWR.n1830 VGND 0.00819f
C22541 VPWR.t1158 VGND 0.0016f
C22542 VPWR.t1162 VGND 0.0016f
C22543 VPWR.n1831 VGND 0.00371f
C22544 VPWR.n1832 VGND 0.00765f
C22545 VPWR.n1833 VGND 0.00445f
C22546 VPWR.t85 VGND 0.004f
C22547 VPWR.n1834 VGND 0.00182f
C22548 VPWR.t3548 VGND 0.00916f
C22549 VPWR.t84 VGND 0.00391f
C22550 VPWR.n1835 VGND 0.018f
C22551 VPWR.n1836 VGND 0.0104f
C22552 VPWR.n1837 VGND 0.00764f
C22553 VPWR.n1838 VGND 0.00262f
C22554 VPWR.t1160 VGND 0.00591f
C22555 VPWR.t648 VGND 0.00387f
C22556 VPWR.n1839 VGND 0.00837f
C22557 VPWR.t1714 VGND 0.00632f
C22558 VPWR.n1840 VGND 0.00123f
C22559 VPWR.t2762 VGND 0.00239f
C22560 VPWR.t3436 VGND 0.00911f
C22561 VPWR.t484 VGND 0.00391f
C22562 VPWR.n1841 VGND 0.0253f
C22563 VPWR.t485 VGND 0.00391f
C22564 VPWR.n1843 VGND 0.0138f
C22565 VPWR.t1511 VGND 6.73e-19
C22566 VPWR.t3012 VGND 6.73e-19
C22567 VPWR.n1844 VGND 0.00157f
C22568 VPWR.t1900 VGND 9.96e-19
C22569 VPWR.t2009 VGND 4.13e-19
C22570 VPWR.n1845 VGND 0.00507f
C22571 VPWR.n1846 VGND 0.0116f
C22572 VPWR.n1847 VGND 0.024f
C22573 VPWR.n1848 VGND 0.00123f
C22574 VPWR.t1949 VGND 0.00598f
C22575 VPWR.n1849 VGND 0.00834f
C22576 VPWR.t3279 VGND 0.00663f
C22577 VPWR.n1850 VGND 0.00878f
C22578 VPWR.t1491 VGND 0.00597f
C22579 VPWR.n1851 VGND 0.00154f
C22580 VPWR.t856 VGND 0.0016f
C22581 VPWR.t854 VGND 0.0016f
C22582 VPWR.n1852 VGND 0.00379f
C22583 VPWR.n1853 VGND 0.0078f
C22584 VPWR.n1854 VGND 0.00137f
C22585 VPWR.t852 VGND 0.00654f
C22586 VPWR.n1855 VGND 0.0106f
C22587 VPWR.n1856 VGND 5.41e-19
C22588 VPWR.n1857 VGND 5.71e-19
C22589 VPWR.n1858 VGND 3.29e-19
C22590 VPWR.n1859 VGND 3.95e-19
C22591 VPWR.n1860 VGND 4.17e-19
C22592 VPWR.n1861 VGND 2.85e-19
C22593 VPWR.n1862 VGND 6.54e-19
C22594 VPWR.n1863 VGND 8.67e-19
C22595 VPWR.n1864 VGND 0.00139f
C22596 VPWR.n1865 VGND 9.06e-19
C22597 VPWR.n1866 VGND 5.92e-19
C22598 VPWR.n1867 VGND 5.05e-19
C22599 VPWR.n1868 VGND 4.17e-19
C22600 VPWR.n1869 VGND 5.48e-19
C22601 VPWR.n1871 VGND 8.67e-19
C22602 VPWR.n1872 VGND 6.54e-19
C22603 VPWR.n1873 VGND 9.06e-19
C22604 VPWR.n1874 VGND 5.05e-19
C22605 VPWR.n1875 VGND 8.11e-19
C22606 VPWR.n1876 VGND 3.95e-19
C22607 VPWR.n1877 VGND 9.96e-19
C22608 VPWR.n1878 VGND 9.68e-19
C22609 VPWR.n1879 VGND 5.12e-19
C22610 VPWR.n1880 VGND 0.00166f
C22611 VPWR.n1881 VGND 3.13e-19
C22612 VPWR.n1882 VGND 6.26e-19
C22613 VPWR.n1883 VGND 5.12e-19
C22614 VPWR.n1884 VGND 3.95e-19
C22615 VPWR.n1885 VGND 7.68e-19
C22616 VPWR.n1886 VGND 3.95e-19
C22617 VPWR.n1887 VGND 6.26e-19
C22618 VPWR.t1279 VGND 0.00483f
C22619 VPWR.t2318 VGND 0.0048f
C22620 VPWR.n1888 VGND 0.00698f
C22621 VPWR.n1889 VGND 0.0129f
C22622 VPWR.t1402 VGND 0.00586f
C22623 VPWR.t3330 VGND 0.00529f
C22624 VPWR.n1890 VGND 0.00489f
C22625 VPWR.t3332 VGND 0.00219f
C22626 VPWR.t3122 VGND 0.00166f
C22627 VPWR.n1891 VGND 0.00445f
C22628 VPWR.n1892 VGND 0.00774f
C22629 VPWR.t1510 VGND 0.0218f
C22630 VPWR.t3011 VGND 0.0232f
C22631 VPWR.t483 VGND 0.0159f
C22632 VPWR.t1899 VGND 0.0183f
C22633 VPWR.t2008 VGND 0.0154f
C22634 VPWR.t1948 VGND 0.0151f
C22635 VPWR.t3278 VGND 0.022f
C22636 VPWR.t2603 VGND 0.0141f
C22637 VPWR.t3280 VGND 0.0143f
C22638 VPWR.t1191 VGND 0.0154f
C22639 VPWR.t1121 VGND 0.0149f
C22640 VPWR.t1986 VGND 0.0114f
C22641 VPWR.t1119 VGND 0.0359f
C22642 VPWR.t2010 VGND 0.0334f
C22643 VPWR.t1115 VGND 0.0451f
C22644 VPWR.t1737 VGND 0.0386f
C22645 VPWR.t1033 VGND 0.00571f
C22646 VPWR.t855 VGND 0.0121f
C22647 VPWR.t851 VGND 0.0141f
C22648 VPWR.t853 VGND 0.0168f
C22649 VPWR.t1750 VGND 0.0282f
C22650 VPWR.t1749 VGND 0.0279f
C22651 VPWR.t1278 VGND 0.0156f
C22652 VPWR.t2317 VGND 0.0232f
C22653 VPWR.t1728 VGND 0.018f
C22654 VPWR.t2227 VGND 0.0123f
C22655 VPWR.t1730 VGND 0.0107f
C22656 VPWR.t1401 VGND 0.0208f
C22657 VPWR.t3329 VGND 0.0235f
C22658 VPWR.t1741 VGND 0.00109f
C22659 VPWR.t3039 VGND 5.47e-19
C22660 VPWR.n1893 VGND 0.0069f
C22661 VPWR.n1894 VGND 0.0071f
C22662 VPWR.n1895 VGND 0.0127f
C22663 VPWR.n1896 VGND 0.0131f
C22664 VPWR.t614 VGND 0.00387f
C22665 VPWR.n1897 VGND 0.00837f
C22666 VPWR.n1898 VGND 0.00513f
C22667 VPWR.n1899 VGND 0.00129f
C22668 VPWR.t1044 VGND 0.00131f
C22669 VPWR.t1394 VGND 4.27e-19
C22670 VPWR.n1900 VGND 0.00672f
C22671 VPWR.t2865 VGND 0.0067f
C22672 VPWR.n1901 VGND 0.0151f
C22673 VPWR.t3475 VGND 0.0289f
C22674 VPWR.t613 VGND 0.00387f
C22675 VPWR.n1902 VGND 0.0604f
C22676 VPWR.n1903 VGND 0.0146f
C22677 VPWR.n1904 VGND 0.0117f
C22678 VPWR.t3498 VGND 0.00911f
C22679 VPWR.t698 VGND 0.00391f
C22680 VPWR.n1905 VGND 0.0253f
C22681 VPWR.t697 VGND 0.00391f
C22682 VPWR.n1907 VGND 0.0138f
C22683 VPWR.n1908 VGND 0.00376f
C22684 VPWR.n1909 VGND 0.00182f
C22685 VPWR.t1458 VGND 0.0016f
C22686 VPWR.t3291 VGND 0.0016f
C22687 VPWR.n1910 VGND 0.00376f
C22688 VPWR.t1456 VGND 0.00634f
C22689 VPWR.n1911 VGND 0.00899f
C22690 VPWR.t2945 VGND 0.00631f
C22691 VPWR.n1912 VGND 0.00177f
C22692 VPWR.n1913 VGND 0.00152f
C22693 VPWR.n1914 VGND 0.00179f
C22694 VPWR.n1915 VGND 0.00186f
C22695 VPWR.n1916 VGND 0.00172f
C22696 VPWR.n1917 VGND 0.00475f
C22697 VPWR.t1404 VGND 0.00225f
C22698 VPWR.t2943 VGND 0.00225f
C22699 VPWR.n1918 VGND 0.00514f
C22700 VPWR.n1919 VGND 0.00635f
C22701 VPWR.n1920 VGND 0.00524f
C22702 VPWR.t3008 VGND 0.00527f
C22703 VPWR.n1921 VGND 0.00595f
C22704 VPWR.n1922 VGND 0.00524f
C22705 VPWR.t2947 VGND 0.0016f
C22706 VPWR.t2941 VGND 0.0016f
C22707 VPWR.n1923 VGND 0.00383f
C22708 VPWR.n1924 VGND 0.00621f
C22709 VPWR.n1925 VGND 0.00524f
C22710 VPWR.n1926 VGND 0.00524f
C22711 VPWR.n1927 VGND 0.00393f
C22712 VPWR.t2229 VGND 0.00208f
C22713 VPWR.t2930 VGND 0.0016f
C22714 VPWR.n1928 VGND 0.00422f
C22715 VPWR.n1929 VGND 0.00578f
C22716 VPWR.n1930 VGND 0.0068f
C22717 VPWR.n1931 VGND 0.00892f
C22718 VPWR.n1932 VGND 0.00112f
C22719 VPWR.n1933 VGND 0.00393f
C22720 VPWR.t3297 VGND 0.0016f
C22721 VPWR.t3295 VGND 0.0016f
C22722 VPWR.n1934 VGND 0.00367f
C22723 VPWR.n1935 VGND 0.00626f
C22724 VPWR.n1936 VGND 0.00119f
C22725 VPWR.n1937 VGND 0.00524f
C22726 VPWR.t1042 VGND 7.22e-19
C22727 VPWR.t2064 VGND 9.22e-19
C22728 VPWR.n1938 VGND 0.00189f
C22729 VPWR.n1939 VGND 0.00348f
C22730 VPWR.n1940 VGND 0.00116f
C22731 VPWR.n1941 VGND 0.00524f
C22732 VPWR.t3289 VGND 0.0016f
C22733 VPWR.t3293 VGND 0.0016f
C22734 VPWR.n1942 VGND 0.00379f
C22735 VPWR.n1943 VGND 0.00819f
C22736 VPWR.n1944 VGND 0.00524f
C22737 VPWR.n1945 VGND 0.00103f
C22738 VPWR.n1946 VGND 0.00524f
C22739 VPWR.t3299 VGND 0.00655f
C22740 VPWR.n1947 VGND 0.0111f
C22741 VPWR.n1948 VGND 0.00393f
C22742 VPWR.n1949 VGND 0.00199f
C22743 VPWR.n1950 VGND 0.00275f
C22744 VPWR.n1951 VGND 0.00996f
C22745 VPWR.n1952 VGND 0.00545f
C22746 VPWR.n1953 VGND 0.0113f
C22747 VPWR.n1954 VGND 0.00699f
C22748 VPWR.n1955 VGND 0.00524f
C22749 VPWR.n1956 VGND 0.00524f
C22750 VPWR.n1957 VGND 0.0031f
C22751 VPWR.n1958 VGND 0.00199f
C22752 VPWR.t401 VGND 0.00387f
C22753 VPWR.t3396 VGND 0.0231f
C22754 VPWR.n1959 VGND 0.0138f
C22755 VPWR.n1960 VGND 0.00393f
C22756 VPWR.t2060 VGND 0.00136f
C22757 VPWR.t2872 VGND 0.00136f
C22758 VPWR.n1961 VGND 0.00317f
C22759 VPWR.n1962 VGND 0.0188f
C22760 VPWR.t402 VGND 0.00387f
C22761 VPWR.n1963 VGND 0.00837f
C22762 VPWR.t2979 VGND 0.00676f
C22763 VPWR.t1218 VGND 0.00239f
C22764 VPWR.n1964 VGND 0.0136f
C22765 VPWR.n1965 VGND 7.88e-19
C22766 VPWR.n1966 VGND 3.95e-19
C22767 VPWR.n1967 VGND 5.05e-19
C22768 VPWR.n1968 VGND 5.05e-19
C22769 VPWR.n1969 VGND 0.00139f
C22770 VPWR.n1970 VGND 9.06e-19
C22771 VPWR.n1971 VGND 9e-19
C22772 VPWR.n1972 VGND 0.00138f
C22773 VPWR.n1973 VGND 6.14e-19
C22774 VPWR.n1974 VGND 5.48e-19
C22775 VPWR.n1975 VGND 0.00138f
C22776 VPWR.n1976 VGND 0.0994f
C22777 VPWR.n1977 VGND 7.39e-19
C22778 VPWR.n1978 VGND 4.11e-19
C22779 VPWR.n1979 VGND 6.54e-19
C22780 VPWR.n1980 VGND 8.67e-19
C22781 VPWR.n1981 VGND 4.17e-19
C22782 VPWR.n1982 VGND 3.51e-19
C22783 VPWR.n1983 VGND 4.61e-19
C22784 VPWR.n1984 VGND 4.39e-19
C22785 VPWR.n1985 VGND 3.29e-19
C22786 VPWR.n1986 VGND 5.27e-19
C22787 VPWR.n1987 VGND 2.85e-19
C22788 VPWR.n1988 VGND 2.85e-19
C22789 VPWR.n1989 VGND 4.17e-19
C22790 VPWR.n1990 VGND 4.11e-19
C22791 VPWR.t2467 VGND 0.00235f
C22792 VPWR.n1992 VGND 0.00665f
C22793 VPWR.n1993 VGND 0.00127f
C22794 VPWR.n1994 VGND 0.00441f
C22795 VPWR.t3373 VGND 0.0289f
C22796 VPWR.t313 VGND 0.00387f
C22797 VPWR.n1995 VGND 0.0604f
C22798 VPWR.n1996 VGND 0.0135f
C22799 VPWR.n1997 VGND 0.0117f
C22800 VPWR.n1998 VGND 0.0146f
C22801 VPWR.t2510 VGND 6.73e-19
C22802 VPWR.t2021 VGND 9.96e-19
C22803 VPWR.n1999 VGND 0.00176f
C22804 VPWR.t448 VGND 0.0463f
C22805 VPWR.t3176 VGND 0.0124f
C22806 VPWR.t2191 VGND 0.0148f
C22807 VPWR.t2030 VGND 0.0144f
C22808 VPWR.t2189 VGND 0.0156f
C22809 VPWR.t2195 VGND 0.0195f
C22810 VPWR.t2193 VGND 0.0255f
C22811 VPWR.t2335 VGND 0.0215f
C22812 VPWR.t1673 VGND 0.0411f
C22813 VPWR.t1755 VGND 0.02f
C22814 VPWR.t101 VGND 0.0154f
C22815 VPWR.t163 VGND 0.0926f
C22816 VPWR.t1775 VGND 0.025f
C22817 VPWR.t1945 VGND 0.0305f
C22818 VPWR.t312 VGND 0.0448f
C22819 VPWR.t2466 VGND 0.0438f
C22820 VPWR.t1506 VGND 0.0321f
C22821 VPWR.t1944 VGND 0.0227f
C22822 VPWR.t2020 VGND 0.0337f
C22823 VPWR.t2509 VGND 0.0164f
C22824 VPWR.n2000 VGND 0.0162f
C22825 VPWR.t1810 VGND 0.00453f
C22826 VPWR.n2001 VGND 0.0138f
C22827 VPWR.n2002 VGND 0.00912f
C22828 VPWR.n2003 VGND 0.0111f
C22829 VPWR.t381 VGND 0.00387f
C22830 VPWR.n2004 VGND 0.00613f
C22831 VPWR.n2005 VGND 0.00525f
C22832 VPWR.t1786 VGND 0.00239f
C22833 VPWR.n2006 VGND 0.00421f
C22834 VPWR.t1241 VGND 0.0016f
C22835 VPWR.t1247 VGND 0.0016f
C22836 VPWR.n2007 VGND 0.00368f
C22837 VPWR.t1243 VGND 0.00655f
C22838 VPWR.n2008 VGND 0.0108f
C22839 VPWR.t860 VGND 0.00624f
C22840 VPWR.n2009 VGND 0.0159f
C22841 VPWR.t3503 VGND 0.00911f
C22842 VPWR.t527 VGND 0.00391f
C22843 VPWR.n2010 VGND 0.0253f
C22844 VPWR.t526 VGND 0.00391f
C22845 VPWR.n2012 VGND 0.0138f
C22846 VPWR.t3486 VGND 0.00911f
C22847 VPWR.t629 VGND 0.00391f
C22848 VPWR.n2013 VGND 0.0253f
C22849 VPWR.t630 VGND 0.00391f
C22850 VPWR.n2015 VGND 0.0138f
C22851 VPWR.n2016 VGND 0.00888f
C22852 VPWR.t1983 VGND 0.00631f
C22853 VPWR.t3527 VGND 0.0179f
C22854 VPWR.n2017 VGND 0.0195f
C22855 VPWR.n2018 VGND 0.0139f
C22856 VPWR.n2019 VGND 0.0179f
C22857 VPWR.t357 VGND 0.0046f
C22858 VPWR.t611 VGND 0.00387f
C22859 VPWR.n2020 VGND 0.0115f
C22860 VPWR.n2021 VGND 0.00681f
C22861 VPWR.n2022 VGND 0.0066f
C22862 VPWR.n2023 VGND 0.00392f
C22863 VPWR.t3364 VGND 0.00911f
C22864 VPWR.t280 VGND 0.00391f
C22865 VPWR.n2024 VGND 0.0253f
C22866 VPWR.t281 VGND 0.00391f
C22867 VPWR.n2026 VGND 0.0138f
C22868 VPWR.t2623 VGND 6.73e-19
C22869 VPWR.t2495 VGND 0.00102f
C22870 VPWR.n2027 VGND 0.0018f
C22871 VPWR.t3539 VGND 0.00911f
C22872 VPWR.t52 VGND 0.00391f
C22873 VPWR.n2028 VGND 0.0253f
C22874 VPWR.t53 VGND 0.00391f
C22875 VPWR.n2030 VGND 0.0138f
C22876 VPWR.n2031 VGND 0.0125f
C22877 VPWR.n2032 VGND 0.00199f
C22878 VPWR.t1569 VGND 0.0124f
C22879 VPWR.t1572 VGND 0.00166f
C22880 VPWR.t1568 VGND 0.00166f
C22881 VPWR.n2033 VGND 0.00345f
C22882 VPWR.n2034 VGND 0.00438f
C22883 VPWR.t1570 VGND 0.00695f
C22884 VPWR.n2035 VGND 0.00819f
C22885 VPWR.t3037 VGND 0.00692f
C22886 VPWR.n2036 VGND 0.0106f
C22887 VPWR.n2037 VGND 3.95e-19
C22888 VPWR.n2038 VGND 7.68e-19
C22889 VPWR.n2039 VGND 5.05e-19
C22890 VPWR.n2040 VGND 1.76e-19
C22891 VPWR.n2041 VGND 2.28e-19
C22892 VPWR.t2465 VGND 0.00166f
C22893 VPWR.t1080 VGND 0.00166f
C22894 VPWR.n2042 VGND 0.00389f
C22895 VPWR.n2043 VGND 0.00538f
C22896 VPWR.n2044 VGND 0.00113f
C22897 VPWR.n2045 VGND 0.00379f
C22898 VPWR.n2046 VGND 0.00179f
C22899 VPWR.t1078 VGND 0.00602f
C22900 VPWR.t266 VGND 0.00387f
C22901 VPWR.n2047 VGND 0.00822f
C22902 VPWR.n2048 VGND 0.00638f
C22903 VPWR.n2049 VGND 0.00457f
C22904 VPWR.n2050 VGND 0.0031f
C22905 VPWR.n2051 VGND 0.00524f
C22906 VPWR.n2052 VGND 0.00524f
C22907 VPWR.t265 VGND 0.00387f
C22908 VPWR.t3412 VGND 0.0179f
C22909 VPWR.t1072 VGND 0.00166f
C22910 VPWR.t1076 VGND 0.00166f
C22911 VPWR.n2053 VGND 0.00379f
C22912 VPWR.n2054 VGND 0.0129f
C22913 VPWR.n2055 VGND 0.0114f
C22914 VPWR.n2056 VGND 0.00389f
C22915 VPWR.n2057 VGND 0.0173f
C22916 VPWR.n2058 VGND 0.00493f
C22917 VPWR.n2059 VGND 0.00457f
C22918 VPWR.n2060 VGND 0.00393f
C22919 VPWR.n2061 VGND 0.0031f
C22920 VPWR.t2689 VGND 0.00102f
C22921 VPWR.t1013 VGND 0.00102f
C22922 VPWR.n2062 VGND 0.00221f
C22923 VPWR.n2063 VGND 0.00124f
C22924 VPWR.n2064 VGND 0.00444f
C22925 VPWR.n2065 VGND 0.00524f
C22926 VPWR.t2459 VGND 0.00166f
C22927 VPWR.t2461 VGND 0.00166f
C22928 VPWR.n2066 VGND 0.00359f
C22929 VPWR.n2067 VGND 0.00538f
C22930 VPWR.n2068 VGND 9.96e-19
C22931 VPWR.n2069 VGND 0.00524f
C22932 VPWR.n2070 VGND 0.00147f
C22933 VPWR.n2071 VGND 0.00524f
C22934 VPWR.t1877 VGND 0.00234f
C22935 VPWR.t2463 VGND 0.00166f
C22936 VPWR.t2457 VGND 0.00166f
C22937 VPWR.n2072 VGND 0.00353f
C22938 VPWR.n2073 VGND 0.00502f
C22939 VPWR.n2074 VGND 0.00342f
C22940 VPWR.n2075 VGND 0.00115f
C22941 VPWR.n2076 VGND 0.00524f
C22942 VPWR.t2455 VGND 0.00166f
C22943 VPWR.t2451 VGND 0.00166f
C22944 VPWR.n2077 VGND 0.00359f
C22945 VPWR.n2078 VGND 0.0057f
C22946 VPWR.n2079 VGND 0.00108f
C22947 VPWR.n2080 VGND 0.00524f
C22948 VPWR.n2081 VGND 0.00125f
C22949 VPWR.n2082 VGND 0.00524f
C22950 VPWR.t2443 VGND 0.0016f
C22951 VPWR.t2453 VGND 0.00166f
C22952 VPWR.n2083 VGND 0.00353f
C22953 VPWR.n2084 VGND 0.00634f
C22954 VPWR.n2085 VGND 0.00527f
C22955 VPWR.n2086 VGND 9.54e-19
C22956 VPWR.n2087 VGND 0.00524f
C22957 VPWR.t2435 VGND 0.00166f
C22958 VPWR.t2437 VGND 0.00166f
C22959 VPWR.n2088 VGND 0.00353f
C22960 VPWR.n2089 VGND 0.00496f
C22961 VPWR.t995 VGND 6.73e-19
C22962 VPWR.t1736 VGND 9.96e-19
C22963 VPWR.n2090 VGND 0.00176f
C22964 VPWR.n2091 VGND 0.00423f
C22965 VPWR.n2092 VGND 5.71e-19
C22966 VPWR.n2093 VGND 0.00524f
C22967 VPWR.n2094 VGND 0.00147f
C22968 VPWR.n2095 VGND 0.00524f
C22969 VPWR.t2439 VGND 0.00166f
C22970 VPWR.t2445 VGND 0.00166f
C22971 VPWR.n2096 VGND 0.00353f
C22972 VPWR.t2653 VGND 0.00453f
C22973 VPWR.n2097 VGND 0.00565f
C22974 VPWR.n2098 VGND 0.00527f
C22975 VPWR.n2099 VGND 0.00524f
C22976 VPWR.n2100 VGND 0.00154f
C22977 VPWR.n2101 VGND 0.00503f
C22978 VPWR.n2102 VGND 3.29e-19
C22979 VPWR.n2103 VGND 5.71e-19
C22980 VPWR.n2104 VGND 5.92e-19
C22981 VPWR.n2105 VGND 5.05e-19
C22982 VPWR.n2106 VGND 8.67e-19
C22983 VPWR.n2107 VGND 6.54e-19
C22984 VPWR.n2108 VGND 9.06e-19
C22985 VPWR.n2109 VGND 0.00139f
C22986 VPWR.n2110 VGND 9.06e-19
C22987 VPWR.n2111 VGND 8.11e-19
C22988 VPWR.n2112 VGND 3.95e-19
C22989 VPWR.t847 VGND 0.00102f
C22990 VPWR.t2910 VGND 0.00154f
C22991 VPWR.n2113 VGND 0.00483f
C22992 VPWR.n2114 VGND 0.00671f
C22993 VPWR.n2115 VGND 0.00433f
C22994 VPWR.t539 VGND 0.046f
C22995 VPWR.t1211 VGND 0.0154f
C22996 VPWR.t1213 VGND 0.00604f
C22997 VPWR.t2276 VGND 0.0141f
C22998 VPWR.t1215 VGND 0.0144f
C22999 VPWR.t2278 VGND 0.0153f
C23000 VPWR.t2272 VGND 0.0258f
C23001 VPWR.t2274 VGND 0.0052f
C23002 VPWR.t1886 VGND 0.017f
C23003 VPWR.t2533 VGND 0.0253f
C23004 VPWR.t1313 VGND 0.0358f
C23005 VPWR.t1759 VGND 0.0151f
C23006 VPWR.t460 VGND 0.0109f
C23007 VPWR.t1536 VGND 0.02f
C23008 VPWR.t1000 VGND 0.0151f
C23009 VPWR.t336 VGND 0.0264f
C23010 VPWR.t178 VGND 0.0211f
C23011 VPWR.t1526 VGND 0.0153f
C23012 VPWR.t1897 VGND 0.0252f
C23013 VPWR.t947 VGND 0.0154f
C23014 VPWR.t2169 VGND 0.0196f
C23015 VPWR.t2364 VGND 0.0141f
C23016 VPWR.t1745 VGND 0.0112f
C23017 VPWR.t2968 VGND 0.0311f
C23018 VPWR.t3135 VGND 0.0203f
C23019 VPWR.t412 VGND 0.0141f
C23020 VPWR.t2165 VGND 0.0232f
C23021 VPWR.t2895 VGND 0.021f
C23022 VPWR.t3254 VGND 0.00632f
C23023 VPWR.t3256 VGND 0.00676f
C23024 VPWR.n2116 VGND 0.0165f
C23025 VPWR.t3465 VGND 0.00911f
C23026 VPWR.t581 VGND 0.00391f
C23027 VPWR.n2117 VGND 0.0253f
C23028 VPWR.t582 VGND 0.00391f
C23029 VPWR.n2119 VGND 0.0138f
C23030 VPWR.n2120 VGND 0.00762f
C23031 VPWR.t94 VGND 0.0046f
C23032 VPWR.n2121 VGND 0.00407f
C23033 VPWR.t1902 VGND 0.00527f
C23034 VPWR.n2122 VGND 0.00619f
C23035 VPWR.t2598 VGND 0.00102f
C23036 VPWR.t1019 VGND 0.00102f
C23037 VPWR.n2123 VGND 0.00221f
C23038 VPWR.n2124 VGND 0.00591f
C23039 VPWR.t359 VGND 0.00387f
C23040 VPWR.t3382 VGND 0.0231f
C23041 VPWR.n2125 VGND 0.00179f
C23042 VPWR.t3466 VGND 0.0179f
C23043 VPWR.t583 VGND 0.00395f
C23044 VPWR.n2126 VGND 0.028f
C23045 VPWR.t584 VGND 0.00432f
C23046 VPWR.n2127 VGND 0.0103f
C23047 VPWR.n2128 VGND 0.0355f
C23048 VPWR.n2129 VGND 0.0103f
C23049 VPWR.t360 VGND 0.00399f
C23050 VPWR.n2130 VGND 0.0073f
C23051 VPWR.n2131 VGND 0.0153f
C23052 VPWR.n2132 VGND 0.0031f
C23053 VPWR.n2133 VGND 0.00524f
C23054 VPWR.n2134 VGND 0.00524f
C23055 VPWR.n2135 VGND 0.00393f
C23056 VPWR.n2136 VGND 0.0384f
C23057 VPWR.n2137 VGND 0.00837f
C23058 VPWR.n2138 VGND 0.00525f
C23059 VPWR.n2139 VGND 0.00179f
C23060 VPWR.n2140 VGND 0.00137f
C23061 VPWR.n2141 VGND 0.0031f
C23062 VPWR.n2142 VGND 0.00524f
C23063 VPWR.n2143 VGND 0.00524f
C23064 VPWR.n2144 VGND 0.00131f
C23065 VPWR.n2145 VGND 0.00524f
C23066 VPWR.t1148 VGND 0.0016f
C23067 VPWR.t1340 VGND 0.00208f
C23068 VPWR.n2146 VGND 0.00411f
C23069 VPWR.n2147 VGND 0.00513f
C23070 VPWR.t2107 VGND 0.00234f
C23071 VPWR.n2148 VGND 0.00391f
C23072 VPWR.n2149 VGND 2.92e-19
C23073 VPWR.n2150 VGND 0.00524f
C23074 VPWR.n2151 VGND 0.00475f
C23075 VPWR.n2152 VGND 0.00165f
C23076 VPWR.n2153 VGND 0.00274f
C23077 VPWR.n2154 VGND 0.0031f
C23078 VPWR.n2155 VGND 0.00639f
C23079 VPWR.n2156 VGND 0.00524f
C23080 VPWR.n2157 VGND 0.00506f
C23081 VPWR.n2158 VGND 0.00524f
C23082 VPWR.t979 VGND 6.73e-19
C23083 VPWR.t1154 VGND 9.96e-19
C23084 VPWR.n2159 VGND 0.00176f
C23085 VPWR.n2160 VGND 0.00658f
C23086 VPWR.n2161 VGND 0.00484f
C23087 VPWR.n2162 VGND 0.00524f
C23088 VPWR.n2163 VGND 0.00553f
C23089 VPWR.n2164 VGND 0.00524f
C23090 VPWR.t2928 VGND 0.00453f
C23091 VPWR.n2165 VGND 0.00799f
C23092 VPWR.n2166 VGND 0.00438f
C23093 VPWR.n2167 VGND 0.00524f
C23094 VPWR.n2168 VGND 0.0066f
C23095 VPWR.n2169 VGND 0.00524f
C23096 VPWR.t3555 VGND 0.0592f
C23097 VPWR.n2170 VGND 0.0356f
C23098 VPWR.n2171 VGND 0.00484f
C23099 VPWR.n2172 VGND 0.00524f
C23100 VPWR.n2173 VGND 0.00459f
C23101 VPWR.n2174 VGND 0.00524f
C23102 VPWR.t973 VGND 6.73e-19
C23103 VPWR.t3252 VGND 0.00127f
C23104 VPWR.n2175 VGND 0.00203f
C23105 VPWR.n2176 VGND 0.00594f
C23106 VPWR.n2177 VGND 0.00377f
C23107 VPWR.n2178 VGND 0.00524f
C23108 VPWR.n2179 VGND 0.00535f
C23109 VPWR.n2180 VGND 0.00524f
C23110 VPWR.t93 VGND 0.0046f
C23111 VPWR.t2367 VGND 0.00239f
C23112 VPWR.n2181 VGND 0.00636f
C23113 VPWR.n2182 VGND 0.00202f
C23114 VPWR.n2183 VGND 0.00233f
C23115 VPWR.n2184 VGND 0.00393f
C23116 VPWR.n2185 VGND 0.00444f
C23117 VPWR.n2186 VGND 0.00199f
C23118 VPWR.t2896 VGND 5.02e-19
C23119 VPWR.t2166 VGND 0.00135f
C23120 VPWR.n2187 VGND 0.00622f
C23121 VPWR.t3402 VGND 0.0179f
C23122 VPWR.n2188 VGND 0.0149f
C23123 VPWR.t2969 VGND 5.02e-19
C23124 VPWR.t1746 VGND 0.00135f
C23125 VPWR.n2189 VGND 0.00633f
C23126 VPWR.n2190 VGND 0.00138f
C23127 VPWR.n2191 VGND 5.41e-19
C23128 VPWR.n2192 VGND 2.85e-19
C23129 VPWR.n2193 VGND 6.54e-19
C23130 VPWR.n2194 VGND 8.67e-19
C23131 VPWR.n2195 VGND 0.0839f
C23132 VPWR.n2196 VGND 0.0057f
C23133 VPWR.n2197 VGND 6.54e-19
C23134 VPWR.n2198 VGND 8.67e-19
C23135 VPWR.n2199 VGND 4.39e-19
C23136 VPWR.n2200 VGND 3.29e-19
C23137 VPWR.n2201 VGND 5.27e-19
C23138 VPWR.n2202 VGND 2.85e-19
C23139 VPWR.n2203 VGND 2.85e-19
C23140 VPWR.n2204 VGND 4.17e-19
C23141 VPWR.n2205 VGND 5.71e-19
C23142 VPWR.n2206 VGND 4.17e-19
C23143 VPWR.n2207 VGND 3.51e-19
C23144 VPWR.n2208 VGND 4.61e-19
C23145 VPWR.n2209 VGND 4.17e-19
C23146 VPWR.n2210 VGND 4.83e-19
C23147 VPWR.n2211 VGND 4.61e-19
C23148 VPWR.n2212 VGND 3.73e-19
C23149 VPWR.n2213 VGND 2.41e-19
C23150 VPWR.t997 VGND 0.00455f
C23151 VPWR.n2214 VGND 0.00727f
C23152 VPWR.t2882 VGND 0.00242f
C23153 VPWR.t2025 VGND 0.00695f
C23154 VPWR.t3517 VGND 0.00911f
C23155 VPWR.t567 VGND 0.00391f
C23156 VPWR.n2215 VGND 0.0253f
C23157 VPWR.t566 VGND 0.00391f
C23158 VPWR.n2217 VGND 0.0138f
C23159 VPWR.n2218 VGND 0.00345f
C23160 VPWR.t3378 VGND 0.00911f
C23161 VPWR.t328 VGND 0.00391f
C23162 VPWR.n2219 VGND 0.0253f
C23163 VPWR.t329 VGND 0.00391f
C23164 VPWR.n2221 VGND 0.0138f
C23165 VPWR.n2222 VGND 0.011f
C23166 VPWR.n2223 VGND 0.00786f
C23167 VPWR.n2224 VGND 0.00393f
C23168 VPWR.t2310 VGND 0.00136f
C23169 VPWR.t1146 VGND 0.00136f
C23170 VPWR.n2225 VGND 0.00328f
C23171 VPWR.n2226 VGND 0.00727f
C23172 VPWR.n2227 VGND 0.00524f
C23173 VPWR.n2228 VGND 0.0031f
C23174 VPWR.t2027 VGND 0.00166f
C23175 VPWR.t2029 VGND 0.00166f
C23176 VPWR.n2229 VGND 0.00345f
C23177 VPWR.n2230 VGND 0.00469f
C23178 VPWR.n2231 VGND 0.00152f
C23179 VPWR.n2232 VGND 0.00393f
C23180 VPWR.t1648 VGND 0.00676f
C23181 VPWR.t2023 VGND 0.00225f
C23182 VPWR.t815 VGND 0.00166f
C23183 VPWR.n2233 VGND 0.00438f
C23184 VPWR.n2234 VGND 0.00631f
C23185 VPWR.n2235 VGND 0.0087f
C23186 VPWR.n2236 VGND 9.68e-19
C23187 VPWR.n2237 VGND 0.00524f
C23188 VPWR.n2238 VGND 0.0031f
C23189 VPWR.n2239 VGND 9.48e-19
C23190 VPWR.n2240 VGND 0.00484f
C23191 VPWR.n2241 VGND 0.00117f
C23192 VPWR.n2242 VGND 0.00393f
C23193 VPWR.t961 VGND 6.73e-19
C23194 VPWR.t1646 VGND 0.00127f
C23195 VPWR.n2243 VGND 0.00203f
C23196 VPWR.n2244 VGND 0.00324f
C23197 VPWR.n2245 VGND 0.00106f
C23198 VPWR.n2246 VGND 0.00524f
C23199 VPWR.t913 VGND 0.00102f
C23200 VPWR.t858 VGND 0.00154f
C23201 VPWR.n2247 VGND 0.00483f
C23202 VPWR.n2248 VGND 0.00658f
C23203 VPWR.n2249 VGND 0.00125f
C23204 VPWR.n2250 VGND 0.00524f
C23205 VPWR.n2251 VGND 0.00186f
C23206 VPWR.n2252 VGND 0.00524f
C23207 VPWR.n2253 VGND 0.00178f
C23208 VPWR.n2254 VGND 0.0031f
C23209 VPWR.n2255 VGND 0.00393f
C23210 VPWR.n2256 VGND 0.00333f
C23211 VPWR.n2257 VGND 0.00118f
C23212 VPWR.t977 VGND 6.73e-19
C23213 VPWR.t2300 VGND 9.96e-19
C23214 VPWR.n2258 VGND 0.00176f
C23215 VPWR.n2259 VGND 0.00421f
C23216 VPWR.n2260 VGND 0.00136f
C23217 VPWR.n2261 VGND 0.00393f
C23218 VPWR.t2705 VGND 0.00166f
C23219 VPWR.t868 VGND 0.00166f
C23220 VPWR.n2262 VGND 0.0037f
C23221 VPWR.n2263 VGND 0.0061f
C23222 VPWR.n2264 VGND 5.14e-19
C23223 VPWR.n2265 VGND 0.00524f
C23224 VPWR.n2266 VGND 0.00184f
C23225 VPWR.n2267 VGND 0.00524f
C23226 VPWR.n2268 VGND 0.0015f
C23227 VPWR.n2269 VGND 0.0039f
C23228 VPWR.n2270 VGND 9e-19
C23229 VPWR.n2271 VGND 0.00138f
C23230 VPWR.n2272 VGND 9.06e-19
C23231 VPWR.n2273 VGND 5.48e-19
C23232 VPWR.n2274 VGND 6.14e-19
C23233 VPWR.n2275 VGND 0.00138f
C23234 VPWR.n2276 VGND 0.0023f
C23235 VPWR.t2708 VGND 0.00598f
C23236 VPWR.n2277 VGND 0.00856f
C23237 VPWR.n2278 VGND 0.00139f
C23238 VPWR.n2279 VGND 4.45e-19
C23239 VPWR.n2280 VGND 4.27e-19
C23240 VPWR.n2281 VGND 6.83e-19
C23241 VPWR.n2282 VGND 3.7e-19
C23242 VPWR.n2283 VGND 9.68e-19
C23243 VPWR.n2284 VGND 9.96e-19
C23244 VPWR.n2285 VGND 5.41e-19
C23245 VPWR.n2286 VGND 7.4e-19
C23246 VPWR.n2287 VGND 3.13e-19
C23247 VPWR.t1625 VGND 0.00238f
C23248 VPWR.n2288 VGND 0.00468f
C23249 VPWR.n2289 VGND 2.31e-19
C23250 VPWR.n2290 VGND 4.81e-19
C23251 VPWR.n2291 VGND 2.56e-19
C23252 VPWR.t915 VGND 0.00102f
C23253 VPWR.t1027 VGND 0.00102f
C23254 VPWR.n2292 VGND 0.00218f
C23255 VPWR.n2293 VGND 0.015f
C23256 VPWR.n2294 VGND 0.00524f
C23257 VPWR.n2295 VGND 0.0117f
C23258 VPWR.t3334 VGND 0.0289f
C23259 VPWR.t200 VGND 0.00387f
C23260 VPWR.n2296 VGND 0.0604f
C23261 VPWR.n2297 VGND 0.0146f
C23262 VPWR.t2693 VGND 0.00136f
C23263 VPWR.t2904 VGND 0.00136f
C23264 VPWR.n2298 VGND 0.00317f
C23265 VPWR.t201 VGND 0.00387f
C23266 VPWR.t3301 VGND 0.00676f
C23267 VPWR.n2299 VGND 0.00944f
C23268 VPWR.n2300 VGND 0.0031f
C23269 VPWR.t327 VGND 0.0515f
C23270 VPWR.t2309 VGND 0.0405f
C23271 VPWR.t2024 VGND 0.0148f
C23272 VPWR.t1145 VGND 0.0144f
C23273 VPWR.t2026 VGND 0.0109f
C23274 VPWR.t2028 VGND 0.0191f
C23275 VPWR.t2022 VGND 0.0159f
C23276 VPWR.t1647 VGND 0.0161f
C23277 VPWR.t814 VGND 0.0257f
C23278 VPWR.t2881 VGND 0.0245f
C23279 VPWR.t960 VGND 0.0206f
C23280 VPWR.t857 VGND 0.0181f
C23281 VPWR.t1645 VGND 0.0163f
C23282 VPWR.t912 VGND 0.0141f
C23283 VPWR.t2305 VGND 0.0121f
C23284 VPWR.t870 VGND 0.0144f
C23285 VPWR.t916 VGND 0.0178f
C23286 VPWR.t996 VGND 0.0311f
C23287 VPWR.t976 VGND 0.021f
C23288 VPWR.t2704 VGND 0.0163f
C23289 VPWR.t2299 VGND 0.0144f
C23290 VPWR.t867 VGND 0.0208f
C23291 VPWR.t911 VGND 0.017f
C23292 VPWR.t917 VGND 0.0193f
C23293 VPWR.t2306 VGND 0.0289f
C23294 VPWR.t2707 VGND 0.0154f
C23295 VPWR.t1624 VGND 0.0112f
C23296 VPWR.t914 VGND 0.0509f
C23297 VPWR.t1026 VGND 0.025f
C23298 VPWR.t199 VGND 0.0206f
C23299 VPWR.t2692 VGND 0.0305f
C23300 VPWR.t2903 VGND 0.0257f
C23301 VPWR.t3300 VGND 0.0126f
C23302 VPWR.t1874 VGND 0.0311f
C23303 VPWR.t2016 VGND 0.0109f
C23304 VPWR.t2883 VGND 0.0052f
C23305 VPWR.t1618 VGND 0.0153f
C23306 VPWR.t871 VGND 0.0311f
C23307 VPWR.t1344 VGND 0.0109f
C23308 VPWR.t2101 VGND 0.0148f
C23309 VPWR.t1619 VGND 0.0148f
C23310 VPWR.t1926 VGND 0.0213f
C23311 VPWR.t2886 VGND 0.0109f
C23312 VPWR.t1024 VGND 0.0151f
C23313 VPWR.t2261 VGND 0.0148f
C23314 VPWR.t1337 VGND 0.0161f
C23315 VPWR.t1922 VGND 0.0361f
C23316 VPWR.t1928 VGND 0.0235f
C23317 VPWR.t2283 VGND 0.0321f
C23318 VPWR.t2263 VGND 0.0401f
C23319 VPWR.t1821 VGND 0.0398f
C23320 VPWR.t974 VGND 0.0242f
C23321 VPWR.t291 VGND 0.0331f
C23322 VPWR.t2081 VGND 0.0418f
C23323 VPWR.t2260 VGND 0.0311f
C23324 VPWR.t2282 VGND 0.0285f
C23325 VPWR.t3302 VGND 0.0322f
C23326 VPWR.t958 VGND 0.027f
C23327 VPWR.t2256 VGND 0.0339f
C23328 VPWR.n2301 VGND 0.0396f
C23329 VPWR.n2302 VGND 0.00902f
C23330 VPWR.t292 VGND 0.0046f
C23331 VPWR.t959 VGND 6.73e-19
C23332 VPWR.t3303 VGND 0.00127f
C23333 VPWR.n2303 VGND 0.00203f
C23334 VPWR.n2304 VGND 0.00572f
C23335 VPWR.n2305 VGND 0.00123f
C23336 VPWR.t293 VGND 0.0046f
C23337 VPWR.n2306 VGND 0.00407f
C23338 VPWR.t1923 VGND 0.0016f
C23339 VPWR.t1338 VGND 0.00208f
C23340 VPWR.n2307 VGND 0.00422f
C23341 VPWR.n2308 VGND 0.00613f
C23342 VPWR.t2262 VGND 0.00102f
C23343 VPWR.t1025 VGND 0.00102f
C23344 VPWR.n2309 VGND 0.00221f
C23345 VPWR.n2310 VGND 0.00577f
C23346 VPWR.n2311 VGND 0.00114f
C23347 VPWR.t2887 VGND 0.00527f
C23348 VPWR.n2312 VGND 0.00615f
C23349 VPWR.t1927 VGND 0.0016f
C23350 VPWR.t1345 VGND 0.00208f
C23351 VPWR.n2313 VGND 0.00422f
C23352 VPWR.n2314 VGND 0.00644f
C23353 VPWR.t872 VGND 0.00527f
C23354 VPWR.t2017 VGND 0.00136f
C23355 VPWR.t1875 VGND 0.00136f
C23356 VPWR.n2315 VGND 0.00328f
C23357 VPWR.n2316 VGND 0.0079f
C23358 VPWR.n2317 VGND 0.00202f
C23359 VPWR.n2318 VGND 0.00134f
C23360 VPWR.n2319 VGND 0.00262f
C23361 VPWR.n2320 VGND 0.00262f
C23362 VPWR.n2321 VGND 0.00179f
C23363 VPWR.n2322 VGND 0.00152f
C23364 VPWR.n2323 VGND 0.00149f
C23365 VPWR.n2324 VGND 0.00333f
C23366 VPWR.n2325 VGND 0.00393f
C23367 VPWR.n2326 VGND 0.0065f
C23368 VPWR.n2327 VGND 0.00135f
C23369 VPWR.n2328 VGND 0.0031f
C23370 VPWR.n2329 VGND 0.00524f
C23371 VPWR.n2330 VGND 0.00393f
C23372 VPWR.n2331 VGND 0.0031f
C23373 VPWR.n2332 VGND 0.00524f
C23374 VPWR.n2333 VGND 0.00524f
C23375 VPWR.n2334 VGND 0.00475f
C23376 VPWR.n2335 VGND 0.00116f
C23377 VPWR.t1929 VGND 0.00235f
C23378 VPWR.n2336 VGND 0.00493f
C23379 VPWR.n2337 VGND 0.00102f
C23380 VPWR.n2338 VGND 0.0031f
C23381 VPWR.n2339 VGND 0.00639f
C23382 VPWR.n2340 VGND 0.00524f
C23383 VPWR.n2341 VGND 0.0066f
C23384 VPWR.n2342 VGND 0.00524f
C23385 VPWR.n2343 VGND 0.0066f
C23386 VPWR.n2344 VGND 0.00524f
C23387 VPWR.n2345 VGND 0.00506f
C23388 VPWR.n2346 VGND 0.00524f
C23389 VPWR.t975 VGND 6.73e-19
C23390 VPWR.t1822 VGND 9.96e-19
C23391 VPWR.n2347 VGND 0.00176f
C23392 VPWR.n2348 VGND 0.00658f
C23393 VPWR.n2349 VGND 0.00484f
C23394 VPWR.n2350 VGND 0.00524f
C23395 VPWR.n2351 VGND 0.00553f
C23396 VPWR.n2352 VGND 0.00524f
C23397 VPWR.t3365 VGND 0.0592f
C23398 VPWR.n2353 VGND 0.0356f
C23399 VPWR.t2082 VGND 0.00453f
C23400 VPWR.n2354 VGND 0.00799f
C23401 VPWR.n2355 VGND 0.00262f
C23402 VPWR.n2356 VGND 0.00524f
C23403 VPWR.n2357 VGND 0.00506f
C23404 VPWR.n2358 VGND 0.00524f
C23405 VPWR.n2359 VGND 0.0066f
C23406 VPWR.n2360 VGND 0.00524f
C23407 VPWR.n2361 VGND 0.00614f
C23408 VPWR.n2362 VGND 0.00524f
C23409 VPWR.n2363 VGND 0.00393f
C23410 VPWR.n2364 VGND 0.00269f
C23411 VPWR.n2365 VGND 0.00107f
C23412 VPWR.n2366 VGND 0.00333f
C23413 VPWR.t2257 VGND 0.00242f
C23414 VPWR.n2367 VGND 0.00484f
C23415 VPWR.n2368 VGND 9.48e-19
C23416 VPWR.n2369 VGND 0.00393f
C23417 VPWR.n2370 VGND 0.00199f
C23418 VPWR.n2371 VGND 0.00179f
C23419 VPWR.n2372 VGND 0.00521f
C23420 VPWR.n2373 VGND 0.00837f
C23421 VPWR.n2374 VGND 0.0133f
C23422 VPWR.n2375 VGND 0.0192f
C23423 VPWR.n2376 VGND 0.0113f
C23424 VPWR.n2377 VGND 0.00393f
C23425 VPWR.n2378 VGND 0.00513f
C23426 VPWR.n2379 VGND 5.27e-19
C23427 VPWR.n2380 VGND 3.95e-19
C23428 VPWR.n2381 VGND 5.05e-19
C23429 VPWR.n2382 VGND 5.05e-19
C23430 VPWR.n2383 VGND 8.67e-19
C23431 VPWR.n2384 VGND 6.54e-19
C23432 VPWR.n2385 VGND 9.06e-19
C23433 VPWR.n2386 VGND 0.0994f
C23434 VPWR.n2388 VGND 0.00139f
C23435 VPWR.n2389 VGND 5.48e-19
C23436 VPWR.n2390 VGND 3.07e-19
C23437 VPWR.n2391 VGND 0.00138f
C23438 VPWR.n2392 VGND 0.0058f
C23439 VPWR.n2393 VGND 0.00124f
C23440 VPWR.n2394 VGND 2.92e-19
C23441 VPWR.n2395 VGND 7.65e-19
C23442 VPWR.n2396 VGND 6.83e-19
C23443 VPWR.n2397 VGND 4.84e-19
C23444 VPWR.n2398 VGND 1.99e-19
C23445 VPWR.n2399 VGND 8.26e-19
C23446 VPWR.n2400 VGND 4.83e-19
C23447 VPWR.n2401 VGND 4.61e-19
C23448 VPWR.n2402 VGND 4.11e-19
C23449 VPWR.n2403 VGND 4.11e-19
C23450 VPWR.n2404 VGND 7.39e-19
C23451 VPWR.n2405 VGND 5.19e-19
C23452 VPWR.n2406 VGND 7.39e-19
C23453 VPWR.n2407 VGND 4.11e-19
C23454 VPWR.n2408 VGND 4.11e-19
C23455 VPWR.n2410 VGND 0.1f
C23456 VPWR.n2411 VGND 0.1f
C23457 VPWR.n2412 VGND 8.67e-19
C23458 VPWR.n2413 VGND 6.54e-19
C23459 VPWR.n2414 VGND 9.06e-19
C23460 VPWR.n2415 VGND 0.00139f
C23461 VPWR.n2416 VGND 5.27e-19
C23462 VPWR.n2417 VGND 3.95e-19
C23463 VPWR.n2418 VGND 5.05e-19
C23464 VPWR.n2419 VGND 5.05e-19
C23465 VPWR.n2420 VGND 3.07e-19
C23466 VPWR.n2421 VGND 5.48e-19
C23467 VPWR.t3577 VGND 0.0179f
C23468 VPWR.t338 VGND 0.00399f
C23469 VPWR.n2423 VGND 0.0129f
C23470 VPWR.n2424 VGND 0.00475f
C23471 VPWR.t1537 VGND 0.00136f
C23472 VPWR.t1001 VGND 0.00136f
C23473 VPWR.n2425 VGND 0.00317f
C23474 VPWR.t3377 VGND 0.0179f
C23475 VPWR.n2426 VGND 0.00513f
C23476 VPWR.n2427 VGND 0.00524f
C23477 VPWR.t1314 VGND 0.00136f
C23478 VPWR.t1760 VGND 0.00136f
C23479 VPWR.n2428 VGND 0.00317f
C23480 VPWR.t3425 VGND 0.0179f
C23481 VPWR.t1887 VGND 0.00136f
C23482 VPWR.t2534 VGND 0.00136f
C23483 VPWR.n2429 VGND 0.00317f
C23484 VPWR.n2430 VGND 0.00653f
C23485 VPWR.t2279 VGND 0.00166f
C23486 VPWR.t2273 VGND 0.00166f
C23487 VPWR.n2431 VGND 0.00345f
C23488 VPWR.n2432 VGND 0.00131f
C23489 VPWR.t1212 VGND 0.00166f
C23490 VPWR.t2277 VGND 0.00225f
C23491 VPWR.n2433 VGND 0.0045f
C23492 VPWR.t3513 VGND 0.00911f
C23493 VPWR.t726 VGND 0.00391f
C23494 VPWR.n2434 VGND 0.0253f
C23495 VPWR.t725 VGND 0.00391f
C23496 VPWR.n2436 VGND 0.0138f
C23497 VPWR.t3450 VGND 0.00911f
C23498 VPWR.t540 VGND 0.00391f
C23499 VPWR.n2437 VGND 0.0253f
C23500 VPWR.t541 VGND 0.00391f
C23501 VPWR.n2439 VGND 0.0138f
C23502 VPWR.n2440 VGND 0.0112f
C23503 VPWR.n2441 VGND 0.00345f
C23504 VPWR.n2442 VGND 0.00179f
C23505 VPWR.n2443 VGND 0.00179f
C23506 VPWR.t1214 VGND 0.00646f
C23507 VPWR.n2444 VGND 0.0137f
C23508 VPWR.n2445 VGND 0.00121f
C23509 VPWR.n2446 VGND 0.00475f
C23510 VPWR.n2447 VGND 0.00393f
C23511 VPWR.t1216 VGND 0.00647f
C23512 VPWR.n2448 VGND 0.0104f
C23513 VPWR.t2275 VGND 0.00682f
C23514 VPWR.n2449 VGND 0.00711f
C23515 VPWR.n2450 VGND 0.00151f
C23516 VPWR.n2451 VGND 0.00179f
C23517 VPWR.n2452 VGND 0.00344f
C23518 VPWR.n2453 VGND 0.00393f
C23519 VPWR.n2454 VGND 0.00199f
C23520 VPWR.n2455 VGND 0.00173f
C23521 VPWR.n2456 VGND 0.00525f
C23522 VPWR.t461 VGND 0.00387f
C23523 VPWR.n2457 VGND 0.00493f
C23524 VPWR.n2458 VGND 0.0173f
C23525 VPWR.n2459 VGND 0.0158f
C23526 VPWR.t462 VGND 0.00387f
C23527 VPWR.n2460 VGND 0.00837f
C23528 VPWR.n2461 VGND 0.0133f
C23529 VPWR.n2462 VGND 0.0031f
C23530 VPWR.n2463 VGND 0.00179f
C23531 VPWR.n2464 VGND 0.00179f
C23532 VPWR.n2465 VGND 0.00513f
C23533 VPWR.t337 VGND 0.00387f
C23534 VPWR.n2466 VGND 0.00493f
C23535 VPWR.n2467 VGND 0.0173f
C23536 VPWR.n2468 VGND 0.0158f
C23537 VPWR.n2469 VGND 0.0126f
C23538 VPWR.n2470 VGND 0.00393f
C23539 VPWR.n2471 VGND 0.00179f
C23540 VPWR.n2472 VGND 0.00443f
C23541 VPWR.t179 VGND 0.00387f
C23542 VPWR.n2473 VGND 0.00493f
C23543 VPWR.n2474 VGND 0.0173f
C23544 VPWR.n2475 VGND 0.0103f
C23545 VPWR.n2476 VGND 0.00393f
C23546 VPWR.t1527 VGND 0.00166f
C23547 VPWR.t1898 VGND 0.00166f
C23548 VPWR.n2477 VGND 0.0037f
C23549 VPWR.t180 VGND 0.00387f
C23550 VPWR.n2478 VGND 0.00247f
C23551 VPWR.n2479 VGND 0.00628f
C23552 VPWR.n2480 VGND 0.0111f
C23553 VPWR.n2481 VGND 0.00702f
C23554 VPWR.n2482 VGND 0.0039f
C23555 VPWR.n2483 VGND 5.41e-19
C23556 VPWR.n2484 VGND 5.12e-19
C23557 VPWR.n2485 VGND 3.7e-19
C23558 VPWR.n2486 VGND 4.39e-19
C23559 VPWR.n2487 VGND 3.29e-19
C23560 VPWR.n2488 VGND 2.85e-19
C23561 VPWR.n2489 VGND 5.27e-19
C23562 VPWR.n2490 VGND 7.47e-19
C23563 VPWR.n2491 VGND 0.00453f
C23564 VPWR.n2492 VGND 4.27e-19
C23565 VPWR.n2493 VGND 1.14e-19
C23566 VPWR.n2494 VGND 4.27e-19
C23567 VPWR.n2495 VGND 0.00153f
C23568 VPWR.n2496 VGND 0.00206f
C23569 VPWR.n2497 VGND 0.00138f
C23570 VPWR.n2498 VGND 9e-19
C23571 VPWR.n2499 VGND 6.14e-19
C23572 VPWR.n2500 VGND 9.06e-19
C23573 VPWR.n2501 VGND 5.48e-19
C23574 VPWR.n2502 VGND 0.00138f
C23575 VPWR.n2503 VGND 0.0057f
C23576 VPWR.n2505 VGND 4.83e-19
C23577 VPWR.n2506 VGND 4.61e-19
C23578 VPWR.n2507 VGND 3.73e-19
C23579 VPWR.n2508 VGND 2.41e-19
C23580 VPWR.n2509 VGND 4.83e-19
C23581 VPWR.n2510 VGND 4.61e-19
C23582 VPWR.n2511 VGND 4.11e-19
C23583 VPWR.n2512 VGND 4.11e-19
C23584 VPWR.n2513 VGND 7.39e-19
C23585 VPWR.n2514 VGND 5.19e-19
C23586 VPWR.n2515 VGND 7.39e-19
C23587 VPWR.n2516 VGND 4.11e-19
C23588 VPWR.n2517 VGND 4.11e-19
C23589 VPWR.n2518 VGND 4.17e-19
C23590 VPWR.n2519 VGND 4.61e-19
C23591 VPWR.n2520 VGND 3.51e-19
C23592 VPWR.n2521 VGND 4.17e-19
C23593 VPWR.n2522 VGND 4.17e-19
C23594 VPWR.n2523 VGND 5.71e-19
C23595 VPWR.n2524 VGND 7.4e-19
C23596 VPWR.n2525 VGND 7.64e-19
C23597 VPWR.n2526 VGND 3.13e-19
C23598 VPWR.n2527 VGND 1.71e-19
C23599 VPWR.n2528 VGND 2.56e-19
C23600 VPWR.n2529 VGND 4.55e-19
C23601 VPWR.t2170 VGND 0.00261f
C23602 VPWR.n2530 VGND 0.00525f
C23603 VPWR.n2531 VGND 3.93e-19
C23604 VPWR.n2532 VGND 2.56e-19
C23605 VPWR.n2533 VGND 9.68e-19
C23606 VPWR.n2534 VGND 3.13e-19
C23607 VPWR.n2535 VGND 4.84e-19
C23608 VPWR.n2536 VGND 6.83e-19
C23609 VPWR.n2537 VGND 4.64e-19
C23610 VPWR.n2538 VGND 4.84e-19
C23611 VPWR.n2539 VGND 1.41e-19
C23612 VPWR.n2540 VGND 4.27e-19
C23613 VPWR.t2365 VGND 0.00587f
C23614 VPWR.n2541 VGND 0.00626f
C23615 VPWR.n2542 VGND 9.07e-20
C23616 VPWR.n2543 VGND 4.27e-19
C23617 VPWR.n2544 VGND 9.28e-19
C23618 VPWR.n2545 VGND 9.6e-19
C23619 VPWR.n2546 VGND 0.00217f
C23620 VPWR.n2547 VGND 0.00237f
C23621 VPWR.n2548 VGND 0.00102f
C23622 VPWR.n2549 VGND 0.00696f
C23623 VPWR.n2550 VGND 0.00102f
C23624 VPWR.n2551 VGND 0.00393f
C23625 VPWR.n2552 VGND 0.00333f
C23626 VPWR.n2553 VGND 0.00173f
C23627 VPWR.t413 VGND 0.00387f
C23628 VPWR.t3136 VGND 0.00261f
C23629 VPWR.n2554 VGND 0.00762f
C23630 VPWR.n2555 VGND 0.00441f
C23631 VPWR.n2556 VGND 0.00525f
C23632 VPWR.n2557 VGND 0.00179f
C23633 VPWR.n2558 VGND 0.0031f
C23634 VPWR.n2559 VGND 0.00524f
C23635 VPWR.n2560 VGND 0.00475f
C23636 VPWR.n2561 VGND 0.0103f
C23637 VPWR.n2562 VGND 0.0106f
C23638 VPWR.n2563 VGND 0.0119f
C23639 VPWR.t414 VGND 0.00387f
C23640 VPWR.n2564 VGND 0.00463f
C23641 VPWR.n2565 VGND 0.00487f
C23642 VPWR.n2566 VGND 0.00991f
C23643 VPWR.n2567 VGND 0.0412f
C23644 VPWR.t3253 VGND 0.0309f
C23645 VPWR.t580 VGND 0.0141f
C23646 VPWR.t3255 VGND 0.0183f
C23647 VPWR.t2366 VGND 0.0399f
C23648 VPWR.t972 VGND 0.0322f
C23649 VPWR.t3251 VGND 0.0322f
C23650 VPWR.t1879 VGND 0.0285f
C23651 VPWR.t2596 VGND 0.0253f
C23652 VPWR.t92 VGND 0.0166f
C23653 VPWR.t2927 VGND 0.0388f
C23654 VPWR.t978 VGND 0.0493f
C23655 VPWR.t1153 VGND 0.0398f
C23656 VPWR.t2595 VGND 0.0327f
C23657 VPWR.t1878 VGND 0.0206f
C23658 VPWR.t1147 VGND 0.0154f
C23659 VPWR.t2106 VGND 0.0154f
C23660 VPWR.t1339 VGND 0.029f
C23661 VPWR.t1901 VGND 0.0316f
C23662 VPWR.t2597 VGND 0.0299f
C23663 VPWR.t1018 VGND 0.0154f
C23664 VPWR.t1620 VGND 0.0109f
C23665 VPWR.t869 VGND 0.0154f
C23666 VPWR.t358 VGND 0.0618f
C23667 VPWR.t2761 VGND 0.0111f
C23668 VPWR.t2931 VGND 0.00504f
C23669 VPWR.t3197 VGND 0.0154f
C23670 VPWR.t3199 VGND 0.0311f
C23671 VPWR.t1713 VGND 0.0248f
C23672 VPWR.t1711 VGND 0.0282f
C23673 VPWR.t764 VGND 0.0164f
C23674 VPWR.t646 VGND 0.0141f
C23675 VPWR.t766 VGND 0.0358f
C23676 VPWR.t83 VGND 0.026f
C23677 VPWR.t1159 VGND 0.028f
C23678 VPWR.t1161 VGND 0.0178f
C23679 VPWR.t753 VGND 0.0141f
C23680 VPWR.t1157 VGND 0.0121f
C23681 VPWR.t2322 VGND 0.0141f
C23682 VPWR.t1163 VGND 0.0163f
C23683 VPWR.t1504 VGND 0.0141f
C23684 VPWR.t1530 VGND 0.0312f
C23685 VPWR.t2407 VGND 0.0114f
C23686 VPWR.t749 VGND 0.0158f
C23687 VPWR.t848 VGND 0.0141f
C23688 VPWR.t754 VGND 0.0159f
C23689 VPWR.t751 VGND 0.0282f
C23690 VPWR.t756 VGND 0.0163f
C23691 VPWR.t1858 VGND 0.0141f
C23692 VPWR.t1681 VGND 0.0159f
C23693 VPWR.t1528 VGND 0.00906f
C23694 VPWR.t1679 VGND 0.0159f
C23695 VPWR.t1680 VGND 0.0151f
C23696 VPWR.t1682 VGND 0.0178f
C23697 VPWR.t1905 VGND 0.0277f
C23698 VPWR.t846 VGND 0.0134f
C23699 VPWR.t2909 VGND 0.018f
C23700 VPWR.n2568 VGND 0.0191f
C23701 VPWR.n2569 VGND 0.00929f
C23702 VPWR.n2570 VGND 0.00199f
C23703 VPWR.n2571 VGND 0.00199f
C23704 VPWR.n2572 VGND 0.00125f
C23705 VPWR.n2573 VGND 0.00186f
C23706 VPWR.n2574 VGND 0.00393f
C23707 VPWR.n2575 VGND 0.0031f
C23708 VPWR.n2576 VGND 0.00175f
C23709 VPWR.n2577 VGND 9.28e-19
C23710 VPWR.n2578 VGND 0.00128f
C23711 VPWR.n2579 VGND 2.85e-19
C23712 VPWR.n2580 VGND 1.71e-19
C23713 VPWR.n2581 VGND 2.28e-19
C23714 VPWR.n2582 VGND 9.28e-19
C23715 VPWR.n2583 VGND 6.26e-19
C23716 VPWR.n2584 VGND 4.84e-19
C23717 VPWR.n2585 VGND 5.98e-19
C23718 VPWR.n2586 VGND 5.12e-19
C23719 VPWR.n2587 VGND 7.12e-19
C23720 VPWR.n2588 VGND 5.98e-19
C23721 VPWR.n2589 VGND 2.56e-19
C23722 VPWR.n2590 VGND 1.76e-19
C23723 VPWR.n2591 VGND 3.95e-19
C23724 VPWR.n2592 VGND 7.68e-19
C23725 VPWR.n2593 VGND 5.05e-19
C23726 VPWR.n2594 VGND 1.76e-19
C23727 VPWR.n2595 VGND 5.48e-19
C23728 VPWR.n2597 VGND 0.1f
C23729 VPWR.n2598 VGND 0.1f
C23730 VPWR.n2599 VGND 6.54e-19
C23731 VPWR.n2600 VGND 8.67e-19
C23732 VPWR.n2601 VGND 4.83e-19
C23733 VPWR.n2602 VGND 2.85e-19
C23734 VPWR.n2603 VGND 3.95e-19
C23735 VPWR.n2604 VGND 3.95e-19
C23736 VPWR.n2605 VGND 4.17e-19
C23737 VPWR.n2606 VGND 2.85e-19
C23738 VPWR.n2607 VGND 2.85e-19
C23739 VPWR.n2608 VGND 4.11e-19
C23740 VPWR.n2609 VGND 4.11e-19
C23741 VPWR.n2610 VGND 7.39e-19
C23742 VPWR.n2611 VGND 5.19e-19
C23743 VPWR.n2612 VGND 7.39e-19
C23744 VPWR.n2613 VGND 4.11e-19
C23745 VPWR.n2614 VGND 3.95e-19
C23746 VPWR.n2615 VGND 4.61e-19
C23747 VPWR.n2616 VGND 2.41e-19
C23748 VPWR.n2617 VGND 3.95e-19
C23749 VPWR.n2618 VGND 5.05e-19
C23750 VPWR.n2619 VGND 4.17e-19
C23751 VPWR.n2620 VGND 6.14e-19
C23752 VPWR.n2621 VGND 4.39e-19
C23753 VPWR.n2622 VGND 1.76e-19
C23754 VPWR.n2623 VGND 3.07e-19
C23755 VPWR.n2624 VGND 4.11e-19
C23756 VPWR.n2626 VGND 9.06e-19
C23757 VPWR.n2627 VGND 5.48e-19
C23758 VPWR.n2628 VGND 0.00138f
C23759 VPWR.n2629 VGND 0.0057f
C23760 VPWR.n2630 VGND 0.0994f
C23761 VPWR.n2632 VGND 0.00139f
C23762 VPWR.n2633 VGND 5.48e-19
C23763 VPWR.n2634 VGND 4.17e-19
C23764 VPWR.n2635 VGND 0.00137f
C23765 VPWR.n2636 VGND 0.00218f
C23766 VPWR.t2447 VGND 0.00166f
C23767 VPWR.t2449 VGND 0.00166f
C23768 VPWR.n2637 VGND 0.00359f
C23769 VPWR.n2638 VGND 0.00523f
C23770 VPWR.n2639 VGND 0.00119f
C23771 VPWR.n2640 VGND 6.8e-19
C23772 VPWR.n2641 VGND 5.69e-19
C23773 VPWR.n2642 VGND 0.00131f
C23774 VPWR.n2643 VGND 9.96e-19
C23775 VPWR.n2644 VGND 4.27e-19
C23776 VPWR.n2645 VGND 5.12e-19
C23777 VPWR.n2646 VGND 5.41e-19
C23778 VPWR.n2647 VGND 7.76e-19
C23779 VPWR.n2648 VGND 5.41e-19
C23780 VPWR.n2649 VGND 1.31e-19
C23781 VPWR.n2650 VGND 3.7e-19
C23782 VPWR.n2651 VGND 1.21e-19
C23783 VPWR.n2652 VGND 3.42e-19
C23784 VPWR.n2653 VGND 7.46e-19
C23785 VPWR.n2654 VGND 3.7e-19
C23786 VPWR.n2655 VGND 6.26e-19
C23787 VPWR.n2656 VGND 6.55e-19
C23788 VPWR.n2657 VGND 5.41e-19
C23789 VPWR.n2658 VGND 9.96e-19
C23790 VPWR.n2659 VGND 9.68e-19
C23791 VPWR.n2660 VGND 5.41e-19
C23792 VPWR.t971 VGND 6.73e-19
C23793 VPWR.t3035 VGND 0.00127f
C23794 VPWR.n2661 VGND 0.00203f
C23795 VPWR.t2441 VGND 0.00556f
C23796 VPWR.n2662 VGND 0.00617f
C23797 VPWR.n2663 VGND 0.0028f
C23798 VPWR.n2664 VGND 9.88e-19
C23799 VPWR.n2665 VGND 3.13e-19
C23800 VPWR.n2666 VGND 5.98e-19
C23801 VPWR.n2667 VGND 5.12e-19
C23802 VPWR.n2668 VGND 7.12e-19
C23803 VPWR.n2669 VGND 5.98e-19
C23804 VPWR.n2670 VGND 3.13e-19
C23805 VPWR.n2671 VGND 1.77e-19
C23806 VPWR.n2672 VGND 3.95e-19
C23807 VPWR.n2673 VGND 8.11e-19
C23808 VPWR.n2674 VGND 9.28e-19
C23809 VPWR.n2675 VGND 4.84e-19
C23810 VPWR.n2676 VGND 1.71e-19
C23811 VPWR.n2677 VGND 2.28e-19
C23812 VPWR.n2678 VGND 2.85e-19
C23813 VPWR.n2679 VGND 5.75e-19
C23814 VPWR.n2680 VGND 0.00259f
C23815 VPWR.t1574 VGND 0.00225f
C23816 VPWR.t3057 VGND 0.00166f
C23817 VPWR.n2681 VGND 0.00438f
C23818 VPWR.n2682 VGND 0.00608f
C23819 VPWR.t2786 VGND 0.00239f
C23820 VPWR.n2683 VGND 0.00411f
C23821 VPWR.n2684 VGND 4.13e-19
C23822 VPWR.n2685 VGND 0.00495f
C23823 VPWR.n2686 VGND 0.00524f
C23824 VPWR.n2687 VGND 0.00393f
C23825 VPWR.n2688 VGND 0.00199f
C23826 VPWR.n2689 VGND 0.0096f
C23827 VPWR.n2690 VGND 0.0182f
C23828 VPWR.t1571 VGND 0.023f
C23829 VPWR.t1567 VGND 0.0149f
C23830 VPWR.t3036 VGND 0.0144f
C23831 VPWR.t1573 VGND 0.03f
C23832 VPWR.t3056 VGND 0.0222f
C23833 VPWR.t2785 VGND 0.0111f
C23834 VPWR.t970 VGND 0.0237f
C23835 VPWR.t2440 VGND 0.0181f
C23836 VPWR.t3034 VGND 0.0144f
C23837 VPWR.t2446 VGND 0.0141f
C23838 VPWR.t2917 VGND 0.0144f
C23839 VPWR.t2448 VGND 0.0144f
C23840 VPWR.t2686 VGND 0.0144f
C23841 VPWR.t2438 VGND 0.0166f
C23842 VPWR.t2652 VGND 0.0144f
C23843 VPWR.t2444 VGND 0.0235f
C23844 VPWR.t2434 VGND 0.024f
C23845 VPWR.t994 VGND 0.0144f
C23846 VPWR.t2436 VGND 0.0163f
C23847 VPWR.t1735 VGND 0.0144f
C23848 VPWR.t2442 VGND 0.0173f
C23849 VPWR.t2452 VGND 0.0205f
C23850 VPWR.t2687 VGND 0.0144f
C23851 VPWR.t2454 VGND 0.0166f
C23852 VPWR.t2918 VGND 0.0144f
C23853 VPWR.t2450 VGND 0.0154f
C23854 VPWR.t1876 VGND 0.0144f
C23855 VPWR.t2462 VGND 0.0195f
C23856 VPWR.t2456 VGND 0.0289f
C23857 VPWR.t2458 VGND 0.0253f
C23858 VPWR.t2688 VGND 0.0144f
C23859 VPWR.t2460 VGND 0.0141f
C23860 VPWR.t1012 VGND 0.0144f
C23861 VPWR.t2464 VGND 0.0109f
C23862 VPWR.t1079 VGND 0.0218f
C23863 VPWR.t1071 VGND 0.0284f
C23864 VPWR.t264 VGND 0.0144f
C23865 VPWR.t1075 VGND 0.0149f
C23866 VPWR.t1077 VGND 0.0227f
C23867 VPWR.t2622 VGND 0.0126f
C23868 VPWR.t51 VGND 0.0164f
C23869 VPWR.t2494 VGND 0.0183f
C23870 VPWR.t2759 VGND 0.0126f
C23871 VPWR.t1809 VGND 0.0369f
C23872 VPWR.t1947 VGND 0.0211f
C23873 VPWR.t379 VGND 0.0144f
C23874 VPWR.t1507 VGND 0.024f
C23875 VPWR.t2961 VGND 0.0322f
C23876 VPWR.t2507 VGND 0.0272f
C23877 VPWR.t1785 VGND 0.0109f
C23878 VPWR.t3058 VGND 0.0218f
C23879 VPWR.t2905 VGND 0.03f
C23880 VPWR.t2907 VGND 0.0143f
C23881 VPWR.t2963 VGND 0.0208f
C23882 VPWR.t3119 VGND 0.0336f
C23883 VPWR.t3123 VGND 0.0218f
C23884 VPWR.t288 VGND 0.0141f
C23885 VPWR.t1248 VGND 0.0205f
C23886 VPWR.t1244 VGND 0.0282f
C23887 VPWR.t1250 VGND 0.0282f
C23888 VPWR.t1246 VGND 0.0282f
C23889 VPWR.t1240 VGND 0.0183f
C23890 VPWR.t1242 VGND 0.0151f
C23891 VPWR.t1459 VGND 0.0109f
C23892 VPWR.t3125 VGND 0.0121f
C23893 VPWR.t1399 VGND 0.0198f
C23894 VPWR.t1203 VGND 0.028f
C23895 VPWR.t3127 VGND 0.0258f
C23896 VPWR.t1988 VGND 0.0193f
C23897 VPWR.t1453 VGND 0.0183f
C23898 VPWR.t525 VGND 0.0163f
C23899 VPWR.t861 VGND 0.0228f
C23900 VPWR.t859 VGND 0.0222f
C23901 VPWR.n2691 VGND 0.0244f
C23902 VPWR.t628 VGND 0.0572f
C23903 VPWR.t2582 VGND 0.053f
C23904 VPWR.t2578 VGND 0.0282f
C23905 VPWR.t2574 VGND 0.0164f
C23906 VPWR.t116 VGND 0.0141f
C23907 VPWR.t2580 VGND 0.0258f
C23908 VPWR.t2584 VGND 0.0282f
C23909 VPWR.t2576 VGND 0.0282f
C23910 VPWR.t1984 VGND 0.0282f
C23911 VPWR.t1982 VGND 0.0279f
C23912 VPWR.t609 VGND 0.0621f
C23913 VPWR.t355 VGND 0.0262f
C23914 VPWR.t1907 VGND 0.0149f
C23915 VPWR.t1343 VGND 0.0319f
C23916 VPWR.t1495 VGND 0.0376f
C23917 VPWR.t1195 VGND 0.0363f
C23918 VPWR.t1117 VGND 0.0374f
C23919 VPWR.t2484 VGND 0.0287f
C23920 VPWR.t279 VGND 0.0264f
C23921 VPWR.t2331 VGND 0.0309f
C23922 VPWR.n2692 VGND 0.0334f
C23923 VPWR.n2693 VGND 0.00944f
C23924 VPWR.t2332 VGND 0.00549f
C23925 VPWR.t2760 VGND 0.00202f
C23926 VPWR.n2694 VGND 0.00345f
C23927 VPWR.n2695 VGND 0.00701f
C23928 VPWR.n2696 VGND 0.00949f
C23929 VPWR.n2697 VGND 0.00179f
C23930 VPWR.t356 VGND 0.0046f
C23931 VPWR.t2485 VGND 0.00267f
C23932 VPWR.t1118 VGND 0.00308f
C23933 VPWR.n2698 VGND 0.00622f
C23934 VPWR.n2699 VGND 0.00888f
C23935 VPWR.n2700 VGND 0.00184f
C23936 VPWR.n2701 VGND 0.00233f
C23937 VPWR.n2702 VGND 0.00393f
C23938 VPWR.n2703 VGND 0.00553f
C23939 VPWR.n2704 VGND 0.00524f
C23940 VPWR.n2705 VGND 0.00578f
C23941 VPWR.n2706 VGND 0.00524f
C23942 VPWR.t1196 VGND 0.00267f
C23943 VPWR.t1496 VGND 0.00267f
C23944 VPWR.n2707 VGND 0.00542f
C23945 VPWR.n2708 VGND 0.00651f
C23946 VPWR.n2709 VGND 0.00258f
C23947 VPWR.n2710 VGND 0.00524f
C23948 VPWR.t3383 VGND 0.0592f
C23949 VPWR.n2711 VGND 0.0356f
C23950 VPWR.n2712 VGND 0.00484f
C23951 VPWR.n2713 VGND 0.00524f
C23952 VPWR.n2714 VGND 0.0066f
C23953 VPWR.n2715 VGND 0.00524f
C23954 VPWR.n2716 VGND 0.00393f
C23955 VPWR.n2717 VGND 0.00199f
C23956 VPWR.n2718 VGND 0.00629f
C23957 VPWR.t610 VGND 0.00387f
C23958 VPWR.n2719 VGND 0.00612f
C23959 VPWR.n2720 VGND 0.00796f
C23960 VPWR.n2721 VGND 0.00393f
C23961 VPWR.n2722 VGND 0.00524f
C23962 VPWR.n2723 VGND 0.00524f
C23963 VPWR.n2724 VGND 0.0031f
C23964 VPWR.n2725 VGND 0.00182f
C23965 VPWR.n2726 VGND 0.00255f
C23966 VPWR.t117 VGND 0.0046f
C23967 VPWR.n2727 VGND 0.00285f
C23968 VPWR.n2728 VGND 0.00758f
C23969 VPWR.n2729 VGND 0.00452f
C23970 VPWR.n2730 VGND 0.00473f
C23971 VPWR.n2731 VGND 0.00506f
C23972 VPWR.n2732 VGND 0.00504f
C23973 VPWR.n2733 VGND 5.92e-19
C23974 VPWR.n2734 VGND 5.05e-19
C23975 VPWR.n2735 VGND 0.1f
C23976 VPWR.n2736 VGND 0.1f
C23977 VPWR.n2737 VGND 6.54e-19
C23978 VPWR.n2738 VGND 8.67e-19
C23979 VPWR.n2739 VGND 5.71e-19
C23980 VPWR.n2740 VGND 3.29e-19
C23981 VPWR.n2741 VGND 3.95e-19
C23982 VPWR.n2742 VGND 4.17e-19
C23983 VPWR.n2743 VGND 2.85e-19
C23984 VPWR.n2744 VGND 4.17e-19
C23985 VPWR.n2745 VGND 5.05e-19
C23986 VPWR.n2746 VGND 4.83e-19
C23987 VPWR.n2747 VGND 2.85e-19
C23988 VPWR.n2748 VGND 3.95e-19
C23989 VPWR.n2749 VGND 2.85e-19
C23990 VPWR.n2750 VGND 6.14e-19
C23991 VPWR.n2751 VGND 4.39e-19
C23992 VPWR.n2752 VGND 1.76e-19
C23993 VPWR.n2753 VGND 4.83e-19
C23994 VPWR.n2754 VGND 2.41e-19
C23995 VPWR.n2755 VGND 3.73e-19
C23996 VPWR.n2756 VGND 3.07e-19
C23997 VPWR.n2757 VGND 4.11e-19
C23998 VPWR.n2758 VGND 4.11e-19
C23999 VPWR.n2759 VGND 7.39e-19
C24000 VPWR.n2760 VGND 5.19e-19
C24001 VPWR.n2761 VGND 7.39e-19
C24002 VPWR.n2762 VGND 4.11e-19
C24003 VPWR.n2763 VGND 4.11e-19
C24004 VPWR.n2765 VGND 7.39e-19
C24005 VPWR.n2766 VGND 4.11e-19
C24006 VPWR.n2767 VGND 6.54e-19
C24007 VPWR.n2768 VGND 8.67e-19
C24008 VPWR.n2769 VGND 5.05e-19
C24009 VPWR.n2770 VGND 4.17e-19
C24010 VPWR.n2771 VGND 6.14e-19
C24011 VPWR.n2772 VGND 4.39e-19
C24012 VPWR.n2773 VGND 1.76e-19
C24013 VPWR.n2774 VGND 3.95e-19
C24014 VPWR.n2775 VGND 3.95e-19
C24015 VPWR.n2776 VGND 4.83e-19
C24016 VPWR.n2777 VGND 2.41e-19
C24017 VPWR.n2778 VGND 3.73e-19
C24018 VPWR.n2779 VGND 3.07e-19
C24019 VPWR.n2780 VGND 4.11e-19
C24020 VPWR.n2782 VGND 0.362f
C24021 VPWR.n2783 VGND 0.00138f
C24022 VPWR.n2784 VGND 0.00456f
C24023 VPWR.t2695 VGND 0.00676f
C24024 VPWR.n2785 VGND 0.0119f
C24025 VPWR.t3547 VGND 0.0592f
C24026 VPWR.n2786 VGND 0.0353f
C24027 VPWR.n2787 VGND 0.0019f
C24028 VPWR.t645 VGND 0.0046f
C24029 VPWR.n2788 VGND 0.00299f
C24030 VPWR.n2789 VGND 0.00282f
C24031 VPWR.t2518 VGND 6.73e-19
C24032 VPWR.t2817 VGND 9.96e-19
C24033 VPWR.n2790 VGND 0.00176f
C24034 VPWR.n2791 VGND 0.00421f
C24035 VPWR.n2792 VGND 0.00146f
C24036 VPWR.t153 VGND 0.0046f
C24037 VPWR.n2793 VGND 0.00407f
C24038 VPWR.n2794 VGND 0.00237f
C24039 VPWR.t71 VGND 0.00399f
C24040 VPWR.n2795 VGND 0.00683f
C24041 VPWR.n2796 VGND 0.00142f
C24042 VPWR.n2797 VGND 0.00393f
C24043 VPWR.n2798 VGND 0.00333f
C24044 VPWR.n2799 VGND 0.00175f
C24045 VPWR.t247 VGND 0.0046f
C24046 VPWR.n2800 VGND 0.00407f
C24047 VPWR.n2801 VGND 0.00269f
C24048 VPWR.n2802 VGND 0.00393f
C24049 VPWR.n2803 VGND 0.00639f
C24050 VPWR.n2804 VGND 0.00524f
C24051 VPWR.t1132 VGND 0.00234f
C24052 VPWR.n2805 VGND 0.00628f
C24053 VPWR.n2806 VGND 0.00398f
C24054 VPWR.n2807 VGND 0.00524f
C24055 VPWR.n2808 VGND 0.00438f
C24056 VPWR.n2809 VGND 0.00524f
C24057 VPWR.t3407 VGND 0.0592f
C24058 VPWR.n2810 VGND 0.0356f
C24059 VPWR.n2811 VGND 0.00484f
C24060 VPWR.n2812 VGND 0.00524f
C24061 VPWR.t1977 VGND 0.00102f
C24062 VPWR.t1762 VGND 0.00102f
C24063 VPWR.n2813 VGND 0.00217f
C24064 VPWR.n2814 VGND 0.0071f
C24065 VPWR.n2815 VGND 0.00337f
C24066 VPWR.n2816 VGND 0.00524f
C24067 VPWR.t70 VGND 0.00387f
C24068 VPWR.n2817 VGND 0.0107f
C24069 VPWR.n2818 VGND 0.00796f
C24070 VPWR.n2819 VGND 0.00622f
C24071 VPWR.n2820 VGND 0.0031f
C24072 VPWR.n2821 VGND 0.00393f
C24073 VPWR.t3558 VGND 0.0231f
C24074 VPWR.n2822 VGND 0.043f
C24075 VPWR.n2823 VGND 0.00524f
C24076 VPWR.n2824 VGND 0.00524f
C24077 VPWR.n2825 VGND 0.00524f
C24078 VPWR.n2826 VGND 0.0185f
C24079 VPWR.n2827 VGND 0.0179f
C24080 VPWR.t248 VGND 0.0046f
C24081 VPWR.n2828 VGND 0.01f
C24082 VPWR.n2829 VGND 0.011f
C24083 VPWR.n2830 VGND 0.0031f
C24084 VPWR.n2831 VGND 0.00262f
C24085 VPWR.n2832 VGND 0.00432f
C24086 VPWR.t1255 VGND 0.00676f
C24087 VPWR.n2833 VGND 0.00899f
C24088 VPWR.t152 VGND 0.0046f
C24089 VPWR.n2834 VGND 0.00407f
C24090 VPWR.n2835 VGND 0.00194f
C24091 VPWR.n2836 VGND 0.00393f
C24092 VPWR.t2971 VGND 0.00239f
C24093 VPWR.n2837 VGND 0.00658f
C24094 VPWR.n2838 VGND 0.00434f
C24095 VPWR.n2839 VGND 0.00524f
C24096 VPWR.n2840 VGND 0.00535f
C24097 VPWR.n2841 VGND 0.00524f
C24098 VPWR.t2528 VGND 6.73e-19
C24099 VPWR.t1257 VGND 0.00127f
C24100 VPWR.n2842 VGND 0.00203f
C24101 VPWR.n2843 VGND 0.0044f
C24102 VPWR.n2844 VGND 0.00377f
C24103 VPWR.n2845 VGND 0.00524f
C24104 VPWR.t3582 VGND 0.0592f
C24105 VPWR.n2846 VGND 0.0351f
C24106 VPWR.n2847 VGND 0.00484f
C24107 VPWR.n2848 VGND 0.00524f
C24108 VPWR.n2849 VGND 0.0066f
C24109 VPWR.n2850 VGND 0.00524f
C24110 VPWR.n2851 VGND 0.0066f
C24111 VPWR.n2852 VGND 0.00524f
C24112 VPWR.t1450 VGND 0.00453f
C24113 VPWR.n2853 VGND 0.00799f
C24114 VPWR.n2854 VGND 0.00438f
C24115 VPWR.n2855 VGND 0.00524f
C24116 VPWR.n2856 VGND 0.00553f
C24117 VPWR.n2857 VGND 0.00524f
C24118 VPWR.t2522 VGND 6.73e-19
C24119 VPWR.t926 VGND 9.96e-19
C24120 VPWR.n2858 VGND 0.00176f
C24121 VPWR.n2859 VGND 0.00658f
C24122 VPWR.n2860 VGND 0.00484f
C24123 VPWR.n2861 VGND 0.00524f
C24124 VPWR.n2862 VGND 0.00484f
C24125 VPWR.n2863 VGND 0.00524f
C24126 VPWR.n2864 VGND 0.0031f
C24127 VPWR.n2865 VGND 0.00138f
C24128 VPWR.n2866 VGND 1.71e-19
C24129 VPWR.n2867 VGND 3.95e-19
C24130 VPWR.n2868 VGND 5.27e-19
C24131 VPWR.n2869 VGND 4.61e-19
C24132 VPWR.n2870 VGND 0.00138f
C24133 VPWR.n2871 VGND 5.05e-19
C24134 VPWR.n2872 VGND 5.05e-19
C24135 VPWR.n2873 VGND 3.07e-19
C24136 VPWR.n2874 VGND 4.31e-19
C24137 VPWR.n2875 VGND 4.5e-19
C24138 VPWR.n2876 VGND 5.74e-19
C24139 VPWR.n2877 VGND 6.54e-19
C24140 VPWR.n2878 VGND 8.67e-19
C24141 VPWR.n2879 VGND 0.0976f
C24142 VPWR.n2880 VGND 0.00389f
C24143 VPWR.n2881 VGND 4.11e-19
C24144 VPWR.n2882 VGND 8.67e-19
C24145 VPWR.n2883 VGND 4.11e-19
C24146 VPWR.n2884 VGND 0.00138f
C24147 VPWR.n2885 VGND 9e-19
C24148 VPWR.t341 VGND 0.0046f
C24149 VPWR.t622 VGND 0.00387f
C24150 VPWR.n2886 VGND 0.0115f
C24151 VPWR.t683 VGND 0.0046f
C24152 VPWR.t214 VGND 0.0046f
C24153 VPWR.n2887 VGND 0.011f
C24154 VPWR.n2888 VGND 0.00721f
C24155 VPWR.t684 VGND 0.0046f
C24156 VPWR.t215 VGND 0.0046f
C24157 VPWR.n2889 VGND 0.00721f
C24158 VPWR.t3490 VGND 0.00911f
C24159 VPWR.t473 VGND 0.00391f
C24160 VPWR.n2890 VGND 0.0253f
C24161 VPWR.t472 VGND 0.00391f
C24162 VPWR.n2892 VGND 0.0138f
C24163 VPWR.n2893 VGND 0.00548f
C24164 VPWR.t3349 VGND 0.00911f
C24165 VPWR.t217 VGND 0.00391f
C24166 VPWR.n2894 VGND 0.0253f
C24167 VPWR.t218 VGND 0.00391f
C24168 VPWR.n2896 VGND 0.0138f
C24169 VPWR.n2897 VGND 0.0112f
C24170 VPWR.n2898 VGND 0.00403f
C24171 VPWR.n2899 VGND 0.0031f
C24172 VPWR.n2900 VGND 0.011f
C24173 VPWR.n2901 VGND 0.00524f
C24174 VPWR.n2902 VGND 0.0113f
C24175 VPWR.n2903 VGND 0.00524f
C24176 VPWR.n2904 VGND 0.0113f
C24177 VPWR.n2905 VGND 0.00524f
C24178 VPWR.n2906 VGND 0.0113f
C24179 VPWR.n2907 VGND 0.00524f
C24180 VPWR.n2908 VGND 0.0113f
C24181 VPWR.n2909 VGND 0.00524f
C24182 VPWR.n2910 VGND 0.0113f
C24183 VPWR.n2911 VGND 0.00524f
C24184 VPWR.t3389 VGND 0.0592f
C24185 VPWR.t3510 VGND 0.0592f
C24186 VPWR.n2912 VGND 0.0703f
C24187 VPWR.n2913 VGND 0.00833f
C24188 VPWR.n2914 VGND 0.00524f
C24189 VPWR.n2915 VGND 0.0087f
C24190 VPWR.n2916 VGND 0.00524f
C24191 VPWR.n2917 VGND 0.0113f
C24192 VPWR.n2918 VGND 0.00524f
C24193 VPWR.n2919 VGND 0.00524f
C24194 VPWR.n2920 VGND 0.00393f
C24195 VPWR.n2921 VGND 0.00418f
C24196 VPWR.n2922 VGND 0.00679f
C24197 VPWR.n2923 VGND 0.0031f
C24198 VPWR.n2924 VGND 0.0179f
C24199 VPWR.n2925 VGND 0.00524f
C24200 VPWR.n2926 VGND 0.0185f
C24201 VPWR.n2927 VGND 0.00524f
C24202 VPWR.n2928 VGND 0.0185f
C24203 VPWR.n2929 VGND 0.00524f
C24204 VPWR.t3532 VGND 0.0231f
C24205 VPWR.n2930 VGND 0.00708f
C24206 VPWR.n2931 VGND 9.04e-19
C24207 VPWR.t621 VGND 0.00387f
C24208 VPWR.n2932 VGND 0.0029f
C24209 VPWR.n2933 VGND 0.00865f
C24210 VPWR.n2934 VGND 0.0421f
C24211 VPWR.n2935 VGND 0.00387f
C24212 VPWR.n2936 VGND 8.83e-19
C24213 VPWR.n2937 VGND 0.00273f
C24214 VPWR.n2938 VGND 9.68e-19
C24215 VPWR.n2939 VGND 4.27e-19
C24216 VPWR.n2940 VGND 2.56e-19
C24217 VPWR.n2941 VGND 6.1e-19
C24218 VPWR.n2942 VGND 0.00289f
C24219 VPWR.n2943 VGND 3.42e-19
C24220 VPWR.n2944 VGND 4.83e-19
C24221 VPWR.n2945 VGND 4.17e-19
C24222 VPWR.n2946 VGND 5.71e-19
C24223 VPWR.n2947 VGND 6.26e-19
C24224 VPWR.n2948 VGND 1.99e-19
C24225 VPWR.n2949 VGND 4.17e-19
C24226 VPWR.n2950 VGND 4.39e-19
C24227 VPWR.n2951 VGND 3.29e-19
C24228 VPWR.n2952 VGND 5.27e-19
C24229 VPWR.n2953 VGND 2.85e-19
C24230 VPWR.n2954 VGND 2.85e-19
C24231 VPWR.n2955 VGND 4.17e-19
C24232 VPWR.n2956 VGND 4.61e-19
C24233 VPWR.n2957 VGND 3.51e-19
C24234 VPWR.n2958 VGND 5.12e-19
C24235 VPWR.n2959 VGND 5.41e-19
C24236 VPWR.n2960 VGND 3.7e-19
C24237 VPWR.n2961 VGND 6.83e-19
C24238 VPWR.n2962 VGND 4.27e-19
C24239 VPWR.n2963 VGND 8.54e-20
C24240 VPWR.n2964 VGND 4.27e-19
C24241 VPWR.n2965 VGND 0.00156f
C24242 VPWR.n2966 VGND 0.00203f
C24243 VPWR.n2967 VGND 0.00138f
C24244 VPWR.n2968 VGND 6.14e-19
C24245 VPWR.n2969 VGND 4.31e-19
C24246 VPWR.n2970 VGND 6.54e-19
C24247 VPWR.n2971 VGND 7.02e-19
C24248 VPWR.n2972 VGND 3.21e-19
C24249 VPWR.n2973 VGND 0.0173f
C24250 VPWR.n2974 VGND 0.365f
C24251 VPWR.n2975 VGND 0.365f
C24252 VPWR.n2976 VGND 0.0166f
C24253 VPWR.n2977 VGND 0.187f
C24254 VPWR.n2978 VGND 9.06e-19
C24255 VPWR.n2979 VGND 9e-19
C24256 VPWR.n2980 VGND 0.00138f
C24257 VPWR.n2981 VGND 6.14e-19
C24258 VPWR.n2982 VGND 5.48e-19
C24259 VPWR.n2983 VGND 0.00138f
C24260 VPWR.n2984 VGND 0.0562f
C24261 VPWR.n2985 VGND 0.00139f
C24262 VPWR.n2986 VGND 8.67e-19
C24263 VPWR.n2987 VGND 6.54e-19
C24264 VPWR.n2988 VGND 9.06e-19
C24265 VPWR.t147 VGND 0.00396f
C24266 VPWR.n2989 VGND 0.0107f
C24267 VPWR.n2990 VGND 0.00944f
C24268 VPWR.t3384 VGND 0.00911f
C24269 VPWR.t105 VGND 0.00391f
C24270 VPWR.n2991 VGND 0.0253f
C24271 VPWR.t106 VGND 0.00391f
C24272 VPWR.n2993 VGND 0.0126f
C24273 VPWR.t1891 VGND 0.00631f
C24274 VPWR.n2994 VGND 0.00646f
C24275 VPWR.n2995 VGND 0.00219f
C24276 VPWR.t1889 VGND 0.00645f
C24277 VPWR.t777 VGND 0.00643f
C24278 VPWR.t556 VGND 0.0046f
C24279 VPWR.n2996 VGND 0.00644f
C24280 VPWR.t366 VGND 0.00398f
C24281 VPWR.n2997 VGND 0.0163f
C24282 VPWR.n2998 VGND 0.0177f
C24283 VPWR.n2999 VGND 6.26e-19
C24284 VPWR.n3000 VGND 3.95e-19
C24285 VPWR.n3001 VGND 7.68e-19
C24286 VPWR.n3002 VGND 5.05e-19
C24287 VPWR.n3003 VGND 9.06e-19
C24288 VPWR.n3004 VGND 0.0562f
C24289 VPWR.n3006 VGND 0.00934f
C24290 VPWR.n3007 VGND 0.0963f
C24291 VPWR.n3008 VGND 0.0952f
C24292 VPWR.n3009 VGND 3.95e-19
C24293 VPWR.n3010 VGND 4.17e-19
C24294 VPWR.n3011 VGND 2.85e-19
C24295 VPWR.n3012 VGND 4.83e-19
C24296 VPWR.n3013 VGND 2.85e-19
C24297 VPWR.n3014 VGND 3.95e-19
C24298 VPWR.n3015 VGND 2.85e-19
C24299 VPWR.n3016 VGND 4.11e-19
C24300 VPWR.n3017 VGND 4.11e-19
C24301 VPWR.n3018 VGND 7.39e-19
C24302 VPWR.n3019 VGND 5.19e-19
C24303 VPWR.n3020 VGND 7.39e-19
C24304 VPWR.n3021 VGND 4.11e-19
C24305 VPWR.n3022 VGND 5.05e-19
C24306 VPWR.n3023 VGND 4.17e-19
C24307 VPWR.n3024 VGND 6.14e-19
C24308 VPWR.n3025 VGND 4.39e-19
C24309 VPWR.n3026 VGND 1.76e-19
C24310 VPWR.t183 VGND 0.00462f
C24311 VPWR.n3027 VGND 0.0093f
C24312 VPWR.t3393 VGND 0.00911f
C24313 VPWR.t129 VGND 0.00391f
C24314 VPWR.n3028 VGND 0.0253f
C24315 VPWR.t130 VGND 0.00391f
C24316 VPWR.n3030 VGND 0.0138f
C24317 VPWR.n3031 VGND 0.00854f
C24318 VPWR.t182 VGND 0.00463f
C24319 VPWR.t299 VGND 0.004f
C24320 VPWR.n3032 VGND 0.00482f
C24321 VPWR.t3454 VGND 0.0182f
C24322 VPWR.t298 VGND 0.00387f
C24323 VPWR.n3033 VGND 0.0244f
C24324 VPWR.n3034 VGND 0.0153f
C24325 VPWR.n3035 VGND 0.00859f
C24326 VPWR.n3036 VGND 0.0125f
C24327 VPWR.t97 VGND 0.00398f
C24328 VPWR.n3037 VGND 0.007f
C24329 VPWR.n3038 VGND 0.0345f
C24330 VPWR.n3039 VGND 0.00123f
C24331 VPWR.n3040 VGND 0.00123f
C24332 VPWR.t1642 VGND 0.00136f
C24333 VPWR.t787 VGND 0.00136f
C24334 VPWR.n3041 VGND 0.00328f
C24335 VPWR.n3042 VGND 0.00789f
C24336 VPWR.t666 VGND 0.0046f
C24337 VPWR.t2164 VGND 0.00261f
C24338 VPWR.n3043 VGND 0.00794f
C24339 VPWR.t90 VGND 0.00387f
C24340 VPWR.t3353 VGND 0.0282f
C24341 VPWR.n3044 VGND 0.0137f
C24342 VPWR.n3045 VGND 0.0512f
C24343 VPWR.n3046 VGND 0.0135f
C24344 VPWR.n3047 VGND 0.0107f
C24345 VPWR.n3048 VGND 0.00796f
C24346 VPWR.t667 VGND 0.0046f
C24347 VPWR.n3049 VGND 0.01f
C24348 VPWR.t2392 VGND 0.00643f
C24349 VPWR.n3050 VGND 0.0132f
C24350 VPWR.t3208 VGND 0.00651f
C24351 VPWR.t2390 VGND -2.18e-20
C24352 VPWR.t3183 VGND 0.00137f
C24353 VPWR.n3051 VGND 0.00618f
C24354 VPWR.n3052 VGND 0.0119f
C24355 VPWR.t91 VGND 0.00387f
C24356 VPWR.n3053 VGND 0.00202f
C24357 VPWR.n3054 VGND 0.00499f
C24358 VPWR.n3055 VGND 0.00813f
C24359 VPWR.t3204 VGND 0.00631f
C24360 VPWR.t3408 VGND 0.00911f
C24361 VPWR.t254 VGND 0.00391f
C24362 VPWR.n3056 VGND 0.0253f
C24363 VPWR.t253 VGND 0.00391f
C24364 VPWR.n3058 VGND 0.0126f
C24365 VPWR.n3059 VGND 0.0115f
C24366 VPWR.n3060 VGND 0.00262f
C24367 VPWR.n3061 VGND 0.0117f
C24368 VPWR.t3357 VGND 0.0289f
C24369 VPWR.t96 VGND 0.00387f
C24370 VPWR.n3062 VGND 0.0547f
C24371 VPWR.n3063 VGND 0.0106f
C24372 VPWR.n3064 VGND 0.0167f
C24373 VPWR.t3525 VGND 0.0289f
C24374 VPWR.t490 VGND 0.00387f
C24375 VPWR.n3065 VGND 0.0604f
C24376 VPWR.n3066 VGND 0.0212f
C24377 VPWR.t491 VGND 0.00398f
C24378 VPWR.n3067 VGND 0.0317f
C24379 VPWR.n3068 VGND 0.0172f
C24380 VPWR.n3069 VGND 0.00618f
C24381 VPWR.n3070 VGND 0.00442f
C24382 VPWR.n3071 VGND 0.00996f
C24383 VPWR.n3072 VGND 0.00131f
C24384 VPWR.n3073 VGND 0.00199f
C24385 VPWR.n3074 VGND 0.00179f
C24386 VPWR.n3075 VGND 0.0031f
C24387 VPWR.n3076 VGND 0.00524f
C24388 VPWR.n3077 VGND 0.00475f
C24389 VPWR.n3078 VGND 0.00702f
C24390 VPWR.n3079 VGND 0.0136f
C24391 VPWR.n3080 VGND 0.00904f
C24392 VPWR.n3081 VGND 0.0031f
C24393 VPWR.n3082 VGND 0.0179f
C24394 VPWR.n3083 VGND 0.00524f
C24395 VPWR.n3084 VGND 0.00524f
C24396 VPWR.n3085 VGND 0.00524f
C24397 VPWR.n3086 VGND 0.00393f
C24398 VPWR.n3087 VGND 0.00199f
C24399 VPWR.n3088 VGND 0.00629f
C24400 VPWR.n3089 VGND 0.0047f
C24401 VPWR.n3090 VGND 0.00288f
C24402 VPWR.n3091 VGND 5.92e-19
C24403 VPWR.n3092 VGND 5.05e-19
C24404 VPWR.n3093 VGND 9.06e-19
C24405 VPWR.n3094 VGND 0.0562f
C24406 VPWR.n3095 VGND 0.00139f
C24407 VPWR.n3096 VGND 8.67e-19
C24408 VPWR.n3097 VGND 6.54e-19
C24409 VPWR.n3098 VGND 9.06e-19
C24410 VPWR.n3099 VGND 8.11e-19
C24411 VPWR.n3100 VGND 3.95e-19
C24412 VPWR.n3101 VGND 1.76e-19
C24413 VPWR.n3102 VGND 3.95e-19
C24414 VPWR.n3103 VGND 3.95e-19
C24415 VPWR.n3104 VGND 7.68e-19
C24416 VPWR.n3105 VGND 5.05e-19
C24417 VPWR.n3106 VGND 1.76e-19
C24418 VPWR.n3107 VGND 5.48e-19
C24419 VPWR.n3109 VGND 0.0976f
C24420 VPWR.n3110 VGND 0.00389f
C24421 VPWR.n3112 VGND 0.00138f
C24422 VPWR.n3113 VGND 8.11e-19
C24423 VPWR.n3114 VGND 3.95e-19
C24424 VPWR.n3115 VGND 1.76e-19
C24425 VPWR.n3116 VGND 7.68e-19
C24426 VPWR.n3117 VGND 5.05e-19
C24427 VPWR.n3118 VGND 1.76e-19
C24428 VPWR.n3119 VGND 4.31e-19
C24429 VPWR.n3120 VGND 4.5e-19
C24430 VPWR.n3121 VGND 6.54e-19
C24431 VPWR.n3122 VGND 7.02e-19
C24432 VPWR.n3123 VGND 3.21e-19
C24433 VPWR.n3124 VGND 0.367f
C24434 VPWR.n3125 VGND 0.0173f
C24435 VPWR.n3126 VGND 0.0976f
C24436 VPWR.n3127 VGND 0.00389f
C24437 VPWR.n3129 VGND 0.00139f
C24438 VPWR.n3130 VGND 0.00138f
C24439 VPWR.n3131 VGND 9e-19
C24440 VPWR.n3132 VGND 6.14e-19
C24441 VPWR.n3133 VGND 6.54e-19
C24442 VPWR.n3134 VGND 9.06e-19
C24443 VPWR.n3135 VGND 5.48e-19
C24444 VPWR.n3136 VGND 8.67e-19
C24445 VPWR.n3137 VGND 6.54e-19
C24446 VPWR.n3138 VGND 9.06e-19
C24447 VPWR.n3139 VGND 3.73e-19
C24448 VPWR.n3140 VGND 5.27e-19
C24449 VPWR.n3141 VGND 3.95e-19
C24450 VPWR.n3142 VGND 5.05e-19
C24451 VPWR.n3143 VGND 5.05e-19
C24452 VPWR.t171 VGND 0.0046f
C24453 VPWR.n3144 VGND 0.004f
C24454 VPWR.t1716 VGND -2.18e-20
C24455 VPWR.t1469 VGND 0.00137f
C24456 VPWR.n3145 VGND 0.00618f
C24457 VPWR.n3146 VGND 0.00587f
C24458 VPWR.t3522 VGND 0.00911f
C24459 VPWR.t590 VGND 0.00391f
C24460 VPWR.n3147 VGND 0.0253f
C24461 VPWR.t589 VGND 0.00391f
C24462 VPWR.n3149 VGND 0.0138f
C24463 VPWR.t3358 VGND 0.0597f
C24464 VPWR.t149 VGND 0.0046f
C24465 VPWR.n3150 VGND 0.011f
C24466 VPWR.n3151 VGND 0.00644f
C24467 VPWR.t100 VGND 0.0046f
C24468 VPWR.n3152 VGND 0.00644f
C24469 VPWR.t150 VGND 0.0046f
C24470 VPWR.n3153 VGND 0.00407f
C24471 VPWR.n3154 VGND 0.00135f
C24472 VPWR.t829 VGND 0.00651f
C24473 VPWR.n3155 VGND 0.0082f
C24474 VPWR.t1999 VGND 0.00166f
C24475 VPWR.t2097 VGND 0.00166f
C24476 VPWR.n3156 VGND 0.0037f
C24477 VPWR.t1156 VGND 0.00137f
C24478 VPWR.t3004 VGND -2.18e-20
C24479 VPWR.n3157 VGND 0.00618f
C24480 VPWR.n3158 VGND 0.00641f
C24481 VPWR.n3159 VGND 0.00525f
C24482 VPWR.t3002 VGND 0.00663f
C24483 VPWR.n3160 VGND 0.00878f
C24484 VPWR.t1840 VGND 0.00598f
C24485 VPWR.n3161 VGND 0.00834f
C24486 VPWR.n3162 VGND 0.0031f
C24487 VPWR.n3163 VGND 0.00393f
C24488 VPWR.n3164 VGND 0.00393f
C24489 VPWR.n3165 VGND 0.00154f
C24490 VPWR.n3166 VGND 0.00524f
C24491 VPWR.n3167 VGND 0.00475f
C24492 VPWR.n3168 VGND 9.48e-19
C24493 VPWR.n3169 VGND 0.00164f
C24494 VPWR.n3170 VGND 0.00179f
C24495 VPWR.n3171 VGND 0.0031f
C24496 VPWR.n3172 VGND 0.00393f
C24497 VPWR.n3173 VGND 0.00262f
C24498 VPWR.t831 VGND 0.0065f
C24499 VPWR.n3174 VGND 0.00756f
C24500 VPWR.n3175 VGND 0.00253f
C24501 VPWR.n3176 VGND 0.0031f
C24502 VPWR.t797 VGND 0.00102f
C24503 VPWR.t2587 VGND 0.00154f
C24504 VPWR.n3177 VGND 0.00483f
C24505 VPWR.n3178 VGND 0.00908f
C24506 VPWR.n3179 VGND 0.00423f
C24507 VPWR.n3180 VGND 0.00524f
C24508 VPWR.n3181 VGND 0.00545f
C24509 VPWR.n3182 VGND 0.00524f
C24510 VPWR.n3183 VGND 0.00475f
C24511 VPWR.n3184 VGND 0.00642f
C24512 VPWR.n3185 VGND 0.00535f
C24513 VPWR.n3186 VGND 0.0031f
C24514 VPWR.n3187 VGND 0.011f
C24515 VPWR.n3188 VGND 0.00524f
C24516 VPWR.n3189 VGND 0.0113f
C24517 VPWR.n3190 VGND 0.00524f
C24518 VPWR.t3397 VGND 0.0592f
C24519 VPWR.n3191 VGND 0.038f
C24520 VPWR.n3192 VGND 0.00833f
C24521 VPWR.n3193 VGND 0.00524f
C24522 VPWR.n3194 VGND 0.0087f
C24523 VPWR.n3195 VGND 0.00524f
C24524 VPWR.n3196 VGND 0.0113f
C24525 VPWR.n3197 VGND 0.00524f
C24526 VPWR.n3198 VGND 0.00524f
C24527 VPWR.n3199 VGND 0.00393f
C24528 VPWR.n3200 VGND 0.00396f
C24529 VPWR.n3201 VGND 0.034f
C24530 VPWR.n3202 VGND 0.0055f
C24531 VPWR.n3203 VGND 0.00333f
C24532 VPWR.n3204 VGND 0.00393f
C24533 VPWR.n3205 VGND 0.0066f
C24534 VPWR.n3206 VGND 0.00639f
C24535 VPWR.n3207 VGND 0.0031f
C24536 VPWR.t99 VGND 0.0046f
C24537 VPWR.n3208 VGND 0.00407f
C24538 VPWR.n3209 VGND 0.00196f
C24539 VPWR.n3210 VGND 0.00393f
C24540 VPWR.n3211 VGND 0.00281f
C24541 VPWR.n3212 VGND 0.00199f
C24542 VPWR.t1718 VGND 0.00643f
C24543 VPWR.t154 VGND 0.053f
C24544 VPWR.t2735 VGND 0.054f
C24545 VPWR.t187 VGND 0.0144f
C24546 VPWR.t2737 VGND 0.0153f
C24547 VPWR.t2731 VGND 0.0252f
C24548 VPWR.t2733 VGND 0.0198f
C24549 VPWR.t3073 VGND 0.017f
C24550 VPWR.t3178 VGND 0.0111f
C24551 VPWR.t2588 VGND 0.0151f
C24552 VPWR.t3273 VGND 0.0211f
C24553 VPWR.t1441 VGND 0.0297f
C24554 VPWR.t1439 VGND 0.0205f
C24555 VPWR.t3143 VGND 0.0159f
C24556 VPWR.t2794 VGND 0.0141f
C24557 VPWR.t962 VGND 0.0109f
C24558 VPWR.t3271 VGND 0.0258f
C24559 VPWR.t2818 VGND 0.0163f
C24560 VPWR.t282 VGND 0.0144f
C24561 VPWR.t1276 VGND 0.0183f
C24562 VPWR.t1141 VGND 0.0436f
C24563 VPWR.t964 VGND 0.0493f
C24564 VPWR.t1903 VGND 0.0398f
C24565 VPWR.t1277 VGND 0.0376f
C24566 VPWR.t169 VGND 0.0166f
C24567 VPWR.t2819 VGND 0.018f
C24568 VPWR.t2925 VGND 0.0603f
C24569 VPWR.t1274 VGND 0.0589f
C24570 VPWR.t1020 VGND 0.025f
C24571 VPWR.t1839 VGND 0.042f
C24572 VPWR.t3001 VGND 0.0316f
C24573 VPWR.t795 VGND 0.0141f
C24574 VPWR.t3003 VGND 0.0143f
C24575 VPWR.t2096 VGND 0.0154f
C24576 VPWR.t1998 VGND 0.0149f
C24577 VPWR.t1155 VGND 0.00571f
C24578 VPWR.t828 VGND 0.0253f
C24579 VPWR.t830 VGND 0.0196f
C24580 VPWR.t2100 VGND 0.0144f
C24581 VPWR.t796 VGND 0.0284f
C24582 VPWR.t2586 VGND 0.0473f
C24583 VPWR.t148 VGND 0.0878f
C24584 VPWR.t98 VGND 0.0973f
C24585 VPWR.t1468 VGND 0.0269f
C24586 VPWR.t1715 VGND 0.02f
C24587 VPWR.t1717 VGND 0.0183f
C24588 VPWR.t588 VGND 0.0237f
C24589 VPWR.n3213 VGND 0.0315f
C24590 VPWR.n3214 VGND 0.0162f
C24591 VPWR.n3215 VGND 0.00788f
C24592 VPWR.n3216 VGND 0.00237f
C24593 VPWR.n3217 VGND 0.0031f
C24594 VPWR.t1275 VGND 0.00102f
C24595 VPWR.t1021 VGND 0.00102f
C24596 VPWR.n3218 VGND 0.00217f
C24597 VPWR.n3219 VGND 0.00688f
C24598 VPWR.n3220 VGND 0.00337f
C24599 VPWR.n3221 VGND 0.00524f
C24600 VPWR.n3222 VGND 0.0066f
C24601 VPWR.n3223 VGND 0.00524f
C24602 VPWR.n3224 VGND 0.00592f
C24603 VPWR.n3225 VGND 0.00524f
C24604 VPWR.t2926 VGND 0.00234f
C24605 VPWR.n3226 VGND 0.00628f
C24606 VPWR.n3227 VGND 0.00398f
C24607 VPWR.n3228 VGND 0.00524f
C24608 VPWR.n3229 VGND 0.0066f
C24609 VPWR.n3230 VGND 0.00524f
C24610 VPWR.n3231 VGND 0.00632f
C24611 VPWR.n3232 VGND 0.00449f
C24612 VPWR.t284 VGND 0.00391f
C24613 VPWR.n3233 VGND 0.00833f
C24614 VPWR.t3274 VGND 0.00692f
C24615 VPWR.t1442 VGND 0.0066f
C24616 VPWR.n3234 VGND 0.00152f
C24617 VPWR.t2734 VGND 0.00225f
C24618 VPWR.t3074 VGND 0.00166f
C24619 VPWR.n3235 VGND 0.0045f
C24620 VPWR.t2738 VGND 0.00166f
C24621 VPWR.t2732 VGND 0.00166f
C24622 VPWR.n3236 VGND 0.00341f
C24623 VPWR.t3414 VGND 0.0179f
C24624 VPWR.n3237 VGND 0.017f
C24625 VPWR.n3238 VGND 0.0103f
C24626 VPWR.n3239 VGND 0.00702f
C24627 VPWR.n3240 VGND 0.00912f
C24628 VPWR.t189 VGND 0.00387f
C24629 VPWR.n3241 VGND 0.00822f
C24630 VPWR.t3371 VGND 0.00911f
C24631 VPWR.t156 VGND 0.00391f
C24632 VPWR.n3242 VGND 0.0253f
C24633 VPWR.t155 VGND 0.00391f
C24634 VPWR.n3244 VGND 0.0138f
C24635 VPWR.n3245 VGND 0.00345f
C24636 VPWR.t3476 VGND 0.00911f
C24637 VPWR.t342 VGND 0.00391f
C24638 VPWR.n3246 VGND 0.0253f
C24639 VPWR.t343 VGND 0.00391f
C24640 VPWR.n3248 VGND 0.0138f
C24641 VPWR.n3249 VGND 0.0112f
C24642 VPWR.t188 VGND 0.00387f
C24643 VPWR.t2736 VGND 0.00682f
C24644 VPWR.n3250 VGND 0.00917f
C24645 VPWR.n3251 VGND 0.00232f
C24646 VPWR.n3252 VGND 0.00487f
C24647 VPWR.n3253 VGND 0.00393f
C24648 VPWR.n3254 VGND 0.00524f
C24649 VPWR.n3255 VGND 0.00524f
C24650 VPWR.n3256 VGND 0.0031f
C24651 VPWR.n3257 VGND 0.00473f
C24652 VPWR.n3258 VGND 0.00747f
C24653 VPWR.n3259 VGND 0.00393f
C24654 VPWR.t3179 VGND 0.00136f
C24655 VPWR.t2589 VGND 0.00136f
C24656 VPWR.n3260 VGND 0.00328f
C24657 VPWR.n3261 VGND 0.00765f
C24658 VPWR.n3262 VGND 0.0031f
C24659 VPWR.n3263 VGND 0.00179f
C24660 VPWR.n3264 VGND 0.00199f
C24661 VPWR.n3265 VGND 0.0015f
C24662 VPWR.n3266 VGND 0.0177f
C24663 VPWR.n3267 VGND 0.00393f
C24664 VPWR.t3144 VGND 0.00239f
C24665 VPWR.n3268 VGND 0.00414f
C24666 VPWR.n3269 VGND 0.00102f
C24667 VPWR.n3270 VGND 0.00524f
C24668 VPWR.t1440 VGND -2.18e-20
C24669 VPWR.t2795 VGND 0.00137f
C24670 VPWR.n3271 VGND 0.00618f
C24671 VPWR.n3272 VGND 0.00607f
C24672 VPWR.n3273 VGND 8.77e-19
C24673 VPWR.n3274 VGND 0.00524f
C24674 VPWR.t283 VGND 0.00391f
C24675 VPWR.t3452 VGND 0.00886f
C24676 VPWR.n3275 VGND 0.0116f
C24677 VPWR.n3276 VGND 0.0146f
C24678 VPWR.n3277 VGND 0.00317f
C24679 VPWR.n3278 VGND 0.00471f
C24680 VPWR.t963 VGND 6.73e-19
C24681 VPWR.t3272 VGND 0.00127f
C24682 VPWR.n3279 VGND 0.00207f
C24683 VPWR.n3280 VGND 0.00499f
C24684 VPWR.n3281 VGND 0.0031f
C24685 VPWR.n3282 VGND 0.00393f
C24686 VPWR.n3283 VGND 0.00524f
C24687 VPWR.n3284 VGND 0.0031f
C24688 VPWR.n3285 VGND 0.00515f
C24689 VPWR.t170 VGND 0.0046f
C24690 VPWR.t1142 VGND 0.00453f
C24691 VPWR.n3286 VGND 0.00778f
C24692 VPWR.n3287 VGND 0.00184f
C24693 VPWR.n3288 VGND 0.00256f
C24694 VPWR.n3289 VGND 0.00393f
C24695 VPWR.n3290 VGND 0.00506f
C24696 VPWR.n3291 VGND 0.0039f
C24697 VPWR.n3292 VGND 0.00206f
C24698 VPWR.n3293 VGND 0.0033f
C24699 VPWR.n3294 VGND 0.00153f
C24700 VPWR.n3295 VGND 6.1e-19
C24701 VPWR.n3296 VGND 4.27e-19
C24702 VPWR.n3297 VGND 1.14e-19
C24703 VPWR.t965 VGND 6.73e-19
C24704 VPWR.t1904 VGND 9.96e-19
C24705 VPWR.n3298 VGND 0.00176f
C24706 VPWR.n3299 VGND 0.0064f
C24707 VPWR.n3300 VGND 0.00154f
C24708 VPWR.n3301 VGND 4.27e-19
C24709 VPWR.n3302 VGND 6.83e-19
C24710 VPWR.n3303 VGND 3.7e-19
C24711 VPWR.n3304 VGND 9.68e-19
C24712 VPWR.n3305 VGND 9.96e-19
C24713 VPWR.n3306 VGND 5.41e-19
C24714 VPWR.n3307 VGND 7.4e-19
C24715 VPWR.n3308 VGND 6.1e-19
C24716 VPWR.n3309 VGND 0.00176f
C24717 VPWR.n3310 VGND 3.13e-19
C24718 VPWR.n3311 VGND 2.56e-19
C24719 VPWR.n3312 VGND 4.55e-19
C24720 VPWR.n3313 VGND 0.00176f
C24721 VPWR.n3314 VGND 9.68e-19
C24722 VPWR.n3315 VGND 9.96e-19
C24723 VPWR.n3316 VGND 3.13e-19
C24724 VPWR.n3317 VGND 4.84e-19
C24725 VPWR.n3318 VGND 6.83e-19
C24726 VPWR.t3405 VGND 0.0592f
C24727 VPWR.n3319 VGND 0.0345f
C24728 VPWR.n3320 VGND 0.00129f
C24729 VPWR.n3321 VGND 4.84e-19
C24730 VPWR.n3322 VGND 5.38e-19
C24731 VPWR.n3323 VGND 4.27e-19
C24732 VPWR.n3324 VGND 5.38e-19
C24733 VPWR.n3325 VGND 4.27e-19
C24734 VPWR.n3326 VGND 0.0033f
C24735 VPWR.n3327 VGND 9.54e-19
C24736 VPWR.n3328 VGND 0.00219f
C24737 VPWR.n3329 VGND 0.00138f
C24738 VPWR.n3330 VGND 3.07e-19
C24739 VPWR.n3331 VGND 5.48e-19
C24740 VPWR.n3332 VGND 0.00138f
C24741 VPWR.n3333 VGND 8.67e-19
C24742 VPWR.n3334 VGND 4.83e-19
C24743 VPWR.n3335 VGND 4.61e-19
C24744 VPWR.n3336 VGND 2.41e-19
C24745 VPWR.n3337 VGND 4.83e-19
C24746 VPWR.n3338 VGND 4.61e-19
C24747 VPWR.n3339 VGND 4.11e-19
C24748 VPWR.n3340 VGND 4.11e-19
C24749 VPWR.n3341 VGND 7.39e-19
C24750 VPWR.n3342 VGND 5.19e-19
C24751 VPWR.n3343 VGND 7.39e-19
C24752 VPWR.n3344 VGND 4.11e-19
C24753 VPWR.n3345 VGND 4.39e-19
C24754 VPWR.n3346 VGND 3.29e-19
C24755 VPWR.n3347 VGND 5.27e-19
C24756 VPWR.n3348 VGND 2.85e-19
C24757 VPWR.n3349 VGND 2.85e-19
C24758 VPWR.n3350 VGND 4.17e-19
C24759 VPWR.n3351 VGND 5.71e-19
C24760 VPWR.n3352 VGND 4.17e-19
C24761 VPWR.n3353 VGND 3.51e-19
C24762 VPWR.n3354 VGND 4.61e-19
C24763 VPWR.n3355 VGND 4.17e-19
C24764 VPWR.n3356 VGND 4.11e-19
C24765 VPWR.n3357 VGND 0.0562f
C24766 VPWR.n3359 VGND 0.0057f
C24767 VPWR.n3361 VGND 0.0952f
C24768 VPWR.n3362 VGND 0.0963f
C24769 VPWR.n3363 VGND 0.00934f
C24770 VPWR.n3365 VGND 7.02e-19
C24771 VPWR.n3366 VGND 0.00138f
C24772 VPWR.n3367 VGND 5.05e-19
C24773 VPWR.n3368 VGND 5.05e-19
C24774 VPWR.n3369 VGND 2.63e-19
C24775 VPWR.n3370 VGND 0.00121f
C24776 VPWR.t942 VGND 0.0065f
C24777 VPWR.n3371 VGND 0.00754f
C24778 VPWR.t3443 VGND 0.00911f
C24779 VPWR.t351 VGND 0.00391f
C24780 VPWR.n3372 VGND 0.0253f
C24781 VPWR.t350 VGND 0.00391f
C24782 VPWR.n3374 VGND 0.0138f
C24783 VPWR.t3567 VGND 0.00911f
C24784 VPWR.t81 VGND 0.00391f
C24785 VPWR.n3375 VGND 0.0253f
C24786 VPWR.t82 VGND 0.00391f
C24787 VPWR.n3377 VGND 0.0138f
C24788 VPWR.n3378 VGND 0.0109f
C24789 VPWR.t3212 VGND 0.00682f
C24790 VPWR.t3214 VGND 0.00166f
C24791 VPWR.t3216 VGND 0.00166f
C24792 VPWR.n3379 VGND 0.00341f
C24793 VPWR.n3380 VGND 0.0101f
C24794 VPWR.n3381 VGND 0.00345f
C24795 VPWR.n3382 VGND 0.00444f
C24796 VPWR.t3398 VGND 0.00911f
C24797 VPWR.t353 VGND 0.00391f
C24798 VPWR.n3383 VGND 0.0253f
C24799 VPWR.t354 VGND 0.00391f
C24800 VPWR.n3385 VGND 0.0138f
C24801 VPWR.n3386 VGND 0.00765f
C24802 VPWR.n3387 VGND 0.0015f
C24803 VPWR.n3388 VGND 0.00393f
C24804 VPWR.t2074 VGND 0.00136f
C24805 VPWR.t1168 VGND 0.00136f
C24806 VPWR.n3389 VGND 0.00317f
C24807 VPWR.t3210 VGND 0.00225f
C24808 VPWR.t2667 VGND 0.00166f
C24809 VPWR.n3390 VGND 0.00438f
C24810 VPWR.n3391 VGND 0.00635f
C24811 VPWR.n3392 VGND 0.00649f
C24812 VPWR.n3393 VGND 0.00524f
C24813 VPWR.n3394 VGND 0.0031f
C24814 VPWR.n3395 VGND 0.00173f
C24815 VPWR.t419 VGND 0.00387f
C24816 VPWR.n3396 VGND 0.00493f
C24817 VPWR.n3397 VGND 0.00525f
C24818 VPWR.n3398 VGND 0.00393f
C24819 VPWR.n3399 VGND 0.00524f
C24820 VPWR.n3400 VGND 0.00524f
C24821 VPWR.t2677 VGND 0.00102f
C24822 VPWR.t1790 VGND 0.00154f
C24823 VPWR.n3401 VGND 0.00483f
C24824 VPWR.t3418 VGND 0.0179f
C24825 VPWR.n3402 VGND 0.0173f
C24826 VPWR.n3403 VGND 0.00792f
C24827 VPWR.n3404 VGND 0.0127f
C24828 VPWR.n3405 VGND 0.00882f
C24829 VPWR.t420 VGND 0.00387f
C24830 VPWR.n3406 VGND 0.00837f
C24831 VPWR.n3407 VGND 0.00504f
C24832 VPWR.n3408 VGND 0.0031f
C24833 VPWR.n3409 VGND 0.00179f
C24834 VPWR.n3410 VGND 0.00179f
C24835 VPWR.n3411 VGND 0.00127f
C24836 VPWR.t1535 VGND 0.00136f
C24837 VPWR.t1997 VGND 0.00136f
C24838 VPWR.n3412 VGND 0.00328f
C24839 VPWR.t938 VGND 0.00645f
C24840 VPWR.n3413 VGND 0.0138f
C24841 VPWR.n3414 VGND 0.00262f
C24842 VPWR.n3415 VGND 0.00262f
C24843 VPWR.n3416 VGND 0.00199f
C24844 VPWR.t781 VGND 0.00166f
C24845 VPWR.t2885 VGND 0.00166f
C24846 VPWR.n3417 VGND 0.00381f
C24847 VPWR.n3418 VGND 0.00759f
C24848 VPWR.t55 VGND 0.00387f
C24849 VPWR.n3419 VGND 0.00837f
C24850 VPWR.n3420 VGND 0.00476f
C24851 VPWR.n3421 VGND 0.00393f
C24852 VPWR.t3343 VGND 0.0231f
C24853 VPWR.n3422 VGND 0.0068f
C24854 VPWR.n3423 VGND 0.0374f
C24855 VPWR.n3424 VGND 0.0039f
C24856 VPWR.n3425 VGND 0.00138f
C24857 VPWR.n3426 VGND 7.39e-19
C24858 VPWR.n3427 VGND 4.11e-19
C24859 VPWR.n3428 VGND 9e-19
C24860 VPWR.n3429 VGND 4.39e-19
C24861 VPWR.n3430 VGND 3.29e-19
C24862 VPWR.n3431 VGND 5.27e-19
C24863 VPWR.n3432 VGND 2.85e-19
C24864 VPWR.n3433 VGND 2.85e-19
C24865 VPWR.n3434 VGND 4.17e-19
C24866 VPWR.n3435 VGND 3.51e-19
C24867 VPWR.n3436 VGND 4.61e-19
C24868 VPWR.n3437 VGND 4.17e-19
C24869 VPWR.n3438 VGND 4.11e-19
C24870 VPWR.n3439 VGND 8.67e-19
C24871 VPWR.n3440 VGND 6.54e-19
C24872 VPWR.n3441 VGND 5.74e-19
C24873 VPWR.n3442 VGND 4.5e-19
C24874 VPWR.n3443 VGND 4.31e-19
C24875 VPWR.n3444 VGND 6.14e-19
C24876 VPWR.n3445 VGND 0.00138f
C24877 VPWR.n3446 VGND 0.00206f
C24878 VPWR.n3447 VGND 0.00153f
C24879 VPWR.n3448 VGND 4.27e-19
C24880 VPWR.n3449 VGND 1.14e-19
C24881 VPWR.t1925 VGND 0.00587f
C24882 VPWR.n3450 VGND 0.00716f
C24883 VPWR.n3451 VGND 3.74e-19
C24884 VPWR.n3452 VGND 0.0068f
C24885 VPWR.n3453 VGND 4.27e-19
C24886 VPWR.n3454 VGND 6.83e-19
C24887 VPWR.n3455 VGND 3.7e-19
C24888 VPWR.n3456 VGND 9.68e-19
C24889 VPWR.n3457 VGND 9.96e-19
C24890 VPWR.n3458 VGND 5.41e-19
C24891 VPWR.n3459 VGND 7.4e-19
C24892 VPWR.n3460 VGND 0.00127f
C24893 VPWR.n3461 VGND 0.00658f
C24894 VPWR.n3462 VGND 3.13e-19
C24895 VPWR.n3463 VGND 2.56e-19
C24896 VPWR.n3464 VGND 4.55e-19
C24897 VPWR.n3465 VGND 0.00575f
C24898 VPWR.n3466 VGND 2.56e-19
C24899 VPWR.n3467 VGND 5.71e-19
C24900 VPWR.n3468 VGND 4.17e-19
C24901 VPWR.n3469 VGND 4.83e-19
C24902 VPWR.n3470 VGND 4.61e-19
C24903 VPWR.n3471 VGND 5.19e-19
C24904 VPWR.n3472 VGND 7.39e-19
C24905 VPWR.n3473 VGND 4.11e-19
C24906 VPWR.n3474 VGND 6.54e-19
C24907 VPWR.n3475 VGND 8.67e-19
C24908 VPWR.n3476 VGND 4.11e-19
C24909 VPWR.n3477 VGND 4.61e-19
C24910 VPWR.n3478 VGND 3.95e-19
C24911 VPWR.n3479 VGND 5.27e-19
C24912 VPWR.n3480 VGND 3.73e-19
C24913 VPWR.n3481 VGND 2.41e-19
C24914 VPWR.n3482 VGND 4.83e-19
C24915 VPWR.n3483 VGND 8.26e-19
C24916 VPWR.n3484 VGND 1.99e-19
C24917 VPWR.n3485 VGND 4.84e-19
C24918 VPWR.n3486 VGND 6.83e-19
C24919 VPWR.n3487 VGND 0.00516f
C24920 VPWR.n3488 VGND 4.84e-19
C24921 VPWR.n3489 VGND 0.00112f
C24922 VPWR.n3490 VGND 4.27e-19
C24923 VPWR.n3491 VGND 0.00112f
C24924 VPWR.n3492 VGND 4.27e-19
C24925 VPWR.n3493 VGND 0.00643f
C24926 VPWR.n3494 VGND 6.26e-19
C24927 VPWR.t56 VGND 0.00387f
C24928 VPWR.n3495 VGND 0.00777f
C24929 VPWR.t932 VGND 5.02e-19
C24930 VPWR.t3194 VGND 0.00135f
C24931 VPWR.n3496 VGND 0.00622f
C24932 VPWR.n3497 VGND 0.0064f
C24933 VPWR.t2168 VGND 0.00265f
C24934 VPWR.n3498 VGND 0.0015f
C24935 VPWR.t955 VGND 0.00692f
C24936 VPWR.n3499 VGND 0.0109f
C24937 VPWR.n3500 VGND 0.00907f
C24938 VPWR.t3553 VGND 0.0179f
C24939 VPWR.n3501 VGND 0.0168f
C24940 VPWR.n3502 VGND 0.0103f
C24941 VPWR.n3503 VGND 0.0133f
C24942 VPWR.t35 VGND 0.00387f
C24943 VPWR.n3504 VGND 0.00837f
C24944 VPWR.t126 VGND 0.0046f
C24945 VPWR.t928 VGND 0.00453f
C24946 VPWR.n3505 VGND 0.00778f
C24947 VPWR.n3506 VGND 0.00184f
C24948 VPWR.t1753 VGND 0.00102f
C24949 VPWR.t1017 VGND 0.00102f
C24950 VPWR.n3507 VGND 0.00217f
C24951 VPWR.n3508 VGND 0.00688f
C24952 VPWR.t127 VGND 0.0046f
C24953 VPWR.n3509 VGND 0.004f
C24954 VPWR.t3489 VGND 0.00911f
C24955 VPWR.t468 VGND 0.00391f
C24956 VPWR.n3510 VGND 0.0253f
C24957 VPWR.t467 VGND 0.00391f
C24958 VPWR.n3512 VGND 0.0138f
C24959 VPWR.n3513 VGND 0.00441f
C24960 VPWR.t2813 VGND 0.0024f
C24961 VPWR.t1152 VGND 0.00678f
C24962 VPWR.n3514 VGND 0.0129f
C24963 VPWR.t987 VGND 6.73e-19
C24964 VPWR.t1150 VGND 0.00127f
C24965 VPWR.n3515 VGND 0.00207f
C24966 VPWR.n3516 VGND 0.00496f
C24967 VPWR.t2099 VGND 0.00527f
C24968 VPWR.n3517 VGND 0.0065f
C24969 VPWR.n3518 VGND 0.00199f
C24970 VPWR.t989 VGND 6.73e-19
C24971 VPWR.t1931 VGND 9.96e-19
C24972 VPWR.n3519 VGND 0.00176f
C24973 VPWR.n3520 VGND 0.00421f
C24974 VPWR.t80 VGND 0.053f
C24975 VPWR.t3211 VGND 0.0463f
C24976 VPWR.t352 VGND 0.0144f
C24977 VPWR.t3213 VGND 0.0183f
C24978 VPWR.t3215 VGND 0.0191f
C24979 VPWR.t3209 VGND 0.0159f
C24980 VPWR.t2073 VGND 0.0161f
C24981 VPWR.t2666 VGND 0.0148f
C24982 VPWR.t1167 VGND 0.0111f
C24983 VPWR.t1789 VGND 0.0358f
C24984 VPWR.t418 VGND 0.0163f
C24985 VPWR.t2676 VGND 0.0237f
C24986 VPWR.t2888 VGND 0.0144f
C24987 VPWR.t941 VGND 0.0154f
C24988 VPWR.t937 VGND 0.0052f
C24989 VPWR.t1534 VGND 0.0112f
C24990 VPWR.t1996 VGND 0.0211f
C24991 VPWR.t780 VGND 0.026f
C24992 VPWR.t2884 VGND 0.0193f
C24993 VPWR.t2678 VGND 0.0458f
C24994 VPWR.t1924 VGND 0.0322f
C24995 VPWR.t54 VGND 0.0112f
C24996 VPWR.t931 VGND 0.0154f
C24997 VPWR.t933 VGND 0.0153f
C24998 VPWR.t3193 VGND 0.0148f
C24999 VPWR.t2061 VGND 0.0141f
C25000 VPWR.t2167 VGND 0.026f
C25001 VPWR.t954 VGND 0.0311f
C25002 VPWR.n3521 VGND 0.0292f
C25003 VPWR.t2826 VGND 0.018f
C25004 VPWR.t980 VGND 0.0275f
C25005 VPWR.t952 VGND 0.0267f
C25006 VPWR.t33 VGND 0.0141f
C25007 VPWR.t1143 VGND 0.02f
C25008 VPWR.t1754 VGND 0.0205f
C25009 VPWR.t927 VGND 0.0436f
C25010 VPWR.t968 VGND 0.0493f
C25011 VPWR.t3158 VGND 0.0398f
C25012 VPWR.t1751 VGND 0.0376f
C25013 VPWR.t125 VGND 0.0166f
C25014 VPWR.t1144 VGND 0.018f
C25015 VPWR.t2470 VGND 0.0603f
C25016 VPWR.t1752 VGND 0.0589f
C25017 VPWR.t1016 VGND 0.025f
C25018 VPWR.t1151 VGND 0.028f
C25019 VPWR.t466 VGND 0.0257f
C25020 VPWR.t2812 VGND 0.0154f
C25021 VPWR.t1906 VGND 0.00906f
C25022 VPWR.t986 VGND 0.0141f
C25023 VPWR.t1621 VGND 0.0181f
C25024 VPWR.t1149 VGND 0.022f
C25025 VPWR.t2532 VGND 0.0233f
C25026 VPWR.t2098 VGND 0.0144f
C25027 VPWR.t2564 VGND 0.0158f
C25028 VPWR.t1341 VGND 0.0166f
C25029 VPWR.t2783 VGND 0.0154f
C25030 VPWR.t2354 VGND 0.0329f
C25031 VPWR.t2796 VGND 0.0369f
C25032 VPWR.t1974 VGND 0.0311f
C25033 VPWR.t2913 VGND 0.0285f
C25034 VPWR.t2696 VGND 0.0322f
C25035 VPWR.t2505 VGND 0.0223f
C25036 VPWR.t643 VGND 0.0141f
C25037 VPWR.t1387 VGND 0.046f
C25038 VPWR.t2694 VGND 0.0567f
C25039 VPWR.t1292 VGND 0.0571f
C25040 VPWR.t24 VGND 0.0361f
C25041 VPWR.t2011 VGND 0.0351f
C25042 VPWR.t2511 VGND 0.0322f
C25043 VPWR.t1294 VGND 0.0322f
C25044 VPWR.t2741 VGND 0.0285f
C25045 VPWR.t2399 VGND 0.0302f
C25046 VPWR.t3174 VGND 0.026f
C25047 VPWR.t506 VGND 0.0331f
C25048 VPWR.t2519 VGND 0.0242f
C25049 VPWR.t3231 VGND 0.0282f
C25050 VPWR.t2402 VGND 0.018f
C25051 VPWR.t550 VGND 0.0046f
C25052 VPWR.n3522 VGND 0.00407f
C25053 VPWR.n3523 VGND 0.00237f
C25054 VPWR.t1015 VGND 0.00102f
C25055 VPWR.t2401 VGND 0.00102f
C25056 VPWR.n3524 VGND 0.00217f
C25057 VPWR.n3525 VGND 0.00653f
C25058 VPWR.t533 VGND 0.00387f
C25059 VPWR.n3526 VGND 0.00837f
C25060 VPWR.n3527 VGND 5.92e-19
C25061 VPWR.n3528 VGND 5.05e-19
C25062 VPWR.n3529 VGND 0.00138f
C25063 VPWR.n3530 VGND 4.31e-19
C25064 VPWR.n3531 VGND 4.17e-19
C25065 VPWR.n3532 VGND 0.00137f
C25066 VPWR.t967 VGND 6.73e-19
C25067 VPWR.t1138 VGND 0.00127f
C25068 VPWR.n3533 VGND 0.00207f
C25069 VPWR.n3534 VGND 0.00451f
C25070 VPWR.n3535 VGND 0.00199f
C25071 VPWR.n3536 VGND 0.00142f
C25072 VPWR.n3537 VGND 0.0015f
C25073 VPWR.n3538 VGND 0.00393f
C25074 VPWR.t1140 VGND 0.00692f
C25075 VPWR.n3539 VGND 0.0108f
C25076 VPWR.n3540 VGND 0.00495f
C25077 VPWR.n3541 VGND 6.65e-19
C25078 VPWR.n3542 VGND 0.00259f
C25079 VPWR.n3543 VGND 2.85e-19
C25080 VPWR.n3544 VGND 1.21e-19
C25081 VPWR.n3545 VGND 2.28e-19
C25082 VPWR.t2952 VGND 0.00242f
C25083 VPWR.n3546 VGND 0.00478f
C25084 VPWR.n3547 VGND 6.26e-19
C25085 VPWR.n3548 VGND 5.12e-19
C25086 VPWR.n3549 VGND 3.13e-19
C25087 VPWR.n3550 VGND 0.00122f
C25088 VPWR.n3551 VGND 0.00108f
C25089 VPWR.n3552 VGND 5.12e-19
C25090 VPWR.n3553 VGND 5.98e-19
C25091 VPWR.t3224 VGND 0.00238f
C25092 VPWR.n3554 VGND 0.0045f
C25093 VPWR.n3555 VGND 3.13e-19
C25094 VPWR.n3556 VGND 5.41e-19
C25095 VPWR.n3557 VGND 9.68e-19
C25096 VPWR.n3558 VGND 9.96e-19
C25097 VPWR.n3559 VGND 5.41e-19
C25098 VPWR.n3560 VGND 6.55e-19
C25099 VPWR.n3561 VGND 6.26e-19
C25100 VPWR.n3562 VGND 5.8e-19
C25101 VPWR.n3563 VGND 3.12e-19
C25102 VPWR.n3564 VGND 7.31e-19
C25103 VPWR.n3565 VGND 5.41e-19
C25104 VPWR.n3566 VGND 5.12e-19
C25105 VPWR.n3567 VGND 4.27e-19
C25106 VPWR.n3568 VGND 9.96e-19
C25107 VPWR.n3569 VGND 0.00131f
C25108 VPWR.n3570 VGND 5.69e-19
C25109 VPWR.n3571 VGND 0.00116f
C25110 VPWR.n3572 VGND 6.8e-19
C25111 VPWR.n3573 VGND 0.00218f
C25112 VPWR.t2566 VGND 0.00102f
C25113 VPWR.t1029 VGND 0.00102f
C25114 VPWR.n3574 VGND 0.00221f
C25115 VPWR.n3575 VGND 0.00627f
C25116 VPWR.n3576 VGND 0.00503f
C25117 VPWR.n3577 VGND 0.0031f
C25118 VPWR.n3578 VGND 0.00137f
C25119 VPWR.t532 VGND 0.00387f
C25120 VPWR.t2404 VGND 0.00453f
C25121 VPWR.t3464 VGND 0.0231f
C25122 VPWR.t993 VGND 6.73e-19
C25123 VPWR.t2281 VGND 9.96e-19
C25124 VPWR.n3579 VGND 0.00176f
C25125 VPWR.n3580 VGND 0.0102f
C25126 VPWR.n3581 VGND 0.0101f
C25127 VPWR.n3582 VGND 0.0366f
C25128 VPWR.n3583 VGND 0.0111f
C25129 VPWR.n3584 VGND 0.00374f
C25130 VPWR.n3585 VGND 0.00525f
C25131 VPWR.n3586 VGND 0.00393f
C25132 VPWR.n3587 VGND 0.00524f
C25133 VPWR.n3588 VGND 0.00524f
C25134 VPWR.n3589 VGND 0.0105f
C25135 VPWR.n3590 VGND 0.00524f
C25136 VPWR.n3591 VGND 0.0133f
C25137 VPWR.n3592 VGND 0.00524f
C25138 VPWR.n3593 VGND 0.0031f
C25139 VPWR.n3594 VGND 0.00515f
C25140 VPWR.t549 VGND 0.0046f
C25141 VPWR.n3595 VGND 0.00407f
C25142 VPWR.n3596 VGND 0.00256f
C25143 VPWR.n3597 VGND 0.00393f
C25144 VPWR.t2744 VGND 0.00234f
C25145 VPWR.n3598 VGND 0.00628f
C25146 VPWR.n3599 VGND 0.00377f
C25147 VPWR.n3600 VGND 0.00524f
C25148 VPWR.n3601 VGND 0.00592f
C25149 VPWR.n3602 VGND 0.00524f
C25150 VPWR.n3603 VGND 0.00506f
C25151 VPWR.n3604 VGND 0.00524f
C25152 VPWR.t3470 VGND 0.0592f
C25153 VPWR.n3605 VGND 0.0356f
C25154 VPWR.t2360 VGND 0.00102f
C25155 VPWR.t1011 VGND 0.00102f
C25156 VPWR.n3606 VGND 0.00217f
C25157 VPWR.n3607 VGND 0.0071f
C25158 VPWR.n3608 VGND 0.00161f
C25159 VPWR.n3609 VGND 0.00524f
C25160 VPWR.n3610 VGND 0.0031f
C25161 VPWR.n3611 VGND 0.00179f
C25162 VPWR.n3612 VGND 0.00653f
C25163 VPWR.n3613 VGND 0.0071f
C25164 VPWR.n3614 VGND 0.00337f
C25165 VPWR.n3615 VGND 0.00475f
C25166 VPWR.n3616 VGND 0.0066f
C25167 VPWR.n3617 VGND 0.00524f
C25168 VPWR.n3618 VGND 0.00592f
C25169 VPWR.n3619 VGND 0.00524f
C25170 VPWR.t1446 VGND 0.00234f
C25171 VPWR.n3620 VGND 0.00628f
C25172 VPWR.n3621 VGND 0.00377f
C25173 VPWR.n3622 VGND 0.00524f
C25174 VPWR.n3623 VGND 0.0031f
C25175 VPWR.t507 VGND 0.00387f
C25176 VPWR.n3624 VGND 0.00493f
C25177 VPWR.t3175 VGND 0.00453f
C25178 VPWR.t3232 VGND 9.96e-19
C25179 VPWR.t2520 VGND 6.73e-19
C25180 VPWR.n3625 VGND 0.00176f
C25181 VPWR.t3456 VGND 0.0179f
C25182 VPWR.n3626 VGND 0.0141f
C25183 VPWR.n3627 VGND 0.00672f
C25184 VPWR.n3628 VGND 0.0101f
C25185 VPWR.n3629 VGND 0.0115f
C25186 VPWR.n3630 VGND 0.0111f
C25187 VPWR.t508 VGND 0.00387f
C25188 VPWR.n3631 VGND 0.00374f
C25189 VPWR.t25 VGND 0.0046f
C25190 VPWR.n3632 VGND 0.00407f
C25191 VPWR.t1293 VGND 0.00676f
C25192 VPWR.n3633 VGND 0.0119f
C25193 VPWR.t644 VGND 0.00462f
C25194 VPWR.n3634 VGND 0.00542f
C25195 VPWR.n3635 VGND 0.0103f
C25196 VPWR.n3636 VGND 0.00279f
C25197 VPWR.n3637 VGND 0.00384f
C25198 VPWR.t26 VGND 0.00462f
C25199 VPWR.n3638 VGND 0.0103f
C25200 VPWR.n3639 VGND 0.0056f
C25201 VPWR.n3640 VGND 0.00333f
C25202 VPWR.n3641 VGND 0.00393f
C25203 VPWR.n3642 VGND 0.0066f
C25204 VPWR.n3643 VGND 0.00642f
C25205 VPWR.n3644 VGND 0.00393f
C25206 VPWR.n3645 VGND 0.00348f
C25207 VPWR.n3646 VGND 0.00524f
C25208 VPWR.t2012 VGND 0.00239f
C25209 VPWR.n3647 VGND 0.00658f
C25210 VPWR.n3648 VGND 0.00456f
C25211 VPWR.n3649 VGND 0.00524f
C25212 VPWR.t3550 VGND 0.0592f
C25213 VPWR.n3650 VGND 0.0356f
C25214 VPWR.n3651 VGND 0.00359f
C25215 VPWR.n3652 VGND 0.00524f
C25216 VPWR.t1295 VGND 0.00127f
C25217 VPWR.t2512 VGND 6.73e-19
C25218 VPWR.n3653 VGND 0.00203f
C25219 VPWR.n3654 VGND 0.00594f
C25220 VPWR.n3655 VGND 0.00222f
C25221 VPWR.n3656 VGND 0.00524f
C25222 VPWR.n3657 VGND 0.00614f
C25223 VPWR.n3658 VGND 0.00524f
C25224 VPWR.n3659 VGND 0.00639f
C25225 VPWR.n3660 VGND 0.00524f
C25226 VPWR.n3661 VGND 0.00393f
C25227 VPWR.n3662 VGND 0.00256f
C25228 VPWR.n3663 VGND 0.00515f
C25229 VPWR.n3664 VGND 0.0031f
C25230 VPWR.n3665 VGND 0.00524f
C25231 VPWR.n3666 VGND 0.00524f
C25232 VPWR.n3667 VGND 0.00393f
C25233 VPWR.n3668 VGND 0.00525f
C25234 VPWR.n3669 VGND 0.00143f
C25235 VPWR.n3670 VGND 0.00199f
C25236 VPWR.n3671 VGND 0.00282f
C25237 VPWR.n3672 VGND 0.0102f
C25238 VPWR.n3673 VGND 0.0204f
C25239 VPWR.t2742 VGND 0.0126f
C25240 VPWR.t1445 VGND 0.0579f
C25241 VPWR.t2400 VGND 0.0589f
C25242 VPWR.t1014 VGND 0.0193f
C25243 VPWR.t548 VGND 0.0154f
C25244 VPWR.t1010 VGND 0.025f
C25245 VPWR.t2359 VGND 0.0589f
C25246 VPWR.t2743 VGND 0.0603f
C25247 VPWR.t1499 VGND 0.0228f
C25248 VPWR.t2358 VGND 0.0327f
C25249 VPWR.t2280 VGND 0.0322f
C25250 VPWR.t531 VGND 0.0163f
C25251 VPWR.t992 VGND 0.0406f
C25252 VPWR.t2403 VGND 0.0436f
C25253 VPWR.t2361 VGND 0.0109f
C25254 VPWR.t1028 VGND 0.0144f
C25255 VPWR.t1498 VGND 0.0141f
C25256 VPWR.t2565 VGND 0.0141f
C25257 VPWR.t1137 VGND 0.0277f
C25258 VPWR.t966 VGND 0.0322f
C25259 VPWR.t2951 VGND 0.0171f
C25260 VPWR.t3223 VGND 0.0185f
C25261 VPWR.t2531 VGND 0.0321f
C25262 VPWR.t2567 VGND 0.0176f
C25263 VPWR.t1139 VGND 0.022f
C25264 VPWR.t1930 VGND 0.0178f
C25265 VPWR.t988 VGND 0.0164f
C25266 VPWR.n3674 VGND 0.0272f
C25267 VPWR.n3675 VGND 0.00941f
C25268 VPWR.n3676 VGND 0.00155f
C25269 VPWR.n3677 VGND 0.00393f
C25270 VPWR.t1342 VGND 0.00208f
C25271 VPWR.t2355 VGND 0.0016f
C25272 VPWR.n3678 VGND 0.00411f
C25273 VPWR.t2784 VGND 0.00453f
C25274 VPWR.n3679 VGND 0.00552f
C25275 VPWR.n3680 VGND 0.0045f
C25276 VPWR.n3681 VGND 0.00103f
C25277 VPWR.n3682 VGND 0.00524f
C25278 VPWR.n3683 VGND 0.0015f
C25279 VPWR.n3684 VGND 0.00524f
C25280 VPWR.n3685 VGND 0.00524f
C25281 VPWR.n3686 VGND 0.00111f
C25282 VPWR.n3687 VGND 0.00524f
C25283 VPWR.n3688 VGND 0.00475f
C25284 VPWR.n3689 VGND 0.00179f
C25285 VPWR.n3690 VGND 0.00105f
C25286 VPWR.n3691 VGND 0.00856f
C25287 VPWR.n3692 VGND 0.00237f
C25288 VPWR.n3693 VGND 0.0031f
C25289 VPWR.n3694 VGND 0.00337f
C25290 VPWR.n3695 VGND 0.00524f
C25291 VPWR.n3696 VGND 0.0066f
C25292 VPWR.n3697 VGND 0.00524f
C25293 VPWR.n3698 VGND 0.00592f
C25294 VPWR.n3699 VGND 0.00524f
C25295 VPWR.t2471 VGND 0.00234f
C25296 VPWR.n3700 VGND 0.00628f
C25297 VPWR.n3701 VGND 0.00398f
C25298 VPWR.n3702 VGND 0.00524f
C25299 VPWR.n3703 VGND 0.0066f
C25300 VPWR.n3704 VGND 0.00524f
C25301 VPWR.n3705 VGND 0.0066f
C25302 VPWR.n3706 VGND 0.00524f
C25303 VPWR.t3576 VGND 0.0592f
C25304 VPWR.n3707 VGND 0.0356f
C25305 VPWR.n3708 VGND 0.00484f
C25306 VPWR.n3709 VGND 0.00524f
C25307 VPWR.n3710 VGND 0.00352f
C25308 VPWR.n3711 VGND 0.00524f
C25309 VPWR.t969 VGND 6.73e-19
C25310 VPWR.t3159 VGND 9.96e-19
C25311 VPWR.n3712 VGND 0.00176f
C25312 VPWR.n3713 VGND 0.00658f
C25313 VPWR.n3714 VGND 0.00484f
C25314 VPWR.n3715 VGND 0.00524f
C25315 VPWR.n3716 VGND 0.00553f
C25316 VPWR.n3717 VGND 0.00524f
C25317 VPWR.n3718 VGND 0.00393f
C25318 VPWR.n3719 VGND 0.00256f
C25319 VPWR.n3720 VGND 0.00515f
C25320 VPWR.n3721 VGND 0.0031f
C25321 VPWR.n3722 VGND 0.00524f
C25322 VPWR.n3723 VGND 0.00524f
C25323 VPWR.t34 VGND 0.00387f
C25324 VPWR.t981 VGND 6.73e-19
C25325 VPWR.t953 VGND 0.00127f
C25326 VPWR.n3724 VGND 0.00203f
C25327 VPWR.n3725 VGND 0.00563f
C25328 VPWR.n3726 VGND 0.00247f
C25329 VPWR.n3727 VGND 0.00525f
C25330 VPWR.n3728 VGND 0.00393f
C25331 VPWR.t2827 VGND 0.00239f
C25332 VPWR.n3729 VGND 0.00421f
C25333 VPWR.n3730 VGND 0.00137f
C25334 VPWR.n3731 VGND 0.00199f
C25335 VPWR.n3732 VGND 0.00199f
C25336 VPWR.n3733 VGND 0.00333f
C25337 VPWR.n3734 VGND 0.00393f
C25338 VPWR.n3735 VGND 0.00179f
C25339 VPWR.n3736 VGND 0.00104f
C25340 VPWR.n3737 VGND 0.00608f
C25341 VPWR.n3738 VGND 0.00118f
C25342 VPWR.n3739 VGND 0.00393f
C25343 VPWR.t934 VGND 0.00136f
C25344 VPWR.t2062 VGND 0.00136f
C25345 VPWR.n3740 VGND 0.00317f
C25346 VPWR.n3741 VGND 0.00693f
C25347 VPWR.n3742 VGND 0.00475f
C25348 VPWR.n3743 VGND 0.00179f
C25349 VPWR.n3744 VGND 0.00122f
C25350 VPWR.n3745 VGND 0.00525f
C25351 VPWR.n3746 VGND 0.00174f
C25352 VPWR.n3747 VGND 9.42e-19
C25353 VPWR.n3748 VGND 0.00131f
C25354 VPWR.n3749 VGND 5.98e-19
C25355 VPWR.n3750 VGND 2.85e-19
C25356 VPWR.n3751 VGND 4.55e-19
C25357 VPWR.n3752 VGND 1.76e-19
C25358 VPWR.n3753 VGND 3.07e-19
C25359 VPWR.n3754 VGND 4.31e-19
C25360 VPWR.n3755 VGND 3.21e-19
C25361 VPWR.n3756 VGND 0.0247f
C25362 VPWR.n3757 VGND 0.37f
C25363 VPWR.n3758 VGND 0.364f
C25364 VPWR.n3759 VGND 0.366f
C25365 VPWR.n3760 VGND 5.19e-19
C25366 VPWR.n3761 VGND 7.39e-19
C25367 VPWR.n3762 VGND 4.11e-19
C25368 VPWR.n3763 VGND 4.83e-19
C25369 VPWR.n3764 VGND 2.85e-19
C25370 VPWR.n3765 VGND 3.95e-19
C25371 VPWR.n3766 VGND 5.71e-19
C25372 VPWR.n3767 VGND 3.29e-19
C25373 VPWR.n3768 VGND 3.95e-19
C25374 VPWR.n3769 VGND 4.17e-19
C25375 VPWR.n3770 VGND 2.85e-19
C25376 VPWR.n3771 VGND 2.85e-19
C25377 VPWR.n3772 VGND 8.67e-19
C25378 VPWR.n3773 VGND 4.11e-19
C25379 VPWR.n3774 VGND 0.00571f
C25380 VPWR.n3775 VGND 5.74e-19
C25381 VPWR.n3776 VGND 6.54e-19
C25382 VPWR.n3777 VGND 8.67e-19
C25383 VPWR.n3778 VGND 7.39e-19
C25384 VPWR.n3779 VGND 4.11e-19
C25385 VPWR.n3780 VGND 3.95e-19
C25386 VPWR.n3781 VGND 3.95e-19
C25387 VPWR.n3782 VGND 4.61e-19
C25388 VPWR.n3783 VGND 2.41e-19
C25389 VPWR.n3784 VGND 3.95e-19
C25390 VPWR.n3785 VGND 5.05e-19
C25391 VPWR.n3786 VGND 4.17e-19
C25392 VPWR.n3787 VGND 6.14e-19
C25393 VPWR.n3788 VGND 4.39e-19
C25394 VPWR.n3789 VGND 1.76e-19
C25395 VPWR.n3790 VGND 3.07e-19
C25396 VPWR.n3791 VGND 4.11e-19
C25397 VPWR.n3793 VGND 0.00934f
C25398 VPWR.n3794 VGND 0.0963f
C25399 VPWR.n3795 VGND 0.0952f
C25400 VPWR.n3796 VGND 4.61e-19
C25401 VPWR.n3797 VGND 2.41e-19
C25402 VPWR.n3798 VGND 3.95e-19
C25403 VPWR.n3799 VGND 6.14e-19
C25404 VPWR.n3800 VGND 4.39e-19
C25405 VPWR.n3801 VGND 1.76e-19
C25406 VPWR.n3802 VGND 3.07e-19
C25407 VPWR.n3803 VGND 4.11e-19
C25408 VPWR.n3804 VGND 4.11e-19
C25409 VPWR.n3805 VGND 7.39e-19
C25410 VPWR.n3806 VGND 5.19e-19
C25411 VPWR.n3807 VGND 7.39e-19
C25412 VPWR.n3808 VGND 4.11e-19
C25413 VPWR.n3809 VGND 4.17e-19
C25414 VPWR.n3810 VGND 5.05e-19
C25415 VPWR.n3811 VGND 4.83e-19
C25416 VPWR.n3812 VGND 2.85e-19
C25417 VPWR.n3813 VGND 3.95e-19
C25418 VPWR.n3814 VGND 5.71e-19
C25419 VPWR.n3815 VGND 3.29e-19
C25420 VPWR.n3816 VGND 3.95e-19
C25421 VPWR.n3817 VGND 4.17e-19
C25422 VPWR.n3818 VGND 2.85e-19
C25423 VPWR.n3819 VGND 2.85e-19
C25424 VPWR.n3820 VGND 6.54e-19
C25425 VPWR.n3821 VGND 8.67e-19
C25426 VPWR.n3822 VGND 4.11e-19
C25427 VPWR.n3824 VGND 0.0057f
C25428 VPWR.n3825 VGND 0.00138f
C25429 VPWR.n3826 VGND 5.48e-19
C25430 VPWR.n3827 VGND 4.17e-19
C25431 VPWR.n3828 VGND 0.00138f
C25432 VPWR.n3829 VGND 0.0022f
C25433 VPWR.t3586 VGND 0.0592f
C25434 VPWR.n3830 VGND 0.0352f
C25435 VPWR.n3831 VGND 0.00344f
C25436 VPWR.n3832 VGND 6.78e-19
C25437 VPWR.n3833 VGND 5.69e-19
C25438 VPWR.n3834 VGND 0.00131f
C25439 VPWR.n3835 VGND 9.96e-19
C25440 VPWR.n3836 VGND 4.27e-19
C25441 VPWR.n3837 VGND 5.12e-19
C25442 VPWR.n3838 VGND 5.41e-19
C25443 VPWR.n3839 VGND 0.00176f
C25444 VPWR.n3840 VGND 5.41e-19
C25445 VPWR.n3841 VGND 4.66e-19
C25446 VPWR.n3842 VGND 3.7e-19
C25447 VPWR.n3843 VGND 4.31e-19
C25448 VPWR.n3844 VGND 3.42e-19
C25449 VPWR.n3845 VGND 0.00172f
C25450 VPWR.n3846 VGND 3.7e-19
C25451 VPWR.n3847 VGND 6.26e-19
C25452 VPWR.n3848 VGND 6.55e-19
C25453 VPWR.n3849 VGND 5.41e-19
C25454 VPWR.n3850 VGND 9.96e-19
C25455 VPWR.n3851 VGND 9.68e-19
C25456 VPWR.n3852 VGND 5.41e-19
C25457 VPWR.t2078 VGND 0.00135f
C25458 VPWR.t1180 VGND 5.02e-19
C25459 VPWR.n3853 VGND 0.00622f
C25460 VPWR.n3854 VGND 0.00834f
C25461 VPWR.n3855 VGND 0.00456f
C25462 VPWR.n3856 VGND 3.13e-19
C25463 VPWR.n3857 VGND 5.98e-19
C25464 VPWR.n3858 VGND 5.12e-19
C25465 VPWR.n3859 VGND 0.00108f
C25466 VPWR.n3860 VGND 0.00122f
C25467 VPWR.n3861 VGND 3.13e-19
C25468 VPWR.n3862 VGND 5.12e-19
C25469 VPWR.n3863 VGND 0.0033f
C25470 VPWR.n3864 VGND 6.26e-19
C25471 VPWR.n3865 VGND 6.1e-19
C25472 VPWR.n3866 VGND 2.28e-19
C25473 VPWR.n3867 VGND 2.85e-19
C25474 VPWR.n3868 VGND 0.00128f
C25475 VPWR.n3869 VGND 0.00309f
C25476 VPWR.n3870 VGND 0.00371f
C25477 VPWR.n3871 VGND 0.00227f
C25478 VPWR.n3872 VGND 0.00262f
C25479 VPWR.n3873 VGND 0.00285f
C25480 VPWR.n3874 VGND 0.00179f
C25481 VPWR.n3875 VGND 0.00199f
C25482 VPWR.n3876 VGND 0.018f
C25483 VPWR.n3877 VGND 0.0382f
C25484 VPWR.t1641 VGND 0.0156f
C25485 VPWR.t786 VGND 0.0433f
C25486 VPWR.t1179 VGND 0.0571f
C25487 VPWR.t2077 VGND 0.0322f
C25488 VPWR.t2163 VGND 0.0311f
C25489 VPWR.t665 VGND 0.0151f
C25490 VPWR.t89 VGND 0.0775f
C25491 VPWR.t2391 VGND 0.0349f
C25492 VPWR.t2389 VGND 0.0255f
C25493 VPWR.t3182 VGND 0.0154f
C25494 VPWR.t3207 VGND 0.0151f
C25495 VPWR.t3203 VGND 0.0438f
C25496 VPWR.t252 VGND 0.0576f
C25497 VPWR.t489 VGND 0.0618f
C25498 VPWR.t95 VGND 0.0126f
C25499 VPWR.t273 VGND 0.0463f
C25500 VPWR.t2957 VGND 0.0257f
C25501 VPWR.t3304 VGND 0.0354f
C25502 VPWR.t732 VGND 0.0415f
C25503 VPWR.t585 VGND 0.067f
C25504 VPWR.t3087 VGND 0.0264f
C25505 VPWR.t1958 VGND 0.0141f
C25506 VPWR.t3089 VGND 0.0141f
C25507 VPWR.t1954 VGND 0.00571f
C25508 VPWR.t1743 VGND 0.0154f
C25509 VPWR.t406 VGND 0.0878f
C25510 VPWR.t480 VGND 0.0975f
C25511 VPWR.n3878 VGND 0.0295f
C25512 VPWR.t145 VGND 0.0126f
C25513 VPWR.t104 VGND 0.0421f
C25514 VPWR.t1890 VGND 0.028f
C25515 VPWR.t1888 VGND 0.0109f
C25516 VPWR.t2039 VGND 0.00554f
C25517 VPWR.t778 VGND 0.0154f
C25518 VPWR.t776 VGND 0.0309f
C25519 VPWR.t625 VGND 0.0878f
C25520 VPWR.t554 VGND 0.0975f
C25521 VPWR.t364 VGND 0.0569f
C25522 VPWR.t685 VGND 0.0665f
C25523 VPWR.n3879 VGND 0.054f
C25524 VPWR.t2765 VGND 0.0272f
C25525 VPWR.t1872 VGND 0.0305f
C25526 VPWR.t1870 VGND 0.0289f
C25527 VPWR.t1868 VGND 0.0289f
C25528 VPWR.t1866 VGND 0.0317f
C25529 VPWR.t427 VGND 0.0222f
C25530 VPWR.t727 VGND 0.0926f
C25531 VPWR.t128 VGND 0.0463f
C25532 VPWR.t181 VGND 0.0111f
C25533 VPWR.t1113 VGND 0.0166f
C25534 VPWR.t1805 VGND 0.0305f
C25535 VPWR.t1803 VGND 0.0289f
C25536 VPWR.t1801 VGND 0.0289f
C25537 VPWR.t1807 VGND 0.0366f
C25538 VPWR.t297 VGND 0.0492f
C25539 VPWR.n3880 VGND 0.0499f
C25540 VPWR.n3881 VGND 0.0131f
C25541 VPWR.n3882 VGND 0.00199f
C25542 VPWR.n3883 VGND 0.00442f
C25543 VPWR.n3884 VGND 0.00179f
C25544 VPWR.n3885 VGND 0.00249f
C25545 VPWR.n3886 VGND 0.00578f
C25546 VPWR.t1808 VGND 0.00682f
C25547 VPWR.n3887 VGND 0.00948f
C25548 VPWR.n3888 VGND 0.00265f
C25549 VPWR.n3889 VGND 0.00393f
C25550 VPWR.n3890 VGND 0.00621f
C25551 VPWR.n3891 VGND 0.00524f
C25552 VPWR.t1802 VGND 0.00166f
C25553 VPWR.t1804 VGND 0.00166f
C25554 VPWR.n3892 VGND 0.00341f
C25555 VPWR.n3893 VGND 0.00445f
C25556 VPWR.n3894 VGND 0.00337f
C25557 VPWR.n3895 VGND 0.00524f
C25558 VPWR.t3380 VGND 0.0592f
C25559 VPWR.n3896 VGND 0.0355f
C25560 VPWR.n3897 VGND 0.00463f
C25561 VPWR.n3898 VGND 0.00524f
C25562 VPWR.t1806 VGND 0.00225f
C25563 VPWR.t1114 VGND 0.00166f
C25564 VPWR.n3899 VGND 0.00438f
C25565 VPWR.n3900 VGND 0.00872f
C25566 VPWR.n3901 VGND 0.00352f
C25567 VPWR.n3902 VGND 0.00524f
C25568 VPWR.n3903 VGND 0.0153f
C25569 VPWR.n3904 VGND 0.00556f
C25570 VPWR.n3905 VGND 0.0031f
C25571 VPWR.n3906 VGND 0.00442f
C25572 VPWR.n3907 VGND 0.00279f
C25573 VPWR.n3908 VGND 0.00529f
C25574 VPWR.n3909 VGND 0.00793f
C25575 VPWR.t728 VGND 0.00387f
C25576 VPWR.n3910 VGND 0.0169f
C25577 VPWR.n3911 VGND 0.00679f
C25578 VPWR.t428 VGND 0.0046f
C25579 VPWR.n3912 VGND 0.00569f
C25580 VPWR.n3913 VGND 0.00907f
C25581 VPWR.n3914 VGND 0.00475f
C25582 VPWR.t3351 VGND 0.0156f
C25583 VPWR.n3915 VGND 0.00623f
C25584 VPWR.n3916 VGND 0.0237f
C25585 VPWR.n3917 VGND 0.00507f
C25586 VPWR.n3918 VGND 0.018f
C25587 VPWR.n3919 VGND 0.0136f
C25588 VPWR.n3920 VGND 0.00524f
C25589 VPWR.n3921 VGND 0.0185f
C25590 VPWR.n3922 VGND 0.00504f
C25591 VPWR.n3923 VGND 3.29e-19
C25592 VPWR.n3924 VGND 5.71e-19
C25593 VPWR.n3925 VGND 5.92e-19
C25594 VPWR.n3926 VGND 5.05e-19
C25595 VPWR.n3927 VGND 0.00139f
C25596 VPWR.n3928 VGND 8.67e-19
C25597 VPWR.n3929 VGND 6.54e-19
C25598 VPWR.n3930 VGND 9.06e-19
C25599 VPWR.n3931 VGND 5.48e-19
C25600 VPWR.n3932 VGND 4.17e-19
C25601 VPWR.n3933 VGND 0.00137f
C25602 VPWR.n3934 VGND 0.00218f
C25603 VPWR.t3478 VGND 0.0592f
C25604 VPWR.n3935 VGND 0.00131f
C25605 VPWR.n3936 VGND 0.00131f
C25606 VPWR.n3937 VGND 0.00432f
C25607 VPWR.n3938 VGND 0.0406f
C25608 VPWR.n3939 VGND 0.0142f
C25609 VPWR.n3940 VGND 6.99e-19
C25610 VPWR.n3941 VGND 5.98e-19
C25611 VPWR.n3942 VGND 0.00131f
C25612 VPWR.n3943 VGND 9.96e-19
C25613 VPWR.n3944 VGND 4.27e-19
C25614 VPWR.n3945 VGND 5.12e-19
C25615 VPWR.n3946 VGND 5.41e-19
C25616 VPWR.n3947 VGND 5.12e-19
C25617 VPWR.n3948 VGND 3.7e-19
C25618 VPWR.n3949 VGND 3.7e-19
C25619 VPWR.n3950 VGND 3.7e-19
C25620 VPWR.n3951 VGND 6.26e-19
C25621 VPWR.n3952 VGND 6.55e-19
C25622 VPWR.n3953 VGND 5.41e-19
C25623 VPWR.n3954 VGND 9.96e-19
C25624 VPWR.n3955 VGND 9.68e-19
C25625 VPWR.n3956 VGND 5.12e-19
C25626 VPWR.n3957 VGND 0.00834f
C25627 VPWR.t729 VGND 0.00387f
C25628 VPWR.n3958 VGND 0.00944f
C25629 VPWR.n3959 VGND 0.00772f
C25630 VPWR.n3960 VGND 3.13e-19
C25631 VPWR.n3961 VGND 4.84e-19
C25632 VPWR.n3962 VGND 6.83e-19
C25633 VPWR.n3963 VGND 2.28e-19
C25634 VPWR.n3964 VGND 3.95e-19
C25635 VPWR.n3965 VGND 4.83e-19
C25636 VPWR.n3966 VGND 2.41e-19
C25637 VPWR.n3967 VGND 3.73e-19
C25638 VPWR.n3968 VGND 3.07e-19
C25639 VPWR.n3969 VGND 6.54e-19
C25640 VPWR.n3970 VGND 8.67e-19
C25641 VPWR.n3971 VGND 4.11e-19
C25642 VPWR.n3973 VGND 0.0057f
C25643 VPWR.n3974 VGND 0.00138f
C25644 VPWR.n3975 VGND 5.48e-19
C25645 VPWR.n3976 VGND 1.76e-19
C25646 VPWR.n3977 VGND 8.11e-19
C25647 VPWR.n3978 VGND 3.95e-19
C25648 VPWR.n3979 VGND 1.77e-19
C25649 VPWR.n3980 VGND 3.13e-19
C25650 VPWR.n3981 VGND 5.12e-19
C25651 VPWR.n3982 VGND 0.00302f
C25652 VPWR.n3983 VGND 5.98e-19
C25653 VPWR.n3984 VGND 6.1e-19
C25654 VPWR.n3985 VGND 2.28e-19
C25655 VPWR.n3986 VGND 3.14e-19
C25656 VPWR.t1867 VGND 0.00682f
C25657 VPWR.n3987 VGND 0.00948f
C25658 VPWR.n3988 VGND 0.00256f
C25659 VPWR.n3989 VGND 0.00621f
C25660 VPWR.n3990 VGND 0.00492f
C25661 VPWR.t1869 VGND 0.00166f
C25662 VPWR.t1871 VGND 0.00166f
C25663 VPWR.n3991 VGND 0.00341f
C25664 VPWR.n3992 VGND 0.00599f
C25665 VPWR.n3993 VGND 0.00337f
C25666 VPWR.n3994 VGND 0.00524f
C25667 VPWR.n3995 VGND 0.00632f
C25668 VPWR.n3996 VGND 0.00524f
C25669 VPWR.t1873 VGND 0.00225f
C25670 VPWR.t2766 VGND 0.00166f
C25671 VPWR.n3997 VGND 0.00438f
C25672 VPWR.n3998 VGND 0.00872f
C25673 VPWR.n3999 VGND 0.0033f
C25674 VPWR.n4000 VGND 0.00524f
C25675 VPWR.t429 VGND 0.0046f
C25676 VPWR.n4001 VGND 0.00407f
C25677 VPWR.n4002 VGND 0.00237f
C25678 VPWR.n4003 VGND 0.0031f
C25679 VPWR.n4004 VGND 0.00199f
C25680 VPWR.n4005 VGND 0.00313f
C25681 VPWR.n4006 VGND 0.00634f
C25682 VPWR.n4007 VGND 0.00671f
C25683 VPWR.t686 VGND 0.00387f
C25684 VPWR.n4008 VGND 0.0161f
C25685 VPWR.n4009 VGND 0.00961f
C25686 VPWR.t365 VGND 0.00387f
C25687 VPWR.t3335 VGND 0.0264f
C25688 VPWR.n4010 VGND 0.0288f
C25689 VPWR.t3447 VGND 0.0282f
C25690 VPWR.n4011 VGND 0.0256f
C25691 VPWR.n4012 VGND 0.019f
C25692 VPWR.n4013 VGND 0.0548f
C25693 VPWR.n4014 VGND 0.0128f
C25694 VPWR.n4015 VGND 0.0216f
C25695 VPWR.n4016 VGND 0.00819f
C25696 VPWR.n4017 VGND 0.00488f
C25697 VPWR.n4018 VGND 0.00393f
C25698 VPWR.n4019 VGND 0.00524f
C25699 VPWR.n4020 VGND 0.00524f
C25700 VPWR.n4021 VGND 0.00524f
C25701 VPWR.n4022 VGND 0.0248f
C25702 VPWR.n4023 VGND 0.00524f
C25703 VPWR.t687 VGND 0.00387f
C25704 VPWR.n4024 VGND 0.0143f
C25705 VPWR.n4025 VGND 0.0156f
C25706 VPWR.n4026 VGND 0.0031f
C25707 VPWR.n4027 VGND 0.00279f
C25708 VPWR.n4028 VGND 0.00634f
C25709 VPWR.t555 VGND 0.00462f
C25710 VPWR.n4029 VGND 0.0102f
C25711 VPWR.t626 VGND 0.0046f
C25712 VPWR.t3546 VGND 0.0592f
C25713 VPWR.n4030 VGND 0.038f
C25714 VPWR.n4031 VGND 0.00833f
C25715 VPWR.n4032 VGND 0.00644f
C25716 VPWR.n4033 VGND 0.00413f
C25717 VPWR.n4034 VGND 0.00393f
C25718 VPWR.n4035 VGND 0.00524f
C25719 VPWR.n4036 VGND 0.00833f
C25720 VPWR.n4037 VGND 0.00524f
C25721 VPWR.n4038 VGND 0.0087f
C25722 VPWR.n4039 VGND 0.00524f
C25723 VPWR.t3535 VGND 0.0592f
C25724 VPWR.n4040 VGND 0.038f
C25725 VPWR.n4041 VGND 0.00833f
C25726 VPWR.n4042 VGND 0.00524f
C25727 VPWR.n4043 VGND 0.0113f
C25728 VPWR.n4044 VGND 0.00524f
C25729 VPWR.n4045 VGND 0.0113f
C25730 VPWR.n4046 VGND 0.00524f
C25731 VPWR.n4047 VGND 0.0113f
C25732 VPWR.n4048 VGND 0.00524f
C25733 VPWR.n4049 VGND 0.011f
C25734 VPWR.n4050 VGND 0.00524f
C25735 VPWR.n4051 VGND 0.0031f
C25736 VPWR.n4052 VGND 0.00527f
C25737 VPWR.n4053 VGND 0.0101f
C25738 VPWR.t627 VGND 0.0046f
C25739 VPWR.n4054 VGND 0.00407f
C25740 VPWR.n4055 VGND 0.00316f
C25741 VPWR.n4056 VGND 0.00475f
C25742 VPWR.n4057 VGND 0.0031f
C25743 VPWR.n4058 VGND 0.00262f
C25744 VPWR.t779 VGND -2.18e-20
C25745 VPWR.t2040 VGND 0.00137f
C25746 VPWR.n4059 VGND 0.00629f
C25747 VPWR.n4060 VGND 0.0139f
C25748 VPWR.n4061 VGND 0.00155f
C25749 VPWR.n4062 VGND 0.00262f
C25750 VPWR.n4063 VGND 0.00262f
C25751 VPWR.n4064 VGND 9.68e-19
C25752 VPWR.n4065 VGND 0.00609f
C25753 VPWR.n4066 VGND 0.00393f
C25754 VPWR.t3367 VGND 0.0179f
C25755 VPWR.t146 VGND 0.00395f
C25756 VPWR.n4067 VGND 0.0261f
C25757 VPWR.n4068 VGND 0.0196f
C25758 VPWR.n4069 VGND 0.00111f
C25759 VPWR.n4070 VGND 0.0031f
C25760 VPWR.n4071 VGND 0.00199f
C25761 VPWR.n4072 VGND 0.00179f
C25762 VPWR.n4073 VGND 0.00341f
C25763 VPWR.t481 VGND 0.00463f
C25764 VPWR.n4074 VGND 0.00571f
C25765 VPWR.t407 VGND 0.0046f
C25766 VPWR.n4075 VGND 0.00644f
C25767 VPWR.n4076 VGND 0.00413f
C25768 VPWR.n4077 VGND 0.00393f
C25769 VPWR.n4078 VGND 0.011f
C25770 VPWR.n4079 VGND 0.00524f
C25771 VPWR.n4080 VGND 0.0087f
C25772 VPWR.n4081 VGND 0.00524f
C25773 VPWR.t3521 VGND 0.0592f
C25774 VPWR.n4082 VGND 0.038f
C25775 VPWR.t3461 VGND 0.0592f
C25776 VPWR.n4083 VGND 0.0376f
C25777 VPWR.n4084 VGND 0.00567f
C25778 VPWR.n4085 VGND 0.00452f
C25779 VPWR.t482 VGND 0.0046f
C25780 VPWR.n4086 VGND 0.00644f
C25781 VPWR.t408 VGND 0.0046f
C25782 VPWR.t1955 VGND 0.00645f
C25783 VPWR.t1744 VGND 0.00137f
C25784 VPWR.t3090 VGND -2.18e-20
C25785 VPWR.n4087 VGND 0.00629f
C25786 VPWR.n4088 VGND 0.0138f
C25787 VPWR.t1959 VGND 0.00631f
C25788 VPWR.n4089 VGND 0.00646f
C25789 VPWR.t3088 VGND 0.00643f
C25790 VPWR.n4090 VGND 0.00199f
C25791 VPWR.n4091 VGND 0.0145f
C25792 VPWR.n4092 VGND 0.00524f
C25793 VPWR.t3579 VGND 0.0291f
C25794 VPWR.t733 VGND 0.00387f
C25795 VPWR.n4093 VGND 0.0649f
C25796 VPWR.n4094 VGND 0.0176f
C25797 VPWR.t3305 VGND 0.00136f
C25798 VPWR.t2958 VGND 0.00136f
C25799 VPWR.n4095 VGND 0.00317f
C25800 VPWR.t734 VGND 0.00387f
C25801 VPWR.t3415 VGND 0.00911f
C25802 VPWR.t275 VGND 0.00391f
C25803 VPWR.n4096 VGND 0.0253f
C25804 VPWR.t274 VGND 0.00391f
C25805 VPWR.n4098 VGND 0.0138f
C25806 VPWR.n4099 VGND 0.0031f
C25807 VPWR.n4100 VGND 0.00444f
C25808 VPWR.t3340 VGND 0.00911f
C25809 VPWR.t701 VGND 0.00391f
C25810 VPWR.n4101 VGND 0.0253f
C25811 VPWR.t702 VGND 0.00391f
C25812 VPWR.n4103 VGND 0.0138f
C25813 VPWR.n4104 VGND 0.0112f
C25814 VPWR.n4105 VGND 0.00487f
C25815 VPWR.n4106 VGND 0.00837f
C25816 VPWR.n4107 VGND 0.0188f
C25817 VPWR.n4108 VGND 0.0116f
C25818 VPWR.n4109 VGND 0.00393f
C25819 VPWR.n4110 VGND 0.00804f
C25820 VPWR.n4111 VGND 0.0192f
C25821 VPWR.n4112 VGND 0.0145f
C25822 VPWR.t3554 VGND 0.0223f
C25823 VPWR.n4113 VGND 0.0202f
C25824 VPWR.t587 VGND 0.00387f
C25825 VPWR.n4114 VGND 0.0274f
C25826 VPWR.t586 VGND 0.00387f
C25827 VPWR.n4115 VGND 0.00782f
C25828 VPWR.n4116 VGND 0.0157f
C25829 VPWR.n4117 VGND 0.00374f
C25830 VPWR.n4118 VGND 0.00362f
C25831 VPWR.n4119 VGND 0.00758f
C25832 VPWR.n4120 VGND 6.05e-20
C25833 VPWR.n4121 VGND 0.00393f
C25834 VPWR.n4122 VGND 0.00141f
C25835 VPWR.n4123 VGND 0.00475f
C25836 VPWR.n4124 VGND 0.00262f
C25837 VPWR.n4125 VGND 0.00262f
C25838 VPWR.n4126 VGND 0.00241f
C25839 VPWR.n4127 VGND 0.0039f
C25840 VPWR.n4128 VGND 0.00512f
C25841 VPWR.n4129 VGND 0.0031f
C25842 VPWR.n4130 VGND 0.011f
C25843 VPWR.n4131 VGND 0.00524f
C25844 VPWR.n4132 VGND 0.0113f
C25845 VPWR.n4133 VGND 0.00524f
C25846 VPWR.n4134 VGND 0.0105f
C25847 VPWR.n4135 VGND 0.00387f
C25848 VPWR.n4136 VGND 0.00203f
C25849 VPWR.n4137 VGND 0.00567f
C25850 VPWR.n4138 VGND 0.00156f
C25851 VPWR.n4139 VGND 4.27e-19
C25852 VPWR.n4140 VGND 8.54e-20
C25853 VPWR.n4141 VGND 0.00105f
C25854 VPWR.n4142 VGND 0.00555f
C25855 VPWR.n4143 VGND 4.27e-19
C25856 VPWR.n4144 VGND 6.83e-19
C25857 VPWR.n4145 VGND 3.7e-19
C25858 VPWR.n4146 VGND 9.68e-19
C25859 VPWR.n4147 VGND 9.96e-19
C25860 VPWR.n4148 VGND 5.41e-19
C25861 VPWR.n4149 VGND 7.4e-19
C25862 VPWR.n4150 VGND 0.00105f
C25863 VPWR.n4151 VGND 0.00549f
C25864 VPWR.n4152 VGND 3.42e-19
C25865 VPWR.n4153 VGND 2.56e-19
C25866 VPWR.n4154 VGND 4.27e-19
C25867 VPWR.n4155 VGND 0.00469f
C25868 VPWR.n4156 VGND 9.68e-19
C25869 VPWR.n4157 VGND 9.96e-19
C25870 VPWR.n4158 VGND 3.13e-19
C25871 VPWR.n4159 VGND 4.84e-19
C25872 VPWR.n4160 VGND 6.83e-19
C25873 VPWR.n4161 VGND 0.00426f
C25874 VPWR.n4162 VGND 4.84e-19
C25875 VPWR.n4163 VGND 9.87e-19
C25876 VPWR.n4164 VGND 4.55e-19
C25877 VPWR.n4165 VGND 9.25e-19
C25878 VPWR.n4166 VGND 4.27e-19
C25879 VPWR.n4167 VGND 0.00265f
C25880 VPWR.n4168 VGND 9.25e-19
C25881 VPWR.n4169 VGND 0.00222f
C25882 VPWR.n4170 VGND 0.00138f
C25883 VPWR.n4171 VGND 5.27e-19
C25884 VPWR.n4172 VGND 3.95e-19
C25885 VPWR.n4173 VGND 5.05e-19
C25886 VPWR.n4174 VGND 5.05e-19
C25887 VPWR.n4175 VGND 3.07e-19
C25888 VPWR.n4176 VGND 5.48e-19
C25889 VPWR.n4178 VGND 0.0057f
C25890 VPWR.n4179 VGND 3.73e-19
C25891 VPWR.n4180 VGND 2.41e-19
C25892 VPWR.n4181 VGND 4.83e-19
C25893 VPWR.n4182 VGND 4.83e-19
C25894 VPWR.n4183 VGND 4.61e-19
C25895 VPWR.n4184 VGND 4.61e-19
C25896 VPWR.n4185 VGND 4.11e-19
C25897 VPWR.n4186 VGND 4.11e-19
C25898 VPWR.n4187 VGND 7.39e-19
C25899 VPWR.n4188 VGND 5.19e-19
C25900 VPWR.n4189 VGND 7.39e-19
C25901 VPWR.n4190 VGND 4.11e-19
C25902 VPWR.n4191 VGND 4.17e-19
C25903 VPWR.n4192 VGND 5.71e-19
C25904 VPWR.n4193 VGND 4.17e-19
C25905 VPWR.n4194 VGND 3.51e-19
C25906 VPWR.n4195 VGND 4.61e-19
C25907 VPWR.n4196 VGND 4.39e-19
C25908 VPWR.n4197 VGND 3.29e-19
C25909 VPWR.n4198 VGND 5.27e-19
C25910 VPWR.n4199 VGND 2.85e-19
C25911 VPWR.n4200 VGND 2.85e-19
C25912 VPWR.n4201 VGND 4.17e-19
C25913 VPWR.n4202 VGND 6.54e-19
C25914 VPWR.n4203 VGND 8.67e-19
C25915 VPWR.n4204 VGND 4.11e-19
C25916 VPWR.n4206 VGND 0.0952f
C25917 VPWR.n4207 VGND 0.0963f
C25918 VPWR.n4208 VGND 0.00934f
C25919 VPWR.n4210 VGND 0.00571f
C25920 VPWR.n4212 VGND 7.39e-19
C25921 VPWR.n4213 VGND 5.19e-19
C25922 VPWR.n4214 VGND 7.39e-19
C25923 VPWR.n4215 VGND 4.11e-19
C25924 VPWR.n4216 VGND 4.11e-19
C25925 VPWR.n4217 VGND 4.61e-19
C25926 VPWR.n4218 VGND 4.83e-19
C25927 VPWR.n4219 VGND 2.41e-19
C25928 VPWR.n4220 VGND 3.73e-19
C25929 VPWR.n4221 VGND 4.84e-19
C25930 VPWR.n4222 VGND 6.55e-19
C25931 VPWR.n4223 VGND 0.00248f
C25932 VPWR.n4224 VGND 2.56e-19
C25933 VPWR.n4225 VGND 5.74e-19
C25934 VPWR.n4226 VGND 4.55e-19
C25935 VPWR.n4227 VGND 5.38e-19
C25936 VPWR.n4228 VGND 4.27e-19
C25937 VPWR.n4229 VGND 0.00154f
C25938 VPWR.n4230 VGND 9.25e-19
C25939 VPWR.n4231 VGND 0.00222f
C25940 VPWR.t2382 VGND 0.00102f
C25941 VPWR.t1772 VGND 0.00102f
C25942 VPWR.n4232 VGND 0.00217f
C25943 VPWR.t3386 VGND 0.0592f
C25944 VPWR.n4233 VGND 0.0353f
C25945 VPWR.n4234 VGND 0.00555f
C25946 VPWR.n4235 VGND 0.00337f
C25947 VPWR.n4236 VGND 0.00452f
C25948 VPWR.n4237 VGND 0.0066f
C25949 VPWR.n4238 VGND 0.00524f
C25950 VPWR.n4239 VGND 0.00592f
C25951 VPWR.n4240 VGND 0.00524f
C25952 VPWR.t340 VGND 0.0046f
C25953 VPWR.t3320 VGND 0.00234f
C25954 VPWR.n4241 VGND 0.00607f
C25955 VPWR.n4242 VGND 0.00145f
C25956 VPWR.n4243 VGND 0.00269f
C25957 VPWR.n4244 VGND 0.00393f
C25958 VPWR.n4245 VGND 0.00199f
C25959 VPWR.n4246 VGND 0.00282f
C25960 VPWR.n4247 VGND 0.0102f
C25961 VPWR.t216 VGND 0.0463f
C25962 VPWR.t213 VGND 0.185f
C25963 VPWR.t620 VGND 0.0878f
C25964 VPWR.t339 VGND 0.0515f
C25965 VPWR.t1771 VGND 0.025f
C25966 VPWR.t2381 VGND 0.0589f
C25967 VPWR.t3319 VGND 0.0525f
C25968 VPWR.t741 VGND 0.018f
C25969 VPWR.n4248 VGND 0.0204f
C25970 VPWR.t2383 VGND 0.0126f
C25971 VPWR.t925 VGND 0.0336f
C25972 VPWR.t2521 VGND 0.0493f
C25973 VPWR.t1449 VGND 0.0497f
C25974 VPWR.t2384 VGND 0.0211f
C25975 VPWR.t151 VGND 0.0144f
C25976 VPWR.t740 VGND 0.024f
C25977 VPWR.t1256 VGND 0.0322f
C25978 VPWR.t2527 VGND 0.0322f
C25979 VPWR.t2970 VGND 0.0502f
C25980 VPWR.t1254 VGND 0.0413f
C25981 VPWR.t69 VGND 0.0772f
C25982 VPWR.t246 VGND 0.0109f
C25983 VPWR.t1761 VGND 0.0144f
C25984 VPWR.t1976 VGND 0.0589f
C25985 VPWR.t1131 VGND 0.0603f
C25986 VPWR.t2914 VGND 0.0321f
C25987 VPWR.t1975 VGND 0.0227f
C25988 VPWR.t2816 VGND 0.0337f
C25989 VPWR.t2517 VGND 0.0164f
C25990 VPWR.n4249 VGND 0.0162f
C25991 VPWR.n4250 VGND 0.00931f
C25992 VPWR.n4251 VGND 0.00274f
C25993 VPWR.n4252 VGND 0.0031f
C25994 VPWR.t2797 VGND 0.00453f
C25995 VPWR.n4253 VGND 0.00778f
C25996 VPWR.n4254 VGND 0.00438f
C25997 VPWR.n4255 VGND 0.00524f
C25998 VPWR.n4256 VGND 0.0066f
C25999 VPWR.n4257 VGND 0.00524f
C26000 VPWR.n4258 VGND 0.0066f
C26001 VPWR.n4259 VGND 0.00524f
C26002 VPWR.n4260 VGND 0.00614f
C26003 VPWR.n4261 VGND 0.00492f
C26004 VPWR.t2506 VGND 6.73e-19
C26005 VPWR.t2697 VGND 0.00127f
C26006 VPWR.n4262 VGND 0.00203f
C26007 VPWR.n4263 VGND 0.00554f
C26008 VPWR.n4264 VGND 4.66e-19
C26009 VPWR.n4265 VGND 0.00256f
C26010 VPWR.n4266 VGND 3.14e-19
C26011 VPWR.n4267 VGND 6.1e-19
C26012 VPWR.n4268 VGND 2.28e-19
C26013 VPWR.n4269 VGND 0.0033f
C26014 VPWR.n4270 VGND 5.98e-19
C26015 VPWR.n4271 VGND 5.12e-19
C26016 VPWR.n4272 VGND 3.13e-19
C26017 VPWR.n4273 VGND 0.00122f
C26018 VPWR.n4274 VGND 0.00108f
C26019 VPWR.n4275 VGND 5.12e-19
C26020 VPWR.n4276 VGND 6.26e-19
C26021 VPWR.t1388 VGND 0.00239f
C26022 VPWR.n4277 VGND 0.00611f
C26023 VPWR.n4278 VGND 0.00513f
C26024 VPWR.n4279 VGND 3.13e-19
C26025 VPWR.n4280 VGND 5.12e-19
C26026 VPWR.n4281 VGND 9.68e-19
C26027 VPWR.n4282 VGND 9.96e-19
C26028 VPWR.n4283 VGND 5.41e-19
C26029 VPWR.n4284 VGND 6.55e-19
C26030 VPWR.n4285 VGND 6.26e-19
C26031 VPWR.n4286 VGND 0.00115f
C26032 VPWR.n4287 VGND 3.7e-19
C26033 VPWR.n4288 VGND 4.66e-19
C26034 VPWR.n4289 VGND 3.7e-19
C26035 VPWR.n4290 VGND 4.66e-19
C26036 VPWR.n4291 VGND 3.7e-19
C26037 VPWR.n4292 VGND 0.00154f
C26038 VPWR.n4293 VGND 5.12e-19
C26039 VPWR.n4294 VGND 5.41e-19
C26040 VPWR.n4295 VGND 5.12e-19
C26041 VPWR.n4296 VGND 4.27e-19
C26042 VPWR.n4297 VGND 9.96e-19
C26043 VPWR.n4298 VGND 0.00131f
C26044 VPWR.n4299 VGND 5.98e-19
C26045 VPWR.n4300 VGND 6.99e-19
C26046 VPWR.n4301 VGND 0.00218f
C26047 VPWR.n4302 VGND 0.00137f
C26048 VPWR.n4303 VGND 5.92e-19
C26049 VPWR.n4304 VGND 5.05e-19
C26050 VPWR.n4305 VGND 4.17e-19
C26051 VPWR.n4306 VGND 4.31e-19
C26052 VPWR.n4307 VGND 7.02e-19
C26053 VPWR.n4308 VGND 3.21e-19
C26054 VPWR.n4309 VGND 0.00138f
C26055 VPWR.n4310 VGND 7.68e-19
C26056 VPWR.n4311 VGND 5.05e-19
C26057 VPWR.n4312 VGND 8.11e-19
C26058 VPWR.n4313 VGND 3.95e-19
C26059 VPWR.n4314 VGND 1.76e-19
C26060 VPWR.n4315 VGND 1.76e-19
C26061 VPWR.n4316 VGND 4.31e-19
C26062 VPWR.n4317 VGND 7.02e-19
C26063 VPWR.n4318 VGND 3.21e-19
C26064 VPWR.n4319 VGND 0.00571f
C26065 VPWR.n4320 VGND 6.54e-19
C26066 VPWR.n4321 VGND 8.67e-19
C26067 VPWR.n4322 VGND 5.19e-19
C26068 VPWR.n4323 VGND 7.39e-19
C26069 VPWR.n4324 VGND 4.11e-19
C26070 VPWR.n4325 VGND 5.71e-19
C26071 VPWR.n4326 VGND 3.29e-19
C26072 VPWR.n4327 VGND 3.95e-19
C26073 VPWR.n4328 VGND 4.17e-19
C26074 VPWR.n4329 VGND 2.85e-19
C26075 VPWR.n4330 VGND 4.83e-19
C26076 VPWR.n4331 VGND 2.85e-19
C26077 VPWR.n4332 VGND 3.95e-19
C26078 VPWR.n4333 VGND 2.85e-19
C26079 VPWR.n4334 VGND 4.11e-19
C26080 VPWR.n4336 VGND 0.00389f
C26081 VPWR.n4337 VGND 0.0976f
C26082 VPWR.n4338 VGND 0.0994f
C26083 VPWR.n4339 VGND 8.67e-19
C26084 VPWR.n4340 VGND 6.54e-19
C26085 VPWR.n4341 VGND 9.06e-19
C26086 VPWR.n4342 VGND 0.00139f
C26087 VPWR.n4343 VGND 3.95e-19
C26088 VPWR.n4344 VGND 3.95e-19
C26089 VPWR.n4345 VGND 7.68e-19
C26090 VPWR.n4346 VGND 5.05e-19
C26091 VPWR.n4347 VGND 8.11e-19
C26092 VPWR.n4348 VGND 3.95e-19
C26093 VPWR.n4349 VGND 1.76e-19
C26094 VPWR.n4350 VGND 1.76e-19
C26095 VPWR.n4351 VGND 5.48e-19
C26096 VPWR.n4353 VGND 0.0057f
C26097 VPWR.n4354 VGND 0.00138f
C26098 VPWR.n4355 VGND 9.06e-19
C26099 VPWR.n4356 VGND 5.48e-19
C26100 VPWR.n4357 VGND 4.17e-19
C26101 VPWR.n4358 VGND 0.00138f
C26102 VPWR.n4359 VGND 0.00218f
C26103 VPWR.t1985 VGND 0.0016f
C26104 VPWR.t2577 VGND 0.0016f
C26105 VPWR.n4360 VGND 0.00365f
C26106 VPWR.n4361 VGND 0.0074f
C26107 VPWR.t3363 VGND 0.0592f
C26108 VPWR.n4362 VGND 0.0353f
C26109 VPWR.n4363 VGND 0.0033f
C26110 VPWR.n4364 VGND 6.99e-19
C26111 VPWR.n4365 VGND 5.98e-19
C26112 VPWR.n4366 VGND 0.00131f
C26113 VPWR.n4367 VGND 9.96e-19
C26114 VPWR.n4368 VGND 4.27e-19
C26115 VPWR.n4369 VGND 5.12e-19
C26116 VPWR.n4370 VGND 5.41e-19
C26117 VPWR.n4371 VGND 0.00154f
C26118 VPWR.n4372 VGND 5.12e-19
C26119 VPWR.n4373 VGND 4.66e-19
C26120 VPWR.n4374 VGND 3.7e-19
C26121 VPWR.n4375 VGND 4.66e-19
C26122 VPWR.n4376 VGND 3.7e-19
C26123 VPWR.t2585 VGND 0.0016f
C26124 VPWR.t2581 VGND 0.0016f
C26125 VPWR.n4377 VGND 0.00367f
C26126 VPWR.n4378 VGND 0.00863f
C26127 VPWR.n4379 VGND 8.25e-19
C26128 VPWR.n4380 VGND 3.7e-19
C26129 VPWR.n4381 VGND 6.26e-19
C26130 VPWR.n4382 VGND 6.55e-19
C26131 VPWR.n4383 VGND 5.41e-19
C26132 VPWR.n4384 VGND 9.96e-19
C26133 VPWR.n4385 VGND 9.68e-19
C26134 VPWR.n4386 VGND 5.12e-19
C26135 VPWR.n4387 VGND 0.00545f
C26136 VPWR.n4388 VGND 3.13e-19
C26137 VPWR.n4389 VGND 6.26e-19
C26138 VPWR.n4390 VGND 5.12e-19
C26139 VPWR.n4391 VGND 0.00108f
C26140 VPWR.n4392 VGND 0.00122f
C26141 VPWR.n4393 VGND 3.13e-19
C26142 VPWR.n4394 VGND 5.12e-19
C26143 VPWR.n4395 VGND 0.0033f
C26144 VPWR.n4396 VGND 5.98e-19
C26145 VPWR.n4397 VGND 5.74e-19
C26146 VPWR.n4398 VGND 2.28e-19
C26147 VPWR.n4399 VGND 3.14e-19
C26148 VPWR.t2575 VGND 0.0016f
C26149 VPWR.t2579 VGND 0.0016f
C26150 VPWR.n4400 VGND 0.00367f
C26151 VPWR.n4401 VGND 0.00619f
C26152 VPWR.n4402 VGND 0.00294f
C26153 VPWR.n4403 VGND 0.00256f
C26154 VPWR.n4404 VGND 0.00599f
C26155 VPWR.n4405 VGND 0.00492f
C26156 VPWR.t2583 VGND 0.00634f
C26157 VPWR.n4406 VGND 0.0121f
C26158 VPWR.t118 VGND 0.00462f
C26159 VPWR.n4407 VGND 0.0148f
C26160 VPWR.n4408 VGND 0.00248f
C26161 VPWR.n4409 VGND 0.00393f
C26162 VPWR.n4410 VGND 0.00444f
C26163 VPWR.n4411 VGND 0.00199f
C26164 VPWR.n4412 VGND 0.00444f
C26165 VPWR.t1454 VGND 0.00102f
C26166 VPWR.t862 VGND 0.00154f
C26167 VPWR.n4413 VGND 0.00486f
C26168 VPWR.n4414 VGND 0.0126f
C26169 VPWR.t1989 VGND 6.73e-19
C26170 VPWR.t3128 VGND 6.73e-19
C26171 VPWR.n4415 VGND 0.00143f
C26172 VPWR.n4416 VGND 0.00449f
C26173 VPWR.n4417 VGND 0.00587f
C26174 VPWR.n4418 VGND 0.00158f
C26175 VPWR.n4419 VGND 0.00393f
C26176 VPWR.n4420 VGND 0.00524f
C26177 VPWR.t1400 VGND 0.00102f
C26178 VPWR.t1204 VGND 0.00154f
C26179 VPWR.n4421 VGND 0.00495f
C26180 VPWR.n4422 VGND 0.00826f
C26181 VPWR.n4423 VGND 0.00524f
C26182 VPWR.t3126 VGND 0.00278f
C26183 VPWR.n4424 VGND 0.00994f
C26184 VPWR.n4425 VGND 0.0031f
C26185 VPWR.n4426 VGND 0.00179f
C26186 VPWR.n4427 VGND 0.00199f
C26187 VPWR.n4428 VGND 0.0012f
C26188 VPWR.n4429 VGND 0.00862f
C26189 VPWR.t289 VGND 0.00387f
C26190 VPWR.t3420 VGND 0.0282f
C26191 VPWR.t1251 VGND 0.0016f
C26192 VPWR.t1245 VGND 0.0016f
C26193 VPWR.n4430 VGND 0.00367f
C26194 VPWR.n4431 VGND 0.00882f
C26195 VPWR.n4432 VGND 0.00908f
C26196 VPWR.n4433 VGND 0.0469f
C26197 VPWR.n4434 VGND 0.01f
C26198 VPWR.n4435 VGND 0.00837f
C26199 VPWR.n4436 VGND 0.00254f
C26200 VPWR.n4437 VGND 0.00393f
C26201 VPWR.n4438 VGND 0.00524f
C26202 VPWR.n4439 VGND 0.00524f
C26203 VPWR.t1249 VGND 0.0016f
C26204 VPWR.t3124 VGND 0.0016f
C26205 VPWR.n4440 VGND 0.00365f
C26206 VPWR.n4441 VGND 0.011f
C26207 VPWR.n4442 VGND 0.0101f
C26208 VPWR.n4443 VGND 0.00524f
C26209 VPWR.n4444 VGND 0.0105f
C26210 VPWR.n4445 VGND 0.00524f
C26211 VPWR.t3120 VGND 0.00631f
C26212 VPWR.n4446 VGND 0.0114f
C26213 VPWR.n4447 VGND 0.00942f
C26214 VPWR.n4448 VGND 0.00524f
C26215 VPWR.n4449 VGND 0.00307f
C26216 VPWR.n4450 VGND 0.0108f
C26217 VPWR.t290 VGND 0.00387f
C26218 VPWR.n4451 VGND 0.00837f
C26219 VPWR.n4452 VGND 0.00488f
C26220 VPWR.n4453 VGND 0.00179f
C26221 VPWR.t2908 VGND 0.00663f
C26222 VPWR.n4454 VGND 0.00874f
C26223 VPWR.n4455 VGND 0.00393f
C26224 VPWR.t2964 VGND 0.00692f
C26225 VPWR.n4456 VGND 0.0106f
C26226 VPWR.n4457 VGND 0.00524f
C26227 VPWR.t2906 VGND -2.18e-20
C26228 VPWR.t3059 VGND 0.00137f
C26229 VPWR.n4458 VGND 0.00618f
C26230 VPWR.n4459 VGND 0.00617f
C26231 VPWR.n4460 VGND 4.23e-19
C26232 VPWR.n4461 VGND 0.00524f
C26233 VPWR.n4462 VGND 0.0031f
C26234 VPWR.n4463 VGND 0.00137f
C26235 VPWR.t380 VGND 0.00387f
C26236 VPWR.t2508 VGND 6.73e-19
C26237 VPWR.t2962 VGND 0.00127f
C26238 VPWR.n4464 VGND 0.00203f
C26239 VPWR.n4465 VGND 0.00906f
C26240 VPWR.n4466 VGND 0.00247f
C26241 VPWR.n4467 VGND 0.00525f
C26242 VPWR.n4468 VGND 0.00393f
C26243 VPWR.t3395 VGND 0.0231f
C26244 VPWR.n4469 VGND 0.0378f
C26245 VPWR.n4470 VGND 0.00524f
C26246 VPWR.n4471 VGND 0.0138f
C26247 VPWR.n4472 VGND 0.00524f
C26248 VPWR.n4473 VGND 0.00524f
C26249 VPWR.n4474 VGND 0.00524f
C26250 VPWR.n4475 VGND 0.0031f
C26251 VPWR.n4476 VGND 0.00199f
C26252 VPWR.n4477 VGND 0.00929f
C26253 VPWR.n4478 VGND 0.00421f
C26254 VPWR.n4479 VGND 0.00142f
C26255 VPWR.n4480 VGND 0.00393f
C26256 VPWR.n4481 VGND 0.00156f
C26257 VPWR.n4482 VGND 0.00333f
C26258 VPWR.n4483 VGND 0.00631f
C26259 VPWR.n4484 VGND 0.00673f
C26260 VPWR.t314 VGND 0.00387f
C26261 VPWR.n4485 VGND 0.00293f
C26262 VPWR.t165 VGND 0.00387f
C26263 VPWR.n4486 VGND 0.0107f
C26264 VPWR.t1756 VGND 0.00136f
C26265 VPWR.t1674 VGND 0.00136f
C26266 VPWR.n4487 VGND 0.00317f
C26267 VPWR.n4488 VGND 0.0121f
C26268 VPWR.t2336 VGND 0.00166f
C26269 VPWR.t2194 VGND 0.00225f
C26270 VPWR.n4489 VGND 0.00438f
C26271 VPWR.t103 VGND 0.0046f
C26272 VPWR.n4490 VGND 0.00385f
C26273 VPWR.n4491 VGND 0.0085f
C26274 VPWR.n4492 VGND 0.00352f
C26275 VPWR.t2196 VGND 0.00166f
C26276 VPWR.t2190 VGND 0.00166f
C26277 VPWR.n4493 VGND 0.00345f
C26278 VPWR.t2031 VGND 0.00136f
C26279 VPWR.t3177 VGND 0.00136f
C26280 VPWR.n4494 VGND 0.00328f
C26281 VPWR.n4495 VGND 0.00727f
C26282 VPWR.t2192 VGND 0.00695f
C26283 VPWR.n4496 VGND 0.00786f
C26284 VPWR.t3568 VGND 0.00911f
C26285 VPWR.t692 VGND 0.00391f
C26286 VPWR.n4497 VGND 0.0253f
C26287 VPWR.t691 VGND 0.00391f
C26288 VPWR.n4499 VGND 0.0138f
C26289 VPWR.t3422 VGND 0.00911f
C26290 VPWR.t449 VGND 0.00391f
C26291 VPWR.n4500 VGND 0.0253f
C26292 VPWR.t450 VGND 0.00391f
C26293 VPWR.n4502 VGND 0.0138f
C26294 VPWR.n4503 VGND 0.011f
C26295 VPWR.n4504 VGND 0.00444f
C26296 VPWR.n4505 VGND 0.0031f
C26297 VPWR.n4506 VGND 0.00524f
C26298 VPWR.n4507 VGND 0.00475f
C26299 VPWR.n4508 VGND 0.00465f
C26300 VPWR.n4509 VGND 0.0024f
C26301 VPWR.n4510 VGND 0.0031f
C26302 VPWR.n4511 VGND 0.00475f
C26303 VPWR.n4512 VGND 0.00179f
C26304 VPWR.n4513 VGND 0.0066f
C26305 VPWR.n4514 VGND 0.0066f
C26306 VPWR.n4515 VGND 0.00393f
C26307 VPWR.n4516 VGND 0.00475f
C26308 VPWR.n4517 VGND 0.00179f
C26309 VPWR.n4518 VGND 0.00629f
C26310 VPWR.n4519 VGND 0.00796f
C26311 VPWR.n4520 VGND 0.0031f
C26312 VPWR.t3562 VGND 0.0592f
C26313 VPWR.n4521 VGND 0.0416f
C26314 VPWR.n4522 VGND 0.013f
C26315 VPWR.n4523 VGND 0.00524f
C26316 VPWR.n4524 VGND 0.0142f
C26317 VPWR.n4525 VGND 0.00524f
C26318 VPWR.n4526 VGND 0.00524f
C26319 VPWR.n4527 VGND 0.00524f
C26320 VPWR.t102 VGND 0.0046f
C26321 VPWR.t164 VGND 0.00387f
C26322 VPWR.n4528 VGND 0.0184f
C26323 VPWR.t3376 VGND 0.0228f
C26324 VPWR.n4529 VGND 0.0164f
C26325 VPWR.n4530 VGND 0.0182f
C26326 VPWR.n4531 VGND 0.00875f
C26327 VPWR.n4532 VGND 0.0115f
C26328 VPWR.n4533 VGND 0.00342f
C26329 VPWR.n4534 VGND 0.00393f
C26330 VPWR.n4535 VGND 0.00179f
C26331 VPWR.n4536 VGND 0.0055f
C26332 VPWR.n4537 VGND 0.00837f
C26333 VPWR.n4538 VGND 0.0123f
C26334 VPWR.n4539 VGND 0.00174f
C26335 VPWR.n4540 VGND 0.00203f
C26336 VPWR.n4541 VGND 0.00156f
C26337 VPWR.n4542 VGND 4.27e-19
C26338 VPWR.n4543 VGND 8.54e-20
C26339 VPWR.t1946 VGND 0.00102f
C26340 VPWR.t1776 VGND 0.00102f
C26341 VPWR.n4544 VGND 0.00217f
C26342 VPWR.n4545 VGND 0.00484f
C26343 VPWR.n4546 VGND 3.74e-19
C26344 VPWR.n4547 VGND 0.00673f
C26345 VPWR.n4548 VGND 4.27e-19
C26346 VPWR.n4549 VGND 6.83e-19
C26347 VPWR.n4550 VGND 3.7e-19
C26348 VPWR.n4551 VGND 9.68e-19
C26349 VPWR.n4552 VGND 9.96e-19
C26350 VPWR.n4553 VGND 5.41e-19
C26351 VPWR.n4554 VGND 7.4e-19
C26352 VPWR.n4555 VGND 3.42e-19
C26353 VPWR.n4556 VGND 2.56e-19
C26354 VPWR.n4557 VGND 4.27e-19
C26355 VPWR.n4558 VGND 9.68e-19
C26356 VPWR.n4559 VGND 9.96e-19
C26357 VPWR.n4560 VGND 3.13e-19
C26358 VPWR.n4561 VGND 4.84e-19
C26359 VPWR.n4562 VGND 6.83e-19
C26360 VPWR.n4563 VGND 7.73e-19
C26361 VPWR.n4564 VGND 2.84e-19
C26362 VPWR.n4565 VGND 0.00123f
C26363 VPWR.n4566 VGND 0.00584f
C26364 VPWR.n4567 VGND 0.00138f
C26365 VPWR.n4568 VGND 3.95e-19
C26366 VPWR.n4569 VGND 5.05e-19
C26367 VPWR.n4570 VGND 5.05e-19
C26368 VPWR.n4571 VGND 3.07e-19
C26369 VPWR.n4572 VGND 9.06e-19
C26370 VPWR.n4573 VGND 5.48e-19
C26371 VPWR.n4574 VGND 0.00138f
C26372 VPWR.n4575 VGND 0.0057f
C26373 VPWR.n4576 VGND 6.54e-19
C26374 VPWR.n4577 VGND 8.67e-19
C26375 VPWR.n4578 VGND 5.19e-19
C26376 VPWR.n4579 VGND 7.39e-19
C26377 VPWR.n4580 VGND 4.11e-19
C26378 VPWR.n4581 VGND 5.27e-19
C26379 VPWR.n4582 VGND 3.73e-19
C26380 VPWR.n4583 VGND 2.41e-19
C26381 VPWR.n4584 VGND 4.83e-19
C26382 VPWR.n4585 VGND 5.71e-19
C26383 VPWR.n4586 VGND 4.17e-19
C26384 VPWR.n4587 VGND 4.83e-19
C26385 VPWR.n4588 VGND 4.61e-19
C26386 VPWR.n4589 VGND 4.61e-19
C26387 VPWR.n4590 VGND 4.11e-19
C26388 VPWR.n4592 VGND 0.1f
C26389 VPWR.n4593 VGND 0.1f
C26390 VPWR.n4594 VGND 0.1f
C26391 VPWR.n4595 VGND 0.1f
C26392 VPWR.n4596 VGND 6.54e-19
C26393 VPWR.n4597 VGND 8.67e-19
C26394 VPWR.n4598 VGND 3.51e-19
C26395 VPWR.n4599 VGND 4.61e-19
C26396 VPWR.n4600 VGND 5.27e-19
C26397 VPWR.n4601 VGND 2.85e-19
C26398 VPWR.n4602 VGND 2.85e-19
C26399 VPWR.n4603 VGND 4.17e-19
C26400 VPWR.n4604 VGND 4.11e-19
C26401 VPWR.n4605 VGND 4.11e-19
C26402 VPWR.n4606 VGND 7.39e-19
C26403 VPWR.n4607 VGND 5.19e-19
C26404 VPWR.n4608 VGND 7.39e-19
C26405 VPWR.n4609 VGND 4.11e-19
C26406 VPWR.n4610 VGND 5.27e-19
C26407 VPWR.n4611 VGND 3.73e-19
C26408 VPWR.n4612 VGND 2.41e-19
C26409 VPWR.n4613 VGND 4.83e-19
C26410 VPWR.n4614 VGND 4.17e-19
C26411 VPWR.n4615 VGND 5.71e-19
C26412 VPWR.n4616 VGND 4.17e-19
C26413 VPWR.n4617 VGND 4.83e-19
C26414 VPWR.n4618 VGND 4.61e-19
C26415 VPWR.n4619 VGND 4.61e-19
C26416 VPWR.n4620 VGND 4.11e-19
C26417 VPWR.n4622 VGND 8.67e-19
C26418 VPWR.n4623 VGND 6.54e-19
C26419 VPWR.n4624 VGND 9.06e-19
C26420 VPWR.n4625 VGND 3.29e-19
C26421 VPWR.n4626 VGND 4.39e-19
C26422 VPWR.n4627 VGND 9e-19
C26423 VPWR.n4628 VGND 0.00138f
C26424 VPWR.n4629 VGND 6.14e-19
C26425 VPWR.n4630 VGND 5.48e-19
C26426 VPWR.n4631 VGND 0.00138f
C26427 VPWR.n4632 VGND 0.0057f
C26428 VPWR.n4633 VGND 0.00139f
C26429 VPWR.n4634 VGND 9.06e-19
C26430 VPWR.t517 VGND 0.00404f
C26431 VPWR.n4635 VGND 0.00212f
C26432 VPWR.t1434 VGND 0.00558f
C26433 VPWR.t593 VGND 0.00387f
C26434 VPWR.n4636 VGND 0.0114f
C26435 VPWR.n4637 VGND 0.00516f
C26436 VPWR.t3541 VGND 0.0176f
C26437 VPWR.n4638 VGND 0.0114f
C26438 VPWR.t592 VGND 0.00387f
C26439 VPWR.n4639 VGND 0.00791f
C26440 VPWR.n4640 VGND 0.0101f
C26441 VPWR.n4641 VGND 0.00717f
C26442 VPWR.n4642 VGND 0.0123f
C26443 VPWR.t3441 VGND 0.00916f
C26444 VPWR.t516 VGND 0.00391f
C26445 VPWR.n4643 VGND 0.0189f
C26446 VPWR.n4644 VGND 0.0106f
C26447 VPWR.n4645 VGND 0.00675f
C26448 VPWR.n4646 VGND 0.00199f
C26449 VPWR.t2320 VGND 0.0235f
C26450 VPWR.t2915 VGND 0.0141f
C26451 VPWR.t2327 VGND 0.0148f
C26452 VPWR.t1031 VGND 0.0141f
C26453 VPWR.t2618 VGND 0.0109f
C26454 VPWR.t2610 VGND 0.0156f
C26455 VPWR.t773 VGND 0.0171f
C26456 VPWR.t2860 VGND 0.0149f
C26457 VPWR.t1610 VGND 0.017f
C26458 VPWR.t1612 VGND 0.0258f
C26459 VPWR.t2612 VGND 0.0193f
C26460 VPWR.t2620 VGND 0.0282f
C26461 VPWR.t1492 VGND 0.0282f
C26462 VPWR.t1490 VGND 0.0468f
C26463 VPWR.t2319 VGND 0.0468f
C26464 VPWR.t2326 VGND 0.0173f
C26465 VPWR.t243 VGND 0.0141f
C26466 VPWR.t3164 VGND 0.025f
C26467 VPWR.t3163 VGND 0.0457f
C26468 VPWR.t3191 VGND 0.0628f
C26469 VPWR.t1972 VGND 0.0331f
C26470 VPWR.t2230 VGND 0.0307f
C26471 VPWR.t2923 VGND 0.0144f
C26472 VPWR.t1385 VGND 0.0141f
C26473 VPWR.t2763 VGND 0.0175f
C26474 VPWR.t2236 VGND 0.0163f
C26475 VPWR.t2616 VGND 0.0121f
C26476 VPWR.t1675 VGND 0.0156f
C26477 VPWR.n4647 VGND 0.00157f
C26478 VPWR.t3014 VGND 0.00586f
C26479 VPWR.n4648 VGND 0.0067f
C26480 VPWR.t1676 VGND 0.00235f
C26481 VPWR.n4649 VGND 2.85e-19
C26482 VPWR.n4650 VGND 0.00186f
C26483 VPWR.n4651 VGND 3.7e-19
C26484 VPWR.n4652 VGND 1.14e-19
C26485 VPWR.n4653 VGND 4.83e-19
C26486 VPWR.n4654 VGND 4.17e-19
C26487 VPWR.n4655 VGND 5.05e-19
C26488 VPWR.n4656 VGND 6.26e-19
C26489 VPWR.n4657 VGND 5.41e-19
C26490 VPWR.n4658 VGND 9.96e-19
C26491 VPWR.n4659 VGND 9.68e-19
C26492 VPWR.n4660 VGND 5.12e-19
C26493 VPWR.t1973 VGND 0.00255f
C26494 VPWR.t2231 VGND 0.00349f
C26495 VPWR.n4661 VGND 0.00938f
C26496 VPWR.n4662 VGND 0.00778f
C26497 VPWR.n4663 VGND 3.13e-19
C26498 VPWR.n4664 VGND 6.26e-19
C26499 VPWR.n4665 VGND 5.12e-19
C26500 VPWR.n4666 VGND 0.00108f
C26501 VPWR.n4667 VGND 0.00122f
C26502 VPWR.n4668 VGND 3.13e-19
C26503 VPWR.n4669 VGND 5.12e-19
C26504 VPWR.n4670 VGND 5.98e-19
C26505 VPWR.t2924 VGND 0.00543f
C26506 VPWR.n4671 VGND 0.00501f
C26507 VPWR.n4672 VGND 8.39e-20
C26508 VPWR.n4673 VGND 4.58e-19
C26509 VPWR.n4674 VGND 0.00256f
C26510 VPWR.n4675 VGND 0.00147f
C26511 VPWR.n4676 VGND 0.00492f
C26512 VPWR.t2617 VGND 0.00102f
C26513 VPWR.t2764 VGND 0.00154f
C26514 VPWR.n4677 VGND 0.00478f
C26515 VPWR.t1386 VGND 9.22e-19
C26516 VPWR.t2237 VGND 9.22e-19
C26517 VPWR.n4678 VGND 0.00201f
C26518 VPWR.n4679 VGND 0.00637f
C26519 VPWR.n4680 VGND 0.00447f
C26520 VPWR.n4681 VGND 9.58e-19
C26521 VPWR.n4682 VGND 0.00524f
C26522 VPWR.n4683 VGND 0.00307f
C26523 VPWR.n4684 VGND 0.00146f
C26524 VPWR.n4685 VGND 0.00579f
C26525 VPWR.n4686 VGND 0.00179f
C26526 VPWR.n4687 VGND 0.00199f
C26527 VPWR.t3016 VGND 0.0065f
C26528 VPWR.n4688 VGND 0.00757f
C26529 VPWR.t3010 VGND 0.00632f
C26530 VPWR.n4689 VGND 0.007f
C26531 VPWR.t1332 VGND 0.00483f
C26532 VPWR.t1398 VGND 0.0048f
C26533 VPWR.n4690 VGND 0.00698f
C26534 VPWR.n4691 VGND 0.00186f
C26535 VPWR.t1396 VGND 6.73e-19
C26536 VPWR.t2121 VGND 0.00343f
C26537 VPWR.n4692 VGND 0.00264f
C26538 VPWR.t2863 VGND 0.00633f
C26539 VPWR.n4693 VGND 0.00967f
C26540 VPWR.n4694 VGND 0.00297f
C26541 VPWR.t1324 VGND 3.74e-19
C26542 VPWR.t2123 VGND 0.00964f
C26543 VPWR.n4695 VGND 0.00544f
C26544 VPWR.n4696 VGND 0.00715f
C26545 VPWR.n4697 VGND 0.00104f
C26546 VPWR.t1060 VGND 0.00614f
C26547 VPWR.n4698 VGND 0.00142f
C26548 VPWR.t1414 VGND 0.00166f
C26549 VPWR.t1438 VGND 0.00166f
C26550 VPWR.n4699 VGND 0.00358f
C26551 VPWR.t2117 VGND 0.00231f
C26552 VPWR.t1134 VGND 0.00231f
C26553 VPWR.n4700 VGND 0.00529f
C26554 VPWR.n4701 VGND 0.0115f
C26555 VPWR.n4702 VGND 9.76e-19
C26556 VPWR.t1410 VGND 0.00166f
C26557 VPWR.t1422 VGND 0.0016f
C26558 VPWR.n4703 VGND 0.00353f
C26559 VPWR.n4704 VGND 0.00636f
C26560 VPWR.n4705 VGND 0.00128f
C26561 VPWR.t2661 VGND 0.00751f
C26562 VPWR.t1416 VGND 0.00166f
C26563 VPWR.t1418 VGND 0.00166f
C26564 VPWR.n4706 VGND 0.00359f
C26565 VPWR.n4707 VGND 0.00596f
C26566 VPWR.n4708 VGND 0.0089f
C26567 VPWR.t1420 VGND 0.00166f
C26568 VPWR.t1424 VGND 0.00166f
C26569 VPWR.n4709 VGND 0.00359f
C26570 VPWR.n4710 VGND 0.00578f
C26571 VPWR.n4711 VGND 0.00606f
C26572 VPWR.t1428 VGND 0.00166f
C26573 VPWR.t1430 VGND 0.00166f
C26574 VPWR.n4712 VGND 0.00355f
C26575 VPWR.n4713 VGND 0.00906f
C26576 VPWR.n4714 VGND 0.00722f
C26577 VPWR.n4715 VGND 0.00199f
C26578 VPWR.n4716 VGND 0.00393f
C26579 VPWR.n4717 VGND 0.00524f
C26580 VPWR.n4718 VGND 0.00524f
C26581 VPWR.n4719 VGND 0.00524f
C26582 VPWR.n4720 VGND 0.00123f
C26583 VPWR.n4721 VGND 0.00524f
C26584 VPWR.n4722 VGND 0.00475f
C26585 VPWR.n4723 VGND 0.00179f
C26586 VPWR.n4724 VGND 0.00112f
C26587 VPWR.t1408 VGND 0.00166f
C26588 VPWR.t1412 VGND 0.00166f
C26589 VPWR.n4725 VGND 0.00359f
C26590 VPWR.n4726 VGND 0.0057f
C26591 VPWR.n4727 VGND 0.00118f
C26592 VPWR.n4728 VGND 0.00393f
C26593 VPWR.t1426 VGND 0.00166f
C26594 VPWR.t1436 VGND 0.00166f
C26595 VPWR.n4729 VGND 0.00353f
C26596 VPWR.n4730 VGND 0.00522f
C26597 VPWR.t1678 VGND 0.00152f
C26598 VPWR.t2615 VGND 6.73e-19
C26599 VPWR.n4731 VGND 0.00226f
C26600 VPWR.n4732 VGND 0.00386f
C26601 VPWR.n4733 VGND 3.32e-19
C26602 VPWR.n4734 VGND 0.00524f
C26603 VPWR.n4735 VGND 0.00524f
C26604 VPWR.t1066 VGND 0.00166f
C26605 VPWR.t1432 VGND 0.00166f
C26606 VPWR.n4736 VGND 0.00388f
C26607 VPWR.t1943 VGND 6.73e-19
C26608 VPWR.t2350 VGND 7.22e-19
C26609 VPWR.n4737 VGND 0.00143f
C26610 VPWR.n4738 VGND 0.00305f
C26611 VPWR.n4739 VGND 0.00646f
C26612 VPWR.n4740 VGND 0.00524f
C26613 VPWR.n4741 VGND 0.0018f
C26614 VPWR.n4742 VGND 0.00524f
C26615 VPWR.t1068 VGND 0.00166f
C26616 VPWR.t1070 VGND 0.00166f
C26617 VPWR.n4743 VGND 0.00379f
C26618 VPWR.n4744 VGND 0.00503f
C26619 VPWR.n4745 VGND 9.88e-19
C26620 VPWR.n4746 VGND 0.00524f
C26621 VPWR.n4747 VGND 0.00475f
C26622 VPWR.n4748 VGND 0.00179f
C26623 VPWR.n4749 VGND 0.00827f
C26624 VPWR.n4750 VGND 6.76e-19
C26625 VPWR.n4751 VGND 0.00342f
C26626 VPWR.n4752 VGND 0.00179f
C26627 VPWR.n4753 VGND 0.00182f
C26628 VPWR.n4754 VGND 0.00179f
C26629 VPWR.n4755 VGND 0.00199f
C26630 VPWR.n4756 VGND 0.00133f
C26631 VPWR.n4757 VGND 0.0129f
C26632 VPWR.n4758 VGND 5.44e-19
C26633 VPWR.n4759 VGND 0.0031f
C26634 VPWR.n4760 VGND 0.00158f
C26635 VPWR.n4761 VGND 0.00524f
C26636 VPWR.n4762 VGND 0.00393f
C26637 VPWR.n4763 VGND 0.00199f
C26638 VPWR.n4764 VGND 0.00904f
C26639 VPWR.n4765 VGND 0.024f
C26640 VPWR.t3013 VGND 0.0233f
C26641 VPWR.t1845 VGND 0.0158f
C26642 VPWR.t3015 VGND 0.0146f
C26643 VPWR.t3009 VGND 0.0176f
C26644 VPWR.t1397 VGND 0.0112f
C26645 VPWR.t1331 VGND 0.0158f
C26646 VPWR.t1742 VGND 0.0154f
C26647 VPWR.t2862 VGND 0.00504f
C26648 VPWR.t1395 VGND 0.0193f
C26649 VPWR.t2120 VGND 0.0228f
C26650 VPWR.t2122 VGND 0.00537f
C26651 VPWR.t1059 VGND 0.0154f
C26652 VPWR.t1067 VGND 0.0277f
C26653 VPWR.t1323 VGND 0.0144f
C26654 VPWR.t1069 VGND 0.0156f
C26655 VPWR.t1065 VGND 0.0146f
C26656 VPWR.t1942 VGND 0.0144f
C26657 VPWR.t1431 VGND 0.0144f
C26658 VPWR.t2349 VGND 0.0143f
C26659 VPWR.t1677 VGND 0.0143f
C26660 VPWR.t1425 VGND 0.0146f
C26661 VPWR.t1435 VGND 0.0196f
C26662 VPWR.t2614 VGND 0.0144f
C26663 VPWR.t1407 VGND 0.0237f
C26664 VPWR.t1411 VGND 0.0171f
C26665 VPWR.t2116 VGND 0.0117f
C26666 VPWR.t1413 VGND 0.0149f
C26667 VPWR.t1437 VGND 0.0176f
C26668 VPWR.t1133 VGND 0.0144f
C26669 VPWR.t1409 VGND 0.0141f
C26670 VPWR.t2868 VGND 0.0143f
C26671 VPWR.t1421 VGND 0.0161f
C26672 VPWR.t1739 VGND 0.0144f
C26673 VPWR.t1415 VGND 0.0193f
C26674 VPWR.t2660 VGND 0.0144f
C26675 VPWR.t1417 VGND 0.0193f
C26676 VPWR.t1419 VGND 0.024f
C26677 VPWR.t1423 VGND 0.0193f
C26678 VPWR.t1427 VGND 0.0289f
C26679 VPWR.t1429 VGND 0.0168f
C26680 VPWR.t591 VGND 0.0144f
C26681 VPWR.t1433 VGND 0.026f
C26682 VPWR.t324 VGND 0.0463f
C26683 VPWR.t2562 VGND 0.0269f
C26684 VPWR.t2560 VGND 0.0289f
C26685 VPWR.t2558 VGND 0.0289f
C26686 VPWR.t2556 VGND 0.0305f
C26687 VPWR.t770 VGND 0.0215f
C26688 VPWR.t385 VGND 0.0158f
C26689 VPWR.t875 VGND 0.0408f
C26690 VPWR.t3162 VGND 0.0171f
C26691 VPWR.t3169 VGND 0.0154f
C26692 VPWR.t3050 VGND 0.0255f
C26693 VPWR.t3111 VGND 0.0358f
C26694 VPWR.t21 VGND 0.0569f
C26695 VPWR.t190 VGND 0.0821f
C26696 VPWR.t515 VGND 0.018f
C26697 VPWR.n4766 VGND 0.0316f
C26698 VPWR.n4767 VGND 0.0143f
C26699 VPWR.n4768 VGND 0.00199f
C26700 VPWR.n4769 VGND 0.00179f
C26701 VPWR.n4770 VGND 0.00252f
C26702 VPWR.t22 VGND 0.00463f
C26703 VPWR.n4771 VGND 0.00569f
C26704 VPWR.t191 VGND 0.00387f
C26705 VPWR.n4772 VGND 0.0107f
C26706 VPWR.n4773 VGND 0.00669f
C26707 VPWR.n4774 VGND 0.00393f
C26708 VPWR.n4775 VGND 0.0135f
C26709 VPWR.n4776 VGND 0.00524f
C26710 VPWR.t3581 VGND 0.0282f
C26711 VPWR.n4777 VGND 0.0512f
C26712 VPWR.t3355 VGND 0.0592f
C26713 VPWR.n4778 VGND 0.00694f
C26714 VPWR.n4779 VGND 0.00161f
C26715 VPWR.n4780 VGND 0.00151f
C26716 VPWR.n4781 VGND 0.00432f
C26717 VPWR.n4782 VGND 0.0409f
C26718 VPWR.n4783 VGND 0.00935f
C26719 VPWR.n4784 VGND 0.00452f
C26720 VPWR.t192 VGND 0.00387f
C26721 VPWR.n4785 VGND 0.0107f
C26722 VPWR.t23 VGND 0.0046f
C26723 VPWR.n4786 VGND 0.00396f
C26724 VPWR.t386 VGND 0.0046f
C26725 VPWR.n4787 VGND 0.00407f
C26726 VPWR.t3480 VGND 0.0592f
C26727 VPWR.t876 VGND 0.00633f
C26728 VPWR.n4788 VGND 0.0103f
C26729 VPWR.n4789 VGND 0.0354f
C26730 VPWR.n4790 VGND 0.00506f
C26731 VPWR.n4791 VGND 0.0066f
C26732 VPWR.t2563 VGND 0.00682f
C26733 VPWR.n4792 VGND 0.00926f
C26734 VPWR.t387 VGND 0.0046f
C26735 VPWR.n4793 VGND 0.00113f
C26736 VPWR.t3375 VGND 0.00911f
C26737 VPWR.t326 VGND 0.00391f
C26738 VPWR.n4794 VGND 0.0253f
C26739 VPWR.t325 VGND 0.00391f
C26740 VPWR.n4796 VGND 0.0138f
C26741 VPWR.n4797 VGND 0.00444f
C26742 VPWR.t3571 VGND 0.00911f
C26743 VPWR.t658 VGND 0.00391f
C26744 VPWR.n4798 VGND 0.0253f
C26745 VPWR.t659 VGND 0.00391f
C26746 VPWR.n4800 VGND 0.0138f
C26747 VPWR.n4801 VGND 0.0112f
C26748 VPWR.n4802 VGND 0.00237f
C26749 VPWR.n4803 VGND 0.0031f
C26750 VPWR.n4804 VGND 0.00624f
C26751 VPWR.n4805 VGND 0.00524f
C26752 VPWR.t2559 VGND 0.00166f
C26753 VPWR.t2561 VGND 0.00166f
C26754 VPWR.n4806 VGND 0.00341f
C26755 VPWR.n4807 VGND 0.00599f
C26756 VPWR.n4808 VGND 0.00334f
C26757 VPWR.n4809 VGND 0.00524f
C26758 VPWR.n4810 VGND 0.00635f
C26759 VPWR.n4811 VGND 0.00524f
C26760 VPWR.t771 VGND 0.00166f
C26761 VPWR.t2557 VGND 0.00225f
C26762 VPWR.n4812 VGND 0.00438f
C26763 VPWR.n4813 VGND 0.00872f
C26764 VPWR.n4814 VGND 0.00352f
C26765 VPWR.n4815 VGND 0.00475f
C26766 VPWR.n4816 VGND 0.00179f
C26767 VPWR.n4817 VGND 0.00199f
C26768 VPWR.n4818 VGND 0.0066f
C26769 VPWR.n4819 VGND 0.00352f
C26770 VPWR.n4820 VGND 0.00393f
C26771 VPWR.n4821 VGND 0.00473f
C26772 VPWR.n4822 VGND 0.00182f
C26773 VPWR.n4823 VGND 0.0066f
C26774 VPWR.n4824 VGND 0.00639f
C26775 VPWR.n4825 VGND 0.00199f
C26776 VPWR.n4826 VGND 0.00262f
C26777 VPWR.n4827 VGND 0.00259f
C26778 VPWR.n4828 VGND 0.00264f
C26779 VPWR.n4829 VGND 0.0031f
C26780 VPWR.t3112 VGND 0.00184f
C26781 VPWR.t3051 VGND 0.00166f
C26782 VPWR.n4830 VGND 0.00358f
C26783 VPWR.n4831 VGND 0.00504f
C26784 VPWR.n4832 VGND 0.00341f
C26785 VPWR.n4833 VGND 0.00524f
C26786 VPWR.n4834 VGND 0.00393f
C26787 VPWR.n4835 VGND 0.00629f
C26788 VPWR.n4836 VGND 0.00796f
C26789 VPWR.n4837 VGND 0.0031f
C26790 VPWR.n4838 VGND 0.00905f
C26791 VPWR.n4839 VGND 0.00171f
C26792 VPWR.n4840 VGND 0.00925f
C26793 VPWR.n4841 VGND 0.0165f
C26794 VPWR.n4842 VGND 0.00387f
C26795 VPWR.n4843 VGND 0.00203f
C26796 VPWR.n4844 VGND 0.00156f
C26797 VPWR.n4845 VGND 4.27e-19
C26798 VPWR.n4846 VGND 8.54e-20
C26799 VPWR.n4847 VGND 4.27e-19
C26800 VPWR.n4848 VGND 6.83e-19
C26801 VPWR.n4849 VGND 3.7e-19
C26802 VPWR.n4850 VGND 9.68e-19
C26803 VPWR.n4851 VGND 9.96e-19
C26804 VPWR.n4852 VGND 5.41e-19
C26805 VPWR.n4853 VGND 7.4e-19
C26806 VPWR.n4854 VGND 0.00171f
C26807 VPWR.n4855 VGND 0.00895f
C26808 VPWR.n4856 VGND 3.42e-19
C26809 VPWR.n4857 VGND 2.56e-19
C26810 VPWR.n4858 VGND 4.27e-19
C26811 VPWR.n4859 VGND 0.00764f
C26812 VPWR.n4860 VGND 9.68e-19
C26813 VPWR.n4861 VGND 9.96e-19
C26814 VPWR.n4862 VGND 3.13e-19
C26815 VPWR.n4863 VGND 4.84e-19
C26816 VPWR.n4864 VGND 6.83e-19
C26817 VPWR.n4865 VGND 4.84e-19
C26818 VPWR.n4866 VGND 4.55e-19
C26819 VPWR.n4867 VGND 4.27e-19
C26820 VPWR.n4868 VGND 9.25e-19
C26821 VPWR.n4869 VGND 0.00222f
C26822 VPWR.n4870 VGND 0.00138f
C26823 VPWR.n4871 VGND 3.95e-19
C26824 VPWR.n4872 VGND 5.05e-19
C26825 VPWR.n4873 VGND 5.05e-19
C26826 VPWR.n4874 VGND 3.07e-19
C26827 VPWR.n4875 VGND 5.48e-19
C26828 VPWR.n4877 VGND 0.0194f
C26829 VPWR.n4878 VGND 0.0976f
C26830 VPWR.n4879 VGND 0.0839f
C26831 VPWR.n4880 VGND 6.54e-19
C26832 VPWR.n4881 VGND 8.67e-19
C26833 VPWR.n4882 VGND 3.51e-19
C26834 VPWR.n4883 VGND 4.61e-19
C26835 VPWR.n4884 VGND 5.27e-19
C26836 VPWR.n4885 VGND 2.85e-19
C26837 VPWR.n4886 VGND 2.85e-19
C26838 VPWR.n4887 VGND 4.17e-19
C26839 VPWR.n4888 VGND 4.11e-19
C26840 VPWR.n4889 VGND 4.11e-19
C26841 VPWR.n4890 VGND 7.39e-19
C26842 VPWR.n4891 VGND 5.19e-19
C26843 VPWR.n4892 VGND 7.39e-19
C26844 VPWR.n4893 VGND 4.11e-19
C26845 VPWR.n4894 VGND 5.27e-19
C26846 VPWR.n4895 VGND 3.73e-19
C26847 VPWR.n4896 VGND 2.41e-19
C26848 VPWR.n4897 VGND 4.83e-19
C26849 VPWR.n4898 VGND 4.17e-19
C26850 VPWR.n4899 VGND 5.71e-19
C26851 VPWR.n4900 VGND 4.17e-19
C26852 VPWR.n4901 VGND 4.83e-19
C26853 VPWR.n4902 VGND 4.61e-19
C26854 VPWR.n4903 VGND 4.61e-19
C26855 VPWR.n4904 VGND 4.11e-19
C26856 VPWR.n4906 VGND 8.67e-19
C26857 VPWR.n4907 VGND 6.54e-19
C26858 VPWR.n4908 VGND 9.06e-19
C26859 VPWR.n4909 VGND 3.29e-19
C26860 VPWR.n4910 VGND 4.39e-19
C26861 VPWR.n4911 VGND 9e-19
C26862 VPWR.t41 VGND 0.00387f
C26863 VPWR.n4912 VGND 0.00837f
C26864 VPWR.t2950 VGND 0.00453f
C26865 VPWR.n4913 VGND 0.00552f
C26866 VPWR.t404 VGND 0.00387f
C26867 VPWR.t3400 VGND 0.0179f
C26868 VPWR.t2226 VGND 0.00102f
C26869 VPWR.t1764 VGND 0.00102f
C26870 VPWR.n4914 VGND 0.00217f
C26871 VPWR.n4915 VGND 0.0102f
C26872 VPWR.n4916 VGND 0.00702f
C26873 VPWR.n4917 VGND 0.0103f
C26874 VPWR.n4918 VGND 0.0173f
C26875 VPWR.n4919 VGND 0.00493f
C26876 VPWR.n4920 VGND 0.00457f
C26877 VPWR.t2433 VGND 0.00238f
C26878 VPWR.t405 VGND 0.00387f
C26879 VPWR.n4921 VGND 0.00822f
C26880 VPWR.t3563 VGND 0.00911f
C26881 VPWR.t124 VGND 0.00391f
C26882 VPWR.n4922 VGND 0.0253f
C26883 VPWR.t123 VGND 0.00391f
C26884 VPWR.n4924 VGND 0.0138f
C26885 VPWR.n4925 VGND 0.00444f
C26886 VPWR.t3494 VGND 0.00911f
C26887 VPWR.t663 VGND 0.00391f
C26888 VPWR.n4926 VGND 0.0253f
C26889 VPWR.t664 VGND 0.00391f
C26890 VPWR.n4928 VGND 0.0138f
C26891 VPWR.n4929 VGND 0.0112f
C26892 VPWR.n4930 VGND 0.00487f
C26893 VPWR.n4931 VGND 0.0031f
C26894 VPWR.n4932 VGND 0.00524f
C26895 VPWR.n4933 VGND 0.00524f
C26896 VPWR.n4934 VGND 0.00393f
C26897 VPWR.n4935 VGND 0.00199f
C26898 VPWR.n4936 VGND 0.00541f
C26899 VPWR.n4937 VGND 0.00179f
C26900 VPWR.n4938 VGND 0.0031f
C26901 VPWR.n4939 VGND 0.00186f
C26902 VPWR.n4940 VGND 0.00524f
C26903 VPWR.n4941 VGND 0.00185f
C26904 VPWR.n4942 VGND 0.00524f
C26905 VPWR.t1494 VGND 0.00524f
C26906 VPWR.n4943 VGND 0.00489f
C26907 VPWR.n4944 VGND 5.04e-19
C26908 VPWR.n4945 VGND 0.00524f
C26909 VPWR.t2514 VGND 6.73e-19
C26910 VPWR.t837 VGND 9.96e-19
C26911 VPWR.n4946 VGND 0.00176f
C26912 VPWR.n4947 VGND 0.00421f
C26913 VPWR.n4948 VGND 0.00136f
C26914 VPWR.n4949 VGND 0.00524f
C26915 VPWR.t2035 VGND 0.0016f
C26916 VPWR.t2803 VGND 0.00208f
C26917 VPWR.n4950 VGND 0.00411f
C26918 VPWR.n4951 VGND 0.00482f
C26919 VPWR.n4952 VGND 0.00103f
C26920 VPWR.n4953 VGND 0.00524f
C26921 VPWR.n4954 VGND 0.00393f
C26922 VPWR.n4955 VGND 0.0011f
C26923 VPWR.n4956 VGND 0.00525f
C26924 VPWR.n4957 VGND 0.0031f
C26925 VPWR.n4958 VGND 0.0133f
C26926 VPWR.n4959 VGND 0.00524f
C26927 VPWR.n4960 VGND 0.0128f
C26928 VPWR.n4961 VGND 0.00524f
C26929 VPWR.t2524 VGND 6.73e-19
C26930 VPWR.t2977 VGND 0.00127f
C26931 VPWR.n4962 VGND 0.00203f
C26932 VPWR.n4963 VGND 0.00951f
C26933 VPWR.n4964 VGND 0.00538f
C26934 VPWR.n4965 VGND 0.00524f
C26935 VPWR.n4966 VGND 0.00387f
C26936 VPWR.n4967 VGND 6.83e-19
C26937 VPWR.n4968 VGND 4.84e-19
C26938 VPWR.n4969 VGND 3.13e-19
C26939 VPWR.n4970 VGND 9.96e-19
C26940 VPWR.n4971 VGND 9.68e-19
C26941 VPWR.n4972 VGND 4.7e-19
C26942 VPWR.n4973 VGND 2.14e-19
C26943 VPWR.n4974 VGND 3.42e-19
C26944 VPWR.n4975 VGND 7.4e-19
C26945 VPWR.n4976 VGND 5.41e-19
C26946 VPWR.n4977 VGND 9.96e-19
C26947 VPWR.n4978 VGND 9.68e-19
C26948 VPWR.n4979 VGND 3.7e-19
C26949 VPWR.n4980 VGND 6.83e-19
C26950 VPWR.n4981 VGND 4.27e-19
C26951 VPWR.n4982 VGND 4.61e-19
C26952 VPWR.n4983 VGND 0.00136f
C26953 VPWR.n4984 VGND 0.00229f
C26954 VPWR.n4985 VGND 0.00138f
C26955 VPWR.n4986 VGND 6.14e-19
C26956 VPWR.n4987 VGND 5.48e-19
C26957 VPWR.n4988 VGND 0.00138f
C26958 VPWR.n4989 VGND 0.0057f
C26959 VPWR.n4991 VGND 9.06e-19
C26960 VPWR.n4992 VGND 5.48e-19
C26961 VPWR.n4993 VGND 3.07e-19
C26962 VPWR.n4994 VGND 1.76e-19
C26963 VPWR.n4995 VGND 2.63e-19
C26964 VPWR.n4996 VGND 9.42e-19
C26965 VPWR.n4997 VGND 8.27e-19
C26966 VPWR.n4998 VGND 6.26e-19
C26967 VPWR.n4999 VGND 3.42e-19
C26968 VPWR.n5000 VGND 4.84e-19
C26969 VPWR.n5001 VGND 9.15e-19
C26970 VPWR.n5002 VGND 2.62e-19
C26971 VPWR.t3538 VGND 0.0289f
C26972 VPWR.t40 VGND 0.00387f
C26973 VPWR.n5003 VGND 0.0604f
C26974 VPWR.n5004 VGND 0.0146f
C26975 VPWR.n5005 VGND 0.0117f
C26976 VPWR.n5006 VGND 0.00992f
C26977 VPWR.n5007 VGND 0.00487f
C26978 VPWR.n5008 VGND 0.0031f
C26979 VPWR.n5009 VGND 0.00475f
C26980 VPWR.n5010 VGND 0.00179f
C26981 VPWR.n5011 VGND 0.00333f
C26982 VPWR.n5012 VGND 0.0138f
C26983 VPWR.n5013 VGND 0.0384f
C26984 VPWR.n5014 VGND 0.00837f
C26985 VPWR.n5015 VGND 0.0132f
C26986 VPWR.t122 VGND 0.0463f
C26987 VPWR.t1763 VGND 0.025f
C26988 VPWR.t2225 VGND 0.0151f
C26989 VPWR.t403 VGND 0.0371f
C26990 VPWR.t2432 VGND 0.0151f
C26991 VPWR.t1951 VGND 0.0109f
C26992 VPWR.t2013 VGND 0.0166f
C26993 VPWR.t2224 VGND 0.0141f
C26994 VPWR.t874 VGND 0.0235f
C26995 VPWR.t836 VGND 0.0312f
C26996 VPWR.t1493 VGND 0.0163f
C26997 VPWR.t2513 VGND 0.0158f
C26998 VPWR.t2802 VGND 0.023f
C26999 VPWR.t2034 VGND 0.0255f
C27000 VPWR.t2949 VGND 0.0206f
C27001 VPWR.t2223 VGND 0.0205f
C27002 VPWR.t1950 VGND 0.0285f
C27003 VPWR.t2976 VGND 0.0322f
C27004 VPWR.t2523 VGND 0.0223f
C27005 VPWR.t39 VGND 0.0141f
C27006 VPWR.t1217 VGND 0.046f
C27007 VPWR.t2978 VGND 0.0567f
C27008 VPWR.t2871 VGND 0.0257f
C27009 VPWR.t2059 VGND 0.02f
C27010 VPWR.t400 VGND 0.0153f
C27011 VPWR.n5016 VGND 0.05f
C27012 VPWR.t1740 VGND 0.0425f
C27013 VPWR.t3038 VGND 0.0329f
C27014 VPWR.t612 VGND 0.0153f
C27015 VPWR.t1497 VGND 0.0144f
C27016 VPWR.t2864 VGND 0.0425f
C27017 VPWR.t1393 VGND 0.0217f
C27018 VPWR.t1043 VGND 0.0203f
C27019 VPWR.t2351 VGND 0.026f
C27020 VPWR.t3298 VGND 0.0248f
C27021 VPWR.t3292 VGND 0.0252f
C27022 VPWR.t1136 VGND 0.0141f
C27023 VPWR.t3288 VGND 0.0121f
C27024 VPWR.t2063 VGND 0.0141f
C27025 VPWR.t3294 VGND 0.0161f
C27026 VPWR.t1041 VGND 0.0141f
C27027 VPWR.t3296 VGND 0.0171f
C27028 VPWR.t3290 VGND 0.0253f
C27029 VPWR.t1457 VGND 0.017f
C27030 VPWR.t1455 VGND 0.0154f
C27031 VPWR.t696 VGND 0.0138f
C27032 VPWR.t2929 VGND 0.027f
C27033 VPWR.t2944 VGND 0.0146f
C27034 VPWR.t2940 VGND 0.0149f
C27035 VPWR.t2228 VGND 0.0141f
C27036 VPWR.t2946 VGND 0.0158f
C27037 VPWR.t3007 VGND 0.0141f
C27038 VPWR.t2942 VGND 0.0294f
C27039 VPWR.t1403 VGND 0.0196f
C27040 VPWR.t1040 VGND 0.0141f
C27041 VPWR.t1193 VGND 0.0141f
C27042 VPWR.t3064 VGND 0.00705f
C27043 VPWR.t1135 VGND 0.0154f
C27044 VPWR.t2866 VGND 0.0111f
C27045 VPWR.t3121 VGND 0.00621f
C27046 VPWR.t3331 VGND 0.0181f
C27047 VPWR.n5017 VGND 0.0179f
C27048 VPWR.n5018 VGND 0.00984f
C27049 VPWR.n5019 VGND 0.00199f
C27050 VPWR.n5020 VGND 0.00262f
C27051 VPWR.n5021 VGND 1.21e-19
C27052 VPWR.n5022 VGND 0.00687f
C27053 VPWR.n5023 VGND 0.00179f
C27054 VPWR.n5024 VGND 0.00307f
C27055 VPWR.n5025 VGND 0.00179f
C27056 VPWR.n5026 VGND 0.00524f
C27057 VPWR.t1729 VGND 0.00633f
C27058 VPWR.n5027 VGND 0.00969f
C27059 VPWR.n5028 VGND 5.85e-19
C27060 VPWR.n5029 VGND 0.00393f
C27061 VPWR.n5030 VGND 0.00285f
C27062 VPWR.n5031 VGND 0.00122f
C27063 VPWR.n5032 VGND 9.28e-19
C27064 VPWR.n5033 VGND 4.27e-19
C27065 VPWR.n5034 VGND 3.14e-19
C27066 VPWR.n5035 VGND 1.71e-19
C27067 VPWR.n5036 VGND 2.28e-19
C27068 VPWR.n5037 VGND 9.28e-19
C27069 VPWR.n5038 VGND 5.98e-19
C27070 VPWR.n5039 VGND 5.12e-19
C27071 VPWR.n5040 VGND 3.13e-19
C27072 VPWR.n5041 VGND 1.77e-19
C27073 VPWR.n5042 VGND 1.76e-19
C27074 VPWR.n5043 VGND 5.48e-19
C27075 VPWR.n5044 VGND 0.00138f
C27076 VPWR.n5045 VGND 0.0057f
C27077 VPWR.n5047 VGND 6.14e-19
C27078 VPWR.n5048 VGND 4.39e-19
C27079 VPWR.n5049 VGND 1.76e-19
C27080 VPWR.n5050 VGND 4.83e-19
C27081 VPWR.n5051 VGND 2.41e-19
C27082 VPWR.n5052 VGND 3.73e-19
C27083 VPWR.n5053 VGND 3.07e-19
C27084 VPWR.n5054 VGND 4.11e-19
C27085 VPWR.n5055 VGND 4.11e-19
C27086 VPWR.n5056 VGND 7.39e-19
C27087 VPWR.n5057 VGND 5.19e-19
C27088 VPWR.n5058 VGND 7.39e-19
C27089 VPWR.n5059 VGND 4.11e-19
C27090 VPWR.n5060 VGND 4.11e-19
C27091 VPWR.n5061 VGND 2.85e-19
C27092 VPWR.n5062 VGND 3.95e-19
C27093 VPWR.n5063 VGND 2.85e-19
C27094 VPWR.n5064 VGND 4.83e-19
C27095 VPWR.n5065 VGND 4.17e-19
C27096 VPWR.n5066 VGND 5.05e-19
C27097 VPWR.n5067 VGND 6.55e-19
C27098 VPWR.n5068 VGND 6.26e-19
C27099 VPWR.n5069 VGND 8.97e-19
C27100 VPWR.n5070 VGND 3.7e-19
C27101 VPWR.n5071 VGND 1.31e-19
C27102 VPWR.n5072 VGND 3.7e-19
C27103 VPWR.n5073 VGND 1.31e-19
C27104 VPWR.n5074 VGND 3.7e-19
C27105 VPWR.n5075 VGND 6.55e-19
C27106 VPWR.n5076 VGND 5.12e-19
C27107 VPWR.n5077 VGND 5.41e-19
C27108 VPWR.n5078 VGND 5.12e-19
C27109 VPWR.n5079 VGND 4.27e-19
C27110 VPWR.n5080 VGND 2.85e-19
C27111 VPWR.n5081 VGND 0.00125f
C27112 VPWR.n5082 VGND 5.98e-19
C27113 VPWR.n5083 VGND 6.99e-19
C27114 VPWR.n5084 VGND 0.00218f
C27115 VPWR.n5085 VGND 0.00453f
C27116 VPWR.n5086 VGND 0.00182f
C27117 VPWR.n5087 VGND 0.00199f
C27118 VPWR.n5088 VGND 0.00186f
C27119 VPWR.n5089 VGND 0.00154f
C27120 VPWR.n5090 VGND 0.00484f
C27121 VPWR.t1116 VGND 0.0048f
C27122 VPWR.t1738 VGND 0.00483f
C27123 VPWR.n5091 VGND 0.00727f
C27124 VPWR.t2052 VGND 0.00483f
C27125 VPWR.t2288 VGND 0.0048f
C27126 VPWR.n5092 VGND 0.00727f
C27127 VPWR.n5093 VGND 0.0276f
C27128 VPWR.n5094 VGND 0.00699f
C27129 VPWR.n5095 VGND 0.00166f
C27130 VPWR.n5096 VGND 0.00698f
C27131 VPWR.n5097 VGND 0.00146f
C27132 VPWR.n5098 VGND 0.00524f
C27133 VPWR.n5099 VGND 0.00393f
C27134 VPWR.t1120 VGND 0.00597f
C27135 VPWR.n5100 VGND 0.0142f
C27136 VPWR.n5101 VGND 0.00158f
C27137 VPWR.n5102 VGND 0.0031f
C27138 VPWR.t1192 VGND 0.00166f
C27139 VPWR.t1122 VGND 0.00166f
C27140 VPWR.n5103 VGND 0.0037f
C27141 VPWR.t3281 VGND -2.18e-20
C27142 VPWR.t1987 VGND 0.00137f
C27143 VPWR.n5104 VGND 0.00618f
C27144 VPWR.n5105 VGND 0.00641f
C27145 VPWR.n5106 VGND 0.00525f
C27146 VPWR.n5107 VGND 9.48e-19
C27147 VPWR.n5108 VGND 0.00524f
C27148 VPWR.n5109 VGND 0.00154f
C27149 VPWR.n5110 VGND 0.00524f
C27150 VPWR.n5111 VGND 0.00393f
C27151 VPWR.n5112 VGND 0.00199f
C27152 VPWR.n5113 VGND 0.00179f
C27153 VPWR.n5114 VGND 0.00442f
C27154 VPWR.n5115 VGND 0.0186f
C27155 VPWR.n5116 VGND 0.00199f
C27156 VPWR.n5117 VGND 0.00182f
C27157 VPWR.t3198 VGND 0.00219f
C27158 VPWR.t2932 VGND 0.00166f
C27159 VPWR.n5118 VGND 0.00445f
C27160 VPWR.n5119 VGND 0.0114f
C27161 VPWR.n5120 VGND 0.00113f
C27162 VPWR.n5121 VGND 0.00333f
C27163 VPWR.n5122 VGND 0.00393f
C27164 VPWR.t3200 VGND 0.00532f
C27165 VPWR.n5123 VGND 0.00667f
C27166 VPWR.n5124 VGND 0.0111f
C27167 VPWR.n5125 VGND 6.73e-19
C27168 VPWR.n5126 VGND 0.00307f
C27169 VPWR.n5127 VGND 0.0126f
C27170 VPWR.n5128 VGND 0.00524f
C27171 VPWR.n5129 VGND 0.00524f
C27172 VPWR.n5130 VGND 0.00524f
C27173 VPWR.t3487 VGND 0.0231f
C27174 VPWR.t647 VGND 0.00387f
C27175 VPWR.n5131 VGND 0.00837f
C27176 VPWR.t767 VGND 0.00593f
C27177 VPWR.t765 VGND 0.0016f
C27178 VPWR.t1712 VGND 0.0016f
C27179 VPWR.n5132 VGND 0.00363f
C27180 VPWR.n5133 VGND 0.00967f
C27181 VPWR.n5134 VGND 0.00762f
C27182 VPWR.n5135 VGND 0.0124f
C27183 VPWR.n5136 VGND 0.012f
C27184 VPWR.n5137 VGND 0.0328f
C27185 VPWR.n5138 VGND 0.00393f
C27186 VPWR.n5139 VGND 0.00179f
C27187 VPWR.n5140 VGND 0.00199f
C27188 VPWR.n5141 VGND 0.0148f
C27189 VPWR.n5142 VGND 0.00103f
C27190 VPWR.n5143 VGND 0.0031f
C27191 VPWR.n5144 VGND 0.00524f
C27192 VPWR.t2323 VGND 0.00102f
C27193 VPWR.t1505 VGND 0.00154f
C27194 VPWR.n5145 VGND 0.00483f
C27195 VPWR.n5146 VGND 0.00645f
C27196 VPWR.n5147 VGND 0.00102f
C27197 VPWR.n5148 VGND 0.00524f
C27198 VPWR.t1531 VGND 0.0016f
C27199 VPWR.t1164 VGND 0.0016f
C27200 VPWR.n5149 VGND 0.00327f
C27201 VPWR.n5150 VGND 0.00351f
C27202 VPWR.n5151 VGND 0.00119f
C27203 VPWR.n5152 VGND 0.00524f
C27204 VPWR.n5153 VGND 0.00393f
C27205 VPWR.n5154 VGND 0.00186f
C27206 VPWR.n5155 VGND 0.00154f
C27207 VPWR.n5156 VGND 0.00307f
C27208 VPWR.n5157 VGND 0.00524f
C27209 VPWR.n5158 VGND 0.00103f
C27210 VPWR.n5159 VGND 0.00502f
C27211 VPWR.n5160 VGND 0.0022f
C27212 VPWR.n5161 VGND 6.78e-19
C27213 VPWR.n5162 VGND 5.69e-19
C27214 VPWR.n5163 VGND 0.00131f
C27215 VPWR.n5164 VGND 9.96e-19
C27216 VPWR.n5165 VGND 4.27e-19
C27217 VPWR.n5166 VGND 5.12e-19
C27218 VPWR.n5167 VGND 5.41e-19
C27219 VPWR.n5168 VGND 7.31e-19
C27220 VPWR.n5169 VGND 3.12e-19
C27221 VPWR.n5170 VGND 5.8e-19
C27222 VPWR.n5171 VGND 6.26e-19
C27223 VPWR.n5172 VGND 6.55e-19
C27224 VPWR.n5173 VGND 5.41e-19
C27225 VPWR.n5174 VGND 9.96e-19
C27226 VPWR.n5175 VGND 5.98e-19
C27227 VPWR.n5176 VGND 5.12e-19
C27228 VPWR.n5177 VGND 3.95e-19
C27229 VPWR.n5178 VGND 5.05e-19
C27230 VPWR.n5179 VGND 4.17e-19
C27231 VPWR.n5180 VGND 6.14e-19
C27232 VPWR.n5181 VGND 4.39e-19
C27233 VPWR.n5182 VGND 1.76e-19
C27234 VPWR.n5183 VGND 3.07e-19
C27235 VPWR.n5184 VGND 4.83e-19
C27236 VPWR.n5185 VGND 2.85e-19
C27237 VPWR.n5186 VGND 3.95e-19
C27238 VPWR.n5187 VGND 3.95e-19
C27239 VPWR.n5188 VGND 4.17e-19
C27240 VPWR.n5189 VGND 2.85e-19
C27241 VPWR.n5190 VGND 2.85e-19
C27242 VPWR.n5191 VGND 4.11e-19
C27243 VPWR.n5192 VGND 4.11e-19
C27244 VPWR.n5193 VGND 7.39e-19
C27245 VPWR.n5194 VGND 5.19e-19
C27246 VPWR.n5195 VGND 7.39e-19
C27247 VPWR.n5196 VGND 4.11e-19
C27248 VPWR.n5197 VGND 4.11e-19
C27249 VPWR.n5199 VGND 0.0839f
C27250 VPWR.n5200 VGND 0.0976f
C27251 VPWR.n5201 VGND 1.01f
C27252 VPWR.n5202 VGND 0.564f
C27253 VPWR.n5203 VGND 0.746f
C27254 VPWR.n5204 VGND 0.0976f
C27255 VPWR.n5205 VGND 0.0194f
C27256 VPWR.n5206 VGND 0.00139f
C27257 VPWR.n5207 VGND 9.06e-19
C27258 VPWR.n5208 VGND 5.92e-19
C27259 VPWR.n5209 VGND 5.05e-19
C27260 VPWR.n5210 VGND 4.17e-19
C27261 VPWR.n5211 VGND 5.48e-19
C27262 VPWR.n5213 VGND 8.67e-19
C27263 VPWR.n5214 VGND 6.54e-19
C27264 VPWR.n5215 VGND 9.06e-19
C27265 VPWR.n5216 VGND 3.95e-19
C27266 VPWR.n5217 VGND 3.95e-19
C27267 VPWR.n5218 VGND 7.68e-19
C27268 VPWR.n5219 VGND 5.05e-19
C27269 VPWR.n5220 VGND 8.11e-19
C27270 VPWR.n5221 VGND 3.95e-19
C27271 VPWR.n5222 VGND 1.77e-19
C27272 VPWR.n5223 VGND 1.76e-19
C27273 VPWR.n5224 VGND 5.48e-19
C27274 VPWR.n5225 VGND 0.00138f
C27275 VPWR.n5226 VGND 0.0057f
C27276 VPWR.n5228 VGND 6.14e-19
C27277 VPWR.n5229 VGND 4.39e-19
C27278 VPWR.n5230 VGND 1.76e-19
C27279 VPWR.n5231 VGND 4.83e-19
C27280 VPWR.n5232 VGND 2.41e-19
C27281 VPWR.n5233 VGND 3.73e-19
C27282 VPWR.n5234 VGND 3.07e-19
C27283 VPWR.n5235 VGND 4.11e-19
C27284 VPWR.n5236 VGND 4.11e-19
C27285 VPWR.n5237 VGND 7.39e-19
C27286 VPWR.n5238 VGND 5.19e-19
C27287 VPWR.n5239 VGND 7.39e-19
C27288 VPWR.n5240 VGND 4.11e-19
C27289 VPWR.n5241 VGND 4.11e-19
C27290 VPWR.n5242 VGND 2.85e-19
C27291 VPWR.n5243 VGND 2.85e-19
C27292 VPWR.n5244 VGND 4.17e-19
C27293 VPWR.n5245 VGND 5.41e-19
C27294 VPWR.n5246 VGND 5.12e-19
C27295 VPWR.n5247 VGND 4.27e-19
C27296 VPWR.n5248 VGND 2.85e-19
C27297 VPWR.n5249 VGND 0.00125f
C27298 VPWR.n5250 VGND 5.98e-19
C27299 VPWR.t3192 VGND 0.00236f
C27300 VPWR.n5251 VGND 0.0065f
C27301 VPWR.n5252 VGND 0.0042f
C27302 VPWR.n5253 VGND 6.99e-19
C27303 VPWR.n5254 VGND 0.00218f
C27304 VPWR.n5255 VGND 0.00535f
C27305 VPWR.n5256 VGND 0.00504f
C27306 VPWR.n5257 VGND 0.0066f
C27307 VPWR.n5258 VGND 0.00524f
C27308 VPWR.n5259 VGND 0.0066f
C27309 VPWR.n5260 VGND 0.00524f
C27310 VPWR.n5261 VGND 0.0066f
C27311 VPWR.n5262 VGND 0.00524f
C27312 VPWR.n5263 VGND 0.0066f
C27313 VPWR.n5264 VGND 0.00524f
C27314 VPWR.t3346 VGND 0.0592f
C27315 VPWR.n5265 VGND 0.0356f
C27316 VPWR.n5266 VGND 0.00484f
C27317 VPWR.n5267 VGND 0.00524f
C27318 VPWR.n5268 VGND 0.00506f
C27319 VPWR.n5269 VGND 0.00524f
C27320 VPWR.n5270 VGND 0.0066f
C27321 VPWR.n5271 VGND 0.00524f
C27322 VPWR.n5272 VGND 0.00639f
C27323 VPWR.n5273 VGND 0.00524f
C27324 VPWR.n5274 VGND 0.00393f
C27325 VPWR.n5275 VGND 0.00255f
C27326 VPWR.n5276 VGND 0.00147f
C27327 VPWR.n5277 VGND 0.00179f
C27328 VPWR.n5278 VGND 0.00199f
C27329 VPWR.n5279 VGND 0.00393f
C27330 VPWR.n5280 VGND 0.00473f
C27331 VPWR.n5281 VGND 0.00182f
C27332 VPWR.n5282 VGND 0.00564f
C27333 VPWR.n5283 VGND 0.00126f
C27334 VPWR.n5284 VGND 0.0031f
C27335 VPWR.n5285 VGND 0.00524f
C27336 VPWR.n5286 VGND 0.00143f
C27337 VPWR.n5287 VGND 0.00393f
C27338 VPWR.n5288 VGND 0.00199f
C27339 VPWR.n5289 VGND 0.00907f
C27340 VPWR.n5290 VGND 0.00168f
C27341 VPWR.n5291 VGND 0.00182f
C27342 VPWR.n5292 VGND 0.00333f
C27343 VPWR.n5293 VGND 0.00393f
C27344 VPWR.n5294 VGND 0.00179f
C27345 VPWR.t2330 VGND 0.00647f
C27346 VPWR.n5295 VGND 0.0142f
C27347 VPWR.n5296 VGND 0.00121f
C27348 VPWR.n5297 VGND 0.00307f
C27349 VPWR.n5298 VGND 0.00524f
C27350 VPWR.n5299 VGND 0.00121f
C27351 VPWR.n5300 VGND 0.00524f
C27352 VPWR.n5301 VGND 0.00524f
C27353 VPWR.n5302 VGND 0.00524f
C27354 VPWR.t2129 VGND 0.00166f
C27355 VPWR.t2131 VGND 0.00166f
C27356 VPWR.n5303 VGND 0.00359f
C27357 VPWR.n5304 VGND 0.00536f
C27358 VPWR.n5305 VGND 9.86e-19
C27359 VPWR.n5306 VGND 0.00524f
C27360 VPWR.t1237 VGND 0.0016f
C27361 VPWR.t2176 VGND 0.00214f
C27362 VPWR.n5307 VGND 0.00419f
C27363 VPWR.n5308 VGND 0.00645f
C27364 VPWR.n5309 VGND 5.29e-19
C27365 VPWR.n5310 VGND 0.00524f
C27366 VPWR.n5311 VGND 0.00393f
C27367 VPWR.n5312 VGND 0.00136f
C27368 VPWR.n5313 VGND 0.00783f
C27369 VPWR.n5314 VGND 4.25e-19
C27370 VPWR.n5315 VGND 0.00393f
C27371 VPWR.n5316 VGND 0.00478f
C27372 VPWR.n5317 VGND 0.00151f
C27373 VPWR.n5318 VGND 9.64e-19
C27374 VPWR.n5319 VGND 0.00177f
C27375 VPWR.n5320 VGND 0.00444f
C27376 VPWR.n5321 VGND 0.00307f
C27377 VPWR.n5322 VGND 0.00502f
C27378 VPWR.n5323 VGND 0.0022f
C27379 VPWR.n5324 VGND 0.00138f
C27380 VPWR.n5325 VGND 4.17e-19
C27381 VPWR.n5326 VGND 5.48e-19
C27382 VPWR.n5327 VGND 0.00138f
C27383 VPWR.n5328 VGND 0.0057f
C27384 VPWR.n5329 VGND 6.54e-19
C27385 VPWR.n5330 VGND 8.67e-19
C27386 VPWR.n5331 VGND 3.95e-19
C27387 VPWR.n5332 VGND 4.61e-19
C27388 VPWR.n5333 VGND 2.41e-19
C27389 VPWR.n5334 VGND 3.95e-19
C27390 VPWR.n5335 VGND 5.05e-19
C27391 VPWR.n5336 VGND 4.17e-19
C27392 VPWR.n5337 VGND 6.14e-19
C27393 VPWR.n5338 VGND 4.39e-19
C27394 VPWR.n5339 VGND 1.76e-19
C27395 VPWR.n5340 VGND 3.07e-19
C27396 VPWR.n5341 VGND 4.83e-19
C27397 VPWR.n5342 VGND 2.85e-19
C27398 VPWR.n5343 VGND 3.95e-19
C27399 VPWR.n5344 VGND 3.95e-19
C27400 VPWR.n5345 VGND 4.17e-19
C27401 VPWR.n5346 VGND 2.85e-19
C27402 VPWR.n5347 VGND 2.85e-19
C27403 VPWR.n5348 VGND 4.11e-19
C27404 VPWR.n5349 VGND 4.11e-19
C27405 VPWR.n5350 VGND 7.39e-19
C27406 VPWR.n5351 VGND 5.19e-19
C27407 VPWR.n5352 VGND 7.39e-19
C27408 VPWR.n5353 VGND 4.11e-19
C27409 VPWR.n5354 VGND 4.11e-19
C27410 VPWR.n5356 VGND 0.1f
C27411 VPWR.n5357 VGND 0.1f
C27412 VPWR.n5358 VGND 0.00139f
C27413 VPWR.n5359 VGND 9.06e-19
C27414 VPWR.n5360 VGND 8.11e-19
C27415 VPWR.n5361 VGND 3.95e-19
C27416 VPWR.n5362 VGND 1.76e-19
C27417 VPWR.n5363 VGND 3.95e-19
C27418 VPWR.n5364 VGND 7.68e-19
C27419 VPWR.n5365 VGND 5.05e-19
C27420 VPWR.n5366 VGND 1.76e-19
C27421 VPWR.n5367 VGND 5.48e-19
C27422 VPWR.n5369 VGND 8.67e-19
C27423 VPWR.n5370 VGND 6.54e-19
C27424 VPWR.n5371 VGND 9.06e-19
C27425 VPWR.n5372 VGND 3.29e-19
C27426 VPWR.n5373 VGND 5.71e-19
C27427 VPWR.n5374 VGND 5.92e-19
C27428 VPWR.n5375 VGND 5.05e-19
C27429 VPWR.n5376 VGND 4.17e-19
C27430 VPWR.n5377 VGND 5.48e-19
C27431 VPWR.n5378 VGND 0.00138f
C27432 VPWR.n5379 VGND 0.0057f
C27433 VPWR.n5381 VGND 4.11e-19
C27434 VPWR.n5382 VGND 4.11e-19
C27435 VPWR.n5383 VGND 7.39e-19
C27436 VPWR.n5384 VGND 5.19e-19
C27437 VPWR.n5385 VGND 7.39e-19
C27438 VPWR.n5386 VGND 4.11e-19
C27439 VPWR.n5387 VGND 4.11e-19
C27440 VPWR.n5388 VGND 2.85e-19
C27441 VPWR.n5389 VGND 2.85e-19
C27442 VPWR.n5390 VGND 3.95e-19
C27443 VPWR.n5391 VGND 4.17e-19
C27444 VPWR.n5392 VGND 3.99e-19
C27445 VPWR.n5393 VGND 5.12e-19
C27446 VPWR.n5394 VGND 4.27e-19
C27447 VPWR.n5395 VGND 2.56e-19
C27448 VPWR.n5396 VGND 0.00128f
C27449 VPWR.n5397 VGND 5.69e-19
C27450 VPWR.n5398 VGND 0.00174f
C27451 VPWR.n5399 VGND 6.78e-19
C27452 VPWR.n5400 VGND 0.0022f
C27453 VPWR.t1523 VGND 5.02e-19
C27454 VPWR.t2178 VGND 0.00135f
C27455 VPWR.n5401 VGND 0.00633f
C27456 VPWR.n5402 VGND 0.00696f
C27457 VPWR.n5403 VGND 0.00102f
C27458 VPWR.n5404 VGND 0.00502f
C27459 VPWR.n5405 VGND 0.0011f
C27460 VPWR.n5406 VGND 0.00524f
C27461 VPWR.t2542 VGND 0.00131f
C27462 VPWR.t2076 VGND 4.27e-19
C27463 VPWR.n5407 VGND 0.00672f
C27464 VPWR.n5408 VGND 0.00391f
C27465 VPWR.n5409 VGND 9.48e-19
C27466 VPWR.n5410 VGND 0.00524f
C27467 VPWR.n5411 VGND 0.00307f
C27468 VPWR.n5412 VGND 7.56e-19
C27469 VPWR.n5413 VGND 0.0141f
C27470 VPWR.n5414 VGND 0.00393f
C27471 VPWR.n5415 VGND 0.00134f
C27472 VPWR.n5416 VGND 0.00524f
C27473 VPWR.t2544 VGND 0.00225f
C27474 VPWR.t1640 VGND 0.00202f
C27475 VPWR.n5417 VGND 0.00473f
C27476 VPWR.n5418 VGND 0.00526f
C27477 VPWR.n5419 VGND 0.0012f
C27478 VPWR.n5420 VGND 0.00524f
C27479 VPWR.t1635 VGND 0.00196f
C27480 VPWR.t2546 VGND 0.00196f
C27481 VPWR.n5421 VGND 0.00402f
C27482 VPWR.n5422 VGND 0.00423f
C27483 VPWR.n5423 VGND 0.00107f
C27484 VPWR.n5424 VGND 0.00524f
C27485 VPWR.n5425 VGND 9.58e-19
C27486 VPWR.n5426 VGND 0.00524f
C27487 VPWR.t1638 VGND 0.00557f
C27488 VPWR.t3047 VGND 0.00496f
C27489 VPWR.n5427 VGND 0.00845f
C27490 VPWR.t3045 VGND 0.00208f
C27491 VPWR.t3006 VGND 0.00202f
C27492 VPWR.n5428 VGND 0.00536f
C27493 VPWR.n5429 VGND 0.0194f
C27494 VPWR.n5430 VGND 0.00524f
C27495 VPWR.n5431 VGND 0.00307f
C27496 VPWR.n5432 VGND 0.00146f
C27497 VPWR.t3041 VGND 0.0016f
C27498 VPWR.t2338 VGND 0.0016f
C27499 VPWR.n5433 VGND 0.00363f
C27500 VPWR.n5434 VGND 0.00343f
C27501 VPWR.n5435 VGND 9.88e-19
C27502 VPWR.n5436 VGND 0.00199f
C27503 VPWR.n5437 VGND 0.00618f
C27504 VPWR.n5438 VGND 0.00333f
C27505 VPWR.n5439 VGND 0.00393f
C27506 VPWR.n5440 VGND 0.0113f
C27507 VPWR.n5441 VGND 0.0138f
C27508 VPWR.t2956 VGND 0.00261f
C27509 VPWR.n5442 VGND 0.0111f
C27510 VPWR.n5443 VGND 0.00979f
C27511 VPWR.n5444 VGND 0.00179f
C27512 VPWR.n5445 VGND 0.00262f
C27513 VPWR.n5446 VGND 0.00525f
C27514 VPWR.t2799 VGND 0.00117f
C27515 VPWR.n5447 VGND 0.00331f
C27516 VPWR.t906 VGND 4.34e-19
C27517 VPWR.n5448 VGND 0.0027f
C27518 VPWR.n5449 VGND 1.85e-19
C27519 VPWR.n5450 VGND 0.00336f
C27520 VPWR.n5451 VGND 0.00114f
C27521 VPWR.n5452 VGND 0.00149f
C27522 VPWR.n5453 VGND 0.00925f
C27523 VPWR.n5454 VGND 0.00199f
C27524 VPWR.n5455 VGND 0.00393f
C27525 VPWR.n5456 VGND 0.00393f
C27526 VPWR.n5457 VGND 0.00187f
C27527 VPWR.t295 VGND 0.00387f
C27528 VPWR.n5458 VGND 0.00493f
C27529 VPWR.n5459 VGND 0.0173f
C27530 VPWR.n5460 VGND 0.0103f
C27531 VPWR.t296 VGND 0.00387f
C27532 VPWR.n5461 VGND 0.0055f
C27533 VPWR.n5462 VGND 0.00837f
C27534 VPWR.n5463 VGND 0.0133f
C27535 VPWR.n5464 VGND 0.00393f
C27536 VPWR.n5465 VGND 0.0031f
C27537 VPWR.n5466 VGND 0.00295f
C27538 VPWR.t546 VGND 0.00387f
C27539 VPWR.t368 VGND 0.0046f
C27540 VPWR.n5467 VGND 0.0115f
C27541 VPWR.n5468 VGND 0.00342f
C27542 VPWR.n5469 VGND 0.00393f
C27543 VPWR.n5470 VGND 0.0136f
C27544 VPWR.n5471 VGND 0.00524f
C27545 VPWR.t3448 VGND 0.0274f
C27546 VPWR.n5472 VGND 0.0287f
C27547 VPWR.n5473 VGND 0.0233f
C27548 VPWR.n5474 VGND 0.0136f
C27549 VPWR.n5475 VGND 0.00524f
C27550 VPWR.n5476 VGND 0.0142f
C27551 VPWR.n5477 VGND 0.00524f
C27552 VPWR.t3485 VGND 0.0592f
C27553 VPWR.n5478 VGND 0.0416f
C27554 VPWR.n5479 VGND 0.0136f
C27555 VPWR.n5480 VGND 0.00524f
C27556 VPWR.n5481 VGND 0.00524f
C27557 VPWR.n5482 VGND 0.00524f
C27558 VPWR.n5483 VGND 0.0031f
C27559 VPWR.n5484 VGND 0.00179f
C27560 VPWR.n5485 VGND 0.00629f
C27561 VPWR.n5486 VGND 0.0121f
C27562 VPWR.n5487 VGND 0.00475f
C27563 VPWR.n5488 VGND 0.00393f
C27564 VPWR.n5489 VGND 0.0056f
C27565 VPWR.n5490 VGND 0.0058f
C27566 VPWR.n5491 VGND 0.00147f
C27567 VPWR.n5492 VGND 0.00179f
C27568 VPWR.n5493 VGND 0.00265f
C27569 VPWR.n5494 VGND 0.00556f
C27570 VPWR.n5495 VGND 0.00639f
C27571 VPWR.n5496 VGND 0.00453f
C27572 VPWR.n5497 VGND 0.00305f
C27573 VPWR.n5498 VGND 3.7e-19
C27574 VPWR.n5499 VGND 4.66e-19
C27575 VPWR.n5500 VGND 3.7e-19
C27576 VPWR.n5501 VGND 4.66e-19
C27577 VPWR.n5502 VGND 3.7e-19
C27578 VPWR.n5503 VGND 0.00154f
C27579 VPWR.n5504 VGND 5.12e-19
C27580 VPWR.n5505 VGND 5.41e-19
C27581 VPWR.n5506 VGND 5.12e-19
C27582 VPWR.n5507 VGND 4.27e-19
C27583 VPWR.n5508 VGND 2.85e-19
C27584 VPWR.n5509 VGND 0.00125f
C27585 VPWR.n5510 VGND 5.98e-19
C27586 VPWR.t1384 VGND 0.00633f
C27587 VPWR.n5511 VGND 0.0121f
C27588 VPWR.t3500 VGND 0.0592f
C27589 VPWR.n5512 VGND 0.0353f
C27590 VPWR.n5513 VGND 0.00197f
C27591 VPWR.n5514 VGND 6.99e-19
C27592 VPWR.n5515 VGND 0.00218f
C27593 VPWR.n5516 VGND 0.00137f
C27594 VPWR.n5517 VGND 5.92e-19
C27595 VPWR.n5518 VGND 5.05e-19
C27596 VPWR.n5519 VGND 4.17e-19
C27597 VPWR.n5520 VGND 5.48e-19
C27598 VPWR.n5522 VGND 8.67e-19
C27599 VPWR.n5523 VGND 6.54e-19
C27600 VPWR.n5524 VGND 9.06e-19
C27601 VPWR.n5525 VGND 3.95e-19
C27602 VPWR.n5526 VGND 3.95e-19
C27603 VPWR.n5527 VGND 7.68e-19
C27604 VPWR.n5528 VGND 5.05e-19
C27605 VPWR.n5529 VGND 8.11e-19
C27606 VPWR.n5530 VGND 3.95e-19
C27607 VPWR.n5531 VGND 1.77e-19
C27608 VPWR.n5532 VGND 1.76e-19
C27609 VPWR.n5533 VGND 5.48e-19
C27610 VPWR.n5534 VGND 0.00138f
C27611 VPWR.n5535 VGND 0.0057f
C27612 VPWR.n5537 VGND 6.14e-19
C27613 VPWR.n5538 VGND 4.39e-19
C27614 VPWR.n5539 VGND 1.76e-19
C27615 VPWR.n5540 VGND 4.83e-19
C27616 VPWR.n5541 VGND 2.41e-19
C27617 VPWR.n5542 VGND 3.73e-19
C27618 VPWR.n5543 VGND 3.07e-19
C27619 VPWR.n5544 VGND 4.11e-19
C27620 VPWR.n5545 VGND 4.11e-19
C27621 VPWR.n5546 VGND 7.39e-19
C27622 VPWR.n5547 VGND 5.19e-19
C27623 VPWR.n5548 VGND 7.39e-19
C27624 VPWR.n5549 VGND 4.11e-19
C27625 VPWR.n5550 VGND 4.11e-19
C27626 VPWR.n5551 VGND 2.85e-19
C27627 VPWR.n5552 VGND 3.95e-19
C27628 VPWR.n5553 VGND 2.85e-19
C27629 VPWR.n5554 VGND 4.83e-19
C27630 VPWR.n5555 VGND 4.17e-19
C27631 VPWR.n5556 VGND 5.05e-19
C27632 VPWR.n5557 VGND 6.55e-19
C27633 VPWR.n5558 VGND 5.41e-19
C27634 VPWR.n5559 VGND 9.96e-19
C27635 VPWR.n5560 VGND 9.68e-19
C27636 VPWR.n5561 VGND 5.12e-19
C27637 VPWR.t3076 VGND 0.00676f
C27638 VPWR.n5562 VGND 0.0115f
C27639 VPWR.n5563 VGND 0.00323f
C27640 VPWR.n5564 VGND 3.13e-19
C27641 VPWR.n5565 VGND 6.26e-19
C27642 VPWR.n5566 VGND 5.12e-19
C27643 VPWR.n5567 VGND 0.00108f
C27644 VPWR.n5568 VGND 0.00122f
C27645 VPWR.n5569 VGND 3.13e-19
C27646 VPWR.n5570 VGND 5.12e-19
C27647 VPWR.n5571 VGND 0.0033f
C27648 VPWR.n5572 VGND 5.98e-19
C27649 VPWR.n5573 VGND 6.1e-19
C27650 VPWR.n5574 VGND 2.28e-19
C27651 VPWR.n5575 VGND 3.14e-19
C27652 VPWR.n5576 VGND 0.00126f
C27653 VPWR.n5577 VGND 0.00256f
C27654 VPWR.t2912 VGND 0.00239f
C27655 VPWR.n5578 VGND 0.00618f
C27656 VPWR.n5579 VGND 0.00535f
C27657 VPWR.n5580 VGND 0.00492f
C27658 VPWR.t2829 VGND 6.73e-19
C27659 VPWR.t3078 VGND 0.00127f
C27660 VPWR.n5581 VGND 0.00203f
C27661 VPWR.n5582 VGND 0.00594f
C27662 VPWR.n5583 VGND 0.00377f
C27663 VPWR.n5584 VGND 0.00524f
C27664 VPWR.n5585 VGND 0.00614f
C27665 VPWR.n5586 VGND 0.00524f
C27666 VPWR.n5587 VGND 0.00639f
C27667 VPWR.n5588 VGND 0.00524f
C27668 VPWR.n5589 VGND 0.0031f
C27669 VPWR.n5590 VGND 0.00282f
C27670 VPWR.n5591 VGND 0.00918f
C27671 VPWR.n5592 VGND 0.00562f
C27672 VPWR.n5593 VGND 0.00126f
C27673 VPWR.n5594 VGND 0.00199f
C27674 VPWR.n5595 VGND 0.00903f
C27675 VPWR.n5596 VGND 0.0113f
C27676 VPWR.n5597 VGND 0.0104f
C27677 VPWR.t2469 VGND 0.00234f
C27678 VPWR.n5598 VGND 0.00986f
C27679 VPWR.n5599 VGND 0.00829f
C27680 VPWR.n5600 VGND 0.00524f
C27681 VPWR.n5601 VGND 0.0119f
C27682 VPWR.n5602 VGND 0.00524f
C27683 VPWR.n5603 VGND 0.0031f
C27684 VPWR.n5604 VGND 0.00483f
C27685 VPWR.n5605 VGND 0.00592f
C27686 VPWR.n5606 VGND 0.00755f
C27687 VPWR.n5607 VGND 0.00152f
C27688 VPWR.n5608 VGND 0.00179f
C27689 VPWR.n5609 VGND 0.00186f
C27690 VPWR.n5610 VGND 0.00393f
C27691 VPWR.n5611 VGND 0.00333f
C27692 VPWR.n5612 VGND 0.00135f
C27693 VPWR.n5613 VGND 0.00748f
C27694 VPWR.t322 VGND 0.0046f
C27695 VPWR.n5614 VGND 0.00407f
C27696 VPWR.n5615 VGND 0.00135f
C27697 VPWR.n5616 VGND 0.00393f
C27698 VPWR.n5617 VGND 0.00639f
C27699 VPWR.n5618 VGND 0.00524f
C27700 VPWR.n5619 VGND 0.0031f
C27701 VPWR.n5620 VGND 0.00182f
C27702 VPWR.n5621 VGND 0.00506f
C27703 VPWR.n5622 VGND 0.0356f
C27704 VPWR.n5623 VGND 0.00463f
C27705 VPWR.n5624 VGND 0.00473f
C27706 VPWR.n5625 VGND 0.00393f
C27707 VPWR.n5626 VGND 0.00199f
C27708 VPWR.n5627 VGND 0.00629f
C27709 VPWR.t46 VGND 0.00387f
C27710 VPWR.n5628 VGND 0.0107f
C27711 VPWR.n5629 VGND 0.00796f
C27712 VPWR.n5630 VGND 0.00393f
C27713 VPWR.t3372 VGND 0.0231f
C27714 VPWR.n5631 VGND 0.043f
C27715 VPWR.n5632 VGND 0.00524f
C27716 VPWR.n5633 VGND 0.00524f
C27717 VPWR.n5634 VGND 0.00524f
C27718 VPWR.n5635 VGND 0.0031f
C27719 VPWR.n5636 VGND 0.0125f
C27720 VPWR.t47 VGND 0.004f
C27721 VPWR.n5637 VGND 0.00668f
C27722 VPWR.n5638 VGND 0.00249f
C27723 VPWR.n5639 VGND 0.00262f
C27724 VPWR.n5640 VGND 0.00199f
C27725 VPWR.n5641 VGND 0.00179f
C27726 VPWR.n5642 VGND 0.0066f
C27727 VPWR.n5643 VGND 0.00506f
C27728 VPWR.n5644 VGND 0.00475f
C27729 VPWR.t3392 VGND 0.0592f
C27730 VPWR.n5645 VGND 0.0356f
C27731 VPWR.t3168 VGND 0.00102f
C27732 VPWR.t1198 VGND 0.00154f
C27733 VPWR.n5646 VGND 0.00483f
C27734 VPWR.n5647 VGND 0.00908f
C27735 VPWR.n5648 VGND 0.00269f
C27736 VPWR.n5649 VGND 0.00524f
C27737 VPWR.n5650 VGND 0.00545f
C27738 VPWR.n5651 VGND 0.00524f
C27739 VPWR.n5652 VGND 0.00635f
C27740 VPWR.n5653 VGND 0.0039f
C27741 VPWR.n5654 VGND 3.95e-19
C27742 VPWR.n5655 VGND 5.05e-19
C27743 VPWR.n5656 VGND 5.05e-19
C27744 VPWR.n5657 VGND 0.00139f
C27745 VPWR.n5658 VGND 9.06e-19
C27746 VPWR.n5659 VGND 5.48e-19
C27747 VPWR.n5660 VGND 3.07e-19
C27748 VPWR.n5661 VGND 1.76e-19
C27749 VPWR.n5662 VGND 2.63e-19
C27750 VPWR.n5663 VGND 9.42e-19
C27751 VPWR.n5664 VGND 0.00131f
C27752 VPWR.n5665 VGND 6.26e-19
C27753 VPWR.n5666 VGND 3.42e-19
C27754 VPWR.n5667 VGND 4.84e-19
C27755 VPWR.n5668 VGND 0.0033f
C27756 VPWR.n5669 VGND 5.98e-19
C27757 VPWR.n5670 VGND 5.38e-19
C27758 VPWR.n5671 VGND 4.27e-19
C27759 VPWR.n5672 VGND 5.74e-19
C27760 VPWR.n5673 VGND 4.55e-19
C27761 VPWR.n5674 VGND 0.00248f
C27762 VPWR.n5675 VGND 4.84e-19
C27763 VPWR.n5676 VGND 6.83e-19
C27764 VPWR.n5677 VGND 4.84e-19
C27765 VPWR.n5678 VGND 3.13e-19
C27766 VPWR.n5679 VGND 9.96e-19
C27767 VPWR.n5680 VGND 0.00258f
C27768 VPWR.n5681 VGND 9.68e-19
C27769 VPWR.n5682 VGND 4.27e-19
C27770 VPWR.n5683 VGND 2.56e-19
C27771 VPWR.t2892 VGND 0.00676f
C27772 VPWR.n5684 VGND 0.00917f
C27773 VPWR.n5685 VGND 2.15e-19
C27774 VPWR.n5686 VGND 0.00319f
C27775 VPWR.n5687 VGND 3.42e-19
C27776 VPWR.n5688 VGND 7.4e-19
C27777 VPWR.n5689 VGND 5.41e-19
C27778 VPWR.n5690 VGND 9.96e-19
C27779 VPWR.n5691 VGND 9.68e-19
C27780 VPWR.n5692 VGND 3.7e-19
C27781 VPWR.n5693 VGND 6.83e-19
C27782 VPWR.n5694 VGND 0.00323f
C27783 VPWR.n5695 VGND 4.27e-19
C27784 VPWR.n5696 VGND 8.54e-20
C27785 VPWR.n5697 VGND 6.1e-19
C27786 VPWR.n5698 VGND 4.27e-19
C27787 VPWR.n5699 VGND 0.00126f
C27788 VPWR.n5700 VGND 0.00156f
C27789 VPWR.n5701 VGND 0.00203f
C27790 VPWR.n5702 VGND 0.00138f
C27791 VPWR.n5703 VGND 6.14e-19
C27792 VPWR.n5704 VGND 5.48e-19
C27793 VPWR.n5705 VGND 0.00138f
C27794 VPWR.n5706 VGND 0.0057f
C27795 VPWR.n5707 VGND 6.54e-19
C27796 VPWR.n5708 VGND 8.67e-19
C27797 VPWR.n5709 VGND 3.51e-19
C27798 VPWR.n5710 VGND 4.61e-19
C27799 VPWR.n5711 VGND 5.27e-19
C27800 VPWR.n5712 VGND 2.85e-19
C27801 VPWR.n5713 VGND 2.85e-19
C27802 VPWR.n5714 VGND 4.17e-19
C27803 VPWR.n5715 VGND 4.11e-19
C27804 VPWR.n5716 VGND 4.11e-19
C27805 VPWR.n5717 VGND 7.39e-19
C27806 VPWR.n5718 VGND 5.19e-19
C27807 VPWR.n5719 VGND 7.39e-19
C27808 VPWR.n5720 VGND 4.11e-19
C27809 VPWR.n5721 VGND 5.27e-19
C27810 VPWR.n5722 VGND 3.73e-19
C27811 VPWR.n5723 VGND 2.41e-19
C27812 VPWR.n5724 VGND 4.83e-19
C27813 VPWR.n5725 VGND 4.17e-19
C27814 VPWR.n5726 VGND 5.71e-19
C27815 VPWR.n5727 VGND 4.17e-19
C27816 VPWR.n5728 VGND 4.83e-19
C27817 VPWR.n5729 VGND 4.61e-19
C27818 VPWR.n5730 VGND 4.61e-19
C27819 VPWR.n5731 VGND 4.11e-19
C27820 VPWR.n5733 VGND 0.1f
C27821 VPWR.n5734 VGND 0.1f
C27822 VPWR.n5736 VGND 9.06e-19
C27823 VPWR.n5737 VGND 5.48e-19
C27824 VPWR.n5738 VGND 3.07e-19
C27825 VPWR.n5739 VGND 1.76e-19
C27826 VPWR.n5740 VGND 2.63e-19
C27827 VPWR.n5741 VGND 9.42e-19
C27828 VPWR.n5742 VGND 8.27e-19
C27829 VPWR.n5743 VGND 0.0031f
C27830 VPWR.n5744 VGND 0.00517f
C27831 VPWR.n5745 VGND 8.14e-19
C27832 VPWR.n5746 VGND 5.98e-19
C27833 VPWR.n5747 VGND 1.51e-19
C27834 VPWR.n5748 VGND 4.27e-19
C27835 VPWR.n5749 VGND 1.61e-19
C27836 VPWR.n5750 VGND 4.55e-19
C27837 VPWR.n5751 VGND 4.94e-19
C27838 VPWR.n5752 VGND 2.56e-19
C27839 VPWR.n5753 VGND 6.55e-19
C27840 VPWR.n5754 VGND 5.27e-19
C27841 VPWR.n5755 VGND 2.41e-19
C27842 VPWR.n5756 VGND 3.73e-19
C27843 VPWR.n5757 VGND 4.84e-19
C27844 VPWR.n5758 VGND 1.71e-19
C27845 VPWR.n5759 VGND 8.83e-19
C27846 VPWR.n5760 VGND 9.68e-19
C27847 VPWR.n5761 VGND 4.7e-19
C27848 VPWR.t2776 VGND 0.00692f
C27849 VPWR.n5762 VGND 0.0108f
C27850 VPWR.n5763 VGND 2.14e-19
C27851 VPWR.n5764 VGND 3.42e-19
C27852 VPWR.n5765 VGND 3.29e-19
C27853 VPWR.n5766 VGND 4.39e-19
C27854 VPWR.n5767 VGND 9e-19
C27855 VPWR.n5768 VGND 8.67e-19
C27856 VPWR.n5769 VGND 6.54e-19
C27857 VPWR.n5770 VGND 9.06e-19
C27858 VPWR.n5771 VGND 0.00138f
C27859 VPWR.n5772 VGND 5.48e-19
C27860 VPWR.n5773 VGND 6.14e-19
C27861 VPWR.t2530 VGND 0.00166f
C27862 VPWR.t1265 VGND 0.00225f
C27863 VPWR.n5774 VGND 0.00438f
C27864 VPWR.t1376 VGND 6.73e-19
C27865 VPWR.t2774 VGND 0.00127f
C27866 VPWR.n5775 VGND 0.00203f
C27867 VPWR.n5776 VGND 0.0035f
C27868 VPWR.n5777 VGND 0.00555f
C27869 VPWR.t1259 VGND 0.00166f
C27870 VPWR.t1261 VGND 0.00166f
C27871 VPWR.n5778 VGND 0.00345f
C27872 VPWR.n5779 VGND 0.00502f
C27873 VPWR.t1263 VGND 0.00682f
C27874 VPWR.n5780 VGND 0.00711f
C27875 VPWR.t2357 VGND 0.00453f
C27876 VPWR.t880 VGND 0.00654f
C27877 VPWR.t2975 VGND 0.00238f
C27878 VPWR.n5781 VGND 0.0053f
C27879 VPWR.t1815 VGND 0.00102f
C27880 VPWR.t1766 VGND 0.00102f
C27881 VPWR.n5782 VGND 0.00221f
C27882 VPWR.n5783 VGND 0.00563f
C27883 VPWR.t1652 VGND 0.00137f
C27884 VPWR.t3238 VGND -2.18e-20
C27885 VPWR.n5784 VGND 0.00629f
C27886 VPWR.t3240 VGND 0.00663f
C27887 VPWR.n5785 VGND 0.00848f
C27888 VPWR.t3533 VGND 0.00911f
C27889 VPWR.t739 VGND 0.00391f
C27890 VPWR.n5786 VGND 0.0253f
C27891 VPWR.t738 VGND 0.00391f
C27892 VPWR.n5788 VGND 0.0138f
C27893 VPWR.t3387 VGND 0.00911f
C27894 VPWR.t504 VGND 0.00391f
C27895 VPWR.n5789 VGND 0.0253f
C27896 VPWR.t505 VGND 0.00391f
C27897 VPWR.n5791 VGND 0.0138f
C27898 VPWR.n5792 VGND 0.0109f
C27899 VPWR.n5793 VGND 0.00444f
C27900 VPWR.n5794 VGND 0.0031f
C27901 VPWR.n5795 VGND 0.00524f
C27902 VPWR.n5796 VGND 0.00475f
C27903 VPWR.n5797 VGND 0.00759f
C27904 VPWR.n5798 VGND 0.00115f
C27905 VPWR.n5799 VGND 0.00179f
C27906 VPWR.n5800 VGND 0.00307f
C27907 VPWR.n5801 VGND 0.0014f
C27908 VPWR.n5802 VGND 0.00524f
C27909 VPWR.n5803 VGND 0.00393f
C27910 VPWR.n5804 VGND 0.0111f
C27911 VPWR.n5805 VGND 0.00158f
C27912 VPWR.n5806 VGND 0.0031f
C27913 VPWR.n5807 VGND 0.00142f
C27914 VPWR.n5808 VGND 0.00524f
C27915 VPWR.t3106 VGND 0.00184f
C27916 VPWR.t1800 VGND 0.00166f
C27917 VPWR.n5809 VGND 0.00358f
C27918 VPWR.t1382 VGND 6.73e-19
C27919 VPWR.t1273 VGND 9.96e-19
C27920 VPWR.n5810 VGND 0.00176f
C27921 VPWR.n5811 VGND 0.00418f
C27922 VPWR.n5812 VGND 0.00239f
C27923 VPWR.n5813 VGND 9.58e-19
C27924 VPWR.n5814 VGND 0.00524f
C27925 VPWR.n5815 VGND 0.00393f
C27926 VPWR.n5816 VGND 0.00155f
C27927 VPWR.n5817 VGND 0.00562f
C27928 VPWR.n5818 VGND 4.03e-19
C27929 VPWR.n5819 VGND 0.00393f
C27930 VPWR.n5820 VGND 0.00151f
C27931 VPWR.n5821 VGND 0.00524f
C27932 VPWR.n5822 VGND 0.00524f
C27933 VPWR.n5823 VGND 0.00145f
C27934 VPWR.n5824 VGND 0.00524f
C27935 VPWR.n5825 VGND 0.00475f
C27936 VPWR.n5826 VGND 9.88e-19
C27937 VPWR.n5827 VGND 0.00117f
C27938 VPWR.n5828 VGND 0.00154f
C27939 VPWR.n5829 VGND 9.06e-19
C27940 VPWR.n5830 VGND 0.00138f
C27941 VPWR.n5831 VGND 5.98e-19
C27942 VPWR.t1005 VGND 0.00242f
C27943 VPWR.n5832 VGND 0.00484f
C27944 VPWR.n5833 VGND 7.12e-19
C27945 VPWR.n5834 VGND 5.04e-20
C27946 VPWR.n5835 VGND 4.27e-19
C27947 VPWR.n5836 VGND 8.54e-20
C27948 VPWR.n5837 VGND 6.65e-19
C27949 VPWR.n5838 VGND 4.27e-19
C27950 VPWR.n5839 VGND 6.83e-19
C27951 VPWR.n5840 VGND 3.7e-19
C27952 VPWR.n5841 VGND 9.68e-19
C27953 VPWR.n5842 VGND 9.96e-19
C27954 VPWR.n5843 VGND 5.41e-19
C27955 VPWR.n5844 VGND 7.4e-19
C27956 VPWR.n5845 VGND 5.71e-19
C27957 VPWR.n5846 VGND 4.17e-19
C27958 VPWR.n5847 VGND 4.83e-19
C27959 VPWR.n5848 VGND 4.61e-19
C27960 VPWR.n5849 VGND 4.61e-19
C27961 VPWR.n5850 VGND 4.11e-19
C27962 VPWR.n5852 VGND 0.071f
C27963 VPWR.n5853 VGND 0.0976f
C27964 VPWR.n5854 VGND 0.564f
C27965 VPWR.n5855 VGND 0.746f
C27966 VPWR.n5856 VGND 0.0976f
C27967 VPWR.n5857 VGND 0.0323f
C27968 VPWR.n5858 VGND 0.00139f
C27969 VPWR.n5859 VGND 9.06e-19
C27970 VPWR.t1224 VGND 7.22e-19
C27971 VPWR.t1281 VGND 9.22e-19
C27972 VPWR.n5860 VGND 0.00189f
C27973 VPWR.n5861 VGND 0.00152f
C27974 VPWR.n5862 VGND 0.00231f
C27975 VPWR.t3097 VGND 0.0321f
C27976 VPWR.t3095 VGND 0.0186f
C27977 VPWR.t1480 VGND 0.0144f
C27978 VPWR.t3093 VGND 0.0141f
C27979 VPWR.t1478 VGND 0.0144f
C27980 VPWR.t3091 VGND 0.0141f
C27981 VPWR.t1482 VGND 0.0161f
C27982 VPWR.t3310 VGND 0.0141f
C27983 VPWR.t1484 VGND 0.00537f
C27984 VPWR.t3265 VGND 0.0153f
C27985 VPWR.t1186 VGND 0.0217f
C27986 VPWR.t1225 VGND 0.0305f
C27987 VPWR.t219 VGND 0.0173f
C27988 VPWR.t3312 VGND 0.041f
C27989 VPWR.t2413 VGND 0.048f
C27990 VPWR.t1280 VGND 0.026f
C27991 VPWR.t1223 VGND 0.026f
C27992 VPWR.t1321 VGND 0.0386f
C27993 VPWR.t1219 VGND 0.0154f
C27994 VPWR.t1952 VGND 0.0052f
C27995 VPWR.t1221 VGND 0.0154f
C27996 VPWR.t568 VGND 0.0723f
C27997 VPWR.t397 VGND 0.0695f
C27998 VPWR.n5863 VGND 0.0705f
C27999 VPWR.n5864 VGND 0.00639f
C28000 VPWR.t140 VGND 0.00387f
C28001 VPWR.n5865 VGND 0.00542f
C28002 VPWR.t636 VGND 0.004f
C28003 VPWR.n5866 VGND 0.00705f
C28004 VPWR.t2249 VGND 0.00632f
C28005 VPWR.t3432 VGND 0.0289f
C28006 VPWR.t635 VGND 0.00387f
C28007 VPWR.n5867 VGND 0.0604f
C28008 VPWR.n5868 VGND 0.0146f
C28009 VPWR.t3575 VGND 0.0179f
C28010 VPWR.t694 VGND 0.00395f
C28011 VPWR.n5869 VGND 0.028f
C28012 VPWR.t695 VGND 0.00432f
C28013 VPWR.n5870 VGND 0.0303f
C28014 VPWR.n5871 VGND 0.0117f
C28015 VPWR.n5872 VGND 0.00966f
C28016 VPWR.t1547 VGND 0.0053f
C28017 VPWR.n5873 VGND 0.00394f
C28018 VPWR.t3552 VGND 0.00911f
C28019 VPWR.t232 VGND 0.00391f
C28020 VPWR.n5874 VGND 0.0253f
C28021 VPWR.t233 VGND 0.00391f
C28022 VPWR.n5876 VGND 0.0138f
C28023 VPWR.t3055 VGND 0.00166f
C28024 VPWR.t1545 VGND 0.00219f
C28025 VPWR.n5877 VGND 0.00445f
C28026 VPWR.n5878 VGND 0.00259f
C28027 VPWR.t2386 VGND 0.00597f
C28028 VPWR.n5879 VGND 0.0141f
C28029 VPWR.n5880 VGND 3.29e-19
C28030 VPWR.n5881 VGND 5.71e-19
C28031 VPWR.n5882 VGND 5.92e-19
C28032 VPWR.n5883 VGND 5.05e-19
C28033 VPWR.n5884 VGND 8.67e-19
C28034 VPWR.n5885 VGND 6.54e-19
C28035 VPWR.n5886 VGND 9.06e-19
C28036 VPWR.n5887 VGND 0.0323f
C28037 VPWR.n5889 VGND 6.54e-19
C28038 VPWR.n5890 VGND 8.67e-19
C28039 VPWR.n5891 VGND 3.95e-19
C28040 VPWR.n5892 VGND 4.61e-19
C28041 VPWR.n5893 VGND 2.41e-19
C28042 VPWR.n5894 VGND 3.95e-19
C28043 VPWR.n5895 VGND 5.05e-19
C28044 VPWR.n5896 VGND 4.17e-19
C28045 VPWR.n5897 VGND 6.14e-19
C28046 VPWR.n5898 VGND 4.39e-19
C28047 VPWR.n5899 VGND 1.76e-19
C28048 VPWR.n5900 VGND 3.07e-19
C28049 VPWR.n5901 VGND 4.83e-19
C28050 VPWR.n5902 VGND 2.85e-19
C28051 VPWR.n5903 VGND 3.95e-19
C28052 VPWR.n5904 VGND 3.95e-19
C28053 VPWR.n5905 VGND 4.17e-19
C28054 VPWR.n5906 VGND 2.85e-19
C28055 VPWR.n5907 VGND 2.85e-19
C28056 VPWR.n5908 VGND 4.11e-19
C28057 VPWR.n5909 VGND 4.11e-19
C28058 VPWR.n5910 VGND 7.39e-19
C28059 VPWR.n5911 VGND 5.19e-19
C28060 VPWR.n5912 VGND 7.39e-19
C28061 VPWR.n5913 VGND 4.11e-19
C28062 VPWR.n5914 VGND 4.11e-19
C28063 VPWR.n5916 VGND 8.67e-19
C28064 VPWR.n5917 VGND 6.54e-19
C28065 VPWR.n5918 VGND 9.06e-19
C28066 VPWR.n5919 VGND 3.29e-19
C28067 VPWR.n5920 VGND 5.71e-19
C28068 VPWR.n5921 VGND 5.92e-19
C28069 VPWR.n5922 VGND 5.05e-19
C28070 VPWR.n5923 VGND 6.78e-19
C28071 VPWR.t115 VGND 0.00387f
C28072 VPWR.n5924 VGND 0.00837f
C28073 VPWR.t194 VGND 0.00387f
C28074 VPWR.t3421 VGND 0.0231f
C28075 VPWR.t1615 VGND 0.00234f
C28076 VPWR.n5925 VGND 0.00986f
C28077 VPWR.n5926 VGND 0.00829f
C28078 VPWR.n5927 VGND 0.0384f
C28079 VPWR.n5928 VGND 0.00837f
C28080 VPWR.n5929 VGND 0.00525f
C28081 VPWR.t195 VGND 0.00387f
C28082 VPWR.n5930 VGND 0.0083f
C28083 VPWR.t1961 VGND 0.00102f
C28084 VPWR.t1917 VGND 0.00102f
C28085 VPWR.n5931 VGND 0.00208f
C28086 VPWR.n5932 VGND 0.00294f
C28087 VPWR.n5933 VGND 0.00134f
C28088 VPWR.t2553 VGND 0.00676f
C28089 VPWR.n5934 VGND 0.00956f
C28090 VPWR.n5935 VGND 0.0216f
C28091 VPWR.t2849 VGND 6.73e-19
C28092 VPWR.t2551 VGND 0.00127f
C28093 VPWR.n5936 VGND 0.00203f
C28094 VPWR.t499 VGND 0.00387f
C28095 VPWR.n5937 VGND 0.00493f
C28096 VPWR.n5938 VGND 0.00525f
C28097 VPWR.t2394 VGND 0.00453f
C28098 VPWR.t3451 VGND 0.0179f
C28099 VPWR.n5939 VGND 0.0173f
C28100 VPWR.n5940 VGND 0.0103f
C28101 VPWR.n5941 VGND 0.00912f
C28102 VPWR.n5942 VGND 0.0111f
C28103 VPWR.t500 VGND 0.00387f
C28104 VPWR.n5943 VGND 0.00613f
C28105 VPWR.t10 VGND 0.0046f
C28106 VPWR.t2833 VGND 6.73e-19
C28107 VPWR.t2207 VGND 9.96e-19
C28108 VPWR.n5944 VGND 0.00176f
C28109 VPWR.n5945 VGND 0.00636f
C28110 VPWR.n5946 VGND 0.00231f
C28111 VPWR.t2489 VGND 0.00102f
C28112 VPWR.t1832 VGND 0.00102f
C28113 VPWR.n5947 VGND 0.00217f
C28114 VPWR.n5948 VGND 0.0071f
C28115 VPWR.t11 VGND 0.0046f
C28116 VPWR.n5949 VGND 0.00407f
C28117 VPWR.n5950 VGND 0.00137f
C28118 VPWR.t2683 VGND 0.00166f
C28119 VPWR.t3114 VGND 0.00184f
C28120 VPWR.n5951 VGND 0.00361f
C28121 VPWR.t1176 VGND 0.00692f
C28122 VPWR.n5952 VGND 0.0128f
C28123 VPWR.n5953 VGND 4.83e-19
C28124 VPWR.n5954 VGND 2.41e-19
C28125 VPWR.n5955 VGND 3.73e-19
C28126 VPWR.n5956 VGND 6.54e-19
C28127 VPWR.n5957 VGND 8.67e-19
C28128 VPWR.n5958 VGND 0.00139f
C28129 VPWR.n5959 VGND 9.06e-19
C28130 VPWR.n5960 VGND 0.00137f
C28131 VPWR.n5961 VGND 5.92e-19
C28132 VPWR.t2573 VGND 0.00102f
C28133 VPWR.t2090 VGND 0.00102f
C28134 VPWR.n5962 VGND 0.00217f
C28135 VPWR.n5963 VGND 0.00688f
C28136 VPWR.t168 VGND 0.0046f
C28137 VPWR.n5964 VGND 0.004f
C28138 VPWR.n5965 VGND 0.00199f
C28139 VPWR.n5966 VGND 0.011f
C28140 VPWR.t705 VGND 0.0046f
C28141 VPWR.n5967 VGND 0.00644f
C28142 VPWR.n5968 VGND 0.00535f
C28143 VPWR.t488 VGND 0.00462f
C28144 VPWR.n5969 VGND 0.0148f
C28145 VPWR.n5970 VGND 0.00861f
C28146 VPWR.n5971 VGND 6.26e-19
C28147 VPWR.n5972 VGND 3.95e-19
C28148 VPWR.n5973 VGND 4.61e-19
C28149 VPWR.n5974 VGND 2.41e-19
C28150 VPWR.n5975 VGND 3.95e-19
C28151 VPWR.n5976 VGND 6.54e-19
C28152 VPWR.n5977 VGND 8.67e-19
C28153 VPWR.n5978 VGND 8.11e-19
C28154 VPWR.n5979 VGND 3.95e-19
C28155 VPWR.n5980 VGND 1.77e-19
C28156 VPWR.n5981 VGND 3.95e-19
C28157 VPWR.n5982 VGND 7.68e-19
C28158 VPWR.n5983 VGND 5.05e-19
C28159 VPWR.n5984 VGND 1.76e-19
C28160 VPWR.n5985 VGND 9.06e-19
C28161 VPWR.n5986 VGND 5.48e-19
C28162 VPWR.n5987 VGND 0.00138f
C28163 VPWR.n5988 VGND 0.0057f
C28164 VPWR.n5989 VGND 4.83e-19
C28165 VPWR.n5990 VGND 2.85e-19
C28166 VPWR.n5991 VGND 3.95e-19
C28167 VPWR.n5992 VGND 4.17e-19
C28168 VPWR.n5993 VGND 2.85e-19
C28169 VPWR.n5994 VGND 2.85e-19
C28170 VPWR.n5995 VGND 4.11e-19
C28171 VPWR.n5996 VGND 8.67e-19
C28172 VPWR.n5997 VGND 6.54e-19
C28173 VPWR.n5998 VGND 9.06e-19
C28174 VPWR.n5999 VGND 0.00139f
C28175 VPWR.n6000 VGND 3.95e-19
C28176 VPWR.n6001 VGND 3.29e-19
C28177 VPWR.n6002 VGND 5.71e-19
C28178 VPWR.n6003 VGND 5.92e-19
C28179 VPWR.n6004 VGND 5.05e-19
C28180 VPWR.t3369 VGND 0.0592f
C28181 VPWR.n6005 VGND 0.038f
C28182 VPWR.n6006 VGND 0.00833f
C28183 VPWR.n6007 VGND 0.00503f
C28184 VPWR.n6008 VGND 0.0106f
C28185 VPWR.t714 VGND 0.0046f
C28186 VPWR.n6009 VGND 0.00644f
C28187 VPWR.t2316 VGND 0.00239f
C28188 VPWR.n6010 VGND 0.00421f
C28189 VPWR.t1356 VGND 0.00692f
C28190 VPWR.t2500 VGND 0.00102f
C28191 VPWR.t2203 VGND 0.00154f
C28192 VPWR.n6011 VGND 0.00483f
C28193 VPWR.n6012 VGND 0.00887f
C28194 VPWR.t305 VGND 0.0046f
C28195 VPWR.n6013 VGND 0.00192f
C28196 VPWR.n6014 VGND 0.00556f
C28197 VPWR.t3472 VGND 0.00911f
C28198 VPWR.t334 VGND 0.00391f
C28199 VPWR.n6015 VGND 0.0253f
C28200 VPWR.t335 VGND 0.00391f
C28201 VPWR.n6017 VGND 0.0138f
C28202 VPWR.t32 VGND 0.0046f
C28203 VPWR.n6018 VGND 0.00644f
C28204 VPWR.t633 VGND 0.0046f
C28205 VPWR.n6019 VGND 0.00644f
C28206 VPWR.n6020 VGND 0.0113f
C28207 VPWR.n6021 VGND 0.00524f
C28208 VPWR.n6022 VGND 0.0113f
C28209 VPWR.n6023 VGND 0.00524f
C28210 VPWR.n6024 VGND 0.011f
C28211 VPWR.n6025 VGND 0.00524f
C28212 VPWR.n6026 VGND 0.0031f
C28213 VPWR.n6027 VGND 0.00516f
C28214 VPWR.t304 VGND 0.0046f
C28215 VPWR.n6028 VGND 0.0106f
C28216 VPWR.n6029 VGND 0.00644f
C28217 VPWR.n6030 VGND 0.00512f
C28218 VPWR.n6031 VGND 0.00475f
C28219 VPWR.n6032 VGND 0.00524f
C28220 VPWR.n6033 VGND 0.0031f
C28221 VPWR.n6034 VGND 0.00535f
C28222 VPWR.t3424 VGND 0.0592f
C28223 VPWR.n6035 VGND 0.0356f
C28224 VPWR.n6036 VGND 0.00487f
C28225 VPWR.n6037 VGND 0.00475f
C28226 VPWR.t2973 VGND 0.00136f
C28227 VPWR.t2233 VGND 0.00136f
C28228 VPWR.n6038 VGND 0.00317f
C28229 VPWR.n6039 VGND 0.0103f
C28230 VPWR.n6040 VGND 0.00524f
C28231 VPWR.n6041 VGND 0.0031f
C28232 VPWR.n6042 VGND 0.00442f
C28233 VPWR.n6043 VGND 0.00854f
C28234 VPWR.n6044 VGND 0.0164f
C28235 VPWR.n6045 VGND 0.00556f
C28236 VPWR.n6046 VGND 0.00393f
C28237 VPWR.n6047 VGND 0.00545f
C28238 VPWR.n6048 VGND 0.00524f
C28239 VPWR.n6049 VGND 0.0031f
C28240 VPWR.n6050 VGND 0.00274f
C28241 VPWR.n6051 VGND 0.0014f
C28242 VPWR.n6052 VGND 0.00475f
C28243 VPWR.n6053 VGND 0.0031f
C28244 VPWR.n6054 VGND 0.0109f
C28245 VPWR.n6055 VGND 0.00102f
C28246 VPWR.n6056 VGND 0.00199f
C28247 VPWR.t2835 VGND 6.73e-19
C28248 VPWR.t1358 VGND 0.00127f
C28249 VPWR.n6057 VGND 0.00207f
C28250 VPWR.n6058 VGND 0.00499f
C28251 VPWR.t2851 VGND 6.73e-19
C28252 VPWR.t1881 VGND 9.96e-19
C28253 VPWR.n6059 VGND 0.00176f
C28254 VPWR.n6060 VGND 0.0101f
C28255 VPWR.n6061 VGND 0.0102f
C28256 VPWR.n6062 VGND 0.0101f
C28257 VPWR.t599 VGND 0.00387f
C28258 VPWR.n6063 VGND 0.00837f
C28259 VPWR.t2220 VGND 0.00632f
C28260 VPWR.n6064 VGND 0.007f
C28261 VPWR.t2243 VGND 0.00234f
C28262 VPWR.n6065 VGND 0.00525f
C28263 VPWR.t3061 VGND 0.00102f
C28264 VPWR.t1836 VGND 0.00102f
C28265 VPWR.n6066 VGND 0.00217f
C28266 VPWR.t3435 VGND 0.0179f
C28267 VPWR.t238 VGND 0.00387f
C28268 VPWR.n6067 VGND 0.00493f
C28269 VPWR.n6068 VGND 0.0173f
C28270 VPWR.n6069 VGND 0.00359f
C28271 VPWR.n6070 VGND 0.0107f
C28272 VPWR.t239 VGND 0.00387f
C28273 VPWR.n6071 VGND 0.00133f
C28274 VPWR.n6072 VGND 0.00179f
C28275 VPWR.n6073 VGND 0.00179f
C28276 VPWR.n6074 VGND 0.00525f
C28277 VPWR.n6075 VGND 0.00837f
C28278 VPWR.n6076 VGND 0.0132f
C28279 VPWR.n6077 VGND 0.0031f
C28280 VPWR.n6078 VGND 0.00524f
C28281 VPWR.n6079 VGND 0.00393f
C28282 VPWR.n6080 VGND 0.00199f
C28283 VPWR.n6081 VGND 0.00154f
C28284 VPWR.n6082 VGND 0.00391f
C28285 VPWR.n6083 VGND 2.12e-19
C28286 VPWR.n6084 VGND 0.0031f
C28287 VPWR.n6085 VGND 0.00158f
C28288 VPWR.n6086 VGND 0.00524f
C28289 VPWR.n6087 VGND 0.00393f
C28290 VPWR.t2218 VGND 0.0065f
C28291 VPWR.n6088 VGND 0.00754f
C28292 VPWR.n6089 VGND 0.00504f
C28293 VPWR.n6090 VGND 0.0031f
C28294 VPWR.n6091 VGND 0.00524f
C28295 VPWR.n6092 VGND 0.00524f
C28296 VPWR.n6093 VGND 0.0115f
C28297 VPWR.n6094 VGND 0.00524f
C28298 VPWR.t2728 VGND 0.00453f
C28299 VPWR.n6095 VGND 0.0116f
C28300 VPWR.n6096 VGND 0.00912f
C28301 VPWR.n6097 VGND 0.00524f
C28302 VPWR.t3561 VGND 0.0282f
C28303 VPWR.n6098 VGND 0.0489f
C28304 VPWR.n6099 VGND 0.0102f
C28305 VPWR.n6100 VGND 0.00524f
C28306 VPWR.n6101 VGND 0.01f
C28307 VPWR.n6102 VGND 0.00524f
C28308 VPWR.t598 VGND 0.00387f
C28309 VPWR.n6103 VGND 0.00837f
C28310 VPWR.n6104 VGND 0.00471f
C28311 VPWR.n6105 VGND 0.00393f
C28312 VPWR.n6106 VGND 0.00199f
C28313 VPWR.n6107 VGND 0.00199f
C28314 VPWR.n6108 VGND 0.00943f
C28315 VPWR.t2900 VGND 0.0299f
C28316 VPWR.t3026 VGND 0.0237f
C28317 VPWR.t563 VGND 0.0163f
C28318 VPWR.t2246 VGND 0.0356f
C28319 VPWR.t3141 VGND 0.0154f
C28320 VPWR.t1348 VGND 0.0109f
C28321 VPWR.t1827 VGND 0.0144f
C28322 VPWR.t1171 VGND 0.0146f
C28323 VPWR.t3109 VGND 0.0213f
C28324 VPWR.t2869 VGND 0.026f
C28325 VPWR.t255 VGND 0.0154f
C28326 VPWR.t3021 VGND 0.0295f
C28327 VPWR.t1173 VGND 0.0232f
C28328 VPWR.t3195 VGND 0.0109f
C28329 VPWR.t2244 VGND 0.0163f
C28330 VPWR.t3115 VGND 0.0148f
C28331 VPWR.t1980 VGND 0.0282f
C28332 VPWR.t1205 VGND 0.0215f
C28333 VPWR.t1174 VGND 0.0211f
C28334 VPWR.t617 VGND 0.0144f
C28335 VPWR.t3020 VGND 0.024f
C28336 VPWR.t1557 VGND 0.0258f
C28337 VPWR.t1377 VGND 0.0112f
C28338 VPWR.t2295 VGND 0.0141f
C28339 VPWR.t3018 VGND 0.0141f
C28340 VPWR.t2293 VGND 0.0258f
C28341 VPWR.t1555 VGND 0.0337f
C28342 VPWR.n6109 VGND 0.0399f
C28343 VPWR.t240 VGND 0.0151f
C28344 VPWR.t3142 VGND 0.0299f
C28345 VPWR.t1346 VGND 0.0284f
C28346 VPWR.t1608 VGND 0.0322f
C28347 VPWR.t3101 VGND 0.0262f
C28348 VPWR.t2501 VGND 0.0294f
C28349 VPWR.t1885 VGND 0.0185f
C28350 VPWR.t877 VGND 0.00587f
C28351 VPWR.t1185 VGND 0.0153f
C28352 VPWR.t237 VGND 0.0109f
C28353 VPWR.t1835 VGND 0.0144f
C28354 VPWR.t3060 VGND 0.0358f
C28355 VPWR.t2242 VGND 0.0112f
C28356 VPWR.t2219 VGND 0.0154f
C28357 VPWR.t793 VGND 0.0141f
C28358 VPWR.t2217 VGND 0.0166f
C28359 VPWR.t3062 VGND 0.021f
C28360 VPWR.t1880 VGND 0.0336f
C28361 VPWR.t2850 VGND 0.0396f
C28362 VPWR.t597 VGND 0.0331f
C28363 VPWR.t2727 VGND 0.0264f
C28364 VPWR.t3063 VGND 0.0311f
C28365 VPWR.t794 VGND 0.0285f
C28366 VPWR.t1357 VGND 0.0262f
C28367 VPWR.t2834 VGND 0.018f
C28368 VPWR.n6110 VGND 0.0176f
C28369 VPWR.t2315 VGND 0.0129f
C28370 VPWR.t1355 VGND 0.0178f
C28371 VPWR.t1884 VGND 0.0196f
C28372 VPWR.t2499 VGND 0.0131f
C28373 VPWR.t2202 VGND 0.0463f
C28374 VPWR.t333 VGND 0.0415f
C28375 VPWR.t303 VGND 0.028f
C28376 VPWR.t2232 VGND 0.0257f
C28377 VPWR.t2972 VGND 0.0354f
C28378 VPWR.t30 VGND 0.0878f
C28379 VPWR.t631 VGND 0.0975f
C28380 VPWR.n6111 VGND 0.0653f
C28381 VPWR.n6112 VGND 0.011f
C28382 VPWR.t212 VGND 0.0046f
C28383 VPWR.n6113 VGND 0.00644f
C28384 VPWR.n6114 VGND 0.00535f
C28385 VPWR.t3388 VGND 0.0612f
C28386 VPWR.n6115 VGND 0.011f
C28387 VPWR.t544 VGND 0.0046f
C28388 VPWR.n6116 VGND 0.00644f
C28389 VPWR.n6117 VGND 0.011f
C28390 VPWR.t530 VGND 0.0046f
C28391 VPWR.n6118 VGND 0.00644f
C28392 VPWR.t529 VGND 0.0046f
C28393 VPWR.n6119 VGND 0.0101f
C28394 VPWR.t543 VGND 0.0046f
C28395 VPWR.n6120 VGND 0.011f
C28396 VPWR.n6121 VGND 0.00644f
C28397 VPWR.n6122 VGND 0.00205f
C28398 VPWR.t3504 VGND 0.0578f
C28399 VPWR.n6123 VGND 0.0317f
C28400 VPWR.n6124 VGND 0.0019f
C28401 VPWR.n6125 VGND 0.0113f
C28402 VPWR.n6126 VGND 0.0118f
C28403 VPWR.t15 VGND 0.053f
C28404 VPWR.t2185 VGND 0.0463f
C28405 VPWR.t0 VGND 0.0144f
C28406 VPWR.t2181 VGND 0.0183f
C28407 VPWR.t2183 VGND 0.0191f
C28408 VPWR.t2179 VGND 0.0305f
C28409 VPWR.t2014 VGND 0.0272f
C28410 VPWR.t3069 VGND 0.0196f
C28411 VPWR.t3071 VGND 0.0302f
C28412 VPWR.t424 VGND 0.0423f
C28413 VPWR.t75 VGND 0.0618f
C28414 VPWR.t660 VGND 0.0975f
C28415 VPWR.t306 VGND 0.0878f
C28416 VPWR.t712 VGND 0.0878f
C28417 VPWR.t210 VGND 0.0975f
C28418 VPWR.t542 VGND 0.0878f
C28419 VPWR.t528 VGND 0.0975f
C28420 VPWR.t309 VGND 0.0618f
C28421 VPWR.n6127 VGND 0.034f
C28422 VPWR.n6128 VGND 0.0145f
C28423 VPWR.t307 VGND 0.0046f
C28424 VPWR.n6129 VGND 0.00126f
C28425 VPWR.n6130 VGND 0.0053f
C28426 VPWR.n6131 VGND 9.6e-19
C28427 VPWR.n6132 VGND 3.73e-19
C28428 VPWR.n6133 VGND 5.27e-19
C28429 VPWR.n6134 VGND 3.95e-19
C28430 VPWR.n6135 VGND 5.05e-19
C28431 VPWR.n6136 VGND 5.05e-19
C28432 VPWR.n6137 VGND 9.06e-19
C28433 VPWR.n6138 VGND 0.0057f
C28434 VPWR.n6139 VGND 6.54e-19
C28435 VPWR.n6140 VGND 8.67e-19
C28436 VPWR.n6141 VGND 4.39e-19
C28437 VPWR.n6142 VGND 3.29e-19
C28438 VPWR.n6143 VGND 5.27e-19
C28439 VPWR.n6144 VGND 2.85e-19
C28440 VPWR.n6145 VGND 2.85e-19
C28441 VPWR.n6146 VGND 4.17e-19
C28442 VPWR.n6147 VGND 5.71e-19
C28443 VPWR.n6148 VGND 4.17e-19
C28444 VPWR.n6149 VGND 3.51e-19
C28445 VPWR.n6150 VGND 4.61e-19
C28446 VPWR.n6151 VGND 4.17e-19
C28447 VPWR.n6152 VGND 4.83e-19
C28448 VPWR.n6153 VGND 4.61e-19
C28449 VPWR.n6154 VGND 3.73e-19
C28450 VPWR.n6155 VGND 2.41e-19
C28451 VPWR.t3530 VGND 0.0289f
C28452 VPWR.t572 VGND 0.00387f
C28453 VPWR.n6156 VGND 0.0547f
C28454 VPWR.t227 VGND 0.00398f
C28455 VPWR.n6157 VGND 0.0317f
C28456 VPWR.t2665 VGND 0.00651f
C28457 VPWR.n6158 VGND 0.0077f
C28458 VPWR.t2663 VGND 0.00634f
C28459 VPWR.t3431 VGND 0.0289f
C28460 VPWR.t226 VGND 0.00387f
C28461 VPWR.n6159 VGND 0.0604f
C28462 VPWR.n6160 VGND 0.0212f
C28463 VPWR.n6161 VGND 0.0117f
C28464 VPWR.t819 VGND 0.0065f
C28465 VPWR.t2045 VGND 0.00682f
C28466 VPWR.t2049 VGND 0.00166f
C28467 VPWR.t2051 VGND 0.00166f
C28468 VPWR.n6162 VGND 0.00341f
C28469 VPWR.n6163 VGND 0.0101f
C28470 VPWR.n6164 VGND 0.00444f
C28471 VPWR.t3542 VGND 0.00911f
C28472 VPWR.t552 VGND 0.00391f
C28473 VPWR.n6165 VGND 0.0253f
C28474 VPWR.t553 VGND 0.00391f
C28475 VPWR.n6167 VGND 0.0138f
C28476 VPWR.t3518 VGND 0.00911f
C28477 VPWR.t521 VGND 0.00391f
C28478 VPWR.n6168 VGND 0.0253f
C28479 VPWR.t520 VGND 0.00391f
C28480 VPWR.n6170 VGND 0.0138f
C28481 VPWR.n6171 VGND 0.00345f
C28482 VPWR.t3455 VGND 0.00911f
C28483 VPWR.t301 VGND 0.00391f
C28484 VPWR.n6172 VGND 0.0253f
C28485 VPWR.t302 VGND 0.00391f
C28486 VPWR.n6174 VGND 0.0138f
C28487 VPWR.n6175 VGND 0.0109f
C28488 VPWR.n6176 VGND 0.00748f
C28489 VPWR.n6177 VGND 0.00696f
C28490 VPWR.n6178 VGND 0.00393f
C28491 VPWR.t2047 VGND 0.00225f
C28492 VPWR.t2287 VGND 0.00166f
C28493 VPWR.n6179 VGND 0.0045f
C28494 VPWR.n6180 VGND 0.00727f
C28495 VPWR.n6181 VGND 0.00524f
C28496 VPWR.t817 VGND 0.00651f
C28497 VPWR.n6182 VGND 0.00774f
C28498 VPWR.n6183 VGND 0.0031f
C28499 VPWR.n6184 VGND 0.00179f
C28500 VPWR.n6185 VGND 0.00392f
C28501 VPWR.n6186 VGND 0.0169f
C28502 VPWR.n6187 VGND 0.00313f
C28503 VPWR.n6188 VGND 0.00618f
C28504 VPWR.n6189 VGND 0.0172f
C28505 VPWR.n6190 VGND 0.0167f
C28506 VPWR.n6191 VGND 0.0107f
C28507 VPWR.t446 VGND 0.0046f
C28508 VPWR.n6192 VGND 0.01f
C28509 VPWR.n6193 VGND 0.0112f
C28510 VPWR.n6194 VGND 0.00393f
C28511 VPWR.n6195 VGND 0.00865f
C28512 VPWR.n6196 VGND 0.00171f
C28513 VPWR.n6197 VGND 0.00925f
C28514 VPWR.n6198 VGND 0.0166f
C28515 VPWR.n6199 VGND 0.0039f
C28516 VPWR.n6200 VGND 9e-19
C28517 VPWR.n6201 VGND 0.00138f
C28518 VPWR.n6202 VGND 9.06e-19
C28519 VPWR.n6203 VGND 5.48e-19
C28520 VPWR.n6204 VGND 6.14e-19
C28521 VPWR.n6205 VGND 0.00138f
C28522 VPWR.n6206 VGND 0.00206f
C28523 VPWR.n6207 VGND 0.00153f
C28524 VPWR.n6208 VGND 4.27e-19
C28525 VPWR.n6209 VGND 1.14e-19
C28526 VPWR.n6210 VGND 4.27e-19
C28527 VPWR.n6211 VGND 6.83e-19
C28528 VPWR.n6212 VGND 3.7e-19
C28529 VPWR.n6213 VGND 9.68e-19
C28530 VPWR.n6214 VGND 9.96e-19
C28531 VPWR.n6215 VGND 5.41e-19
C28532 VPWR.n6216 VGND 7.4e-19
C28533 VPWR.t573 VGND 0.00387f
C28534 VPWR.n6217 VGND 0.0102f
C28535 VPWR.n6218 VGND 0.00171f
C28536 VPWR.n6219 VGND 6.03e-19
C28537 VPWR.n6220 VGND 3.13e-19
C28538 VPWR.n6221 VGND 2.56e-19
C28539 VPWR.n6222 VGND 4.55e-19
C28540 VPWR.n6223 VGND 0.0049f
C28541 VPWR.n6224 VGND 2.56e-19
C28542 VPWR.n6225 VGND 0.0109f
C28543 VPWR.t447 VGND 0.0046f
C28544 VPWR.n6226 VGND 0.00644f
C28545 VPWR.t300 VGND 0.053f
C28546 VPWR.t2044 VGND 0.0463f
C28547 VPWR.t551 VGND 0.0144f
C28548 VPWR.t2048 VGND 0.0183f
C28549 VPWR.t2050 VGND 0.0191f
C28550 VPWR.t2046 VGND 0.0163f
C28551 VPWR.t818 VGND 0.0159f
C28552 VPWR.t816 VGND 0.0143f
C28553 VPWR.t2286 VGND 0.0112f
C28554 VPWR.t2664 VGND 0.0196f
C28555 VPWR.t2662 VGND 0.0564f
C28556 VPWR.t225 VGND 0.0616f
C28557 VPWR.t571 VGND 0.0618f
C28558 VPWR.t445 VGND 0.0975f
C28559 VPWR.t57 VGND 0.0878f
C28560 VPWR.t486 VGND 0.0878f
C28561 VPWR.t703 VGND 0.0975f
C28562 VPWR.t330 VGND 0.0618f
C28563 VPWR.t1817 VGND 0.0257f
C28564 VPWR.t2674 VGND 0.0354f
C28565 VPWR.t285 VGND 0.0183f
C28566 VPWR.t347 VGND 0.0358f
C28567 VPWR.t2824 VGND 0.0253f
C28568 VPWR.t2822 VGND 0.0351f
C28569 VPWR.t160 VGND 0.0492f
C28570 VPWR.n6227 VGND 0.0547f
C28571 VPWR.t59 VGND 0.00462f
C28572 VPWR.n6228 VGND 0.0148f
C28573 VPWR.n6229 VGND 0.00854f
C28574 VPWR.t2823 VGND 0.00631f
C28575 VPWR.n6230 VGND 0.00884f
C28576 VPWR.t2825 VGND 0.00632f
C28577 VPWR.n6231 VGND 0.00937f
C28578 VPWR.t3434 VGND 0.0592f
C28579 VPWR.t287 VGND 0.00462f
C28580 VPWR.n6232 VGND 0.00793f
C28581 VPWR.t3471 VGND 0.0111f
C28582 VPWR.n6233 VGND 0.0205f
C28583 VPWR.n6234 VGND 0.00719f
C28584 VPWR.t332 VGND 0.00387f
C28585 VPWR.n6235 VGND 0.0186f
C28586 VPWR.t331 VGND 0.00387f
C28587 VPWR.n6236 VGND 0.0163f
C28588 VPWR.n6237 VGND 0.00638f
C28589 VPWR.n6238 VGND 0.0132f
C28590 VPWR.n6239 VGND 0.0115f
C28591 VPWR.n6240 VGND 0.0118f
C28592 VPWR.n6241 VGND 0.0031f
C28593 VPWR.n6242 VGND 0.00524f
C28594 VPWR.n6243 VGND 0.0113f
C28595 VPWR.n6244 VGND 0.00524f
C28596 VPWR.t3524 VGND 0.0592f
C28597 VPWR.n6245 VGND 0.038f
C28598 VPWR.n6246 VGND 0.00833f
C28599 VPWR.n6247 VGND 0.00524f
C28600 VPWR.n6248 VGND 0.0087f
C28601 VPWR.n6249 VGND 0.00524f
C28602 VPWR.n6250 VGND 0.0113f
C28603 VPWR.n6251 VGND 0.00524f
C28604 VPWR.n6252 VGND 0.011f
C28605 VPWR.n6253 VGND 0.00524f
C28606 VPWR.t704 VGND 0.00461f
C28607 VPWR.t3578 VGND 0.0578f
C28608 VPWR.n6254 VGND 0.0317f
C28609 VPWR.n6255 VGND 0.0101f
C28610 VPWR.n6256 VGND 0.0113f
C28611 VPWR.n6257 VGND 0.00247f
C28612 VPWR.t487 VGND 0.0046f
C28613 VPWR.n6258 VGND 0.00644f
C28614 VPWR.n6259 VGND 0.00148f
C28615 VPWR.n6260 VGND 0.00393f
C28616 VPWR.n6261 VGND 0.00723f
C28617 VPWR.n6262 VGND 0.00279f
C28618 VPWR.n6263 VGND 0.00529f
C28619 VPWR.n6264 VGND 0.0103f
C28620 VPWR.n6265 VGND 0.00556f
C28621 VPWR.n6266 VGND 0.0031f
C28622 VPWR.t2675 VGND 0.00136f
C28623 VPWR.t1818 VGND 0.00136f
C28624 VPWR.n6267 VGND 0.00317f
C28625 VPWR.n6268 VGND 0.0121f
C28626 VPWR.n6269 VGND 0.00524f
C28627 VPWR.n6270 VGND 0.00393f
C28628 VPWR.n6271 VGND 0.0066f
C28629 VPWR.n6272 VGND 0.0066f
C28630 VPWR.n6273 VGND 0.0031f
C28631 VPWR.t3483 VGND 0.00911f
C28632 VPWR.t348 VGND 0.00391f
C28633 VPWR.n6274 VGND 0.0253f
C28634 VPWR.t349 VGND 0.00391f
C28635 VPWR.n6276 VGND 0.0126f
C28636 VPWR.n6277 VGND 0.0108f
C28637 VPWR.n6278 VGND 0.00524f
C28638 VPWR.n6279 VGND 0.00393f
C28639 VPWR.n6280 VGND 0.00484f
C28640 VPWR.n6281 VGND 0.0356f
C28641 VPWR.n6282 VGND 0.00183f
C28642 VPWR.n6283 VGND 0.0031f
C28643 VPWR.n6284 VGND 0.00639f
C28644 VPWR.n6285 VGND 0.00524f
C28645 VPWR.n6286 VGND 0.00393f
C28646 VPWR.n6287 VGND 0.0024f
C28647 VPWR.t286 VGND 0.00463f
C28648 VPWR.n6288 VGND 0.00578f
C28649 VPWR.n6289 VGND 0.00859f
C28650 VPWR.t3403 VGND 0.0182f
C28651 VPWR.t161 VGND 0.00387f
C28652 VPWR.n6290 VGND 0.0244f
C28653 VPWR.n6291 VGND 0.0153f
C28654 VPWR.t162 VGND 0.004f
C28655 VPWR.n6292 VGND 0.00482f
C28656 VPWR.n6293 VGND 0.00249f
C28657 VPWR.n6294 VGND 0.00262f
C28658 VPWR.n6295 VGND 0.00442f
C28659 VPWR.n6296 VGND 0.00282f
C28660 VPWR.n6297 VGND 0.0134f
C28661 VPWR.n6298 VGND 0.00535f
C28662 VPWR.n6299 VGND 0.0031f
C28663 VPWR.n6300 VGND 0.011f
C28664 VPWR.n6301 VGND 0.00524f
C28665 VPWR.n6302 VGND 0.0113f
C28666 VPWR.n6303 VGND 0.00524f
C28667 VPWR.t3354 VGND 0.0592f
C28668 VPWR.n6304 VGND 0.038f
C28669 VPWR.n6305 VGND 0.00833f
C28670 VPWR.n6306 VGND 0.00524f
C28671 VPWR.n6307 VGND 0.0087f
C28672 VPWR.n6308 VGND 0.00524f
C28673 VPWR.n6309 VGND 0.0113f
C28674 VPWR.n6310 VGND 0.00524f
C28675 VPWR.n6311 VGND 0.00451f
C28676 VPWR.n6312 VGND 5.27e-19
C28677 VPWR.n6313 VGND 3.95e-19
C28678 VPWR.n6314 VGND 5.05e-19
C28679 VPWR.n6315 VGND 5.05e-19
C28680 VPWR.n6316 VGND 8.67e-19
C28681 VPWR.n6317 VGND 6.54e-19
C28682 VPWR.n6318 VGND 9.06e-19
C28683 VPWR.n6319 VGND 0.0057f
C28684 VPWR.n6320 VGND 6.54e-19
C28685 VPWR.n6321 VGND 8.67e-19
C28686 VPWR.n6322 VGND 4.39e-19
C28687 VPWR.n6323 VGND 3.29e-19
C28688 VPWR.n6324 VGND 5.27e-19
C28689 VPWR.n6325 VGND 2.85e-19
C28690 VPWR.n6326 VGND 2.85e-19
C28691 VPWR.n6327 VGND 4.17e-19
C28692 VPWR.n6328 VGND 5.41e-19
C28693 VPWR.n6329 VGND 3.42e-19
C28694 VPWR.n6330 VGND 5.27e-19
C28695 VPWR.n6331 VGND 3.95e-19
C28696 VPWR.n6332 VGND 5.05e-19
C28697 VPWR.n6333 VGND 5.05e-19
C28698 VPWR.n6334 VGND 8.67e-19
C28699 VPWR.n6335 VGND 6.54e-19
C28700 VPWR.n6336 VGND 9.06e-19
C28701 VPWR.n6337 VGND 0.0323f
C28702 VPWR.n6339 VGND 0.00139f
C28703 VPWR.n6340 VGND 5.48e-19
C28704 VPWR.n6341 VGND 3.07e-19
C28705 VPWR.n6342 VGND 5.98e-19
C28706 VPWR.t1503 VGND 8.82e-19
C28707 VPWR.t1289 VGND 0.00144f
C28708 VPWR.n6343 VGND 0.00521f
C28709 VPWR.n6344 VGND 0.00571f
C28710 VPWR.t2198 VGND 0.00638f
C28711 VPWR.n6345 VGND 0.00967f
C28712 VPWR.n6346 VGND 2.52e-19
C28713 VPWR.t1291 VGND 0.00148f
C28714 VPWR.t1692 VGND 9.71e-19
C28715 VPWR.n6347 VGND 0.00364f
C28716 VPWR.n6348 VGND 0.00728f
C28717 VPWR.n6349 VGND 9.78e-19
C28718 VPWR.n6350 VGND 0.00199f
C28719 VPWR.t86 VGND 0.053f
C28720 VPWR.t2713 VGND 0.054f
C28721 VPWR.t276 VGND 0.0144f
C28722 VPWR.t2715 VGND 0.0153f
C28723 VPWR.t2709 VGND 0.0252f
C28724 VPWR.t2711 VGND 0.0154f
C28725 VPWR.t745 VGND 0.0112f
C28726 VPWR.t2418 VGND 0.0111f
C28727 VPWR.t2199 VGND 0.028f
C28728 VPWR.t267 VGND 0.0364f
C28729 VPWR.t812 VGND 0.0205f
C28730 VPWR.t2991 VGND 0.0253f
C28731 VPWR.t2593 VGND 0.0143f
C28732 VPWR.t2041 VGND 0.0163f
C28733 VPWR.t2416 VGND 0.025f
C28734 VPWR.t2201 VGND 0.0186f
C28735 VPWR.t3249 VGND 0.0178f
C28736 VPWR.t3145 VGND 0.0203f
C28737 VPWR.t1329 VGND 0.0257f
C28738 VPWR.t706 VGND 0.0309f
C28739 VPWR.t1502 VGND 0.0181f
C28740 VPWR.t1288 VGND 0.0185f
C28741 VPWR.t2197 VGND 0.0146f
C28742 VPWR.t2094 VGND 0.029f
C28743 VPWR.t1290 VGND 0.0208f
C28744 VPWR.t1656 VGND 0.0161f
C28745 VPWR.t1691 VGND 0.0129f
C28746 VPWR.t2999 VGND 0.0307f
C28747 VPWR.t784 VGND 0.0309f
C28748 VPWR.t1856 VGND 0.0116f
C28749 VPWR.t1239 VGND 0.0126f
C28750 VPWR.n6351 VGND 0.0066f
C28751 VPWR.t3350 VGND 0.0592f
C28752 VPWR.t1444 VGND 0.00136f
C28753 VPWR.t1644 VGND 0.00136f
C28754 VPWR.n6352 VGND 0.00317f
C28755 VPWR.t392 VGND 0.0046f
C28756 VPWR.n6353 VGND 0.00407f
C28757 VPWR.t2994 VGND 0.00131f
C28758 VPWR.t2037 VGND 4.27e-19
C28759 VPWR.n6354 VGND 0.00672f
C28760 VPWR.n6355 VGND 0.00674f
C28761 VPWR.t135 VGND 0.0046f
C28762 VPWR.n6356 VGND 0.004f
C28763 VPWR.t50 VGND 0.00387f
C28764 VPWR.n6357 VGND 0.00837f
C28765 VPWR.t1702 VGND 9.71e-19
C28766 VPWR.t3138 VGND 9.22e-19
C28767 VPWR.n6358 VGND 0.00197f
C28768 VPWR.t1202 VGND 6.73e-19
C28769 VPWR.t1200 VGND 6.73e-19
C28770 VPWR.n6359 VGND 0.00142f
C28771 VPWR.n6360 VGND 0.00777f
C28772 VPWR.t3493 VGND 0.0289f
C28773 VPWR.t49 VGND 0.00387f
C28774 VPWR.n6361 VGND 0.0604f
C28775 VPWR.n6362 VGND 0.0146f
C28776 VPWR.n6363 VGND 0.0117f
C28777 VPWR.n6364 VGND 0.0104f
C28778 VPWR.n6365 VGND 0.00199f
C28779 VPWR.n6366 VGND 0.00899f
C28780 VPWR.n6367 VGND 0.0113f
C28781 VPWR.n6368 VGND 0.0104f
C28782 VPWR.n6369 VGND 0.0136f
C28783 VPWR.n6370 VGND 0.00524f
C28784 VPWR.t2730 VGND 0.00469f
C28785 VPWR.n6371 VGND 0.0113f
C28786 VPWR.n6372 VGND 0.00658f
C28787 VPWR.n6373 VGND 0.00524f
C28788 VPWR.n6374 VGND 0.0031f
C28789 VPWR.n6375 VGND 0.00483f
C28790 VPWR.n6376 VGND 0.00169f
C28791 VPWR.t2936 VGND 0.00102f
C28792 VPWR.t1919 VGND 0.00102f
C28793 VPWR.n6377 VGND 0.00208f
C28794 VPWR.n6378 VGND 0.00292f
C28795 VPWR.t134 VGND 0.0046f
C28796 VPWR.n6379 VGND 0.00392f
C28797 VPWR.n6380 VGND 0.00115f
C28798 VPWR.n6381 VGND 0.00115f
C28799 VPWR.n6382 VGND 0.00393f
C28800 VPWR.n6383 VGND 0.0031f
C28801 VPWR.n6384 VGND 0.00639f
C28802 VPWR.n6385 VGND 0.0066f
C28803 VPWR.n6386 VGND 0.00199f
C28804 VPWR.n6387 VGND 0.00506f
C28805 VPWR.n6388 VGND 0.00393f
C28806 VPWR.t3516 VGND 0.0592f
C28807 VPWR.n6389 VGND 0.0356f
C28808 VPWR.n6390 VGND 0.00319f
C28809 VPWR.n6391 VGND 0.00524f
C28810 VPWR.t2988 VGND 7.22e-19
C28811 VPWR.t1824 VGND 9.22e-19
C28812 VPWR.n6392 VGND 0.00189f
C28813 VPWR.n6393 VGND 0.00612f
C28814 VPWR.n6394 VGND 0.00495f
C28815 VPWR.n6395 VGND 0.00524f
C28816 VPWR.n6396 VGND 0.0066f
C28817 VPWR.n6397 VGND 0.00524f
C28818 VPWR.n6398 VGND 0.0066f
C28819 VPWR.n6399 VGND 0.00524f
C28820 VPWR.n6400 VGND 0.0066f
C28821 VPWR.n6401 VGND 0.00524f
C28822 VPWR.n6402 VGND 0.0066f
C28823 VPWR.n6403 VGND 0.00524f
C28824 VPWR.n6404 VGND 0.00337f
C28825 VPWR.n6405 VGND 0.00524f
C28826 VPWR.n6406 VGND 0.00307f
C28827 VPWR.n6407 VGND 0.00264f
C28828 VPWR.n6408 VGND 0.00259f
C28829 VPWR.n6409 VGND 0.00199f
C28830 VPWR.n6410 VGND 0.00179f
C28831 VPWR.n6411 VGND 0.00639f
C28832 VPWR.n6412 VGND 0.0121f
C28833 VPWR.n6413 VGND 0.00475f
C28834 VPWR.n6414 VGND 0.00393f
C28835 VPWR.n6415 VGND 0.00506f
C28836 VPWR.n6416 VGND 0.0356f
C28837 VPWR.n6417 VGND 0.00484f
C28838 VPWR.n6418 VGND 0.00393f
C28839 VPWR.n6419 VGND 0.00333f
C28840 VPWR.n6420 VGND 0.00199f
C28841 VPWR.t437 VGND 0.00387f
C28842 VPWR.n6421 VGND 0.0107f
C28843 VPWR.n6422 VGND 0.00796f
C28844 VPWR.n6423 VGND 0.00122f
C28845 VPWR.n6424 VGND 8.11e-19
C28846 VPWR.n6425 VGND 3.95e-19
C28847 VPWR.n6426 VGND 3.95e-19
C28848 VPWR.n6427 VGND 7.68e-19
C28849 VPWR.n6428 VGND 5.05e-19
C28850 VPWR.n6429 VGND 0.00139f
C28851 VPWR.n6430 VGND 9.06e-19
C28852 VPWR.n6431 VGND 5.48e-19
C28853 VPWR.n6432 VGND 1.76e-19
C28854 VPWR.n6433 VGND 1.76e-19
C28855 VPWR.n6434 VGND 3.13e-19
C28856 VPWR.n6435 VGND 5.12e-19
C28857 VPWR.n6436 VGND 6.26e-19
C28858 VPWR.n6437 VGND 2.28e-19
C28859 VPWR.n6438 VGND 2.85e-19
C28860 VPWR.n6439 VGND 0.00259f
C28861 VPWR.t3492 VGND 0.0231f
C28862 VPWR.n6440 VGND 0.00925f
C28863 VPWR.n6441 VGND 0.0419f
C28864 VPWR.n6442 VGND 0.00495f
C28865 VPWR.n6443 VGND 0.00393f
C28866 VPWR.n6444 VGND 0.00199f
C28867 VPWR.n6445 VGND 0.00629f
C28868 VPWR.n6446 VGND 0.0147f
C28869 VPWR.t2779 VGND 0.0154f
C28870 VPWR.t2800 VGND 0.0413f
C28871 VPWR.t2000 VGND 0.0183f
C28872 VPWR.t139 VGND 0.0153f
C28873 VPWR.t3042 VGND 0.0358f
C28874 VPWR.t2250 VGND 0.0408f
C28875 VPWR.t2248 VGND 0.0196f
C28876 VPWR.t634 VGND 0.0154f
C28877 VPWR.t693 VGND 0.0618f
C28878 VPWR.t231 VGND 0.026f
C28879 VPWR.t1546 VGND 0.0222f
C28880 VPWR.t1544 VGND 0.0201f
C28881 VPWR.t3054 VGND 0.0107f
C28882 VPWR.t2001 VGND 0.00537f
C28883 VPWR.t3086 VGND 0.0154f
C28884 VPWR.t2385 VGND 0.0309f
C28885 VPWR.t436 VGND 0.0621f
C28886 VPWR.n6447 VGND 0.0292f
C28887 VPWR.t391 VGND 0.0124f
C28888 VPWR.t1643 VGND 0.0567f
C28889 VPWR.t1443 VGND 0.02f
C28890 VPWR.t2036 VGND 0.0217f
C28891 VPWR.t2993 VGND 0.0356f
C28892 VPWR.t2093 VGND 0.0532f
C28893 VPWR.t1654 VGND 0.0413f
C28894 VPWR.t133 VGND 0.0121f
C28895 VPWR.t1823 VGND 0.0228f
C28896 VPWR.t2987 VGND 0.0448f
C28897 VPWR.t1918 VGND 0.0222f
C28898 VPWR.t2935 VGND 0.02f
C28899 VPWR.t2729 VGND 0.042f
C28900 VPWR.t1238 VGND 0.0304f
C28901 VPWR.t2937 VGND 0.0149f
C28902 VPWR.t48 VGND 0.0201f
C28903 VPWR.t3137 VGND 0.0371f
C28904 VPWR.t1701 VGND 0.0319f
C28905 VPWR.t1199 VGND 0.0282f
C28906 VPWR.t1201 VGND 0.0158f
C28907 VPWR.t2934 VGND 0.018f
C28908 VPWR.n6448 VGND 0.0219f
C28909 VPWR.n6449 VGND 0.0102f
C28910 VPWR.n6450 VGND 0.00102f
C28911 VPWR.n6451 VGND 0.00484f
C28912 VPWR.t1857 VGND 0.00233f
C28913 VPWR.t785 VGND 0.00569f
C28914 VPWR.t3000 VGND 0.00557f
C28915 VPWR.n6452 VGND 0.00785f
C28916 VPWR.n6453 VGND 0.0212f
C28917 VPWR.n6454 VGND 0.00699f
C28918 VPWR.n6455 VGND 0.00698f
C28919 VPWR.n6456 VGND 0.00139f
C28920 VPWR.n6457 VGND 0.00524f
C28921 VPWR.n6458 VGND 0.00182f
C28922 VPWR.n6459 VGND 0.00524f
C28923 VPWR.n6460 VGND 0.00387f
C28924 VPWR.n6461 VGND 0.00131f
C28925 VPWR.n6462 VGND 9.42e-19
C28926 VPWR.n6463 VGND 2.63e-19
C28927 VPWR.n6464 VGND 1.76e-19
C28928 VPWR.n6465 VGND 2.28e-19
C28929 VPWR.n6466 VGND 0.00402f
C28930 VPWR.n6467 VGND 4.84e-19
C28931 VPWR.n6468 VGND 0.00105f
C28932 VPWR.n6469 VGND 4.27e-19
C28933 VPWR.t708 VGND 0.00387f
C28934 VPWR.n6470 VGND 0.00202f
C28935 VPWR.n6471 VGND 6.73e-19
C28936 VPWR.n6472 VGND 4.27e-19
C28937 VPWR.n6473 VGND 0.00516f
C28938 VPWR.n6474 VGND 4.84e-19
C28939 VPWR.n6475 VGND 6.83e-19
C28940 VPWR.n6476 VGND 4.84e-19
C28941 VPWR.n6477 VGND 3.13e-19
C28942 VPWR.n6478 VGND 9.96e-19
C28943 VPWR.n6479 VGND 0.00575f
C28944 VPWR.n6480 VGND 9.68e-19
C28945 VPWR.n6481 VGND 4.55e-19
C28946 VPWR.n6482 VGND 2.56e-19
C28947 VPWR.n6483 VGND 0.00127f
C28948 VPWR.n6484 VGND 0.00152f
C28949 VPWR.t3428 VGND 0.00911f
C28950 VPWR.t269 VGND 0.00391f
C28951 VPWR.n6485 VGND 0.0253f
C28952 VPWR.t268 VGND 0.00391f
C28953 VPWR.n6487 VGND 0.0138f
C28954 VPWR.t2706 VGND 5.02e-19
C28955 VPWR.t2200 VGND 0.00135f
C28956 VPWR.n6488 VGND 0.00626f
C28957 VPWR.n6489 VGND 0.0146f
C28958 VPWR.t2419 VGND 0.00261f
C28959 VPWR.t2712 VGND 0.00225f
C28960 VPWR.t746 VGND 0.00166f
C28961 VPWR.n6490 VGND 0.00438f
C28962 VPWR.n6491 VGND 0.00623f
C28963 VPWR.t3366 VGND 0.00911f
C28964 VPWR.t88 VGND 0.00391f
C28965 VPWR.n6492 VGND 0.0253f
C28966 VPWR.t87 VGND 0.00391f
C28967 VPWR.n6494 VGND 0.0138f
C28968 VPWR.n6495 VGND 0.00345f
C28969 VPWR.t3419 VGND 0.00911f
C28970 VPWR.t615 VGND 0.00391f
C28971 VPWR.n6496 VGND 0.0253f
C28972 VPWR.t616 VGND 0.00391f
C28973 VPWR.n6498 VGND 0.0138f
C28974 VPWR.n6499 VGND 0.0112f
C28975 VPWR.t277 VGND 0.00387f
C28976 VPWR.t2714 VGND 0.00682f
C28977 VPWR.n6500 VGND 0.00917f
C28978 VPWR.n6501 VGND 0.00232f
C28979 VPWR.n6502 VGND 0.00487f
C28980 VPWR.n6503 VGND 0.00393f
C28981 VPWR.n6504 VGND 0.00524f
C28982 VPWR.n6505 VGND 0.00524f
C28983 VPWR.t2716 VGND 0.00166f
C28984 VPWR.t2710 VGND 0.00166f
C28985 VPWR.n6506 VGND 0.00341f
C28986 VPWR.t3570 VGND 0.0179f
C28987 VPWR.n6507 VGND 0.017f
C28988 VPWR.n6508 VGND 0.0103f
C28989 VPWR.n6509 VGND 0.00702f
C28990 VPWR.n6510 VGND 0.00912f
C28991 VPWR.t278 VGND 0.00387f
C28992 VPWR.n6511 VGND 0.00822f
C28993 VPWR.n6512 VGND 0.00518f
C28994 VPWR.n6513 VGND 0.0031f
C28995 VPWR.n6514 VGND 0.00179f
C28996 VPWR.n6515 VGND 4.54e-19
C28997 VPWR.n6516 VGND 0.00556f
C28998 VPWR.n6517 VGND 0.00117f
C28999 VPWR.n6518 VGND 0.00262f
C29000 VPWR.n6519 VGND 0.00444f
C29001 VPWR.n6520 VGND 0.00199f
C29002 VPWR.n6521 VGND 0.00125f
C29003 VPWR.t813 VGND 0.00166f
C29004 VPWR.t2992 VGND 0.00166f
C29005 VPWR.n6522 VGND 0.00381f
C29006 VPWR.n6523 VGND 0.00759f
C29007 VPWR.n6524 VGND 0.00393f
C29008 VPWR.n6525 VGND 8.47e-19
C29009 VPWR.n6526 VGND 0.00524f
C29010 VPWR.t2417 VGND 0.00102f
C29011 VPWR.t2594 VGND 0.00154f
C29012 VPWR.n6527 VGND 0.00495f
C29013 VPWR.n6528 VGND 0.00783f
C29014 VPWR.n6529 VGND 0.00524f
C29015 VPWR.t3250 VGND 0.00598f
C29016 VPWR.n6530 VGND 0.00861f
C29017 VPWR.n6531 VGND 0.00524f
C29018 VPWR.n6532 VGND 0.0031f
C29019 VPWR.n6533 VGND 0.00199f
C29020 VPWR.n6534 VGND 0.00152f
C29021 VPWR.n6535 VGND 0.00292f
C29022 VPWR.t3146 VGND 0.00136f
C29023 VPWR.t1330 VGND 0.00136f
C29024 VPWR.n6536 VGND 0.00279f
C29025 VPWR.n6537 VGND 0.00448f
C29026 VPWR.t707 VGND 0.00387f
C29027 VPWR.t3457 VGND 0.0179f
C29028 VPWR.n6538 VGND 0.00344f
C29029 VPWR.n6539 VGND 0.0164f
C29030 VPWR.n6540 VGND 0.00478f
C29031 VPWR.n6541 VGND 0.00177f
C29032 VPWR.n6542 VGND 0.00232f
C29033 VPWR.n6543 VGND 0.00259f
C29034 VPWR.n6544 VGND 9e-19
C29035 VPWR.n6545 VGND 0.00138f
C29036 VPWR.n6546 VGND 9.06e-19
C29037 VPWR.n6547 VGND 5.48e-19
C29038 VPWR.n6548 VGND 6.14e-19
C29039 VPWR.n6549 VGND 0.00138f
C29040 VPWR.n6550 VGND 0.00206f
C29041 VPWR.n6551 VGND 0.00153f
C29042 VPWR.n6552 VGND 4.27e-19
C29043 VPWR.n6553 VGND 1.14e-19
C29044 VPWR.n6554 VGND 5.41e-19
C29045 VPWR.n6555 VGND 5.12e-19
C29046 VPWR.n6556 VGND 3.7e-19
C29047 VPWR.n6557 VGND 6.83e-19
C29048 VPWR.n6558 VGND 4.27e-19
C29049 VPWR.n6559 VGND 0.00127f
C29050 VPWR.n6560 VGND 0.00127f
C29051 VPWR.n6561 VGND 0.0056f
C29052 VPWR.n6562 VGND 3.13e-19
C29053 VPWR.n6563 VGND 7.4e-19
C29054 VPWR.n6564 VGND 5.71e-19
C29055 VPWR.n6565 VGND 4.17e-19
C29056 VPWR.n6566 VGND 3.51e-19
C29057 VPWR.n6567 VGND 4.61e-19
C29058 VPWR.n6568 VGND 4.17e-19
C29059 VPWR.n6569 VGND 4.83e-19
C29060 VPWR.n6570 VGND 4.61e-19
C29061 VPWR.n6571 VGND 3.73e-19
C29062 VPWR.n6572 VGND 2.41e-19
C29063 VPWR.n6573 VGND 4.83e-19
C29064 VPWR.n6574 VGND 4.61e-19
C29065 VPWR.n6575 VGND 4.11e-19
C29066 VPWR.n6576 VGND 4.11e-19
C29067 VPWR.n6577 VGND 7.39e-19
C29068 VPWR.n6578 VGND 5.19e-19
C29069 VPWR.n6579 VGND 7.39e-19
C29070 VPWR.n6580 VGND 4.11e-19
C29071 VPWR.n6581 VGND 4.11e-19
C29072 VPWR.n6583 VGND 0.1f
C29073 VPWR.n6584 VGND 0.1f
C29074 VPWR.n6586 VGND 0.0066f
C29075 VPWR.n6587 VGND 0.00175f
C29076 VPWR.t3328 VGND 0.00695f
C29077 VPWR.n6588 VGND 0.00819f
C29078 VPWR.t3444 VGND 0.00911f
C29079 VPWR.t79 VGND 0.00391f
C29080 VPWR.n6589 VGND 0.0253f
C29081 VPWR.t78 VGND 0.00391f
C29082 VPWR.n6591 VGND 0.0138f
C29083 VPWR.t3559 VGND 0.00911f
C29084 VPWR.t73 VGND 0.00391f
C29085 VPWR.n6592 VGND 0.0253f
C29086 VPWR.t74 VGND 0.00391f
C29087 VPWR.n6594 VGND 0.0138f
C29088 VPWR.n6595 VGND 0.011f
C29089 VPWR.n6596 VGND 0.00345f
C29090 VPWR.n6597 VGND 0.00199f
C29091 VPWR.n6598 VGND 0.00179f
C29092 VPWR.n6599 VGND 0.00111f
C29093 VPWR.t3322 VGND 0.00166f
C29094 VPWR.t3324 VGND 0.00166f
C29095 VPWR.n6600 VGND 0.00344f
C29096 VPWR.t2043 VGND 6.73e-19
C29097 VPWR.t1782 VGND 0.00102f
C29098 VPWR.n6601 VGND 0.00183f
C29099 VPWR.n6602 VGND 0.00857f
C29100 VPWR.n6603 VGND 0.00475f
C29101 VPWR.n6604 VGND 0.00148f
C29102 VPWR.n6605 VGND 0.00524f
C29103 VPWR.t3326 VGND 0.00225f
C29104 VPWR.t2372 VGND 0.00166f
C29105 VPWR.n6606 VGND 0.00438f
C29106 VPWR.n6607 VGND 0.00635f
C29107 VPWR.n6608 VGND 5.04e-19
C29108 VPWR.n6609 VGND 0.00524f
C29109 VPWR.t811 VGND 0.00204f
C29110 VPWR.t2939 VGND 0.0055f
C29111 VPWR.n6610 VGND 0.00336f
C29112 VPWR.n6611 VGND 0.00848f
C29113 VPWR.n6612 VGND 0.00141f
C29114 VPWR.n6613 VGND 0.0031f
C29115 VPWR.n6614 VGND 0.00199f
C29116 VPWR.n6615 VGND 0.00179f
C29117 VPWR.n6616 VGND 0.00269f
C29118 VPWR.t601 VGND 0.0046f
C29119 VPWR.n6617 VGND 0.00407f
C29120 VPWR.n6618 VGND 0.00632f
C29121 VPWR.n6619 VGND 0.00475f
C29122 VPWR.t2990 VGND 0.0016f
C29123 VPWR.t2996 VGND 0.0016f
C29124 VPWR.n6620 VGND 0.00369f
C29125 VPWR.n6621 VGND 0.00624f
C29126 VPWR.n6622 VGND 0.00337f
C29127 VPWR.n6623 VGND 0.00524f
C29128 VPWR.n6624 VGND 0.00506f
C29129 VPWR.n6625 VGND 0.00524f
C29130 VPWR.t3148 VGND 0.00533f
C29131 VPWR.t3459 VGND 0.0592f
C29132 VPWR.n6626 VGND 0.035f
C29133 VPWR.n6627 VGND 0.00444f
C29134 VPWR.n6628 VGND 0.00395f
C29135 VPWR.n6629 VGND 0.00524f
C29136 VPWR.n6630 VGND 0.0066f
C29137 VPWR.n6631 VGND 0.00524f
C29138 VPWR.n6632 VGND 0.00393f
C29139 VPWR.n6633 VGND 0.00199f
C29140 VPWR.n6634 VGND 0.00641f
C29141 VPWR.t675 VGND 0.0046f
C29142 VPWR.n6635 VGND 0.00644f
C29143 VPWR.n6636 VGND 0.0053f
C29144 VPWR.n6637 VGND 0.00393f
C29145 VPWR.n6638 VGND 0.0102f
C29146 VPWR.n6639 VGND 0.0039f
C29147 VPWR.n6640 VGND 0.0109f
C29148 VPWR.t676 VGND 0.0046f
C29149 VPWR.n6641 VGND 0.00644f
C29150 VPWR.t72 VGND 0.046f
C29151 VPWR.t3327 VGND 0.0158f
C29152 VPWR.t2042 VGND 0.00571f
C29153 VPWR.t3321 VGND 0.0149f
C29154 VPWR.t3323 VGND 0.0159f
C29155 VPWR.t1781 VGND 0.0144f
C29156 VPWR.t3325 VGND 0.0148f
C29157 VPWR.t810 VGND 0.0161f
C29158 VPWR.t2371 VGND 0.0253f
C29159 VPWR.t2938 VGND 0.0151f
C29160 VPWR.t3149 VGND 0.0206f
C29161 VPWR.t2989 VGND 0.0282f
C29162 VPWR.t2995 VGND 0.0282f
C29163 VPWR.t3147 VGND 0.0457f
C29164 VPWR.t1302 VGND 0.0332f
C29165 VPWR.t600 VGND 0.0274f
C29166 VPWR.t674 VGND 0.0975f
C29167 VPWR.t107 VGND 0.0878f
C29168 VPWR.n6642 VGND 0.034f
C29169 VPWR.n6643 VGND 0.00556f
C29170 VPWR.t109 VGND 0.00462f
C29171 VPWR.n6644 VGND 0.0103f
C29172 VPWR.n6645 VGND 0.00529f
C29173 VPWR.t1465 VGND 0.00148f
C29174 VPWR.t1704 VGND 9.71e-19
C29175 VPWR.n6646 VGND 0.00358f
C29176 VPWR.n6647 VGND 0.00829f
C29177 VPWR.t375 VGND 0.0046f
C29178 VPWR.n6648 VGND 0.00123f
C29179 VPWR.t440 VGND 0.0046f
C29180 VPWR.n6649 VGND 0.00407f
C29181 VPWR.t1521 VGND 0.00461f
C29182 VPWR.n6650 VGND 0.00352f
C29183 VPWR.t441 VGND 0.0046f
C29184 VPWR.n6651 VGND 0.00396f
C29185 VPWR.n6652 VGND 0.00116f
C29186 VPWR.t3515 VGND 0.00911f
C29187 VPWR.t132 VGND 0.00391f
C29188 VPWR.n6653 VGND 0.0253f
C29189 VPWR.t131 VGND 0.00391f
C29190 VPWR.n6655 VGND 0.0138f
C29191 VPWR.t3080 VGND 0.00102f
C29192 VPWR.t1915 VGND 0.00102f
C29193 VPWR.n6656 VGND 0.00218f
C29194 VPWR.n6657 VGND 0.0124f
C29195 VPWR.t261 VGND 0.0926f
C29196 VPWR.t373 VGND 0.0331f
C29197 VPWR.t1282 VGND 0.0441f
C29198 VPWR.t1466 VGND 0.0475f
C29199 VPWR.t1464 VGND 0.0436f
C29200 VPWR.t1703 VGND 0.0356f
C29201 VPWR.t3133 VGND 0.0436f
C29202 VPWR.t1843 VGND 0.0302f
C29203 VPWR.t3081 VGND 0.0309f
C29204 VPWR.t893 VGND 0.0269f
C29205 VPWR.t891 VGND 0.019f
C29206 VPWR.t439 VGND 0.0141f
C29207 VPWR.t1707 VGND 0.027f
C29208 VPWR.t865 VGND 0.0379f
C29209 VPWR.t3082 VGND 0.0342f
C29210 VPWR.t1844 VGND 0.0304f
C29211 VPWR.t1520 VGND 0.0265f
C29212 VPWR.t2848 VGND 0.0126f
C29213 VPWR.t1721 VGND 0.0183f
C29214 VPWR.t522 VGND 0.0361f
C29215 VPWR.t2552 VGND 0.028f
C29216 VPWR.t1916 VGND 0.0154f
C29217 VPWR.t1960 VGND 0.0415f
C29218 VPWR.t193 VGND 0.0448f
C29219 VPWR.t1614 VGND 0.0284f
C29220 VPWR.t3308 VGND 0.0321f
C29221 VPWR.t1962 VGND 0.0232f
C29222 VPWR.t2702 VGND 0.0178f
C29223 VPWR.t900 VGND 0.0163f
C29224 VPWR.t1687 VGND 0.0121f
C29225 VPWR.t2680 VGND 0.028f
C29226 VPWR.t2717 VGND 0.0213f
C29227 VPWR.t1819 VGND 0.0217f
C29228 VPWR.t1963 VGND 0.026f
C29229 VPWR.t3309 VGND 0.0191f
C29230 VPWR.t1669 VGND 0.0322f
C29231 VPWR.t1689 VGND 0.0322f
C29232 VPWR.t1524 VGND 0.0196f
C29233 VPWR.t113 VGND 0.0361f
C29234 VPWR.t1671 VGND 0.0446f
C29235 VPWR.t1667 VGND 0.0361f
C29236 VPWR.t1914 VGND 0.0222f
C29237 VPWR.t3079 VGND 0.0228f
C29238 VPWR.n6658 VGND 0.0251f
C29239 VPWR.n6659 VGND 5.69e-19
C29240 VPWR.n6660 VGND 0.00131f
C29241 VPWR.n6661 VGND 9.96e-19
C29242 VPWR.n6662 VGND 4.27e-19
C29243 VPWR.n6663 VGND 5.12e-19
C29244 VPWR.n6664 VGND 5.41e-19
C29245 VPWR.n6665 VGND 7.35e-19
C29246 VPWR.t3534 VGND 0.0289f
C29247 VPWR.t114 VGND 0.00387f
C29248 VPWR.n6666 VGND 0.0604f
C29249 VPWR.n6667 VGND 0.0116f
C29250 VPWR.n6668 VGND 0.0117f
C29251 VPWR.t1668 VGND 0.00632f
C29252 VPWR.t1672 VGND 0.00676f
C29253 VPWR.t1525 VGND 0.00234f
C29254 VPWR.n6669 VGND 0.00258f
C29255 VPWR.n6670 VGND 0.0173f
C29256 VPWR.n6671 VGND 0.00966f
C29257 VPWR.n6672 VGND 2.95e-19
C29258 VPWR.n6673 VGND 5.93e-19
C29259 VPWR.n6674 VGND 6.26e-19
C29260 VPWR.n6675 VGND 6.55e-19
C29261 VPWR.n6676 VGND 5.41e-19
C29262 VPWR.n6677 VGND 9.96e-19
C29263 VPWR.n6678 VGND 9.68e-19
C29264 VPWR.n6679 VGND 5.41e-19
C29265 VPWR.n6680 VGND 3.13e-19
C29266 VPWR.n6681 VGND 5.98e-19
C29267 VPWR.n6682 VGND 5.12e-19
C29268 VPWR.n6683 VGND 0.00108f
C29269 VPWR.n6684 VGND 0.00122f
C29270 VPWR.n6685 VGND 3.13e-19
C29271 VPWR.n6686 VGND 5.12e-19
C29272 VPWR.n6687 VGND 6.26e-19
C29273 VPWR.n6688 VGND 4.61e-20
C29274 VPWR.n6689 VGND 4.67e-19
C29275 VPWR.n6690 VGND 0.00128f
C29276 VPWR.n6691 VGND 0.00179f
C29277 VPWR.n6692 VGND 0.00279f
C29278 VPWR.n6693 VGND 0.00282f
C29279 VPWR.n6694 VGND 0.00961f
C29280 VPWR.n6695 VGND 0.00142f
C29281 VPWR.n6696 VGND 0.00115f
C29282 VPWR.n6697 VGND 0.0031f
C29283 VPWR.n6698 VGND 0.00639f
C29284 VPWR.n6699 VGND 0.00524f
C29285 VPWR.n6700 VGND 0.0066f
C29286 VPWR.n6701 VGND 0.00524f
C29287 VPWR.n6702 VGND 0.0066f
C29288 VPWR.n6703 VGND 0.00524f
C29289 VPWR.t1708 VGND 9.71e-19
C29290 VPWR.t866 VGND 9.22e-19
C29291 VPWR.n6704 VGND 0.00196f
C29292 VPWR.n6705 VGND 0.00666f
C29293 VPWR.n6706 VGND 0.00452f
C29294 VPWR.n6707 VGND 0.00524f
C29295 VPWR.n6708 VGND 0.00538f
C29296 VPWR.n6709 VGND 0.00524f
C29297 VPWR.t894 VGND 6.73e-19
C29298 VPWR.t892 VGND 6.73e-19
C29299 VPWR.n6710 VGND 0.00141f
C29300 VPWR.n6711 VGND 0.00621f
C29301 VPWR.n6712 VGND 0.0042f
C29302 VPWR.n6713 VGND 0.00524f
C29303 VPWR.t3501 VGND 0.0592f
C29304 VPWR.n6714 VGND 0.0356f
C29305 VPWR.n6715 VGND 0.00395f
C29306 VPWR.n6716 VGND 0.00524f
C29307 VPWR.n6717 VGND 0.00506f
C29308 VPWR.n6718 VGND 0.00524f
C29309 VPWR.n6719 VGND 0.00617f
C29310 VPWR.n6720 VGND 0.00524f
C29311 VPWR.t3134 VGND 0.00231f
C29312 VPWR.n6721 VGND 0.00736f
C29313 VPWR.n6722 VGND 0.00352f
C29314 VPWR.n6723 VGND 0.00524f
C29315 VPWR.n6724 VGND 0.00475f
C29316 VPWR.n6725 VGND 0.00259f
C29317 VPWR.n6726 VGND 0.00264f
C29318 VPWR.n6727 VGND 0.0031f
C29319 VPWR.n6728 VGND 0.00614f
C29320 VPWR.n6729 VGND 0.00524f
C29321 VPWR.n6730 VGND 0.0066f
C29322 VPWR.n6731 VGND 0.00524f
C29323 VPWR.t1283 VGND 8.82e-19
C29324 VPWR.t1467 VGND 0.00144f
C29325 VPWR.n6732 VGND 0.00521f
C29326 VPWR.n6733 VGND 0.00825f
C29327 VPWR.n6734 VGND 0.00409f
C29328 VPWR.n6735 VGND 0.00524f
C29329 VPWR.n6736 VGND 0.00581f
C29330 VPWR.n6737 VGND 0.00524f
C29331 VPWR.n6738 VGND 0.00629f
C29332 VPWR.n6739 VGND 0.00393f
C29333 VPWR.t263 VGND 0.00387f
C29334 VPWR.n6740 VGND 0.0107f
C29335 VPWR.n6741 VGND 0.00796f
C29336 VPWR.n6742 VGND 0.0031f
C29337 VPWR.t3362 VGND 0.0592f
C29338 VPWR.n6743 VGND 0.0416f
C29339 VPWR.n6744 VGND 0.013f
C29340 VPWR.n6745 VGND 0.00524f
C29341 VPWR.n6746 VGND 0.0142f
C29342 VPWR.n6747 VGND 0.00524f
C29343 VPWR.n6748 VGND 0.00524f
C29344 VPWR.n6749 VGND 0.00524f
C29345 VPWR.n6750 VGND 0.00793f
C29346 VPWR.t262 VGND 0.00387f
C29347 VPWR.n6751 VGND 0.0169f
C29348 VPWR.n6752 VGND 0.00679f
C29349 VPWR.t374 VGND 0.0046f
C29350 VPWR.t3368 VGND 0.0156f
C29351 VPWR.n6753 VGND 0.00623f
C29352 VPWR.n6754 VGND 0.0237f
C29353 VPWR.n6755 VGND 0.00507f
C29354 VPWR.n6756 VGND 0.0185f
C29355 VPWR.n6757 VGND 0.0136f
C29356 VPWR.n6758 VGND 0.018f
C29357 VPWR.n6759 VGND 0.00569f
C29358 VPWR.n6760 VGND 0.00907f
C29359 VPWR.n6761 VGND 0.00475f
C29360 VPWR.n6762 VGND 0.00279f
C29361 VPWR.n6763 VGND 0.00199f
C29362 VPWR.n6764 VGND 0.00282f
C29363 VPWR.n6765 VGND 0.0145f
C29364 VPWR.n6766 VGND 0.00535f
C29365 VPWR.n6767 VGND 0.0031f
C29366 VPWR.n6768 VGND 0.011f
C29367 VPWR.n6769 VGND 0.00524f
C29368 VPWR.n6770 VGND 0.0113f
C29369 VPWR.n6771 VGND 0.00524f
C29370 VPWR.t3537 VGND 0.0592f
C29371 VPWR.n6772 VGND 0.038f
C29372 VPWR.n6773 VGND 0.00833f
C29373 VPWR.n6774 VGND 0.00524f
C29374 VPWR.n6775 VGND 0.0087f
C29375 VPWR.n6776 VGND 0.00524f
C29376 VPWR.n6777 VGND 0.0113f
C29377 VPWR.n6778 VGND 0.00524f
C29378 VPWR.n6779 VGND 0.00451f
C29379 VPWR.n6780 VGND 5.27e-19
C29380 VPWR.n6781 VGND 3.95e-19
C29381 VPWR.n6782 VGND 5.05e-19
C29382 VPWR.n6783 VGND 5.05e-19
C29383 VPWR.n6784 VGND 8.67e-19
C29384 VPWR.n6785 VGND 6.54e-19
C29385 VPWR.n6786 VGND 9.06e-19
C29386 VPWR.n6787 VGND 0.00139f
C29387 VPWR.n6788 VGND 5.48e-19
C29388 VPWR.n6789 VGND 3.07e-19
C29389 VPWR.n6790 VGND 0.00138f
C29390 VPWR.n6791 VGND 0.00217f
C29391 VPWR.t108 VGND 0.0046f
C29392 VPWR.n6792 VGND 0.00126f
C29393 VPWR.n6793 VGND 0.0053f
C29394 VPWR.n6794 VGND 9.6e-19
C29395 VPWR.n6795 VGND 8.02e-19
C29396 VPWR.n6796 VGND 4.27e-19
C29397 VPWR.n6797 VGND 9.25e-19
C29398 VPWR.n6798 VGND 4.27e-19
C29399 VPWR.t3508 VGND 0.0612f
C29400 VPWR.n6799 VGND 0.0318f
C29401 VPWR.n6800 VGND 0.00248f
C29402 VPWR.n6801 VGND 4.84e-19
C29403 VPWR.n6802 VGND 6.83e-19
C29404 VPWR.n6803 VGND 4.84e-19
C29405 VPWR.n6804 VGND 3.13e-19
C29406 VPWR.n6805 VGND 9.68e-19
C29407 VPWR.n6806 VGND 0.00314f
C29408 VPWR.n6807 VGND 2.56e-19
C29409 VPWR.n6808 VGND 4.55e-19
C29410 VPWR.n6809 VGND 2.56e-19
C29411 VPWR.t602 VGND 0.0046f
C29412 VPWR.n6810 VGND 0.00613f
C29413 VPWR.n6811 VGND 0.00105f
C29414 VPWR.n6812 VGND 3.7e-19
C29415 VPWR.n6813 VGND 3.13e-19
C29416 VPWR.n6814 VGND 7.4e-19
C29417 VPWR.n6815 VGND 5.41e-19
C29418 VPWR.n6816 VGND 9.96e-19
C29419 VPWR.n6817 VGND 9.68e-19
C29420 VPWR.n6818 VGND 3.7e-19
C29421 VPWR.n6819 VGND 6.83e-19
C29422 VPWR.n6820 VGND 0.00105f
C29423 VPWR.n6821 VGND 0.0053f
C29424 VPWR.n6822 VGND 4.27e-19
C29425 VPWR.n6823 VGND 1.14e-19
C29426 VPWR.n6824 VGND 4.27e-19
C29427 VPWR.n6825 VGND 0.00567f
C29428 VPWR.n6826 VGND 0.00153f
C29429 VPWR.n6827 VGND 0.00206f
C29430 VPWR.n6828 VGND 0.00138f
C29431 VPWR.n6829 VGND 9e-19
C29432 VPWR.n6830 VGND 6.14e-19
C29433 VPWR.n6831 VGND 9.06e-19
C29434 VPWR.n6832 VGND 5.48e-19
C29435 VPWR.n6833 VGND 0.00138f
C29436 VPWR.n6834 VGND 0.0057f
C29437 VPWR.n6835 VGND 6.54e-19
C29438 VPWR.n6836 VGND 8.67e-19
C29439 VPWR.n6837 VGND 4.39e-19
C29440 VPWR.n6838 VGND 3.29e-19
C29441 VPWR.n6839 VGND 5.27e-19
C29442 VPWR.n6840 VGND 2.85e-19
C29443 VPWR.n6841 VGND 2.85e-19
C29444 VPWR.n6842 VGND 4.17e-19
C29445 VPWR.n6843 VGND 5.71e-19
C29446 VPWR.n6844 VGND 4.17e-19
C29447 VPWR.n6845 VGND 3.51e-19
C29448 VPWR.n6846 VGND 4.61e-19
C29449 VPWR.n6847 VGND 4.17e-19
C29450 VPWR.n6848 VGND 4.83e-19
C29451 VPWR.n6849 VGND 4.61e-19
C29452 VPWR.n6850 VGND 3.73e-19
C29453 VPWR.n6851 VGND 2.41e-19
C29454 VPWR.n6852 VGND 4.83e-19
C29455 VPWR.n6853 VGND 4.61e-19
C29456 VPWR.n6854 VGND 4.11e-19
C29457 VPWR.n6855 VGND 4.11e-19
C29458 VPWR.n6856 VGND 7.39e-19
C29459 VPWR.n6857 VGND 5.19e-19
C29460 VPWR.n6858 VGND 7.39e-19
C29461 VPWR.n6859 VGND 4.11e-19
C29462 VPWR.n6860 VGND 4.11e-19
C29463 VPWR.n6862 VGND 0.1f
C29464 VPWR.n6863 VGND 0.1f
C29465 VPWR.n6865 VGND 0.00139f
C29466 VPWR.n6866 VGND 5.48e-19
C29467 VPWR.n6867 VGND 3.07e-19
C29468 VPWR.n6868 VGND 0.00138f
C29469 VPWR.n6869 VGND 0.00217f
C29470 VPWR.t58 VGND 0.0046f
C29471 VPWR.n6870 VGND 0.00126f
C29472 VPWR.n6871 VGND 0.0053f
C29473 VPWR.n6872 VGND 9.6e-19
C29474 VPWR.n6873 VGND 8.02e-19
C29475 VPWR.n6874 VGND 4.27e-19
C29476 VPWR.n6875 VGND 9.25e-19
C29477 VPWR.n6876 VGND 4.27e-19
C29478 VPWR.t3507 VGND 0.0612f
C29479 VPWR.n6877 VGND 0.0319f
C29480 VPWR.n6878 VGND 0.00225f
C29481 VPWR.n6879 VGND 4.84e-19
C29482 VPWR.n6880 VGND 6.83e-19
C29483 VPWR.n6881 VGND 4.84e-19
C29484 VPWR.n6882 VGND 1.99e-19
C29485 VPWR.n6883 VGND 8.26e-19
C29486 VPWR.n6884 VGND 4.83e-19
C29487 VPWR.n6885 VGND 4.61e-19
C29488 VPWR.n6886 VGND 4.11e-19
C29489 VPWR.n6887 VGND 4.11e-19
C29490 VPWR.n6888 VGND 7.39e-19
C29491 VPWR.n6889 VGND 5.19e-19
C29492 VPWR.n6890 VGND 7.39e-19
C29493 VPWR.n6891 VGND 4.11e-19
C29494 VPWR.n6892 VGND 4.11e-19
C29495 VPWR.n6894 VGND 0.0581f
C29496 VPWR.n6895 VGND 0.59f
C29497 VPWR.n6896 VGND 0.0452f
C29498 VPWR.n6897 VGND 0.00626f
C29499 VPWR.n6898 VGND 6.54e-19
C29500 VPWR.n6899 VGND 8.67e-19
C29501 VPWR.n6900 VGND 4.11e-19
C29502 VPWR.n6901 VGND 7.39e-19
C29503 VPWR.n6902 VGND 5.19e-19
C29504 VPWR.n6903 VGND 7.39e-19
C29505 VPWR.n6904 VGND 4.11e-19
C29506 VPWR.n6905 VGND 4.39e-19
C29507 VPWR.n6906 VGND 3.29e-19
C29508 VPWR.n6907 VGND 5.27e-19
C29509 VPWR.n6908 VGND 2.85e-19
C29510 VPWR.n6909 VGND 2.85e-19
C29511 VPWR.n6910 VGND 4.17e-19
C29512 VPWR.n6911 VGND 5.71e-19
C29513 VPWR.n6912 VGND 4.17e-19
C29514 VPWR.n6913 VGND 3.51e-19
C29515 VPWR.n6914 VGND 4.61e-19
C29516 VPWR.n6915 VGND 4.17e-19
C29517 VPWR.n6916 VGND 4.11e-19
C29518 VPWR.n6918 VGND 0.00138f
C29519 VPWR.n6919 VGND 9e-19
C29520 VPWR.n6920 VGND 6.14e-19
C29521 VPWR.n6921 VGND 9.06e-19
C29522 VPWR.n6922 VGND 5.48e-19
C29523 VPWR.n6923 VGND 0.00138f
C29524 VPWR.n6924 VGND 0.0057f
C29525 VPWR.n6925 VGND 4.83e-19
C29526 VPWR.n6926 VGND 4.61e-19
C29527 VPWR.n6927 VGND 2.41e-19
C29528 VPWR.n6928 VGND 4.83e-19
C29529 VPWR.n6929 VGND 4.61e-19
C29530 VPWR.n6930 VGND 4.11e-19
C29531 VPWR.n6931 VGND 8.67e-19
C29532 VPWR.n6932 VGND 6.54e-19
C29533 VPWR.n6933 VGND 9.06e-19
C29534 VPWR.n6934 VGND 0.00139f
C29535 VPWR.n6935 VGND 3.73e-19
C29536 VPWR.n6936 VGND 5.27e-19
C29537 VPWR.n6937 VGND 3.95e-19
C29538 VPWR.n6938 VGND 5.05e-19
C29539 VPWR.n6939 VGND 5.05e-19
C29540 VPWR.n6940 VGND 0.00632f
C29541 VPWR.t144 VGND 0.0046f
C29542 VPWR.n6941 VGND 0.00407f
C29543 VPWR.t2058 VGND 0.00663f
C29544 VPWR.n6942 VGND 0.00884f
C29545 VPWR.t718 VGND 0.0301f
C29546 VPWR.t2379 VGND 0.0311f
C29547 VPWR.t2375 VGND 0.0164f
C29548 VPWR.t2377 VGND 0.0164f
C29549 VPWR.t2373 VGND 0.0173f
C29550 VPWR.t742 VGND 0.0154f
C29551 VPWR.t1488 VGND 0.0197f
C29552 VPWR.t1486 VGND 0.017f
C29553 VPWR.t939 VGND 0.0152f
C29554 VPWR.t640 VGND 0.0263f
C29555 VPWR.t142 VGND 0.105f
C29556 VPWR.n6943 VGND 0.0243f
C29557 VPWR.t2056 VGND -2.18e-20
C29558 VPWR.t2821 VGND 0.00137f
C29559 VPWR.n6944 VGND 0.00629f
C29560 VPWR.n6945 VGND 0.0079f
C29561 VPWR.t434 VGND 0.00387f
C29562 VPWR.t3430 VGND 0.0179f
C29563 VPWR.n6946 VGND 0.0133f
C29564 VPWR.n6947 VGND 0.0103f
C29565 VPWR.n6948 VGND 0.0173f
C29566 VPWR.n6949 VGND 0.00493f
C29567 VPWR.n6950 VGND 0.00525f
C29568 VPWR.t435 VGND 0.00387f
C29569 VPWR.n6951 VGND 0.00837f
C29570 VPWR.t120 VGND 0.0046f
C29571 VPWR.n6952 VGND 0.00407f
C29572 VPWR.t2304 VGND 0.00663f
C29573 VPWR.n6953 VGND 0.00913f
C29574 VPWR.n6954 VGND 0.00156f
C29575 VPWR.t2057 VGND 0.0214f
C29576 VPWR.t2055 VGND 0.017f
C29577 VPWR.t2820 VGND 0.0152f
C29578 VPWR.t433 VGND 0.0352f
C29579 VPWR.t119 VGND 0.105f
C29580 VPWR.t826 VGND 0.012f
C29581 VPWR.t2301 VGND 0.017f
C29582 VPWR.t2303 VGND 0.0319f
C29583 VPWR.n6955 VGND 0.03f
C29584 VPWR.t669 VGND 0.0046f
C29585 VPWR.n6956 VGND 0.00371f
C29586 VPWR.n6957 VGND 3.95e-19
C29587 VPWR.n6958 VGND 3.29e-19
C29588 VPWR.n6959 VGND 5.71e-19
C29589 VPWR.n6960 VGND 5.92e-19
C29590 VPWR.n6961 VGND 5.05e-19
C29591 VPWR.n6962 VGND 4.83e-19
C29592 VPWR.n6963 VGND 2.85e-19
C29593 VPWR.n6964 VGND 3.95e-19
C29594 VPWR.n6965 VGND 4.17e-19
C29595 VPWR.n6966 VGND 2.85e-19
C29596 VPWR.n6967 VGND 2.85e-19
C29597 VPWR.n6968 VGND 4.11e-19
C29598 VPWR.n6969 VGND 8.67e-19
C29599 VPWR.n6970 VGND 6.54e-19
C29600 VPWR.n6971 VGND 9.06e-19
C29601 VPWR.n6972 VGND 0.00626f
C29602 VPWR.n6973 VGND 6.54e-19
C29603 VPWR.n6974 VGND 8.67e-19
C29604 VPWR.n6975 VGND 4.11e-19
C29605 VPWR.n6976 VGND 7.39e-19
C29606 VPWR.n6977 VGND 5.19e-19
C29607 VPWR.n6978 VGND 7.39e-19
C29608 VPWR.n6979 VGND 4.11e-19
C29609 VPWR.n6980 VGND 3.95e-19
C29610 VPWR.n6981 VGND 4.61e-19
C29611 VPWR.n6982 VGND 2.41e-19
C29612 VPWR.n6983 VGND 3.95e-19
C29613 VPWR.n6984 VGND 5.05e-19
C29614 VPWR.n6985 VGND 4.17e-19
C29615 VPWR.n6986 VGND 6.14e-19
C29616 VPWR.n6987 VGND 4.39e-19
C29617 VPWR.n6988 VGND 1.76e-19
C29618 VPWR.n6989 VGND 3.07e-19
C29619 VPWR.n6990 VGND 4.11e-19
C29620 VPWR.n6992 VGND 8.11e-19
C29621 VPWR.n6993 VGND 3.95e-19
C29622 VPWR.n6994 VGND 1.77e-19
C29623 VPWR.n6995 VGND 3.95e-19
C29624 VPWR.n6996 VGND 7.68e-19
C29625 VPWR.n6997 VGND 5.05e-19
C29626 VPWR.n6998 VGND 1.76e-19
C29627 VPWR.n6999 VGND 9.06e-19
C29628 VPWR.n7000 VGND 5.48e-19
C29629 VPWR.n7001 VGND 0.00138f
C29630 VPWR.n7002 VGND 0.0057f
C29631 VPWR.n7003 VGND 6.54e-19
C29632 VPWR.n7004 VGND 8.67e-19
C29633 VPWR.n7005 VGND 4.11e-19
C29634 VPWR.n7006 VGND 7.39e-19
C29635 VPWR.n7007 VGND 5.19e-19
C29636 VPWR.n7008 VGND 7.39e-19
C29637 VPWR.n7009 VGND 4.11e-19
C29638 VPWR.n7010 VGND 3.95e-19
C29639 VPWR.n7011 VGND 4.61e-19
C29640 VPWR.n7012 VGND 2.41e-19
C29641 VPWR.n7013 VGND 3.95e-19
C29642 VPWR.n7014 VGND 5.05e-19
C29643 VPWR.n7015 VGND 4.17e-19
C29644 VPWR.n7016 VGND 6.14e-19
C29645 VPWR.n7017 VGND 4.39e-19
C29646 VPWR.n7018 VGND 1.76e-19
C29647 VPWR.n7019 VGND 3.07e-19
C29648 VPWR.n7020 VGND 4.11e-19
C29649 VPWR.n7022 VGND 0.1f
C29650 VPWR.n7023 VGND 0.1f
C29651 VPWR.n7025 VGND 0.00139f
C29652 VPWR.n7026 VGND 5.48e-19
C29653 VPWR.n7027 VGND 4.17e-19
C29654 VPWR.n7028 VGND 0.00137f
C29655 VPWR.n7029 VGND 0.0066f
C29656 VPWR.t670 VGND 0.0046f
C29657 VPWR.n7030 VGND 0.00407f
C29658 VPWR.t3206 VGND 0.00137f
C29659 VPWR.t3242 VGND -2.18e-20
C29660 VPWR.n7031 VGND 0.00629f
C29661 VPWR.n7032 VGND 0.0079f
C29662 VPWR.t3244 VGND 0.00663f
C29663 VPWR.n7033 VGND 0.00913f
C29664 VPWR.t578 VGND 0.00387f
C29665 VPWR.n7034 VGND 0.0127f
C29666 VPWR.n7035 VGND 0.0109f
C29667 VPWR.t3482 VGND 0.0156f
C29668 VPWR.n7036 VGND 0.00597f
C29669 VPWR.n7037 VGND 0.0228f
C29670 VPWR.n7038 VGND 0.00971f
C29671 VPWR.n7039 VGND 0.0109f
C29672 VPWR.n7040 VGND 0.011f
C29673 VPWR.n7041 VGND 0.00846f
C29674 VPWR.t579 VGND 0.00387f
C29675 VPWR.t431 VGND 0.00387f
C29676 VPWR.t3429 VGND 0.0179f
C29677 VPWR.n7042 VGND 0.0103f
C29678 VPWR.n7043 VGND 0.0173f
C29679 VPWR.n7044 VGND 0.00493f
C29680 VPWR.n7045 VGND 0.00487f
C29681 VPWR.t668 VGND 0.105f
C29682 VPWR.t3205 VGND 0.012f
C29683 VPWR.t3241 VGND 0.017f
C29684 VPWR.t3243 VGND 0.0228f
C29685 VPWR.t577 VGND 0.0703f
C29686 VPWR.n7046 VGND 0.0102f
C29687 VPWR.t175 VGND 0.0333f
C29688 VPWR.t2476 VGND 0.0311f
C29689 VPWR.t2472 VGND 0.0164f
C29690 VPWR.t2478 VGND 0.0164f
C29691 VPWR.t2474 VGND 0.0173f
C29692 VPWR.t3139 VGND 0.0122f
C29693 VPWR.t1476 VGND 0.0238f
C29694 VPWR.t1472 VGND 0.0164f
C29695 VPWR.t1470 VGND 0.0164f
C29696 VPWR.t1474 VGND 0.0173f
C29697 VPWR.t1956 VGND 0.0122f
C29698 VPWR.t1268 VGND 0.023f
C29699 VPWR.t1266 VGND 0.017f
C29700 VPWR.t2901 VGND 0.012f
C29701 VPWR.t469 VGND 0.0717f
C29702 VPWR.n7047 VGND 0.00487f
C29703 VPWR.n7048 VGND 0.00186f
C29704 VPWR.t456 VGND 0.0046f
C29705 VPWR.n7049 VGND 0.00407f
C29706 VPWR.t29 VGND 0.00387f
C29707 VPWR.n7050 VGND 0.00837f
C29708 VPWR.n7051 VGND 5.98e-19
C29709 VPWR.t2072 VGND 0.00695f
C29710 VPWR.n7052 VGND 0.0084f
C29711 VPWR.n7053 VGND 8.39e-20
C29712 VPWR.n7054 VGND 4.58e-19
C29713 VPWR.n7055 VGND 0.00256f
C29714 VPWR.n7056 VGND 0.00122f
C29715 VPWR.n7057 VGND 0.00492f
C29716 VPWR.t2066 VGND 0.00166f
C29717 VPWR.t2068 VGND 0.00166f
C29718 VPWR.n7058 VGND 0.00345f
C29719 VPWR.n7059 VGND 0.00502f
C29720 VPWR.n7060 VGND 0.00524f
C29721 VPWR.n7061 VGND 0.00121f
C29722 VPWR.n7062 VGND 0.00524f
C29723 VPWR.t2070 VGND 0.00225f
C29724 VPWR.t2292 VGND 0.00166f
C29725 VPWR.n7063 VGND 0.0045f
C29726 VPWR.n7064 VGND 0.00778f
C29727 VPWR.n7065 VGND 0.00524f
C29728 VPWR.n7066 VGND 0.00131f
C29729 VPWR.n7067 VGND 0.0031f
C29730 VPWR.n7068 VGND 0.00199f
C29731 VPWR.n7069 VGND 0.00199f
C29732 VPWR.n7070 VGND 0.00143f
C29733 VPWR.t28 VGND 0.00387f
C29734 VPWR.t3551 VGND 0.0179f
C29735 VPWR.n7071 VGND 0.0133f
C29736 VPWR.n7072 VGND 0.0103f
C29737 VPWR.n7073 VGND 0.0173f
C29738 VPWR.n7074 VGND 0.00493f
C29739 VPWR.n7075 VGND 0.00525f
C29740 VPWR.n7076 VGND 0.00393f
C29741 VPWR.n7077 VGND 0.00524f
C29742 VPWR.n7078 VGND 0.00524f
C29743 VPWR.n7079 VGND 0.0031f
C29744 VPWR.n7080 VGND 0.00515f
C29745 VPWR.t455 VGND 0.0046f
C29746 VPWR.n7081 VGND 0.00407f
C29747 VPWR.n7082 VGND 0.00256f
C29748 VPWR.n7083 VGND 0.00393f
C29749 VPWR.n7084 VGND 0.00639f
C29750 VPWR.n7085 VGND 0.00524f
C29751 VPWR.n7086 VGND 0.0066f
C29752 VPWR.n7087 VGND 0.00524f
C29753 VPWR.n7088 VGND 0.00506f
C29754 VPWR.n7089 VGND 0.00524f
C29755 VPWR.t3437 VGND 0.0592f
C29756 VPWR.n7090 VGND 0.0356f
C29757 VPWR.n7091 VGND 0.00484f
C29758 VPWR.n7092 VGND 0.00524f
C29759 VPWR.n7093 VGND 0.0066f
C29760 VPWR.n7094 VGND 0.00524f
C29761 VPWR.n7095 VGND 0.0066f
C29762 VPWR.n7096 VGND 0.00524f
C29763 VPWR.n7097 VGND 0.0066f
C29764 VPWR.n7098 VGND 0.00524f
C29765 VPWR.n7099 VGND 0.0066f
C29766 VPWR.n7100 VGND 0.00524f
C29767 VPWR.n7101 VGND 0.0066f
C29768 VPWR.n7102 VGND 0.00524f
C29769 VPWR.n7103 VGND 0.00639f
C29770 VPWR.n7104 VGND 0.00524f
C29771 VPWR.n7105 VGND 0.0031f
C29772 VPWR.n7106 VGND 0.0024f
C29773 VPWR.t886 VGND 0.00654f
C29774 VPWR.n7107 VGND 0.011f
C29775 VPWR.n7108 VGND 0.00475f
C29776 VPWR.n7109 VGND 0.00146f
C29777 VPWR.n7110 VGND 0.00524f
C29778 VPWR.n7111 VGND 0.00307f
C29779 VPWR.n7112 VGND 0.00179f
C29780 VPWR.n7113 VGND 0.00159f
C29781 VPWR.t1893 VGND 0.00137f
C29782 VPWR.t845 VGND -2.18e-20
C29783 VPWR.n7114 VGND 0.00629f
C29784 VPWR.n7115 VGND 0.0079f
C29785 VPWR.n7116 VGND 0.00475f
C29786 VPWR.n7117 VGND 0.00121f
C29787 VPWR.n7118 VGND 0.00524f
C29788 VPWR.t843 VGND 0.00663f
C29789 VPWR.t13 VGND 0.00391f
C29790 VPWR.t3545 VGND 0.00886f
C29791 VPWR.t14 VGND 0.00391f
C29792 VPWR.n7119 VGND 0.00833f
C29793 VPWR.n7120 VGND 0.0116f
C29794 VPWR.n7121 VGND 0.0146f
C29795 VPWR.n7122 VGND 0.00317f
C29796 VPWR.n7123 VGND 0.00488f
C29797 VPWR.n7124 VGND 0.00909f
C29798 VPWR.n7125 VGND 0.00393f
C29799 VPWR.n7126 VGND 0.00393f
C29800 VPWR.n7127 VGND 0.00524f
C29801 VPWR.n7128 VGND 0.0031f
C29802 VPWR.n7129 VGND 0.00199f
C29803 VPWR.t470 VGND 0.00387f
C29804 VPWR.n7130 VGND 0.00846f
C29805 VPWR.n7131 VGND 0.00688f
C29806 VPWR.n7132 VGND 9.25e-19
C29807 VPWR.n7133 VGND 5.05e-19
C29808 VPWR.n7134 VGND 5.05e-19
C29809 VPWR.n7135 VGND 0.00138f
C29810 VPWR.n7136 VGND 0.00626f
C29811 VPWR.n7137 VGND 0.1f
C29812 VPWR.n7138 VGND 0.1f
C29813 VPWR.n7140 VGND 0.0057f
C29814 VPWR.n7142 VGND 0.00139f
C29815 VPWR.n7143 VGND 5.27e-19
C29816 VPWR.n7144 VGND 3.29e-19
C29817 VPWR.n7145 VGND 4.39e-19
C29818 VPWR.n7146 VGND 9e-19
C29819 VPWR.t1269 VGND 0.00663f
C29820 VPWR.n7147 VGND 0.00913f
C29821 VPWR.t1471 VGND 0.00166f
C29822 VPWR.t1473 VGND 0.00166f
C29823 VPWR.n7148 VGND 0.00345f
C29824 VPWR.n7149 VGND 0.00502f
C29825 VPWR.t1477 VGND 0.00695f
C29826 VPWR.n7150 VGND 0.00848f
C29827 VPWR.t3140 VGND 0.00166f
C29828 VPWR.t2475 VGND 0.00225f
C29829 VPWR.n7151 VGND 0.0045f
C29830 VPWR.n7152 VGND 0.00778f
C29831 VPWR.t2479 VGND 0.00166f
C29832 VPWR.t2473 VGND 0.00166f
C29833 VPWR.n7153 VGND 0.00345f
C29834 VPWR.n7154 VGND 0.00502f
C29835 VPWR.t2477 VGND 0.00695f
C29836 VPWR.n7155 VGND 0.0084f
C29837 VPWR.t176 VGND 0.00391f
C29838 VPWR.t3337 VGND 0.00886f
C29839 VPWR.t177 VGND 0.00391f
C29840 VPWR.n7156 VGND 0.0125f
C29841 VPWR.n7157 VGND 0.0116f
C29842 VPWR.n7158 VGND 0.0146f
C29843 VPWR.n7159 VGND 0.00317f
C29844 VPWR.n7160 VGND 0.00503f
C29845 VPWR.n7161 VGND 0.00338f
C29846 VPWR.n7162 VGND 0.00524f
C29847 VPWR.n7163 VGND 0.00393f
C29848 VPWR.n7164 VGND 0.00393f
C29849 VPWR.n7165 VGND 0.00122f
C29850 VPWR.n7166 VGND 0.00524f
C29851 VPWR.n7167 VGND 0.00524f
C29852 VPWR.n7168 VGND 0.00121f
C29853 VPWR.n7169 VGND 0.00524f
C29854 VPWR.n7170 VGND 0.00475f
C29855 VPWR.n7171 VGND 0.00179f
C29856 VPWR.n7172 VGND 0.0016f
C29857 VPWR.n7173 VGND 0.00167f
C29858 VPWR.n7174 VGND 0.00199f
C29859 VPWR.n7175 VGND 0.00393f
C29860 VPWR.n7176 VGND 0.00122f
C29861 VPWR.n7177 VGND 0.00524f
C29862 VPWR.n7178 VGND 0.00524f
C29863 VPWR.n7179 VGND 0.00121f
C29864 VPWR.n7180 VGND 0.00524f
C29865 VPWR.n7181 VGND 0.00475f
C29866 VPWR.t1957 VGND 0.00166f
C29867 VPWR.t1475 VGND 0.00225f
C29868 VPWR.n7182 VGND 0.0045f
C29869 VPWR.n7183 VGND 0.00778f
C29870 VPWR.n7184 VGND 0.00132f
C29871 VPWR.n7185 VGND 0.00179f
C29872 VPWR.n7186 VGND 0.00393f
C29873 VPWR.n7187 VGND 0.00121f
C29874 VPWR.n7188 VGND 0.00524f
C29875 VPWR.n7189 VGND 0.00475f
C29876 VPWR.t2902 VGND 0.00137f
C29877 VPWR.t1267 VGND -2.18e-20
C29878 VPWR.n7190 VGND 0.00629f
C29879 VPWR.n7191 VGND 0.0079f
C29880 VPWR.n7192 VGND 0.00136f
C29881 VPWR.n7193 VGND 0.00154f
C29882 VPWR.n7194 VGND 9.06e-19
C29883 VPWR.n7195 VGND 0.00112f
C29884 VPWR.n7196 VGND 4.27e-19
C29885 VPWR.n7197 VGND 0.0012f
C29886 VPWR.n7198 VGND 4.55e-19
C29887 VPWR.n7199 VGND 0.00516f
C29888 VPWR.n7200 VGND 4.84e-19
C29889 VPWR.n7201 VGND 6.83e-19
C29890 VPWR.n7202 VGND 4.84e-19
C29891 VPWR.n7203 VGND 3.13e-19
C29892 VPWR.n7204 VGND 9.96e-19
C29893 VPWR.n7205 VGND 0.00568f
C29894 VPWR.n7206 VGND 9.68e-19
C29895 VPWR.n7207 VGND 4.27e-19
C29896 VPWR.n7208 VGND 2.56e-19
C29897 VPWR.n7209 VGND 0.00127f
C29898 VPWR.n7210 VGND 0.00643f
C29899 VPWR.n7211 VGND 3.42e-19
C29900 VPWR.n7212 VGND 7.4e-19
C29901 VPWR.n7213 VGND 5.41e-19
C29902 VPWR.n7214 VGND 9.96e-19
C29903 VPWR.n7215 VGND 9.68e-19
C29904 VPWR.n7216 VGND 3.7e-19
C29905 VPWR.n7217 VGND 6.83e-19
C29906 VPWR.t471 VGND 0.00387f
C29907 VPWR.n7218 VGND 0.008f
C29908 VPWR.n7219 VGND 0.00127f
C29909 VPWR.n7220 VGND 4.48e-19
C29910 VPWR.n7221 VGND 4.27e-19
C29911 VPWR.n7222 VGND 8.54e-20
C29912 VPWR.n7223 VGND 4.27e-19
C29913 VPWR.n7224 VGND 0.00387f
C29914 VPWR.n7225 VGND 4.84e-19
C29915 VPWR.n7226 VGND 8.26e-19
C29916 VPWR.n7227 VGND 0.00138f
C29917 VPWR.n7228 VGND 6.14e-19
C29918 VPWR.n7229 VGND 5.48e-19
C29919 VPWR.n7230 VGND 9.06e-19
C29920 VPWR.n7231 VGND 6.54e-19
C29921 VPWR.n7232 VGND 8.67e-19
C29922 VPWR.n7233 VGND 4.17e-19
C29923 VPWR.n7234 VGND 5.71e-19
C29924 VPWR.n7235 VGND 4.17e-19
C29925 VPWR.n7236 VGND 3.51e-19
C29926 VPWR.n7237 VGND 4.61e-19
C29927 VPWR.n7238 VGND 2.85e-19
C29928 VPWR.n7239 VGND 2.85e-19
C29929 VPWR.n7240 VGND 4.17e-19
C29930 VPWR.n7241 VGND 4.11e-19
C29931 VPWR.n7242 VGND 4.11e-19
C29932 VPWR.n7243 VGND 7.39e-19
C29933 VPWR.n7244 VGND 5.19e-19
C29934 VPWR.n7245 VGND 7.39e-19
C29935 VPWR.n7246 VGND 4.11e-19
C29936 VPWR.n7247 VGND 3.95e-19
C29937 VPWR.n7248 VGND 5.27e-19
C29938 VPWR.n7249 VGND 3.73e-19
C29939 VPWR.n7250 VGND 2.41e-19
C29940 VPWR.n7251 VGND 4.83e-19
C29941 VPWR.n7252 VGND 4.83e-19
C29942 VPWR.n7253 VGND 4.61e-19
C29943 VPWR.n7254 VGND 4.61e-19
C29944 VPWR.n7255 VGND 4.11e-19
C29945 VPWR.n7256 VGND 8.67e-19
C29946 VPWR.n7257 VGND 6.54e-19
C29947 VPWR.n7258 VGND 9.06e-19
C29948 VPWR.n7259 VGND 5.48e-19
C29949 VPWR.n7260 VGND 3.07e-19
C29950 VPWR.n7261 VGND 0.00138f
C29951 VPWR.n7262 VGND 0.00222f
C29952 VPWR.n7263 VGND 0.013f
C29953 VPWR.n7264 VGND 0.00452f
C29954 VPWR.n7265 VGND 0.0127f
C29955 VPWR.n7266 VGND 0.00956f
C29956 VPWR.n7267 VGND 0.00524f
C29957 VPWR.t3442 VGND 0.0156f
C29958 VPWR.n7268 VGND 0.00597f
C29959 VPWR.n7269 VGND 0.0228f
C29960 VPWR.n7270 VGND 0.00971f
C29961 VPWR.n7271 VGND 0.0109f
C29962 VPWR.n7272 VGND 0.00524f
C29963 VPWR.n7273 VGND 0.011f
C29964 VPWR.n7274 VGND 0.0109f
C29965 VPWR.n7275 VGND 0.00524f
C29966 VPWR.n7276 VGND 0.00393f
C29967 VPWR.n7277 VGND 0.00684f
C29968 VPWR.n7278 VGND 0.0102f
C29969 VPWR.n7279 VGND 0.0503f
C29970 VPWR.t12 VGND 0.0326f
C29971 VPWR.t842 VGND 0.0302f
C29972 VPWR.t844 VGND 0.017f
C29973 VPWR.t1892 VGND 0.012f
C29974 VPWR.t2038 VGND 0.0129f
C29975 VPWR.t885 VGND 0.0201f
C29976 VPWR.t454 VGND 0.105f
C29977 VPWR.t27 VGND 0.0352f
C29978 VPWR.n7280 VGND 0.0211f
C29979 VPWR.t2291 VGND 0.0154f
C29980 VPWR.t2069 VGND 0.0173f
C29981 VPWR.t2067 VGND 0.0164f
C29982 VPWR.t2065 VGND 0.0164f
C29983 VPWR.t2071 VGND 0.0208f
C29984 VPWR.t557 VGND 0.0263f
C29985 VPWR.t2966 VGND 0.0146f
C29986 VPWR.t832 VGND 0.0201f
C29987 VPWR.t512 VGND 0.0352f
C29988 VPWR.t2221 VGND 0.0154f
C29989 VPWR.t2264 VGND 0.0173f
C29990 VPWR.t2268 VGND 0.0164f
C29991 VPWR.t2266 VGND 0.0164f
C29992 VPWR.t2270 VGND 0.0208f
C29993 VPWR.t430 VGND 0.0366f
C29994 VPWR.n7281 VGND 0.0328f
C29995 VPWR.n7282 VGND 0.0133f
C29996 VPWR.t432 VGND 0.00387f
C29997 VPWR.n7283 VGND 0.00837f
C29998 VPWR.t2267 VGND 0.00166f
C29999 VPWR.t2269 VGND 0.00166f
C30000 VPWR.n7284 VGND 0.00345f
C30001 VPWR.n7285 VGND 0.00502f
C30002 VPWR.t2265 VGND 0.00225f
C30003 VPWR.t2222 VGND 0.00166f
C30004 VPWR.n7286 VGND 0.0045f
C30005 VPWR.n7287 VGND 0.00778f
C30006 VPWR.t513 VGND 0.00387f
C30007 VPWR.n7288 VGND 0.00493f
C30008 VPWR.n7289 VGND 0.00525f
C30009 VPWR.t3458 VGND 0.0179f
C30010 VPWR.n7290 VGND 0.0173f
C30011 VPWR.n7291 VGND 0.0103f
C30012 VPWR.n7292 VGND 0.0133f
C30013 VPWR.t514 VGND 0.00387f
C30014 VPWR.n7293 VGND 0.00837f
C30015 VPWR.t833 VGND 0.00136f
C30016 VPWR.t2967 VGND 0.00136f
C30017 VPWR.n7294 VGND 0.00328f
C30018 VPWR.n7295 VGND 0.0079f
C30019 VPWR.t558 VGND 0.00391f
C30020 VPWR.t3473 VGND 0.00886f
C30021 VPWR.n7296 VGND 9.71e-19
C30022 VPWR.n7297 VGND 0.00516f
C30023 VPWR.n7298 VGND 0.0138f
C30024 VPWR.n7299 VGND 0.00317f
C30025 VPWR.n7300 VGND 7.68e-19
C30026 VPWR.n7301 VGND 3.95e-19
C30027 VPWR.n7302 VGND 3.95e-19
C30028 VPWR.n7303 VGND 4.83e-19
C30029 VPWR.n7304 VGND 2.41e-19
C30030 VPWR.n7305 VGND 3.73e-19
C30031 VPWR.n7306 VGND 3.07e-19
C30032 VPWR.n7307 VGND 1.76e-19
C30033 VPWR.n7308 VGND 4.39e-19
C30034 VPWR.n7309 VGND 6.14e-19
C30035 VPWR.n7310 VGND 4.17e-19
C30036 VPWR.n7311 VGND 5.05e-19
C30037 VPWR.n7312 VGND 4.83e-19
C30038 VPWR.n7313 VGND 2.85e-19
C30039 VPWR.n7314 VGND 3.95e-19
C30040 VPWR.n7315 VGND 2.85e-19
C30041 VPWR.n7316 VGND 2.85e-19
C30042 VPWR.n7317 VGND 4.17e-19
C30043 VPWR.n7318 VGND 3.95e-19
C30044 VPWR.n7319 VGND 3.29e-19
C30045 VPWR.n7320 VGND 5.71e-19
C30046 VPWR.n7321 VGND 5.92e-19
C30047 VPWR.n7322 VGND 5.05e-19
C30048 VPWR.n7323 VGND 4.17e-19
C30049 VPWR.n7324 VGND 0.00138f
C30050 VPWR.n7325 VGND 8.32e-19
C30051 VPWR.n7326 VGND 2.28e-19
C30052 VPWR.n7327 VGND 4.84e-19
C30053 VPWR.n7328 VGND 9.71e-19
C30054 VPWR.n7329 VGND 0.0062f
C30055 VPWR.t559 VGND 0.00391f
C30056 VPWR.n7330 VGND 0.00736f
C30057 VPWR.n7331 VGND 0.00503f
C30058 VPWR.n7332 VGND 3.13e-19
C30059 VPWR.n7333 VGND 5.12e-19
C30060 VPWR.n7334 VGND 9.68e-19
C30061 VPWR.n7335 VGND 9.96e-19
C30062 VPWR.n7336 VGND 5.41e-19
C30063 VPWR.n7337 VGND 6.55e-19
C30064 VPWR.n7338 VGND 6.26e-19
C30065 VPWR.n7339 VGND 3.7e-19
C30066 VPWR.n7340 VGND 3.7e-19
C30067 VPWR.n7341 VGND 3.7e-19
C30068 VPWR.n7342 VGND 5.12e-19
C30069 VPWR.n7343 VGND 5.41e-19
C30070 VPWR.n7344 VGND 5.12e-19
C30071 VPWR.n7345 VGND 4.27e-19
C30072 VPWR.n7346 VGND 9.96e-19
C30073 VPWR.n7347 VGND 0.00131f
C30074 VPWR.n7348 VGND 5.98e-19
C30075 VPWR.n7349 VGND 6.99e-19
C30076 VPWR.n7350 VGND 0.00525f
C30077 VPWR.n7351 VGND 0.00139f
C30078 VPWR.n7352 VGND 0.0031f
C30079 VPWR.n7353 VGND 0.00524f
C30080 VPWR.n7354 VGND 0.00393f
C30081 VPWR.n7355 VGND 0.00139f
C30082 VPWR.n7356 VGND 0.00525f
C30083 VPWR.n7357 VGND 0.0031f
C30084 VPWR.n7358 VGND 0.00524f
C30085 VPWR.n7359 VGND 0.00524f
C30086 VPWR.n7360 VGND 0.00393f
C30087 VPWR.n7361 VGND 0.00199f
C30088 VPWR.n7362 VGND 0.00173f
C30089 VPWR.n7363 VGND 0.0016f
C30090 VPWR.n7364 VGND 0.0031f
C30091 VPWR.n7365 VGND 0.00524f
C30092 VPWR.n7366 VGND 0.00121f
C30093 VPWR.n7367 VGND 0.00524f
C30094 VPWR.n7368 VGND 0.00524f
C30095 VPWR.n7369 VGND 0.00122f
C30096 VPWR.n7370 VGND 0.00524f
C30097 VPWR.n7371 VGND 0.00393f
C30098 VPWR.t2271 VGND 0.00695f
C30099 VPWR.n7372 VGND 0.0084f
C30100 VPWR.n7373 VGND 0.00503f
C30101 VPWR.n7374 VGND 0.0031f
C30102 VPWR.n7375 VGND 0.00524f
C30103 VPWR.n7376 VGND 0.00524f
C30104 VPWR.n7377 VGND 0.00393f
C30105 VPWR.n7378 VGND 0.00199f
C30106 VPWR.n7379 VGND 0.0102f
C30107 VPWR.n7380 VGND 0.00487f
C30108 VPWR.n7381 VGND 0.00837f
C30109 VPWR.n7382 VGND 0.0133f
C30110 VPWR.n7383 VGND 0.00524f
C30111 VPWR.n7384 VGND 0.0138f
C30112 VPWR.n7385 VGND 0.00524f
C30113 VPWR.n7386 VGND 0.0135f
C30114 VPWR.n7387 VGND 0.00524f
C30115 VPWR.n7388 VGND 0.00956f
C30116 VPWR.n7389 VGND 0.00524f
C30117 VPWR.n7390 VGND 0.00524f
C30118 VPWR.n7391 VGND 0.00524f
C30119 VPWR.n7392 VGND 0.00393f
C30120 VPWR.n7393 VGND 0.00724f
C30121 VPWR.n7394 VGND 0.00144f
C30122 VPWR.n7395 VGND 0.00199f
C30123 VPWR.n7396 VGND 0.00393f
C30124 VPWR.n7397 VGND 0.00121f
C30125 VPWR.n7398 VGND 0.00524f
C30126 VPWR.n7399 VGND 0.00475f
C30127 VPWR.n7400 VGND 0.00262f
C30128 VPWR.n7401 VGND 0.00149f
C30129 VPWR.n7402 VGND 0.00274f
C30130 VPWR.n7403 VGND 0.0031f
C30131 VPWR.n7404 VGND 0.00639f
C30132 VPWR.n7405 VGND 0.00524f
C30133 VPWR.n7406 VGND 0.0066f
C30134 VPWR.n7407 VGND 0.00524f
C30135 VPWR.n7408 VGND 0.0066f
C30136 VPWR.n7409 VGND 0.00524f
C30137 VPWR.n7410 VGND 0.0066f
C30138 VPWR.n7411 VGND 0.00524f
C30139 VPWR.n7412 VGND 0.0066f
C30140 VPWR.n7413 VGND 0.00524f
C30141 VPWR.n7414 VGND 0.00503f
C30142 VPWR.n7415 VGND 0.00218f
C30143 VPWR.t3506 VGND 0.0592f
C30144 VPWR.n7416 VGND 0.0352f
C30145 VPWR.n7417 VGND 0.00484f
C30146 VPWR.n7418 VGND 6.8e-19
C30147 VPWR.n7419 VGND 5.69e-19
C30148 VPWR.n7420 VGND 0.00131f
C30149 VPWR.n7421 VGND 9.96e-19
C30150 VPWR.n7422 VGND 4.27e-19
C30151 VPWR.n7423 VGND 5.12e-19
C30152 VPWR.n7424 VGND 5.41e-19
C30153 VPWR.n7425 VGND 0.00176f
C30154 VPWR.n7426 VGND 5.41e-19
C30155 VPWR.n7427 VGND 4.66e-19
C30156 VPWR.n7428 VGND 3.7e-19
C30157 VPWR.n7429 VGND 4.31e-19
C30158 VPWR.n7430 VGND 3.42e-19
C30159 VPWR.n7431 VGND 0.00323f
C30160 VPWR.n7432 VGND 3.7e-19
C30161 VPWR.n7433 VGND 6.26e-19
C30162 VPWR.n7434 VGND 6.55e-19
C30163 VPWR.n7435 VGND 5.41e-19
C30164 VPWR.n7436 VGND 9.96e-19
C30165 VPWR.n7437 VGND 9.68e-19
C30166 VPWR.n7438 VGND 5.41e-19
C30167 VPWR.n7439 VGND 0.00592f
C30168 VPWR.n7440 VGND 3.13e-19
C30169 VPWR.n7441 VGND 5.98e-19
C30170 VPWR.n7442 VGND 5.12e-19
C30171 VPWR.n7443 VGND 0.00108f
C30172 VPWR.n7444 VGND 0.00122f
C30173 VPWR.n7445 VGND 3.13e-19
C30174 VPWR.n7446 VGND 5.12e-19
C30175 VPWR.n7447 VGND 0.0033f
C30176 VPWR.n7448 VGND 6.26e-19
C30177 VPWR.n7449 VGND 6.1e-19
C30178 VPWR.n7450 VGND 2.28e-19
C30179 VPWR.n7451 VGND 2.85e-19
C30180 VPWR.n7452 VGND 0.00309f
C30181 VPWR.n7453 VGND 0.00259f
C30182 VPWR.n7454 VGND 0.00364f
C30183 VPWR.n7455 VGND 0.00269f
C30184 VPWR.n7456 VGND 0.00175f
C30185 VPWR.n7457 VGND 0.00333f
C30186 VPWR.n7458 VGND 0.00393f
C30187 VPWR.n7459 VGND 0.00199f
C30188 VPWR.n7460 VGND 0.0102f
C30189 VPWR.n7461 VGND 0.00156f
C30190 VPWR.n7462 VGND 0.00333f
C30191 VPWR.n7463 VGND 0.00157f
C30192 VPWR.n7464 VGND 0.00393f
C30193 VPWR.n7465 VGND 0.00393f
C30194 VPWR.n7466 VGND 0.00121f
C30195 VPWR.n7467 VGND 0.00524f
C30196 VPWR.n7468 VGND 0.00475f
C30197 VPWR.t827 VGND 0.00137f
C30198 VPWR.t2302 VGND -2.18e-20
C30199 VPWR.n7469 VGND 0.00629f
C30200 VPWR.n7470 VGND 0.0079f
C30201 VPWR.n7471 VGND 0.00149f
C30202 VPWR.n7472 VGND 0.00262f
C30203 VPWR.t121 VGND 0.0046f
C30204 VPWR.n7473 VGND 0.00407f
C30205 VPWR.n7474 VGND 0.00274f
C30206 VPWR.n7475 VGND 0.0031f
C30207 VPWR.n7476 VGND 0.00639f
C30208 VPWR.n7477 VGND 0.00524f
C30209 VPWR.n7478 VGND 0.0066f
C30210 VPWR.n7479 VGND 0.00524f
C30211 VPWR.n7480 VGND 0.0066f
C30212 VPWR.n7481 VGND 0.00524f
C30213 VPWR.n7482 VGND 0.0066f
C30214 VPWR.n7483 VGND 0.00524f
C30215 VPWR.n7484 VGND 0.0066f
C30216 VPWR.n7485 VGND 0.00524f
C30217 VPWR.n7486 VGND 0.0066f
C30218 VPWR.n7487 VGND 0.00524f
C30219 VPWR.t3574 VGND 0.0592f
C30220 VPWR.n7488 VGND 0.0356f
C30221 VPWR.n7489 VGND 0.00484f
C30222 VPWR.n7490 VGND 0.00524f
C30223 VPWR.n7491 VGND 0.00506f
C30224 VPWR.n7492 VGND 0.00524f
C30225 VPWR.n7493 VGND 0.0066f
C30226 VPWR.n7494 VGND 0.00524f
C30227 VPWR.n7495 VGND 0.00639f
C30228 VPWR.n7496 VGND 0.00524f
C30229 VPWR.n7497 VGND 0.00393f
C30230 VPWR.n7498 VGND 0.00256f
C30231 VPWR.n7499 VGND 0.00515f
C30232 VPWR.n7500 VGND 0.0031f
C30233 VPWR.n7501 VGND 0.00524f
C30234 VPWR.n7502 VGND 0.00524f
C30235 VPWR.n7503 VGND 0.00393f
C30236 VPWR.n7504 VGND 0.00199f
C30237 VPWR.n7505 VGND 0.00173f
C30238 VPWR.n7506 VGND 0.00159f
C30239 VPWR.n7507 VGND 0.0031f
C30240 VPWR.n7508 VGND 0.00524f
C30241 VPWR.n7509 VGND 0.00121f
C30242 VPWR.n7510 VGND 0.00524f
C30243 VPWR.n7511 VGND 0.00393f
C30244 VPWR.n7512 VGND 0.00282f
C30245 VPWR.n7513 VGND 0.00993f
C30246 VPWR.n7514 VGND 0.00237f
C30247 VPWR.n7515 VGND 0.0031f
C30248 VPWR.n7516 VGND 0.00639f
C30249 VPWR.n7517 VGND 0.00524f
C30250 VPWR.n7518 VGND 0.0066f
C30251 VPWR.n7519 VGND 0.00524f
C30252 VPWR.n7520 VGND 0.0066f
C30253 VPWR.n7521 VGND 0.00524f
C30254 VPWR.n7522 VGND 0.0066f
C30255 VPWR.n7523 VGND 0.00524f
C30256 VPWR.n7524 VGND 0.0066f
C30257 VPWR.n7525 VGND 0.00524f
C30258 VPWR.n7526 VGND 0.00451f
C30259 VPWR.t642 VGND 0.00391f
C30260 VPWR.n7527 VGND 0.00833f
C30261 VPWR.t720 VGND 0.00391f
C30262 VPWR.n7528 VGND 0.00317f
C30263 VPWR.t719 VGND 0.00391f
C30264 VPWR.t3526 VGND 0.00886f
C30265 VPWR.n7529 VGND 0.0146f
C30266 VPWR.n7530 VGND 0.0116f
C30267 VPWR.n7531 VGND 0.0125f
C30268 VPWR.n7532 VGND 0.00475f
C30269 VPWR.n7533 VGND 0.00393f
C30270 VPWR.n7534 VGND 0.00503f
C30271 VPWR.t2380 VGND 0.00695f
C30272 VPWR.n7535 VGND 0.0084f
C30273 VPWR.n7536 VGND 0.00393f
C30274 VPWR.n7537 VGND 0.00122f
C30275 VPWR.n7538 VGND 0.00524f
C30276 VPWR.t2376 VGND 0.00166f
C30277 VPWR.t2378 VGND 0.00166f
C30278 VPWR.n7539 VGND 0.00345f
C30279 VPWR.n7540 VGND 0.00502f
C30280 VPWR.n7541 VGND 0.00524f
C30281 VPWR.n7542 VGND 0.00121f
C30282 VPWR.n7543 VGND 0.00524f
C30283 VPWR.t2374 VGND 0.00225f
C30284 VPWR.t743 VGND 0.00166f
C30285 VPWR.n7544 VGND 0.0045f
C30286 VPWR.n7545 VGND 0.00778f
C30287 VPWR.n7546 VGND 0.00524f
C30288 VPWR.n7547 VGND 0.0031f
C30289 VPWR.n7548 VGND 0.0016f
C30290 VPWR.n7549 VGND 0.00186f
C30291 VPWR.n7550 VGND 0.00393f
C30292 VPWR.n7551 VGND 0.00333f
C30293 VPWR.n7552 VGND 0.00157f
C30294 VPWR.t1489 VGND 0.00663f
C30295 VPWR.n7553 VGND 0.00913f
C30296 VPWR.n7554 VGND 0.00393f
C30297 VPWR.n7555 VGND 0.00121f
C30298 VPWR.n7556 VGND 0.00524f
C30299 VPWR.t1487 VGND -2.18e-20
C30300 VPWR.t940 VGND 0.00137f
C30301 VPWR.n7557 VGND 0.00629f
C30302 VPWR.n7558 VGND 0.0079f
C30303 VPWR.n7559 VGND 0.00524f
C30304 VPWR.t641 VGND 0.00391f
C30305 VPWR.t3497 VGND 0.00886f
C30306 VPWR.n7560 VGND 0.0116f
C30307 VPWR.n7561 VGND 0.0146f
C30308 VPWR.n7562 VGND 0.00317f
C30309 VPWR.n7563 VGND 0.00525f
C30310 VPWR.n7564 VGND 0.00146f
C30311 VPWR.n7565 VGND 0.0031f
C30312 VPWR.n7566 VGND 0.00393f
C30313 VPWR.n7567 VGND 0.00524f
C30314 VPWR.n7568 VGND 0.0031f
C30315 VPWR.n7569 VGND 0.00515f
C30316 VPWR.t143 VGND 0.0046f
C30317 VPWR.n7570 VGND 0.00407f
C30318 VPWR.n7571 VGND 0.00256f
C30319 VPWR.n7572 VGND 0.00393f
C30320 VPWR.n7573 VGND 0.00592f
C30321 VPWR.n7574 VGND 0.0039f
C30322 VPWR.n7575 VGND 0.00206f
C30323 VPWR.n7576 VGND 0.0033f
C30324 VPWR.n7577 VGND 0.00153f
C30325 VPWR.n7578 VGND 6.1e-19
C30326 VPWR.n7579 VGND 4.27e-19
C30327 VPWR.n7580 VGND 1.14e-19
C30328 VPWR.n7581 VGND 0.00326f
C30329 VPWR.n7582 VGND 4.27e-19
C30330 VPWR.n7583 VGND 6.83e-19
C30331 VPWR.n7584 VGND 3.7e-19
C30332 VPWR.n7585 VGND 9.68e-19
C30333 VPWR.n7586 VGND 9.96e-19
C30334 VPWR.n7587 VGND 5.41e-19
C30335 VPWR.n7588 VGND 7.4e-19
C30336 VPWR.n7589 VGND 6.1e-19
C30337 VPWR.n7590 VGND 0.00316f
C30338 VPWR.n7591 VGND 3.13e-19
C30339 VPWR.n7592 VGND 2.56e-19
C30340 VPWR.n7593 VGND 4.55e-19
C30341 VPWR.n7594 VGND 0.00176f
C30342 VPWR.n7595 VGND 9.68e-19
C30343 VPWR.n7596 VGND 9.96e-19
C30344 VPWR.n7597 VGND 3.13e-19
C30345 VPWR.n7598 VGND 4.84e-19
C30346 VPWR.n7599 VGND 6.83e-19
C30347 VPWR.t3580 VGND 0.0592f
C30348 VPWR.n7600 VGND 0.0345f
C30349 VPWR.n7601 VGND 0.00129f
C30350 VPWR.n7602 VGND 4.84e-19
C30351 VPWR.n7603 VGND 5.38e-19
C30352 VPWR.n7604 VGND 4.27e-19
C30353 VPWR.n7605 VGND 5.38e-19
C30354 VPWR.n7606 VGND 4.27e-19
C30355 VPWR.n7607 VGND 0.0033f
C30356 VPWR.n7608 VGND 9.6e-19
C30357 VPWR.n7609 VGND 0.00217f
C30358 VPWR.n7610 VGND 0.00138f
C30359 VPWR.n7611 VGND 3.07e-19
C30360 VPWR.n7612 VGND 5.48e-19
C30361 VPWR.n7614 VGND 0.1f
C30362 VPWR.n7615 VGND 0.1f
C30363 VPWR.n7616 VGND 6.54e-19
C30364 VPWR.n7617 VGND 8.67e-19
C30365 VPWR.n7618 VGND 4.39e-19
C30366 VPWR.n7619 VGND 3.29e-19
C30367 VPWR.n7620 VGND 5.27e-19
C30368 VPWR.n7621 VGND 2.85e-19
C30369 VPWR.n7622 VGND 2.85e-19
C30370 VPWR.n7623 VGND 4.17e-19
C30371 VPWR.n7624 VGND 5.71e-19
C30372 VPWR.n7625 VGND 4.17e-19
C30373 VPWR.n7626 VGND 3.51e-19
C30374 VPWR.n7627 VGND 4.61e-19
C30375 VPWR.n7628 VGND 4.17e-19
C30376 VPWR.n7629 VGND 4.11e-19
C30377 VPWR.n7630 VGND 7.39e-19
C30378 VPWR.n7631 VGND 5.19e-19
C30379 VPWR.n7632 VGND 7.39e-19
C30380 VPWR.n7633 VGND 4.11e-19
C30381 VPWR.n7634 VGND 4.11e-19
C30382 VPWR.t3347 VGND 0.0289f
C30383 VPWR.t76 VGND 0.00387f
C30384 VPWR.n7636 VGND 0.0547f
C30385 VPWR.t426 VGND 0.00462f
C30386 VPWR.n7637 VGND 0.0192f
C30387 VPWR.t3072 VGND 0.00631f
C30388 VPWR.n7638 VGND 0.00884f
C30389 VPWR.t3499 VGND 0.0592f
C30390 VPWR.t3070 VGND 0.00632f
C30391 VPWR.n7639 VGND 0.0066f
C30392 VPWR.t3338 VGND 0.00911f
C30393 VPWR.t17 VGND 0.00391f
C30394 VPWR.n7640 VGND 0.0253f
C30395 VPWR.t16 VGND 0.00391f
C30396 VPWR.n7642 VGND 0.0138f
C30397 VPWR.t3528 VGND 0.00911f
C30398 VPWR.t501 VGND 0.00391f
C30399 VPWR.n7643 VGND 0.0253f
C30400 VPWR.t502 VGND 0.00391f
C30401 VPWR.n7645 VGND 0.0138f
C30402 VPWR.n7646 VGND 0.0109f
C30403 VPWR.t2186 VGND 0.00682f
C30404 VPWR.t2182 VGND 0.00166f
C30405 VPWR.t2184 VGND 0.00166f
C30406 VPWR.n7647 VGND 0.00341f
C30407 VPWR.n7648 VGND 0.0101f
C30408 VPWR.n7649 VGND 0.00345f
C30409 VPWR.n7650 VGND 0.00444f
C30410 VPWR.t3360 VGND 0.00911f
C30411 VPWR.t1 VGND 0.00391f
C30412 VPWR.n7651 VGND 0.0253f
C30413 VPWR.t2 VGND 0.00391f
C30414 VPWR.n7653 VGND 0.0138f
C30415 VPWR.n7654 VGND 0.00762f
C30416 VPWR.t425 VGND 0.0046f
C30417 VPWR.n7655 VGND 0.00385f
C30418 VPWR.n7656 VGND 0.00233f
C30419 VPWR.n7657 VGND 0.00393f
C30420 VPWR.t2180 VGND 0.00225f
C30421 VPWR.t2015 VGND 0.00166f
C30422 VPWR.n7658 VGND 0.00438f
C30423 VPWR.n7659 VGND 0.0085f
C30424 VPWR.n7660 VGND 0.00352f
C30425 VPWR.n7661 VGND 0.00524f
C30426 VPWR.n7662 VGND 0.0031f
C30427 VPWR.n7663 VGND 0.00179f
C30428 VPWR.n7664 VGND 0.00337f
C30429 VPWR.n7665 VGND 0.00783f
C30430 VPWR.n7666 VGND 0.0355f
C30431 VPWR.n7667 VGND 0.0047f
C30432 VPWR.n7668 VGND 0.00475f
C30433 VPWR.n7669 VGND 0.00393f
C30434 VPWR.n7670 VGND 0.00344f
C30435 VPWR.n7671 VGND 0.0066f
C30436 VPWR.n7672 VGND 0.00393f
C30437 VPWR.n7673 VGND 0.00556f
C30438 VPWR.n7674 VGND 0.00333f
C30439 VPWR.n7675 VGND 0.00618f
C30440 VPWR.n7676 VGND 0.0119f
C30441 VPWR.n7677 VGND 0.0167f
C30442 VPWR.n7678 VGND 0.0107f
C30443 VPWR.t661 VGND 0.0046f
C30444 VPWR.n7679 VGND 0.01f
C30445 VPWR.n7680 VGND 0.0112f
C30446 VPWR.n7681 VGND 0.00475f
C30447 VPWR.n7682 VGND 0.00865f
C30448 VPWR.n7683 VGND 0.00171f
C30449 VPWR.n7684 VGND 0.00925f
C30450 VPWR.n7685 VGND 0.0166f
C30451 VPWR.n7686 VGND 0.0039f
C30452 VPWR.n7687 VGND 8.02e-19
C30453 VPWR.n7688 VGND 4.27e-19
C30454 VPWR.n7689 VGND 9.25e-19
C30455 VPWR.n7690 VGND 4.27e-19
C30456 VPWR.t3584 VGND 0.0612f
C30457 VPWR.n7691 VGND 0.0319f
C30458 VPWR.n7692 VGND 0.00225f
C30459 VPWR.n7693 VGND 4.84e-19
C30460 VPWR.n7694 VGND 6.83e-19
C30461 VPWR.n7695 VGND 4.84e-19
C30462 VPWR.n7696 VGND 1.99e-19
C30463 VPWR.n7697 VGND 4.83e-19
C30464 VPWR.n7698 VGND 4.61e-19
C30465 VPWR.n7699 VGND 6.54e-19
C30466 VPWR.n7700 VGND 8.67e-19
C30467 VPWR.n7701 VGND 4.11e-19
C30468 VPWR.n7702 VGND 4.61e-19
C30469 VPWR.n7703 VGND 2.41e-19
C30470 VPWR.n7704 VGND 4.83e-19
C30471 VPWR.n7705 VGND 8.26e-19
C30472 VPWR.n7706 VGND 0.0049f
C30473 VPWR.n7707 VGND 2.56e-19
C30474 VPWR.n7708 VGND 4.55e-19
C30475 VPWR.n7709 VGND 2.56e-19
C30476 VPWR.t77 VGND 0.00387f
C30477 VPWR.n7710 VGND 0.0102f
C30478 VPWR.n7711 VGND 0.00171f
C30479 VPWR.n7712 VGND 6.03e-19
C30480 VPWR.n7713 VGND 3.13e-19
C30481 VPWR.n7714 VGND 7.4e-19
C30482 VPWR.n7715 VGND 5.41e-19
C30483 VPWR.n7716 VGND 9.96e-19
C30484 VPWR.n7717 VGND 9.68e-19
C30485 VPWR.n7718 VGND 3.7e-19
C30486 VPWR.n7719 VGND 6.83e-19
C30487 VPWR.n7720 VGND 4.27e-19
C30488 VPWR.n7721 VGND 1.14e-19
C30489 VPWR.n7722 VGND 4.27e-19
C30490 VPWR.n7723 VGND 0.00153f
C30491 VPWR.n7724 VGND 0.00206f
C30492 VPWR.n7725 VGND 0.00138f
C30493 VPWR.n7726 VGND 9e-19
C30494 VPWR.n7727 VGND 6.14e-19
C30495 VPWR.n7728 VGND 9.06e-19
C30496 VPWR.n7729 VGND 5.48e-19
C30497 VPWR.n7730 VGND 0.00138f
C30498 VPWR.n7731 VGND 0.0057f
C30499 VPWR.n7733 VGND 0.00139f
C30500 VPWR.n7734 VGND 5.48e-19
C30501 VPWR.n7735 VGND 3.07e-19
C30502 VPWR.n7736 VGND 0.00138f
C30503 VPWR.n7737 VGND 0.00217f
C30504 VPWR.n7738 VGND 0.0109f
C30505 VPWR.n7739 VGND 0.00451f
C30506 VPWR.n7740 VGND 0.0113f
C30507 VPWR.n7741 VGND 0.00524f
C30508 VPWR.n7742 VGND 0.0087f
C30509 VPWR.n7743 VGND 0.00524f
C30510 VPWR.t3427 VGND 0.0592f
C30511 VPWR.n7744 VGND 0.038f
C30512 VPWR.n7745 VGND 0.00833f
C30513 VPWR.n7746 VGND 0.00524f
C30514 VPWR.n7747 VGND 0.0113f
C30515 VPWR.n7748 VGND 0.00524f
C30516 VPWR.n7749 VGND 0.011f
C30517 VPWR.n7750 VGND 0.00524f
C30518 VPWR.t662 VGND 0.0046f
C30519 VPWR.n7751 VGND 0.00644f
C30520 VPWR.n7752 VGND 0.00535f
C30521 VPWR.n7753 VGND 0.0031f
C30522 VPWR.n7754 VGND 0.00282f
C30523 VPWR.n7755 VGND 0.00199f
C30524 VPWR.n7756 VGND 0.00556f
C30525 VPWR.t308 VGND 0.00462f
C30526 VPWR.n7757 VGND 0.0103f
C30527 VPWR.t3463 VGND 0.0111f
C30528 VPWR.n7758 VGND 0.0205f
C30529 VPWR.t310 VGND 0.00387f
C30530 VPWR.n7759 VGND 0.0163f
C30531 VPWR.n7760 VGND 0.0115f
C30532 VPWR.n7761 VGND 0.00719f
C30533 VPWR.t311 VGND 0.00387f
C30534 VPWR.n7762 VGND 0.0186f
C30535 VPWR.n7763 VGND 0.0132f
C30536 VPWR.n7764 VGND 0.00638f
C30537 VPWR.n7765 VGND 0.00793f
C30538 VPWR.n7766 VGND 0.00529f
C30539 VPWR.n7767 VGND 0.00279f
C30540 VPWR.n7768 VGND 0.00723f
C30541 VPWR.n7769 VGND 0.00393f
C30542 VPWR.n7770 VGND 0.00524f
C30543 VPWR.n7771 VGND 0.0113f
C30544 VPWR.n7772 VGND 0.00524f
C30545 VPWR.n7773 VGND 0.0087f
C30546 VPWR.n7774 VGND 0.00524f
C30547 VPWR.t3540 VGND 0.0592f
C30548 VPWR.n7775 VGND 0.038f
C30549 VPWR.n7776 VGND 0.00833f
C30550 VPWR.n7777 VGND 0.00524f
C30551 VPWR.n7778 VGND 0.0113f
C30552 VPWR.n7779 VGND 0.00524f
C30553 VPWR.n7780 VGND 0.00524f
C30554 VPWR.n7781 VGND 0.0031f
C30555 VPWR.n7782 VGND 0.00516f
C30556 VPWR.t211 VGND 0.0046f
C30557 VPWR.n7783 VGND 0.00644f
C30558 VPWR.n7784 VGND 0.00512f
C30559 VPWR.n7785 VGND 0.00475f
C30560 VPWR.n7786 VGND 0.011f
C30561 VPWR.n7787 VGND 0.00524f
C30562 VPWR.n7788 VGND 0.00524f
C30563 VPWR.n7789 VGND 0.0031f
C30564 VPWR.n7790 VGND 0.00285f
C30565 VPWR.n7791 VGND 0.0351f
C30566 VPWR.t713 VGND 0.0046f
C30567 VPWR.n7792 VGND 0.00644f
C30568 VPWR.n7793 VGND 0.00255f
C30569 VPWR.n7794 VGND 0.00475f
C30570 VPWR.n7795 VGND 0.011f
C30571 VPWR.n7796 VGND 0.00524f
C30572 VPWR.n7797 VGND 0.0113f
C30573 VPWR.n7798 VGND 0.00524f
C30574 VPWR.n7799 VGND 0.0087f
C30575 VPWR.n7800 VGND 0.00524f
C30576 VPWR.t3341 VGND 0.0592f
C30577 VPWR.n7801 VGND 0.038f
C30578 VPWR.n7802 VGND 0.00833f
C30579 VPWR.n7803 VGND 0.00524f
C30580 VPWR.n7804 VGND 0.0113f
C30581 VPWR.n7805 VGND 0.00524f
C30582 VPWR.n7806 VGND 0.00524f
C30583 VPWR.n7807 VGND 0.0031f
C30584 VPWR.n7808 VGND 0.00282f
C30585 VPWR.n7809 VGND 0.0143f
C30586 VPWR.t632 VGND 0.0046f
C30587 VPWR.n7810 VGND 0.00644f
C30588 VPWR.n7811 VGND 0.0053f
C30589 VPWR.n7812 VGND 0.00393f
C30590 VPWR.n7813 VGND 0.00524f
C30591 VPWR.n7814 VGND 0.0031f
C30592 VPWR.n7815 VGND 0.00478f
C30593 VPWR.n7816 VGND 0.00452f
C30594 VPWR.n7817 VGND 0.00211f
C30595 VPWR.n7818 VGND 2.85e-19
C30596 VPWR.n7819 VGND 9.87e-19
C30597 VPWR.n7820 VGND 2.28e-19
C30598 VPWR.t31 VGND 0.0046f
C30599 VPWR.n7821 VGND 0.0012f
C30600 VPWR.n7822 VGND 0.00265f
C30601 VPWR.n7823 VGND 6.26e-19
C30602 VPWR.n7824 VGND 5.12e-19
C30603 VPWR.n7825 VGND 3.13e-19
C30604 VPWR.n7826 VGND 0.00122f
C30605 VPWR.n7827 VGND 0.00108f
C30606 VPWR.n7828 VGND 5.12e-19
C30607 VPWR.n7829 VGND 5.98e-19
C30608 VPWR.t3536 VGND 0.0592f
C30609 VPWR.n7830 VGND 0.0376f
C30610 VPWR.n7831 VGND 0.00759f
C30611 VPWR.n7832 VGND 3.13e-19
C30612 VPWR.n7833 VGND 5.41e-19
C30613 VPWR.n7834 VGND 9.68e-19
C30614 VPWR.n7835 VGND 9.96e-19
C30615 VPWR.n7836 VGND 5.41e-19
C30616 VPWR.n7837 VGND 6.55e-19
C30617 VPWR.n7838 VGND 6.26e-19
C30618 VPWR.n7839 VGND 0.00555f
C30619 VPWR.n7840 VGND 3.7e-19
C30620 VPWR.n7841 VGND 7.4e-19
C30621 VPWR.n7842 VGND 3.42e-19
C30622 VPWR.n7843 VGND 8.02e-19
C30623 VPWR.n7844 VGND 3.7e-19
C30624 VPWR.n7845 VGND 0.00567f
C30625 VPWR.n7846 VGND 5.41e-19
C30626 VPWR.n7847 VGND 5.41e-19
C30627 VPWR.n7848 VGND 5.12e-19
C30628 VPWR.n7849 VGND 4.27e-19
C30629 VPWR.n7850 VGND 9.96e-19
C30630 VPWR.n7851 VGND 0.00131f
C30631 VPWR.n7852 VGND 5.69e-19
C30632 VPWR.n7853 VGND 0.00802f
C30633 VPWR.n7854 VGND 6.8e-19
C30634 VPWR.n7855 VGND 0.00218f
C30635 VPWR.n7856 VGND 0.00137f
C30636 VPWR.n7857 VGND 4.17e-19
C30637 VPWR.n7858 VGND 5.48e-19
C30638 VPWR.n7860 VGND 0.0452f
C30639 VPWR.n7861 VGND 0.0976f
C30640 VPWR.n7862 VGND 0.0581f
C30641 VPWR.n7864 VGND 4.83e-19
C30642 VPWR.n7865 VGND 2.85e-19
C30643 VPWR.n7866 VGND 3.95e-19
C30644 VPWR.n7867 VGND 3.95e-19
C30645 VPWR.n7868 VGND 3.7e-19
C30646 VPWR.n7869 VGND 3.42e-19
C30647 VPWR.n7870 VGND 3.7e-19
C30648 VPWR.n7871 VGND 4.84e-19
C30649 VPWR.n7872 VGND 8.54e-20
C30650 VPWR.n7873 VGND 3.29e-19
C30651 VPWR.n7874 VGND 5.71e-19
C30652 VPWR.n7875 VGND 5.92e-19
C30653 VPWR.n7876 VGND 5.05e-19
C30654 VPWR.n7877 VGND 8.67e-19
C30655 VPWR.n7878 VGND 6.54e-19
C30656 VPWR.n7879 VGND 9.06e-19
C30657 VPWR.n7880 VGND 0.1f
C30658 VPWR.n7881 VGND 0.1f
C30659 VPWR.n7882 VGND 0.00139f
C30660 VPWR.n7883 VGND 9.06e-19
C30661 VPWR.n7884 VGND 8.11e-19
C30662 VPWR.n7885 VGND 3.95e-19
C30663 VPWR.n7886 VGND 1.76e-19
C30664 VPWR.n7887 VGND 3.95e-19
C30665 VPWR.n7888 VGND 7.68e-19
C30666 VPWR.n7889 VGND 5.05e-19
C30667 VPWR.n7890 VGND 1.76e-19
C30668 VPWR.n7891 VGND 5.48e-19
C30669 VPWR.n7893 VGND 0.0057f
C30670 VPWR.n7894 VGND 0.00138f
C30671 VPWR.n7895 VGND 5.48e-19
C30672 VPWR.n7896 VGND 4.17e-19
C30673 VPWR.n7897 VGND 6.55e-19
C30674 VPWR.n7898 VGND 6.26e-19
C30675 VPWR.n7899 VGND 0.00688f
C30676 VPWR.n7900 VGND 0.0125f
C30677 VPWR.t536 VGND 0.00387f
C30678 VPWR.n7901 VGND 0.00837f
C30679 VPWR.t2807 VGND 0.00676f
C30680 VPWR.t4 VGND 0.0046f
C30681 VPWR.n7902 VGND 0.00407f
C30682 VPWR.t5 VGND 0.0046f
C30683 VPWR.n7903 VGND 0.00407f
C30684 VPWR.t3260 VGND 0.00692f
C30685 VPWR.n7904 VGND 0.0109f
C30686 VPWR.t2847 VGND 6.73e-19
C30687 VPWR.t3258 VGND 0.00127f
C30688 VPWR.n7905 VGND 0.00207f
C30689 VPWR.n7906 VGND 0.00464f
C30690 VPWR.t946 VGND 0.00102f
C30691 VPWR.t2092 VGND 0.00102f
C30692 VPWR.n7907 VGND 0.00221f
C30693 VPWR.n7908 VGND 0.00589f
C30694 VPWR.n7909 VGND 0.00121f
C30695 VPWR.n7910 VGND 0.0031f
C30696 VPWR.n7911 VGND 0.00524f
C30697 VPWR.n7912 VGND 0.00524f
C30698 VPWR.n7913 VGND 0.00138f
C30699 VPWR.n7914 VGND 0.00524f
C30700 VPWR.t1993 VGND 0.00234f
C30701 VPWR.t1995 VGND 0.00239f
C30702 VPWR.n7915 VGND 0.00401f
C30703 VPWR.n7916 VGND 0.00333f
C30704 VPWR.n7917 VGND 8.57e-19
C30705 VPWR.n7918 VGND 0.00524f
C30706 VPWR.n7919 VGND 0.00524f
C30707 VPWR.n7920 VGND 0.00475f
C30708 VPWR.n7921 VGND 0.0014f
C30709 VPWR.n7922 VGND 0.00274f
C30710 VPWR.n7923 VGND 0.0031f
C30711 VPWR.n7924 VGND 0.00484f
C30712 VPWR.n7925 VGND 0.00524f
C30713 VPWR.t1706 VGND 6.73e-19
C30714 VPWR.t2981 VGND 9.96e-19
C30715 VPWR.n7926 VGND 0.00176f
C30716 VPWR.n7927 VGND 0.00658f
C30717 VPWR.n7928 VGND 0.00484f
C30718 VPWR.n7929 VGND 0.00524f
C30719 VPWR.n7930 VGND 0.00553f
C30720 VPWR.n7931 VGND 0.00524f
C30721 VPWR.t775 VGND 0.00453f
C30722 VPWR.n7932 VGND 0.00799f
C30723 VPWR.n7933 VGND 0.00438f
C30724 VPWR.n7934 VGND 0.00524f
C30725 VPWR.n7935 VGND 0.0066f
C30726 VPWR.n7936 VGND 0.00524f
C30727 VPWR.n7937 VGND 0.0066f
C30728 VPWR.n7938 VGND 0.00524f
C30729 VPWR.t3344 VGND 0.0592f
C30730 VPWR.n7939 VGND 0.0351f
C30731 VPWR.n7940 VGND 0.00484f
C30732 VPWR.n7941 VGND 0.00524f
C30733 VPWR.t1710 VGND 6.73e-19
C30734 VPWR.t2805 VGND 0.00127f
C30735 VPWR.n7942 VGND 0.00203f
C30736 VPWR.n7943 VGND 0.0044f
C30737 VPWR.n7944 VGND 0.00377f
C30738 VPWR.n7945 VGND 0.00524f
C30739 VPWR.n7946 VGND 0.00535f
C30740 VPWR.n7947 VGND 0.00524f
C30741 VPWR.t2983 VGND 0.00239f
C30742 VPWR.n7948 VGND 0.00658f
C30743 VPWR.n7949 VGND 0.00434f
C30744 VPWR.n7950 VGND 0.00524f
C30745 VPWR.n7951 VGND 0.00393f
C30746 VPWR.n7952 VGND 0.00194f
C30747 VPWR.n7953 VGND 0.00927f
C30748 VPWR.n7954 VGND 0.00513f
C30749 VPWR.n7955 VGND 0.00179f
C30750 VPWR.n7956 VGND 6.26e-19
C30751 VPWR.n7957 VGND 6.8e-19
C30752 VPWR.n7958 VGND 5.05e-19
C30753 VPWR.n7959 VGND 6.58e-20
C30754 VPWR.n7960 VGND 1.33e-19
C30755 VPWR.n7961 VGND 5.69e-19
C30756 VPWR.n7962 VGND 0.00128f
C30757 VPWR.n7963 VGND 2.56e-19
C30758 VPWR.n7964 VGND 4.27e-19
C30759 VPWR.n7965 VGND 5.12e-19
C30760 VPWR.n7966 VGND 3.7e-19
C30761 VPWR.n7967 VGND 4.17e-19
C30762 VPWR.n7968 VGND 2.85e-19
C30763 VPWR.n7969 VGND 2.85e-19
C30764 VPWR.n7970 VGND 4.11e-19
C30765 VPWR.n7971 VGND 4.11e-19
C30766 VPWR.n7972 VGND 7.39e-19
C30767 VPWR.n7973 VGND 5.19e-19
C30768 VPWR.n7974 VGND 7.39e-19
C30769 VPWR.n7975 VGND 4.11e-19
C30770 VPWR.n7976 VGND 4.11e-19
C30771 VPWR.n7977 VGND 3.07e-19
C30772 VPWR.n7978 VGND 1.76e-19
C30773 VPWR.n7979 VGND 4.39e-19
C30774 VPWR.n7980 VGND 6.14e-19
C30775 VPWR.n7981 VGND 4.17e-19
C30776 VPWR.n7982 VGND 5.05e-19
C30777 VPWR.n7983 VGND 6.55e-19
C30778 VPWR.n7984 VGND 5.41e-19
C30779 VPWR.n7985 VGND 9.96e-19
C30780 VPWR.n7986 VGND 9.68e-19
C30781 VPWR.n7987 VGND 5.41e-19
C30782 VPWR.t1297 VGND 0.00136f
C30783 VPWR.t1865 VGND 0.00136f
C30784 VPWR.n7988 VGND 0.00317f
C30785 VPWR.t535 VGND 0.00389f
C30786 VPWR.t3519 VGND 0.029f
C30787 VPWR.n7989 VGND 0.0437f
C30788 VPWR.n7990 VGND 0.0123f
C30789 VPWR.n7991 VGND 0.0206f
C30790 VPWR.n7992 VGND 0.00899f
C30791 VPWR.n7993 VGND 9.71e-19
C30792 VPWR.n7994 VGND 8.97e-19
C30793 VPWR.n7995 VGND 0.00673f
C30794 VPWR.n7996 VGND 0.0159f
C30795 VPWR.n7997 VGND 3.13e-19
C30796 VPWR.n7998 VGND 5.98e-19
C30797 VPWR.n7999 VGND 5.12e-19
C30798 VPWR.n8000 VGND 0.00108f
C30799 VPWR.n8001 VGND 0.00122f
C30800 VPWR.n8002 VGND 3.13e-19
C30801 VPWR.n8003 VGND 5.12e-19
C30802 VPWR.n8004 VGND 6.26e-19
C30803 VPWR.n8005 VGND 0.00407f
C30804 VPWR.n8006 VGND 4.61e-20
C30805 VPWR.n8007 VGND 4.67e-19
C30806 VPWR.n8008 VGND 0.00211f
C30807 VPWR.n8009 VGND 0.00442f
C30808 VPWR.n8010 VGND 0.00282f
C30809 VPWR.n8011 VGND 0.0134f
C30810 VPWR.n8012 VGND 0.0653f
C30811 VPWR.t534 VGND 0.0206f
C30812 VPWR.t1296 VGND 0.0151f
C30813 VPWR.t1864 VGND 0.0257f
C30814 VPWR.t2806 VGND 0.0413f
C30815 VPWR.t2982 VGND 0.0502f
C30816 VPWR.t1709 VGND 0.0322f
C30817 VPWR.t2804 VGND 0.0322f
C30818 VPWR.t2879 VGND 0.024f
C30819 VPWR.t3 VGND 0.0144f
C30820 VPWR.t944 VGND 0.0211f
C30821 VPWR.t774 VGND 0.0497f
C30822 VPWR.t1705 VGND 0.0493f
C30823 VPWR.t2980 VGND 0.0336f
C30824 VPWR.t943 VGND 0.0206f
C30825 VPWR.t3259 VGND 0.0166f
C30826 VPWR.t2880 VGND 0.0176f
C30827 VPWR.t1992 VGND 0.0339f
C30828 VPWR.t1994 VGND 0.0326f
C30829 VPWR.t2846 VGND 0.0264f
C30830 VPWR.t945 VGND 0.0181f
C30831 VPWR.t3257 VGND 0.0141f
C30832 VPWR.t2091 VGND 0.0141f
C30833 VPWR.t2672 VGND 0.0109f
C30834 VPWR.t2571 VGND 0.0126f
C30835 VPWR.t361 VGND 0.0415f
C30836 VPWR.t574 VGND 0.0666f
C30837 VPWR.t2498 VGND 0.025f
C30838 VPWR.t1551 VGND 0.02f
C30839 VPWR.t2679 VGND 0.025f
C30840 VPWR.t1549 VGND 0.0144f
C30841 VPWR.t1350 VGND 0.0161f
C30842 VPWR.t1848 VGND 0.0309f
C30843 VPWR.t2496 VGND 0.0154f
C30844 VPWR.t782 VGND 0.0158f
C30845 VPWR.t1846 VGND 0.0205f
C30846 VPWR.t1990 VGND 0.0311f
C30847 VPWR.t2089 VGND 0.025f
C30848 VPWR.t2572 VGND 0.0589f
C30849 VPWR.t2079 VGND 0.0603f
C30850 VPWR.t2673 VGND 0.018f
C30851 VPWR.t166 VGND 0.0166f
C30852 VPWR.t2570 VGND 0.0376f
C30853 VPWR.t1389 VGND 0.0398f
C30854 VPWR.t2842 VGND 0.0493f
C30855 VPWR.t2313 VGND 0.0465f
C30856 VPWR.n8013 VGND 0.0204f
C30857 VPWR.n8014 VGND 0.0102f
C30858 VPWR.t167 VGND 0.0046f
C30859 VPWR.t2314 VGND 0.00453f
C30860 VPWR.n8015 VGND 0.00778f
C30861 VPWR.n8016 VGND 0.00184f
C30862 VPWR.n8017 VGND 0.00233f
C30863 VPWR.n8018 VGND 0.00393f
C30864 VPWR.n8019 VGND 0.00553f
C30865 VPWR.n8020 VGND 0.00524f
C30866 VPWR.t2843 VGND 6.73e-19
C30867 VPWR.t1390 VGND 9.96e-19
C30868 VPWR.n8021 VGND 0.00176f
C30869 VPWR.n8022 VGND 0.00658f
C30870 VPWR.n8023 VGND 0.00484f
C30871 VPWR.n8024 VGND 0.00524f
C30872 VPWR.n8025 VGND 0.00352f
C30873 VPWR.n8026 VGND 0.00524f
C30874 VPWR.t3404 VGND 0.0592f
C30875 VPWR.n8027 VGND 0.0356f
C30876 VPWR.n8028 VGND 0.00484f
C30877 VPWR.n8029 VGND 0.00524f
C30878 VPWR.n8030 VGND 0.0066f
C30879 VPWR.n8031 VGND 0.00524f
C30880 VPWR.n8032 VGND 0.0066f
C30881 VPWR.n8033 VGND 0.00524f
C30882 VPWR.t2080 VGND 0.00234f
C30883 VPWR.n8034 VGND 0.00628f
C30884 VPWR.n8035 VGND 0.00398f
C30885 VPWR.n8036 VGND 0.00524f
C30886 VPWR.n8037 VGND 0.00592f
C30887 VPWR.n8038 VGND 0.00524f
C30888 VPWR.n8039 VGND 0.0066f
C30889 VPWR.n8040 VGND 0.00524f
C30890 VPWR.n8041 VGND 0.00337f
C30891 VPWR.n8042 VGND 0.00524f
C30892 VPWR.n8043 VGND 0.0031f
C30893 VPWR.n8044 VGND 0.00274f
C30894 VPWR.n8045 VGND 0.0014f
C30895 VPWR.n8046 VGND 0.00393f
C30896 VPWR.n8047 VGND 0.00333f
C30897 VPWR.t1991 VGND 0.0016f
C30898 VPWR.t1847 VGND 0.00208f
C30899 VPWR.n8048 VGND 0.00422f
C30900 VPWR.n8049 VGND 0.00644f
C30901 VPWR.n8050 VGND 0.00135f
C30902 VPWR.n8051 VGND 0.00393f
C30903 VPWR.t783 VGND 0.0016f
C30904 VPWR.t1849 VGND 0.00208f
C30905 VPWR.n8052 VGND 0.00419f
C30906 VPWR.t2497 VGND 0.00527f
C30907 VPWR.n8053 VGND 0.0106f
C30908 VPWR.n8054 VGND 0.00524f
C30909 VPWR.n8055 VGND 0.00114f
C30910 VPWR.n8056 VGND 0.00524f
C30911 VPWR.t1351 VGND 0.00527f
C30912 VPWR.n8057 VGND 0.0065f
C30913 VPWR.n8058 VGND 0.00504f
C30914 VPWR.n8059 VGND 0.00218f
C30915 VPWR.n8060 VGND 0.0013f
C30916 VPWR.n8061 VGND 6.99e-19
C30917 VPWR.n8062 VGND 4.84e-19
C30918 VPWR.n8063 VGND 0.00309f
C30919 VPWR.n8064 VGND 3.7e-19
C30920 VPWR.t362 VGND 0.0046f
C30921 VPWR.n8065 VGND 0.00113f
C30922 VPWR.n8066 VGND 2.15e-19
C30923 VPWR.n8067 VGND 3.7e-19
C30924 VPWR.n8068 VGND 4.66e-19
C30925 VPWR.n8069 VGND 3.7e-19
C30926 VPWR.n8070 VGND 0.0022f
C30927 VPWR.n8071 VGND 5.12e-19
C30928 VPWR.n8072 VGND 5.41e-19
C30929 VPWR.n8073 VGND 5.12e-19
C30930 VPWR.n8074 VGND 4.27e-19
C30931 VPWR.n8075 VGND 2.85e-19
C30932 VPWR.n8076 VGND 8.26e-19
C30933 VPWR.n8077 VGND 5.05e-19
C30934 VPWR.n8078 VGND 4.17e-19
C30935 VPWR.n8079 VGND 5.48e-19
C30936 VPWR.n8081 VGND 0.1f
C30937 VPWR.n8082 VGND 0.1f
C30938 VPWR.n8083 VGND 0.1f
C30939 VPWR.n8084 VGND 0.1f
C30940 VPWR.n8085 VGND 0.00139f
C30941 VPWR.n8086 VGND 9.06e-19
C30942 VPWR.n8087 VGND 5.92e-19
C30943 VPWR.n8088 VGND 5.05e-19
C30944 VPWR.n8089 VGND 4.17e-19
C30945 VPWR.n8090 VGND 5.48e-19
C30946 VPWR.n8092 VGND 8.67e-19
C30947 VPWR.n8093 VGND 6.54e-19
C30948 VPWR.n8094 VGND 9.06e-19
C30949 VPWR.n8095 VGND 3.95e-19
C30950 VPWR.n8096 VGND 3.95e-19
C30951 VPWR.n8097 VGND 7.68e-19
C30952 VPWR.n8098 VGND 5.05e-19
C30953 VPWR.n8099 VGND 8.11e-19
C30954 VPWR.n8100 VGND 3.95e-19
C30955 VPWR.n8101 VGND 9.68e-19
C30956 VPWR.n8102 VGND 5.12e-19
C30957 VPWR.n8103 VGND 0.00105f
C30958 VPWR.n8104 VGND 3.13e-19
C30959 VPWR.n8105 VGND 5.12e-19
C30960 VPWR.n8106 VGND 1.99e-19
C30961 VPWR.n8107 VGND 0.00108f
C30962 VPWR.n8108 VGND 0.00122f
C30963 VPWR.t882 VGND 0.00654f
C30964 VPWR.n8109 VGND 0.0107f
C30965 VPWR.t372 VGND 0.00387f
C30966 VPWR.n8110 VGND 0.00613f
C30967 VPWR.n8111 VGND 0.00199f
C30968 VPWR.t2845 VGND 6.73e-19
C30969 VPWR.t1130 VGND 9.96e-19
C30970 VPWR.n8112 VGND 0.00176f
C30971 VPWR.n8113 VGND 0.00421f
C30972 VPWR.t2550 VGND 0.018f
C30973 VPWR.t2809 VGND 0.0252f
C30974 VPWR.t2486 VGND 0.0253f
C30975 VPWR.t498 VGND 0.0166f
C30976 VPWR.t2393 VGND 0.026f
C30977 VPWR.t2832 VGND 0.029f
C30978 VPWR.t2206 VGND 0.0398f
C30979 VPWR.t2487 VGND 0.0401f
C30980 VPWR.t2808 VGND 0.0321f
C30981 VPWR.t907 VGND 0.0284f
C30982 VPWR.t9 VGND 0.0448f
C30983 VPWR.t2488 VGND 0.046f
C30984 VPWR.t1831 VGND 0.025f
C30985 VPWR.t899 VGND 0.0203f
C30986 VPWR.t2682 VGND 0.0148f
C30987 VPWR.t1175 VGND 0.0149f
C30988 VPWR.t3113 VGND 0.0361f
C30989 VPWR.t1500 VGND 0.0267f
C30990 VPWR.t2368 VGND 0.0089f
C30991 VPWR.t2830 VGND 0.0121f
C30992 VPWR.t881 VGND 0.0181f
C30993 VPWR.t1177 VGND 0.024f
C30994 VPWR.t999 VGND 0.0285f
C30995 VPWR.t1932 VGND 0.0253f
C30996 VPWR.t370 VGND 0.0166f
C30997 VPWR.t824 VGND 0.026f
C30998 VPWR.t2157 VGND 0.00102f
C30999 VPWR.t2555 VGND 0.00154f
C31000 VPWR.n8114 VGND 0.00486f
C31001 VPWR.n8115 VGND 0.0117f
C31002 VPWR.n8116 VGND 0.0171f
C31003 VPWR.n8117 VGND 0.00121f
C31004 VPWR.t2752 VGND 6.73e-19
C31005 VPWR.t1354 VGND 9.96e-19
C31006 VPWR.n8118 VGND 0.00176f
C31007 VPWR.n8119 VGND 0.0101f
C31008 VPWR.n8120 VGND 0.0102f
C31009 VPWR.n8121 VGND 0.0101f
C31010 VPWR.t68 VGND 0.00387f
C31011 VPWR.n8122 VGND 0.00837f
C31012 VPWR.n8123 VGND 0.00525f
C31013 VPWR.t2298 VGND 0.00239f
C31014 VPWR.t1366 VGND 6.73e-19
C31015 VPWR.t2790 VGND 0.00127f
C31016 VPWR.n8124 VGND 0.00204f
C31017 VPWR.n8125 VGND 0.00705f
C31018 VPWR.t1935 VGND 0.00102f
C31019 VPWR.t2086 VGND 0.00102f
C31020 VPWR.n8126 VGND 0.00221f
C31021 VPWR.n8127 VGND 0.00179f
C31022 VPWR.n8128 VGND 0.00142f
C31023 VPWR.n8129 VGND 0.00186f
C31024 VPWR.n8130 VGND 0.00475f
C31025 VPWR.n8131 VGND 0.00149f
C31026 VPWR.n8132 VGND 0.00524f
C31027 VPWR.t2685 VGND 0.00527f
C31028 VPWR.n8133 VGND 0.00644f
C31029 VPWR.n8134 VGND 0.00524f
C31030 VPWR.t2922 VGND 0.00238f
C31031 VPWR.n8135 VGND 0.0048f
C31032 VPWR.n8136 VGND 0.00524f
C31033 VPWR.t1851 VGND 0.00208f
C31034 VPWR.t2205 VGND 0.0016f
C31035 VPWR.n8137 VGND 0.00422f
C31036 VPWR.n8138 VGND 0.006f
C31037 VPWR.n8139 VGND 0.00524f
C31038 VPWR.n8140 VGND 0.00393f
C31039 VPWR.n8141 VGND 0.00119f
C31040 VPWR.n8142 VGND 0.00592f
C31041 VPWR.n8143 VGND 0.00393f
C31042 VPWR.n8144 VGND 0.0031f
C31043 VPWR.n8145 VGND 0.00444f
C31044 VPWR.t3543 VGND 0.00911f
C31045 VPWR.t7 VGND 0.00391f
C31046 VPWR.n8146 VGND 0.0253f
C31047 VPWR.t8 VGND 0.00391f
C31048 VPWR.n8148 VGND 0.0138f
C31049 VPWR.t2792 VGND 0.00692f
C31050 VPWR.n8149 VGND 0.0103f
C31051 VPWR.n8150 VGND 0.00789f
C31052 VPWR.t67 VGND 0.00387f
C31053 VPWR.n8151 VGND 0.00837f
C31054 VPWR.n8152 VGND 0.00471f
C31055 VPWR.n8153 VGND 0.00393f
C31056 VPWR.n8154 VGND 0.01f
C31057 VPWR.n8155 VGND 0.00524f
C31058 VPWR.t3556 VGND 0.0282f
C31059 VPWR.n8156 VGND 0.0489f
C31060 VPWR.n8157 VGND 0.0102f
C31061 VPWR.n8158 VGND 0.00524f
C31062 VPWR.t2960 VGND 0.00453f
C31063 VPWR.n8159 VGND 0.0116f
C31064 VPWR.n8160 VGND 0.00912f
C31065 VPWR.n8161 VGND 0.00524f
C31066 VPWR.n8162 VGND 0.0115f
C31067 VPWR.n8163 VGND 0.00524f
C31068 VPWR.n8164 VGND 0.00524f
C31069 VPWR.n8165 VGND 0.00524f
C31070 VPWR.n8166 VGND 0.0031f
C31071 VPWR.n8167 VGND 0.00179f
C31072 VPWR.n8168 VGND 0.00173f
C31073 VPWR.n8169 VGND 0.00179f
C31074 VPWR.n8170 VGND 0.00475f
C31075 VPWR.t1607 VGND 0.00238f
C31076 VPWR.n8171 VGND 0.00494f
C31077 VPWR.n8172 VGND 0.00524f
C31078 VPWR.t2160 VGND 0.00527f
C31079 VPWR.n8173 VGND 0.00606f
C31080 VPWR.n8174 VGND 0.00524f
C31081 VPWR.n8175 VGND 0.00119f
C31082 VPWR.n8176 VGND 0.00524f
C31083 VPWR.t1009 VGND 0.00102f
C31084 VPWR.t1834 VGND 0.00102f
C31085 VPWR.n8177 VGND 0.00221f
C31086 VPWR.t2429 VGND 0.00208f
C31087 VPWR.t2933 VGND 0.0016f
C31088 VPWR.n8178 VGND 0.00419f
C31089 VPWR.n8179 VGND 0.0104f
C31090 VPWR.n8180 VGND 0.00524f
C31091 VPWR.n8181 VGND 0.0031f
C31092 VPWR.n8182 VGND 0.00622f
C31093 VPWR.n8183 VGND 0.00199f
C31094 VPWR.n8184 VGND 0.00994f
C31095 VPWR.t196 VGND 0.0463f
C31096 VPWR.t1825 VGND 0.0111f
C31097 VPWR.t2480 VGND 0.0141f
C31098 VPWR.t2113 VGND 0.0141f
C31099 VPWR.t2482 VGND 0.0161f
C31100 VPWR.t3129 VGND 0.0211f
C31101 VPWR.t2893 VGND 0.0237f
C31102 VPWR.t3181 VGND 0.0321f
C31103 VPWR.t2112 VGND 0.021f
C31104 VPWR.t889 VGND 0.0164f
C31105 VPWR.t3275 VGND 0.0171f
C31106 VPWR.t840 VGND 0.0156f
C31107 VPWR.t1367 VGND 0.026f
C31108 VPWR.t409 VGND 0.0331f
C31109 VPWR.t2814 VGND 0.0264f
C31110 VPWR.t2115 VGND 0.026f
C31111 VPWR.t3180 VGND 0.0116f
C31112 VPWR.t3132 VGND 0.0141f
C31113 VPWR.t2856 VGND 0.0144f
C31114 VPWR.t2161 VGND 0.0181f
C31115 VPWR.t2753 VGND 0.0149f
C31116 VPWR.t3103 VGND 0.0141f
C31117 VPWR.t2568 VGND 0.0208f
C31118 VPWR.t2858 VGND 0.0467f
C31119 VPWR.t560 VGND 0.0151f
C31120 VPWR.t3131 VGND 0.0299f
C31121 VPWR.t2156 VGND 0.0284f
C31122 VPWR.t2554 VGND 0.0347f
C31123 VPWR.n8185 VGND 0.0348f
C31124 VPWR.t1833 VGND 0.025f
C31125 VPWR.t1008 VGND 0.0154f
C31126 VPWR.t2428 VGND 0.0171f
C31127 VPWR.t2159 VGND 0.0435f
C31128 VPWR.t1606 VGND 0.0312f
C31129 VPWR.t1550 VGND 0.0154f
C31130 VPWR.t1970 VGND 0.0141f
C31131 VPWR.t3190 VGND 0.00739f
C31132 VPWR.t1006 VGND 0.0154f
C31133 VPWR.t1353 VGND 0.0336f
C31134 VPWR.t2751 VGND 0.0396f
C31135 VPWR.t66 VGND 0.0331f
C31136 VPWR.t2959 VGND 0.0264f
C31137 VPWR.t1007 VGND 0.0311f
C31138 VPWR.t1971 VGND 0.0285f
C31139 VPWR.t2789 VGND 0.0258f
C31140 VPWR.t1365 VGND 0.0183f
C31141 VPWR.t6 VGND 0.0141f
C31142 VPWR.t2297 VGND 0.028f
C31143 VPWR.t2791 VGND 0.0109f
C31144 VPWR.t2085 VGND 0.0148f
C31145 VPWR.t1934 VGND 0.0309f
C31146 VPWR.t2204 VGND 0.0322f
C31147 VPWR.t1850 VGND 0.028f
C31148 VPWR.t2921 VGND 0.0158f
C31149 VPWR.t2684 VGND 0.0154f
C31150 VPWR.t998 VGND 0.0289f
C31151 VPWR.t1933 VGND 0.019f
C31152 VPWR.t1552 VGND 0.0164f
C31153 VPWR.t2158 VGND 0.0193f
C31154 VPWR.t1129 VGND 0.0181f
C31155 VPWR.t2844 VGND 0.0164f
C31156 VPWR.n8186 VGND 0.0162f
C31157 VPWR.n8187 VGND 0.00929f
C31158 VPWR.n8188 VGND 0.00525f
C31159 VPWR.n8189 VGND 0.0031f
C31160 VPWR.n8190 VGND 0.00524f
C31161 VPWR.n8191 VGND 0.00524f
C31162 VPWR.t371 VGND 0.00387f
C31163 VPWR.t3460 VGND 0.0179f
C31164 VPWR.t825 VGND 0.00453f
C31165 VPWR.n8192 VGND 0.0111f
C31166 VPWR.n8193 VGND 0.00912f
C31167 VPWR.n8194 VGND 0.0103f
C31168 VPWR.n8195 VGND 0.0173f
C31169 VPWR.n8196 VGND 0.00493f
C31170 VPWR.n8197 VGND 0.0049f
C31171 VPWR.n8198 VGND 0.00393f
C31172 VPWR.n8199 VGND 0.00362f
C31173 VPWR.n8200 VGND 0.00256f
C31174 VPWR.n8201 VGND 4.58e-19
C31175 VPWR.t2831 VGND 6.73e-19
C31176 VPWR.t1178 VGND 0.00127f
C31177 VPWR.n8202 VGND 0.00207f
C31178 VPWR.n8203 VGND 0.00456f
C31179 VPWR.n8204 VGND 8.39e-20
C31180 VPWR.n8205 VGND 5.98e-19
C31181 VPWR.n8206 VGND 5.12e-19
C31182 VPWR.n8207 VGND 3.13e-19
C31183 VPWR.n8208 VGND 1.77e-19
C31184 VPWR.n8209 VGND 1.76e-19
C31185 VPWR.n8210 VGND 5.48e-19
C31186 VPWR.n8211 VGND 0.00138f
C31187 VPWR.n8212 VGND 0.0057f
C31188 VPWR.n8214 VGND 5.71e-19
C31189 VPWR.n8215 VGND 3.29e-19
C31190 VPWR.n8216 VGND 3.95e-19
C31191 VPWR.n8217 VGND 4.17e-19
C31192 VPWR.n8218 VGND 2.85e-19
C31193 VPWR.n8219 VGND 4.17e-19
C31194 VPWR.n8220 VGND 5.05e-19
C31195 VPWR.n8221 VGND 4.83e-19
C31196 VPWR.n8222 VGND 2.85e-19
C31197 VPWR.n8223 VGND 3.95e-19
C31198 VPWR.n8224 VGND 2.85e-19
C31199 VPWR.n8225 VGND 4.11e-19
C31200 VPWR.n8226 VGND 4.11e-19
C31201 VPWR.n8227 VGND 7.39e-19
C31202 VPWR.n8228 VGND 5.19e-19
C31203 VPWR.n8229 VGND 7.39e-19
C31204 VPWR.n8230 VGND 4.11e-19
C31205 VPWR.n8231 VGND 4.11e-19
C31206 VPWR.n8232 VGND 3.07e-19
C31207 VPWR.n8233 VGND 1.76e-19
C31208 VPWR.n8234 VGND 4.39e-19
C31209 VPWR.n8235 VGND 6.14e-19
C31210 VPWR.n8236 VGND 7.97e-19
C31211 VPWR.n8237 VGND 3.13e-19
C31212 VPWR.n8238 VGND 6.55e-19
C31213 VPWR.n8239 VGND 6.26e-19
C31214 VPWR.n8240 VGND 3.7e-19
C31215 VPWR.n8241 VGND 1.21e-19
C31216 VPWR.t1501 VGND 0.00242f
C31217 VPWR.n8242 VGND 0.00484f
C31218 VPWR.n8243 VGND 1.31e-19
C31219 VPWR.n8244 VGND 6.09e-19
C31220 VPWR.n8245 VGND 6.65e-19
C31221 VPWR.n8246 VGND 5.12e-19
C31222 VPWR.n8247 VGND 5.41e-19
C31223 VPWR.n8248 VGND 5.12e-19
C31224 VPWR.n8249 VGND 4.27e-19
C31225 VPWR.n8250 VGND 9.96e-19
C31226 VPWR.n8251 VGND 0.00131f
C31227 VPWR.n8252 VGND 5.98e-19
C31228 VPWR.n8253 VGND 6.99e-19
C31229 VPWR.n8254 VGND 0.00218f
C31230 VPWR.n8255 VGND 0.00456f
C31231 VPWR.n8256 VGND 0.0014f
C31232 VPWR.n8257 VGND 0.00274f
C31233 VPWR.n8258 VGND 0.00179f
C31234 VPWR.n8259 VGND 0.00199f
C31235 VPWR.n8260 VGND 0.00639f
C31236 VPWR.n8261 VGND 0.00653f
C31237 VPWR.n8262 VGND 0.0031f
C31238 VPWR.n8263 VGND 0.00337f
C31239 VPWR.n8264 VGND 0.00524f
C31240 VPWR.n8265 VGND 0.0066f
C31241 VPWR.n8266 VGND 0.00524f
C31242 VPWR.n8267 VGND 0.00592f
C31243 VPWR.n8268 VGND 0.00524f
C31244 VPWR.t908 VGND 0.00234f
C31245 VPWR.n8269 VGND 0.00628f
C31246 VPWR.n8270 VGND 0.00398f
C31247 VPWR.n8271 VGND 0.00524f
C31248 VPWR.t3544 VGND 0.0592f
C31249 VPWR.n8272 VGND 0.0356f
C31250 VPWR.n8273 VGND 0.00484f
C31251 VPWR.n8274 VGND 0.00524f
C31252 VPWR.n8275 VGND 0.00506f
C31253 VPWR.n8276 VGND 0.00524f
C31254 VPWR.n8277 VGND 0.0066f
C31255 VPWR.n8278 VGND 0.00524f
C31256 VPWR.n8279 VGND 0.00506f
C31257 VPWR.n8280 VGND 0.00524f
C31258 VPWR.n8281 VGND 0.00393f
C31259 VPWR.n8282 VGND 0.00256f
C31260 VPWR.n8283 VGND 0.00515f
C31261 VPWR.n8284 VGND 0.0031f
C31262 VPWR.n8285 VGND 0.00524f
C31263 VPWR.n8286 VGND 0.00524f
C31264 VPWR.n8287 VGND 0.00393f
C31265 VPWR.n8288 VGND 0.00199f
C31266 VPWR.n8289 VGND 0.0016f
C31267 VPWR.n8290 VGND 0.00356f
C31268 VPWR.n8291 VGND 0.00911f
C31269 VPWR.n8292 VGND 0.00199f
C31270 VPWR.n8293 VGND 0.0015f
C31271 VPWR.n8294 VGND 0.0031f
C31272 VPWR.t3462 VGND 0.00911f
C31273 VPWR.t523 VGND 0.00391f
C31274 VPWR.n8295 VGND 0.0253f
C31275 VPWR.t524 VGND 0.00391f
C31276 VPWR.n8297 VGND 0.0126f
C31277 VPWR.t1722 VGND 0.00239f
C31278 VPWR.n8298 VGND 0.00421f
C31279 VPWR.n8299 VGND 0.00551f
C31280 VPWR.n8300 VGND 0.00524f
C31281 VPWR.n8301 VGND 9.68e-19
C31282 VPWR.n8302 VGND 0.00393f
C31283 VPWR.n8303 VGND 0.00179f
C31284 VPWR.n8304 VGND 0.00146f
C31285 VPWR.n8305 VGND 0.00292f
C31286 VPWR.n8306 VGND 0.00224f
C31287 VPWR.n8307 VGND 0.0031f
C31288 VPWR.n8308 VGND 0.0133f
C31289 VPWR.n8309 VGND 0.00524f
C31290 VPWR.n8310 VGND 0.0123f
C31291 VPWR.n8311 VGND 0.00524f
C31292 VPWR.n8312 VGND 0.00524f
C31293 VPWR.n8313 VGND 0.00524f
C31294 VPWR.n8314 VGND 0.00393f
C31295 VPWR.n8315 VGND 0.00199f
C31296 VPWR.n8316 VGND 0.00173f
C31297 VPWR.n8317 VGND 0.00109f
C31298 VPWR.n8318 VGND 0.0031f
C31299 VPWR.t1688 VGND 6.73e-19
C31300 VPWR.t2703 VGND 9.96e-19
C31301 VPWR.n8319 VGND 0.0018f
C31302 VPWR.n8320 VGND 0.00483f
C31303 VPWR.n8321 VGND 0.00103f
C31304 VPWR.n8322 VGND 0.00524f
C31305 VPWR.t2681 VGND 0.00102f
C31306 VPWR.t2718 VGND 0.00154f
C31307 VPWR.n8323 VGND 0.00483f
C31308 VPWR.n8324 VGND 0.00641f
C31309 VPWR.n8325 VGND 0.00125f
C31310 VPWR.n8326 VGND 0.00524f
C31311 VPWR.t1820 VGND 0.00453f
C31312 VPWR.n8327 VGND 0.0053f
C31313 VPWR.n8328 VGND 0.00123f
C31314 VPWR.n8329 VGND 0.00524f
C31315 VPWR.n8330 VGND 0.00393f
C31316 VPWR.n8331 VGND 0.00173f
C31317 VPWR.n8332 VGND 0.00525f
C31318 VPWR.n8333 VGND 0.0031f
C31319 VPWR.n8334 VGND 0.0123f
C31320 VPWR.n8335 VGND 0.00524f
C31321 VPWR.t1690 VGND 6.73e-19
C31322 VPWR.t1670 VGND 0.00127f
C31323 VPWR.n8336 VGND 0.00203f
C31324 VPWR.n8337 VGND 0.00951f
C31325 VPWR.n8338 VGND 0.00785f
C31326 VPWR.n8339 VGND 0.00524f
C31327 VPWR.n8340 VGND 0.0048f
C31328 VPWR.n8341 VGND 0.00994f
C31329 VPWR.n8342 VGND 0.00502f
C31330 VPWR.n8343 VGND 0.0022f
C31331 VPWR.n8344 VGND 0.00138f
C31332 VPWR.n8345 VGND 4.17e-19
C31333 VPWR.n8346 VGND 5.48e-19
C31334 VPWR.n8347 VGND 0.00138f
C31335 VPWR.n8348 VGND 0.0057f
C31336 VPWR.n8349 VGND 0.00139f
C31337 VPWR.n8350 VGND 9.06e-19
C31338 VPWR.n8351 VGND 8.11e-19
C31339 VPWR.n8352 VGND 3.95e-19
C31340 VPWR.n8353 VGND 1.76e-19
C31341 VPWR.n8354 VGND 3.95e-19
C31342 VPWR.n8355 VGND 7.68e-19
C31343 VPWR.n8356 VGND 5.05e-19
C31344 VPWR.n8357 VGND 1.76e-19
C31345 VPWR.n8358 VGND 5.48e-19
C31346 VPWR.n8360 VGND 0.1f
C31347 VPWR.n8361 VGND 0.1f
C31348 VPWR.n8362 VGND 6.54e-19
C31349 VPWR.n8363 VGND 8.67e-19
C31350 VPWR.n8364 VGND 3.95e-19
C31351 VPWR.n8365 VGND 4.61e-19
C31352 VPWR.n8366 VGND 2.41e-19
C31353 VPWR.n8367 VGND 3.95e-19
C31354 VPWR.n8368 VGND 0.00108f
C31355 VPWR.n8369 VGND 5.12e-19
C31356 VPWR.n8370 VGND 5.98e-19
C31357 VPWR.n8371 VGND 0.00171f
C31358 VPWR.n8372 VGND 0.00864f
C31359 VPWR.t393 VGND 0.0046f
C31360 VPWR.n8373 VGND 0.00931f
C31361 VPWR.t438 VGND 0.00398f
C31362 VPWR.n8374 VGND 0.015f
C31363 VPWR.n8375 VGND 0.013f
C31364 VPWR.n8376 VGND 3.13e-19
C31365 VPWR.n8377 VGND 4.84e-19
C31366 VPWR.n8378 VGND 6.26e-19
C31367 VPWR.n8379 VGND 9.96e-19
C31368 VPWR.n8380 VGND 5.41e-19
C31369 VPWR.n8381 VGND 4.84e-19
C31370 VPWR.n8382 VGND 8.54e-20
C31371 VPWR.n8383 VGND 5.69e-19
C31372 VPWR.n8384 VGND 0.00131f
C31373 VPWR.n8385 VGND 9.96e-19
C31374 VPWR.n8386 VGND 4.27e-19
C31375 VPWR.n8387 VGND 5.12e-19
C31376 VPWR.n8388 VGND 5.41e-19
C31377 VPWR.n8389 VGND 7.35e-19
C31378 VPWR.n8390 VGND 2.95e-19
C31379 VPWR.n8391 VGND 5.93e-19
C31380 VPWR.n8392 VGND 6.26e-19
C31381 VPWR.n8393 VGND 6.55e-19
C31382 VPWR.n8394 VGND 5.05e-19
C31383 VPWR.n8395 VGND 4.17e-19
C31384 VPWR.n8396 VGND 6.14e-19
C31385 VPWR.n8397 VGND 4.39e-19
C31386 VPWR.n8398 VGND 1.76e-19
C31387 VPWR.n8399 VGND 3.07e-19
C31388 VPWR.n8400 VGND 4.83e-19
C31389 VPWR.n8401 VGND 2.85e-19
C31390 VPWR.n8402 VGND 3.95e-19
C31391 VPWR.n8403 VGND 3.95e-19
C31392 VPWR.n8404 VGND 4.17e-19
C31393 VPWR.n8405 VGND 2.85e-19
C31394 VPWR.n8406 VGND 2.85e-19
C31395 VPWR.n8407 VGND 4.11e-19
C31396 VPWR.n8408 VGND 4.11e-19
C31397 VPWR.n8409 VGND 7.39e-19
C31398 VPWR.n8410 VGND 5.19e-19
C31399 VPWR.n8411 VGND 7.39e-19
C31400 VPWR.n8412 VGND 4.11e-19
C31401 VPWR.n8413 VGND 4.11e-19
C31402 VPWR.n8415 VGND 0.0057f
C31403 VPWR.n8416 VGND 0.00138f
C31404 VPWR.n8417 VGND 5.48e-19
C31405 VPWR.n8418 VGND 4.17e-19
C31406 VPWR.n8419 VGND 1.33e-19
C31407 VPWR.n8420 VGND 6.58e-20
C31408 VPWR.n8421 VGND 0.00118f
C31409 VPWR.n8422 VGND 8.05e-19
C31410 VPWR.n8423 VGND 0.00123f
C31411 VPWR.n8424 VGND 0.00774f
C31412 VPWR.n8425 VGND 0.0128f
C31413 VPWR.n8426 VGND 0.00179f
C31414 VPWR.n8427 VGND 0.00618f
C31415 VPWR.n8428 VGND 0.00179f
C31416 VPWR.n8429 VGND 0.00456f
C31417 VPWR.n8430 VGND 0.0129f
C31418 VPWR.t2251 VGND 0.00631f
C31419 VPWR.n8431 VGND 0.0103f
C31420 VPWR.n8432 VGND 0.0124f
C31421 VPWR.n8433 VGND 0.0133f
C31422 VPWR.n8434 VGND 0.00475f
C31423 VPWR.n8435 VGND 0.00393f
C31424 VPWR.n8436 VGND 0.00179f
C31425 VPWR.n8437 VGND 0.0031f
C31426 VPWR.n8438 VGND 0.00264f
C31427 VPWR.n8439 VGND 0.00646f
C31428 VPWR.t3043 VGND 0.00586f
C31429 VPWR.t3379 VGND 0.0225f
C31430 VPWR.n8440 VGND 0.0158f
C31431 VPWR.n8441 VGND 0.0138f
C31432 VPWR.n8442 VGND 0.0116f
C31433 VPWR.n8443 VGND 0.0148f
C31434 VPWR.n8444 VGND 0.00811f
C31435 VPWR.n8445 VGND 0.00516f
C31436 VPWR.n8446 VGND 0.00393f
C31437 VPWR.n8447 VGND 0.00524f
C31438 VPWR.n8448 VGND 0.00524f
C31439 VPWR.n8449 VGND 0.0107f
C31440 VPWR.n8450 VGND 0.00524f
C31441 VPWR.t2780 VGND 0.00172f
C31442 VPWR.n8451 VGND 0.00611f
C31443 VPWR.t2801 VGND 0.00166f
C31444 VPWR.n8452 VGND 0.00605f
C31445 VPWR.n8453 VGND 1.45e-19
C31446 VPWR.n8454 VGND 0.00718f
C31447 VPWR.n8455 VGND 0.00324f
C31448 VPWR.n8456 VGND 0.00888f
C31449 VPWR.t141 VGND 0.00387f
C31450 VPWR.n8457 VGND 0.00456f
C31451 VPWR.n8458 VGND 0.00283f
C31452 VPWR.n8459 VGND 0.00262f
C31453 VPWR.n8460 VGND 0.0031f
C31454 VPWR.t398 VGND 0.0046f
C31455 VPWR.n8461 VGND 0.00407f
C31456 VPWR.n8462 VGND 0.0023f
C31457 VPWR.n8463 VGND 0.00179f
C31458 VPWR.n8464 VGND 0.00199f
C31459 VPWR.n8465 VGND 0.00199f
C31460 VPWR.n8466 VGND 0.0143f
C31461 VPWR.t569 VGND 0.00387f
C31462 VPWR.n8467 VGND 0.00642f
C31463 VPWR.n8468 VGND 0.00796f
C31464 VPWR.n8469 VGND 0.00393f
C31465 VPWR.t3477 VGND 0.0592f
C31466 VPWR.n8470 VGND 0.041f
C31467 VPWR.n8471 VGND 0.00915f
C31468 VPWR.n8472 VGND 0.00524f
C31469 VPWR.t3411 VGND 0.0282f
C31470 VPWR.n8473 VGND 0.0512f
C31471 VPWR.n8474 VGND 0.0137f
C31472 VPWR.n8475 VGND 0.00524f
C31473 VPWR.n8476 VGND 0.0185f
C31474 VPWR.n8477 VGND 0.00524f
C31475 VPWR.n8478 VGND 0.0185f
C31476 VPWR.n8479 VGND 0.00524f
C31477 VPWR.n8480 VGND 0.00524f
C31478 VPWR.n8481 VGND 0.00524f
C31479 VPWR.n8482 VGND 0.0185f
C31480 VPWR.n8483 VGND 0.0179f
C31481 VPWR.t570 VGND 0.00387f
C31482 VPWR.n8484 VGND 0.0107f
C31483 VPWR.t399 VGND 0.0046f
C31484 VPWR.n8485 VGND 0.00379f
C31485 VPWR.n8486 VGND 0.00772f
C31486 VPWR.n8487 VGND 0.0031f
C31487 VPWR.n8488 VGND 0.00179f
C31488 VPWR.n8489 VGND 0.00262f
C31489 VPWR.t1222 VGND 0.00136f
C31490 VPWR.t1953 VGND 0.00136f
C31491 VPWR.n8490 VGND 0.00328f
C31492 VPWR.n8491 VGND 0.00757f
C31493 VPWR.t1220 VGND 0.00136f
C31494 VPWR.t1322 VGND 0.00136f
C31495 VPWR.n8492 VGND 0.00328f
C31496 VPWR.n8493 VGND 0.00757f
C31497 VPWR.n8494 VGND 0.00344f
C31498 VPWR.n8495 VGND 0.00262f
C31499 VPWR.n8496 VGND 0.00199f
C31500 VPWR.n8497 VGND 0.00139f
C31501 VPWR.n8498 VGND 0.00391f
C31502 VPWR.t220 VGND 0.00387f
C31503 VPWR.n8499 VGND 0.00846f
C31504 VPWR.n8500 VGND 0.00647f
C31505 VPWR.n8501 VGND 0.00393f
C31506 VPWR.n8502 VGND 0.011f
C31507 VPWR.n8503 VGND 0.0109f
C31508 VPWR.n8504 VGND 0.00524f
C31509 VPWR.t3409 VGND 0.0156f
C31510 VPWR.n8505 VGND 0.00597f
C31511 VPWR.n8506 VGND 0.0228f
C31512 VPWR.n8507 VGND 0.00971f
C31513 VPWR.n8508 VGND 0.0109f
C31514 VPWR.n8509 VGND 0.00524f
C31515 VPWR.n8510 VGND 0.0127f
C31516 VPWR.n8511 VGND 0.00956f
C31517 VPWR.n8512 VGND 0.00524f
C31518 VPWR.n8513 VGND 0.0135f
C31519 VPWR.n8514 VGND 0.00504f
C31520 VPWR.n8515 VGND 6.55e-19
C31521 VPWR.n8516 VGND 5.71e-19
C31522 VPWR.n8517 VGND 3.29e-19
C31523 VPWR.n8518 VGND 3.95e-19
C31524 VPWR.n8519 VGND 4.17e-19
C31525 VPWR.n8520 VGND 2.85e-19
C31526 VPWR.n8521 VGND 6.54e-19
C31527 VPWR.n8522 VGND 8.67e-19
C31528 VPWR.n8523 VGND 3.13e-19
C31529 VPWR.n8524 VGND 7.97e-19
C31530 VPWR.n8525 VGND 6.14e-19
C31531 VPWR.n8526 VGND 4.39e-19
C31532 VPWR.n8527 VGND 1.76e-19
C31533 VPWR.n8528 VGND 4.83e-19
C31534 VPWR.n8529 VGND 2.41e-19
C31535 VPWR.n8530 VGND 9.68e-19
C31536 VPWR.n8531 VGND 3.95e-19
C31537 VPWR.n8532 VGND 7.68e-19
C31538 VPWR.n8533 VGND 3.95e-19
C31539 VPWR.n8534 VGND 6.83e-19
C31540 VPWR.n8535 VGND 1.99e-19
C31541 VPWR.n8536 VGND 4.84e-19
C31542 VPWR.t221 VGND 0.00387f
C31543 VPWR.n8537 VGND 0.0074f
C31544 VPWR.n8538 VGND 0.00501f
C31545 VPWR.n8539 VGND 3.13e-19
C31546 VPWR.n8540 VGND 5.12e-19
C31547 VPWR.n8541 VGND 3.73e-19
C31548 VPWR.n8542 VGND 3.07e-19
C31549 VPWR.n8543 VGND 4.11e-19
C31550 VPWR.n8544 VGND 4.11e-19
C31551 VPWR.n8545 VGND 7.39e-19
C31552 VPWR.n8546 VGND 5.19e-19
C31553 VPWR.n8547 VGND 7.39e-19
C31554 VPWR.n8548 VGND 4.11e-19
C31555 VPWR.n8549 VGND 4.11e-19
C31556 VPWR.n8550 VGND 2.85e-19
C31557 VPWR.n8551 VGND 3.95e-19
C31558 VPWR.n8552 VGND 2.85e-19
C31559 VPWR.n8553 VGND 4.17e-19
C31560 VPWR.n8554 VGND 5.05e-19
C31561 VPWR.n8555 VGND 4.83e-19
C31562 VPWR.n8556 VGND 0.0062f
C31563 VPWR.n8557 VGND 3.7e-19
C31564 VPWR.n8558 VGND 3.7e-19
C31565 VPWR.n8559 VGND 3.7e-19
C31566 VPWR.n8560 VGND 5.12e-19
C31567 VPWR.n8561 VGND 5.41e-19
C31568 VPWR.n8562 VGND 5.12e-19
C31569 VPWR.n8563 VGND 4.27e-19
C31570 VPWR.n8564 VGND 9.96e-19
C31571 VPWR.n8565 VGND 0.00131f
C31572 VPWR.n8566 VGND 5.98e-19
C31573 VPWR.t1226 VGND 0.00131f
C31574 VPWR.t1187 VGND 4.27e-19
C31575 VPWR.n8567 VGND 0.00672f
C31576 VPWR.n8568 VGND 9.71e-19
C31577 VPWR.n8569 VGND 9.71e-19
C31578 VPWR.n8570 VGND 0.00673f
C31579 VPWR.n8571 VGND 0.00978f
C31580 VPWR.n8572 VGND 0.00702f
C31581 VPWR.n8573 VGND 6.99e-19
C31582 VPWR.n8574 VGND 0.00218f
C31583 VPWR.n8575 VGND 0.00137f
C31584 VPWR.n8576 VGND 5.92e-19
C31585 VPWR.n8577 VGND 5.05e-19
C31586 VPWR.n8578 VGND 4.17e-19
C31587 VPWR.n8579 VGND 5.48e-19
C31588 VPWR.n8581 VGND 0.0057f
C31589 VPWR.n8582 VGND 0.00138f
C31590 VPWR.n8583 VGND 5.48e-19
C31591 VPWR.n8584 VGND 1.76e-19
C31592 VPWR.n8585 VGND 8.11e-19
C31593 VPWR.n8586 VGND 3.95e-19
C31594 VPWR.n8587 VGND 1.77e-19
C31595 VPWR.n8588 VGND 3.13e-19
C31596 VPWR.n8589 VGND 5.12e-19
C31597 VPWR.n8590 VGND 5.98e-19
C31598 VPWR.n8591 VGND 4.27e-19
C31599 VPWR.n8592 VGND 4.58e-19
C31600 VPWR.n8593 VGND 8.39e-20
C31601 VPWR.t3266 VGND 0.0016f
C31602 VPWR.t1485 VGND 0.0016f
C31603 VPWR.n8594 VGND 0.00377f
C31604 VPWR.n8595 VGND 0.006f
C31605 VPWR.t3311 VGND 0.00166f
C31606 VPWR.t3092 VGND 0.00225f
C31607 VPWR.n8596 VGND 0.0045f
C31608 VPWR.t1483 VGND 0.0016f
C31609 VPWR.t1479 VGND 0.0016f
C31610 VPWR.n8597 VGND 0.00379f
C31611 VPWR.n8598 VGND 0.00755f
C31612 VPWR.n8599 VGND 0.00697f
C31613 VPWR.n8600 VGND 0.00475f
C31614 VPWR.n8601 VGND 0.00524f
C31615 VPWR.t3094 VGND 0.00166f
C31616 VPWR.t3096 VGND 0.00166f
C31617 VPWR.n8602 VGND 0.00345f
C31618 VPWR.t1481 VGND 0.00655f
C31619 VPWR.n8603 VGND 0.00997f
C31620 VPWR.n8604 VGND 0.00419f
C31621 VPWR.n8605 VGND 0.00524f
C31622 VPWR.n8606 VGND 0.00393f
C31623 VPWR.n8607 VGND 5.44e-19
C31624 VPWR.t3098 VGND 0.00695f
C31625 VPWR.n8608 VGND 0.00844f
C31626 VPWR.n8609 VGND 0.00262f
C31627 VPWR.n8610 VGND 0.00199f
C31628 VPWR.t650 VGND 0.00387f
C31629 VPWR.t3564 VGND 0.0282f
C31630 VPWR.n8611 VGND 0.0102f
C31631 VPWR.n8612 VGND 0.0489f
C31632 VPWR.n8613 VGND 0.01f
C31633 VPWR.n8614 VGND 0.00837f
C31634 VPWR.n8615 VGND 0.00471f
C31635 VPWR.t3356 VGND 0.00911f
C31636 VPWR.t62 VGND 0.00391f
C31637 VPWR.n8616 VGND 0.0253f
C31638 VPWR.t61 VGND 0.00391f
C31639 VPWR.n8618 VGND 0.0138f
C31640 VPWR.t651 VGND 0.00387f
C31641 VPWR.n8619 VGND 0.00837f
C31642 VPWR.t1684 VGND 0.00102f
C31643 VPWR.t1774 VGND 0.00102f
C31644 VPWR.n8620 VGND 0.00221f
C31645 VPWR.n8621 VGND 0.00598f
C31646 VPWR.t3566 VGND 0.0289f
C31647 VPWR.t656 VGND 0.00387f
C31648 VPWR.n8622 VGND 0.0604f
C31649 VPWR.n8623 VGND 0.0146f
C31650 VPWR.n8624 VGND 0.0117f
C31651 VPWR.t1784 VGND 0.0016f
C31652 VPWR.t2427 VGND 0.00208f
C31653 VPWR.n8625 VGND 0.00413f
C31654 VPWR.n8626 VGND 0.0155f
C31655 VPWR.n8627 VGND 0.0137f
C31656 VPWR.n8628 VGND 0.0133f
C31657 VPWR.t657 VGND 0.00387f
C31658 VPWR.n8629 VGND 0.00837f
C31659 VPWR.n8630 VGND 0.00333f
C31660 VPWR.n8631 VGND 0.00393f
C31661 VPWR.n8632 VGND 0.00156f
C31662 VPWR.n8633 VGND 0.00525f
C31663 VPWR.n8634 VGND 0.0031f
C31664 VPWR.n8635 VGND 0.00524f
C31665 VPWR.n8636 VGND 0.00524f
C31666 VPWR.t3187 VGND 0.00524f
C31667 VPWR.n8637 VGND 0.0108f
C31668 VPWR.n8638 VGND 0.00448f
C31669 VPWR.n8639 VGND 0.00869f
C31670 VPWR.n8640 VGND 0.00719f
C31671 VPWR.n8641 VGND 0.00179f
C31672 VPWR.n8642 VGND 0.00199f
C31673 VPWR.n8643 VGND 0.00154f
C31674 VPWR.n8644 VGND 0.0031f
C31675 VPWR.n8645 VGND 0.00166f
C31676 VPWR.n8646 VGND 0.00524f
C31677 VPWR.t3185 VGND 0.00102f
C31678 VPWR.t2259 VGND 0.00154f
C31679 VPWR.n8647 VGND 0.00483f
C31680 VPWR.n8648 VGND 0.00671f
C31681 VPWR.t2691 VGND 0.00234f
C31682 VPWR.n8649 VGND 0.00391f
C31683 VPWR.n8650 VGND 5.14e-19
C31684 VPWR.n8651 VGND 0.00524f
C31685 VPWR.n8652 VGND 0.00153f
C31686 VPWR.n8653 VGND 0.00524f
C31687 VPWR.n8654 VGND 0.00393f
C31688 VPWR.n8655 VGND 0.00173f
C31689 VPWR.n8656 VGND 0.00525f
C31690 VPWR.n8657 VGND 0.0031f
C31691 VPWR.n8658 VGND 0.0101f
C31692 VPWR.n8659 VGND 0.00524f
C31693 VPWR.t2855 VGND 6.73e-19
C31694 VPWR.t3031 VGND 9.96e-19
C31695 VPWR.n8660 VGND 0.00176f
C31696 VPWR.n8661 VGND 0.0102f
C31697 VPWR.n8662 VGND 0.0101f
C31698 VPWR.n8663 VGND 0.00524f
C31699 VPWR.n8664 VGND 0.0115f
C31700 VPWR.n8665 VGND 0.00524f
C31701 VPWR.t3277 VGND 0.00453f
C31702 VPWR.n8666 VGND 0.0116f
C31703 VPWR.n8667 VGND 0.00912f
C31704 VPWR.n8668 VGND 0.00524f
C31705 VPWR.n8669 VGND 0.00524f
C31706 VPWR.n8670 VGND 0.00524f
C31707 VPWR.n8671 VGND 0.00393f
C31708 VPWR.n8672 VGND 0.00444f
C31709 VPWR.t1662 VGND 0.00239f
C31710 VPWR.t2853 VGND 6.73e-19
C31711 VPWR.t1732 VGND 0.00127f
C31712 VPWR.n8673 VGND 0.00204f
C31713 VPWR.n8674 VGND 0.00705f
C31714 VPWR.n8675 VGND 0.00815f
C31715 VPWR.n8676 VGND 0.00873f
C31716 VPWR.n8677 VGND 0.0396f
C31717 VPWR.t1661 VGND 0.0309f
C31718 VPWR.t60 VGND 0.0141f
C31719 VPWR.t2852 VGND 0.0183f
C31720 VPWR.t1731 VGND 0.0258f
C31721 VPWR.t1792 VGND 0.0285f
C31722 VPWR.t1685 VGND 0.0311f
C31723 VPWR.t3276 VGND 0.0264f
C31724 VPWR.t649 VGND 0.0331f
C31725 VPWR.t2854 VGND 0.0396f
C31726 VPWR.t3030 VGND 0.0336f
C31727 VPWR.t1686 VGND 0.0228f
C31728 VPWR.t1791 VGND 0.0248f
C31729 VPWR.t2258 VGND 0.0154f
C31730 VPWR.t2690 VGND 0.0163f
C31731 VPWR.t3184 VGND 0.0211f
C31732 VPWR.t3235 VGND 0.0299f
C31733 VPWR.t1683 VGND 0.0151f
C31734 VPWR.t1773 VGND 0.0158f
C31735 VPWR.t1783 VGND 0.0361f
C31736 VPWR.t2426 VGND 0.0305f
C31737 VPWR.t655 VGND 0.0158f
C31738 VPWR.t3186 VGND 0.0319f
C31739 VPWR.t1553 VGND 0.0453f
C31740 VPWR.t1797 VGND 0.025f
C31741 VPWR.t3107 VGND 0.0311f
C31742 VPWR.t3188 VGND 0.0124f
C31743 VPWR.t222 VGND 0.0463f
C31744 VPWR.t2343 VGND 0.026f
C31745 VPWR.t688 VGND 0.0144f
C31746 VPWR.t2341 VGND 0.0153f
C31747 VPWR.t2347 VGND 0.0289f
C31748 VPWR.t2345 VGND 0.0205f
C31749 VPWR.t3233 VGND 0.0109f
C31750 VPWR.t1829 VGND 0.00537f
C31751 VPWR.t820 VGND 0.0153f
C31752 VPWR.t3221 VGND 0.0446f
C31753 VPWR.t887 VGND 0.0154f
C31754 VPWR.t2768 VGND 0.0121f
C31755 VPWR.t1227 VGND 0.00722f
C31756 VPWR.t823 VGND 0.0156f
C31757 VPWR.t2018 VGND 0.0336f
C31758 VPWR.t2755 VGND 0.0242f
C31759 VPWR.t258 VGND 0.0331f
C31760 VPWR.t1757 VGND 0.0418f
C31761 VPWR.t822 VGND 0.0264f
C31762 VPWR.t2767 VGND 0.0151f
C31763 VPWR.t2006 VGND 0.0178f
C31764 VPWR.t1798 VGND 0.0181f
C31765 VPWR.t2745 VGND 0.0121f
C31766 VPWR.t1649 VGND 0.0141f
C31767 VPWR.t2289 VGND 0.0163f
C31768 VPWR.t909 VGND 0.0361f
C31769 VPWR.t2004 VGND 0.0309f
C31770 VPWR.t3236 VGND 0.0183f
C31771 VPWR.n8678 VGND 0.0182f
C31772 VPWR.n8679 VGND 0.01f
C31773 VPWR.n8680 VGND 0.00199f
C31774 VPWR.n8681 VGND 0.00179f
C31775 VPWR.n8682 VGND 0.00202f
C31776 VPWR.n8683 VGND 0.0015f
C31777 VPWR.n8684 VGND 0.0109f
C31778 VPWR.n8685 VGND 0.00393f
C31779 VPWR.t2290 VGND 0.00239f
C31780 VPWR.n8686 VGND 0.00388f
C31781 VPWR.n8687 VGND 0.00102f
C31782 VPWR.n8688 VGND 0.00524f
C31783 VPWR.t1650 VGND 0.00102f
C31784 VPWR.t910 VGND 0.00154f
C31785 VPWR.n8689 VGND 0.00483f
C31786 VPWR.n8690 VGND 0.00636f
C31787 VPWR.n8691 VGND 0.00113f
C31788 VPWR.n8692 VGND 0.00452f
C31789 VPWR.n8693 VGND 3.95e-19
C31790 VPWR.n8694 VGND 5.05e-19
C31791 VPWR.n8695 VGND 5.05e-19
C31792 VPWR.n8696 VGND 0.00139f
C31793 VPWR.n8697 VGND 0.0323f
C31794 VPWR.n8699 VGND 9.06e-19
C31795 VPWR.n8700 VGND 5.48e-19
C31796 VPWR.n8701 VGND 3.07e-19
C31797 VPWR.n8702 VGND 0.00138f
C31798 VPWR.n8703 VGND 0.00222f
C31799 VPWR.n8704 VGND 0.00124f
C31800 VPWR.n8705 VGND 2.62e-19
C31801 VPWR.n8706 VGND 7.88e-19
C31802 VPWR.n8707 VGND 6.83e-19
C31803 VPWR.n8708 VGND 4.84e-19
C31804 VPWR.n8709 VGND 3.13e-19
C31805 VPWR.n8710 VGND 9.96e-19
C31806 VPWR.n8711 VGND 5.44e-19
C31807 VPWR.n8712 VGND 9.68e-19
C31808 VPWR.n8713 VGND 4.27e-19
C31809 VPWR.n8714 VGND 1.71e-19
C31810 VPWR.n8715 VGND 2.56e-19
C31811 VPWR.n8716 VGND 8.97e-19
C31812 VPWR.n8717 VGND 3.42e-19
C31813 VPWR.n8718 VGND 4.27e-19
C31814 VPWR.n8719 VGND 3.99e-19
C31815 VPWR.n8720 VGND 3.51e-19
C31816 VPWR.n8721 VGND 5.12e-19
C31817 VPWR.n8722 VGND 5.41e-19
C31818 VPWR.n8723 VGND 3.29e-19
C31819 VPWR.n8724 VGND 4.39e-19
C31820 VPWR.n8725 VGND 9e-19
C31821 VPWR.n8726 VGND 8.67e-19
C31822 VPWR.n8727 VGND 6.54e-19
C31823 VPWR.n8728 VGND 9.06e-19
C31824 VPWR.n8729 VGND 0.00138f
C31825 VPWR.n8730 VGND 5.48e-19
C31826 VPWR.n8731 VGND 6.14e-19
C31827 VPWR.t260 VGND 0.00387f
C31828 VPWR.n8732 VGND 0.00837f
C31829 VPWR.n8733 VGND 0.00179f
C31830 VPWR.t888 VGND 0.00633f
C31831 VPWR.n8734 VGND 0.00969f
C31832 VPWR.t3222 VGND 0.00234f
C31833 VPWR.t3234 VGND 0.00166f
C31834 VPWR.t2346 VGND 0.00225f
C31835 VPWR.n8735 VGND 0.0045f
C31836 VPWR.n8736 VGND 0.00745f
C31837 VPWR.t821 VGND 0.00102f
C31838 VPWR.t1830 VGND 0.00102f
C31839 VPWR.n8737 VGND 0.00221f
C31840 VPWR.t2344 VGND 0.00682f
C31841 VPWR.n8738 VGND 0.0126f
C31842 VPWR.t690 VGND 0.00387f
C31843 VPWR.n8739 VGND 0.00224f
C31844 VPWR.t3410 VGND 0.00911f
C31845 VPWR.t224 VGND 0.00391f
C31846 VPWR.n8740 VGND 0.0253f
C31847 VPWR.t223 VGND 0.00391f
C31848 VPWR.n8742 VGND 0.0138f
C31849 VPWR.n8743 VGND 0.00444f
C31850 VPWR.t3469 VGND 0.00911f
C31851 VPWR.t723 VGND 0.00391f
C31852 VPWR.n8744 VGND 0.0253f
C31853 VPWR.t724 VGND 0.00391f
C31854 VPWR.n8746 VGND 0.0138f
C31855 VPWR.n8747 VGND 0.0112f
C31856 VPWR.n8748 VGND 0.00487f
C31857 VPWR.n8749 VGND 0.0031f
C31858 VPWR.n8750 VGND 0.00524f
C31859 VPWR.n8751 VGND 0.00524f
C31860 VPWR.t689 VGND 0.00387f
C31861 VPWR.t3573 VGND 0.0179f
C31862 VPWR.t2348 VGND 0.00166f
C31863 VPWR.t2342 VGND 0.00166f
C31864 VPWR.n8752 VGND 0.00341f
C31865 VPWR.n8753 VGND 0.013f
C31866 VPWR.n8754 VGND 0.00695f
C31867 VPWR.n8755 VGND 0.00613f
C31868 VPWR.n8756 VGND 0.0173f
C31869 VPWR.n8757 VGND 0.00493f
C31870 VPWR.n8758 VGND 0.00473f
C31871 VPWR.n8759 VGND 0.00393f
C31872 VPWR.n8760 VGND 0.00262f
C31873 VPWR.n8761 VGND 0.00179f
C31874 VPWR.n8762 VGND 0.00602f
C31875 VPWR.n8763 VGND 0.00154f
C31876 VPWR.n8764 VGND 0.00333f
C31877 VPWR.n8765 VGND 0.00393f
C31878 VPWR.n8766 VGND 0.00166f
C31879 VPWR.n8767 VGND 0.00391f
C31880 VPWR.n8768 VGND 2.52e-19
C31881 VPWR.n8769 VGND 0.00393f
C31882 VPWR.n8770 VGND 0.00473f
C31883 VPWR.n8771 VGND 0.00182f
C31884 VPWR.n8772 VGND 0.00173f
C31885 VPWR.n8773 VGND 0.00525f
C31886 VPWR.n8774 VGND 0.0031f
C31887 VPWR.n8775 VGND 0.0101f
C31888 VPWR.n8776 VGND 0.00524f
C31889 VPWR.t2756 VGND 6.73e-19
C31890 VPWR.t2019 VGND 9.96e-19
C31891 VPWR.n8777 VGND 0.00176f
C31892 VPWR.n8778 VGND 0.0102f
C31893 VPWR.n8779 VGND 0.0101f
C31894 VPWR.n8780 VGND 0.00524f
C31895 VPWR.n8781 VGND 0.0115f
C31896 VPWR.n8782 VGND 0.00524f
C31897 VPWR.t3565 VGND 0.0231f
C31898 VPWR.t1758 VGND 0.00453f
C31899 VPWR.n8783 VGND 0.0116f
C31900 VPWR.n8784 VGND 0.0337f
C31901 VPWR.n8785 VGND 0.00524f
C31902 VPWR.t259 VGND 0.00387f
C31903 VPWR.n8786 VGND 0.00837f
C31904 VPWR.n8787 VGND 0.00508f
C31905 VPWR.n8788 VGND 0.00367f
C31906 VPWR.n8789 VGND 9.06e-19
C31907 VPWR.n8790 VGND 0.00138f
C31908 VPWR.n8791 VGND 6.26e-19
C31909 VPWR.n8792 VGND 8.32e-19
C31910 VPWR.n8793 VGND 6.83e-19
C31911 VPWR.n8794 VGND 1.71e-19
C31912 VPWR.n8795 VGND 4.27e-19
C31913 VPWR.n8796 VGND 8.54e-20
C31914 VPWR.n8797 VGND 9.07e-19
C31915 VPWR.n8798 VGND 4.27e-19
C31916 VPWR.n8799 VGND 6.83e-19
C31917 VPWR.n8800 VGND 3.7e-19
C31918 VPWR.n8801 VGND 2.85e-19
C31919 VPWR.n8802 VGND 2.85e-19
C31920 VPWR.n8803 VGND 4.17e-19
C31921 VPWR.n8804 VGND 4.11e-19
C31922 VPWR.n8805 VGND 4.11e-19
C31923 VPWR.n8806 VGND 7.39e-19
C31924 VPWR.n8807 VGND 5.19e-19
C31925 VPWR.n8808 VGND 7.39e-19
C31926 VPWR.n8809 VGND 4.11e-19
C31927 VPWR.n8810 VGND 5.27e-19
C31928 VPWR.n8811 VGND 3.73e-19
C31929 VPWR.n8812 VGND 2.41e-19
C31930 VPWR.n8813 VGND 4.83e-19
C31931 VPWR.n8814 VGND 4.17e-19
C31932 VPWR.n8815 VGND 5.71e-19
C31933 VPWR.n8816 VGND 4.17e-19
C31934 VPWR.n8817 VGND 4.83e-19
C31935 VPWR.n8818 VGND 4.61e-19
C31936 VPWR.n8819 VGND 4.61e-19
C31937 VPWR.n8820 VGND 4.11e-19
C31938 VPWR.n8822 VGND 0.1f
C31939 VPWR.n8823 VGND 0.1f
C31940 VPWR.n8825 VGND 9.06e-19
C31941 VPWR.n8826 VGND 5.48e-19
C31942 VPWR.n8827 VGND 3.07e-19
C31943 VPWR.n8828 VGND 1.76e-19
C31944 VPWR.n8829 VGND 2.63e-19
C31945 VPWR.n8830 VGND 9.42e-19
C31946 VPWR.n8831 VGND 6.27e-19
C31947 VPWR.n8832 VGND 0.00199f
C31948 VPWR.n8833 VGND 0.0108f
C31949 VPWR.n8834 VGND 0.00688f
C31950 VPWR.n8835 VGND 5.98e-19
C31951 VPWR.n8836 VGND 0.00112f
C31952 VPWR.n8837 VGND 4.27e-19
C31953 VPWR.n8838 VGND 0.0012f
C31954 VPWR.n8839 VGND 4.55e-19
C31955 VPWR.n8840 VGND 0.00516f
C31956 VPWR.n8841 VGND 4.84e-19
C31957 VPWR.n8842 VGND 6.83e-19
C31958 VPWR.n8843 VGND 4.84e-19
C31959 VPWR.n8844 VGND 3.13e-19
C31960 VPWR.n8845 VGND 9.96e-19
C31961 VPWR.n8846 VGND 0.00538f
C31962 VPWR.n8847 VGND 9.68e-19
C31963 VPWR.n8848 VGND 4.27e-19
C31964 VPWR.n8849 VGND 2.56e-19
C31965 VPWR.t2859 VGND 0.00676f
C31966 VPWR.n8850 VGND 0.00976f
C31967 VPWR.n8851 VGND 4.48e-19
C31968 VPWR.n8852 VGND 0.00643f
C31969 VPWR.n8853 VGND 3.42e-19
C31970 VPWR.n8854 VGND 3.29e-19
C31971 VPWR.n8855 VGND 4.39e-19
C31972 VPWR.n8856 VGND 9e-19
C31973 VPWR.n8857 VGND 8.67e-19
C31974 VPWR.n8858 VGND 6.54e-19
C31975 VPWR.n8859 VGND 9.06e-19
C31976 VPWR.n8860 VGND 0.00138f
C31977 VPWR.n8861 VGND 5.48e-19
C31978 VPWR.n8862 VGND 6.14e-19
C31979 VPWR.t410 VGND 0.00387f
C31980 VPWR.t3413 VGND 0.0179f
C31981 VPWR.t2815 VGND 0.00453f
C31982 VPWR.n8863 VGND 0.0111f
C31983 VPWR.n8864 VGND 0.0116f
C31984 VPWR.n8865 VGND 0.00568f
C31985 VPWR.n8866 VGND 0.0173f
C31986 VPWR.n8867 VGND 0.00493f
C31987 VPWR.t411 VGND 0.00387f
C31988 VPWR.n8868 VGND 0.00837f
C31989 VPWR.n8869 VGND 0.00146f
C31990 VPWR.t890 VGND 0.00654f
C31991 VPWR.n8870 VGND 0.0111f
C31992 VPWR.t2894 VGND 0.00238f
C31993 VPWR.n8871 VGND 0.0053f
C31994 VPWR.t2114 VGND 0.00102f
C31995 VPWR.t1826 VGND 0.00102f
C31996 VPWR.n8872 VGND 0.00221f
C31997 VPWR.n8873 VGND 0.00563f
C31998 VPWR.t2481 VGND 0.00663f
C31999 VPWR.n8874 VGND 0.00848f
C32000 VPWR.t3509 VGND 0.00911f
C32001 VPWR.t209 VGND 0.00391f
C32002 VPWR.n8875 VGND 0.0253f
C32003 VPWR.t208 VGND 0.00391f
C32004 VPWR.n8877 VGND 0.0138f
C32005 VPWR.t3345 VGND 0.00911f
C32006 VPWR.t197 VGND 0.00391f
C32007 VPWR.n8878 VGND 0.0253f
C32008 VPWR.t198 VGND 0.00391f
C32009 VPWR.n8880 VGND 0.0138f
C32010 VPWR.n8881 VGND 0.0109f
C32011 VPWR.n8882 VGND 0.00444f
C32012 VPWR.n8883 VGND 0.0031f
C32013 VPWR.n8884 VGND 0.00524f
C32014 VPWR.n8885 VGND 0.00475f
C32015 VPWR.t3130 VGND 0.00137f
C32016 VPWR.t2483 VGND -2.18e-20
C32017 VPWR.n8886 VGND 0.00629f
C32018 VPWR.n8887 VGND 0.00759f
C32019 VPWR.n8888 VGND 0.00115f
C32020 VPWR.n8889 VGND 0.00179f
C32021 VPWR.n8890 VGND 0.00333f
C32022 VPWR.n8891 VGND 0.00152f
C32023 VPWR.n8892 VGND 0.00393f
C32024 VPWR.n8893 VGND 0.00393f
C32025 VPWR.n8894 VGND 0.00473f
C32026 VPWR.n8895 VGND 0.00182f
C32027 VPWR.n8896 VGND 0.00115f
C32028 VPWR.t1368 VGND 6.73e-19
C32029 VPWR.t841 VGND 9.96e-19
C32030 VPWR.n8897 VGND 0.00178f
C32031 VPWR.n8898 VGND 0.00661f
C32032 VPWR.n8899 VGND 0.00248f
C32033 VPWR.n8900 VGND 0.0031f
C32034 VPWR.n8901 VGND 0.00524f
C32035 VPWR.n8902 VGND 0.00524f
C32036 VPWR.n8903 VGND 0.00393f
C32037 VPWR.n8904 VGND 0.00525f
C32038 VPWR.n8905 VGND 0.00173f
C32039 VPWR.n8906 VGND 0.0031f
C32040 VPWR.n8907 VGND 0.00172f
C32041 VPWR.n8908 VGND 0.00524f
C32042 VPWR.t3104 VGND 0.00184f
C32043 VPWR.t2162 VGND 0.00166f
C32044 VPWR.n8909 VGND 0.00358f
C32045 VPWR.t2754 VGND 6.73e-19
C32046 VPWR.t2857 VGND 0.00127f
C32047 VPWR.n8910 VGND 0.00203f
C32048 VPWR.n8911 VGND 0.00353f
C32049 VPWR.n8912 VGND 0.00208f
C32050 VPWR.n8913 VGND 9.58e-19
C32051 VPWR.n8914 VGND 0.00524f
C32052 VPWR.n8915 VGND 0.00125f
C32053 VPWR.n8916 VGND 0.00367f
C32054 VPWR.n8917 VGND 9.06e-19
C32055 VPWR.n8918 VGND 0.00138f
C32056 VPWR.n8919 VGND 8.26e-19
C32057 VPWR.t2569 VGND 0.0024f
C32058 VPWR.n8920 VGND 0.00522f
C32059 VPWR.n8921 VGND 0.00228f
C32060 VPWR.n8922 VGND 4.84e-19
C32061 VPWR.n8923 VGND 4.27e-19
C32062 VPWR.n8924 VGND 8.54e-20
C32063 VPWR.t562 VGND 0.00387f
C32064 VPWR.n8925 VGND 0.008f
C32065 VPWR.n8926 VGND 0.00127f
C32066 VPWR.n8927 VGND 4.48e-19
C32067 VPWR.n8928 VGND 4.27e-19
C32068 VPWR.n8929 VGND 6.83e-19
C32069 VPWR.n8930 VGND 3.7e-19
C32070 VPWR.n8931 VGND 9.68e-19
C32071 VPWR.n8932 VGND 9.96e-19
C32072 VPWR.n8933 VGND 5.41e-19
C32073 VPWR.n8934 VGND 7.4e-19
C32074 VPWR.n8935 VGND 5.71e-19
C32075 VPWR.n8936 VGND 4.17e-19
C32076 VPWR.n8937 VGND 4.83e-19
C32077 VPWR.n8938 VGND 4.61e-19
C32078 VPWR.n8939 VGND 4.61e-19
C32079 VPWR.n8940 VGND 4.11e-19
C32080 VPWR.n8942 VGND 0.1f
C32081 VPWR.n8943 VGND 0.1f
C32082 VPWR.n8944 VGND 7.39e-19
C32083 VPWR.n8945 VGND 4.11e-19
C32084 VPWR.n8946 VGND 4.17e-19
C32085 VPWR.n8947 VGND 3.51e-19
C32086 VPWR.n8948 VGND 4.61e-19
C32087 VPWR.n8949 VGND 4.39e-19
C32088 VPWR.n8950 VGND 3.29e-19
C32089 VPWR.n8951 VGND 5.27e-19
C32090 VPWR.n8952 VGND 2.85e-19
C32091 VPWR.n8953 VGND 2.85e-19
C32092 VPWR.n8954 VGND 4.17e-19
C32093 VPWR.n8955 VGND 6.54e-19
C32094 VPWR.n8956 VGND 8.67e-19
C32095 VPWR.n8957 VGND 4.11e-19
C32096 VPWR.n8959 VGND 0.0057f
C32097 VPWR.n8960 VGND 0.00138f
C32098 VPWR.n8961 VGND 9.06e-19
C32099 VPWR.n8962 VGND 5.48e-19
C32100 VPWR.n8963 VGND 3.07e-19
C32101 VPWR.n8964 VGND 0.00138f
C32102 VPWR.n8965 VGND 0.00222f
C32103 VPWR.t2109 VGND 0.00676f
C32104 VPWR.t3374 VGND 0.0289f
C32105 VPWR.t64 VGND 0.00387f
C32106 VPWR.n8966 VGND 0.0604f
C32107 VPWR.n8967 VGND 0.0143f
C32108 VPWR.n8968 VGND 0.013f
C32109 VPWR.n8969 VGND 0.00665f
C32110 VPWR.n8970 VGND 0.00452f
C32111 VPWR.n8971 VGND 0.00393f
C32112 VPWR.n8972 VGND 0.00199f
C32113 VPWR.n8973 VGND 0.00394f
C32114 VPWR.n8974 VGND 0.00179f
C32115 VPWR.t346 VGND 0.0046f
C32116 VPWR.n8975 VGND 0.00407f
C32117 VPWR.t3481 VGND 0.0592f
C32118 VPWR.t1666 VGND 0.00102f
C32119 VPWR.t2103 VGND 0.00102f
C32120 VPWR.n8976 VGND 0.00217f
C32121 VPWR.n8977 VGND 0.00555f
C32122 VPWR.n8978 VGND 0.0355f
C32123 VPWR.t363 VGND 0.0046f
C32124 VPWR.n8979 VGND 0.00407f
C32125 VPWR.n8980 VGND 0.00393f
C32126 VPWR.n8981 VGND 0.00323f
C32127 VPWR.n8982 VGND 0.00524f
C32128 VPWR.n8983 VGND 0.0031f
C32129 VPWR.n8984 VGND 0.00119f
C32130 VPWR.t1448 VGND 0.0024f
C32131 VPWR.n8985 VGND 0.00564f
C32132 VPWR.t681 VGND 0.0046f
C32133 VPWR.n8986 VGND 0.00407f
C32134 VPWR.n8987 VGND 0.00166f
C32135 VPWR.n8988 VGND 0.00475f
C32136 VPWR.t1360 VGND 6.73e-19
C32137 VPWR.t2493 VGND 0.00127f
C32138 VPWR.n8989 VGND 0.00203f
C32139 VPWR.n8990 VGND 0.00594f
C32140 VPWR.n8991 VGND 0.00355f
C32141 VPWR.n8992 VGND 0.00524f
C32142 VPWR.n8993 VGND 0.00614f
C32143 VPWR.n8994 VGND 0.00524f
C32144 VPWR.n8995 VGND 0.00506f
C32145 VPWR.n8996 VGND 0.00524f
C32146 VPWR.t3333 VGND 0.0592f
C32147 VPWR.n8997 VGND 0.0356f
C32148 VPWR.n8998 VGND 0.00484f
C32149 VPWR.n8999 VGND 0.00524f
C32150 VPWR.t1724 VGND 0.00453f
C32151 VPWR.n9000 VGND 0.00799f
C32152 VPWR.n9001 VGND 0.00438f
C32153 VPWR.n9002 VGND 0.00524f
C32154 VPWR.n9003 VGND 0.00553f
C32155 VPWR.n9004 VGND 0.00524f
C32156 VPWR.t1362 VGND 6.73e-19
C32157 VPWR.t1627 VGND 9.96e-19
C32158 VPWR.n9005 VGND 0.00176f
C32159 VPWR.n9006 VGND 0.00658f
C32160 VPWR.n9007 VGND 0.00484f
C32161 VPWR.n9008 VGND 0.00524f
C32162 VPWR.n9009 VGND 0.00506f
C32163 VPWR.n9010 VGND 0.00524f
C32164 VPWR.n9011 VGND 0.0066f
C32165 VPWR.n9012 VGND 0.00524f
C32166 VPWR.n9013 VGND 0.00639f
C32167 VPWR.n9014 VGND 0.00524f
C32168 VPWR.t682 VGND 0.0046f
C32169 VPWR.n9015 VGND 0.00407f
C32170 VPWR.n9016 VGND 0.00264f
C32171 VPWR.n9017 VGND 0.0031f
C32172 VPWR.t345 VGND 0.0046f
C32173 VPWR.t896 VGND 0.00234f
C32174 VPWR.n9018 VGND 0.00607f
C32175 VPWR.n9019 VGND 0.00145f
C32176 VPWR.n9020 VGND 0.00259f
C32177 VPWR.n9021 VGND 0.00475f
C32178 VPWR.n9022 VGND 0.00592f
C32179 VPWR.n9023 VGND 0.00524f
C32180 VPWR.n9024 VGND 0.0066f
C32181 VPWR.n9025 VGND 0.00524f
C32182 VPWR.n9026 VGND 0.00337f
C32183 VPWR.n9027 VGND 0.00524f
C32184 VPWR.n9028 VGND 0.0031f
C32185 VPWR.n9029 VGND 0.00484f
C32186 VPWR.n9030 VGND 0.00624f
C32187 VPWR.n9031 VGND 0.00393f
C32188 VPWR.t1788 VGND 0.0016f
C32189 VPWR.t2421 VGND 0.00208f
C32190 VPWR.n9032 VGND 0.00411f
C32191 VPWR.n9033 VGND 0.0075f
C32192 VPWR.n9034 VGND 0.00366f
C32193 VPWR.n9035 VGND 0.00524f
C32194 VPWR.n9036 VGND 0.0066f
C32195 VPWR.n9037 VGND 0.00524f
C32196 VPWR.t3029 VGND 0.00524f
C32197 VPWR.n9038 VGND 0.00726f
C32198 VPWR.n9039 VGND 0.00334f
C32199 VPWR.n9040 VGND 0.00524f
C32200 VPWR.n9041 VGND 0.00657f
C32201 VPWR.n9042 VGND 0.00524f
C32202 VPWR.n9043 VGND 0.00639f
C32203 VPWR.n9044 VGND 0.00524f
C32204 VPWR.n9045 VGND 0.0031f
C32205 VPWR.n9046 VGND 0.00237f
C32206 VPWR.n9047 VGND 0.0158f
C32207 VPWR.t477 VGND 0.0462f
C32208 VPWR.t2698 VGND 0.0253f
C32209 VPWR.t2700 VGND 0.0198f
C32210 VPWR.t897 VGND 0.0109f
C32211 VPWR.t2087 VGND 0.0052f
C32212 VPWR.t1335 VGND 0.0154f
C32213 VPWR.t2187 VGND 0.0415f
C32214 VPWR.t205 VGND 0.0154f
C32215 VPWR.t1720 VGND 0.0295f
C32216 VPWR.t1334 VGND 0.0386f
C32217 VPWR.t1181 VGND 0.0151f
C32218 VPWR.t2749 VGND 0.0112f
C32219 VPWR.t1209 VGND 0.0331f
C32220 VPWR.t2877 VGND 0.0316f
C32221 VPWR.t873 VGND 0.0166f
C32222 VPWR.t1333 VGND 0.0143f
C32223 VPWR.t3022 VGND 0.0144f
C32224 VPWR.t1719 VGND 0.0144f
C32225 VPWR.t849 VGND 0.0141f
C32226 VPWR.t2110 VGND 0.0211f
C32227 VPWR.t3117 VGND 0.0205f
C32228 VPWR.t1964 VGND 0.0502f
C32229 VPWR.t2108 VGND 0.0364f
C32230 VPWR.t63 VGND 0.021f
C32231 VPWR.t2424 VGND 0.0405f
C32232 VPWR.t2422 VGND 0.0196f
C32233 VPWR.n9048 VGND 0.0192f
C32234 VPWR.t1352 VGND 0.025f
C32235 VPWR.t1548 VGND 0.0453f
C32236 VPWR.t3028 VGND 0.047f
C32237 VPWR.t2420 VGND 0.0312f
C32238 VPWR.t1787 VGND 0.0158f
C32239 VPWR.t344 VGND 0.0206f
C32240 VPWR.t2102 VGND 0.025f
C32241 VPWR.t1665 VGND 0.0589f
C32242 VPWR.t895 VGND 0.0522f
C32243 VPWR.t2053 VGND 0.0247f
C32244 VPWR.t1663 VGND 0.0401f
C32245 VPWR.t1626 VGND 0.0398f
C32246 VPWR.t1361 VGND 0.0396f
C32247 VPWR.t680 VGND 0.0331f
C32248 VPWR.t1723 VGND 0.0264f
C32249 VPWR.t1664 VGND 0.0311f
C32250 VPWR.t2054 VGND 0.0285f
C32251 VPWR.t2492 VGND 0.0322f
C32252 VPWR.t1359 VGND 0.0322f
C32253 VPWR.t1447 VGND 0.0245f
C32254 VPWR.t2490 VGND 0.0492f
C32255 VPWR.n9049 VGND 0.0396f
C32256 VPWR.n9050 VGND 0.0143f
C32257 VPWR.n9051 VGND 0.00796f
C32258 VPWR.n9052 VGND 0.0031f
C32259 VPWR.n9053 VGND 0.0179f
C32260 VPWR.n9054 VGND 0.00524f
C32261 VPWR.n9055 VGND 0.0185f
C32262 VPWR.n9056 VGND 0.00524f
C32263 VPWR.t3484 VGND 0.0592f
C32264 VPWR.n9057 VGND 0.0416f
C32265 VPWR.n9058 VGND 0.0136f
C32266 VPWR.n9059 VGND 0.00524f
C32267 VPWR.t3531 VGND 0.0231f
C32268 VPWR.n9060 VGND 0.00696f
C32269 VPWR.n9061 VGND 0.00121f
C32270 VPWR.t575 VGND 0.00387f
C32271 VPWR.n9062 VGND 0.0026f
C32272 VPWR.n9063 VGND 0.00864f
C32273 VPWR.n9064 VGND 0.0381f
C32274 VPWR.n9065 VGND 0.00492f
C32275 VPWR.n9066 VGND 0.00256f
C32276 VPWR.n9067 VGND 3.14e-19
C32277 VPWR.n9068 VGND 2.28e-19
C32278 VPWR.n9069 VGND 5.98e-19
C32279 VPWR.n9070 VGND 5.12e-19
C32280 VPWR.n9071 VGND 3.13e-19
C32281 VPWR.n9072 VGND 1.77e-19
C32282 VPWR.n9073 VGND 8.67e-19
C32283 VPWR.n9074 VGND 6.54e-19
C32284 VPWR.n9075 VGND 9.06e-19
C32285 VPWR.n9076 VGND 0.00138f
C32286 VPWR.n9077 VGND 5.48e-19
C32287 VPWR.n9078 VGND 1.76e-19
C32288 VPWR.n9079 VGND 5.05e-19
C32289 VPWR.n9080 VGND 7.68e-19
C32290 VPWR.n9081 VGND 3.95e-19
C32291 VPWR.n9082 VGND 6.83e-19
C32292 VPWR.n9083 VGND 2.28e-19
C32293 VPWR.n9084 VGND 4.84e-19
C32294 VPWR.n9085 VGND 0.00562f
C32295 VPWR.n9086 VGND 3.13e-19
C32296 VPWR.n9087 VGND 5.12e-19
C32297 VPWR.n9088 VGND 9.68e-19
C32298 VPWR.n9089 VGND 9.96e-19
C32299 VPWR.n9090 VGND 5.41e-19
C32300 VPWR.n9091 VGND 6.55e-19
C32301 VPWR.n9092 VGND 5.05e-19
C32302 VPWR.n9093 VGND 4.83e-19
C32303 VPWR.n9094 VGND 2.85e-19
C32304 VPWR.n9095 VGND 3.95e-19
C32305 VPWR.n9096 VGND 2.85e-19
C32306 VPWR.n9097 VGND 4.11e-19
C32307 VPWR.n9099 VGND 0.0581f
C32308 VPWR.n9100 VGND 0.0976f
C32309 VPWR.n9101 VGND 0.746f
C32310 VPWR.n9102 VGND 0.564f
C32311 VPWR.n9103 VGND 0.0976f
C32312 VPWR.n9104 VGND 0.0452f
C32313 VPWR.n9105 VGND 5.19e-19
C32314 VPWR.n9106 VGND 7.39e-19
C32315 VPWR.n9107 VGND 4.11e-19
C32316 VPWR.n9108 VGND 5.71e-19
C32317 VPWR.n9109 VGND 4.17e-19
C32318 VPWR.n9110 VGND 3.51e-19
C32319 VPWR.n9111 VGND 4.61e-19
C32320 VPWR.n9112 VGND 4.39e-19
C32321 VPWR.n9113 VGND 3.29e-19
C32322 VPWR.n9114 VGND 5.27e-19
C32323 VPWR.n9115 VGND 2.85e-19
C32324 VPWR.n9116 VGND 2.85e-19
C32325 VPWR.n9117 VGND 4.17e-19
C32326 VPWR.n9118 VGND 6.54e-19
C32327 VPWR.n9119 VGND 8.67e-19
C32328 VPWR.n9120 VGND 4.11e-19
C32329 VPWR.n9122 VGND 0.0057f
C32330 VPWR.n9123 VGND 0.00138f
C32331 VPWR.n9124 VGND 9.06e-19
C32332 VPWR.n9125 VGND 5.48e-19
C32333 VPWR.n9126 VGND 3.07e-19
C32334 VPWR.n9127 VGND 0.00138f
C32335 VPWR.n9128 VGND 0.00407f
C32336 VPWR.n9129 VGND 0.00464f
C32337 VPWR.n9130 VGND 0.00179f
C32338 VPWR.n9131 VGND 0.00306f
C32339 VPWR.n9132 VGND 0.00368f
C32340 VPWR.t3512 VGND 0.0289f
C32341 VPWR.t452 VGND 0.00387f
C32342 VPWR.n9133 VGND 0.0604f
C32343 VPWR.n9134 VGND 0.0116f
C32344 VPWR.n9135 VGND 0.0117f
C32345 VPWR.t2649 VGND 0.00676f
C32346 VPWR.t1631 VGND 0.00234f
C32347 VPWR.n9136 VGND 0.00258f
C32348 VPWR.n9137 VGND 0.0125f
C32349 VPWR.t673 VGND 0.00399f
C32350 VPWR.n9138 VGND 0.00181f
C32351 VPWR.n9139 VGND 0.0193f
C32352 VPWR.n9140 VGND 0.0116f
C32353 VPWR.n9141 VGND 0.00333f
C32354 VPWR.n9142 VGND 0.00393f
C32355 VPWR.n9143 VGND 0.00199f
C32356 VPWR.n9144 VGND 0.0132f
C32357 VPWR.n9145 VGND 0.00513f
C32358 VPWR.n9146 VGND 0.0031f
C32359 VPWR.n9147 VGND 0.00524f
C32360 VPWR.n9148 VGND 0.00524f
C32361 VPWR.n9149 VGND 0.0114f
C32362 VPWR.n9150 VGND 0.00524f
C32363 VPWR.t3549 VGND 0.0231f
C32364 VPWR.t564 VGND 0.00387f
C32365 VPWR.n9151 VGND 0.00837f
C32366 VPWR.n9152 VGND 0.0384f
C32367 VPWR.n9153 VGND 0.00393f
C32368 VPWR.n9154 VGND 0.00202f
C32369 VPWR.n9155 VGND 0.00179f
C32370 VPWR.n9156 VGND 0.00173f
C32371 VPWR.n9157 VGND 0.0015f
C32372 VPWR.n9158 VGND 0.0031f
C32373 VPWR.n9159 VGND 0.00524f
C32374 VPWR.n9160 VGND 0.00393f
C32375 VPWR.n9161 VGND 0.00141f
C32376 VPWR.n9162 VGND 0.00525f
C32377 VPWR.n9163 VGND 0.0031f
C32378 VPWR.n9164 VGND 0.00524f
C32379 VPWR.n9165 VGND 0.00524f
C32380 VPWR.n9166 VGND 0.00393f
C32381 VPWR.n9167 VGND 0.00525f
C32382 VPWR.n9168 VGND 0.00173f
C32383 VPWR.n9169 VGND 0.00199f
C32384 VPWR.n9170 VGND 0.00142f
C32385 VPWR.n9171 VGND 0.0031f
C32386 VPWR.t1981 VGND 0.00136f
C32387 VPWR.t2245 VGND 0.00136f
C32388 VPWR.n9172 VGND 0.00317f
C32389 VPWR.t3116 VGND 6.73e-19
C32390 VPWR.t3196 VGND 9.96e-19
C32391 VPWR.n9173 VGND 0.00176f
C32392 VPWR.n9174 VGND 0.00421f
C32393 VPWR.n9175 VGND 0.00686f
C32394 VPWR.n9176 VGND 0.00524f
C32395 VPWR.n9177 VGND 0.00393f
C32396 VPWR.n9178 VGND 0.00132f
C32397 VPWR.t1206 VGND 0.00454f
C32398 VPWR.n9179 VGND 0.00798f
C32399 VPWR.n9180 VGND 0.00236f
C32400 VPWR.n9181 VGND 0.0031f
C32401 VPWR.n9182 VGND 0.00524f
C32402 VPWR.n9183 VGND 0.00524f
C32403 VPWR.n9184 VGND 0.00393f
C32404 VPWR.n9185 VGND 0.00509f
C32405 VPWR.n9186 VGND 0.00347f
C32406 VPWR.n9187 VGND 1.51e-19
C32407 VPWR.n9188 VGND 0.0031f
C32408 VPWR.n9189 VGND 0.00148f
C32409 VPWR.n9190 VGND 0.00524f
C32410 VPWR.n9191 VGND 0.00393f
C32411 VPWR.n9192 VGND 8.39e-19
C32412 VPWR.n9193 VGND 0.0051f
C32413 VPWR.n9194 VGND 0.00908f
C32414 VPWR.n9195 VGND 0.00807f
C32415 VPWR.n9196 VGND 0.0133f
C32416 VPWR.n9197 VGND 0.00393f
C32417 VPWR.n9198 VGND 0.00199f
C32418 VPWR.n9199 VGND 0.00199f
C32419 VPWR.n9200 VGND 0.0113f
C32420 VPWR.t3438 VGND 0.0289f
C32421 VPWR.t241 VGND 0.00387f
C32422 VPWR.n9201 VGND 0.0604f
C32423 VPWR.n9202 VGND 0.0146f
C32424 VPWR.n9203 VGND 0.0117f
C32425 VPWR.n9204 VGND 0.0173f
C32426 VPWR.n9205 VGND 6.35e-19
C32427 VPWR.n9206 VGND 6.26e-19
C32428 VPWR.n9207 VGND 3.14e-19
C32429 VPWR.n9208 VGND 1.71e-19
C32430 VPWR.n9209 VGND 2.28e-19
C32431 VPWR.n9210 VGND 9.28e-19
C32432 VPWR.n9211 VGND 5.98e-19
C32433 VPWR.n9212 VGND 5.12e-19
C32434 VPWR.n9213 VGND 3.13e-19
C32435 VPWR.n9214 VGND 1.76e-19
C32436 VPWR.n9215 VGND 1.76e-19
C32437 VPWR.n9216 VGND 5.05e-19
C32438 VPWR.n9217 VGND 7.68e-19
C32439 VPWR.n9218 VGND 3.95e-19
C32440 VPWR.n9219 VGND 5.12e-19
C32441 VPWR.n9220 VGND 6.26e-19
C32442 VPWR.n9221 VGND 0.00162f
C32443 VPWR.n9222 VGND 3.13e-19
C32444 VPWR.n9223 VGND 5.12e-19
C32445 VPWR.n9224 VGND 9.68e-19
C32446 VPWR.n9225 VGND 9.96e-19
C32447 VPWR.n9226 VGND 5.41e-19
C32448 VPWR.n9227 VGND 3.95e-19
C32449 VPWR.n9228 VGND 4.83e-19
C32450 VPWR.n9229 VGND 2.41e-19
C32451 VPWR.n9230 VGND 3.73e-19
C32452 VPWR.n9231 VGND 4.17e-19
C32453 VPWR.n9232 VGND 2.85e-19
C32454 VPWR.n9233 VGND 4.83e-19
C32455 VPWR.n9234 VGND 2.85e-19
C32456 VPWR.n9235 VGND 3.95e-19
C32457 VPWR.n9236 VGND 2.85e-19
C32458 VPWR.n9237 VGND 4.11e-19
C32459 VPWR.n9238 VGND 4.11e-19
C32460 VPWR.n9239 VGND 7.39e-19
C32461 VPWR.n9240 VGND 5.19e-19
C32462 VPWR.n9241 VGND 7.39e-19
C32463 VPWR.n9242 VGND 4.11e-19
C32464 VPWR.n9243 VGND 8.67e-19
C32465 VPWR.n9244 VGND 4.11e-19
C32466 VPWR.n9245 VGND 3.07e-19
C32467 VPWR.n9246 VGND 1.76e-19
C32468 VPWR.n9247 VGND 4.39e-19
C32469 VPWR.n9248 VGND 6.14e-19
C32470 VPWR.n9249 VGND 4.17e-19
C32471 VPWR.n9250 VGND 5.05e-19
C32472 VPWR.n9251 VGND 6.55e-19
C32473 VPWR.n9252 VGND 6.26e-19
C32474 VPWR.n9253 VGND 5.85e-19
C32475 VPWR.t2502 VGND 0.00166f
C32476 VPWR.t3102 VGND 0.00184f
C32477 VPWR.n9254 VGND 0.00362f
C32478 VPWR.n9255 VGND 0.00389f
C32479 VPWR.n9256 VGND 3.1e-19
C32480 VPWR.n9257 VGND 7.27e-19
C32481 VPWR.n9258 VGND 5.41e-19
C32482 VPWR.n9259 VGND 5.12e-19
C32483 VPWR.n9260 VGND 4.27e-19
C32484 VPWR.n9261 VGND 2.85e-19
C32485 VPWR.n9262 VGND 0.00125f
C32486 VPWR.n9263 VGND 5.98e-19
C32487 VPWR.n9264 VGND 6.99e-19
C32488 VPWR.n9265 VGND 0.00169f
C32489 VPWR.n9266 VGND 0.00138f
C32490 VPWR.n9267 VGND 3.95e-19
C32491 VPWR.n9268 VGND 3.29e-19
C32492 VPWR.n9269 VGND 5.71e-19
C32493 VPWR.n9270 VGND 5.92e-19
C32494 VPWR.n9271 VGND 5.05e-19
C32495 VPWR.n9272 VGND 4.17e-19
C32496 VPWR.n9273 VGND 8.67e-19
C32497 VPWR.n9274 VGND 6.54e-19
C32498 VPWR.n9275 VGND 9.06e-19
C32499 VPWR.n9276 VGND 5.48e-19
C32500 VPWR.n9277 VGND 0.00138f
C32501 VPWR.n9278 VGND 0.0057f
C32502 VPWR.n9280 VGND 0.1f
C32503 VPWR.n9281 VGND 0.1f
C32504 VPWR.n9283 VGND 0.00139f
C32505 VPWR.n9284 VGND 5.48e-19
C32506 VPWR.n9285 VGND 1.76e-19
C32507 VPWR.n9286 VGND 8.11e-19
C32508 VPWR.n9287 VGND 3.95e-19
C32509 VPWR.n9288 VGND 1.76e-19
C32510 VPWR.n9289 VGND 3.13e-19
C32511 VPWR.n9290 VGND 6.26e-19
.ends

