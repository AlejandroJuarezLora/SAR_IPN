magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 774 542
<< pwell >>
rect 1 -19 735 163
rect 30 -57 64 -19
<< scnmos >>
rect 93 7 123 137
rect 226 7 256 137
rect 316 7 346 137
rect 436 7 466 137
rect 554 7 584 137
rect 626 7 656 137
<< scpmoshvt >>
rect 93 257 123 457
rect 220 257 250 457
rect 316 257 346 457
rect 436 257 466 457
rect 540 257 570 457
rect 626 257 656 457
<< ndiff >>
rect 27 122 93 137
rect 27 88 35 122
rect 69 88 93 122
rect 27 54 93 88
rect 27 20 35 54
rect 69 20 93 54
rect 27 7 93 20
rect 123 57 226 137
rect 123 23 135 57
rect 169 23 226 57
rect 123 7 226 23
rect 256 7 316 137
rect 346 7 436 137
rect 466 57 554 137
rect 466 23 492 57
rect 526 23 554 57
rect 466 7 554 23
rect 584 7 626 137
rect 656 121 709 137
rect 656 87 667 121
rect 701 87 709 121
rect 656 53 709 87
rect 656 19 667 53
rect 701 19 709 53
rect 656 7 709 19
<< pdiff >>
rect 27 445 93 457
rect 27 411 35 445
rect 69 411 93 445
rect 27 377 93 411
rect 27 343 35 377
rect 69 343 93 377
rect 27 309 93 343
rect 27 275 35 309
rect 69 275 93 309
rect 27 257 93 275
rect 123 445 220 457
rect 123 411 151 445
rect 185 411 220 445
rect 123 377 220 411
rect 123 343 151 377
rect 185 343 220 377
rect 123 257 220 343
rect 250 437 316 457
rect 250 403 266 437
rect 300 403 316 437
rect 250 369 316 403
rect 250 335 266 369
rect 300 335 316 369
rect 250 257 316 335
rect 346 445 436 457
rect 346 411 374 445
rect 408 411 436 445
rect 346 257 436 411
rect 466 445 540 457
rect 466 411 485 445
rect 519 411 540 445
rect 466 377 540 411
rect 466 343 485 377
rect 519 343 540 377
rect 466 257 540 343
rect 570 369 626 457
rect 570 335 581 369
rect 615 335 626 369
rect 570 257 626 335
rect 656 437 709 457
rect 656 403 667 437
rect 701 403 709 437
rect 656 369 709 403
rect 656 335 667 369
rect 701 335 709 369
rect 656 257 709 335
<< ndiffc >>
rect 35 88 69 122
rect 35 20 69 54
rect 135 23 169 57
rect 492 23 526 57
rect 667 87 701 121
rect 667 19 701 53
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 35 275 69 309
rect 151 411 185 445
rect 151 343 185 377
rect 266 403 300 437
rect 266 335 300 369
rect 374 411 408 445
rect 485 411 519 445
rect 485 343 519 377
rect 581 335 615 369
rect 667 403 701 437
rect 667 335 701 369
<< poly >>
rect 93 457 123 483
rect 220 457 250 483
rect 316 457 346 483
rect 436 457 466 483
rect 540 457 570 483
rect 626 457 656 483
rect 93 225 123 257
rect 220 225 250 257
rect 316 225 346 257
rect 436 225 466 257
rect 540 225 570 257
rect 626 225 656 257
rect 93 209 158 225
rect 93 175 114 209
rect 148 175 158 209
rect 93 159 158 175
rect 220 209 274 225
rect 220 175 230 209
rect 264 175 274 209
rect 220 159 274 175
rect 316 209 370 225
rect 316 175 326 209
rect 360 175 370 209
rect 316 159 370 175
rect 412 209 466 225
rect 412 175 422 209
rect 456 175 466 209
rect 412 159 466 175
rect 530 209 584 225
rect 530 175 540 209
rect 574 175 584 209
rect 530 159 584 175
rect 93 137 123 159
rect 226 137 256 159
rect 316 137 346 159
rect 436 137 466 159
rect 554 137 584 159
rect 626 209 680 225
rect 626 175 636 209
rect 670 175 680 209
rect 626 159 680 175
rect 626 137 656 159
rect 93 -19 123 7
rect 226 -19 256 7
rect 316 -19 346 7
rect 436 -19 466 7
rect 554 -19 584 7
rect 626 -19 656 7
<< polycont >>
rect 114 175 148 209
rect 230 175 264 209
rect 326 175 360 209
rect 422 175 456 209
rect 540 175 574 209
rect 636 175 670 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 135 445 201 487
rect 18 411 35 445
rect 69 411 85 445
rect 18 377 85 411
rect 18 343 35 377
rect 69 343 85 377
rect 135 411 151 445
rect 185 411 201 445
rect 135 377 201 411
rect 135 343 151 377
rect 185 343 201 377
rect 18 309 69 343
rect 135 327 201 343
rect 250 437 307 453
rect 250 403 266 437
rect 300 403 307 437
rect 358 445 424 487
rect 358 411 374 445
rect 408 411 424 445
rect 358 403 424 411
rect 469 445 701 453
rect 469 411 485 445
rect 519 437 701 445
rect 519 419 667 437
rect 519 411 535 419
rect 250 369 307 403
rect 469 377 535 411
rect 469 369 485 377
rect 250 335 266 369
rect 300 343 485 369
rect 519 343 535 377
rect 300 335 535 343
rect 581 369 615 385
rect 18 275 35 309
rect 581 293 615 335
rect 667 369 701 403
rect 667 319 701 335
rect 18 122 69 275
rect 141 259 615 293
rect 141 225 175 259
rect 665 225 706 283
rect 114 209 175 225
rect 148 175 175 209
rect 114 159 175 175
rect 214 209 264 225
rect 214 175 230 209
rect 214 159 264 175
rect 306 209 360 225
rect 306 175 326 209
rect 18 88 35 122
rect 141 125 175 159
rect 141 91 253 125
rect 306 93 360 175
rect 398 209 456 225
rect 398 175 422 209
rect 398 93 456 175
rect 490 209 574 225
rect 490 175 540 209
rect 490 92 574 175
rect 636 209 706 225
rect 670 175 706 209
rect 636 159 706 175
rect 18 72 69 88
rect 18 54 85 72
rect 219 57 253 91
rect 651 87 667 121
rect 701 87 717 121
rect 18 20 35 54
rect 69 20 85 54
rect 119 23 135 57
rect 169 23 185 57
rect 219 23 492 57
rect 526 23 542 57
rect 651 53 717 87
rect 119 -23 185 23
rect 651 19 667 53
rect 701 19 717 53
rect 651 -23 717 19
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
<< metal1 >>
rect 0 521 736 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 0 456 736 487
rect 0 -23 736 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
rect 0 -88 736 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 a32o_1
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 30 45 64 79 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 30 113 64 147 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 30 249 64 283 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 30 317 64 351 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 30 385 64 419 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 214 181 248 215 0 FreeSans 200 0 0 0 A3
port 8 nsew
flabel locali s 672 181 706 215 0 FreeSans 200 0 0 0 B2
port 12 nsew
flabel locali s 490 113 524 147 0 FreeSans 200 0 0 0 B1
port 11 nsew
flabel locali s 398 113 432 147 0 FreeSans 200 0 0 0 A1
port 10 nsew
flabel locali s 398 181 432 215 0 FreeSans 200 0 0 0 A1
port 10 nsew
flabel locali s 306 181 340 215 0 FreeSans 200 0 0 0 A2
port 9 nsew
flabel locali s 490 181 524 215 0 FreeSans 200 0 0 0 B1
port 11 nsew
flabel locali s 672 249 706 283 0 FreeSans 200 0 0 0 B2
port 12 nsew
flabel locali s 306 113 340 147 0 FreeSans 200 0 0 0 A2
port 9 nsew
flabel locali s 30 181 64 215 0 FreeSans 200 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 736 504
string path 0.000 -1.000 18.400 -1.000 
<< end >>
