magic
tech sky130B
timestamp 1696364841
<< metal3 >>
rect 0 16 80 20
rect 0 -16 4 16
rect 36 -16 44 16
rect 76 -16 80 16
rect 0 -20 80 -16
<< via3 >>
rect 4 -16 36 16
rect 44 -16 76 16
<< metal4 >>
rect 0 16 80 20
rect 0 -16 4 16
rect 36 -16 44 16
rect 76 -16 80 16
rect 0 -20 80 -16
<< end >>
