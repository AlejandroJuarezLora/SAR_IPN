magic
tech sky130B
timestamp 1696364841
<< metal1 >>
rect 0 -17 3 9
rect 29 -17 32 9
<< via1 >>
rect 3 -17 29 9
<< metal2 >>
rect 3 9 29 12
rect 3 -20 29 -17
<< end >>
