magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 130 542
<< pwell >>
rect 3 -2 89 155
<< psubdiff >>
rect 29 105 63 129
rect 29 24 63 71
<< nsubdiff >>
rect 29 416 63 440
rect 29 323 63 382
rect 29 265 63 289
<< psubdiffcont >>
rect 29 71 63 105
<< nsubdiffcont >>
rect 29 382 63 416
rect 29 289 63 323
<< locali >>
rect 0 487 29 521
rect 63 487 92 521
rect 17 416 75 487
rect 17 382 29 416
rect 63 382 75 416
rect 17 323 75 382
rect 17 289 29 323
rect 63 289 75 323
rect 17 254 75 289
rect 17 105 75 122
rect 17 71 29 105
rect 63 71 75 105
rect 17 -23 75 71
rect 0 -57 29 -23
rect 63 -57 92 -23
<< viali >>
rect 29 487 63 521
rect 29 -57 63 -23
<< metal1 >>
rect 0 521 92 552
rect 0 487 29 521
rect 63 487 92 521
rect 0 456 92 487
rect 0 -23 92 8
rect 0 -57 29 -23
rect 63 -57 92 -23
rect 0 -88 92 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 tapvpwrvgnd_1
flabel metal1 s 22 484 75 513 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 21 -58 72 -20 0 FreeSans 200 0 0 0 VGND
port 3 nsew
<< properties >>
string FIXED_BBOX 0 -40 92 504
<< end >>
