magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_s >>
rect 312 2937 2484 3023
rect 312 2433 398 2937
rect 2398 2433 2484 2937
rect 312 2347 2484 2433
<< nwell >>
rect 302 2337 2494 3033
<< metal1 >>
rect 591 2802 637 3206
rect 962 2957 1008 3214
rect 1380 2802 1426 3206
rect 1806 2957 1852 3214
rect 2159 2802 2205 3206
rect 213 2679 519 2725
rect 213 872 259 2679
rect 709 2670 1308 2730
rect 1498 2670 2087 2730
rect 2277 2679 2591 2725
rect 526 2515 710 2561
rect 1202 2515 1373 2561
rect 1433 2515 1602 2561
rect 2094 2515 2278 2561
rect 591 1794 637 2515
rect 1202 2219 1248 2515
rect 1556 2166 1602 2515
rect 1042 1997 1602 2043
rect 1042 1888 1088 1997
rect 1556 1936 1602 1997
rect 1014 1842 1088 1888
rect 1716 1842 1790 1888
rect 366 1748 637 1794
rect 366 1053 412 1748
rect 1202 1735 1248 1796
rect 1716 1735 1762 1842
rect 2161 1794 2207 2515
rect 2161 1748 2438 1794
rect 1202 1689 1762 1735
rect 575 1526 1366 1572
rect 1320 1282 1366 1526
rect 1438 1526 2229 1572
rect 1438 1282 1484 1526
rect 975 1050 1143 1190
rect 1261 872 1307 1096
rect 213 826 1307 872
rect 1379 620 1425 1096
rect 1497 872 1543 1096
rect 1661 1050 1829 1190
rect 2392 1053 2438 1748
rect 2545 872 2591 2679
rect 1497 826 2591 872
rect 366 388 412 530
rect 1156 450 1261 590
rect 1543 450 1648 590
rect 2392 388 2438 530
rect 366 342 2438 388
rect 1372 -40 1432 342
<< metal2 >>
rect 554 3151 2242 3231
rect 905 1905 985 2640
rect 1195 1926 1255 2311
rect 1549 1926 1609 2311
rect 1819 1905 1899 2640
rect 349 467 429 1180
rect 905 -40 985 1825
rect 1195 1398 1255 1834
rect 1549 1449 1609 1834
rect 1087 308 1167 981
rect 1637 308 1717 981
rect 1087 228 1717 308
rect 1362 -40 1442 228
rect 1819 -40 1899 1825
rect 2375 467 2455 1180
<< metal4 >>
rect 1152 3431 1252 3481
rect 0 3331 1252 3431
rect 1552 3431 1652 3481
rect 1552 3331 2804 3431
rect 0 1599 100 3331
rect 2704 1599 2804 3331
rect 0 1499 748 1599
rect 2056 1499 2804 1599
use gr_contact  gr_contact_0
timestamp 1696364841
transform 0 1 1698 -1 0 3003
box 0 -40 46 295
use gr_contact  gr_contact_1
timestamp 1696364841
transform 0 1 854 -1 0 3003
box 0 -40 46 295
use Guardring_N_1  Guardring_N_1_0
timestamp 1696364841
transform 1 0 -7046 0 1 -886
box 8130 1111 8766 1662
use Guardring_N_4  Guardring_N_4_0
timestamp 1696364841
transform 1 0 -7046 0 1 -886
box 8032 1784 8864 2350
use M1  M1_0
timestamp 1696364841
transform 1 0 555 0 -1 2626
box -124 -238 124 124
use M2  M2_0
timestamp 1696364841
transform 1 0 673 0 -1 2626
box -124 -238 124 124
use M3  M3_0
timestamp 1696364841
transform 1 0 2123 0 -1 2626
box -124 -238 124 124
use M4  M4_0
timestamp 1696364841
transform 1 0 2241 0 -1 2626
box -124 -238 124 124
use Mdiff  Mdiff_0
timestamp 1696364841
transform 1 0 1461 0 -1 449
box -114 -197 114 117
use Mdiff  Mdiff_1
timestamp 1696364841
transform 1 0 1343 0 -1 449
box -114 -197 114 117
use Minn  Minn_0
timestamp 1696364841
transform 1 0 1343 0 1 1221
box -114 -197 114 117
use Minp  Minp_0
timestamp 1696364841
transform 1 0 1461 0 1 1221
box -114 -197 114 117
use Ml1  Ml1_0
timestamp 1696364841
transform -1 0 1225 0 1 1221
box -114 -197 114 117
use Ml2  Ml2_0
timestamp 1696364841
transform -1 0 1579 0 1 1221
box -114 -197 114 117
use Ml3  Ml3_0
timestamp 1696364841
transform 1 0 1344 0 -1 2626
box -124 -238 124 124
use Ml4  Ml4_0
timestamp 1696364841
transform 1 0 1462 0 -1 2626
box -124 -238 124 124
use pguard  pguard_0
timestamp 1696364841
transform 1 0 1398 0 1 2725
box -1096 -388 1096 308
use via1_2  via1_2_0
timestamp 1696364841
transform 1 0 1068 0 1 958
box -6 -46 124 12
use via1_2  via1_2_1
timestamp 1696364841
transform 0 -1 1660 1 0 461
box -6 -46 124 12
use via1_2  via1_2_2
timestamp 1696364841
transform 0 -1 1110 1 0 461
box -6 -46 124 12
use via1_2  via1_2_3
timestamp 1696364841
transform 1 0 1618 0 1 958
box -6 -46 124 12
use via2_1  via2_1_0
timestamp 1696364841
transform 0 -1 389 -1 0 1190
box 0 -40 140 40
use via2_1  via2_1_1
timestamp 1696364841
transform 0 -1 389 -1 0 597
box 0 -40 140 40
use via2_1  via2_1_2
timestamp 1696364841
transform 0 1 2415 -1 0 1190
box 0 -40 140 40
use via2_1  via2_1_3
timestamp 1696364841
transform 0 1 2415 -1 0 597
box 0 -40 140 40
use via2_1  via2_1_4
timestamp 1696364841
transform -1 0 2229 0 -1 1549
box 0 -40 140 40
use via2_1  via2_1_5
timestamp 1696364841
transform 1 0 575 0 -1 1549
box 0 -40 140 40
use via2_1  via2_1_6
timestamp 1696364841
transform -1 0 1197 0 1 941
box 0 -40 140 40
use via2_1  via2_1_7
timestamp 1696364841
transform 0 1 1677 -1 0 590
box 0 -40 140 40
use via2_1  via2_1_8
timestamp 1696364841
transform 0 -1 1127 -1 0 590
box 0 -40 140 40
use via2_1  via2_1_9
timestamp 1696364841
transform 0 1 1859 -1 0 1190
box 0 -40 140 40
use via2_1  via2_1_10
timestamp 1696364841
transform 0 -1 945 -1 0 1190
box 0 -40 140 40
use via2_1  via2_1_11
timestamp 1696364841
transform -1 0 1930 0 -1 1865
box 0 -40 140 40
use via2_1  via2_1_12
timestamp 1696364841
transform -1 0 1014 0 -1 1865
box 0 -40 140 40
use via2_1  via2_1_13
timestamp 1696364841
transform 0 -1 1225 1 0 1796
box 0 -40 140 40
use via2_1  via2_1_14
timestamp 1696364841
transform 0 -1 1579 1 0 1796
box 0 -40 140 40
use via2_1  via2_1_15
timestamp 1696364841
transform 0 1 1225 -1 0 1468
box 0 -40 140 40
use via2_1  via2_1_16
timestamp 1696364841
transform 0 1 1579 -1 0 1468
box 0 -40 140 40
use via2_1  via2_1_17
timestamp 1696364841
transform 0 -1 1225 1 0 2171
box 0 -40 140 40
use via2_1  via2_1_18
timestamp 1696364841
transform 0 -1 1579 1 0 2171
box 0 -40 140 40
use via2_1  via2_1_19
timestamp 1696364841
transform 0 -1 945 1 0 2630
box 0 -40 140 40
use via2_1  via2_1_20
timestamp 1696364841
transform 0 1 1859 1 0 2630
box 0 -40 140 40
use via2_1  via2_1_21
timestamp 1696364841
transform 1 0 1333 0 1 3191
box 0 -40 140 40
use via2_1  via2_1_22
timestamp 1696364841
transform -1 0 1747 0 -1 941
box 0 -40 140 40
use via2_1  via2_1_23
timestamp 1696364841
transform 1 0 544 0 1 3191
box 0 -40 140 40
use via2_1  via2_1_24
timestamp 1696364841
transform 1 0 2112 0 1 3191
box 0 -40 140 40
use via2_1  via2_1_25
timestamp 1696364841
transform 1 0 1759 0 1 3191
box 0 -40 140 40
use via2_1  via2_1_26
timestamp 1696364841
transform 1 0 915 0 1 3191
box 0 -40 140 40
use via23_2  via23_2_0
timestamp 1696364841
transform -1 0 2240 0 -1 1629
box 1 40 161 120
use via23_2  via23_2_1
timestamp 1696364841
transform -1 0 726 0 -1 1629
box 1 40 161 120
use via34  via34_0
timestamp 1696364841
transform -1 0 755 0 -1 1589
box 9 -8 211 88
use via34  via34_1
timestamp 1696364841
transform -1 0 2269 0 -1 1589
box 9 -8 211 88
<< labels >>
flabel metal2 s 554 3151 594 3231 2 FreeSans 44 0 0 0 vdd
port 2 nsew
flabel metal2 s 1362 -40 1442 0 2 FreeSans 44 0 0 0 vss
port 3 nsew
flabel metal2 s 1819 -40 1899 0 2 FreeSans 44 0 0 0 outp
port 4 nsew
flabel metal2 s 905 -40 985 0 2 FreeSans 44 0 0 0 outn
port 5 nsew
flabel metal1 s 1372 -40 1432 -10 2 FreeSans 44 0 0 0 clk
port 7 nsew
flabel metal1 s 1497 826 1543 872 1 FreeSans 44 0 0 0 ip
port 8 nsew
flabel metal1 s 1261 826 1307 872 1 FreeSans 44 0 0 0 in
port 9 nsew
flabel metal1 s 1379 826 1425 872 1 FreeSans 44 0 0 0 diff
port 10 nsew
flabel metal4 s 1552 3431 1652 3481 2 FreeSans 96 0 0 0 vp
port 12 nsew
flabel metal4 s 1152 3431 1252 3481 2 FreeSans 96 0 0 0 vn
port 13 nsew
<< properties >>
string FIXED_BBOX 0 -40 2804 3481
string path 17.450 38.725 1.250 38.725 1.250 84.525 
<< end >>
