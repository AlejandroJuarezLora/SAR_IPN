magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 866 542
<< pwell >>
rect 31 -19 762 163
rect 31 -23 63 -19
rect 29 -57 63 -23
<< scnmos >>
rect 119 7 149 137
rect 210 7 240 137
rect 294 7 324 137
rect 482 7 512 137
rect 566 7 596 137
rect 650 7 680 137
<< scpmoshvt >>
rect 119 257 149 457
rect 215 257 245 457
rect 287 257 317 457
rect 482 257 512 457
rect 554 257 584 457
rect 650 257 680 457
<< ndiff >>
rect 57 123 119 137
rect 57 89 65 123
rect 99 89 119 123
rect 57 55 119 89
rect 57 21 65 55
rect 99 21 119 55
rect 57 7 119 21
rect 149 55 210 137
rect 149 21 165 55
rect 199 21 210 55
rect 149 7 210 21
rect 240 123 294 137
rect 240 89 250 123
rect 284 89 294 123
rect 240 7 294 89
rect 324 55 376 137
rect 324 21 334 55
rect 368 21 376 55
rect 324 7 376 21
rect 430 55 482 137
rect 430 21 438 55
rect 472 21 482 55
rect 430 7 482 21
rect 512 123 566 137
rect 512 89 522 123
rect 556 89 566 123
rect 512 55 566 89
rect 512 21 522 55
rect 556 21 566 55
rect 512 7 566 21
rect 596 123 650 137
rect 596 89 606 123
rect 640 89 650 123
rect 596 55 650 89
rect 596 21 606 55
rect 640 21 650 55
rect 596 7 650 21
rect 680 123 736 137
rect 680 89 690 123
rect 724 89 736 123
rect 680 55 736 89
rect 680 21 690 55
rect 724 21 736 55
rect 680 7 736 21
<< pdiff >>
rect 51 437 119 457
rect 51 403 74 437
rect 108 403 119 437
rect 51 369 119 403
rect 51 335 74 369
rect 108 335 119 369
rect 51 301 119 335
rect 51 267 74 301
rect 108 267 119 301
rect 51 257 119 267
rect 149 437 215 457
rect 149 403 163 437
rect 197 403 215 437
rect 149 369 215 403
rect 149 335 163 369
rect 197 335 215 369
rect 149 257 215 335
rect 245 257 287 457
rect 317 437 482 457
rect 317 403 327 437
rect 361 403 438 437
rect 472 403 482 437
rect 317 369 482 403
rect 317 335 327 369
rect 361 335 438 369
rect 472 335 482 369
rect 317 257 482 335
rect 512 257 554 457
rect 584 437 650 457
rect 584 403 594 437
rect 628 403 650 437
rect 584 369 650 403
rect 584 335 594 369
rect 628 335 650 369
rect 584 257 650 335
rect 680 437 736 457
rect 680 403 694 437
rect 728 403 736 437
rect 680 369 736 403
rect 680 335 694 369
rect 728 335 736 369
rect 680 257 736 335
<< ndiffc >>
rect 65 89 99 123
rect 65 21 99 55
rect 165 21 199 55
rect 250 89 284 123
rect 334 21 368 55
rect 438 21 472 55
rect 522 89 556 123
rect 522 21 556 55
rect 606 89 640 123
rect 606 21 640 55
rect 690 89 724 123
rect 690 21 724 55
<< pdiffc >>
rect 74 403 108 437
rect 74 335 108 369
rect 74 267 108 301
rect 163 403 197 437
rect 163 335 197 369
rect 327 403 361 437
rect 438 403 472 437
rect 327 335 361 369
rect 438 335 472 369
rect 594 403 628 437
rect 594 335 628 369
rect 694 403 728 437
rect 694 335 728 369
<< poly >>
rect 119 457 149 483
rect 215 457 245 483
rect 287 457 317 483
rect 482 457 512 483
rect 554 457 584 483
rect 650 457 680 483
rect 119 225 149 257
rect 215 225 245 257
rect 23 209 149 225
rect 23 175 33 209
rect 67 175 149 209
rect 23 159 149 175
rect 191 209 245 225
rect 191 175 201 209
rect 235 175 245 209
rect 191 159 245 175
rect 287 225 317 257
rect 482 225 512 257
rect 287 209 357 225
rect 287 175 313 209
rect 347 175 357 209
rect 287 159 357 175
rect 438 209 512 225
rect 438 175 448 209
rect 482 175 512 209
rect 438 159 512 175
rect 554 225 584 257
rect 650 225 680 257
rect 554 209 608 225
rect 554 175 564 209
rect 598 175 608 209
rect 554 159 608 175
rect 650 209 721 225
rect 650 175 677 209
rect 711 175 721 209
rect 650 159 721 175
rect 119 137 149 159
rect 210 137 240 159
rect 294 137 324 159
rect 482 137 512 159
rect 566 137 596 159
rect 650 137 680 159
rect 119 -19 149 7
rect 210 -19 240 7
rect 294 -19 324 7
rect 482 -19 512 7
rect 566 -19 596 7
rect 650 -19 680 7
<< polycont >>
rect 33 175 67 209
rect 201 175 235 209
rect 313 175 347 209
rect 448 175 482 209
rect 564 175 598 209
rect 677 175 711 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 828 521
rect 48 437 108 453
rect 48 403 74 437
rect 48 369 108 403
rect 48 335 74 369
rect 48 301 108 335
rect 147 437 197 487
rect 147 403 163 437
rect 147 369 197 403
rect 315 437 476 453
rect 315 403 327 437
rect 361 403 438 437
rect 472 403 476 437
rect 315 369 476 403
rect 578 437 644 487
rect 578 403 594 437
rect 628 403 644 437
rect 578 369 644 403
rect 147 335 163 369
rect 147 319 197 335
rect 231 335 327 369
rect 361 335 438 369
rect 472 335 544 369
rect 48 267 74 301
rect 231 285 265 335
rect 108 267 265 285
rect 48 251 265 267
rect 17 209 83 217
rect 17 175 33 209
rect 67 175 83 209
rect 17 159 83 175
rect 117 125 151 251
rect 299 225 363 301
rect 185 209 251 217
rect 185 175 201 209
rect 235 175 251 209
rect 287 209 363 225
rect 287 175 313 209
rect 347 175 363 209
rect 401 217 476 301
rect 510 285 544 335
rect 578 335 594 369
rect 628 335 644 369
rect 678 437 811 453
rect 678 403 694 437
rect 728 403 811 437
rect 678 369 811 403
rect 678 335 694 369
rect 728 335 811 369
rect 578 319 644 335
rect 510 251 694 285
rect 660 217 694 251
rect 401 209 498 217
rect 401 175 448 209
rect 482 175 498 209
rect 536 209 626 217
rect 536 175 564 209
rect 598 175 626 209
rect 660 209 727 217
rect 660 175 677 209
rect 711 175 727 209
rect 761 141 811 335
rect 49 123 151 125
rect 49 89 65 123
rect 99 89 151 123
rect 232 123 572 141
rect 232 89 250 123
rect 284 107 522 123
rect 284 89 309 107
rect 506 89 522 107
rect 556 89 572 123
rect 49 55 115 89
rect 438 55 472 71
rect 49 21 65 55
rect 99 21 115 55
rect 149 21 165 55
rect 199 21 334 55
rect 368 21 386 55
rect 49 11 115 21
rect 438 -23 472 21
rect 506 55 572 89
rect 506 21 522 55
rect 556 21 572 55
rect 506 14 572 21
rect 606 123 640 141
rect 606 55 640 89
rect 606 -23 640 21
rect 674 123 811 141
rect 674 89 690 123
rect 724 89 811 123
rect 674 55 811 89
rect 674 21 690 55
rect 724 21 811 55
rect 674 13 811 21
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 828 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
<< metal1 >>
rect 0 521 828 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 828 521
rect 0 456 828 487
rect 0 -23 828 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 828 -23
rect 0 -88 828 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 o221a_1
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 401 181 435 215 0 FreeSans 400 0 0 0 A2
port 9 nsew
flabel locali s 765 317 799 351 0 FreeSans 400 0 0 0 X
port 11 nsew
flabel locali s 213 181 247 215 0 FreeSans 400 0 0 0 B1
port 7 nsew
flabel locali s 29 181 63 215 0 FreeSans 400 0 0 0 C1
port 12 nsew
flabel locali s 585 181 619 215 0 FreeSans 400 0 0 0 A1
port 10 nsew
flabel locali s 401 249 435 283 0 FreeSans 400 0 0 0 A2
port 9 nsew
flabel locali s 305 181 339 215 0 FreeSans 400 0 0 0 B2
port 8 nsew
flabel locali s 305 249 339 283 0 FreeSans 400 0 0 0 B2
port 8 nsew
<< properties >>
string FIXED_BBOX 0 -40 828 504
string path 0.000 -1.000 20.700 -1.000 
<< end >>
