* SPICE3 file created from dac_flat.ext - technology: sky130B

.subckt dac_flat ctl_4_ ctl_3_ ctl_2_ ctl_0_ dum ctl_5_ ctl_7_ ctl_6_ vin vdd sample
+ ctl_1_ out vss
X0 ctl_6_.t3 sky130_fd_sc_hd__inv_2_0.A vss.t48 vss.t47 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 out.t29 sw_top_3.en_buf vin.t24 vdd.t65 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X2 out.t80 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 ctl_2_.t3 sky130_fd_sc_hd__inv_2_6.A vss.t3 vss.t2 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4 out.t81 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 out.t82 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 out.t83 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 vss.t17 sample.t0 sw_top_2.en_buf vss.t16 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 out.t84 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 vss.t111 vdd.t146 vss.t110 vss.t109 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X10 out.t49 sw_top_2.net1 vin.t40 vss.t121 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X11 out.t85 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 out.t86 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 out.t87 carray_0.unitcap_39.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 out.t88 carray_0.unitcap_80.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 vin.t19 sw_top_2.en_buf out.t19 vdd.t45 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X16 out.t89 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 out.t90 sky130_fd_sc_hd__inv_2_7.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 out.t18 sw_top_2.en_buf vin.t12 vdd.t44 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X19 out.t91 carray_0.unitcap_247.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 out.t92 carray_0.unitcap_119.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 sw_top_1.en_buf sample.t1 vss.t19 vss.t18 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 out.t93 carray_0.unitcap_144.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 out.t94 carray_0.unitcap_320.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X24 out.t95 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 vss.t21 sky130_fd_sc_hd__inv_2_9.A.t2 ctl_7_.t3 vss.t20 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 out.t96 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 vss.t7 sky130_fd_sc_hd__inv_2_7.A ctl_3_.t3 vss.t6 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 sw_top_0.net1 sw_top_0.en_buf vdd.t21 vdd.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X29 out.t39 sw_top_1.net1 vin.t39 vss.t108 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X30 out.t97 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 out.t98 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 out.t99 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 out.t100 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 vin.t76 sw_top_1.en_buf out.t79 vdd.t141 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X35 vss.t161 sky130_fd_sc_hd__inv_2_4.A ctl_4_.t3 vss.t160 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 out.t101 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 sw_top_1.net1 sw_top_1.en_buf vss.t157 vss.t156 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X38 sw_top_2.en_buf sample.t2 vdd.t87 vdd.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X39 vss.t85 sample.t3 sw_top_0.en_buf vss.t84 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X40 vss.t149 sky130_fd_sc_hd__inv_2_2.A dum.t3 vss.t148 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X41 out.t102 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 out.t103 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 out.t104 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 out.t105 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 out.t106 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 out.t107 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 out.t108 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 vin.t66 sw_top_3.net1 out.t69 vss.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X49 out.t109 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 vss.t56 sw_top_3.en_buf sw_top_3.net1 vss.t55 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X51 out.t110 carray_0.unitcap_12.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 vin.t53 sw_top_0.net1 out.t59 vss.t131 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X53 ctl_3_.t2 sky130_fd_sc_hd__inv_2_7.A vss.t5 vss.t4 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X54 vss.t15 sw_top_0.en_buf sw_top_0.net1 vss.t14 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X55 ctl_1_.t3 sky130_fd_sc_hd__inv_2_3.A vss.t98 vss.t97 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X56 out.t111 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X57 out.t112 sky130_fd_sc_hd__inv_2_9.A.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 out.t113 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 out.t114 carray_0.unitcap_95.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 out.t115 sky130_fd_sc_hd__inv_2_3.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X61 out.t116 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 out.t117 carray_0.unitcap_183.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X63 sw_top_2.net1 sw_top_2.en_buf vss.t44 vss.t43 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X64 out.t118 carray_0.unitcap_40.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X65 out.t119 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 vss.t24 vdd.t147 vss.t23 vss.t22 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X67 out.t120 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 out.t38 sw_top_1.net1 vin.t38 vss.t107 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X69 out.t121 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 out.t122 carray_0.unitcap_216.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 out.t123 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 out.t124 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 out.t125 carray_0.unitcap_120.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 out.t126 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 vdd.t117 vss.t164 vdd.t116 vdd.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X76 sw_top_1.net1 sw_top_1.en_buf vss.t155 vss.t154 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X77 out.t127 sky130_fd_sc_hd__inv_2_7.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 vin.t65 sw_top_3.net1 out.t68 vss.t140 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X79 out.t128 carray_0.unitcap_322.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X80 out.t129 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 out.t130 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 out.t131 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 out.t132 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 out.t28 sw_top_3.en_buf vin.t23 vdd.t64 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X85 vin.t79 sw_top_1.en_buf out.t78 vdd.t140 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X86 vin.t22 sw_top_3.en_buf out.t27 vdd.t63 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X87 out.t133 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 out.t134 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 vss.t13 sw_top_0.en_buf sw_top_0.net1 vss.t12 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X90 vin.t2 sw_top_0.en_buf out.t9 vdd.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X91 out.t135 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 out.t136 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 vdd.t43 sw_top_2.en_buf sw_top_2.net1 vdd.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X94 out.t137 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 out.t48 sw_top_2.net1 vin.t46 vss.t120 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X96 vin.t52 sw_top_0.net1 out.t58 vss.t130 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X97 out.t8 sw_top_0.en_buf vin.t1 vdd.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X98 vdd.t83 sample.t4 sw_top_1.en_buf vdd.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X99 out.t138 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 vin.t45 sw_top_2.net1 out.t47 vss.t119 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X101 out.t139 carray_0.unitcap_64.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X102 out.t140 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X103 out.t141 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 out.t142 carray_0.unitcap_63.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 out.t143 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 out.t144 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 sw_top_2.net1 sw_top_2.en_buf vss.t42 vss.t41 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X108 out.t17 sw_top_2.en_buf vin.t11 vdd.t41 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X109 out.t145 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 out.t146 carray_0.unitcap_15.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 out.t147 carray_0.unitcap_239.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 out.t148 carray_0.unitcap_143.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 sw_top_0.en_buf sample.t5 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X114 out.t149 carray_0.unitcap_160.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 out.t150 sky130_fd_sc_hd__inv_2_6.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 out.t151 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 out.t37 sw_top_1.net1 vin.t37 vss.t106 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X118 vdd.t114 vss.t165 vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X119 out.t152 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 out.t153 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 out.t154 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 out.t155 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 out.t156 carray_0.unitcap_9.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 vin.t64 sw_top_3.net1 out.t67 vss.t139 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X125 sw_top_0.net1 sw_top_0.en_buf vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X126 vss.t73 sample.t6 sw_top_3.en_buf vss.t72 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X127 out.t157 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 out.t158 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 out.t159 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 out.t160 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 out.t161 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 out.t66 sw_top_3.net1 vin.t62 vss.t138 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X133 out.t162 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 out.t163 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X135 out.t164 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 vdd.t40 sw_top_2.en_buf sw_top_2.net1 vdd.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X137 sw_top_1.en_buf sample.t7 vdd.t80 vdd.t79 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X138 out.t165 sky130_fd_sc_hd__inv_2_7.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 out.t166 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 out.t167 carray_0.unitcap_326.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X141 vss.t27 vdd.t148 vss.t26 vss.t25 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X142 out.t168 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 out.t169 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 out.t170 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 ctl_7_.t1 sky130_fd_sc_hd__inv_2_9.A.t3 vdd.t81 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X146 vdd.t92 sky130_fd_sc_hd__inv_2_5.A.t1 ctl_5_.t1 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X147 out.t171 carray_0.unitcap_32.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 out.t172 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 out.t173 carray_0.unitcap_23.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 out.t174 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X151 out.t175 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 ctl_4_.t1 sky130_fd_sc_hd__inv_2_4.A vdd.t143 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X153 out.t176 carray_0.unitcap_240.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 out.t177 carray_0.unitcap_191.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 dum.t1 sky130_fd_sc_hd__inv_2_2.A vdd.t123 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X156 out.t178 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 out.t179 carray_0.unitcap_112.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 out.t180 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 out.t181 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X160 out.t182 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 out.t36 sw_top_1.net1 vin.t36 vss.t105 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X162 vss.t30 vdd.t149 vss.t29 vss.t28 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X163 vin.t78 sw_top_1.en_buf out.t77 vdd.t139 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X164 vdd.t78 sky130_fd_sc_hd__inv_2_8.A ctl_0_.t1 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X165 vin.t35 sw_top_1.net1 out.t35 vss.t104 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X166 vdd.t111 vss.t166 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X167 vss.t143 sample.t8 sw_top_3.en_buf vss.t142 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X168 out.t183 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 out.t184 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 out.t185 sky130_fd_sc_hd__inv_2_6.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 ctl_5_.t0 sky130_fd_sc_hd__inv_2_5.A.t2 vdd.t93 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X172 out.t186 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 vin.t59 sw_top_0.net1 out.t57 vss.t129 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X174 out.t187 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 out.t188 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 out.t189 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 vss.t145 sample.t9 sw_top_0.en_buf vss.t144 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X178 out.t65 sw_top_3.net1 vin.t61 vss.t137 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X179 out.t190 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 out.t191 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 out.t192 carray_0.unitcap_288.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 vin.t0 sw_top_0.en_buf out.t7 vdd.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X183 out.t193 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X184 out.t194 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 out.t26 sw_top_3.en_buf vin.t21 vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X186 out.t195 carray_0.unitcap_88.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 out.t196 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 out.t197 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X189 out.t198 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 out.t199 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 out.t6 sw_top_0.en_buf vin.t8 vdd.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X192 out.t200 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 vin.t44 sw_top_2.net1 out.t46 vss.t118 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X194 vdd.t74 sample.t10 sw_top_1.en_buf vdd.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X195 out.t201 carray_0.unitcap_255.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 out.t202 carray_0.unitcap_176.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 out.t203 carray_0.unitcap_331.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 out.t45 sw_top_2.net1 vin.t43 vss.t117 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X199 out.t204 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 out.t205 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X201 out.t206 carray_0.unitcap_111.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 vin.t10 sw_top_2.en_buf out.t16 vdd.t38 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X203 sw_top_3.en_buf sample.t11 vdd.t76 vdd.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X204 ctl_7_.t2 sky130_fd_sc_hd__inv_2_9.A.t4 vss.t79 vss.t78 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X205 out.t207 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 out.t208 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 out.t209 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 out.t210 carray_0.unitcap_175.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 vin.t34 sw_top_1.net1 out.t34 vss.t103 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X210 vss.t89 sky130_fd_sc_hd__inv_2_5.A.t3 ctl_5_.t3 vss.t88 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X211 vss.t61 vdd.t150 vss.t60 vss.t59 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X212 out.t211 sky130_fd_sc_hd__inv_2_7.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 vss.t153 sw_top_1.en_buf sw_top_1.net1 vss.t152 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X214 vdd.t145 sample.t12 sw_top_2.en_buf vdd.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X215 out.t212 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 out.t213 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 out.t214 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 out.t215 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 ctl_4_.t2 sky130_fd_sc_hd__inv_2_4.A vss.t159 vss.t158 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X220 out.t216 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X221 out.t217 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 out.t218 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 out.t64 sw_top_3.net1 vin.t60 vss.t136 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X224 dum.t2 sky130_fd_sc_hd__inv_2_2.A vss.t147 vss.t146 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X225 sw_top_3.net1 sw_top_3.en_buf vss.t54 vss.t53 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X226 out.t219 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 out.t220 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 out.t221 sky130_fd_sc_hd__inv_2_6.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X229 out.t222 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 out.t223 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 vss.t64 vdd.t151 vss.t63 vss.t62 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X232 sw_top_2.en_buf sample.t13 vss.t163 vss.t162 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X233 vss.t71 sky130_fd_sc_hd__inv_2_8.A ctl_0_.t3 vss.t70 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X234 ctl_5_.t2 sky130_fd_sc_hd__inv_2_5.A.t4 vss.t91 vss.t90 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X235 out.t224 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X236 out.t225 carray_0.unitcap_56.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 out.t226 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 out.t227 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 out.t228 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 out.t229 carray_0.unitcap_8.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 vdd.t108 vss.t167 vdd.t107 vdd.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X242 sw_top_3.en_buf sample.t14 vdd.t70 vdd.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X243 out.t230 carray_0.unitcap_215.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 out.t231 carray_0.unitcap_136.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 out.t232 carray_0.unitcap_232.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 out.t233 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 out.t234 sky130_fd_sc_hd__inv_2_5.A.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 out.t235 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 out.t236 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 out.t237 carray_0.unitcap_55.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X251 sw_top_0.en_buf sample.t15 vdd.t72 vdd.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X252 vdd.t61 sw_top_3.en_buf sw_top_3.net1 vdd.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X253 out.t238 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 vss.t67 vdd.t152 vss.t66 vss.t65 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X255 out.t239 carray_0.unitcap_337.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 out.t240 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 out.t241 carray_0.unitcap_135.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 vin.t77 sw_top_1.en_buf out.t76 vdd.t138 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X259 vss.t151 sw_top_1.en_buf sw_top_1.net1 vss.t150 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X260 out.t63 sw_top_3.net1 vin.t69 vss.t135 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X261 vin.t32 sw_top_1.net1 out.t33 vss.t102 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X262 vdd.t25 sample.t16 sw_top_2.en_buf vdd.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X263 out.t242 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 out.t243 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 out.t244 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 vdd.t105 vss.t168 vdd.t104 vdd.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X267 sw_top_3.net1 sw_top_3.en_buf vss.t52 vss.t51 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X268 out.t245 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 out.t25 sw_top_3.en_buf vin.t20 vdd.t59 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X270 vin.t58 sw_top_0.net1 out.t56 vss.t128 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X271 out.t246 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X272 out.t5 sw_top_0.en_buf vin.t7 vdd.t13 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X273 out.t55 sw_top_0.net1 vin.t57 vss.t127 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X274 out.t247 sky130_fd_sc_hd__inv_2_7.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X275 out.t248 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X276 out.t249 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 out.t250 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 out.t251 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 out.t252 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 out.t253 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 out.t254 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X282 sw_top_1.en_buf sample.t17 vdd.t27 vdd.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X283 out.t255 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X284 out.t44 sw_top_2.net1 vin.t42 vss.t116 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X285 vin.t18 sw_top_2.en_buf out.t15 vdd.t37 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X286 out.t256 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 out.t257 carray_0.unitcap_16.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 out.t258 sky130_fd_sc_hd__inv_2_6.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 out.t259 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 out.t260 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 sw_top_1.net1 sw_top_1.en_buf vdd.t137 vdd.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X292 vdd.t23 sample.t18 sw_top_0.en_buf vdd.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X293 vin.t31 sw_top_1.net1 out.t32 vss.t101 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X294 out.t261 carray_0.unitcap_184.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 out.t262 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 out.t263 carray_0.unitcap_199.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 out.t264 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 out.t265 carray_0.unitcap_31.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 out.t266 carray_0.unitcap_256.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 vdd.t1 sky130_fd_sc_hd__inv_2_6.A ctl_2_.t1 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X301 vdd.t58 sw_top_3.en_buf sw_top_3.net1 vdd.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X302 out.t267 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 out.t268 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 out.t269 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 out.t270 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 out.t271 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 out.t272 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X308 vdd.t12 sw_top_0.en_buf sw_top_0.net1 vdd.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X309 out.t273 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 out.t274 carray_0.unitcap_334.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X311 out.t275 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X312 sw_top_2.net1 sw_top_2.en_buf vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X313 out.t276 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X314 out.t277 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 vin.t27 sw_top_3.en_buf out.t24 vdd.t56 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X316 vdd.t102 vss.t169 vdd.t101 vdd.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X317 sw_top_0.net1 sw_top_0.en_buf vss.t11 vss.t10 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X318 out.t4 sw_top_0.en_buf vin.t6 vdd.t10 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X319 out.t278 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 vdd.t47 sky130_fd_sc_hd__inv_2_0.A ctl_6_.t1 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X321 out.t43 sw_top_2.net1 vin.t41 vss.t115 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X322 out.t279 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 out.t280 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 sw_top_2.en_buf sample.t19 vss.t32 vss.t31 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X325 out.t281 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 out.t282 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 out.t283 carray_0.unitcap_248.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 sw_top_1.net1 sw_top_1.en_buf vdd.t135 vdd.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X329 vdd.t99 vss.t170 vdd.t98 vdd.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X330 out.t284 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 out.t285 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 out.t286 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 out.t287 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X334 out.t288 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 out.t289 carray_0.unitcap_104.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 out.t290 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 out.t291 carray_0.unitcap_79.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 out.t14 sw_top_2.en_buf vin.t17 vdd.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X339 vin.t30 sw_top_1.net1 out.t31 vss.t100 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X340 out.t292 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 out.t293 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 out.t294 carray_0.unitcap_338.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X343 out.t295 carray_0.unitcap_159.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X344 out.t296 carray_0.unitcap_168.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 vdd.t91 sky130_fd_sc_hd__inv_2_3.A ctl_1_.t1 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X346 vdd.t9 sw_top_0.en_buf sw_top_0.net1 vdd.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X347 ctl_0_.t0 sky130_fd_sc_hd__inv_2_8.A vdd.t77 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X348 out.t297 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 out.t298 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 out.t299 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X351 out.t75 sw_top_1.en_buf vin.t72 vdd.t133 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X352 out.t54 sw_top_0.net1 vin.t56 vss.t126 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X353 out.t300 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 out.t301 carray_0.unitcap_10.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 sw_top_2.net1 sw_top_2.en_buf vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X356 vdd.t96 vss.t171 vdd.t95 vdd.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X357 vin.t55 sw_top_0.net1 out.t53 vss.t125 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X358 out.t302 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 out.t303 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 out.t304 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X361 out.t305 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 out.t306 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 out.t307 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 out.t3 sw_top_0.en_buf vin.t5 vdd.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X365 out.t308 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 out.t309 sky130_fd_sc_hd__inv_2_2.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X367 vss.t1 sky130_fd_sc_hd__inv_2_6.A ctl_2_.t2 vss.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X368 out.t52 sw_top_0.net1 vin.t54 vss.t124 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X369 vin.t26 sw_top_3.en_buf out.t23 vdd.t55 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X370 out.t310 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 out.t311 carray_0.unitcap_330.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 out.t312 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 out.t313 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 out.t314 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 vin.t49 sw_top_2.net1 out.t42 vss.t114 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X376 out.t13 sw_top_2.en_buf vin.t16 vdd.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X377 out.t315 carray_0.unitcap_208.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 vss.t40 sw_top_2.en_buf sw_top_2.net1 vss.t39 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X379 vdd.t89 sample.t20 sw_top_3.en_buf vdd.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X380 out.t316 carray_0.unitcap_207.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 out.t317 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 out.t318 carray_0.unitcap_48.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 out.t319 carray_0.unitcap_7.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 vss.t87 sample.t21 sw_top_1.en_buf vss.t86 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X385 vin.t15 sw_top_2.en_buf out.t12 vdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X386 vss.t46 sky130_fd_sc_hd__inv_2_0.A ctl_6_.t2 vss.t45 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X387 out.t320 sky130_fd_sc_hd__inv_2_7.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 out.t30 sw_top_1.net1 vin.t33 vss.t99 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X389 out.t321 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 out.t322 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 out.t323 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 out.t324 carray_0.unitcap_231.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X393 out.t325 carray_0.unitcap_103.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 out.t326 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 out.t327 carray_0.unitcap_128.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 sw_top_0.en_buf sample.t22 vss.t81 vss.t80 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X397 out.t74 sw_top_1.en_buf vin.t71 vdd.t132 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X398 out.t328 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 out.t329 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 out.t330 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 out.t331 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 out.t332 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 vin.t25 sw_top_3.en_buf out.t22 vdd.t54 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X404 out.t333 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 out.t334 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 vss.t96 sky130_fd_sc_hd__inv_2_3.A ctl_1_.t2 vss.t95 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X407 out.t335 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 out.t336 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 out.t337 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 out.t338 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 sw_top_0.net1 sw_top_0.en_buf vss.t9 vss.t8 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X412 out.t339 carray_0.unitcap_13.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 ctl_0_.t2 sky130_fd_sc_hd__inv_2_8.A vss.t69 vss.t68 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X414 vin.t4 sw_top_0.en_buf out.t2 vdd.t6 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X415 out.t340 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 out.t341 sky130_fd_sc_hd__inv_2_9.A.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 out.t342 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 out.t343 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 vin.t48 sw_top_2.net1 out.t41 vss.t113 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X420 out.t344 sky130_fd_sc_hd__inv_2_3.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 out.t345 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 out.t346 carray_0.unitcap_87.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 out.t347 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 sw_top_1.en_buf sample.t23 vss.t83 vss.t82 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X425 vss.t38 sw_top_2.en_buf sw_top_2.net1 vss.t37 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X426 vdd.t119 sample.t24 sw_top_3.en_buf vdd.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X427 out.t348 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 out.t349 carray_0.unitcap_336.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 out.t350 carray_0.unitcap_192.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 out.t351 carray_0.unitcap_151.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 vdd.t121 sample.t25 sw_top_0.en_buf vdd.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X432 out.t352 carray_0.unitcap_24.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 out.t73 sw_top_1.en_buf vin.t70 vdd.t131 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X434 out.t353 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 out.t354 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 out.t355 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 out.t356 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 out.t62 sw_top_3.net1 vin.t68 vss.t134 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X439 vin.t29 sw_top_3.en_buf out.t21 vdd.t53 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X440 out.t51 sw_top_0.net1 vin.t51 vss.t123 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X441 out.t357 sky130_fd_sc_hd__inv_2_7.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 out.t358 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 out.t359 carray_0.unitcap_324.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 out.t360 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 out.t361 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 out.t362 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 out.t363 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 out.t364 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 vin.t47 sw_top_2.net1 out.t40 vss.t112 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X450 out.t365 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 out.t366 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 out.t367 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 out.t11 sw_top_2.en_buf vin.t14 vdd.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.3
X454 vin.t3 sw_top_0.en_buf out.t1 vdd.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.3
X455 out.t368 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 out.t369 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 vin.t13 sw_top_2.en_buf out.t10 vdd.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X458 out.t370 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 out.t371 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 out.t372 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 out.t373 carray_0.unitcap_47.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 vdd.t130 sw_top_1.en_buf sw_top_1.net1 vdd.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X463 out.t374 carray_0.unitcap_72.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 out.t375 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 out.t376 carray_0.unitcap_14.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 out.t377 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 out.t378 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 out.t379 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 out.t380 carray_0.unitcap_223.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 ctl_6_.t0 sky130_fd_sc_hd__inv_2_0.A vdd.t46 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X471 out.t381 carray_0.unitcap_152.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 out.t382 carray_0.unitcap_321.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X473 out.t383 carray_0.unitcap_127.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 vss.t58 sample.t26 sw_top_1.en_buf vss.t57 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X475 out.t72 sw_top_1.en_buf vin.t75 vdd.t128 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X476 sw_top_3.net1 sw_top_3.en_buf vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X477 ctl_2_.t0 sky130_fd_sc_hd__inv_2_6.A vdd.t0 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X478 sw_top_2.en_buf sample.t27 vdd.t68 vdd.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X479 out.t384 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 out.t385 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X481 sw_top_3.en_buf sample.t28 vss.t75 vss.t74 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X482 out.t386 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 out.t387 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 vin.t67 sw_top_3.net1 out.t61 vss.t133 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X485 out.t388 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 out.t20 sw_top_3.en_buf vin.t28 vdd.t50 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X487 out.t389 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 out.t390 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 out.t391 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 out.t392 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 out.t393 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 vdd.t66 sky130_fd_sc_hd__inv_2_9.A.t5 ctl_7_.t0 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X493 vss.t77 sample.t29 sw_top_2.en_buf vss.t76 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X494 vdd.t3 sky130_fd_sc_hd__inv_2_7.A ctl_3_.t1 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X495 out.t394 sky130_fd_sc_hd__inv_2_7.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X496 out.t395 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 out.t396 carray_0.unitcap_328.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 out.t397 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 out.t398 carray_0.unitcap_71.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X500 out.t399 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 out.t400 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 out.t401 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 vdd.t127 sw_top_1.en_buf sw_top_1.net1 vdd.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X504 vdd.t142 sky130_fd_sc_hd__inv_2_4.A ctl_4_.t0 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X505 out.t402 carray_0.unitcap_167.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 vss.t94 vdd.t153 vss.t93 vss.t92 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X507 out.t403 carray_0.unitcap_200.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 out.t404 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 out.t405 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 vdd.t122 sky130_fd_sc_hd__inv_2_2.A dum.t0 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X511 out.t406 carray_0.unitcap_0.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 sw_top_3.net1 sw_top_3.en_buf vdd.t49 vdd.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X513 out.t407 sky130_fd_sc_hd__inv_2_5.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 ctl_3_.t0 sky130_fd_sc_hd__inv_2_7.A vdd.t2 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X515 out.t408 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 out.t409 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 out.t410 carray_0.unitcap_96.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 out.t411 carray_0.unitcap_224.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 out.t71 sw_top_1.en_buf vin.t74 vdd.t125 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X520 ctl_1_.t0 sky130_fd_sc_hd__inv_2_3.A vdd.t90 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X521 out.t412 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 out.t413 carray_0.unitcap_11.cn sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 sw_top_3.en_buf sample.t30 vss.t34 vss.t33 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X524 vin.t73 sw_top_1.en_buf out.t70 vdd.t124 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X525 out.t414 sky130_fd_sc_hd__inv_2_4.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 out.t415 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 out.t416 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 out.t417 sky130_fd_sc_hd__inv_2_9.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 out.t418 sky130_fd_sc_hd__inv_2_0.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 out.t419 sky130_fd_sc_hd__inv_2_8.A sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 out.t50 sw_top_0.net1 vin.t50 vss.t122 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X532 sw_top_0.en_buf sample.t31 vss.t36 vss.t35 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X533 vss.t50 sw_top_3.en_buf sw_top_3.net1 vss.t49 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X534 vin.t9 sw_top_0.en_buf out.t0 vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
X535 vin.t63 sw_top_3.net1 out.t60 vss.t132 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.3
R0 vss.n166 vss.n165 137683
R1 vss.n165 vss.n164 19857.7
R2 vss.n165 vss.n42 11545.9
R3 vss.n169 vss.n40 10267.2
R4 vss.n143 vss.n140 10267.2
R5 vss.n151 vss.n130 10267.2
R6 vss.n159 vss.n121 10267.2
R7 vss.n167 vss.n41 7329.75
R8 vss.n149 vss.n131 6110.51
R9 vss.n157 vss.n42 6110.51
R10 vss.n141 vss.n41 6110.51
R11 vss.n170 vss.n169 5290.03
R12 vss.n144 vss.n143 5290.03
R13 vss.n152 vss.n151 5290.03
R14 vss.n160 vss.n159 5290.03
R15 vss.n170 vss.n38 4820.71
R16 vss.n144 vss.n137 4820.71
R17 vss.n152 vss.n127 4820.71
R18 vss.n160 vss.n118 4820.71
R19 vss.n131 vss.n42 3902.77
R20 vss.n131 vss.n41 3902.77
R21 vss.n167 vss 3595.41
R22 vss.n158 vss.n157 2015.03
R23 vss.n150 vss.n149 2015.03
R24 vss.n142 vss.n141 2015.03
R25 vss.n157 vss.n156 1920.57
R26 vss.n149 vss.n148 1920.57
R27 vss.n141 vss.n35 1920.57
R28 vss.n158 vss.t123 1361.72
R29 vss.n150 vss.t107 1361.72
R30 vss.n142 vss.t120 1361.72
R31 vss.n168 vss.t135 1361.72
R32 vss.n162 vss.t130 1345.97
R33 vss.n154 vss.t102 1345.97
R34 vss.n146 vss.t113 1345.97
R35 vss.n172 vss.t141 1345.97
R36 vss.t130 vss.t127 928.802
R37 vss.t127 vss.t131 928.802
R38 vss.t131 vss.t124 928.802
R39 vss.t124 vss.t125 928.802
R40 vss.t129 vss.t122 928.802
R41 vss.t126 vss.t129 928.802
R42 vss.t128 vss.t126 928.802
R43 vss.t123 vss.t128 928.802
R44 vss.t102 vss.t108 928.802
R45 vss.t108 vss.t103 928.802
R46 vss.t103 vss.t99 928.802
R47 vss.t99 vss.t104 928.802
R48 vss.t100 vss.t105 928.802
R49 vss.t106 vss.t100 928.802
R50 vss.t101 vss.t106 928.802
R51 vss.t107 vss.t101 928.802
R52 vss.t113 vss.t117 928.802
R53 vss.t117 vss.t114 928.802
R54 vss.t114 vss.t121 928.802
R55 vss.t121 vss.t118 928.802
R56 vss.t119 vss.t115 928.802
R57 vss.t116 vss.t119 928.802
R58 vss.t112 vss.t116 928.802
R59 vss.t120 vss.t112 928.802
R60 vss.t141 vss.t136 928.802
R61 vss.t136 vss.t132 928.802
R62 vss.t132 vss.t137 928.802
R63 vss.t137 vss.t133 928.802
R64 vss.t139 vss.t138 928.802
R65 vss.t134 vss.t139 928.802
R66 vss.t140 vss.t134 928.802
R67 vss.t135 vss.t140 928.802
R68 vss.t59 vss 777.63
R69 vss.t92 vss 777.63
R70 vss.t25 vss 777.63
R71 vss.t28 vss 777.63
R72 vss vss.t59 667.384
R73 vss vss.t92 667.384
R74 vss vss.t25 667.384
R75 vss vss.t28 667.384
R76 vss.n156 vss.n155 585
R77 vss.n148 vss.n147 585
R78 vss.n173 vss.n35 585
R79 vss.n164 vss.n163 585
R80 vss.t125 vss.n161 464.401
R81 vss.n161 vss.t122 464.401
R82 vss.t104 vss.n153 464.401
R83 vss.n153 vss.t105 464.401
R84 vss.t118 vss.n145 464.401
R85 vss.n145 vss.t115 464.401
R86 vss.t133 vss.n171 464.401
R87 vss.n171 vss.t138 464.401
R88 vss.n168 vss.n167 401.432
R89 vss.t22 vss.n166 348.457
R90 vss.t62 vss 328.771
R91 vss.t65 vss 328.771
R92 vss.t109 vss 328.771
R93 vss.t14 vss 261.834
R94 vss.t152 vss 261.834
R95 vss.t39 vss 261.834
R96 vss.t49 vss 261.834
R97 vss.t144 vss 248.054
R98 vss.t57 vss 248.054
R99 vss.t76 vss 248.054
R100 vss.t72 vss 248.054
R101 vss vss.t22 214.587
R102 vss vss.t62 214.587
R103 vss vss.t65 214.587
R104 vss vss.t109 214.587
R105 vss.n173 vss.n36 201.282
R106 vss.n147 vss.n134 201.282
R107 vss.n155 vss.n124 201.282
R108 vss.n163 vss.n45 201.282
R109 vss.n182 vss.t34 193.933
R110 vss.n180 vss.t52 193.933
R111 vss.n1 vss.t11 193.933
R112 vss.n3 vss.t81 193.933
R113 vss.n13 vss.t155 193.933
R114 vss.n15 vss.t83 193.933
R115 vss.n25 vss.t42 193.933
R116 vss.n27 vss.t163 193.933
R117 vss.n181 vss.t73 192.982
R118 vss.n223 vss.t50 192.982
R119 vss.n0 vss.t15 192.982
R120 vss.n2 vss.t145 192.982
R121 vss.n323 vss.t153 192.982
R122 vss.n14 vss.t58 192.982
R123 vss.n273 vss.t40 192.982
R124 vss.n26 vss.t77 192.982
R125 vss.n166 vss 187.642
R126 vss.n51 vss.t166 183.082
R127 vss.n11 vss.t170 183.082
R128 vss.n23 vss.t171 183.082
R129 vss.n178 vss.t165 183.082
R130 vss.t8 vss.t14 165.369
R131 vss.t12 vss.t8 165.369
R132 vss.t10 vss.t12 165.369
R133 vss.t35 vss.t144 165.369
R134 vss.t84 vss.t35 165.369
R135 vss.t80 vss.t84 165.369
R136 vss.t156 vss.t152 165.369
R137 vss.t150 vss.t156 165.369
R138 vss.t154 vss.t150 165.369
R139 vss.t18 vss.t57 165.369
R140 vss.t86 vss.t18 165.369
R141 vss.t82 vss.t86 165.369
R142 vss.t43 vss.t39 165.369
R143 vss.t37 vss.t43 165.369
R144 vss.t41 vss.t37 165.369
R145 vss.t31 vss.t76 165.369
R146 vss.t16 vss.t31 165.369
R147 vss.t162 vss.t16 165.369
R148 vss.t53 vss.t49 165.369
R149 vss.t55 vss.t53 165.369
R150 vss.t51 vss.t55 165.369
R151 vss.t74 vss.t72 165.369
R152 vss.t142 vss.t74 165.369
R153 vss.t33 vss.t142 165.369
R154 vss.n173 vss.n34 156.441
R155 vss.n147 vss.n133 156.441
R156 vss.n155 vss.n123 156.441
R157 vss.n163 vss.n44 156.441
R158 vss vss.t10 147.651
R159 vss vss.t80 147.651
R160 vss vss.t154 147.651
R161 vss vss.t82 147.651
R162 vss vss.t41 147.651
R163 vss vss.t162 147.651
R164 vss vss.t51 147.651
R165 vss vss.t33 147.651
R166 vss.n179 vss.t111 121.956
R167 vss.n32 vss.t110 121.956
R168 vss.n202 vss.t29 121.956
R169 vss.n183 vss.t30 121.956
R170 vss.n28 vss.t27 121.956
R171 vss.n252 vss.t26 121.956
R172 vss.n24 vss.t67 121.956
R173 vss.n20 vss.t66 121.956
R174 vss.n16 vss.t94 121.956
R175 vss.n302 vss.t93 121.956
R176 vss.n12 vss.t64 121.956
R177 vss.n8 vss.t63 121.956
R178 vss.n4 vss.t61 121.956
R179 vss.n352 vss.t60 121.956
R180 vss.n52 vss.t24 121.956
R181 vss.n46 vss.t23 121.956
R182 vss.n164 vss.n43 118.069
R183 vss.n156 vss.n122 118.069
R184 vss.n148 vss.n132 118.069
R185 vss.n37 vss.n35 118.069
R186 vss.n104 vss.t149 116.115
R187 vss.n58 vss.t71 116.115
R188 vss.n96 vss.t96 116.115
R189 vss.n62 vss.t1 116.115
R190 vss.n90 vss.t5 116.115
R191 vss.n87 vss.t159 116.115
R192 vss.n82 vss.t91 116.115
R193 vss.n79 vss.t48 116.115
R194 vss.n74 vss.t79 116.115
R195 vss.n368 vss.n367 114.713
R196 vss.n359 vss.n358 114.713
R197 vss.n318 vss.n317 114.713
R198 vss.n309 vss.n308 114.713
R199 vss.n268 vss.n267 114.713
R200 vss.n259 vss.n258 114.713
R201 vss.n218 vss.n217 114.713
R202 vss.n209 vss.n208 114.713
R203 vss.n72 vss.t21 113.677
R204 vss.n106 vss.t147 113.677
R205 vss.n103 vss.t69 113.677
R206 vss.n98 vss.t98 113.677
R207 vss.n95 vss.t3 113.677
R208 vss.n88 vss.t7 113.677
R209 vss.n66 vss.t161 113.677
R210 vss.n80 vss.t89 113.677
R211 vss.n70 vss.t46 113.677
R212 vss.n190 vss.n189 76.0005
R213 vss.n340 vss.n339 76.0005
R214 vss.n290 vss.n289 76.0005
R215 vss.n240 vss.n239 76.0005
R216 vss.n109 vss.n108 48.3595
R217 vss.t4 vss.t0 47.0331
R218 vss.t78 vss 38.9494
R219 vss.t47 vss 38.9494
R220 vss.t90 vss 38.9494
R221 vss.t158 vss 38.2145
R222 vss.n188 vss.t168 34.2973
R223 vss.n238 vss.t167 34.2973
R224 vss.n288 vss.t164 34.2973
R225 vss.n338 vss.t169 34.2973
R226 vss vss.t70 30.6207
R227 vss vss.t148 30.1308
R228 vss vss.t95 29.6409
R229 vss.n105 vss.n104 25.224
R230 vss.n106 vss.n105 25.224
R231 vss.n102 vss.n58 25.224
R232 vss.n103 vss.n102 25.224
R233 vss.n97 vss.n96 25.224
R234 vss.n98 vss.n97 25.224
R235 vss.n94 vss.n62 25.224
R236 vss.n95 vss.n94 25.224
R237 vss.n89 vss.n88 25.224
R238 vss.n90 vss.n89 25.224
R239 vss.n86 vss.n66 25.224
R240 vss.n87 vss.n86 25.224
R241 vss.n81 vss.n80 25.224
R242 vss.n82 vss.n81 25.224
R243 vss.n78 vss.n70 25.224
R244 vss.n79 vss.n78 25.224
R245 vss.n73 vss.n72 25.224
R246 vss.n74 vss.n73 25.224
R247 vss.n367 vss.t9 24.9236
R248 vss.n367 vss.t13 24.9236
R249 vss.n358 vss.t36 24.9236
R250 vss.n358 vss.t85 24.9236
R251 vss.n317 vss.t157 24.9236
R252 vss.n317 vss.t151 24.9236
R253 vss.n308 vss.t19 24.9236
R254 vss.n308 vss.t87 24.9236
R255 vss.n267 vss.t44 24.9236
R256 vss.n267 vss.t38 24.9236
R257 vss.n258 vss.t32 24.9236
R258 vss.n258 vss.t17 24.9236
R259 vss.n217 vss.t54 24.9236
R260 vss.n217 vss.t56 24.9236
R261 vss.n208 vss.t75 24.9236
R262 vss.n208 vss.t143 24.9236
R263 vss.n90 vss.n62 21.8358
R264 vss.t20 vss.t78 20.5773
R265 vss.t45 vss.t47 20.5773
R266 vss.t88 vss.t90 20.5773
R267 vss.t160 vss.t158 20.5773
R268 vss.t6 vss.t4 20.5773
R269 vss.t0 vss.t2 20.5773
R270 vss.t95 vss.t97 20.5773
R271 vss.t70 vss.t68 20.5773
R272 vss.t148 vss.t146 20.5773
R273 vss.n98 vss.n58 20.3299
R274 vss.n82 vss.n66 20.3299
R275 vss.n80 vss.n79 20.3299
R276 vss.n74 vss.n70 20.3299
R277 vss.n104 vss.n103 19.577
R278 vss.n40 vss.n39 19.3358
R279 vss.n140 vss.n139 19.3358
R280 vss.n130 vss.n129 19.3358
R281 vss.n121 vss.n120 19.3358
R282 vss.n224 vss.n223 19.3355
R283 vss.n53 vss.n0 19.3355
R284 vss.n324 vss.n323 19.3355
R285 vss.n274 vss.n273 19.3355
R286 vss.n88 vss.n87 19.2005
R287 vss.n96 vss.n95 18.824
R288 vss.n181 vss.n180 18.0711
R289 vss.n2 vss.n1 18.0711
R290 vss.n14 vss.n13 18.0711
R291 vss.n26 vss.n25 18.0711
R292 vss.n203 vss.n182 17.4103
R293 vss.n353 vss.n3 17.4103
R294 vss.n303 vss.n15 17.4103
R295 vss.n253 vss.n27 17.4103
R296 vss.t2 vss 16.4129
R297 vss.t97 vss 16.4129
R298 vss.t68 vss 16.4129
R299 vss.t146 vss 16.4129
R300 vss.n333 vss.n332 16.0891
R301 vss.n283 vss.n282 16.0891
R302 vss.n233 vss.n232 16.0891
R303 vss.n162 vss.n43 15.7429
R304 vss.n154 vss.n122 15.7429
R305 vss.n146 vss.n132 15.7429
R306 vss.n172 vss.n37 15.7429
R307 vss.n117 vss.n116 12.2372
R308 vss.n175 vss.n174 12.2362
R309 vss.n136 vss.n135 12.2362
R310 vss.n126 vss.n125 12.2362
R311 vss.n36 vss.n33 9.39653
R312 vss.n138 vss.n134 9.39653
R313 vss.n128 vss.n124 9.39653
R314 vss.n119 vss.n45 9.39653
R315 vss.n155 vss.n126 9.3005
R316 vss.n155 vss.n154 9.3005
R317 vss.n147 vss.n136 9.3005
R318 vss.n147 vss.n146 9.3005
R319 vss.n174 vss.n173 9.3005
R320 vss.n173 vss.n172 9.3005
R321 vss.n163 vss.n117 9.3005
R322 vss.n163 vss.n162 9.3005
R323 vss.n165 vss 8.57416
R324 vss vss.t20 8.08423
R325 vss vss.t45 8.08423
R326 vss vss.t88 8.08423
R327 vss vss.t160 8.08423
R328 vss vss.t6 8.08423
R329 vss.n202 vss.n201 5.85582
R330 vss.n352 vss.n351 5.85582
R331 vss.n302 vss.n301 5.85582
R332 vss.n252 vss.n251 5.85582
R333 vss.n47 vss.n46 5.1356
R334 vss.n8 vss.n7 5.0092
R335 vss.n20 vss.n19 5.0092
R336 vss.n32 vss.n31 5.0092
R337 vss.n38 vss.n36 4.97808
R338 vss.n137 vss.n134 4.97808
R339 vss.n127 vss.n124 4.97808
R340 vss.n118 vss.n45 4.97808
R341 vss.n184 vss.n183 4.91351
R342 vss.n189 vss.n188 4.85762
R343 vss.n239 vss.n238 4.85762
R344 vss.n289 vss.n288 4.85762
R345 vss.n339 vss.n338 4.85762
R346 vss.n72 vss 4.67264
R347 vss.n73 vss.n71 4.6505
R348 vss.n75 vss.n74 4.6505
R349 vss.n76 vss.n70 4.6505
R350 vss.n79 vss.n69 4.6505
R351 vss.n80 vss.n68 4.6505
R352 vss.n83 vss.n82 4.6505
R353 vss.n84 vss.n66 4.6505
R354 vss.n87 vss.n65 4.6505
R355 vss.n88 vss.n64 4.6505
R356 vss.n91 vss.n90 4.6505
R357 vss.n92 vss.n62 4.6505
R358 vss.n95 vss.n61 4.6505
R359 vss.n96 vss.n60 4.6505
R360 vss.n99 vss.n98 4.6505
R361 vss.n100 vss.n58 4.6505
R362 vss.n103 vss.n57 4.6505
R363 vss.n104 vss.n56 4.6505
R364 vss.n78 vss.n77 4.6505
R365 vss.n81 vss.n67 4.6505
R366 vss.n86 vss.n85 4.6505
R367 vss.n89 vss.n63 4.6505
R368 vss.n94 vss.n93 4.6505
R369 vss.n97 vss.n59 4.6505
R370 vss.n102 vss.n101 4.6505
R371 vss.n105 vss.n55 4.6505
R372 vss.n107 vss.n106 4.6505
R373 vss.n223 vss.n222 4.6505
R374 vss.n214 vss.n180 4.6505
R375 vss.n213 vss.n181 4.6505
R376 vss.n205 vss.n182 4.6505
R377 vss.n255 vss.n27 4.6505
R378 vss.n263 vss.n26 4.6505
R379 vss.n264 vss.n25 4.6505
R380 vss.n273 vss.n272 4.6505
R381 vss.n305 vss.n15 4.6505
R382 vss.n313 vss.n14 4.6505
R383 vss.n314 vss.n13 4.6505
R384 vss.n323 vss.n322 4.6505
R385 vss.n355 vss.n3 4.6505
R386 vss.n363 vss.n2 4.6505
R387 vss.n364 vss.n1 4.6505
R388 vss.n372 vss.n0 4.6505
R389 vss.n187 vss.n186 4.6505
R390 vss.n192 vss.n191 4.6505
R391 vss.n195 vss.n194 4.6505
R392 vss.n197 vss.n196 4.6505
R393 vss.n199 vss.n198 4.6505
R394 vss.n204 vss.n203 4.6505
R395 vss.n207 vss.n206 4.6505
R396 vss.n210 vss.n209 4.6505
R397 vss.n212 vss.n211 4.6505
R398 vss.n216 vss.n215 4.6505
R399 vss.n219 vss.n218 4.6505
R400 vss.n221 vss.n220 4.6505
R401 vss.n225 vss.n224 4.6505
R402 vss.n232 vss.n231 4.6505
R403 vss.n234 vss.n233 4.6505
R404 vss.n237 vss.n236 4.6505
R405 vss.n242 vss.n241 4.6505
R406 vss.n245 vss.n244 4.6505
R407 vss.n247 vss.n246 4.6505
R408 vss.n249 vss.n248 4.6505
R409 vss.n254 vss.n253 4.6505
R410 vss.n257 vss.n256 4.6505
R411 vss.n260 vss.n259 4.6505
R412 vss.n262 vss.n261 4.6505
R413 vss.n266 vss.n265 4.6505
R414 vss.n269 vss.n268 4.6505
R415 vss.n271 vss.n270 4.6505
R416 vss.n275 vss.n274 4.6505
R417 vss.n282 vss.n281 4.6505
R418 vss.n284 vss.n283 4.6505
R419 vss.n287 vss.n286 4.6505
R420 vss.n292 vss.n291 4.6505
R421 vss.n295 vss.n294 4.6505
R422 vss.n297 vss.n296 4.6505
R423 vss.n299 vss.n298 4.6505
R424 vss.n304 vss.n303 4.6505
R425 vss.n307 vss.n306 4.6505
R426 vss.n310 vss.n309 4.6505
R427 vss.n312 vss.n311 4.6505
R428 vss.n316 vss.n315 4.6505
R429 vss.n319 vss.n318 4.6505
R430 vss.n321 vss.n320 4.6505
R431 vss.n325 vss.n324 4.6505
R432 vss.n332 vss.n331 4.6505
R433 vss.n334 vss.n333 4.6505
R434 vss.n337 vss.n336 4.6505
R435 vss.n342 vss.n341 4.6505
R436 vss.n345 vss.n344 4.6505
R437 vss.n347 vss.n346 4.6505
R438 vss.n349 vss.n348 4.6505
R439 vss.n354 vss.n353 4.6505
R440 vss.n357 vss.n356 4.6505
R441 vss.n360 vss.n359 4.6505
R442 vss.n362 vss.n361 4.6505
R443 vss.n366 vss.n365 4.6505
R444 vss.n369 vss.n368 4.6505
R445 vss.n371 vss.n370 4.6505
R446 vss.n54 vss.n53 4.6505
R447 vss.n51 vss.n50 4.5918
R448 vss.n108 vss 4.19097
R449 vss.n39 vss.n33 3.77398
R450 vss.n139 vss.n138 3.77398
R451 vss.n129 vss.n128 3.77398
R452 vss.n120 vss.n119 3.77398
R453 vss.n229 vss.n177 2.99647
R454 vss.n279 vss.n22 2.99647
R455 vss.n329 vss.n10 2.99647
R456 vss.n115 vss.n113 2.99647
R457 vss.n52 vss.n51 1.18311
R458 vss.n12 vss.n11 1.18311
R459 vss.n24 vss.n23 1.18311
R460 vss.n179 vss.n178 1.18311
R461 vss.n186 vss.n185 1.14023
R462 vss.n336 vss.n335 1.14023
R463 vss.n286 vss.n285 1.14023
R464 vss.n236 vss.n235 1.14023
R465 vss.n49 vss.n48 0.974413
R466 vss.n7 vss.n6 0.974413
R467 vss.n19 vss.n18 0.974413
R468 vss.n31 vss.n30 0.974413
R469 vss.n191 vss.n190 0.833377
R470 vss.n341 vss.n340 0.833377
R471 vss.n291 vss.n290 0.833377
R472 vss.n241 vss.n240 0.833377
R473 vss.n174 vss.n33 0.753441
R474 vss.n138 vss.n136 0.753441
R475 vss.n128 vss.n126 0.753441
R476 vss.n119 vss.n117 0.753441
R477 vss.n127 vss.n122 0.67602
R478 vss.n137 vss.n132 0.67602
R479 vss.n38 vss.n37 0.67602
R480 vss.n118 vss.n43 0.67602
R481 vss.n194 vss.n193 0.526527
R482 vss.n344 vss.n343 0.526527
R483 vss.n294 vss.n293 0.526527
R484 vss.n244 vss.n243 0.526527
R485 vss.n108 vss 0.495181
R486 vss.n53 vss.n52 0.417891
R487 vss.n332 vss.n8 0.417891
R488 vss.n324 vss.n12 0.417891
R489 vss.n282 vss.n20 0.417891
R490 vss.n274 vss.n24 0.417891
R491 vss.n232 vss.n32 0.417891
R492 vss.n224 vss.n179 0.417891
R493 vss.n203 vss.n202 0.409011
R494 vss.n353 vss.n352 0.409011
R495 vss.n303 vss.n302 0.409011
R496 vss.n253 vss.n252 0.409011
R497 vss.n130 vss.n122 0.288252
R498 vss.n140 vss.n132 0.288252
R499 vss.n40 vss.n37 0.288252
R500 vss.n121 vss.n43 0.288252
R501 vss.n333 vss.n4 0.263514
R502 vss.n283 vss.n16 0.263514
R503 vss.n233 vss.n28 0.263514
R504 vss.n50 vss.n49 0.209196
R505 vss.n6 vss.n5 0.209196
R506 vss.n18 vss.n17 0.209196
R507 vss.n30 vss.n29 0.209196
R508 vss.n123 vss.n122 0.134398
R509 vss.n133 vss.n132 0.134398
R510 vss.n37 vss.n34 0.134398
R511 vss.n44 vss.n43 0.134398
R512 vss.n129 vss.n123 0.12657
R513 vss.n139 vss.n133 0.12657
R514 vss.n39 vss.n34 0.12657
R515 vss.n120 vss.n44 0.12657
R516 vss.n75 vss.n71 0.120292
R517 vss.n77 vss.n69 0.120292
R518 vss.n83 vss.n67 0.120292
R519 vss.n85 vss.n65 0.120292
R520 vss.n91 vss.n63 0.120292
R521 vss.n93 vss.n92 0.120292
R522 vss.n93 vss.n61 0.120292
R523 vss.n60 vss.n59 0.120292
R524 vss.n99 vss.n59 0.120292
R525 vss.n101 vss.n100 0.120292
R526 vss.n101 vss.n57 0.120292
R527 vss.n56 vss.n55 0.120292
R528 vss.n107 vss.n55 0.120292
R529 vss.n372 vss.n371 0.120292
R530 vss.n371 vss.n369 0.120292
R531 vss.n369 vss.n366 0.120292
R532 vss.n366 vss.n364 0.120292
R533 vss.n363 vss.n362 0.120292
R534 vss.n362 vss.n360 0.120292
R535 vss.n360 vss.n357 0.120292
R536 vss.n357 vss.n355 0.120292
R537 vss.n354 vss.n350 0.120292
R538 vss.n350 vss.n349 0.120292
R539 vss.n349 vss.n347 0.120292
R540 vss.n347 vss.n345 0.120292
R541 vss.n345 vss.n342 0.120292
R542 vss.n342 vss.n337 0.120292
R543 vss.n337 vss.n334 0.120292
R544 vss.n322 vss.n321 0.120292
R545 vss.n321 vss.n319 0.120292
R546 vss.n319 vss.n316 0.120292
R547 vss.n316 vss.n314 0.120292
R548 vss.n313 vss.n312 0.120292
R549 vss.n312 vss.n310 0.120292
R550 vss.n310 vss.n307 0.120292
R551 vss.n307 vss.n305 0.120292
R552 vss.n304 vss.n300 0.120292
R553 vss.n300 vss.n299 0.120292
R554 vss.n299 vss.n297 0.120292
R555 vss.n297 vss.n295 0.120292
R556 vss.n295 vss.n292 0.120292
R557 vss.n292 vss.n287 0.120292
R558 vss.n287 vss.n284 0.120292
R559 vss.n272 vss.n271 0.120292
R560 vss.n271 vss.n269 0.120292
R561 vss.n269 vss.n266 0.120292
R562 vss.n266 vss.n264 0.120292
R563 vss.n263 vss.n262 0.120292
R564 vss.n262 vss.n260 0.120292
R565 vss.n260 vss.n257 0.120292
R566 vss.n257 vss.n255 0.120292
R567 vss.n254 vss.n250 0.120292
R568 vss.n250 vss.n249 0.120292
R569 vss.n249 vss.n247 0.120292
R570 vss.n247 vss.n245 0.120292
R571 vss.n245 vss.n242 0.120292
R572 vss.n242 vss.n237 0.120292
R573 vss.n237 vss.n234 0.120292
R574 vss.n222 vss.n221 0.120292
R575 vss.n221 vss.n219 0.120292
R576 vss.n219 vss.n216 0.120292
R577 vss.n216 vss.n214 0.120292
R578 vss.n213 vss.n212 0.120292
R579 vss.n212 vss.n210 0.120292
R580 vss.n210 vss.n207 0.120292
R581 vss.n207 vss.n205 0.120292
R582 vss.n204 vss.n200 0.120292
R583 vss.n200 vss.n199 0.120292
R584 vss.n199 vss.n197 0.120292
R585 vss.n197 vss.n195 0.120292
R586 vss.n195 vss.n192 0.120292
R587 vss.n192 vss.n187 0.120292
R588 vss.n187 vss.n184 0.120292
R589 vss.n326 vss.n325 0.116385
R590 vss.n276 vss.n275 0.116385
R591 vss.n226 vss.n225 0.116385
R592 vss vss.n71 0.0981562
R593 vss.n77 vss 0.0981562
R594 vss vss.n67 0.0981562
R595 vss.n85 vss 0.0981562
R596 vss vss.n63 0.0981562
R597 vss.n331 vss.n330 0.0682083
R598 vss.n281 vss.n280 0.0682083
R599 vss.n231 vss.n230 0.0682083
R600 vss.n151 vss.n150 0.067449
R601 vss.n143 vss.n142 0.067449
R602 vss.n169 vss.n168 0.067449
R603 vss.n159 vss.n158 0.067449
R604 vss.n110 vss.n109 0.0643021
R605 vss vss.n75 0.0603958
R606 vss.n76 vss 0.0603958
R607 vss.n69 vss 0.0603958
R608 vss vss.n68 0.0603958
R609 vss vss.n83 0.0603958
R610 vss.n84 vss 0.0603958
R611 vss.n65 vss 0.0603958
R612 vss vss.n91 0.0603958
R613 vss.n92 vss 0.0603958
R614 vss.n100 vss 0.0603958
R615 vss vss.n372 0.0603958
R616 vss.n331 vss 0.0603958
R617 vss.n322 vss 0.0603958
R618 vss.n281 vss 0.0603958
R619 vss.n272 vss 0.0603958
R620 vss.n231 vss 0.0603958
R621 vss.n222 vss 0.0603958
R622 vss vss.n56 0.0577917
R623 vss vss.n354 0.0577917
R624 vss vss.n304 0.0577917
R625 vss vss.n254 0.0577917
R626 vss vss.n204 0.0577917
R627 vss vss.n64 0.0564896
R628 vss vss.n60 0.0551875
R629 vss.n109 vss.n54 0.0525833
R630 vss vss.n363 0.0512812
R631 vss vss.n313 0.0512812
R632 vss vss.n263 0.0512812
R633 vss vss.n213 0.0512812
R634 vss.n177 vss 0.0441068
R635 vss vss.n22 0.0441068
R636 vss vss.n10 0.0441068
R637 vss vss.n115 0.0441068
R638 vss.n113 vss.n112 0.0304479
R639 vss.n329 vss.n328 0.0304479
R640 vss.n279 vss.n278 0.0304479
R641 vss.n229 vss.n228 0.0304479
R642 vss vss.n76 0.0226354
R643 vss.n68 vss 0.0226354
R644 vss vss.n84 0.0226354
R645 vss.n64 vss 0.0226354
R646 vss.n61 vss 0.0226354
R647 vss vss.n99 0.0226354
R648 vss.n57 vss 0.0226354
R649 vss vss.n107 0.0226354
R650 vss.n54 vss 0.0226354
R651 vss.n364 vss 0.0226354
R652 vss.n355 vss 0.0226354
R653 vss.n334 vss 0.0226354
R654 vss.n325 vss 0.0226354
R655 vss.n314 vss 0.0226354
R656 vss.n305 vss 0.0226354
R657 vss.n284 vss 0.0226354
R658 vss.n275 vss 0.0226354
R659 vss.n264 vss 0.0226354
R660 vss.n255 vss 0.0226354
R661 vss.n234 vss 0.0226354
R662 vss.n225 vss 0.0226354
R663 vss.n214 vss 0.0226354
R664 vss.n205 vss 0.0226354
R665 vss.n184 vss 0.0226354
R666 vss.n175 vss 0.0219286
R667 vss.n135 vss 0.0219286
R668 vss.n125 vss 0.0219286
R669 vss.n116 vss 0.0219286
R670 vss.n112 vss.n111 0.0187292
R671 vss.n328 vss.n327 0.0187292
R672 vss.n278 vss.n277 0.0187292
R673 vss.n228 vss.n227 0.0187292
R674 vss.n177 vss.n176 0.0178015
R675 vss.n22 vss.n21 0.0178015
R676 vss.n10 vss.n9 0.0178015
R677 vss.n115 vss.n114 0.0178015
R678 vss vss.n175 0.0149231
R679 vss.n135 vss 0.0149231
R680 vss.n125 vss 0.0149231
R681 vss.n116 vss 0.0149231
R682 vss.n153 vss.n152 0.0145006
R683 vss.n145 vss.n144 0.0145006
R684 vss.n171 vss.n170 0.0145006
R685 vss.n161 vss.n160 0.0145006
R686 vss.n113 vss.n47 0.00440625
R687 vss.n111 vss.n110 0.00440625
R688 vss.n330 vss.n329 0.00440625
R689 vss.n327 vss.n326 0.00440625
R690 vss.n280 vss.n279 0.00440625
R691 vss.n277 vss.n276 0.00440625
R692 vss.n230 vss.n229 0.00440625
R693 vss.n227 vss.n226 0.00440625
R694 ctl_6_ ctl_6_.n0 50.4671
R695 ctl_6_.n2 ctl_6_.t1 26.5955
R696 ctl_6_.n2 ctl_6_.t0 26.5955
R697 ctl_6_.n0 ctl_6_.t2 24.9236
R698 ctl_6_.n0 ctl_6_.t3 24.9236
R699 ctl_6_ ctl_6_.n1 11.2645
R700 ctl_6_.n10 ctl_6_.n9 9.30959
R701 ctl_6_.n3 ctl_6_.n2 8.88979
R702 ctl_6_.n11 ctl_6_.n10 6.78838
R703 ctl_6_.n1 ctl_6_ 6.1445
R704 ctl_6_.n1 ctl_6_ 4.65505
R705 ctl_6_.n9 ctl_6_.n8 3.29747
R706 ctl_6_.n11 ctl_6_ 2.0485
R707 ctl_6_ ctl_6_.n11 1.55202
R708 ctl_6_.n5 ctl_6_ 0.66901
R709 ctl_6_.n8 ctl_6_.n3 0.582318
R710 ctl_6_.n6 ctl_6_.n5 0.0569547
R711 ctl_6_.n7 ctl_6_.n4 0.00635938
R712 ctl_6_.n8 ctl_6_.n7 0.00116875
R713 ctl_6_.n7 ctl_6_.n6 0.00100244
R714 vin.n52 vin.t25 29.3118
R715 vin.n37 vin.t15 29.3118
R716 vin.n22 vin.t79 29.3118
R717 vin.n8 vin.t3 29.3118
R718 vin.n57 vin.t23 29.3084
R719 vin.n42 vin.t14 29.3084
R720 vin.n27 vin.t70 29.3084
R721 vin.n13 vin.t7 29.3084
R722 vin.n50 vin.t21 28.5655
R723 vin.n50 vin.t26 28.5655
R724 vin.n48 vin.t24 28.5655
R725 vin.n48 vin.t27 28.5655
R726 vin.n46 vin.t28 28.5655
R727 vin.n46 vin.t22 28.5655
R728 vin.n44 vin.t20 28.5655
R729 vin.n44 vin.t29 28.5655
R730 vin.n35 vin.t12 28.5655
R731 vin.n35 vin.t10 28.5655
R732 vin.n33 vin.t16 28.5655
R733 vin.n33 vin.t19 28.5655
R734 vin.n31 vin.t17 28.5655
R735 vin.n31 vin.t13 28.5655
R736 vin.n29 vin.t11 28.5655
R737 vin.n29 vin.t18 28.5655
R738 vin.n20 vin.t71 28.5655
R739 vin.n20 vin.t76 28.5655
R740 vin.n18 vin.t72 28.5655
R741 vin.n18 vin.t73 28.5655
R742 vin.n16 vin.t74 28.5655
R743 vin.n16 vin.t78 28.5655
R744 vin.n14 vin.t75 28.5655
R745 vin.n14 vin.t77 28.5655
R746 vin.n6 vin.t1 28.5655
R747 vin.n6 vin.t4 28.5655
R748 vin.n4 vin.t8 28.5655
R749 vin.n4 vin.t0 28.5655
R750 vin.n2 vin.t5 28.5655
R751 vin.n2 vin.t9 28.5655
R752 vin.n0 vin.t6 28.5655
R753 vin.n0 vin.t2 28.5655
R754 vin.n52 vin.t66 18.1397
R755 vin.n57 vin.t69 18.1397
R756 vin.n37 vin.t48 18.1397
R757 vin.n42 vin.t46 18.1397
R758 vin.n22 vin.t32 18.1397
R759 vin.n27 vin.t38 18.1397
R760 vin.n8 vin.t52 18.1397
R761 vin.n13 vin.t51 18.1397
R762 vin.n51 vin.t60 17.4005
R763 vin.n51 vin.t63 17.4005
R764 vin.n49 vin.t61 17.4005
R765 vin.n49 vin.t67 17.4005
R766 vin.n47 vin.t62 17.4005
R767 vin.n47 vin.t64 17.4005
R768 vin.n45 vin.t68 17.4005
R769 vin.n45 vin.t65 17.4005
R770 vin.n36 vin.t43 17.4005
R771 vin.n36 vin.t49 17.4005
R772 vin.n34 vin.t40 17.4005
R773 vin.n34 vin.t44 17.4005
R774 vin.n32 vin.t41 17.4005
R775 vin.n32 vin.t45 17.4005
R776 vin.n30 vin.t42 17.4005
R777 vin.n30 vin.t47 17.4005
R778 vin.n21 vin.t39 17.4005
R779 vin.n21 vin.t34 17.4005
R780 vin.n19 vin.t33 17.4005
R781 vin.n19 vin.t35 17.4005
R782 vin.n17 vin.t36 17.4005
R783 vin.n17 vin.t30 17.4005
R784 vin.n15 vin.t37 17.4005
R785 vin.n15 vin.t31 17.4005
R786 vin.n7 vin.t57 17.4005
R787 vin.n7 vin.t53 17.4005
R788 vin.n5 vin.t54 17.4005
R789 vin.n5 vin.t55 17.4005
R790 vin.n3 vin.t50 17.4005
R791 vin.n3 vin.t59 17.4005
R792 vin.n1 vin.t56 17.4005
R793 vin.n1 vin.t58 17.4005
R794 vin.n62 vin.n61 13.5897
R795 vin.n59 vin 7.61508
R796 vin.n60 vin.n43 6.84826
R797 vin.n61 vin.n28 6.84826
R798 vin.n59 vin.n58 6.83948
R799 vin.n60 vin.n59 6.68453
R800 vin.n61 vin.n60 6.66717
R801 vin.n54 vin.n53 0.811311
R802 vin.n39 vin.n38 0.811311
R803 vin.n24 vin.n23 0.811311
R804 vin.n10 vin.n9 0.811311
R805 vin.n56 vin.n55 0.799575
R806 vin.n41 vin.n40 0.799575
R807 vin.n26 vin.n25 0.799575
R808 vin.n12 vin.n11 0.799575
R809 vin.n55 vin.n54 0.794419
R810 vin.n40 vin.n39 0.794419
R811 vin.n25 vin.n24 0.794419
R812 vin.n11 vin.n10 0.794419
R813 vin.n53 vin.n52 0.787662
R814 vin.n38 vin.n37 0.787662
R815 vin.n23 vin.n22 0.787662
R816 vin.n9 vin.n8 0.787662
R817 vin.n57 vin.n56 0.773526
R818 vin.n42 vin.n41 0.773526
R819 vin.n27 vin.n26 0.773526
R820 vin.n13 vin.n12 0.773526
R821 vin.n53 vin.n50 0.746823
R822 vin.n54 vin.n48 0.746823
R823 vin.n55 vin.n46 0.746823
R824 vin.n38 vin.n35 0.746823
R825 vin.n39 vin.n33 0.746823
R826 vin.n40 vin.n31 0.746823
R827 vin.n23 vin.n20 0.746823
R828 vin.n24 vin.n18 0.746823
R829 vin.n25 vin.n16 0.746823
R830 vin.n9 vin.n6 0.746823
R831 vin.n10 vin.n4 0.746823
R832 vin.n11 vin.n2 0.746823
R833 vin.n56 vin.n44 0.743351
R834 vin.n41 vin.n29 0.743351
R835 vin.n26 vin.n14 0.743351
R836 vin.n12 vin.n0 0.743351
R837 vin.n53 vin.n51 0.739748
R838 vin.n54 vin.n49 0.739748
R839 vin.n55 vin.n47 0.739748
R840 vin.n56 vin.n45 0.739748
R841 vin.n38 vin.n36 0.739748
R842 vin.n39 vin.n34 0.739748
R843 vin.n40 vin.n32 0.739748
R844 vin.n41 vin.n30 0.739748
R845 vin.n23 vin.n21 0.739748
R846 vin.n24 vin.n19 0.739748
R847 vin.n25 vin.n17 0.739748
R848 vin.n26 vin.n15 0.739748
R849 vin.n9 vin.n7 0.739748
R850 vin.n10 vin.n5 0.739748
R851 vin.n11 vin.n3 0.739748
R852 vin.n12 vin.n1 0.739748
R853 vin.n28 vin.n27 0.542884
R854 vin.n58 vin.n57 0.534103
R855 vin.n43 vin.n42 0.532467
R856 vin.n62 vin.n13 0.52205
R857 vin vin.n62 0.0557885
R858 vin.n43 vin 0.0485769
R859 vin.n28 vin 0.0413654
R860 vin.n58 vin 0.0356562
R861 out out.n59 105.326
R862 out out.n14 105.326
R863 out out.n44 105.031
R864 out out.n29 104.98
R865 out.n56 out.n55 86.3387
R866 out.n41 out.n40 86.3387
R867 out.n26 out.n25 86.3387
R868 out.n11 out.n10 86.3387
R869 out.n59 out.n58 85.9532
R870 out.n44 out.n43 85.9532
R871 out.n29 out.n28 85.9532
R872 out.n14 out.n13 85.9532
R873 out.n55 out.n53 84.93
R874 out.n40 out.n38 84.93
R875 out.n25 out.n23 84.93
R876 out.n10 out.n8 84.93
R877 out.n57 out.n49 83.8601
R878 out.n42 out.n34 83.8601
R879 out.n27 out.n19 83.8601
R880 out.n12 out.n4 83.8601
R881 out.n59 out.n45 83.6607
R882 out.n44 out.n30 83.6607
R883 out.n29 out.n15 83.6607
R884 out.n14 out.n0 83.6607
R885 out.n58 out.n47 83.2397
R886 out.n43 out.n32 83.2397
R887 out.n28 out.n17 83.2397
R888 out.n13 out.n2 83.2397
R889 out.n56 out.n51 83.0069
R890 out.n41 out.n36 83.0069
R891 out.n26 out.n21 83.0069
R892 out.n11 out.n6 83.0069
R893 out.n59 out.n46 81.7128
R894 out.n44 out.n31 81.7128
R895 out.n29 out.n16 81.7128
R896 out.n14 out.n1 81.7128
R897 out.n58 out.n48 81.5763
R898 out.n43 out.n33 81.5763
R899 out.n28 out.n18 81.5763
R900 out.n13 out.n3 81.5763
R901 out.n57 out.n50 81.3057
R902 out.n42 out.n35 81.3057
R903 out.n27 out.n20 81.3057
R904 out.n12 out.n5 81.3057
R905 out.n58 out.n57 81.2978
R906 out.n43 out.n42 81.2978
R907 out.n28 out.n27 81.2978
R908 out.n13 out.n12 81.2978
R909 out.n408 out.n407 81.0971
R910 out.n57 out.n56 80.9519
R911 out.n42 out.n41 80.9519
R912 out.n27 out.n26 80.9519
R913 out.n12 out.n11 80.9519
R914 out.n56 out.n52 80.2068
R915 out.n41 out.n37 80.2068
R916 out.n26 out.n22 80.2068
R917 out.n11 out.n7 80.2068
R918 out.n55 out.n54 80.0412
R919 out.n40 out.n39 80.0412
R920 out.n25 out.n24 80.0412
R921 out.n10 out.n9 80.0412
R922 out.n406 out 62.2988
R923 out.n407 out 54.3231
R924 out.n405 out 41.2855
R925 out.n53 out.t21 28.5655
R926 out.n53 out.t28 28.5655
R927 out.n47 out.t23 28.5655
R928 out.n47 out.t29 28.5655
R929 out.n49 out.t24 28.5655
R930 out.n49 out.t20 28.5655
R931 out.n51 out.t27 28.5655
R932 out.n51 out.t25 28.5655
R933 out.n45 out.t22 28.5655
R934 out.n45 out.t26 28.5655
R935 out.n38 out.t15 28.5655
R936 out.n38 out.t11 28.5655
R937 out.n32 out.t16 28.5655
R938 out.n32 out.t13 28.5655
R939 out.n34 out.t19 28.5655
R940 out.n34 out.t14 28.5655
R941 out.n36 out.t10 28.5655
R942 out.n36 out.t17 28.5655
R943 out.n30 out.t12 28.5655
R944 out.n30 out.t18 28.5655
R945 out.n23 out.t76 28.5655
R946 out.n23 out.t73 28.5655
R947 out.n17 out.t79 28.5655
R948 out.n17 out.t75 28.5655
R949 out.n19 out.t70 28.5655
R950 out.n19 out.t71 28.5655
R951 out.n21 out.t77 28.5655
R952 out.n21 out.t72 28.5655
R953 out.n15 out.t78 28.5655
R954 out.n15 out.t74 28.5655
R955 out.n8 out.t9 28.5655
R956 out.n8 out.t5 28.5655
R957 out.n2 out.t2 28.5655
R958 out.n2 out.t6 28.5655
R959 out.n4 out.t7 28.5655
R960 out.n4 out.t3 28.5655
R961 out.n6 out.t0 28.5655
R962 out.n6 out.t4 28.5655
R963 out.n0 out.t1 28.5655
R964 out.n0 out.t8 28.5655
R965 out.n54 out.t68 17.4005
R966 out.n54 out.t63 17.4005
R967 out.n48 out.t60 17.4005
R968 out.n48 out.t65 17.4005
R969 out.n50 out.t61 17.4005
R970 out.n50 out.t66 17.4005
R971 out.n52 out.t67 17.4005
R972 out.n52 out.t62 17.4005
R973 out.n46 out.t69 17.4005
R974 out.n46 out.t64 17.4005
R975 out.n39 out.t40 17.4005
R976 out.n39 out.t48 17.4005
R977 out.n33 out.t42 17.4005
R978 out.n33 out.t49 17.4005
R979 out.n35 out.t46 17.4005
R980 out.n35 out.t43 17.4005
R981 out.n37 out.t47 17.4005
R982 out.n37 out.t44 17.4005
R983 out.n31 out.t41 17.4005
R984 out.n31 out.t45 17.4005
R985 out.n24 out.t32 17.4005
R986 out.n24 out.t38 17.4005
R987 out.n18 out.t34 17.4005
R988 out.n18 out.t30 17.4005
R989 out.n20 out.t35 17.4005
R990 out.n20 out.t36 17.4005
R991 out.n22 out.t31 17.4005
R992 out.n22 out.t37 17.4005
R993 out.n16 out.t33 17.4005
R994 out.n16 out.t39 17.4005
R995 out.n9 out.t56 17.4005
R996 out.n9 out.t51 17.4005
R997 out.n3 out.t59 17.4005
R998 out.n3 out.t52 17.4005
R999 out.n5 out.t53 17.4005
R1000 out.n5 out.t50 17.4005
R1001 out.n7 out.t57 17.4005
R1002 out.n7 out.t54 17.4005
R1003 out.n1 out.t58 17.4005
R1004 out.n1 out.t55 17.4005
R1005 out.n407 out.n406 6.79693
R1006 out.n404 out 6.29528
R1007 out.n406 out.n405 3.67907
R1008 out.n404 out.n403 2.59022
R1009 out.n408 out 1.09764
R1010 out.n405 out.n404 1.08457
R1011 out out.n408 1.06717
R1012 out.n87 out 0.400915
R1013 out.n88 out 0.400915
R1014 out.n89 out 0.400915
R1015 out.n90 out 0.400915
R1016 out.n91 out 0.400915
R1017 out.n92 out 0.400915
R1018 out.n93 out 0.400915
R1019 out.n94 out 0.400915
R1020 out.n95 out 0.400915
R1021 out.n96 out 0.400915
R1022 out.n97 out 0.400915
R1023 out.n98 out 0.400915
R1024 out.n99 out 0.400915
R1025 out.n100 out 0.400915
R1026 out.n101 out 0.400915
R1027 out.n102 out 0.400915
R1028 out.n103 out 0.400915
R1029 out.n104 out 0.400915
R1030 out.n105 out 0.400915
R1031 out.n106 out 0.400915
R1032 out.n107 out 0.400915
R1033 out.n108 out 0.400915
R1034 out.n109 out 0.400915
R1035 out.n110 out 0.400915
R1036 out.n111 out 0.400915
R1037 out.n112 out 0.400915
R1038 out.n113 out 0.400915
R1039 out.n114 out 0.400915
R1040 out.n115 out 0.400915
R1041 out.n116 out 0.400915
R1042 out.n117 out 0.400915
R1043 out.n118 out 0.400915
R1044 out.n119 out 0.400915
R1045 out.n120 out 0.400915
R1046 out.n121 out 0.400915
R1047 out.n122 out 0.400915
R1048 out.n123 out 0.400915
R1049 out.n124 out 0.400915
R1050 out.n125 out 0.400915
R1051 out.n126 out 0.400915
R1052 out.n127 out 0.400915
R1053 out.n128 out 0.400915
R1054 out.n129 out 0.400915
R1055 out.n130 out 0.400915
R1056 out.n131 out 0.400915
R1057 out.n132 out 0.400915
R1058 out.n133 out 0.400915
R1059 out.n134 out 0.400915
R1060 out.n135 out 0.400915
R1061 out.n136 out 0.400915
R1062 out.n137 out 0.400915
R1063 out.n138 out 0.400915
R1064 out.n139 out 0.400915
R1065 out.n140 out 0.400915
R1066 out.n141 out 0.400915
R1067 out.n142 out 0.400915
R1068 out.n143 out 0.400915
R1069 out.n144 out 0.400915
R1070 out.n145 out 0.400915
R1071 out.n146 out 0.400915
R1072 out.n147 out 0.400915
R1073 out.n148 out 0.400915
R1074 out.n149 out 0.400915
R1075 out.n150 out 0.400915
R1076 out.n151 out 0.400915
R1077 out.n152 out 0.400915
R1078 out.n153 out 0.400915
R1079 out.n154 out 0.400915
R1080 out.n155 out 0.400915
R1081 out.n156 out 0.400915
R1082 out.n157 out 0.400915
R1083 out.n158 out 0.400915
R1084 out.n159 out 0.400915
R1085 out.n160 out 0.400915
R1086 out.n161 out 0.400915
R1087 out.n162 out 0.400915
R1088 out.n163 out 0.400915
R1089 out.n164 out 0.400915
R1090 out.n165 out 0.400915
R1091 out.n166 out 0.400915
R1092 out.n167 out 0.400915
R1093 out.n168 out 0.400915
R1094 out.n169 out 0.400915
R1095 out.n170 out 0.400915
R1096 out.n171 out 0.400915
R1097 out.n172 out 0.400915
R1098 out.n173 out 0.400915
R1099 out.n174 out 0.400915
R1100 out.n175 out 0.400915
R1101 out.n176 out 0.400915
R1102 out.n177 out 0.400915
R1103 out.n178 out 0.400915
R1104 out.n179 out 0.400915
R1105 out.n180 out 0.400915
R1106 out.n181 out 0.400915
R1107 out.n182 out 0.400915
R1108 out.n183 out 0.400915
R1109 out.n184 out 0.400915
R1110 out.n185 out 0.400915
R1111 out.n186 out 0.400915
R1112 out.n187 out 0.400915
R1113 out.n188 out 0.400915
R1114 out.n189 out 0.400915
R1115 out.n190 out 0.400915
R1116 out.n191 out 0.400915
R1117 out.n192 out 0.400915
R1118 out.n193 out 0.400915
R1119 out.n194 out 0.400915
R1120 out.n195 out 0.400915
R1121 out.n196 out 0.400915
R1122 out.n197 out 0.400915
R1123 out.n198 out 0.400915
R1124 out.n199 out 0.400915
R1125 out.n200 out 0.400915
R1126 out.n201 out 0.400915
R1127 out.n202 out 0.400915
R1128 out.n203 out 0.400915
R1129 out.n204 out 0.400915
R1130 out.n205 out 0.400915
R1131 out.n206 out 0.400915
R1132 out.n207 out 0.400915
R1133 out.n208 out 0.400915
R1134 out.n209 out 0.400915
R1135 out.n210 out 0.400915
R1136 out.n211 out 0.400915
R1137 out.n212 out 0.400915
R1138 out.n213 out 0.400915
R1139 out.n214 out 0.400915
R1140 out.n215 out 0.400915
R1141 out.n216 out 0.400915
R1142 out.n217 out 0.400915
R1143 out.n218 out 0.400915
R1144 out.n219 out 0.400915
R1145 out.n220 out 0.400915
R1146 out.n221 out 0.400915
R1147 out.n222 out 0.400915
R1148 out.n223 out 0.400915
R1149 out.n224 out 0.400915
R1150 out.n225 out 0.400915
R1151 out.n226 out 0.400915
R1152 out.n227 out 0.400915
R1153 out.n228 out 0.400915
R1154 out.n229 out 0.400915
R1155 out.n230 out 0.400915
R1156 out.n231 out 0.400915
R1157 out.n232 out 0.400915
R1158 out.n233 out 0.400915
R1159 out.n234 out 0.400915
R1160 out.n235 out 0.400915
R1161 out.n236 out 0.400915
R1162 out.n237 out 0.400915
R1163 out.n238 out 0.400915
R1164 out.n239 out 0.400915
R1165 out.n240 out 0.400915
R1166 out.n241 out 0.400915
R1167 out.n242 out 0.400915
R1168 out.n243 out 0.400915
R1169 out.n244 out 0.400915
R1170 out.n245 out 0.400915
R1171 out.n246 out 0.400915
R1172 out.n247 out 0.400915
R1173 out.n248 out 0.400915
R1174 out.n249 out 0.400915
R1175 out.n250 out 0.400915
R1176 out.n251 out 0.400915
R1177 out.n252 out 0.400915
R1178 out.n253 out 0.400915
R1179 out.n254 out 0.400915
R1180 out.n255 out 0.400915
R1181 out.n256 out 0.400915
R1182 out.n257 out 0.400915
R1183 out.n258 out 0.400915
R1184 out.n259 out 0.400915
R1185 out.n260 out 0.400915
R1186 out.n261 out 0.400915
R1187 out.n262 out 0.400915
R1188 out.n263 out 0.400915
R1189 out.n264 out 0.400915
R1190 out.n265 out 0.400915
R1191 out.n266 out 0.400915
R1192 out.n267 out 0.400915
R1193 out.n268 out 0.400915
R1194 out.n269 out 0.400915
R1195 out.n270 out 0.400915
R1196 out.n271 out 0.400915
R1197 out.n272 out 0.400915
R1198 out.n273 out 0.400915
R1199 out.n274 out 0.400915
R1200 out.n275 out 0.400915
R1201 out.n276 out 0.400915
R1202 out.n277 out 0.400915
R1203 out.n278 out 0.400915
R1204 out.n279 out 0.400915
R1205 out.n280 out 0.400915
R1206 out.n281 out 0.400915
R1207 out.n282 out 0.400915
R1208 out.n283 out 0.400915
R1209 out.n284 out 0.400915
R1210 out.n285 out 0.400915
R1211 out.n286 out 0.400915
R1212 out.n287 out 0.400915
R1213 out.n288 out 0.400915
R1214 out.n289 out 0.400915
R1215 out.n290 out 0.400915
R1216 out.n291 out 0.400915
R1217 out.n292 out 0.400915
R1218 out.n293 out 0.400915
R1219 out.n294 out 0.400915
R1220 out.n295 out 0.400915
R1221 out.n296 out 0.400915
R1222 out.n297 out 0.400915
R1223 out.n298 out 0.400915
R1224 out.n299 out 0.400915
R1225 out.n300 out 0.400915
R1226 out.n301 out 0.400915
R1227 out.n302 out 0.400915
R1228 out.n303 out 0.400915
R1229 out out.n307 0.400915
R1230 out out.n308 0.400915
R1231 out out.n309 0.400915
R1232 out out.n310 0.400915
R1233 out out.n311 0.400915
R1234 out out.n312 0.400915
R1235 out out.n313 0.400915
R1236 out out.n314 0.400915
R1237 out out.n315 0.400915
R1238 out out.n316 0.400915
R1239 out out.n317 0.400915
R1240 out out.n318 0.400915
R1241 out out.n319 0.400915
R1242 out out.n320 0.400915
R1243 out out.n321 0.400915
R1244 out out.n322 0.400915
R1245 out out.n323 0.400915
R1246 out out.n324 0.400915
R1247 out out.n325 0.400915
R1248 out out.n326 0.400915
R1249 out out.n327 0.400915
R1250 out out.n328 0.400915
R1251 out out.n329 0.400915
R1252 out out.n330 0.400915
R1253 out out.n331 0.400915
R1254 out out.n332 0.400915
R1255 out out.n333 0.400915
R1256 out out.n334 0.400915
R1257 out out.n335 0.400915
R1258 out out.n336 0.400915
R1259 out out.n337 0.400915
R1260 out out.n338 0.400915
R1261 out out.n339 0.400915
R1262 out.n352 out 0.400915
R1263 out.n353 out 0.400915
R1264 out.n354 out 0.400915
R1265 out.n355 out 0.400915
R1266 out.n356 out 0.400915
R1267 out.n357 out 0.400915
R1268 out.n358 out 0.400915
R1269 out.n359 out 0.400915
R1270 out.n360 out 0.400915
R1271 out.n361 out 0.400915
R1272 out.n362 out 0.400915
R1273 out.n363 out 0.400915
R1274 out.n364 out 0.400915
R1275 out.n365 out 0.400915
R1276 out.n366 out 0.400915
R1277 out.n367 out 0.400915
R1278 out.n368 out 0.400915
R1279 out.n369 out 0.400915
R1280 out.n370 out 0.400915
R1281 out.n371 out 0.400915
R1282 out.n372 out 0.400915
R1283 out.n373 out 0.400915
R1284 out.n374 out 0.400915
R1285 out.n375 out 0.400915
R1286 out.n376 out 0.400915
R1287 out.n377 out 0.400915
R1288 out.n378 out 0.400915
R1289 out.n379 out 0.400915
R1290 out.n380 out 0.400915
R1291 out.n381 out 0.400915
R1292 out.n382 out 0.400915
R1293 out.n383 out 0.400915
R1294 out out.n398 0.400915
R1295 out out.n399 0.400915
R1296 out out.n400 0.400915
R1297 out out.n401 0.400915
R1298 out.n60 out 0.400915
R1299 out.n61 out 0.400915
R1300 out.n62 out 0.400915
R1301 out.n63 out 0.400915
R1302 out.n64 out 0.400915
R1303 out.n65 out 0.400915
R1304 out.n66 out 0.400915
R1305 out.n67 out 0.400915
R1306 out.n68 out 0.400915
R1307 out.n69 out 0.400915
R1308 out.n70 out 0.400915
R1309 out.n71 out 0.400915
R1310 out.n72 out 0.400915
R1311 out.n73 out 0.400915
R1312 out.n74 out 0.400915
R1313 out.n75 out 0.400915
R1314 out.n76 out 0.400915
R1315 out.n77 out 0.400915
R1316 out.n78 out 0.400915
R1317 out.n79 out 0.400915
R1318 out.n80 out 0.400915
R1319 out.n81 out 0.400915
R1320 out.n82 out 0.400915
R1321 out.n83 out 0.400915
R1322 out.n84 out 0.400915
R1323 out.n85 out 0.400915
R1324 out.n351 out.n350 0.398433
R1325 out.n395 out 0.377415
R1326 out.n393 out 0.377415
R1327 out.n391 out 0.377415
R1328 out.n389 out 0.377415
R1329 out.n387 out 0.377415
R1330 out.n385 out 0.377415
R1331 out.n304 out 0.377415
R1332 out out.n397 0.377415
R1333 out out.n86 0.250087
R1334 out.n342 out 0.250087
R1335 out.n343 out 0.250087
R1336 out.n344 out 0.250087
R1337 out.n345 out 0.250087
R1338 out.n346 out 0.250087
R1339 out.n347 out 0.250087
R1340 out.n348 out 0.250087
R1341 out.n349 out 0.250087
R1342 out out.n386 0.250087
R1343 out out.n388 0.250087
R1344 out out.n390 0.250087
R1345 out out.n392 0.250087
R1346 out out.n394 0.250087
R1347 out out.n396 0.250087
R1348 out.n341 out.n340 0.243372
R1349 out.n306 out.n305 0.241767
R1350 out out.n384 0.226587
R1351 out.n403 out.n402 0.210433
R1352 out.n403 out 0.190981
R1353 out out.t150 0.0215188
R1354 out out.t221 0.0215188
R1355 out out.t115 0.0215188
R1356 out out.t344 0.0215188
R1357 out out.t419 0.0215188
R1358 out out.t309 0.0215188
R1359 out out.t185 0.0215188
R1360 out out.t258 0.0215188
R1361 out out.n87 0.0215186
R1362 out out.n88 0.0215186
R1363 out out.n89 0.0215186
R1364 out out.n90 0.0215186
R1365 out out.n91 0.0215186
R1366 out out.n92 0.0215186
R1367 out out.n93 0.0215186
R1368 out out.n94 0.0215186
R1369 out out.n95 0.0215186
R1370 out out.n96 0.0215186
R1371 out out.n97 0.0215186
R1372 out out.n98 0.0215186
R1373 out out.n99 0.0215186
R1374 out out.n100 0.0215186
R1375 out out.n101 0.0215186
R1376 out out.n102 0.0215186
R1377 out out.n103 0.0215186
R1378 out out.n104 0.0215186
R1379 out out.n105 0.0215186
R1380 out out.n106 0.0215186
R1381 out out.n107 0.0215186
R1382 out out.n108 0.0215186
R1383 out out.n109 0.0215186
R1384 out out.n110 0.0215186
R1385 out out.n111 0.0215186
R1386 out out.n112 0.0215186
R1387 out out.n113 0.0215186
R1388 out out.n114 0.0215186
R1389 out out.n115 0.0215186
R1390 out out.n116 0.0215186
R1391 out out.n117 0.0215186
R1392 out out.n118 0.0215186
R1393 out out.n119 0.0215186
R1394 out out.n120 0.0215186
R1395 out out.n121 0.0215186
R1396 out out.n122 0.0215186
R1397 out out.n123 0.0215186
R1398 out out.n124 0.0215186
R1399 out out.n125 0.0215186
R1400 out out.n126 0.0215186
R1401 out out.n127 0.0215186
R1402 out out.n128 0.0215186
R1403 out out.n129 0.0215186
R1404 out out.n130 0.0215186
R1405 out out.n131 0.0215186
R1406 out out.n132 0.0215186
R1407 out out.n133 0.0215186
R1408 out out.n134 0.0215186
R1409 out out.n135 0.0215186
R1410 out out.n136 0.0215186
R1411 out out.n137 0.0215186
R1412 out out.n138 0.0215186
R1413 out out.n139 0.0215186
R1414 out out.n140 0.0215186
R1415 out out.n141 0.0215186
R1416 out out.n142 0.0215186
R1417 out out.n143 0.0215186
R1418 out out.n144 0.0215186
R1419 out out.n145 0.0215186
R1420 out out.n146 0.0215186
R1421 out out.n147 0.0215186
R1422 out out.n148 0.0215186
R1423 out out.n149 0.0215186
R1424 out out.n150 0.0215186
R1425 out out.n151 0.0215186
R1426 out out.n152 0.0215186
R1427 out out.n153 0.0215186
R1428 out out.n154 0.0215186
R1429 out out.n155 0.0215186
R1430 out out.n156 0.0215186
R1431 out out.n157 0.0215186
R1432 out out.n158 0.0215186
R1433 out out.n159 0.0215186
R1434 out out.n160 0.0215186
R1435 out out.n161 0.0215186
R1436 out out.n162 0.0215186
R1437 out out.n163 0.0215186
R1438 out out.n164 0.0215186
R1439 out out.n165 0.0215186
R1440 out out.n166 0.0215186
R1441 out out.n167 0.0215186
R1442 out out.n168 0.0215186
R1443 out out.n169 0.0215186
R1444 out out.n170 0.0215186
R1445 out out.n171 0.0215186
R1446 out out.n172 0.0215186
R1447 out out.n173 0.0215186
R1448 out out.n174 0.0215186
R1449 out out.n175 0.0215186
R1450 out out.n176 0.0215186
R1451 out out.n177 0.0215186
R1452 out out.n178 0.0215186
R1453 out out.n179 0.0215186
R1454 out out.n180 0.0215186
R1455 out out.n181 0.0215186
R1456 out out.n182 0.0215186
R1457 out out.n183 0.0215186
R1458 out out.n184 0.0215186
R1459 out out.n185 0.0215186
R1460 out out.n186 0.0215186
R1461 out out.n187 0.0215186
R1462 out out.n188 0.0215186
R1463 out out.n189 0.0215186
R1464 out out.n190 0.0215186
R1465 out out.n191 0.0215186
R1466 out out.n192 0.0215186
R1467 out out.n193 0.0215186
R1468 out out.n194 0.0215186
R1469 out out.n195 0.0215186
R1470 out out.n196 0.0215186
R1471 out out.n197 0.0215186
R1472 out out.n198 0.0215186
R1473 out out.n199 0.0215186
R1474 out out.n200 0.0215186
R1475 out out.n201 0.0215186
R1476 out out.n202 0.0215186
R1477 out out.n203 0.0215186
R1478 out out.n204 0.0215186
R1479 out out.n205 0.0215186
R1480 out out.n206 0.0215186
R1481 out out.n207 0.0215186
R1482 out out.n208 0.0215186
R1483 out out.n209 0.0215186
R1484 out out.n210 0.0215186
R1485 out out.n211 0.0215186
R1486 out out.n212 0.0215186
R1487 out out.n213 0.0215186
R1488 out out.n214 0.0215186
R1489 out out.n215 0.0215186
R1490 out out.n216 0.0215186
R1491 out out.n217 0.0215186
R1492 out out.n218 0.0215186
R1493 out out.n219 0.0215186
R1494 out out.n220 0.0215186
R1495 out out.n221 0.0215186
R1496 out out.n222 0.0215186
R1497 out out.n223 0.0215186
R1498 out out.n224 0.0215186
R1499 out out.n225 0.0215186
R1500 out out.n226 0.0215186
R1501 out out.n227 0.0215186
R1502 out out.n228 0.0215186
R1503 out out.n229 0.0215186
R1504 out out.n230 0.0215186
R1505 out out.n231 0.0215186
R1506 out out.n232 0.0215186
R1507 out out.n233 0.0215186
R1508 out out.n234 0.0215186
R1509 out out.n235 0.0215186
R1510 out out.n236 0.0215186
R1511 out out.n237 0.0215186
R1512 out out.n238 0.0215186
R1513 out out.n239 0.0215186
R1514 out out.n240 0.0215186
R1515 out out.n241 0.0215186
R1516 out out.n242 0.0215186
R1517 out out.n243 0.0215186
R1518 out out.n244 0.0215186
R1519 out out.n245 0.0215186
R1520 out out.n246 0.0215186
R1521 out out.n247 0.0215186
R1522 out out.n248 0.0215186
R1523 out out.n249 0.0215186
R1524 out out.n250 0.0215186
R1525 out out.n251 0.0215186
R1526 out out.n252 0.0215186
R1527 out out.n253 0.0215186
R1528 out out.n254 0.0215186
R1529 out out.n255 0.0215186
R1530 out out.n256 0.0215186
R1531 out out.n257 0.0215186
R1532 out out.n258 0.0215186
R1533 out out.n259 0.0215186
R1534 out out.n260 0.0215186
R1535 out out.n261 0.0215186
R1536 out out.n262 0.0215186
R1537 out out.n263 0.0215186
R1538 out out.n264 0.0215186
R1539 out out.n265 0.0215186
R1540 out out.n266 0.0215186
R1541 out out.n267 0.0215186
R1542 out out.n268 0.0215186
R1543 out out.n269 0.0215186
R1544 out out.n270 0.0215186
R1545 out out.n271 0.0215186
R1546 out out.n272 0.0215186
R1547 out out.n273 0.0215186
R1548 out out.n274 0.0215186
R1549 out out.n275 0.0215186
R1550 out out.n276 0.0215186
R1551 out out.n277 0.0215186
R1552 out out.n278 0.0215186
R1553 out out.n279 0.0215186
R1554 out out.n280 0.0215186
R1555 out out.n281 0.0215186
R1556 out out.n282 0.0215186
R1557 out out.n283 0.0215186
R1558 out out.n284 0.0215186
R1559 out out.n285 0.0215186
R1560 out out.n286 0.0215186
R1561 out out.n287 0.0215186
R1562 out out.n288 0.0215186
R1563 out out.n289 0.0215186
R1564 out out.n290 0.0215186
R1565 out out.n291 0.0215186
R1566 out out.n292 0.0215186
R1567 out out.n293 0.0215186
R1568 out out.n294 0.0215186
R1569 out out.n295 0.0215186
R1570 out out.n296 0.0215186
R1571 out out.n297 0.0215186
R1572 out out.n298 0.0215186
R1573 out out.n299 0.0215186
R1574 out out.n300 0.0215186
R1575 out out.n301 0.0215186
R1576 out out.n302 0.0215186
R1577 out out.n303 0.0215186
R1578 out.n308 out 0.0215186
R1579 out.n309 out 0.0215186
R1580 out.n310 out 0.0215186
R1581 out.n311 out 0.0215186
R1582 out.n312 out 0.0215186
R1583 out.n313 out 0.0215186
R1584 out.n314 out 0.0215186
R1585 out.n315 out 0.0215186
R1586 out.n316 out 0.0215186
R1587 out.n317 out 0.0215186
R1588 out.n318 out 0.0215186
R1589 out.n319 out 0.0215186
R1590 out.n320 out 0.0215186
R1591 out.n321 out 0.0215186
R1592 out.n322 out 0.0215186
R1593 out.n323 out 0.0215186
R1594 out.n324 out 0.0215186
R1595 out.n325 out 0.0215186
R1596 out.n326 out 0.0215186
R1597 out.n327 out 0.0215186
R1598 out.n328 out 0.0215186
R1599 out.n329 out 0.0215186
R1600 out.n330 out 0.0215186
R1601 out.n331 out 0.0215186
R1602 out.n332 out 0.0215186
R1603 out.n333 out 0.0215186
R1604 out.n334 out 0.0215186
R1605 out.n335 out 0.0215186
R1606 out.n336 out 0.0215186
R1607 out.n337 out 0.0215186
R1608 out.n338 out 0.0215186
R1609 out.n339 out 0.0215186
R1610 out.n340 out 0.0215186
R1611 out out.n351 0.0215186
R1612 out out.n352 0.0215186
R1613 out out.n353 0.0215186
R1614 out out.n354 0.0215186
R1615 out out.n355 0.0215186
R1616 out out.n356 0.0215186
R1617 out out.n357 0.0215186
R1618 out out.n358 0.0215186
R1619 out out.n359 0.0215186
R1620 out out.n360 0.0215186
R1621 out out.n361 0.0215186
R1622 out out.n362 0.0215186
R1623 out out.n363 0.0215186
R1624 out out.n364 0.0215186
R1625 out out.n365 0.0215186
R1626 out out.n366 0.0215186
R1627 out out.n367 0.0215186
R1628 out out.n368 0.0215186
R1629 out out.n369 0.0215186
R1630 out out.n370 0.0215186
R1631 out out.n371 0.0215186
R1632 out out.n372 0.0215186
R1633 out out.n373 0.0215186
R1634 out out.n374 0.0215186
R1635 out out.n375 0.0215186
R1636 out out.n376 0.0215186
R1637 out out.n377 0.0215186
R1638 out out.n378 0.0215186
R1639 out out.n379 0.0215186
R1640 out out.n380 0.0215186
R1641 out out.n381 0.0215186
R1642 out out.n382 0.0215186
R1643 out.n398 out 0.0215186
R1644 out.n399 out 0.0215186
R1645 out.n400 out 0.0215186
R1646 out.n401 out 0.0215186
R1647 out.n402 out 0.0215186
R1648 out out.n60 0.0215186
R1649 out out.n61 0.0215186
R1650 out out.n62 0.0215186
R1651 out out.n63 0.0215186
R1652 out out.n64 0.0215186
R1653 out out.n65 0.0215186
R1654 out out.n66 0.0215186
R1655 out out.n67 0.0215186
R1656 out out.n68 0.0215186
R1657 out out.n69 0.0215186
R1658 out out.n70 0.0215186
R1659 out out.n71 0.0215186
R1660 out out.n72 0.0215186
R1661 out out.n73 0.0215186
R1662 out out.n74 0.0215186
R1663 out out.n75 0.0215186
R1664 out out.n76 0.0215186
R1665 out out.n77 0.0215186
R1666 out out.n78 0.0215186
R1667 out out.n79 0.0215186
R1668 out out.n80 0.0215186
R1669 out out.n81 0.0215186
R1670 out out.n82 0.0215186
R1671 out out.n83 0.0215186
R1672 out out.n84 0.0215186
R1673 out out.n85 0.0215186
R1674 out.n306 out 0.0193292
R1675 out.n384 out 0.0193292
R1676 out out.n341 0.0156801
R1677 out out.n342 0.0156801
R1678 out out.n343 0.0156801
R1679 out out.n344 0.0156801
R1680 out out.n345 0.0156801
R1681 out out.n346 0.0156801
R1682 out out.n347 0.0156801
R1683 out out.n348 0.0156801
R1684 out.n350 out 0.0150963
R1685 out.n397 out.n86 0.0139286
R1686 out.n392 out.n391 0.012177
R1687 out.n394 out.n393 0.012177
R1688 out.n305 out.n304 0.0118851
R1689 out.n386 out.n385 0.0110093
R1690 out.n388 out.n387 0.0110093
R1691 out.n390 out.n389 0.00954969
R1692 out.n396 out.n395 0.00925776
R1693 out.n395 out 0.00692236
R1694 out.n389 out 0.00663044
R1695 out.n385 out 0.00517081
R1696 out.n387 out 0.00517081
R1697 out.n304 out 0.00429503
R1698 out.n391 out 0.00400311
R1699 out.n393 out 0.00400311
R1700 out.n307 out.n306 0.00268944
R1701 out.n384 out.n383 0.00268944
R1702 out.n397 out 0.00225155
R1703 out.n350 out.n349 0.00108385
R1704 out.n87 out.t394 0.000500141
R1705 out.n88 out.t340 0.000500141
R1706 out.n89 out.t284 0.000500141
R1707 out.n90 out.t234 0.000500141
R1708 out.n91 out.t180 0.000500141
R1709 out.n92 out.t84 0.000500141
R1710 out.n93 out.t370 0.000500141
R1711 out.n94 out.t172 0.000500141
R1712 out.n95 out.t119 0.000500141
R1713 out.n96 out.t405 0.000500141
R1714 out.n97 out.t310 0.000500141
R1715 out.n98 out.t256 0.000500141
R1716 out.n99 out.t204 0.000500141
R1717 out.n100 out.t151 0.000500141
R1718 out.n101 out.t95 0.000500141
R1719 out.n102 out.t341 0.000500141
R1720 out.n103 out.t285 0.000500141
R1721 out.n104 out.t235 0.000500141
R1722 out.n105 out.t181 0.000500141
R1723 out.n106 out.t401 0.000500141
R1724 out.n107 out.t306 0.000500141
R1725 out.n108 out.t252 0.000500141
R1726 out.n109 out.t199 0.000500141
R1727 out.n110 out.t145 0.000500141
R1728 out.n111 out.t89 0.000500141
R1729 out.n112 out.t334 0.000500141
R1730 out.n113 out.t280 0.000500141
R1731 out.n114 out.t227 0.000500141
R1732 out.n115 out.t174 0.000500141
R1733 out.n116 out.t120 0.000500141
R1734 out.n117 out.t365 0.000500141
R1735 out.n118 out.t127 0.000500141
R1736 out.n119 out.t414 0.000500141
R1737 out.n120 out.t358 0.000500141
R1738 out.n121 out.t304 0.000500141
R1739 out.n122 out.t250 0.000500141
R1740 out.n123 out.t157 0.000500141
R1741 out.n124 out.t102 0.000500141
R1742 out.n125 out.t243 0.000500141
R1743 out.n126 out.t189 0.000500141
R1744 out.n127 out.t136 0.000500141
R1745 out.n128 out.t384 0.000500141
R1746 out.n129 out.t328 0.000500141
R1747 out.n130 out.t275 0.000500141
R1748 out.n131 out.t222 0.000500141
R1749 out.n132 out.t169 0.000500141
R1750 out.n133 out.t415 0.000500141
R1751 out.n134 out.t360 0.000500141
R1752 out.n135 out.t305 0.000500141
R1753 out.n136 out.t251 0.000500141
R1754 out.n137 out.t131 0.000500141
R1755 out.n138 out.t378 0.000500141
R1756 out.n139 out.t321 0.000500141
R1757 out.n140 out.t272 0.000500141
R1758 out.n141 out.t216 0.000500141
R1759 out.n142 out.t164 0.000500141
R1760 out.n143 out.t408 0.000500141
R1761 out.n144 out.t354 0.000500141
R1762 out.n145 out.t299 0.000500141
R1763 out.n146 out.t245 0.000500141
R1764 out.n147 out.t191 0.000500141
R1765 out.n148 out.t98 0.000500141
R1766 out.n149 out.t357 0.000500141
R1767 out.n150 out.t302 0.000500141
R1768 out.n151 out.t248 0.000500141
R1769 out.n152 out.t197 0.000500141
R1770 out.n153 out.t143 0.000500141
R1771 out.n154 out.t388 0.000500141
R1772 out.n155 out.t333 0.000500141
R1773 out.n156 out.t133 0.000500141
R1774 out.n157 out.t81 0.000500141
R1775 out.n158 out.t369 0.000500141
R1776 out.n159 out.t273 0.000500141
R1777 out.n160 out.t219 0.000500141
R1778 out.n161 out.t168 0.000500141
R1779 out.n162 out.t116 0.000500141
R1780 out.n163 out.t400 0.000500141
R1781 out.n164 out.t303 0.000500141
R1782 out.n165 out.t249 0.000500141
R1783 out.n166 out.t198 0.000500141
R1784 out.n167 out.t144 0.000500141
R1785 out.n168 out.t364 0.000500141
R1786 out.n169 out.t269 0.000500141
R1787 out.n170 out.t214 0.000500141
R1788 out.n171 out.t163 0.000500141
R1789 out.n172 out.t109 0.000500141
R1790 out.n173 out.t393 0.000500141
R1791 out.n174 out.t298 0.000500141
R1792 out.n175 out.t244 0.000500141
R1793 out.n176 out.t190 0.000500141
R1794 out.n177 out.t137 0.000500141
R1795 out.n178 out.t83 0.000500141
R1796 out.n179 out.t330 0.000500141
R1797 out.n180 out.t247 0.000500141
R1798 out.n181 out.t194 0.000500141
R1799 out.n182 out.t140 0.000500141
R1800 out.n183 out.t85 0.000500141
R1801 out.n184 out.t372 0.000500141
R1802 out.n185 out.t278 0.000500141
R1803 out.n186 out.t224 0.000500141
R1804 out.n187 out.t367 0.000500141
R1805 out.n188 out.t313 0.000500141
R1806 out.n189 out.t260 0.000500141
R1807 out.n190 out.t166 0.000500141
R1808 out.n191 out.t113 0.000500141
R1809 out.n192 out.t399 0.000500141
R1810 out.n193 out.t347 0.000500141
R1811 out.n194 out.t290 0.000500141
R1812 out.n195 out.t196 0.000500141
R1813 out.n196 out.t141 0.000500141
R1814 out.n197 out.t86 0.000500141
R1815 out.n198 out.t375 0.000500141
R1816 out.n199 out.t255 0.000500141
R1817 out.n200 out.t161 0.000500141
R1818 out.n201 out.t108 0.000500141
R1819 out.n202 out.t392 0.000500141
R1820 out.n203 out.t338 0.000500141
R1821 out.n204 out.t282 0.000500141
R1822 out.n205 out.t188 0.000500141
R1823 out.n206 out.t135 0.000500141
R1824 out.n207 out.t82 0.000500141
R1825 out.n208 out.t368 0.000500141
R1826 out.n209 out.t314 0.000500141
R1827 out.n210 out.t220 0.000500141
R1828 out.n211 out.t320 0.000500141
R1829 out.n212 out.t268 0.000500141
R1830 out.n213 out.t213 0.000500141
R1831 out.n214 out.t159 0.000500141
R1832 out.n215 out.t107 0.000500141
R1833 out.n216 out.t353 0.000500141
R1834 out.n217 out.t297 0.000500141
R1835 out.n218 out.t97 0.000500141
R1836 out.n219 out.t385 0.000500141
R1837 out.n220 out.t331 0.000500141
R1838 out.n221 out.t238 0.000500141
R1839 out.n222 out.t183 0.000500141
R1840 out.n223 out.t130 0.000500141
R1841 out.n224 out.t418 0.000500141
R1842 out.n225 out.t363 0.000500141
R1843 out.n226 out.t267 0.000500141
R1844 out.n227 out.t212 0.000500141
R1845 out.n228 out.t162 0.000500141
R1846 out.n229 out.t106 0.000500141
R1847 out.n230 out.t326 0.000500141
R1848 out.n231 out.t233 0.000500141
R1849 out.n232 out.t178 0.000500141
R1850 out.n233 out.t123 0.000500141
R1851 out.n234 out.t412 0.000500141
R1852 out.n235 out.t356 0.000500141
R1853 out.n236 out.t262 0.000500141
R1854 out.n237 out.t207 0.000500141
R1855 out.n238 out.t153 0.000500141
R1856 out.n239 out.t101 0.000500141
R1857 out.n240 out.t387 0.000500141
R1858 out.n241 out.t293 0.000500141
R1859 out.n242 out.t211 0.000500141
R1860 out.n243 out.t158 0.000500141
R1861 out.n244 out.t104 0.000500141
R1862 out.n245 out.t389 0.000500141
R1863 out.n246 out.t335 0.000500141
R1864 out.n247 out.t242 0.000500141
R1865 out.n248 out.t187 0.000500141
R1866 out.n249 out.t329 0.000500141
R1867 out.n250 out.t276 0.000500141
R1868 out.n251 out.t223 0.000500141
R1869 out.n252 out.t129 0.000500141
R1870 out.n253 out.t416 0.000500141
R1871 out.n254 out.t362 0.000500141
R1872 out.n255 out.t308 0.000500141
R1873 out.n256 out.t253 0.000500141
R1874 out.n257 out.t160 0.000500141
R1875 out.n258 out.t103 0.000500141
R1876 out.n259 out.t391 0.000500141
R1877 out.n260 out.t337 0.000500141
R1878 out.n261 out.t218 0.000500141
R1879 out.n262 out.t124 0.000500141
R1880 out.n263 out.t409 0.000500141
R1881 out.n264 out.t355 0.000500141
R1882 out.n265 out.t300 0.000500141
R1883 out.n266 out.t246 0.000500141
R1884 out.n267 out.t152 0.000500141
R1885 out.n268 out.t99 0.000500141
R1886 out.n269 out.t386 0.000500141
R1887 out.n270 out.t332 0.000500141
R1888 out.n271 out.t277 0.000500141
R1889 out.n272 out.t184 0.000500141
R1890 out.n273 out.t90 0.000500141
R1891 out.n274 out.t377 0.000500141
R1892 out.n275 out.t322 0.000500141
R1893 out.n276 out.t270 0.000500141
R1894 out.n277 out.t215 0.000500141
R1895 out.n278 out.t121 0.000500141
R1896 out.n279 out.t407 0.000500141
R1897 out.n280 out.t208 0.000500141
R1898 out.n281 out.t154 0.000500141
R1899 out.n282 out.t100 0.000500141
R1900 out.n283 out.t348 0.000500141
R1901 out.n284 out.t292 0.000500141
R1902 out.n285 out.t240 0.000500141
R1903 out.n286 out.t186 0.000500141
R1904 out.n287 out.t132 0.000500141
R1905 out.n288 out.t379 0.000500141
R1906 out.n289 out.t323 0.000500141
R1907 out.n290 out.t271 0.000500141
R1908 out.n291 out.t217 0.000500141
R1909 out.n292 out.t96 0.000500141
R1910 out.n293 out.t343 0.000500141
R1911 out.n294 out.t288 0.000500141
R1912 out.n295 out.t236 0.000500141
R1913 out.n296 out.t182 0.000500141
R1914 out.n297 out.t126 0.000500141
R1915 out.n298 out.t371 0.000500141
R1916 out.n299 out.t317 0.000500141
R1917 out.n300 out.t264 0.000500141
R1918 out.n301 out.t209 0.000500141
R1919 out.n302 out.t155 0.000500141
R1920 out.n303 out.t404 0.000500141
R1921 out.n305 out.t376 0.000500141
R1922 out.n307 out.t146 0.000500141
R1923 out.n308 out.t173 0.000500141
R1924 out.n309 out.t265 0.000500141
R1925 out.n310 out.t319 0.000500141
R1926 out.n311 out.t373 0.000500141
R1927 out.n312 out.t87 0.000500141
R1928 out.n313 out.t142 0.000500141
R1929 out.n314 out.t237 0.000500141
R1930 out.n315 out.t291 0.000500141
R1931 out.n316 out.t346 0.000500141
R1932 out.n317 out.t398 0.000500141
R1933 out.n318 out.t114 0.000500141
R1934 out.n319 out.t206 0.000500141
R1935 out.n320 out.t325 0.000500141
R1936 out.n321 out.t383 0.000500141
R1937 out.n322 out.t92 0.000500141
R1938 out.n323 out.t148 0.000500141
R1939 out.n324 out.t241 0.000500141
R1940 out.n325 out.t295 0.000500141
R1941 out.n326 out.t351 0.000500141
R1942 out.n327 out.t402 0.000500141
R1943 out.n328 out.t117 0.000500141
R1944 out.n329 out.t210 0.000500141
R1945 out.n330 out.t263 0.000500141
R1946 out.n331 out.t316 0.000500141
R1947 out.n332 out.t177 0.000500141
R1948 out.n333 out.t230 0.000500141
R1949 out.n334 out.t324 0.000500141
R1950 out.n335 out.t380 0.000500141
R1951 out.n336 out.t91 0.000500141
R1952 out.n337 out.t147 0.000500141
R1953 out.n338 out.t201 0.000500141
R1954 out.n339 out.t294 0.000500141
R1955 out.n340 out.t349 0.000500141
R1956 out.n341 out.t239 0.000500141
R1957 out.n342 out.t311 0.000500141
R1958 out.n343 out.t203 0.000500141
R1959 out.n344 out.t274 0.000500141
R1960 out.n345 out.t167 0.000500141
R1961 out.n346 out.t396 0.000500141
R1962 out.n347 out.t128 0.000500141
R1963 out.n348 out.t359 0.000500141
R1964 out.n349 out.t94 0.000500141
R1965 out.n351 out.t382 0.000500141
R1966 out.n352 out.t283 0.000500141
R1967 out.n353 out.t232 0.000500141
R1968 out.n354 out.t176 0.000500141
R1969 out.n355 out.t122 0.000500141
R1970 out.n356 out.t411 0.000500141
R1971 out.n357 out.t315 0.000500141
R1972 out.n358 out.t261 0.000500141
R1973 out.n359 out.t403 0.000500141
R1974 out.n360 out.t350 0.000500141
R1975 out.n361 out.t296 0.000500141
R1976 out.n362 out.t202 0.000500141
R1977 out.n363 out.t149 0.000500141
R1978 out.n364 out.t93 0.000500141
R1979 out.n365 out.t381 0.000500141
R1980 out.n366 out.t327 0.000500141
R1981 out.n367 out.t231 0.000500141
R1982 out.n368 out.t179 0.000500141
R1983 out.n369 out.t125 0.000500141
R1984 out.n370 out.t410 0.000500141
R1985 out.n371 out.t289 0.000500141
R1986 out.n372 out.t195 0.000500141
R1987 out.n373 out.t139 0.000500141
R1988 out.n374 out.t88 0.000500141
R1989 out.n375 out.t374 0.000500141
R1990 out.n376 out.t318 0.000500141
R1991 out.n377 out.t225 0.000500141
R1992 out.n378 out.t171 0.000500141
R1993 out.n379 out.t118 0.000500141
R1994 out.n380 out.t406 0.000500141
R1995 out.n381 out.t352 0.000500141
R1996 out.n382 out.t257 0.000500141
R1997 out.n383 out.t229 0.000500141
R1998 out.n386 out.t156 0.000500141
R1999 out.n388 out.t266 0.000500141
R2000 out.n390 out.t192 0.000500141
R2001 out.n392 out.t301 0.000500141
R2002 out.n394 out.t413 0.000500141
R2003 out.n396 out.t339 0.000500141
R2004 out.n86 out.t110 0.000500141
R2005 out.n398 out.t134 0.000500141
R2006 out.n399 out.t228 0.000500141
R2007 out.n400 out.t281 0.000500141
R2008 out.n401 out.t336 0.000500141
R2009 out.n402 out.t390 0.000500141
R2010 out.n60 out.t165 0.000500141
R2011 out.n61 out.t111 0.000500141
R2012 out.n62 out.t395 0.000500141
R2013 out.n63 out.t342 0.000500141
R2014 out.n64 out.t286 0.000500141
R2015 out.n65 out.t193 0.000500141
R2016 out.n66 out.t138 0.000500141
R2017 out.n67 out.t279 0.000500141
R2018 out.n68 out.t226 0.000500141
R2019 out.n69 out.t175 0.000500141
R2020 out.n70 out.t80 0.000500141
R2021 out.n71 out.t366 0.000500141
R2022 out.n72 out.t312 0.000500141
R2023 out.n73 out.t259 0.000500141
R2024 out.n74 out.t205 0.000500141
R2025 out.n75 out.t112 0.000500141
R2026 out.n76 out.t397 0.000500141
R2027 out.n77 out.t345 0.000500141
R2028 out.n78 out.t287 0.000500141
R2029 out.n79 out.t170 0.000500141
R2030 out.n80 out.t417 0.000500141
R2031 out.n81 out.t361 0.000500141
R2032 out.n82 out.t307 0.000500141
R2033 out.n83 out.t254 0.000500141
R2034 out.n84 out.t200 0.000500141
R2035 out.n85 out.t105 0.000500141
R2036 vdd.t100 vdd 895.586
R2037 vdd vdd.t115 895.586
R2038 vdd vdd.t106 895.586
R2039 vdd vdd.t103 895.586
R2040 vdd.n221 vdd.t89 584.644
R2041 vdd.n210 vdd.t61 584.644
R2042 vdd.n184 vdd.t145 584.644
R2043 vdd.n173 vdd.t43 584.644
R2044 vdd.n147 vdd.t74 584.644
R2045 vdd.n136 vdd.t130 584.644
R2046 vdd.n65 vdd.t121 584.644
R2047 vdd.n63 vdd.t12 584.644
R2048 vdd.n261 vdd.t101 459.192
R2049 vdd.n108 vdd.t116 459.192
R2050 vdd.n90 vdd.t107 459.192
R2051 vdd.n72 vdd.t104 459.192
R2052 vdd.n255 vdd 428.521
R2053 vdd.n254 vdd 428.521
R2054 vdd.n253 vdd 428.521
R2055 vdd.n252 vdd 428.521
R2056 vdd vdd.t97 378.64
R2057 vdd vdd.t94 378.64
R2058 vdd vdd.t112 378.64
R2059 vdd.n255 vdd.t100 340.096
R2060 vdd.t115 vdd.n254 340.096
R2061 vdd.t106 vdd.n253 340.096
R2062 vdd.t103 vdd.n252 340.096
R2063 vdd.t11 vdd 301.551
R2064 vdd vdd.t129 301.551
R2065 vdd vdd.t42 301.551
R2066 vdd vdd.t60 301.551
R2067 vdd.t5 vdd.n114 289.37
R2068 vdd.t140 vdd.n96 289.37
R2069 vdd.t30 vdd.n78 289.37
R2070 vdd.t54 vdd.n234 289.37
R2071 vdd.n119 vdd.t13 289.349
R2072 vdd.n101 vdd.t131 289.349
R2073 vdd.n83 vdd.t29 289.349
R2074 vdd.n239 vdd.t64 289.349
R2075 vdd.t120 vdd 285.68
R2076 vdd vdd.t73 285.68
R2077 vdd vdd.t144 285.68
R2078 vdd vdd.t88 285.68
R2079 vdd vdd.t109 247.137
R2080 vdd.t97 vdd 247.137
R2081 vdd.t94 vdd 247.137
R2082 vdd.t112 vdd 247.137
R2083 vdd.n68 vdd.t117 243.03
R2084 vdd.n70 vdd.t108 243.03
R2085 vdd.n250 vdd.t105 243.03
R2086 vdd.n256 vdd.t102 243.03
R2087 vdd.n205 vdd.t113 234.554
R2088 vdd.n208 vdd.t114 234.554
R2089 vdd.n168 vdd.t95 234.554
R2090 vdd.n171 vdd.t96 234.554
R2091 vdd.n131 vdd.t98 234.554
R2092 vdd.n134 vdd.t99 234.554
R2093 vdd.n0 vdd.t110 234.554
R2094 vdd.n3 vdd.t111 234.554
R2095 vdd.t18 vdd.t5 197.359
R2096 vdd.t6 vdd.t18 197.359
R2097 vdd.t14 vdd.t6 197.359
R2098 vdd.t15 vdd.t14 197.359
R2099 vdd.t4 vdd.t7 197.359
R2100 vdd.t10 vdd.t4 197.359
R2101 vdd.t19 vdd.t10 197.359
R2102 vdd.t13 vdd.t19 197.359
R2103 vdd.t132 vdd.t140 197.359
R2104 vdd.t141 vdd.t132 197.359
R2105 vdd.t133 vdd.t141 197.359
R2106 vdd.t124 vdd.t133 197.359
R2107 vdd.t139 vdd.t125 197.359
R2108 vdd.t128 vdd.t139 197.359
R2109 vdd.t138 vdd.t128 197.359
R2110 vdd.t131 vdd.t138 197.359
R2111 vdd.t44 vdd.t30 197.359
R2112 vdd.t38 vdd.t44 197.359
R2113 vdd.t31 vdd.t38 197.359
R2114 vdd.t45 vdd.t31 197.359
R2115 vdd.t28 vdd.t34 197.359
R2116 vdd.t41 vdd.t28 197.359
R2117 vdd.t37 vdd.t41 197.359
R2118 vdd.t29 vdd.t37 197.359
R2119 vdd.t62 vdd.t54 197.359
R2120 vdd.t55 vdd.t62 197.359
R2121 vdd.t65 vdd.t55 197.359
R2122 vdd.t56 vdd.t65 197.359
R2123 vdd.t63 vdd.t50 197.359
R2124 vdd.t59 vdd.t63 197.359
R2125 vdd.t53 vdd.t59 197.359
R2126 vdd.t64 vdd.t53 197.359
R2127 vdd.t16 vdd.t11 190.453
R2128 vdd.t8 vdd.t16 190.453
R2129 vdd.t20 vdd.t8 190.453
R2130 vdd.t71 vdd.t120 190.453
R2131 vdd.t22 vdd.t71 190.453
R2132 vdd.t84 vdd.t22 190.453
R2133 vdd.t129 vdd.t136 190.453
R2134 vdd.t136 vdd.t126 190.453
R2135 vdd.t126 vdd.t134 190.453
R2136 vdd.t73 vdd.t26 190.453
R2137 vdd.t26 vdd.t82 190.453
R2138 vdd.t82 vdd.t79 190.453
R2139 vdd.t42 vdd.t35 190.453
R2140 vdd.t35 vdd.t39 190.453
R2141 vdd.t39 vdd.t32 190.453
R2142 vdd.t144 vdd.t86 190.453
R2143 vdd.t86 vdd.t24 190.453
R2144 vdd.t24 vdd.t67 190.453
R2145 vdd.t60 vdd.t51 190.453
R2146 vdd.t51 vdd.t57 190.453
R2147 vdd.t57 vdd.t48 190.453
R2148 vdd.t88 vdd.t75 190.453
R2149 vdd.t75 vdd.t118 190.453
R2150 vdd.t118 vdd.t69 190.453
R2151 vdd.n252 vdd.n251 185
R2152 vdd.n253 vdd.n71 185
R2153 vdd.n254 vdd.n69 185
R2154 vdd.n257 vdd.n255 185
R2155 vdd.n226 vdd.n225 174.595
R2156 vdd.n215 vdd.n214 174.595
R2157 vdd.n189 vdd.n188 174.595
R2158 vdd.n178 vdd.n177 174.595
R2159 vdd.n152 vdd.n151 174.595
R2160 vdd.n141 vdd.n140 174.595
R2161 vdd.n271 vdd.n270 174.595
R2162 vdd.n280 vdd.n279 174.595
R2163 vdd vdd.t20 170.048
R2164 vdd vdd.t84 170.048
R2165 vdd.t134 vdd 170.048
R2166 vdd.t79 vdd 170.048
R2167 vdd.t32 vdd 170.048
R2168 vdd.t67 vdd 170.048
R2169 vdd.t48 vdd 170.048
R2170 vdd.t69 vdd 170.048
R2171 vdd.n206 vdd.t146 166.282
R2172 vdd.n169 vdd.t152 166.282
R2173 vdd.n132 vdd.t151 166.282
R2174 vdd.n1 vdd.t147 166.282
R2175 vdd.n20 vdd.t122 158.06
R2176 vdd.n18 vdd.t78 158.06
R2177 vdd.n16 vdd.t91 158.06
R2178 vdd.n14 vdd.t1 158.06
R2179 vdd.n13 vdd.t2 158.06
R2180 vdd.n11 vdd.t143 158.06
R2181 vdd.n9 vdd.t93 158.06
R2182 vdd.n7 vdd.t46 158.06
R2183 vdd.n5 vdd.t81 158.06
R2184 vdd.n21 vdd.t123 155.161
R2185 vdd.n12 vdd.t3 155.161
R2186 vdd.n10 vdd.t142 155.161
R2187 vdd.n8 vdd.t92 155.161
R2188 vdd.n6 vdd.t47 155.161
R2189 vdd.n19 vdd.t77 155.16
R2190 vdd.n17 vdd.t90 155.16
R2191 vdd.n15 vdd.t0 155.16
R2192 vdd.n4 vdd.t66 155.16
R2193 vdd.n230 vdd.t70 151.123
R2194 vdd.n220 vdd.t49 151.123
R2195 vdd.n193 vdd.t68 151.123
R2196 vdd.n183 vdd.t33 151.123
R2197 vdd.n156 vdd.t80 151.123
R2198 vdd.n146 vdd.t135 151.123
R2199 vdd.n66 vdd.t85 151.123
R2200 vdd.n64 vdd.t21 151.123
R2201 vdd.n116 vdd.t15 98.6801
R2202 vdd.t7 vdd.n116 98.6801
R2203 vdd.n98 vdd.t124 98.6801
R2204 vdd.t125 vdd.n98 98.6801
R2205 vdd.n80 vdd.t45 98.6801
R2206 vdd.t34 vdd.n80 98.6801
R2207 vdd.n236 vdd.t56 98.6801
R2208 vdd.t50 vdd.n236 98.6801
R2209 vdd.n261 vdd.t150 92.9047
R2210 vdd.n108 vdd.t153 92.9047
R2211 vdd.n90 vdd.t148 92.9047
R2212 vdd.n72 vdd.t149 92.9047
R2213 vdd.n59 vdd.n58 74.3398
R2214 vdd.n225 vdd.t76 26.5955
R2215 vdd.n225 vdd.t119 26.5955
R2216 vdd.n214 vdd.t52 26.5955
R2217 vdd.n214 vdd.t58 26.5955
R2218 vdd.n188 vdd.t87 26.5955
R2219 vdd.n188 vdd.t25 26.5955
R2220 vdd.n177 vdd.t36 26.5955
R2221 vdd.n177 vdd.t40 26.5955
R2222 vdd.n151 vdd.t27 26.5955
R2223 vdd.n151 vdd.t83 26.5955
R2224 vdd.n140 vdd.t137 26.5955
R2225 vdd.n140 vdd.t127 26.5955
R2226 vdd.n270 vdd.t72 26.5955
R2227 vdd.n270 vdd.t23 26.5955
R2228 vdd.n279 vdd.t17 26.5955
R2229 vdd.n279 vdd.t9 26.5955
R2230 vdd.n39 vdd.n12 25.224
R2231 vdd.n43 vdd.n10 25.224
R2232 vdd.n47 vdd.n8 25.224
R2233 vdd.n51 vdd.n6 25.224
R2234 vdd.n55 vdd.n4 25.224
R2235 vdd.n14 vdd.n13 21.8358
R2236 vdd.n210 vdd.n209 21.8029
R2237 vdd.n173 vdd.n172 21.8029
R2238 vdd.n136 vdd.n135 21.8029
R2239 vdd.n63 vdd.n62 21.8029
R2240 vdd.n221 vdd.n220 21.0829
R2241 vdd.n184 vdd.n183 21.0829
R2242 vdd.n147 vdd.n146 21.0829
R2243 vdd.n65 vdd.n64 21.0829
R2244 vdd.n18 vdd.n17 20.3299
R2245 vdd.n10 vdd.n9 20.3299
R2246 vdd.n8 vdd.n7 20.3299
R2247 vdd.n6 vdd.n5 20.3299
R2248 vdd.n20 vdd.n19 19.577
R2249 vdd.n12 vdd.n11 19.2005
R2250 vdd.n16 vdd.n15 18.824
R2251 vdd.n230 vdd.n76 15.4358
R2252 vdd.n193 vdd.n94 15.4358
R2253 vdd.n156 vdd.n112 15.4358
R2254 vdd.n265 vdd.n66 15.4358
R2255 vdd.n204 vdd.n77 14.2735
R2256 vdd.n167 vdd.n95 14.2735
R2257 vdd.n130 vdd.n113 14.2735
R2258 vdd.n124 vdd.n123 4.7293
R2259 vdd.n106 vdd.n105 4.7293
R2260 vdd.n88 vdd.n87 4.7293
R2261 vdd.n244 vdd.n243 4.7293
R2262 vdd.n57 vdd.n4 4.6505
R2263 vdd.n54 vdd.n5 4.6505
R2264 vdd.n53 vdd.n6 4.6505
R2265 vdd.n50 vdd.n7 4.6505
R2266 vdd.n49 vdd.n8 4.6505
R2267 vdd.n46 vdd.n9 4.6505
R2268 vdd.n45 vdd.n10 4.6505
R2269 vdd.n42 vdd.n11 4.6505
R2270 vdd.n41 vdd.n12 4.6505
R2271 vdd.n38 vdd.n13 4.6505
R2272 vdd.n37 vdd.n14 4.6505
R2273 vdd.n34 vdd.n15 4.6505
R2274 vdd.n33 vdd.n16 4.6505
R2275 vdd.n30 vdd.n17 4.6505
R2276 vdd.n29 vdd.n18 4.6505
R2277 vdd.n26 vdd.n19 4.6505
R2278 vdd.n25 vdd.n20 4.6505
R2279 vdd.n52 vdd.n51 4.6505
R2280 vdd.n48 vdd.n47 4.6505
R2281 vdd.n44 vdd.n43 4.6505
R2282 vdd.n40 vdd.n39 4.6505
R2283 vdd.n36 vdd.n35 4.6505
R2284 vdd.n32 vdd.n31 4.6505
R2285 vdd.n28 vdd.n27 4.6505
R2286 vdd.n24 vdd.n23 4.6505
R2287 vdd.n22 vdd.n21 4.6505
R2288 vdd.n56 vdd.n55 4.6505
R2289 vdd.n284 vdd.n63 4.6505
R2290 vdd.n276 vdd.n64 4.6505
R2291 vdd.n275 vdd.n65 4.6505
R2292 vdd.n267 vdd.n66 4.6505
R2293 vdd.n130 vdd.n129 4.6505
R2294 vdd.n137 vdd.n136 4.6505
R2295 vdd.n146 vdd.n145 4.6505
R2296 vdd.n148 vdd.n147 4.6505
R2297 vdd.n157 vdd.n156 4.6505
R2298 vdd.n167 vdd.n166 4.6505
R2299 vdd.n174 vdd.n173 4.6505
R2300 vdd.n183 vdd.n182 4.6505
R2301 vdd.n185 vdd.n184 4.6505
R2302 vdd.n194 vdd.n193 4.6505
R2303 vdd.n204 vdd.n203 4.6505
R2304 vdd.n211 vdd.n210 4.6505
R2305 vdd.n220 vdd.n219 4.6505
R2306 vdd.n222 vdd.n221 4.6505
R2307 vdd.n231 vdd.n230 4.6505
R2308 vdd.n62 vdd.n61 4.6505
R2309 vdd.n283 vdd.n282 4.6505
R2310 vdd.n281 vdd.n280 4.6505
R2311 vdd.n278 vdd.n277 4.6505
R2312 vdd.n274 vdd.n273 4.6505
R2313 vdd.n272 vdd.n271 4.6505
R2314 vdd.n269 vdd.n268 4.6505
R2315 vdd.n259 vdd.n258 4.6505
R2316 vdd.n139 vdd.n138 4.6505
R2317 vdd.n142 vdd.n141 4.6505
R2318 vdd.n144 vdd.n143 4.6505
R2319 vdd.n150 vdd.n149 4.6505
R2320 vdd.n153 vdd.n152 4.6505
R2321 vdd.n155 vdd.n154 4.6505
R2322 vdd.n161 vdd.n160 4.6505
R2323 vdd.n176 vdd.n175 4.6505
R2324 vdd.n179 vdd.n178 4.6505
R2325 vdd.n181 vdd.n180 4.6505
R2326 vdd.n187 vdd.n186 4.6505
R2327 vdd.n190 vdd.n189 4.6505
R2328 vdd.n192 vdd.n191 4.6505
R2329 vdd.n198 vdd.n197 4.6505
R2330 vdd.n213 vdd.n212 4.6505
R2331 vdd.n216 vdd.n215 4.6505
R2332 vdd.n218 vdd.n217 4.6505
R2333 vdd.n224 vdd.n223 4.6505
R2334 vdd.n227 vdd.n226 4.6505
R2335 vdd.n229 vdd.n228 4.6505
R2336 vdd.n249 vdd.n248 4.6505
R2337 vdd.n208 vdd.n207 4.36875
R2338 vdd.n171 vdd.n170 4.36875
R2339 vdd.n134 vdd.n133 4.36875
R2340 vdd.n3 vdd.n2 4.36875
R2341 vdd.n207 vdd.n206 3.50526
R2342 vdd.n170 vdd.n169 3.50526
R2343 vdd.n133 vdd.n132 3.50526
R2344 vdd.n2 vdd.n1 3.50526
R2345 vdd.n124 vdd 3.4052
R2346 vdd.n106 vdd 3.4052
R2347 vdd.n88 vdd 3.4052
R2348 vdd.n244 vdd 3.4052
R2349 vdd.n126 vdd.n125 3.23979
R2350 vdd.n163 vdd.n107 3.23979
R2351 vdd.n200 vdd.n89 3.23979
R2352 vdd.n246 vdd.n245 3.23979
R2353 vdd.n69 vdd.n68 3.08362
R2354 vdd.n71 vdd.n70 3.08362
R2355 vdd.n251 vdd.n250 3.08362
R2356 vdd.n257 vdd.n256 3.08362
R2357 vdd.n110 vdd.n108 2.61352
R2358 vdd.n92 vdd.n90 2.61352
R2359 vdd.n74 vdd.n72 2.61352
R2360 vdd.n263 vdd.n261 2.61352
R2361 vdd.n113 vdd.n67 2.29662
R2362 vdd.n162 vdd.n95 2.29662
R2363 vdd.n199 vdd.n77 2.29662
R2364 vdd.n110 vdd.n109 2.29594
R2365 vdd.n92 vdd.n91 2.29594
R2366 vdd.n74 vdd.n73 2.29594
R2367 vdd.n263 vdd.n262 2.29594
R2368 vdd.n123 vdd.n121 2.19925
R2369 vdd.n105 vdd.n103 2.19925
R2370 vdd.n87 vdd.n85 2.19925
R2371 vdd.n243 vdd.n241 2.19925
R2372 vdd.n112 vdd.n111 1.84013
R2373 vdd.n94 vdd.n93 1.84013
R2374 vdd.n76 vdd.n75 1.84013
R2375 vdd.n265 vdd.n264 1.84013
R2376 vdd.n158 vdd.n112 1.09272
R2377 vdd.n195 vdd.n94 1.09272
R2378 vdd.n232 vdd.n76 1.09272
R2379 vdd.n266 vdd.n265 1.09216
R2380 vdd.n206 vdd.n205 0.863992
R2381 vdd.n169 vdd.n168 0.863992
R2382 vdd.n132 vdd.n131 0.863992
R2383 vdd.n1 vdd.n0 0.863992
R2384 vdd.n123 vdd.n122 0.847933
R2385 vdd.n105 vdd.n104 0.847933
R2386 vdd.n87 vdd.n86 0.847933
R2387 vdd.n243 vdd.n242 0.847933
R2388 vdd.n111 vdd.n110 0.79957
R2389 vdd.n93 vdd.n92 0.79957
R2390 vdd.n75 vdd.n74 0.79957
R2391 vdd.n264 vdd.n263 0.79957
R2392 vdd.n125 vdd 0.783034
R2393 vdd.n107 vdd 0.783034
R2394 vdd.n89 vdd 0.783034
R2395 vdd.n245 vdd 0.783034
R2396 vdd.n58 vdd.n57 0.472161
R2397 vdd.n160 vdd.n69 0.467369
R2398 vdd.n197 vdd.n71 0.467369
R2399 vdd.n251 vdd.n249 0.467369
R2400 vdd.n258 vdd.n257 0.467369
R2401 vdd.n58 vdd 0.3755
R2402 vdd.n205 vdd.n204 0.305262
R2403 vdd.n209 vdd.n208 0.305262
R2404 vdd.n168 vdd.n167 0.305262
R2405 vdd.n172 vdd.n171 0.305262
R2406 vdd.n131 vdd.n130 0.305262
R2407 vdd.n135 vdd.n134 0.305262
R2408 vdd.n62 vdd.n3 0.305262
R2409 vdd.n159 vdd.n158 0.294492
R2410 vdd.n196 vdd.n195 0.294492
R2411 vdd.n233 vdd.n232 0.294492
R2412 vdd.n266 vdd.n260 0.294041
R2413 vdd.n158 vdd 0.234
R2414 vdd.n195 vdd 0.234
R2415 vdd.n232 vdd 0.234
R2416 vdd vdd.n266 0.231541
R2417 vdd.n259 vdd.n67 0.180551
R2418 vdd.n162 vdd.n161 0.180551
R2419 vdd.n199 vdd.n198 0.180551
R2420 vdd.n248 vdd.n247 0.180551
R2421 vdd.n119 vdd.n117 0.134074
R2422 vdd.n101 vdd.n99 0.134074
R2423 vdd.n83 vdd.n81 0.134074
R2424 vdd.n239 vdd.n237 0.134074
R2425 vdd.n56 vdd.n54 0.120292
R2426 vdd.n52 vdd.n50 0.120292
R2427 vdd.n48 vdd.n46 0.120292
R2428 vdd.n44 vdd.n42 0.120292
R2429 vdd.n40 vdd.n38 0.120292
R2430 vdd.n37 vdd.n36 0.120292
R2431 vdd.n36 vdd.n34 0.120292
R2432 vdd.n33 vdd.n32 0.120292
R2433 vdd.n32 vdd.n30 0.120292
R2434 vdd.n29 vdd.n28 0.120292
R2435 vdd.n28 vdd.n26 0.120292
R2436 vdd.n25 vdd.n24 0.120292
R2437 vdd.n24 vdd.n22 0.120292
R2438 vdd.n60 vdd.n59 0.120292
R2439 vdd.n61 vdd.n60 0.120292
R2440 vdd.n284 vdd.n283 0.120292
R2441 vdd.n283 vdd.n281 0.120292
R2442 vdd.n281 vdd.n278 0.120292
R2443 vdd.n278 vdd.n276 0.120292
R2444 vdd.n275 vdd.n274 0.120292
R2445 vdd.n274 vdd.n272 0.120292
R2446 vdd.n272 vdd.n269 0.120292
R2447 vdd.n269 vdd.n267 0.120292
R2448 vdd.n260 vdd.n259 0.120292
R2449 vdd.n129 vdd.n128 0.120292
R2450 vdd.n128 vdd.n127 0.120292
R2451 vdd.n139 vdd.n137 0.120292
R2452 vdd.n142 vdd.n139 0.120292
R2453 vdd.n144 vdd.n142 0.120292
R2454 vdd.n145 vdd.n144 0.120292
R2455 vdd.n150 vdd.n148 0.120292
R2456 vdd.n153 vdd.n150 0.120292
R2457 vdd.n155 vdd.n153 0.120292
R2458 vdd.n157 vdd.n155 0.120292
R2459 vdd.n161 vdd.n159 0.120292
R2460 vdd.n166 vdd.n165 0.120292
R2461 vdd.n165 vdd.n164 0.120292
R2462 vdd.n176 vdd.n174 0.120292
R2463 vdd.n179 vdd.n176 0.120292
R2464 vdd.n181 vdd.n179 0.120292
R2465 vdd.n182 vdd.n181 0.120292
R2466 vdd.n187 vdd.n185 0.120292
R2467 vdd.n190 vdd.n187 0.120292
R2468 vdd.n192 vdd.n190 0.120292
R2469 vdd.n194 vdd.n192 0.120292
R2470 vdd.n198 vdd.n196 0.120292
R2471 vdd.n203 vdd.n202 0.120292
R2472 vdd.n202 vdd.n201 0.120292
R2473 vdd.n213 vdd.n211 0.120292
R2474 vdd.n216 vdd.n213 0.120292
R2475 vdd.n218 vdd.n216 0.120292
R2476 vdd.n219 vdd.n218 0.120292
R2477 vdd.n224 vdd.n222 0.120292
R2478 vdd.n227 vdd.n224 0.120292
R2479 vdd.n229 vdd.n227 0.120292
R2480 vdd.n231 vdd.n229 0.120292
R2481 vdd.n248 vdd.n233 0.120292
R2482 vdd.n119 vdd.n118 0.11303
R2483 vdd.n101 vdd.n100 0.11303
R2484 vdd.n83 vdd.n82 0.11303
R2485 vdd.n239 vdd.n238 0.11303
R2486 vdd vdd.n56 0.0981562
R2487 vdd vdd.n52 0.0981562
R2488 vdd vdd.n48 0.0981562
R2489 vdd vdd.n44 0.0981562
R2490 vdd vdd.n40 0.0981562
R2491 vdd.n126 vdd.n67 0.0748257
R2492 vdd.n163 vdd.n162 0.0748257
R2493 vdd.n200 vdd.n199 0.0748257
R2494 vdd.n247 vdd.n246 0.0748257
R2495 vdd.n121 vdd.n120 0.0671871
R2496 vdd.n103 vdd.n102 0.0671871
R2497 vdd.n85 vdd.n84 0.0671871
R2498 vdd.n241 vdd.n240 0.0671871
R2499 vdd.n54 vdd 0.0603958
R2500 vdd vdd.n53 0.0603958
R2501 vdd.n50 vdd 0.0603958
R2502 vdd vdd.n49 0.0603958
R2503 vdd.n46 vdd 0.0603958
R2504 vdd vdd.n45 0.0603958
R2505 vdd.n42 vdd 0.0603958
R2506 vdd.n38 vdd 0.0603958
R2507 vdd vdd.n37 0.0603958
R2508 vdd vdd.n29 0.0603958
R2509 vdd vdd.n284 0.0603958
R2510 vdd.n129 vdd 0.0603958
R2511 vdd.n137 vdd 0.0603958
R2512 vdd.n166 vdd 0.0603958
R2513 vdd.n174 vdd 0.0603958
R2514 vdd.n203 vdd 0.0603958
R2515 vdd.n211 vdd 0.0603958
R2516 vdd vdd.n25 0.0577917
R2517 vdd vdd.n41 0.0564896
R2518 vdd vdd.n33 0.0551875
R2519 vdd vdd.n275 0.0512812
R2520 vdd.n148 vdd 0.0512812
R2521 vdd.n185 vdd 0.0512812
R2522 vdd.n222 vdd 0.0512812
R2523 vdd.n126 vdd 0.0255
R2524 vdd.n163 vdd 0.0255
R2525 vdd.n200 vdd 0.0255
R2526 vdd.n246 vdd 0.0255
R2527 vdd.n57 vdd 0.0226354
R2528 vdd.n53 vdd 0.0226354
R2529 vdd.n49 vdd 0.0226354
R2530 vdd.n45 vdd 0.0226354
R2531 vdd.n41 vdd 0.0226354
R2532 vdd.n34 vdd 0.0226354
R2533 vdd.n30 vdd 0.0226354
R2534 vdd.n26 vdd 0.0226354
R2535 vdd.n22 vdd 0.0226354
R2536 vdd.n61 vdd 0.0226354
R2537 vdd.n276 vdd 0.0226354
R2538 vdd.n267 vdd 0.0226354
R2539 vdd.n127 vdd 0.0226354
R2540 vdd.n145 vdd 0.0226354
R2541 vdd vdd.n157 0.0226354
R2542 vdd.n164 vdd 0.0226354
R2543 vdd.n182 vdd 0.0226354
R2544 vdd vdd.n194 0.0226354
R2545 vdd.n201 vdd 0.0226354
R2546 vdd.n219 vdd 0.0226354
R2547 vdd vdd.n231 0.0226354
R2548 vdd.n125 vdd.n124 0.0150548
R2549 vdd.n107 vdd.n106 0.0150548
R2550 vdd.n89 vdd.n88 0.0150548
R2551 vdd.n245 vdd.n244 0.0150548
R2552 vdd.n120 vdd.n119 0.0135311
R2553 vdd.n102 vdd.n101 0.0135311
R2554 vdd.n84 vdd.n83 0.0135311
R2555 vdd.n240 vdd.n239 0.0135311
R2556 vdd vdd.n126 0.0083125
R2557 vdd vdd.n163 0.0083125
R2558 vdd vdd.n200 0.0083125
R2559 vdd.n246 vdd 0.0083125
R2560 vdd.n116 vdd.n115 0.00492753
R2561 vdd.n98 vdd.n97 0.00492753
R2562 vdd.n80 vdd.n79 0.00492753
R2563 vdd.n236 vdd.n235 0.00492753
R2564 ctl_2_ ctl_2_.n0 50.4671
R2565 ctl_2_.n5 ctl_2_.t1 25.6264
R2566 ctl_2_.n0 ctl_2_.t2 24.9236
R2567 ctl_2_.n0 ctl_2_.t3 24.9236
R2568 ctl_2_.n4 ctl_2_.n3 15.7605
R2569 ctl_2_ ctl_2_.n1 11.2645
R2570 ctl_2_.n3 ctl_2_.t0 10.8355
R2571 ctl_2_.n14 ctl_2_.n13 9.50353
R2572 ctl_2_.n6 ctl_2_.n5 9.14032
R2573 ctl_2_.n15 ctl_2_.n14 6.78838
R2574 ctl_2_.n1 ctl_2_ 6.1445
R2575 ctl_2_.n1 ctl_2_ 4.65505
R2576 ctl_2_.n6 ctl_2_.n2 3.49141
R2577 ctl_2_.n13 ctl_2_.n12 3.49141
R2578 ctl_2_.n15 ctl_2_ 2.0485
R2579 ctl_2_ ctl_2_.n15 1.55202
R2580 ctl_2_.n5 ctl_2_.n4 0.968982
R2581 ctl_2_.n9 ctl_2_ 0.644086
R2582 ctl_2_.n12 ctl_2_.n6 0.194439
R2583 ctl_2_.n10 ctl_2_.n9 0.0569545
R2584 ctl_2_.n8 ctl_2_.n7 0.0356562
R2585 ctl_2_.n11 ctl_2_.n8 0.00245312
R2586 ctl_2_.n12 ctl_2_.n11 0.0011688
R2587 ctl_2_.n11 ctl_2_.n10 0.00100258
R2588 sky130_fd_sc_hd__inv_2_9.A.n1 sky130_fd_sc_hd__inv_2_9.A.t3 212.081
R2589 sky130_fd_sc_hd__inv_2_9.A.n2 sky130_fd_sc_hd__inv_2_9.A.t5 212.081
R2590 sky130_fd_sc_hd__inv_2_9.A.n1 sky130_fd_sc_hd__inv_2_9.A.t4 139.78
R2591 sky130_fd_sc_hd__inv_2_9.A.n2 sky130_fd_sc_hd__inv_2_9.A.t2 139.78
R2592 sky130_fd_sc_hd__inv_2_9.A.n2 sky130_fd_sc_hd__inv_2_9.A.n1 61.346
R2593 sky130_fd_sc_hd__inv_2_9.A.n3 sky130_fd_sc_hd__inv_2_9.A.n2 38.8554
R2594 sky130_fd_sc_hd__inv_2_9.A sky130_fd_sc_hd__inv_2_9.A.n3 4.85584
R2595 sky130_fd_sc_hd__inv_2_9.A.n3 sky130_fd_sc_hd__inv_2_9.A 1.99263
R2596 sky130_fd_sc_hd__inv_2_9.A.t1 sky130_fd_sc_hd__inv_2_9.A 0.197458
R2597 sky130_fd_sc_hd__inv_2_9.A.n0 sky130_fd_sc_hd__inv_2_9.A 0.18982
R2598 sky130_fd_sc_hd__inv_2_9.A sky130_fd_sc_hd__inv_2_9.A.t1 0.1012
R2599 sky130_fd_sc_hd__inv_2_9.A sky130_fd_sc_hd__inv_2_9.A.n0 0.0316375
R2600 sky130_fd_sc_hd__inv_2_9.A.t1 sky130_fd_sc_hd__inv_2_9.A 0.00959054
R2601 sky130_fd_sc_hd__inv_2_9.A sky130_fd_sc_hd__inv_2_9.A.t0 0.00959054
R2602 sample.n69 sample.t25 212.081
R2603 sample.n71 sample.t15 212.081
R2604 sample.n68 sample.t18 212.081
R2605 sample.n76 sample.t5 212.081
R2606 sample.n48 sample.t10 212.081
R2607 sample.n50 sample.t17 212.081
R2608 sample.n47 sample.t4 212.081
R2609 sample.n55 sample.t7 212.081
R2610 sample.n27 sample.t12 212.081
R2611 sample.n29 sample.t2 212.081
R2612 sample.n26 sample.t16 212.081
R2613 sample.n34 sample.t27 212.081
R2614 sample.n5 sample.t20 212.081
R2615 sample.n7 sample.t11 212.081
R2616 sample.n4 sample.t24 212.081
R2617 sample.n12 sample.t14 212.081
R2618 sample.n69 sample.t9 139.78
R2619 sample.n71 sample.t31 139.78
R2620 sample.n68 sample.t3 139.78
R2621 sample.n76 sample.t22 139.78
R2622 sample.n48 sample.t26 139.78
R2623 sample.n50 sample.t1 139.78
R2624 sample.n47 sample.t21 139.78
R2625 sample.n55 sample.t23 139.78
R2626 sample.n27 sample.t29 139.78
R2627 sample.n29 sample.t19 139.78
R2628 sample.n26 sample.t0 139.78
R2629 sample.n34 sample.t13 139.78
R2630 sample.n5 sample.t6 139.78
R2631 sample.n7 sample.t28 139.78
R2632 sample.n4 sample.t8 139.78
R2633 sample.n12 sample.t30 139.78
R2634 sample.n70 sample 78.3045
R2635 sample.n49 sample 78.3045
R2636 sample.n28 sample 78.3045
R2637 sample.n6 sample 78.3045
R2638 sample.n73 sample.n72 76.0005
R2639 sample.n75 sample.n74 76.0005
R2640 sample.n52 sample.n51 76.0005
R2641 sample.n54 sample.n53 76.0005
R2642 sample.n31 sample.n30 76.0005
R2643 sample.n33 sample.n32 76.0005
R2644 sample.n9 sample.n8 76.0005
R2645 sample.n11 sample.n10 76.0005
R2646 sample.n77 sample.n76 44.8017
R2647 sample.n56 sample.n55 44.8017
R2648 sample.n35 sample.n34 44.8017
R2649 sample.n13 sample.n12 44.8017
R2650 sample.n70 sample.n69 30.6732
R2651 sample.n71 sample.n70 30.6732
R2652 sample.n72 sample.n71 30.6732
R2653 sample.n72 sample.n68 30.6732
R2654 sample.n75 sample.n68 30.6732
R2655 sample.n76 sample.n75 30.6732
R2656 sample.n49 sample.n48 30.6732
R2657 sample.n50 sample.n49 30.6732
R2658 sample.n51 sample.n50 30.6732
R2659 sample.n51 sample.n47 30.6732
R2660 sample.n54 sample.n47 30.6732
R2661 sample.n55 sample.n54 30.6732
R2662 sample.n28 sample.n27 30.6732
R2663 sample.n29 sample.n28 30.6732
R2664 sample.n30 sample.n29 30.6732
R2665 sample.n30 sample.n26 30.6732
R2666 sample.n33 sample.n26 30.6732
R2667 sample.n34 sample.n33 30.6732
R2668 sample.n6 sample.n5 30.6732
R2669 sample.n7 sample.n6 30.6732
R2670 sample.n8 sample.n7 30.6732
R2671 sample.n8 sample.n4 30.6732
R2672 sample.n11 sample.n4 30.6732
R2673 sample.n12 sample.n11 30.6732
R2674 sample.n73 sample 19.2005
R2675 sample.n52 sample 19.2005
R2676 sample.n31 sample 19.2005
R2677 sample.n9 sample 19.2005
R2678 sample.n74 sample 17.1525
R2679 sample.n53 sample 17.1525
R2680 sample.n32 sample 17.1525
R2681 sample.n10 sample 17.1525
R2682 sample sample.n65 12.2885
R2683 sample sample.n44 12.2885
R2684 sample sample.n23 12.2885
R2685 sample sample.n2 12.2885
R2686 sample.n65 sample.n63 9.34456
R2687 sample.n44 sample.n42 9.34456
R2688 sample.n23 sample.n21 9.34456
R2689 sample.n77 sample.n64 9.3005
R2690 sample.n67 sample.n66 9.3005
R2691 sample.n56 sample.n43 9.3005
R2692 sample.n46 sample.n45 9.3005
R2693 sample.n35 sample.n22 9.3005
R2694 sample.n25 sample.n24 9.3005
R2695 sample.n66 sample.n62 9.01011
R2696 sample.n45 sample.n41 9.01011
R2697 sample.n24 sample.n20 9.01011
R2698 sample.n84 sample 8.66513
R2699 sample.n74 sample 6.4005
R2700 sample.n53 sample 6.4005
R2701 sample.n32 sample 6.4005
R2702 sample.n10 sample 6.4005
R2703 sample.n82 sample 6.20782
R2704 sample.n84 sample.n83 5.8694
R2705 sample.n83 sample.n82 5.85111
R2706 sample.n78 sample.n65 4.6085
R2707 sample.n77 sample.n67 4.6085
R2708 sample.n57 sample.n44 4.6085
R2709 sample.n56 sample.n46 4.6085
R2710 sample.n36 sample.n23 4.6085
R2711 sample.n35 sample.n25 4.6085
R2712 sample.n14 sample.n2 4.6085
R2713 sample.n13 sample.n3 4.6085
R2714 sample.n80 sample.n79 4.501
R2715 sample.n59 sample.n58 4.501
R2716 sample.n38 sample.n37 4.501
R2717 sample sample.n73 4.3525
R2718 sample sample.n52 4.3525
R2719 sample sample.n31 4.3525
R2720 sample sample.n9 4.3525
R2721 sample.n67 sample 1.7925
R2722 sample.n46 sample 1.7925
R2723 sample.n25 sample 1.7925
R2724 sample.n3 sample 1.7925
R2725 sample sample.n81 0.973061
R2726 sample sample.n19 0.973061
R2727 sample.n61 sample.n60 0.869402
R2728 sample.n40 sample.n39 0.845012
R2729 sample.n81 sample 0.767327
R2730 sample.n60 sample 0.767327
R2731 sample.n39 sample 0.767327
R2732 sample.n19 sample 0.767327
R2733 sample.n82 sample 0.338915
R2734 sample.n83 sample 0.338915
R2735 sample sample.n84 0.338915
R2736 sample.n78 sample.n77 0.2565
R2737 sample.n57 sample.n56 0.2565
R2738 sample.n36 sample.n35 0.2565
R2739 sample.n14 sample.n13 0.2565
R2740 sample.n40 sample 0.128549
R2741 sample sample.n40 0.122593
R2742 sample.n61 sample 0.104159
R2743 sample sample.n61 0.0993372
R2744 sample.n19 sample.n18 0.0775814
R2745 sample.n81 sample.n80 0.0501101
R2746 sample.n60 sample.n59 0.0501101
R2747 sample.n39 sample.n38 0.0501101
R2748 sample.n66 sample.n64 0.0437692
R2749 sample.n45 sample.n43 0.0437692
R2750 sample.n24 sample.n22 0.0437692
R2751 sample.n17 sample.n1 0.0437692
R2752 sample.n16 sample.n15 0.0437692
R2753 sample.n80 sample.n62 0.0286442
R2754 sample.n59 sample.n41 0.0286442
R2755 sample.n38 sample.n20 0.0286442
R2756 sample.n79 sample.n64 0.00290385
R2757 sample.n58 sample.n43 0.00290385
R2758 sample.n37 sample.n22 0.00290385
R2759 sample.n17 sample.n16 0.00290385
R2760 sample.n63 sample.n62 0.00216539
R2761 sample.n42 sample.n41 0.00216539
R2762 sample.n21 sample.n20 0.00216539
R2763 sample.n18 sample.n17 0.00166462
R2764 sample.n79 sample.n63 0.0015031
R2765 sample.n58 sample.n42 0.0015031
R2766 sample.n37 sample.n21 0.0015031
R2767 sample.n79 sample.n78 0.0011688
R2768 sample.n58 sample.n57 0.0011688
R2769 sample.n37 sample.n36 0.0011688
R2770 sample.n17 sample.n14 0.0011688
R2771 sample.n18 sample.n0 0.00100408
R2772 sky130_fd_sc_hd__inv_2_5.A.n1 sky130_fd_sc_hd__inv_2_5.A.t2 212.081
R2773 sky130_fd_sc_hd__inv_2_5.A.n2 sky130_fd_sc_hd__inv_2_5.A.t1 212.081
R2774 sky130_fd_sc_hd__inv_2_5.A.n4 sky130_fd_sc_hd__inv_2_5.A 152.388
R2775 sky130_fd_sc_hd__inv_2_5.A.n1 sky130_fd_sc_hd__inv_2_5.A.t4 139.78
R2776 sky130_fd_sc_hd__inv_2_5.A.n2 sky130_fd_sc_hd__inv_2_5.A.t3 139.78
R2777 sky130_fd_sc_hd__inv_2_5.A.n3 sky130_fd_sc_hd__inv_2_5.A.n0 73.3576
R2778 sky130_fd_sc_hd__inv_2_5.A.n2 sky130_fd_sc_hd__inv_2_5.A.n1 61.346
R2779 sky130_fd_sc_hd__inv_2_5.A.n3 sky130_fd_sc_hd__inv_2_5.A.n2 25.0059
R2780 sky130_fd_sc_hd__inv_2_5.A.n5 sky130_fd_sc_hd__inv_2_5.A.n4 9.3005
R2781 sky130_fd_sc_hd__inv_2_5.A.n6 sky130_fd_sc_hd__inv_2_5.A 8.80626
R2782 sky130_fd_sc_hd__inv_2_5.A.n4 sky130_fd_sc_hd__inv_2_5.A.n3 6.74837
R2783 sky130_fd_sc_hd__inv_2_5.A sky130_fd_sc_hd__inv_2_5.A.n5 4.08071
R2784 sky130_fd_sc_hd__inv_2_5.A sky130_fd_sc_hd__inv_2_5.A.n0 2.13383
R2785 sky130_fd_sc_hd__inv_2_5.A.n5 sky130_fd_sc_hd__inv_2_5.A.n0 0.776258
R2786 sky130_fd_sc_hd__inv_2_5.A sky130_fd_sc_hd__inv_2_5.A.t0 0.127353
R2787 sky130_fd_sc_hd__inv_2_5.A.n6 sky130_fd_sc_hd__inv_2_5.A 0.0465389
R2788 sky130_fd_sc_hd__inv_2_5.A.t0 sky130_fd_sc_hd__inv_2_5.A.n6 0.0388945
R2789 ctl_7_ ctl_7_.n0 50.4671
R2790 ctl_7_.n9 ctl_7_.t0 26.5955
R2791 ctl_7_.n9 ctl_7_.t1 26.5955
R2792 ctl_7_.n0 ctl_7_.t3 24.9236
R2793 ctl_7_.n0 ctl_7_.t2 24.9236
R2794 ctl_7_.n11 ctl_7_.n10 20.1729
R2795 ctl_7_ ctl_7_.n1 11.2645
R2796 ctl_7_.n10 ctl_7_.n9 8.28289
R2797 ctl_7_.n1 ctl_7_ 6.1445
R2798 ctl_7_.n1 ctl_7_ 4.65505
R2799 ctl_7_.n8 ctl_7_.n7 2.13383
R2800 ctl_7_.n11 ctl_7_ 2.0485
R2801 ctl_7_.n7 ctl_7_.n2 1.74595
R2802 ctl_7_ ctl_7_.n11 1.55202
R2803 ctl_7_.n4 ctl_7_ 0.53918
R2804 ctl_7_.n10 ctl_7_.n8 0.482005
R2805 ctl_7_.n5 ctl_7_.n4 0.0569555
R2806 ctl_7_.n6 ctl_7_.n3 0.0180781
R2807 ctl_7_.n7 ctl_7_.n6 0.00116875
R2808 ctl_7_.n6 ctl_7_.n5 0.00100158
R2809 ctl_3_ ctl_3_.n0 50.4671
R2810 ctl_3_.n2 ctl_3_.t1 26.5955
R2811 ctl_3_.n3 ctl_3_.t0 25.8979
R2812 ctl_3_.n0 ctl_3_.t3 24.9236
R2813 ctl_3_.n0 ctl_3_.t2 24.9236
R2814 ctl_3_ ctl_3_.n1 11.2645
R2815 ctl_3_.n11 ctl_3_.n10 9.11565
R2816 ctl_3_.n4 ctl_3_.n3 8.39596
R2817 ctl_3_.n12 ctl_3_.n11 6.78838
R2818 ctl_3_.n1 ctl_3_ 6.1445
R2819 ctl_3_.n1 ctl_3_ 4.65505
R2820 ctl_3_.n10 ctl_3_.n9 3.29747
R2821 ctl_3_.n12 ctl_3_ 2.0485
R2822 ctl_3_ ctl_3_.n12 1.55202
R2823 ctl_3_.n6 ctl_3_ 0.672135
R2824 ctl_3_.n9 ctl_3_.n4 0.582318
R2825 ctl_3_.n3 ctl_3_.n2 0.240912
R2826 ctl_3_.n7 ctl_3_.n6 0.0569547
R2827 ctl_3_.n8 ctl_3_.n5 0.00635938
R2828 ctl_3_.n9 ctl_3_.n8 0.0011688
R2829 ctl_3_.n8 ctl_3_.n7 0.00100244
R2830 ctl_4_ ctl_4_.n0 50.4671
R2831 ctl_4_.n2 ctl_4_.t0 26.5955
R2832 ctl_4_.n2 ctl_4_.t1 26.5955
R2833 ctl_4_.n0 ctl_4_.t3 24.9236
R2834 ctl_4_.n0 ctl_4_.t2 24.9236
R2835 ctl_4_ ctl_4_.n1 11.2645
R2836 ctl_4_.n12 ctl_4_.n11 9.50353
R2837 ctl_4_.n3 ctl_4_.n2 8.78779
R2838 ctl_4_.n13 ctl_4_.n12 6.78838
R2839 ctl_4_.n1 ctl_4_ 6.1445
R2840 ctl_4_.n1 ctl_4_ 4.65505
R2841 ctl_4_.n11 ctl_4_.n10 3.49141
R2842 ctl_4_.n13 ctl_4_ 2.0485
R2843 ctl_4_ ctl_4_.n13 1.55202
R2844 ctl_4_.n7 ctl_4_ 0.66276
R2845 ctl_4_.n10 ctl_4_.n4 0.194439
R2846 ctl_4_.n4 ctl_4_.n3 0.102503
R2847 ctl_4_.n8 ctl_4_.n7 0.0569545
R2848 ctl_4_.n6 ctl_4_.n5 0.0356562
R2849 ctl_4_.n9 ctl_4_.n6 0.00245312
R2850 ctl_4_.n10 ctl_4_.n9 0.00116875
R2851 ctl_4_.n9 ctl_4_.n8 0.00100258
R2852 dum dum.n0 50.4671
R2853 dum.n3 dum.t0 26.5955
R2854 dum.n4 dum.t1 25.8861
R2855 dum.n0 dum.t3 24.9236
R2856 dum.n0 dum.t2 24.9236
R2857 dum dum.n1 11.2645
R2858 dum.n11 dum.n10 9.50353
R2859 dum.n9 dum.n4 8.76736
R2860 dum.n12 dum.n11 6.78838
R2861 dum.n1 dum 6.1445
R2862 dum.n1 dum 4.65505
R2863 dum.n10 dum.n9 3.68535
R2864 dum.n9 dum.n2 3.49141
R2865 dum.n12 dum 2.0485
R2866 dum dum.n12 1.55202
R2867 dum.n6 dum 0.659635
R2868 dum.n4 dum.n3 0.251928
R2869 dum.n7 dum.n6 0.0569544
R2870 dum.n8 dum.n5 0.0356562
R2871 dum.n9 dum.n8 0.00116875
R2872 dum.n8 dum.n7 0.00100273
R2873 ctl_1_ ctl_1_.n0 50.4671
R2874 ctl_1_.n10 ctl_1_.t1 26.5955
R2875 ctl_1_.n10 ctl_1_.t0 26.5955
R2876 ctl_1_.n0 ctl_1_.t2 24.9236
R2877 ctl_1_.n0 ctl_1_.t3 24.9236
R2878 ctl_1_ ctl_1_.n1 11.2645
R2879 ctl_1_.n13 ctl_1_.n12 9.69747
R2880 ctl_1_.n11 ctl_1_.n10 9.15497
R2881 ctl_1_.n14 ctl_1_.n13 6.78838
R2882 ctl_1_.n1 ctl_1_ 6.1445
R2883 ctl_1_.n1 ctl_1_ 4.65505
R2884 ctl_1_.n12 ctl_1_.n11 3.49141
R2885 ctl_1_.n9 ctl_1_.n2 3.29747
R2886 ctl_1_.n14 ctl_1_ 2.0485
R2887 ctl_1_ ctl_1_.n14 1.55202
R2888 ctl_1_.n6 ctl_1_ 0.63494
R2889 ctl_1_.n11 ctl_1_.n9 0.388379
R2890 ctl_1_.n7 ctl_1_.n6 0.0557885
R2891 ctl_1_.n5 ctl_1_.n4 0.0356562
R2892 ctl_1_.n8 ctl_1_.n3 0.0337031
R2893 ctl_1_.n8 ctl_1_.n5 0.00440625
R2894 ctl_1_.n9 ctl_1_.n8 0.0011688
R2895 ctl_1_.n8 ctl_1_.n7 0.0011687
R2896 ctl_5_ ctl_5_.n0 50.4671
R2897 ctl_5_.n2 ctl_5_.t1 26.5955
R2898 ctl_5_.n2 ctl_5_.t0 26.5955
R2899 ctl_5_.n0 ctl_5_.t3 24.9236
R2900 ctl_5_.n0 ctl_5_.t2 24.9236
R2901 ctl_5_ ctl_5_.n1 11.2645
R2902 ctl_5_.n10 ctl_5_.n9 9.50353
R2903 ctl_5_.n3 ctl_5_.n2 8.78779
R2904 ctl_5_.n11 ctl_5_.n10 6.78838
R2905 ctl_5_.n1 ctl_5_ 6.1445
R2906 ctl_5_.n1 ctl_5_ 4.65505
R2907 ctl_5_.n9 ctl_5_.n8 3.68535
R2908 ctl_5_.n11 ctl_5_ 2.0485
R2909 ctl_5_ ctl_5_.n11 1.55202
R2910 ctl_5_.n5 ctl_5_ 0.659635
R2911 ctl_5_.n8 ctl_5_.n3 0.102503
R2912 ctl_5_.n6 ctl_5_.n5 0.0569544
R2913 ctl_5_.n7 ctl_5_.n4 0.0356562
R2914 ctl_5_.n8 ctl_5_.n7 0.0011687
R2915 ctl_5_.n7 ctl_5_.n6 0.00100273
R2916 ctl_0_ ctl_0_.n0 50.4671
R2917 ctl_0_.n8 ctl_0_.t1 26.5955
R2918 ctl_0_.n9 ctl_0_.t0 25.8861
R2919 ctl_0_.n0 ctl_0_.t3 24.9236
R2920 ctl_0_.n0 ctl_0_.t2 24.9236
R2921 ctl_0_ ctl_0_.n1 11.2645
R2922 ctl_0_.n12 ctl_0_.n11 10.0491
R2923 ctl_0_.n11 ctl_0_.n10 9.81841
R2924 ctl_0_.n10 ctl_0_.n9 8.76736
R2925 ctl_0_.n1 ctl_0_ 6.1445
R2926 ctl_0_.n1 ctl_0_ 4.65505
R2927 ctl_0_.n7 ctl_0_.n2 3.10353
R2928 ctl_0_.n12 ctl_0_ 2.0485
R2929 ctl_0_ ctl_0_.n12 1.55202
R2930 ctl_0_.n10 ctl_0_.n7 0.776258
R2931 ctl_0_.n4 ctl_0_ 0.647135
R2932 ctl_0_.n9 ctl_0_.n8 0.251928
R2933 ctl_0_.n5 ctl_0_.n4 0.0569565
R2934 ctl_0_.n6 ctl_0_.n3 0.03175
R2935 ctl_0_.n7 ctl_0_.n6 0.0011688
R2936 ctl_0_.n6 ctl_0_.n5 0.00100057
C0 sky130_fd_sc_hd__inv_2_0.A ctl_4_ 1.81e-20
C1 carray_0.unitcap_23.cn carray_0.unitcap_31.cn 0.0902f
C2 vin sample 0.0186f
C3 sky130_fd_sc_hd__inv_2_6.A ctl_7_ 3.29e-20
C4 carray_0.unitcap_0.cn out 0.514f
C5 vin vdd 2.51f
C6 sky130_fd_sc_hd__inv_2_7.A sky130_fd_sc_hd__inv_2_3.A 0.251f
C7 out carray_0.unitcap_71.cn 0.51f
C8 sky130_fd_sc_hd__inv_2_4.A carray_0.unitcap_334.cn 0.0418f
C9 sky130_fd_sc_hd__inv_2_4.A vdd 0.215f
C10 sky130_fd_sc_hd__inv_2_2.VPB carray_0.unitcap_331.cn 0.0021f
C11 ctl_4_ ctl_7_ 4.45e-20
C12 ctl_5_ ctl_6_ 0.0689f
C13 carray_0.unitcap_0.cn carray_0.unitcap_40.cn 0.0902f
C14 ctl_0_ dum 0.0679f
C15 carray_0.unitcap_175.cn vdd 0.00397f
C16 sky130_fd_sc_hd__inv_2_9.A sample 3.19f
C17 carray_0.unitcap_8.cn out 0.503f
C18 carray_0.unitcap_71.cn carray_0.unitcap_95.cn 0.0902f
C19 sky130_fd_sc_hd__inv_2_7.A ctl_3_ 0.109f
C20 sky130_fd_sc_hd__inv_2_9.A vdd 3.83f
C21 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_338.cn 0.161f
C22 sw_top_1.en_buf sw_top_2.en_buf 0.00273f
C23 carray_0.unitcap_240.cn carray_0.unitcap_232.cn 0.0902f
C24 carray_0.unitcap_13.cn vin 0.198f
C25 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_215.cn 0.161f
C26 sky130_fd_sc_hd__inv_2_3.A ctl_3_ 5.77e-20
C27 carray_0.unitcap_331.cn ctl_6_ 0.00225f
C28 sw_top_1.en_buf carray_0.unitcap_80.cn 3.18e-20
C29 vdd sample 1.47f
C30 carray_0.unitcap_63.cn carray_0.unitcap_55.cn 0.0902f
C31 carray_0.unitcap_47.cn vin 4.46e-19
C32 sw_top_2.net1 out 0.396f
C33 carray_0.unitcap_11.cn carray_0.unitcap_10.cn 0.18f
C34 sw_top_3.net1 sw_top_2.net1 0.00267f
C35 carray_0.unitcap_334.cn vdd 0.00423f
C36 vdd carray_0.unitcap_338.cn 0.00397f
C37 carray_0.unitcap_337.cn sky130_fd_sc_hd__inv_2_6.A 0.0902f
C38 sky130_fd_sc_hd__inv_2_0.A out 35.4f
C39 sky130_fd_sc_hd__inv_2_2.A dum 0.0966f
C40 carray_0.unitcap_8.cn carray_0.unitcap_16.cn 0.0902f
C41 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_13.cn 0.0902f
C42 sky130_fd_sc_hd__inv_2_7.A ctl_5_ 3.21e-20
C43 carray_0.unitcap_215.cn vdd 0.00397f
C44 ctl_0_ ctl_1_ 0.0679f
C45 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_207.cn 0.161f
C46 out ctl_7_ 0.00175f
C47 carray_0.unitcap_87.cn vin 4.46e-19
C48 sky130_fd_sc_hd__inv_2_8.A carray_0.unitcap_322.cn 0.277f
C49 sky130_fd_sc_hd__inv_2_3.A ctl_5_ 3.18e-21
C50 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_47.cn 0.18f
C51 out carray_0.unitcap_111.cn 0.51f
C52 sky130_fd_sc_hd__inv_2_0.A sky130_fd_sc_hd__inv_2_5.A 2.27f
C53 carray_0.unitcap_322.cn out 0.502f
C54 carray_0.unitcap_31.cn out 0.51f
C55 carray_0.unitcap_207.cn vdd 0.00397f
C56 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_87.cn 0.18f
C57 ctl_3_ ctl_5_ 4.43e-20
C58 sky130_fd_sc_hd__inv_2_5.A ctl_7_ 3.04e-19
C59 carray_0.unitcap_95.cn carray_0.unitcap_111.cn 0.0902f
C60 carray_0.unitcap_255.cn carray_0.unitcap_239.cn 0.0902f
C61 carray_0.unitcap_328.cn ctl_0_ 0.00143f
C62 sky130_fd_sc_hd__inv_2_2.A ctl_1_ 1.05e-20
C63 sky130_fd_sc_hd__inv_2_2.VPB ctl_0_ 0.0101f
C64 carray_0.unitcap_128.cn out 0.514f
C65 carray_0.unitcap_96.cn carray_0.unitcap_120.cn 0.0902f
C66 carray_0.unitcap_216.cn carray_0.unitcap_240.cn 0.0902f
C67 carray_0.unitcap_330.cn carray_0.unitcap_331.cn 0.18f
C68 carray_0.unitcap_9.cn carray_0.unitcap_8.cn 0.18f
C69 carray_0.unitcap_63.cn vin 4.46e-19
C70 carray_0.unitcap_337.cn out 0.505f
C71 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_72.cn 0.18f
C72 ctl_0_ ctl_6_ 3.69e-22
C73 carray_0.unitcap_248.cn out 0.514f
C74 carray_0.unitcap_288.cn out 0.558f
C75 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_63.cn 0.18f
C76 sky130_fd_sc_hd__inv_2_2.A carray_0.unitcap_328.cn 0.00374f
C77 carray_0.unitcap_224.cn out 0.514f
C78 carray_0.unitcap_103.cn out 0.51f
C79 carray_0.unitcap_72.cn sample 0.00155f
C80 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_sc_hd__inv_2_2.A 0.0813f
C81 out carray_0.unitcap_151.cn 0.51f
C82 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_135.cn 0.161f
C83 carray_0.unitcap_72.cn vdd 2.17e-20
C84 carray_0.unitcap_23.cn vin 4.46e-19
C85 sky130_fd_sc_hd__inv_2_4.A ctl_2_ 2.12e-20
C86 ctl_5_ carray_0.unitcap_331.cn 0.00261f
C87 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_112.cn 0.18f
C88 sw_top_1.net1 sw_top_0.en_buf 2.34e-19
C89 carray_0.unitcap_256.cn carray_0.unitcap_288.cn 0.18f
C90 sky130_fd_sc_hd__inv_2_4.A carray_0.unitcap_247.cn 0.18f
C91 sw_top_1.en_buf sw_top_2.net1 2.34e-19
C92 carray_0.unitcap_55.cn out 0.514f
C93 carray_0.unitcap_224.cn sky130_fd_sc_hd__inv_2_5.A 0.18f
C94 sky130_fd_sc_hd__inv_2_6.A sky130_fd_sc_hd__inv_2_4.A 0.227f
C95 sky130_fd_sc_hd__inv_2_0.A ctl_1_ 1.74e-21
C96 sky130_fd_sc_hd__inv_2_9.A ctl_2_ 8.15e-22
C97 vin sw_top_0.en_buf 0.448f
C98 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_152.cn 0.18f
C99 carray_0.unitcap_135.cn vdd 0.00397f
C100 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_23.cn 0.18f
C101 carray_0.unitcap_144.cn out 0.514f
C102 carray_0.unitcap_31.cn carray_0.unitcap_7.cn 0.0902f
C103 sky130_fd_sc_hd__inv_2_7.A ctl_0_ 1.81e-20
C104 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_247.cn 0.161f
C105 ctl_1_ ctl_7_ 5.64e-20
C106 sky130_fd_sc_hd__inv_2_4.A ctl_4_ 0.0998f
C107 sky130_fd_sc_hd__inv_2_6.A sky130_fd_sc_hd__inv_2_9.A 0.135f
C108 ctl_2_ vdd 0.269f
C109 sky130_fd_sc_hd__inv_2_3.A ctl_0_ 0.0384f
C110 sky130_fd_sc_hd__inv_2_9.A sw_top_0.en_buf 0.867f
C111 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_64.cn 0.18f
C112 carray_0.unitcap_56.cn out 0.514f
C113 sky130_fd_sc_hd__inv_2_9.A ctl_4_ 2.07e-21
C114 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_24.cn 0.18f
C115 vdd carray_0.unitcap_247.cn 0.00397f
C116 carray_0.unitcap_104.cn out 0.514f
C117 sky130_fd_sc_hd__inv_2_0.A sky130_fd_sc_hd__inv_2_2.VPB 0.0805f
C118 sample sw_top_0.en_buf 0.408f
C119 carray_0.unitcap_119.cn out 0.51f
C120 sky130_fd_sc_hd__inv_2_6.A vdd 0.146f
C121 sky130_fd_sc_hd__inv_2_6.A carray_0.unitcap_334.cn 0.348f
C122 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_167.cn 0.18f
C123 carray_0.unitcap_64.cn sample 0.00149f
C124 out carray_0.unitcap_183.cn 0.51f
C125 sky130_fd_sc_hd__inv_2_6.A carray_0.unitcap_338.cn 0.18f
C126 ctl_3_ ctl_0_ 2.11e-20
C127 carray_0.unitcap_231.cn carray_0.unitcap_223.cn 0.0902f
C128 carray_0.unitcap_232.cn carray_0.unitcap_248.cn 0.0902f
C129 vdd sw_top_0.en_buf 1.84f
C130 carray_0.unitcap_24.cn sample 0.00149f
C131 carray_0.unitcap_64.cn vdd 1.93e-19
C132 sky130_fd_sc_hd__inv_2_2.A sky130_fd_sc_hd__inv_2_7.A 0.0925f
C133 sky130_fd_sc_hd__inv_2_2.VPB ctl_7_ 0.0103f
C134 carray_0.unitcap_128.cn carray_0.unitcap_152.cn 0.0902f
C135 carray_0.unitcap_334.cn ctl_4_ 0.00253f
C136 ctl_4_ vdd 0.268f
C137 sw_top_1.net1 out 0.381f
C138 carray_0.unitcap_24.cn vdd 3.66e-20
C139 carray_0.unitcap_208.cn carray_0.unitcap_224.cn 0.0902f
C140 sky130_fd_sc_hd__inv_2_4.A sky130_fd_sc_hd__inv_2_8.A 1.66e-19
C141 carray_0.unitcap_32.cn carray_0.unitcap_56.cn 0.0902f
C142 out carray_0.unitcap_160.cn 0.514f
C143 carray_0.unitcap_322.cn carray_0.unitcap_328.cn 0.18f
C144 sky130_fd_sc_hd__inv_2_2.A sky130_fd_sc_hd__inv_2_3.A 0.0424f
C145 vin out 10.3f
C146 sw_top_3.net1 vin 0.392f
C147 sw_top_3.en_buf sw_top_2.en_buf 0.00273f
C148 sky130_fd_sc_hd__inv_2_0.A ctl_6_ 0.0994f
C149 sky130_fd_sc_hd__inv_2_4.A out 8.83f
C150 ctl_5_ ctl_0_ 1.88e-21
C151 carray_0.unitcap_175.cn out 0.51f
C152 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_192.cn 0.18f
C153 ctl_7_ ctl_6_ 0.0628f
C154 sky130_fd_sc_hd__inv_2_2.A ctl_3_ 9.56e-21
C155 sky130_fd_sc_hd__inv_2_9.A out 79.6f
C156 sky130_fd_sc_hd__inv_2_9.A sw_top_3.net1 0.484f
C157 sky130_fd_sc_hd__inv_2_4.A sky130_fd_sc_hd__inv_2_5.A 1.35f
C158 sky130_fd_sc_hd__inv_2_8.A vdd 0.0977f
C159 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_40.cn 0.18f
C160 sample out 0.306f
C161 sw_top_3.net1 sample 0.0344f
C162 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_95.cn 0.18f
C163 carray_0.unitcap_334.cn out 0.501f
C164 sw_top_3.net1 vdd 0.824f
C165 vdd out 2.98f
C166 sky130_fd_sc_hd__inv_2_9.A sky130_fd_sc_hd__inv_2_5.A 0.552f
C167 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_256.cn 0.0902f
C168 carray_0.unitcap_338.cn out 0.51f
C169 sky130_fd_sc_hd__inv_2_0.A sky130_fd_sc_hd__inv_2_7.A 0.325f
C170 carray_0.unitcap_40.cn sample 0.00149f
C171 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_32.cn 0.18f
C172 carray_0.unitcap_215.cn out 0.51f
C173 carray_0.unitcap_152.cn carray_0.unitcap_144.cn 0.0902f
C174 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_16.cn 0.18f
C175 carray_0.unitcap_103.cn carray_0.unitcap_127.cn 0.0902f
C176 carray_0.unitcap_224.cn carray_0.unitcap_216.cn 0.0902f
C177 carray_0.unitcap_40.cn vdd 1.17e-20
C178 sky130_fd_sc_hd__inv_2_0.A sky130_fd_sc_hd__inv_2_3.A 8.44e-21
C179 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_176.cn 0.18f
C180 carray_0.unitcap_256.cn sample 0.107f
C181 out carray_0.unitcap_168.cn 0.514f
C182 carray_0.unitcap_151.cn carray_0.unitcap_167.cn 0.0902f
C183 sky130_fd_sc_hd__inv_2_7.A ctl_7_ 2.42e-20
C184 carray_0.unitcap_320.cn carray_0.unitcap_324.cn 0.18f
C185 carray_0.unitcap_14.cn vin 0.00323f
C186 carray_0.unitcap_32.cn sample 0.00149f
C187 sky130_fd_sc_hd__inv_2_5.A vdd 1.05f
C188 sky130_fd_sc_hd__inv_2_4.A dum 1.8e-21
C189 sample carray_0.unitcap_16.cn 0.00149f
C190 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_330.cn 0.149f
C191 vdd carray_0.unitcap_32.cn 2.58e-19
C192 sky130_fd_sc_hd__inv_2_3.A ctl_7_ 5.64e-21
C193 carray_0.unitcap_13.cn out 0.558f
C194 sky130_fd_sc_hd__inv_2_7.A carray_0.unitcap_322.cn 8.85e-20
C195 sky130_fd_sc_hd__inv_2_5.A carray_0.unitcap_215.cn 0.18f
C196 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_199.cn 0.18f
C197 carray_0.unitcap_207.cn out 0.51f
C198 sky130_fd_sc_hd__inv_2_0.A ctl_3_ 1.11e-20
C199 sky130_fd_sc_hd__inv_2_4.A carray_0.unitcap_232.cn 0.18f
C200 carray_0.unitcap_47.cn out 0.514f
C201 carray_0.unitcap_330.cn ctl_7_ 6.04e-19
C202 sky130_fd_sc_hd__inv_2_3.A carray_0.unitcap_322.cn 0.121f
C203 carray_0.unitcap_14.cn sky130_fd_sc_hd__inv_2_9.A 0.0902f
C204 carray_0.unitcap_7.cn vin 4.46e-19
C205 ctl_3_ ctl_7_ 2.76e-20
C206 carray_0.unitcap_15.cn vin 4.46e-19
C207 sw_top_1.en_buf sw_top_1.net1 0.636f
C208 carray_0.unitcap_87.cn out 0.51f
C209 dum vdd 0.263f
C210 sky130_fd_sc_hd__inv_2_0.A ctl_5_ 0.00136f
C211 sw_top_1.en_buf vin 0.525f
C212 sky130_fd_sc_hd__inv_2_6.A ctl_2_ 0.103f
C213 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_9.cn 0.0902f
C214 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_7.cn 0.18f
C215 sky130_fd_sc_hd__inv_2_4.A ctl_1_ 1.37e-20
C216 sky130_fd_sc_hd__inv_2_8.A carray_0.unitcap_324.cn 0.14f
C217 carray_0.unitcap_88.cn carray_0.unitcap_104.cn 0.0902f
C218 carray_0.unitcap_326.cn vdd 0.00391f
C219 carray_0.unitcap_334.cn carray_0.unitcap_326.cn 0.18f
C220 carray_0.unitcap_127.cn carray_0.unitcap_119.cn 0.0902f
C221 ctl_5_ ctl_7_ 3.49e-19
C222 carray_0.unitcap_200.cn out 0.514f
C223 carray_0.unitcap_324.cn out 0.505f
C224 sky130_fd_sc_hd__inv_2_7.A carray_0.unitcap_248.cn 0.18f
C225 ctl_2_ ctl_4_ 2.49e-19
C226 carray_0.unitcap_9.cn sample 0.00536f
C227 sw_top_3.en_buf sw_top_2.net1 0.00175f
C228 carray_0.unitcap_167.cn carray_0.unitcap_183.cn 0.0902f
C229 sky130_fd_sc_hd__inv_2_9.A ctl_1_ 6.34e-22
C230 carray_0.unitcap_12.cn vin 0.0175f
C231 sw_top_1.en_buf sky130_fd_sc_hd__inv_2_9.A 0.604f
C232 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_255.cn 0.161f
C233 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_331.cn 0.0108f
C234 carray_0.unitcap_337.cn carray_0.unitcap_330.cn 0.18f
C235 carray_0.unitcap_72.cn out 0.514f
C236 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_191.cn 0.161f
C237 sky130_fd_sc_hd__inv_2_2.A carray_0.unitcap_321.cn 0.18f
C238 sky130_fd_sc_hd__inv_2_6.A ctl_4_ 0.0028f
C239 sw_top_1.en_buf sample 0.443f
C240 carray_0.unitcap_63.cn out 0.537f
C241 sky130_fd_sc_hd__inv_2_4.A sky130_fd_sc_hd__inv_2_2.VPB 0.0799f
C242 vdd ctl_1_ 0.269f
C243 carray_0.unitcap_12.cn sky130_fd_sc_hd__inv_2_9.A 0.0902f
C244 sw_top_1.en_buf vdd 1.84f
C245 vdd carray_0.unitcap_255.cn 0.00397f
C246 carray_0.unitcap_255.cn carray_0.unitcap_338.cn 0.0902f
C247 carray_0.unitcap_135.cn out 0.51f
C248 carray_0.unitcap_191.cn vdd 0.00397f
C249 sky130_fd_sc_hd__inv_2_2.A ctl_0_ 0.00127f
C250 carray_0.unitcap_56.cn carray_0.unitcap_48.cn 0.0902f
C251 carray_0.unitcap_112.cn out 0.514f
C252 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_88.cn 0.18f
C253 sky130_fd_sc_hd__inv_2_8.A ctl_2_ 3.25e-19
C254 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_127.cn 0.18f
C255 sky130_fd_sc_hd__inv_2_9.A sky130_fd_sc_hd__inv_2_2.VPB 0.079f
C256 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_167.cn 0.161f
C257 carray_0.unitcap_191.cn carray_0.unitcap_215.cn 0.0902f
C258 carray_0.unitcap_47.cn carray_0.unitcap_7.cn 0.0902f
C259 carray_0.unitcap_337.cn carray_0.unitcap_336.cn 0.18f
C260 ctl_2_ out 0.00201f
C261 sky130_fd_sc_hd__inv_2_4.A ctl_6_ 2.58e-20
C262 carray_0.unitcap_88.cn sample 6.36e-21
C263 carray_0.unitcap_23.cn out 0.512f
C264 sky130_fd_sc_hd__inv_2_6.A sky130_fd_sc_hd__inv_2_8.A 0.00332f
C265 carray_0.unitcap_104.cn carray_0.unitcap_96.cn 0.0902f
C266 carray_0.unitcap_328.cn vdd 0.00361f
C267 carray_0.unitcap_10.cn carray_0.unitcap_288.cn 0.18f
C268 carray_0.unitcap_127.cn vdd 0.00397f
C269 sky130_fd_sc_hd__inv_2_2.VPB vdd 0.432f
C270 sky130_fd_sc_hd__inv_2_2.VPB carray_0.unitcap_334.cn 0.00136f
C271 carray_0.unitcap_247.cn out 0.51f
C272 vdd carray_0.unitcap_167.cn 0.00397f
C273 sw_top_2.en_buf sw_top_2.net1 0.636f
C274 sky130_fd_sc_hd__inv_2_6.A out 2.01f
C275 carray_0.unitcap_207.cn carray_0.unitcap_191.cn 0.0902f
C276 sky130_fd_sc_hd__inv_2_9.A ctl_6_ 0.00149f
C277 sky130_fd_sc_hd__inv_2_8.A ctl_4_ 8.05e-20
C278 out sw_top_0.en_buf 0.709f
C279 carray_0.unitcap_320.cn out 0.496f
C280 carray_0.unitcap_64.cn out 0.514f
C281 carray_0.unitcap_12.cn carray_0.unitcap_13.cn 0.18f
C282 carray_0.unitcap_55.cn carray_0.unitcap_79.cn 0.0902f
C283 ctl_4_ out 0.00223f
C284 carray_0.unitcap_24.cn out 0.514f
C285 carray_0.unitcap_11.cn vin 0.0099f
C286 vdd ctl_6_ 0.271f
C287 sky130_fd_sc_hd__inv_2_6.A sky130_fd_sc_hd__inv_2_5.A 0.0927f
C288 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_48.cn 0.18f
C289 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_159.cn 0.18f
C290 sky130_fd_sc_hd__inv_2_4.A sky130_fd_sc_hd__inv_2_7.A 1.2f
C291 sky130_fd_sc_hd__inv_2_0.A ctl_0_ 6.35e-22
C292 carray_0.unitcap_160.cn carray_0.unitcap_176.cn 0.0902f
C293 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_96.cn 0.18f
C294 sky130_fd_sc_hd__inv_2_5.A ctl_4_ 0.00134f
C295 sky130_fd_sc_hd__inv_2_4.A sky130_fd_sc_hd__inv_2_3.A 1.71e-19
C296 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_11.cn 0.0902f
C297 carray_0.unitcap_48.cn sample 0.00149f
C298 sky130_fd_sc_hd__inv_2_9.A sky130_fd_sc_hd__inv_2_7.A 0.134f
C299 ctl_2_ dum 2.37e-19
C300 carray_0.unitcap_24.cn carray_0.unitcap_16.cn 0.0902f
C301 vdd carray_0.unitcap_48.cn 1.74e-19
C302 carray_0.unitcap_11.cn sample 0.00139f
C303 carray_0.unitcap_192.cn carray_0.unitcap_168.cn 0.0902f
C304 sky130_fd_sc_hd__inv_2_8.A out 0.54f
C305 sky130_fd_sc_hd__inv_2_4.A ctl_3_ 0.00142f
C306 ctl_2_ carray_0.unitcap_326.cn 0.00254f
C307 carray_0.unitcap_11.cn vdd 6.16e-19
C308 sky130_fd_sc_hd__inv_2_6.A dum 4.66e-19
C309 sw_top_0.net1 sw_top_1.net1 0.00267f
C310 carray_0.unitcap_175.cn carray_0.unitcap_199.cn 0.0902f
C311 sw_top_3.net1 out 0.373f
C312 sky130_fd_sc_hd__inv_2_7.A carray_0.unitcap_334.cn 0.0522f
C313 sky130_fd_sc_hd__inv_2_7.A vdd 0.146f
C314 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_330.cn 0.00328f
C315 sw_top_0.net1 vin 0.377f
C316 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_199.cn 0.161f
C317 sky130_fd_sc_hd__inv_2_6.A carray_0.unitcap_326.cn 0.361f
C318 sky130_fd_sc_hd__inv_2_9.A ctl_3_ 4.43e-21
C319 sky130_fd_sc_hd__inv_2_5.A sky130_fd_sc_hd__inv_2_8.A 1.1e-19
C320 sky130_fd_sc_hd__inv_2_3.A carray_0.unitcap_334.cn 2.28e-19
C321 carray_0.unitcap_79.cn vin 4.46e-19
C322 sky130_fd_sc_hd__inv_2_3.A vdd 0.104f
C323 carray_0.unitcap_40.cn out 0.514f
C324 carray_0.unitcap_15.cn carray_0.unitcap_23.cn 0.0902f
C325 carray_0.unitcap_136.cn carray_0.unitcap_128.cn 0.0902f
C326 carray_0.unitcap_321.cn carray_0.unitcap_248.cn 0.0902f
C327 carray_0.unitcap_10.cn vin 0.0025f
C328 out carray_0.unitcap_95.cn 0.51f
C329 sky130_fd_sc_hd__inv_2_4.A ctl_5_ 0.0154f
C330 sky130_fd_sc_hd__inv_2_5.A out 17.5f
C331 ctl_2_ ctl_1_ 0.0686f
C332 carray_0.unitcap_11.cn carray_0.unitcap_13.cn 0.18f
C333 carray_0.unitcap_256.cn out 0.557f
C334 carray_0.unitcap_330.cn vdd 0.058f
C335 sw_top_0.net1 sky130_fd_sc_hd__inv_2_9.A 0.44f
C336 sky130_fd_sc_hd__inv_2_2.A carray_0.unitcap_322.cn 0.00173f
C337 carray_0.unitcap_176.cn carray_0.unitcap_168.cn 0.0902f
C338 carray_0.unitcap_199.cn vdd 0.00397f
C339 carray_0.unitcap_32.cn out 0.514f
C340 ctl_3_ carray_0.unitcap_334.cn 0.00225f
C341 ctl_3_ vdd 0.269f
C342 carray_0.unitcap_16.cn out 0.515f
C343 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_79.cn 0.18f
C344 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_10.cn 0.0902f
C345 sky130_fd_sc_hd__inv_2_9.A ctl_5_ 1.3e-20
C346 sky130_fd_sc_hd__inv_2_6.A ctl_1_ 0.0234f
C347 sw_top_0.net1 sample 0.0138f
C348 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_336.cn 0.161f
C349 sw_top_3.en_buf vin 0.53f
C350 carray_0.unitcap_143.cn carray_0.unitcap_119.cn 0.0902f
C351 carray_0.unitcap_40.cn carray_0.unitcap_32.cn 0.0902f
C352 carray_0.unitcap_159.cn carray_0.unitcap_151.cn 0.0902f
C353 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_231.cn 0.161f
C354 sw_top_0.net1 vdd 0.819f
C355 sw_top_1.en_buf sw_top_0.en_buf 0.00273f
C356 carray_0.unitcap_192.cn carray_0.unitcap_200.cn 0.0902f
C357 sky130_fd_sc_hd__inv_2_4.A carray_0.unitcap_331.cn 0.0404f
C358 sky130_fd_sc_hd__inv_2_8.A dum 0.057f
C359 carray_0.unitcap_10.cn sample 0.00512f
C360 ctl_4_ ctl_1_ 8.03e-21
C361 carray_0.unitcap_39.cn vin 4.46e-19
C362 carray_0.unitcap_10.cn vdd 7.04e-19
C363 ctl_5_ vdd 0.269f
C364 sky130_fd_sc_hd__inv_2_2.VPB ctl_2_ 0.0102f
C365 sw_top_3.en_buf sky130_fd_sc_hd__inv_2_9.A 0.747f
C366 vdd carray_0.unitcap_336.cn 0.00397f
C367 dum out 0.0018f
C368 carray_0.unitcap_14.cn out 0.556f
C369 carray_0.unitcap_338.cn carray_0.unitcap_336.cn 0.0902f
C370 carray_0.unitcap_199.cn carray_0.unitcap_207.cn 0.0902f
C371 carray_0.unitcap_231.cn vdd 0.00397f
C372 sw_top_2.en_buf carray_0.unitcap_56.cn 3.18e-20
C373 sky130_fd_sc_hd__inv_2_6.A carray_0.unitcap_328.cn 0.113f
C374 carray_0.unitcap_232.cn out 0.514f
C375 sky130_fd_sc_hd__inv_2_0.A ctl_7_ 0.0296f
C376 carray_0.unitcap_72.cn carray_0.unitcap_48.cn 0.0902f
C377 carray_0.unitcap_326.cn out 0.501f
C378 sw_top_3.en_buf sample 0.443f
C379 sky130_fd_sc_hd__inv_2_6.A sky130_fd_sc_hd__inv_2_2.VPB 0.0806f
C380 carray_0.unitcap_215.cn carray_0.unitcap_231.cn 0.0902f
C381 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_39.cn 0.18f
C382 carray_0.unitcap_208.cn out 0.514f
C383 carray_0.unitcap_88.cn sw_top_0.en_buf 6.36e-20
C384 sw_top_3.en_buf vdd 1.84f
C385 carray_0.unitcap_88.cn carray_0.unitcap_64.cn 0.0902f
C386 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_143.cn 0.18f
C387 carray_0.unitcap_9.cn out 0.557f
C388 carray_0.unitcap_334.cn carray_0.unitcap_331.cn 0.18f
C389 carray_0.unitcap_331.cn vdd 0.00379f
C390 carray_0.unitcap_7.cn out 0.51f
C391 sky130_fd_sc_hd__inv_2_2.VPB ctl_4_ 0.01f
C392 carray_0.unitcap_15.cn out 0.501f
C393 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_120.cn 0.18f
C394 sky130_fd_sc_hd__inv_2_8.A ctl_1_ 0.00217f
C395 sw_top_2.en_buf sw_top_1.net1 0.00175f
C396 carray_0.unitcap_208.cn sky130_fd_sc_hd__inv_2_5.A 0.18f
C397 sw_top_2.en_buf vin 0.526f
C398 ctl_1_ out 0.00224f
C399 sky130_fd_sc_hd__inv_2_6.A ctl_6_ 1.24e-21
C400 sw_top_1.en_buf out 0.747f
C401 carray_0.unitcap_143.cn vdd 0.00397f
C402 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_128.cn 0.18f
C403 carray_0.unitcap_255.cn out 0.51f
C404 carray_0.unitcap_152.cn out 0.514f
C405 carray_0.unitcap_256.cn carray_0.unitcap_9.cn 0.18f
C406 carray_0.unitcap_79.cn carray_0.unitcap_87.cn 0.0902f
C407 carray_0.unitcap_191.cn out 0.51f
C408 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_223.cn 0.161f
C409 ctl_4_ ctl_6_ 1.99e-19
C410 sw_top_2.en_buf sky130_fd_sc_hd__inv_2_9.A 0.837f
C411 carray_0.unitcap_337.cn sky130_fd_sc_hd__inv_2_0.A 0.13f
C412 sky130_fd_sc_hd__inv_2_8.A carray_0.unitcap_328.cn 0.00461f
C413 carray_0.unitcap_12.cn out 0.556f
C414 sky130_fd_sc_hd__inv_2_5.A ctl_1_ 3.45e-21
C415 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_80.cn 0.18f
C416 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_sc_hd__inv_2_8.A 0.0821f
C417 sky130_fd_sc_hd__inv_2_7.A ctl_2_ 0.00404f
C418 sky130_fd_sc_hd__inv_2_4.A ctl_0_ 5.4e-21
C419 vdd carray_0.unitcap_223.cn 0.00397f
C420 carray_0.unitcap_47.cn carray_0.unitcap_39.cn 0.0902f
C421 sky130_fd_sc_hd__inv_2_5.A carray_0.unitcap_191.cn 0.18f
C422 carray_0.unitcap_328.cn out 0.501f
C423 sw_top_2.en_buf sample 0.443f
C424 carray_0.unitcap_88.cn out 0.514f
C425 sky130_fd_sc_hd__inv_2_4.A carray_0.unitcap_240.cn 0.18f
C426 carray_0.unitcap_127.cn out 0.51f
C427 sky130_fd_sc_hd__inv_2_2.VPB out 0.00887f
C428 carray_0.unitcap_216.cn out 0.514f
C429 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_151.cn 0.18f
C430 carray_0.unitcap_80.cn sample 0.00149f
C431 sky130_fd_sc_hd__inv_2_3.A ctl_2_ 0.00141f
C432 out carray_0.unitcap_167.cn 0.51f
C433 sw_top_2.en_buf vdd 1.84f
C434 sky130_fd_sc_hd__inv_2_6.A sky130_fd_sc_hd__inv_2_7.A 0.613f
C435 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_159.cn 0.161f
C436 carray_0.unitcap_80.cn vdd 6.25e-20
C437 carray_0.unitcap_14.cn carray_0.unitcap_15.cn 0.18f
C438 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_136.cn 0.18f
C439 sky130_fd_sc_hd__inv_2_6.A sky130_fd_sc_hd__inv_2_3.A 0.39f
C440 carray_0.unitcap_103.cn carray_0.unitcap_111.cn 0.0902f
C441 sky130_fd_sc_hd__inv_2_7.A ctl_4_ 0.0154f
C442 sky130_fd_sc_hd__inv_2_4.A carray_0.unitcap_239.cn 0.18f
C443 ctl_3_ ctl_2_ 0.0744f
C444 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_sc_hd__inv_2_5.A 0.081f
C445 carray_0.unitcap_216.cn sky130_fd_sc_hd__inv_2_5.A 0.18f
C446 dum ctl_1_ 3.73e-19
C447 out ctl_6_ 0.00223f
C448 carray_0.unitcap_159.cn vdd 0.00397f
C449 sky130_fd_sc_hd__inv_2_6.A carray_0.unitcap_330.cn 0.0919f
C450 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_144.cn 0.18f
C451 sky130_fd_sc_hd__inv_2_4.A sky130_fd_sc_hd__inv_2_2.A 2.49e-21
C452 ctl_0_ vdd 0.269f
C453 sky130_fd_sc_hd__inv_2_3.A ctl_4_ 6.53e-21
C454 sky130_fd_sc_hd__inv_2_6.A ctl_3_ 0.00386f
C455 carray_0.unitcap_326.cn ctl_1_ 0.00226f
C456 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_239.cn 0.161f
C457 carray_0.unitcap_192.cn out 0.514f
C458 carray_0.unitcap_14.cn carray_0.unitcap_12.cn 0.18f
C459 ctl_3_ ctl_4_ 0.0695f
C460 ctl_2_ ctl_5_ 2.63e-21
C461 sky130_fd_sc_hd__inv_2_5.A ctl_6_ 0.0228f
C462 carray_0.unitcap_48.cn out 0.514f
C463 carray_0.unitcap_328.cn dum 0.00171f
C464 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_0.cn 0.18f
C465 sw_top_0.net1 sw_top_0.en_buf 0.636f
C466 carray_0.unitcap_39.cn carray_0.unitcap_63.cn 0.0902f
C467 vdd carray_0.unitcap_239.cn 0.00397f
C468 sky130_fd_sc_hd__inv_2_2.VPB dum 0.0104f
C469 carray_0.unitcap_96.cn out 0.514f
C470 sky130_fd_sc_hd__inv_2_7.A sky130_fd_sc_hd__inv_2_8.A 0.094f
C471 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_71.cn 0.18f
C472 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_183.cn 0.18f
C473 sky130_fd_sc_hd__inv_2_6.A ctl_5_ 4.49e-21
C474 carray_0.unitcap_11.cn out 0.556f
C475 sky130_fd_sc_hd__inv_2_2.A vdd 0.0829f
C476 carray_0.unitcap_200.cn carray_0.unitcap_184.cn 0.0902f
C477 carray_0.unitcap_326.cn carray_0.unitcap_328.cn 0.18f
C478 sky130_fd_sc_hd__inv_2_7.A out 4.37f
C479 sw_top_1.net1 sw_top_2.net1 0.00267f
C480 sky130_fd_sc_hd__inv_2_3.A sky130_fd_sc_hd__inv_2_8.A 0.409f
C481 carray_0.unitcap_0.cn sample 0.00152f
C482 sky130_fd_sc_hd__inv_2_2.VPB carray_0.unitcap_326.cn 0.00172f
C483 carray_0.unitcap_0.cn vdd 1.03e-19
C484 ctl_5_ ctl_4_ 0.0684f
C485 carray_0.unitcap_143.cn carray_0.unitcap_135.cn 0.0902f
C486 sw_top_2.net1 vin 0.392f
C487 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_160.cn 0.18f
C488 out carray_0.unitcap_176.cn 0.514f
C489 sky130_fd_sc_hd__inv_2_3.A out 1.03f
C490 sky130_fd_sc_hd__inv_2_4.A sky130_fd_sc_hd__inv_2_0.A 0.663f
C491 sky130_fd_sc_hd__inv_2_8.A ctl_3_ 1.53e-19
C492 carray_0.unitcap_120.cn carray_0.unitcap_112.cn 0.0902f
C493 sample carray_0.unitcap_8.cn 0.00149f
C494 sky130_fd_sc_hd__inv_2_6.A carray_0.unitcap_331.cn 0.135f
C495 sky130_fd_sc_hd__inv_2_5.A sky130_fd_sc_hd__inv_2_7.A 0.0883f
C496 carray_0.unitcap_330.cn out 0.502f
C497 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_175.cn 0.18f
C498 carray_0.unitcap_199.cn out 0.51f
C499 ctl_3_ out 0.00214f
C500 carray_0.unitcap_72.cn carray_0.unitcap_80.cn 0.0902f
C501 sky130_fd_sc_hd__inv_2_9.A sw_top_2.net1 0.358f
C502 sky130_fd_sc_hd__inv_2_4.A ctl_7_ 4.24e-20
C503 sky130_fd_sc_hd__inv_2_2.VPB ctl_1_ 0.01f
C504 sky130_fd_sc_hd__inv_2_5.A sky130_fd_sc_hd__inv_2_3.A 1.23e-20
C505 sky130_fd_sc_hd__inv_2_0.A sky130_fd_sc_hd__inv_2_9.A 3.29f
C506 carray_0.unitcap_31.cn vin 4.46e-19
C507 sw_top_2.net1 sample 0.0344f
C508 sky130_fd_sc_hd__inv_2_5.A carray_0.unitcap_330.cn 0.0288f
C509 sw_top_0.net1 out 0.383f
C510 sky130_fd_sc_hd__inv_2_8.A ctl_5_ 5.26e-20
C511 sky130_fd_sc_hd__inv_2_9.A ctl_7_ 0.0967f
C512 sw_top_2.net1 vdd 0.824f
C513 carray_0.unitcap_79.cn out 0.51f
C514 sky130_fd_sc_hd__inv_2_5.A ctl_3_ 3.08e-20
C515 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_111.cn 0.18f
C516 sky130_fd_sc_hd__inv_2_0.A vdd 1f
C517 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_334.cn 0.00107f
C518 carray_0.unitcap_10.cn out 0.557f
C519 ctl_5_ out 0.00193f
C520 carray_0.unitcap_336.cn out 0.496f
C521 sky130_fd_sc_hd__inv_2_7.A dum 8.18e-21
C522 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_31.cn 0.18f
C523 ctl_1_ ctl_6_ 1.88e-21
C524 carray_0.unitcap_231.cn out 0.51f
C525 carray_0.unitcap_223.cn carray_0.unitcap_247.cn 0.0902f
C526 sky130_fd_sc_hd__inv_2_2.VPB carray_0.unitcap_328.cn 0.00245f
C527 vdd ctl_7_ 0.282f
C528 carray_0.unitcap_87.cn carray_0.unitcap_71.cn 0.0902f
C529 carray_0.unitcap_135.cn carray_0.unitcap_159.cn 0.0902f
C530 sky130_fd_sc_hd__inv_2_3.A dum 0.0261f
C531 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_168.cn 0.18f
C532 sky130_fd_sc_hd__inv_2_7.A carray_0.unitcap_326.cn 0.0361f
C533 sky130_fd_sc_hd__inv_2_2.A carray_0.unitcap_324.cn 0.291f
C534 sw_top_3.en_buf sw_top_3.net1 0.636f
C535 sw_top_3.en_buf out 0.453f
C536 sky130_fd_sc_hd__inv_2_5.A ctl_5_ 0.1f
C537 carray_0.unitcap_112.cn carray_0.unitcap_136.cn 0.0902f
C538 sky130_fd_sc_hd__inv_2_3.A carray_0.unitcap_326.cn 0.0955f
C539 carray_0.unitcap_331.cn out 0.501f
C540 sky130_fd_sc_hd__inv_2_5.A carray_0.unitcap_231.cn 0.18f
C541 ctl_2_ ctl_0_ 4.97e-20
C542 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_207.cn 0.18f
C543 ctl_3_ dum 1.05e-20
C544 carray_0.unitcap_321.cn carray_0.unitcap_320.cn 0.0902f
C545 sw_top_3.en_buf carray_0.unitcap_40.cn 6.36e-20
C546 carray_0.unitcap_80.cn carray_0.unitcap_64.cn 0.0902f
C547 carray_0.unitcap_39.cn out 0.537f
C548 sky130_fd_sc_hd__inv_2_2.VPB ctl_6_ 0.0105f
C549 carray_0.unitcap_337.cn sky130_fd_sc_hd__inv_2_9.A 0.14f
C550 sky130_fd_sc_hd__inv_2_7.A ctl_1_ 5.41e-20
C551 carray_0.unitcap_143.cn out 0.51f
C552 sky130_fd_sc_hd__inv_2_6.A ctl_0_ 0.00134f
C553 sky130_fd_sc_hd__inv_2_7.A carray_0.unitcap_255.cn 0.18f
C554 sky130_fd_sc_hd__inv_2_5.A carray_0.unitcap_331.cn 0.0597f
C555 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_288.cn 0.0902f
C556 carray_0.unitcap_120.cn out 0.514f
C557 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_103.cn 0.18f
C558 carray_0.unitcap_55.cn vin 4.46e-19
C559 sky130_fd_sc_hd__inv_2_3.A ctl_1_ 0.0996f
C560 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_151.cn 0.161f
C561 carray_0.unitcap_144.cn carray_0.unitcap_160.cn 0.0902f
C562 ctl_4_ ctl_0_ 2.97e-21
C563 carray_0.unitcap_337.cn vdd 0.0135f
C564 carray_0.unitcap_288.cn sample 0.0938f
C565 sky130_fd_sc_hd__inv_2_2.A ctl_2_ 1.07e-20
C566 carray_0.unitcap_247.cn carray_0.unitcap_239.cn 0.0902f
C567 carray_0.unitcap_288.cn vdd 2.22e-20
C568 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_200.cn 0.18f
C569 carray_0.unitcap_184.cn out 0.514f
C570 carray_0.unitcap_103.cn vdd 0.00397f
C571 ctl_3_ ctl_1_ 5.59e-20
C572 carray_0.unitcap_223.cn out 0.51f
C573 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_55.cn 0.18f
C574 sky130_fd_sc_hd__inv_2_7.A carray_0.unitcap_328.cn 0.007f
C575 vdd carray_0.unitcap_151.cn 0.00397f
C576 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_sc_hd__inv_2_7.A 0.0798f
C577 sky130_fd_sc_hd__inv_2_6.A sky130_fd_sc_hd__inv_2_2.A 4.85e-19
C578 sw_top_2.en_buf sw_top_3.net1 2.34e-19
C579 sw_top_2.en_buf out 0.712f
C580 carray_0.unitcap_321.cn out 0.512f
C581 sky130_fd_sc_hd__inv_2_3.A carray_0.unitcap_328.cn 0.323f
C582 carray_0.unitcap_80.cn out 0.514f
C583 sky130_fd_sc_hd__inv_2_2.A carray_0.unitcap_320.cn 0.109f
C584 sw_top_0.net1 sw_top_1.en_buf 0.00175f
C585 sky130_fd_sc_hd__inv_2_2.VPB sky130_fd_sc_hd__inv_2_3.A 0.0867f
C586 sky130_fd_sc_hd__inv_2_5.A carray_0.unitcap_184.cn 0.18f
C587 sky130_fd_sc_hd__inv_2_5.A carray_0.unitcap_223.cn 0.18f
C588 sky130_fd_sc_hd__inv_2_8.A ctl_0_ 0.108f
C589 carray_0.unitcap_322.cn carray_0.unitcap_324.cn 0.18f
C590 ctl_5_ ctl_1_ 4.37e-20
C591 sky130_fd_sc_hd__inv_2_2.VPB carray_0.unitcap_330.cn 0.00125f
C592 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_56.cn 0.18f
C593 sky130_fd_sc_hd__inv_2_0.A carray_0.unitcap_135.cn 0.18f
C594 carray_0.unitcap_24.cn carray_0.unitcap_0.cn 0.0902f
C595 carray_0.unitcap_159.cn out 0.51f
C596 sky130_fd_sc_hd__inv_2_7.A ctl_6_ 1.56e-20
C597 ctl_0_ out 0.00178f
C598 sw_top_1.net1 vin 0.392f
C599 sky130_fd_sc_hd__inv_2_2.VPB ctl_3_ 0.0103f
C600 carray_0.unitcap_175.cn carray_0.unitcap_183.cn 0.0902f
C601 carray_0.unitcap_136.cn out 0.514f
C602 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_104.cn 0.18f
C603 carray_0.unitcap_240.cn out 0.514f
C604 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_119.cn 0.18f
C605 carray_0.unitcap_56.cn sample 0.00152f
C606 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_183.cn 0.161f
C607 sky130_fd_sc_hd__inv_2_3.A ctl_6_ 1.64e-21
C608 sky130_fd_sc_hd__inv_2_9.A sw_top_1.net1 0.485f
C609 sky130_fd_sc_hd__inv_2_5.A ctl_0_ 1.74e-21
C610 carray_0.unitcap_119.cn vdd 0.00397f
C611 sky130_fd_sc_hd__inv_2_2.A sky130_fd_sc_hd__inv_2_8.A 0.723f
C612 carray_0.unitcap_239.cn out 0.51f
C613 ctl_2_ ctl_7_ 1.59e-20
C614 ctl_3_ ctl_6_ 2.37e-19
C615 vdd carray_0.unitcap_183.cn 0.00397f
C616 sky130_fd_sc_hd__inv_2_2.VPB ctl_5_ 0.0101f
C617 sky130_fd_sc_hd__inv_2_9.A vin 4.52f
C618 sky130_fd_sc_hd__inv_2_6.A sky130_fd_sc_hd__inv_2_0.A 0.359f
C619 sky130_fd_sc_hd__inv_2_4.A sky130_fd_sc_hd__inv_2_9.A 0.29f
C620 sw_top_1.net1 sample 0.0344f
C621 sky130_fd_sc_hd__inv_2_2.A out 0.544f
C622 carray_0.unitcap_208.cn carray_0.unitcap_184.cn 0.0902f
C623 sw_top_1.net1 vdd 0.824f
C624 sky130_fd_sc_hd__inv_2_9.A carray_0.unitcap_175.cn 0.161f
C625 dum vss 0.235f
C626 ctl_0_ vss 0.194f
C627 sample vss 5.86f
C628 ctl_1_ vss 0.194f
C629 ctl_2_ vss 0.198f
C630 ctl_3_ vss 0.196f
C631 ctl_4_ vss 0.196f
C632 ctl_5_ vss 0.199f
C633 out vss 54.2f
C634 vin vss 4.85f
C635 ctl_6_ vss 0.197f
C636 ctl_7_ vss 0.242f
C637 vdd vss 46.4f
C638 carray_0.unitcap_320.cn vss 0.28f
C639 carray_0.unitcap_321.cn vss 0.206f
C640 carray_0.unitcap_248.cn vss 0.204f
C641 carray_0.unitcap_232.cn vss 0.204f
C642 carray_0.unitcap_240.cn vss 0.204f
C643 carray_0.unitcap_216.cn vss 0.204f
C644 carray_0.unitcap_224.cn vss 0.204f
C645 carray_0.unitcap_208.cn vss 0.204f
C646 carray_0.unitcap_184.cn vss 0.204f
C647 carray_0.unitcap_200.cn vss 0.204f
C648 carray_0.unitcap_192.cn vss 0.204f
C649 carray_0.unitcap_168.cn vss 0.204f
C650 carray_0.unitcap_176.cn vss 0.204f
C651 carray_0.unitcap_160.cn vss 0.204f
C652 carray_0.unitcap_144.cn vss 0.204f
C653 carray_0.unitcap_152.cn vss 0.204f
C654 carray_0.unitcap_128.cn vss 0.204f
C655 carray_0.unitcap_136.cn vss 0.204f
C656 carray_0.unitcap_112.cn vss 0.204f
C657 carray_0.unitcap_120.cn vss 0.204f
C658 carray_0.unitcap_96.cn vss 0.204f
C659 carray_0.unitcap_104.cn vss 0.204f
C660 carray_0.unitcap_88.cn vss 0.202f
C661 carray_0.unitcap_64.cn vss 0.202f
C662 carray_0.unitcap_80.cn vss 0.202f
C663 carray_0.unitcap_72.cn vss 0.202f
C664 carray_0.unitcap_48.cn vss 0.202f
C665 carray_0.unitcap_56.cn vss 0.202f
C666 carray_0.unitcap_32.cn vss 0.202f
C667 carray_0.unitcap_40.cn vss 0.202f
C668 carray_0.unitcap_0.cn vss 0.202f
C669 carray_0.unitcap_24.cn vss 0.202f
C670 carray_0.unitcap_16.cn vss 0.201f
C671 carray_0.unitcap_8.cn vss 0.271f
C672 carray_0.unitcap_324.cn vss 0.192f
C673 carray_0.unitcap_9.cn vss 0.189f
C674 carray_0.unitcap_322.cn vss 0.223f
C675 carray_0.unitcap_256.cn vss 0.186f
C676 carray_0.unitcap_328.cn vss 0.195f
C677 carray_0.unitcap_288.cn vss 0.187f
C678 carray_0.unitcap_326.cn vss 0.168f
C679 carray_0.unitcap_10.cn vss 0.189f
C680 carray_0.unitcap_334.cn vss 0.16f
C681 carray_0.unitcap_11.cn vss 0.189f
C682 carray_0.unitcap_331.cn vss 0.177f
C683 carray_0.unitcap_13.cn vss 0.182f
C684 carray_0.unitcap_330.cn vss 0.167f
C685 carray_0.unitcap_12.cn vss 0.189f
C686 carray_0.unitcap_337.cn vss 0.176f
C687 carray_0.unitcap_14.cn vss 0.189f
C688 carray_0.unitcap_336.cn vss 0.265f
C689 carray_0.unitcap_338.cn vss 0.196f
C690 carray_0.unitcap_255.cn vss 0.196f
C691 carray_0.unitcap_239.cn vss 0.196f
C692 carray_0.unitcap_247.cn vss 0.196f
C693 carray_0.unitcap_223.cn vss 0.196f
C694 carray_0.unitcap_231.cn vss 0.196f
C695 carray_0.unitcap_215.cn vss 0.196f
C696 carray_0.unitcap_191.cn vss 0.196f
C697 carray_0.unitcap_207.cn vss 0.196f
C698 carray_0.unitcap_199.cn vss 0.196f
C699 carray_0.unitcap_175.cn vss 0.196f
C700 carray_0.unitcap_183.cn vss 0.196f
C701 carray_0.unitcap_167.cn vss 0.196f
C702 carray_0.unitcap_151.cn vss 0.196f
C703 carray_0.unitcap_159.cn vss 0.196f
C704 carray_0.unitcap_135.cn vss 0.196f
C705 carray_0.unitcap_143.cn vss 0.201f
C706 carray_0.unitcap_119.cn vss 0.201f
C707 carray_0.unitcap_127.cn vss 0.201f
C708 carray_0.unitcap_103.cn vss 0.201f
C709 carray_0.unitcap_111.cn vss 0.201f
C710 carray_0.unitcap_95.cn vss 0.201f
C711 carray_0.unitcap_71.cn vss 0.201f
C712 carray_0.unitcap_87.cn vss 0.201f
C713 carray_0.unitcap_79.cn vss 0.201f
C714 carray_0.unitcap_55.cn vss 0.201f
C715 carray_0.unitcap_63.cn vss 0.199f
C716 carray_0.unitcap_39.cn vss 0.199f
C717 carray_0.unitcap_47.cn vss 0.201f
C718 carray_0.unitcap_7.cn vss 0.201f
C719 carray_0.unitcap_31.cn vss 0.201f
C720 carray_0.unitcap_23.cn vss 0.201f
C721 carray_0.unitcap_15.cn vss 0.271f
C722 sky130_fd_sc_hd__inv_2_2.A vss 1.5f
C723 sky130_fd_sc_hd__inv_2_8.A vss 1.5f
C724 sky130_fd_sc_hd__inv_2_3.A vss 1.37f
C725 sky130_fd_sc_hd__inv_2_6.A vss 1.6f
C726 sw_top_0.net1 vss 1.97f
C727 sky130_fd_sc_hd__inv_2_7.A vss 2.49f
C728 sw_top_1.net1 vss 1.94f
C729 sw_top_2.net1 vss 1.94f
C730 sw_top_3.net1 vss 1.94f
C731 sky130_fd_sc_hd__inv_2_4.A vss 3.91f
C732 sky130_fd_sc_hd__inv_2_5.A vss 25.3f
C733 sw_top_0.en_buf vss 1.59f
C734 sw_top_1.en_buf vss 1.5f
C735 sw_top_2.en_buf vss 1.5f
C736 sw_top_3.en_buf vss 1.7f
C737 sky130_fd_sc_hd__inv_2_0.A vss 13.9f
C738 sky130_fd_sc_hd__inv_2_9.A vss 0.119p
C739 sky130_fd_sc_hd__inv_2_2.VPB vss 2.5f
C740 sky130_fd_sc_hd__inv_2_5.A.n0 vss 0.0012f
C741 sky130_fd_sc_hd__inv_2_5.A.t3 vss 0.00602f
C742 sky130_fd_sc_hd__inv_2_5.A.t1 vss 0.0102f
C743 sky130_fd_sc_hd__inv_2_5.A.t4 vss 0.00602f
C744 sky130_fd_sc_hd__inv_2_5.A.t2 vss 0.0102f
C745 sky130_fd_sc_hd__inv_2_5.A.n1 vss 0.0171f
C746 sky130_fd_sc_hd__inv_2_5.A.n2 vss 0.0176f
C747 sky130_fd_sc_hd__inv_2_5.A.n3 vss 0.00295f
C748 sky130_fd_sc_hd__inv_2_5.A.n4 vss 0.00621f
C749 sky130_fd_sc_hd__inv_2_5.A.n5 vss 0.0419f
C750 sky130_fd_sc_hd__inv_2_5.A.n6 vss 0.625f
C751 sky130_fd_sc_hd__inv_2_5.A.t0 vss 0.48f
C752 sample.n0 vss 0.00939f
C753 sample.n1 vss 0.00497f
C754 sample.n2 vss 0.00687f
C755 sample.n3 vss 0.0026f
C756 sample.t14 vss 0.0175f
C757 sample.t30 vss 0.0103f
C758 sample.t24 vss 0.0175f
C759 sample.t8 vss 0.0103f
C760 sample.n4 vss 0.0252f
C761 sample.t11 vss 0.0175f
C762 sample.t28 vss 0.0103f
C763 sample.t20 vss 0.0175f
C764 sample.t6 vss 0.0103f
C765 sample.n5 vss 0.0236f
C766 sample.n6 vss 0.0118f
C767 sample.n7 vss 0.0252f
C768 sample.n8 vss 0.0115f
C769 sample.n9 vss 0.00957f
C770 sample.n10 vss 0.00957f
C771 sample.n11 vss 0.0115f
C772 sample.n12 vss 0.0293f
C773 sample.n13 vss 0.015f
C774 sample.n14 vss 0.00198f
C775 sample.n15 vss 0.00476f
C776 sample.n16 vss 0.00206f
C777 sample.n17 vss 0.00208f
C778 sample.n18 vss 9.72e-19
C779 sample.n19 vss 0.0652f
C780 sample.n20 vss 0.00939f
C781 sample.n21 vss 0.00495f
C782 sample.n22 vss 0.00206f
C783 sample.n23 vss 0.00689f
C784 sample.n24 vss 0.00476f
C785 sample.n25 vss 0.0026f
C786 sample.t27 vss 0.0175f
C787 sample.t13 vss 0.0103f
C788 sample.t16 vss 0.0175f
C789 sample.t0 vss 0.0103f
C790 sample.n26 vss 0.0252f
C791 sample.t2 vss 0.0175f
C792 sample.t19 vss 0.0103f
C793 sample.t12 vss 0.0175f
C794 sample.t29 vss 0.0103f
C795 sample.n27 vss 0.0236f
C796 sample.n28 vss 0.0118f
C797 sample.n29 vss 0.0252f
C798 sample.n30 vss 0.0115f
C799 sample.n31 vss 0.00957f
C800 sample.n32 vss 0.00957f
C801 sample.n33 vss 0.0115f
C802 sample.n34 vss 0.0293f
C803 sample.n35 vss 0.015f
C804 sample.n36 vss 0.00198f
C805 sample.n37 vss 0.00208f
C806 sample.n38 vss 0.00151f
C807 sample.n39 vss 0.0611f
C808 sample.n40 vss 0.031f
C809 sample.n41 vss 0.00939f
C810 sample.n42 vss 0.00495f
C811 sample.n43 vss 0.00206f
C812 sample.n44 vss 0.00689f
C813 sample.n45 vss 0.00476f
C814 sample.n46 vss 0.0026f
C815 sample.t7 vss 0.0175f
C816 sample.t23 vss 0.0103f
C817 sample.t4 vss 0.0175f
C818 sample.t21 vss 0.0103f
C819 sample.n47 vss 0.0252f
C820 sample.t17 vss 0.0175f
C821 sample.t1 vss 0.0103f
C822 sample.t10 vss 0.0175f
C823 sample.t26 vss 0.0103f
C824 sample.n48 vss 0.0236f
C825 sample.n49 vss 0.0118f
C826 sample.n50 vss 0.0252f
C827 sample.n51 vss 0.0115f
C828 sample.n52 vss 0.00957f
C829 sample.n53 vss 0.00957f
C830 sample.n54 vss 0.0115f
C831 sample.n55 vss 0.0293f
C832 sample.n56 vss 0.015f
C833 sample.n57 vss 0.00198f
C834 sample.n58 vss 0.00208f
C835 sample.n59 vss 0.00151f
C836 sample.n60 vss 0.0618f
C837 sample.n61 vss 0.0303f
C838 sample.n62 vss 0.00939f
C839 sample.n63 vss 0.00495f
C840 sample.n64 vss 0.00206f
C841 sample.n65 vss 0.00689f
C842 sample.n66 vss 0.00476f
C843 sample.n67 vss 0.0026f
C844 sample.t5 vss 0.0175f
C845 sample.t22 vss 0.0103f
C846 sample.t18 vss 0.0175f
C847 sample.t3 vss 0.0103f
C848 sample.n68 vss 0.0252f
C849 sample.t15 vss 0.0175f
C850 sample.t31 vss 0.0103f
C851 sample.t25 vss 0.0175f
C852 sample.t9 vss 0.0103f
C853 sample.n69 vss 0.0236f
C854 sample.n70 vss 0.0118f
C855 sample.n71 vss 0.0252f
C856 sample.n72 vss 0.0115f
C857 sample.n73 vss 0.00957f
C858 sample.n74 vss 0.00957f
C859 sample.n75 vss 0.0115f
C860 sample.n76 vss 0.0293f
C861 sample.n77 vss 0.015f
C862 sample.n78 vss 0.00198f
C863 sample.n79 vss 0.00208f
C864 sample.n80 vss 0.00151f
C865 sample.n81 vss 0.0647f
C866 sample.n82 vss 0.347f
C867 sample.n83 vss 0.337f
C868 sample.n84 vss 0.416f
C869 sky130_fd_sc_hd__inv_2_9.A.t0 vss 0.35f
C870 sky130_fd_sc_hd__inv_2_9.A.t1 vss 0.46f
C871 sky130_fd_sc_hd__inv_2_9.A.n0 vss 0.212f
C872 sky130_fd_sc_hd__inv_2_9.A.t2 vss 0.00674f
C873 sky130_fd_sc_hd__inv_2_9.A.t5 vss 0.0114f
C874 sky130_fd_sc_hd__inv_2_9.A.t4 vss 0.00674f
C875 sky130_fd_sc_hd__inv_2_9.A.t3 vss 0.0114f
C876 sky130_fd_sc_hd__inv_2_9.A.n1 vss 0.0192f
C877 sky130_fd_sc_hd__inv_2_9.A.n2 vss 0.0223f
C878 sky130_fd_sc_hd__inv_2_9.A.n3 vss 0.111f
C879 vdd.t12 vss 0.00692f
C880 vdd.t147 vss 0.0115f
C881 vdd.t110 vss 0.00509f
C882 vdd.n0 vss 0.00954f
C883 vdd.n1 vss 0.0189f
C884 vdd.n2 vss 0.0151f
C885 vdd.t111 vss 0.00509f
C886 vdd.n3 vss 0.0108f
C887 vdd.t66 vss 0.00846f
C888 vdd.n4 vss 0.00907f
C889 vdd.t81 vss 0.00845f
C890 vdd.n5 vss 0.00964f
C891 vdd.t47 vss 0.00846f
C892 vdd.n6 vss 0.0104f
C893 vdd.t46 vss 0.00845f
C894 vdd.n7 vss 0.00964f
C895 vdd.t92 vss 0.00846f
C896 vdd.n8 vss 0.0104f
C897 vdd.t93 vss 0.00845f
C898 vdd.n9 vss 0.00964f
C899 vdd.t142 vss 0.00846f
C900 vdd.n10 vss 0.0104f
C901 vdd.t143 vss 0.00845f
C902 vdd.n11 vss 0.0096f
C903 vdd.t3 vss 0.00846f
C904 vdd.n12 vss 0.0104f
C905 vdd.t2 vss 0.00845f
C906 vdd.n13 vss 0.00969f
C907 vdd.t1 vss 0.00845f
C908 vdd.n14 vss 0.00969f
C909 vdd.t0 vss 0.00846f
C910 vdd.n15 vss 0.0104f
C911 vdd.t91 vss 0.00845f
C912 vdd.n16 vss 0.00958f
C913 vdd.t90 vss 0.00846f
C914 vdd.n17 vss 0.0104f
C915 vdd.t78 vss 0.00845f
C916 vdd.n18 vss 0.00964f
C917 vdd.t77 vss 0.00846f
C918 vdd.n19 vss 0.0104f
C919 vdd.t122 vss 0.00845f
C920 vdd.n20 vss 0.00961f
C921 vdd.t123 vss 0.00846f
C922 vdd.n21 vss 0.00907f
C923 vdd.n22 vss 0.00403f
C924 vdd.n23 vss 0.00176f
C925 vdd.n24 vss 0.00681f
C926 vdd.n25 vss 0.00503f
C927 vdd.n26 vss 0.00403f
C928 vdd.n27 vss 0.00176f
C929 vdd.n28 vss 0.00681f
C930 vdd.n29 vss 0.00511f
C931 vdd.n30 vss 0.00403f
C932 vdd.n31 vss 0.00176f
C933 vdd.n32 vss 0.00681f
C934 vdd.n33 vss 0.00496f
C935 vdd.n34 vss 0.00403f
C936 vdd.n35 vss 0.00176f
C937 vdd.n36 vss 0.00681f
C938 vdd.n37 vss 0.00511f
C939 vdd.n38 vss 0.00511f
C940 vdd.n39 vss 0.00176f
C941 vdd.n40 vss 0.00618f
C942 vdd.n41 vss 0.00222f
C943 vdd.n42 vss 0.00511f
C944 vdd.n43 vss 0.00176f
C945 vdd.n44 vss 0.00618f
C946 vdd.n45 vss 0.00233f
C947 vdd.n46 vss 0.00511f
C948 vdd.n47 vss 0.00176f
C949 vdd.n48 vss 0.00618f
C950 vdd.n49 vss 0.00233f
C951 vdd.n50 vss 0.00511f
C952 vdd.n51 vss 0.00176f
C953 vdd.n52 vss 0.00618f
C954 vdd.n53 vss 0.00233f
C955 vdd.n54 vss 0.00511f
C956 vdd.n55 vss 0.00176f
C957 vdd.n56 vss 0.00618f
C958 vdd.n57 vss 0.0051f
C959 vdd.n58 vss 0.269f
C960 vdd.n59 vss 0.273f
C961 vdd.n60 vss 0.00681f
C962 vdd.n61 vss 0.00403f
C963 vdd.n62 vss 0.00669f
C964 vdd.n63 vss 0.0069f
C965 vdd.t21 vss 0.00847f
C966 vdd.n64 vss 0.0118f
C967 vdd.t121 vss 0.00692f
C968 vdd.n65 vss 0.00668f
C969 vdd.t85 vss 0.00847f
C970 vdd.n66 vss 0.0116f
C971 vdd.n67 vss 0.00526f
C972 vdd.t109 vss 0.0748f
C973 vdd.t11 vss 0.035f
C974 vdd.t16 vss 0.0271f
C975 vdd.t8 vss 0.0271f
C976 vdd.t20 vss 0.0257f
C977 vdd.t120 vss 0.0339f
C978 vdd.t71 vss 0.0271f
C979 vdd.t22 vss 0.0271f
C980 vdd.t84 vss 0.0257f
C981 vdd.t100 vss 0.088f
C982 vdd.t117 vss 0.00518f
C983 vdd.n68 vss 0.0199f
C984 vdd.n69 vss 0.0222f
C985 vdd.t108 vss 0.00518f
C986 vdd.n70 vss 0.0199f
C987 vdd.n71 vss 0.0222f
C988 vdd.t149 vss 0.0375f
C989 vdd.t104 vss 0.00504f
C990 vdd.n72 vss 0.0784f
C991 vdd.n73 vss 0.0191f
C992 vdd.n74 vss 0.0243f
C993 vdd.n75 vss 0.0152f
C994 vdd.n76 vss 0.0156f
C995 vdd.t89 vss 0.00692f
C996 vdd.t61 vss 0.00692f
C997 vdd.t146 vss 0.0115f
C998 vdd.n77 vss 0.00874f
C999 vdd.n78 vss 0.104f
C1000 vdd.t30 vss 0.0637f
C1001 vdd.t44 vss 0.0517f
C1002 vdd.t38 vss 0.0517f
C1003 vdd.t31 vss 0.0517f
C1004 vdd.t45 vss 0.0387f
C1005 vdd.n79 vss 0.0504f
C1006 vdd.n80 vss 0.0258f
C1007 vdd.t34 vss 0.0387f
C1008 vdd.t28 vss 0.0517f
C1009 vdd.t41 vss 0.0517f
C1010 vdd.t37 vss 0.0517f
C1011 vdd.t29 vss 0.0637f
C1012 vdd.n81 vss 0.0251f
C1013 vdd.n82 vss 0.0151f
C1014 vdd.n83 vss 0.0611f
C1015 vdd.n84 vss 0.00106f
C1016 vdd.n85 vss 0.00138f
C1017 vdd.n86 vss 4.18e-19
C1018 vdd.n87 vss 0.001f
C1019 vdd.n88 vss 0.0179f
C1020 vdd.n89 vss 0.0646f
C1021 vdd.t148 vss 0.0375f
C1022 vdd.t107 vss 0.00504f
C1023 vdd.n90 vss 0.0784f
C1024 vdd.n91 vss 0.0191f
C1025 vdd.n92 vss 0.0243f
C1026 vdd.n93 vss 0.0152f
C1027 vdd.n94 vss 0.0156f
C1028 vdd.t145 vss 0.00692f
C1029 vdd.t43 vss 0.00692f
C1030 vdd.t152 vss 0.0115f
C1031 vdd.n95 vss 0.00874f
C1032 vdd.n96 vss 0.104f
C1033 vdd.t140 vss 0.0637f
C1034 vdd.t132 vss 0.0517f
C1035 vdd.t141 vss 0.0517f
C1036 vdd.t133 vss 0.0517f
C1037 vdd.t124 vss 0.0387f
C1038 vdd.n97 vss 0.0504f
C1039 vdd.n98 vss 0.0258f
C1040 vdd.t125 vss 0.0387f
C1041 vdd.t139 vss 0.0517f
C1042 vdd.t128 vss 0.0517f
C1043 vdd.t138 vss 0.0517f
C1044 vdd.t131 vss 0.0637f
C1045 vdd.n99 vss 0.0251f
C1046 vdd.n100 vss 0.0151f
C1047 vdd.n101 vss 0.0611f
C1048 vdd.n102 vss 0.00106f
C1049 vdd.n103 vss 0.00138f
C1050 vdd.n104 vss 4.18e-19
C1051 vdd.n105 vss 0.001f
C1052 vdd.n106 vss 0.0179f
C1053 vdd.n107 vss 0.0646f
C1054 vdd.t153 vss 0.0375f
C1055 vdd.t116 vss 0.00504f
C1056 vdd.n108 vss 0.0784f
C1057 vdd.n109 vss 0.0191f
C1058 vdd.n110 vss 0.0243f
C1059 vdd.n111 vss 0.0152f
C1060 vdd.n112 vss 0.0156f
C1061 vdd.t74 vss 0.00692f
C1062 vdd.t130 vss 0.00692f
C1063 vdd.t151 vss 0.0115f
C1064 vdd.n113 vss 0.00874f
C1065 vdd.n114 vss 0.104f
C1066 vdd.t5 vss 0.0637f
C1067 vdd.t18 vss 0.0517f
C1068 vdd.t6 vss 0.0517f
C1069 vdd.t14 vss 0.0517f
C1070 vdd.t15 vss 0.0387f
C1071 vdd.n115 vss 0.0504f
C1072 vdd.n116 vss 0.0258f
C1073 vdd.t7 vss 0.0387f
C1074 vdd.t4 vss 0.0517f
C1075 vdd.t10 vss 0.0517f
C1076 vdd.t19 vss 0.0517f
C1077 vdd.t13 vss 0.0637f
C1078 vdd.n117 vss 0.0251f
C1079 vdd.n118 vss 0.0151f
C1080 vdd.n119 vss 0.0611f
C1081 vdd.n120 vss 0.00106f
C1082 vdd.n121 vss 0.00138f
C1083 vdd.n122 vss 4.18e-19
C1084 vdd.n123 vss 0.001f
C1085 vdd.n124 vss 0.0179f
C1086 vdd.n125 vss 0.0646f
C1087 vdd.n126 vss 0.016f
C1088 vdd.n127 vss 0.00403f
C1089 vdd.n128 vss 0.00681f
C1090 vdd.n129 vss 0.00511f
C1091 vdd.n130 vss 0.00632f
C1092 vdd.t98 vss 0.00509f
C1093 vdd.n131 vss 0.00412f
C1094 vdd.n132 vss 0.0189f
C1095 vdd.n133 vss 0.0151f
C1096 vdd.t99 vss 0.00509f
C1097 vdd.n134 vss 0.0108f
C1098 vdd.n135 vss 0.00669f
C1099 vdd.n136 vss 0.0069f
C1100 vdd.n137 vss 0.00511f
C1101 vdd.n138 vss 0.00198f
C1102 vdd.n139 vss 0.00681f
C1103 vdd.t137 vss 0.00208f
C1104 vdd.t127 vss 0.00208f
C1105 vdd.n140 vss 0.00472f
C1106 vdd.n141 vss 0.00605f
C1107 vdd.n142 vss 0.00681f
C1108 vdd.n143 vss 0.00198f
C1109 vdd.n144 vss 0.00681f
C1110 vdd.n145 vss 0.00403f
C1111 vdd.t135 vss 0.00847f
C1112 vdd.n146 vss 0.0118f
C1113 vdd.n147 vss 0.00668f
C1114 vdd.n148 vss 0.00485f
C1115 vdd.n149 vss 0.00198f
C1116 vdd.n150 vss 0.00681f
C1117 vdd.t27 vss 0.00208f
C1118 vdd.t83 vss 0.00208f
C1119 vdd.n151 vss 0.00472f
C1120 vdd.n152 vss 0.00605f
C1121 vdd.n153 vss 0.00681f
C1122 vdd.n154 vss 0.00198f
C1123 vdd.n155 vss 0.00681f
C1124 vdd.t80 vss 0.00847f
C1125 vdd.n156 vss 0.0116f
C1126 vdd.n157 vss 0.00403f
C1127 vdd.n158 vss 0.0116f
C1128 vdd.n159 vss 0.0135f
C1129 vdd.n160 vss 0.0132f
C1130 vdd.n161 vss 0.00909f
C1131 vdd.n162 vss 0.00526f
C1132 vdd.n163 vss 0.016f
C1133 vdd.n164 vss 0.00403f
C1134 vdd.n165 vss 0.00681f
C1135 vdd.n166 vss 0.00511f
C1136 vdd.n167 vss 0.00632f
C1137 vdd.t95 vss 0.00509f
C1138 vdd.n168 vss 0.00412f
C1139 vdd.n169 vss 0.0189f
C1140 vdd.n170 vss 0.0151f
C1141 vdd.t96 vss 0.00509f
C1142 vdd.n171 vss 0.0108f
C1143 vdd.n172 vss 0.00669f
C1144 vdd.n173 vss 0.0069f
C1145 vdd.n174 vss 0.00511f
C1146 vdd.n175 vss 0.00198f
C1147 vdd.n176 vss 0.00681f
C1148 vdd.t36 vss 0.00208f
C1149 vdd.t40 vss 0.00208f
C1150 vdd.n177 vss 0.00472f
C1151 vdd.n178 vss 0.00605f
C1152 vdd.n179 vss 0.00681f
C1153 vdd.n180 vss 0.00198f
C1154 vdd.n181 vss 0.00681f
C1155 vdd.n182 vss 0.00403f
C1156 vdd.t33 vss 0.00847f
C1157 vdd.n183 vss 0.0118f
C1158 vdd.n184 vss 0.00668f
C1159 vdd.n185 vss 0.00485f
C1160 vdd.n186 vss 0.00198f
C1161 vdd.n187 vss 0.00681f
C1162 vdd.t87 vss 0.00208f
C1163 vdd.t25 vss 0.00208f
C1164 vdd.n188 vss 0.00472f
C1165 vdd.n189 vss 0.00605f
C1166 vdd.n190 vss 0.00681f
C1167 vdd.n191 vss 0.00198f
C1168 vdd.n192 vss 0.00681f
C1169 vdd.t68 vss 0.00847f
C1170 vdd.n193 vss 0.0116f
C1171 vdd.n194 vss 0.00403f
C1172 vdd.n195 vss 0.0116f
C1173 vdd.n196 vss 0.0135f
C1174 vdd.n197 vss 0.0132f
C1175 vdd.n198 vss 0.00909f
C1176 vdd.n199 vss 0.00526f
C1177 vdd.n200 vss 0.016f
C1178 vdd.n201 vss 0.00403f
C1179 vdd.n202 vss 0.00681f
C1180 vdd.n203 vss 0.00511f
C1181 vdd.n204 vss 0.00632f
C1182 vdd.t113 vss 0.00509f
C1183 vdd.n205 vss 0.00412f
C1184 vdd.n206 vss 0.0189f
C1185 vdd.n207 vss 0.0151f
C1186 vdd.t114 vss 0.00509f
C1187 vdd.n208 vss 0.0108f
C1188 vdd.n209 vss 0.00669f
C1189 vdd.n210 vss 0.0069f
C1190 vdd.n211 vss 0.00511f
C1191 vdd.n212 vss 0.00198f
C1192 vdd.n213 vss 0.00681f
C1193 vdd.t52 vss 0.00208f
C1194 vdd.t58 vss 0.00208f
C1195 vdd.n214 vss 0.00472f
C1196 vdd.n215 vss 0.00605f
C1197 vdd.n216 vss 0.00681f
C1198 vdd.n217 vss 0.00198f
C1199 vdd.n218 vss 0.00681f
C1200 vdd.n219 vss 0.00403f
C1201 vdd.t49 vss 0.00847f
C1202 vdd.n220 vss 0.0118f
C1203 vdd.n221 vss 0.00668f
C1204 vdd.n222 vss 0.00485f
C1205 vdd.n223 vss 0.00198f
C1206 vdd.n224 vss 0.00681f
C1207 vdd.t76 vss 0.00208f
C1208 vdd.t119 vss 0.00208f
C1209 vdd.n225 vss 0.00472f
C1210 vdd.n226 vss 0.00605f
C1211 vdd.n227 vss 0.00681f
C1212 vdd.n228 vss 0.00198f
C1213 vdd.n229 vss 0.00681f
C1214 vdd.t70 vss 0.00847f
C1215 vdd.n230 vss 0.0116f
C1216 vdd.n231 vss 0.00403f
C1217 vdd.n232 vss 0.0116f
C1218 vdd.n233 vss 0.0135f
C1219 vdd.n234 vss 0.104f
C1220 vdd.t54 vss 0.0637f
C1221 vdd.t62 vss 0.0517f
C1222 vdd.t55 vss 0.0517f
C1223 vdd.t65 vss 0.0517f
C1224 vdd.t56 vss 0.0387f
C1225 vdd.n235 vss 0.0504f
C1226 vdd.n236 vss 0.0258f
C1227 vdd.t50 vss 0.0387f
C1228 vdd.t63 vss 0.0517f
C1229 vdd.t59 vss 0.0517f
C1230 vdd.t53 vss 0.0517f
C1231 vdd.t64 vss 0.0637f
C1232 vdd.n237 vss 0.0251f
C1233 vdd.n238 vss 0.0151f
C1234 vdd.n239 vss 0.0611f
C1235 vdd.n240 vss 0.00106f
C1236 vdd.n241 vss 0.00138f
C1237 vdd.n242 vss 4.18e-19
C1238 vdd.n243 vss 0.001f
C1239 vdd.n244 vss 0.0179f
C1240 vdd.n245 vss 0.0646f
C1241 vdd.n246 vss 0.016f
C1242 vdd.n247 vss 0.0111f
C1243 vdd.n248 vss 0.00909f
C1244 vdd.n249 vss 0.0132f
C1245 vdd.t105 vss 0.00518f
C1246 vdd.n250 vss 0.0216f
C1247 vdd.n251 vss 0.0222f
C1248 vdd.n252 vss 0.0597f
C1249 vdd.t103 vss 0.088f
C1250 vdd.t69 vss 0.0257f
C1251 vdd.t118 vss 0.0271f
C1252 vdd.t75 vss 0.0271f
C1253 vdd.t88 vss 0.0339f
C1254 vdd.t48 vss 0.0257f
C1255 vdd.t57 vss 0.0271f
C1256 vdd.t51 vss 0.0271f
C1257 vdd.t60 vss 0.035f
C1258 vdd.t112 vss 0.0446f
C1259 vdd.n253 vss 0.0597f
C1260 vdd.t106 vss 0.088f
C1261 vdd.t67 vss 0.0257f
C1262 vdd.t24 vss 0.0271f
C1263 vdd.t86 vss 0.0271f
C1264 vdd.t144 vss 0.0339f
C1265 vdd.t32 vss 0.0257f
C1266 vdd.t39 vss 0.0271f
C1267 vdd.t35 vss 0.0271f
C1268 vdd.t42 vss 0.035f
C1269 vdd.t94 vss 0.0446f
C1270 vdd.n254 vss 0.0597f
C1271 vdd.t115 vss 0.088f
C1272 vdd.t79 vss 0.0257f
C1273 vdd.t82 vss 0.0271f
C1274 vdd.t26 vss 0.0271f
C1275 vdd.t73 vss 0.0339f
C1276 vdd.t134 vss 0.0257f
C1277 vdd.t126 vss 0.0271f
C1278 vdd.t136 vss 0.0271f
C1279 vdd.t129 vss 0.035f
C1280 vdd.t97 vss 0.0446f
C1281 vdd.n255 vss 0.0597f
C1282 vdd.t102 vss 0.00518f
C1283 vdd.n256 vss 0.0199f
C1284 vdd.n257 vss 0.0222f
C1285 vdd.n258 vss 0.0132f
C1286 vdd.n259 vss 0.00909f
C1287 vdd.n260 vss 0.0135f
C1288 vdd.t150 vss 0.0375f
C1289 vdd.t101 vss 0.00504f
C1290 vdd.n261 vss 0.0784f
C1291 vdd.n262 vss 0.0191f
C1292 vdd.n263 vss 0.0243f
C1293 vdd.n264 vss 0.0152f
C1294 vdd.n265 vss 0.0156f
C1295 vdd.n266 vss 0.0116f
C1296 vdd.n267 vss 0.00403f
C1297 vdd.n268 vss 0.00198f
C1298 vdd.n269 vss 0.00681f
C1299 vdd.t72 vss 0.00208f
C1300 vdd.t23 vss 0.00208f
C1301 vdd.n270 vss 0.00472f
C1302 vdd.n271 vss 0.00605f
C1303 vdd.n272 vss 0.00681f
C1304 vdd.n273 vss 0.00198f
C1305 vdd.n274 vss 0.00681f
C1306 vdd.n275 vss 0.00485f
C1307 vdd.n276 vss 0.00403f
C1308 vdd.n277 vss 0.00198f
C1309 vdd.n278 vss 0.00681f
C1310 vdd.t17 vss 0.00208f
C1311 vdd.t9 vss 0.00208f
C1312 vdd.n279 vss 0.00472f
C1313 vdd.n280 vss 0.00605f
C1314 vdd.n281 vss 0.00681f
C1315 vdd.n282 vss 0.00198f
C1316 vdd.n283 vss 0.00681f
C1317 vdd.n284 vss 0.00511f
C1318 out.t1 vss 0.00463f
C1319 out.t8 vss 0.00463f
C1320 out.n0 vss 0.0301f
C1321 out.t58 vss 0.00463f
C1322 out.t55 vss 0.00463f
C1323 out.n1 vss 0.0299f
C1324 out.t2 vss 0.00463f
C1325 out.t6 vss 0.00463f
C1326 out.n2 vss 0.03f
C1327 out.t59 vss 0.00463f
C1328 out.t52 vss 0.00463f
C1329 out.n3 vss 0.0299f
C1330 out.t7 vss 0.00463f
C1331 out.t3 vss 0.00463f
C1332 out.n4 vss 0.0299f
C1333 out.t53 vss 0.00463f
C1334 out.t50 vss 0.00463f
C1335 out.n5 vss 0.03f
C1336 out.t0 vss 0.00463f
C1337 out.t4 vss 0.00463f
C1338 out.n6 vss 0.0301f
C1339 out.t57 vss 0.00463f
C1340 out.t54 vss 0.00463f
C1341 out.n7 vss 0.0302f
C1342 out.t9 vss 0.00463f
C1343 out.t5 vss 0.00463f
C1344 out.n8 vss 0.0299f
C1345 out.t56 vss 0.00463f
C1346 out.t51 vss 0.00463f
C1347 out.n9 vss 0.0302f
C1348 out.n10 vss 0.0203f
C1349 out.n11 vss 0.0263f
C1350 out.n12 vss 0.0265f
C1351 out.n13 vss 0.0263f
C1352 out.n14 vss 0.0273f
C1353 out.t78 vss 0.00463f
C1354 out.t74 vss 0.00463f
C1355 out.n15 vss 0.0301f
C1356 out.t33 vss 0.00463f
C1357 out.t39 vss 0.00463f
C1358 out.n16 vss 0.0299f
C1359 out.t79 vss 0.00463f
C1360 out.t75 vss 0.00463f
C1361 out.n17 vss 0.03f
C1362 out.t34 vss 0.00463f
C1363 out.t30 vss 0.00463f
C1364 out.n18 vss 0.0299f
C1365 out.t70 vss 0.00463f
C1366 out.t71 vss 0.00463f
C1367 out.n19 vss 0.0299f
C1368 out.t35 vss 0.00463f
C1369 out.t36 vss 0.00463f
C1370 out.n20 vss 0.03f
C1371 out.t77 vss 0.00463f
C1372 out.t72 vss 0.00463f
C1373 out.n21 vss 0.0301f
C1374 out.t31 vss 0.00463f
C1375 out.t37 vss 0.00463f
C1376 out.n22 vss 0.0302f
C1377 out.t76 vss 0.00463f
C1378 out.t73 vss 0.00463f
C1379 out.n23 vss 0.0299f
C1380 out.t32 vss 0.00463f
C1381 out.t38 vss 0.00463f
C1382 out.n24 vss 0.0302f
C1383 out.n25 vss 0.0203f
C1384 out.n26 vss 0.0263f
C1385 out.n27 vss 0.0265f
C1386 out.n28 vss 0.0263f
C1387 out.n29 vss 0.0273f
C1388 out.t12 vss 0.00463f
C1389 out.t18 vss 0.00463f
C1390 out.n30 vss 0.0301f
C1391 out.t41 vss 0.00463f
C1392 out.t45 vss 0.00463f
C1393 out.n31 vss 0.0299f
C1394 out.t16 vss 0.00463f
C1395 out.t13 vss 0.00463f
C1396 out.n32 vss 0.03f
C1397 out.t42 vss 0.00463f
C1398 out.t49 vss 0.00463f
C1399 out.n33 vss 0.0299f
C1400 out.t19 vss 0.00463f
C1401 out.t14 vss 0.00463f
C1402 out.n34 vss 0.0299f
C1403 out.t46 vss 0.00463f
C1404 out.t43 vss 0.00463f
C1405 out.n35 vss 0.03f
C1406 out.t10 vss 0.00463f
C1407 out.t17 vss 0.00463f
C1408 out.n36 vss 0.0301f
C1409 out.t47 vss 0.00463f
C1410 out.t44 vss 0.00463f
C1411 out.n37 vss 0.0302f
C1412 out.t15 vss 0.00463f
C1413 out.t11 vss 0.00463f
C1414 out.n38 vss 0.0299f
C1415 out.t40 vss 0.00463f
C1416 out.t48 vss 0.00463f
C1417 out.n39 vss 0.0302f
C1418 out.n40 vss 0.0203f
C1419 out.n41 vss 0.0263f
C1420 out.n42 vss 0.0265f
C1421 out.n43 vss 0.0263f
C1422 out.n44 vss 0.0273f
C1423 out.t22 vss 0.00463f
C1424 out.t26 vss 0.00463f
C1425 out.n45 vss 0.0301f
C1426 out.t69 vss 0.00463f
C1427 out.t64 vss 0.00463f
C1428 out.n46 vss 0.0299f
C1429 out.t23 vss 0.00463f
C1430 out.t29 vss 0.00463f
C1431 out.n47 vss 0.03f
C1432 out.t60 vss 0.00463f
C1433 out.t65 vss 0.00463f
C1434 out.n48 vss 0.0299f
C1435 out.t24 vss 0.00463f
C1436 out.t20 vss 0.00463f
C1437 out.n49 vss 0.0299f
C1438 out.t61 vss 0.00463f
C1439 out.t66 vss 0.00463f
C1440 out.n50 vss 0.03f
C1441 out.t27 vss 0.00463f
C1442 out.t25 vss 0.00463f
C1443 out.n51 vss 0.0301f
C1444 out.t67 vss 0.00463f
C1445 out.t62 vss 0.00463f
C1446 out.n52 vss 0.0302f
C1447 out.t21 vss 0.00463f
C1448 out.t28 vss 0.00463f
C1449 out.n53 vss 0.0299f
C1450 out.t68 vss 0.00463f
C1451 out.t63 vss 0.00463f
C1452 out.n54 vss 0.0302f
C1453 out.n55 vss 0.0203f
C1454 out.n56 vss 0.0263f
C1455 out.n57 vss 0.0265f
C1456 out.n58 vss 0.0263f
C1457 out.n59 vss 0.0273f
C1458 out.t258 vss 0.375f
C1459 out.t165 vss 0.255f
C1460 out.n60 vss 0.139f
C1461 out.t111 vss 0.255f
C1462 out.n61 vss 0.139f
C1463 out.t395 vss 0.255f
C1464 out.n62 vss 0.139f
C1465 out.t342 vss 0.255f
C1466 out.n63 vss 0.139f
C1467 out.t286 vss 0.255f
C1468 out.n64 vss 0.139f
C1469 out.t193 vss 0.255f
C1470 out.n65 vss 0.139f
C1471 out.t138 vss 0.255f
C1472 out.n66 vss 0.139f
C1473 out.t279 vss 0.255f
C1474 out.n67 vss 0.139f
C1475 out.t226 vss 0.255f
C1476 out.n68 vss 0.139f
C1477 out.t175 vss 0.255f
C1478 out.n69 vss 0.139f
C1479 out.t80 vss 0.255f
C1480 out.n70 vss 0.139f
C1481 out.t366 vss 0.255f
C1482 out.n71 vss 0.139f
C1483 out.t312 vss 0.255f
C1484 out.n72 vss 0.139f
C1485 out.t259 vss 0.255f
C1486 out.n73 vss 0.139f
C1487 out.t205 vss 0.255f
C1488 out.n74 vss 0.139f
C1489 out.t112 vss 0.255f
C1490 out.n75 vss 0.139f
C1491 out.t397 vss 0.255f
C1492 out.n76 vss 0.139f
C1493 out.t345 vss 0.255f
C1494 out.n77 vss 0.139f
C1495 out.t287 vss 0.255f
C1496 out.n78 vss 0.139f
C1497 out.t170 vss 0.255f
C1498 out.n79 vss 0.139f
C1499 out.t417 vss 0.255f
C1500 out.n80 vss 0.139f
C1501 out.t361 vss 0.255f
C1502 out.n81 vss 0.139f
C1503 out.t307 vss 0.255f
C1504 out.n82 vss 0.139f
C1505 out.t254 vss 0.255f
C1506 out.n83 vss 0.139f
C1507 out.t200 vss 0.255f
C1508 out.n84 vss 0.139f
C1509 out.t105 vss 0.255f
C1510 out.n85 vss 0.139f
C1511 out.t390 vss 0.255f
C1512 out.t336 vss 0.255f
C1513 out.t281 vss 0.255f
C1514 out.t228 vss 0.255f
C1515 out.t134 vss 0.255f
C1516 out.t110 vss 0.255f
C1517 out.n86 vss 0.115f
C1518 out.t339 vss 0.255f
C1519 out.t150 vss 0.375f
C1520 out.t394 vss 0.255f
C1521 out.n87 vss 0.139f
C1522 out.t340 vss 0.255f
C1523 out.n88 vss 0.139f
C1524 out.t284 vss 0.255f
C1525 out.n89 vss 0.139f
C1526 out.t234 vss 0.255f
C1527 out.n90 vss 0.139f
C1528 out.t180 vss 0.255f
C1529 out.n91 vss 0.139f
C1530 out.t84 vss 0.255f
C1531 out.n92 vss 0.139f
C1532 out.t370 vss 0.255f
C1533 out.n93 vss 0.139f
C1534 out.t172 vss 0.255f
C1535 out.n94 vss 0.139f
C1536 out.t119 vss 0.255f
C1537 out.n95 vss 0.139f
C1538 out.t405 vss 0.255f
C1539 out.n96 vss 0.139f
C1540 out.t310 vss 0.255f
C1541 out.n97 vss 0.139f
C1542 out.t256 vss 0.255f
C1543 out.n98 vss 0.139f
C1544 out.t204 vss 0.255f
C1545 out.n99 vss 0.139f
C1546 out.t151 vss 0.255f
C1547 out.n100 vss 0.139f
C1548 out.t95 vss 0.255f
C1549 out.n101 vss 0.139f
C1550 out.t341 vss 0.255f
C1551 out.n102 vss 0.139f
C1552 out.t285 vss 0.255f
C1553 out.n103 vss 0.139f
C1554 out.t235 vss 0.255f
C1555 out.n104 vss 0.139f
C1556 out.t181 vss 0.255f
C1557 out.n105 vss 0.139f
C1558 out.t401 vss 0.255f
C1559 out.n106 vss 0.139f
C1560 out.t306 vss 0.255f
C1561 out.n107 vss 0.139f
C1562 out.t252 vss 0.255f
C1563 out.n108 vss 0.139f
C1564 out.t199 vss 0.255f
C1565 out.n109 vss 0.139f
C1566 out.t145 vss 0.255f
C1567 out.n110 vss 0.139f
C1568 out.t89 vss 0.255f
C1569 out.n111 vss 0.139f
C1570 out.t334 vss 0.255f
C1571 out.n112 vss 0.139f
C1572 out.t280 vss 0.255f
C1573 out.n113 vss 0.139f
C1574 out.t227 vss 0.255f
C1575 out.n114 vss 0.139f
C1576 out.t174 vss 0.255f
C1577 out.n115 vss 0.139f
C1578 out.t120 vss 0.255f
C1579 out.n116 vss 0.139f
C1580 out.t365 vss 0.255f
C1581 out.n117 vss 0.139f
C1582 out.t413 vss 0.255f
C1583 out.t221 vss 0.375f
C1584 out.t127 vss 0.255f
C1585 out.n118 vss 0.139f
C1586 out.t414 vss 0.255f
C1587 out.n119 vss 0.139f
C1588 out.t358 vss 0.255f
C1589 out.n120 vss 0.139f
C1590 out.t304 vss 0.255f
C1591 out.n121 vss 0.139f
C1592 out.t250 vss 0.255f
C1593 out.n122 vss 0.139f
C1594 out.t157 vss 0.255f
C1595 out.n123 vss 0.139f
C1596 out.t102 vss 0.255f
C1597 out.n124 vss 0.139f
C1598 out.t243 vss 0.255f
C1599 out.n125 vss 0.139f
C1600 out.t189 vss 0.255f
C1601 out.n126 vss 0.139f
C1602 out.t136 vss 0.255f
C1603 out.n127 vss 0.139f
C1604 out.t384 vss 0.255f
C1605 out.n128 vss 0.139f
C1606 out.t328 vss 0.255f
C1607 out.n129 vss 0.139f
C1608 out.t275 vss 0.255f
C1609 out.n130 vss 0.139f
C1610 out.t222 vss 0.255f
C1611 out.n131 vss 0.139f
C1612 out.t169 vss 0.255f
C1613 out.n132 vss 0.139f
C1614 out.t415 vss 0.255f
C1615 out.n133 vss 0.139f
C1616 out.t360 vss 0.255f
C1617 out.n134 vss 0.139f
C1618 out.t305 vss 0.255f
C1619 out.n135 vss 0.139f
C1620 out.t251 vss 0.255f
C1621 out.n136 vss 0.139f
C1622 out.t131 vss 0.255f
C1623 out.n137 vss 0.139f
C1624 out.t378 vss 0.255f
C1625 out.n138 vss 0.139f
C1626 out.t321 vss 0.255f
C1627 out.n139 vss 0.139f
C1628 out.t272 vss 0.255f
C1629 out.n140 vss 0.139f
C1630 out.t216 vss 0.255f
C1631 out.n141 vss 0.139f
C1632 out.t164 vss 0.255f
C1633 out.n142 vss 0.139f
C1634 out.t408 vss 0.255f
C1635 out.n143 vss 0.139f
C1636 out.t354 vss 0.255f
C1637 out.n144 vss 0.139f
C1638 out.t299 vss 0.255f
C1639 out.n145 vss 0.139f
C1640 out.t245 vss 0.255f
C1641 out.n146 vss 0.139f
C1642 out.t191 vss 0.255f
C1643 out.n147 vss 0.139f
C1644 out.t98 vss 0.255f
C1645 out.n148 vss 0.139f
C1646 out.t301 vss 0.255f
C1647 out.t115 vss 0.375f
C1648 out.t357 vss 0.255f
C1649 out.n149 vss 0.139f
C1650 out.t302 vss 0.255f
C1651 out.n150 vss 0.139f
C1652 out.t248 vss 0.255f
C1653 out.n151 vss 0.139f
C1654 out.t197 vss 0.255f
C1655 out.n152 vss 0.139f
C1656 out.t143 vss 0.255f
C1657 out.n153 vss 0.139f
C1658 out.t388 vss 0.255f
C1659 out.n154 vss 0.139f
C1660 out.t333 vss 0.255f
C1661 out.n155 vss 0.139f
C1662 out.t133 vss 0.255f
C1663 out.n156 vss 0.139f
C1664 out.t81 vss 0.255f
C1665 out.n157 vss 0.139f
C1666 out.t369 vss 0.255f
C1667 out.n158 vss 0.139f
C1668 out.t273 vss 0.255f
C1669 out.n159 vss 0.139f
C1670 out.t219 vss 0.255f
C1671 out.n160 vss 0.139f
C1672 out.t168 vss 0.255f
C1673 out.n161 vss 0.139f
C1674 out.t116 vss 0.255f
C1675 out.n162 vss 0.139f
C1676 out.t400 vss 0.255f
C1677 out.n163 vss 0.139f
C1678 out.t303 vss 0.255f
C1679 out.n164 vss 0.139f
C1680 out.t249 vss 0.255f
C1681 out.n165 vss 0.139f
C1682 out.t198 vss 0.255f
C1683 out.n166 vss 0.139f
C1684 out.t144 vss 0.255f
C1685 out.n167 vss 0.139f
C1686 out.t364 vss 0.255f
C1687 out.n168 vss 0.139f
C1688 out.t269 vss 0.255f
C1689 out.n169 vss 0.139f
C1690 out.t214 vss 0.255f
C1691 out.n170 vss 0.139f
C1692 out.t163 vss 0.255f
C1693 out.n171 vss 0.139f
C1694 out.t109 vss 0.255f
C1695 out.n172 vss 0.139f
C1696 out.t393 vss 0.255f
C1697 out.n173 vss 0.139f
C1698 out.t298 vss 0.255f
C1699 out.n174 vss 0.139f
C1700 out.t244 vss 0.255f
C1701 out.n175 vss 0.139f
C1702 out.t190 vss 0.255f
C1703 out.n176 vss 0.139f
C1704 out.t137 vss 0.255f
C1705 out.n177 vss 0.139f
C1706 out.t83 vss 0.255f
C1707 out.n178 vss 0.139f
C1708 out.t330 vss 0.255f
C1709 out.n179 vss 0.139f
C1710 out.t192 vss 0.255f
C1711 out.t344 vss 0.375f
C1712 out.t247 vss 0.255f
C1713 out.n180 vss 0.139f
C1714 out.t194 vss 0.255f
C1715 out.n181 vss 0.139f
C1716 out.t140 vss 0.255f
C1717 out.n182 vss 0.139f
C1718 out.t85 vss 0.255f
C1719 out.n183 vss 0.139f
C1720 out.t372 vss 0.255f
C1721 out.n184 vss 0.139f
C1722 out.t278 vss 0.255f
C1723 out.n185 vss 0.139f
C1724 out.t224 vss 0.255f
C1725 out.n186 vss 0.139f
C1726 out.t367 vss 0.255f
C1727 out.n187 vss 0.139f
C1728 out.t313 vss 0.255f
C1729 out.n188 vss 0.139f
C1730 out.t260 vss 0.255f
C1731 out.n189 vss 0.139f
C1732 out.t166 vss 0.255f
C1733 out.n190 vss 0.139f
C1734 out.t113 vss 0.255f
C1735 out.n191 vss 0.139f
C1736 out.t399 vss 0.255f
C1737 out.n192 vss 0.139f
C1738 out.t347 vss 0.255f
C1739 out.n193 vss 0.139f
C1740 out.t290 vss 0.255f
C1741 out.n194 vss 0.139f
C1742 out.t196 vss 0.255f
C1743 out.n195 vss 0.139f
C1744 out.t141 vss 0.255f
C1745 out.n196 vss 0.139f
C1746 out.t86 vss 0.255f
C1747 out.n197 vss 0.139f
C1748 out.t375 vss 0.255f
C1749 out.n198 vss 0.139f
C1750 out.t255 vss 0.255f
C1751 out.n199 vss 0.139f
C1752 out.t161 vss 0.255f
C1753 out.n200 vss 0.139f
C1754 out.t108 vss 0.255f
C1755 out.n201 vss 0.139f
C1756 out.t392 vss 0.255f
C1757 out.n202 vss 0.139f
C1758 out.t338 vss 0.255f
C1759 out.n203 vss 0.139f
C1760 out.t282 vss 0.255f
C1761 out.n204 vss 0.139f
C1762 out.t188 vss 0.255f
C1763 out.n205 vss 0.139f
C1764 out.t135 vss 0.255f
C1765 out.n206 vss 0.139f
C1766 out.t82 vss 0.255f
C1767 out.n207 vss 0.139f
C1768 out.t368 vss 0.255f
C1769 out.n208 vss 0.139f
C1770 out.t314 vss 0.255f
C1771 out.n209 vss 0.139f
C1772 out.t220 vss 0.255f
C1773 out.n210 vss 0.139f
C1774 out.t266 vss 0.255f
C1775 out.t419 vss 0.375f
C1776 out.t320 vss 0.255f
C1777 out.n211 vss 0.139f
C1778 out.t268 vss 0.255f
C1779 out.n212 vss 0.139f
C1780 out.t213 vss 0.255f
C1781 out.n213 vss 0.139f
C1782 out.t159 vss 0.255f
C1783 out.n214 vss 0.139f
C1784 out.t107 vss 0.255f
C1785 out.n215 vss 0.139f
C1786 out.t353 vss 0.255f
C1787 out.n216 vss 0.139f
C1788 out.t297 vss 0.255f
C1789 out.n217 vss 0.139f
C1790 out.t97 vss 0.255f
C1791 out.n218 vss 0.139f
C1792 out.t385 vss 0.255f
C1793 out.n219 vss 0.139f
C1794 out.t331 vss 0.255f
C1795 out.n220 vss 0.139f
C1796 out.t238 vss 0.255f
C1797 out.n221 vss 0.139f
C1798 out.t183 vss 0.255f
C1799 out.n222 vss 0.139f
C1800 out.t130 vss 0.255f
C1801 out.n223 vss 0.139f
C1802 out.t418 vss 0.255f
C1803 out.n224 vss 0.139f
C1804 out.t363 vss 0.255f
C1805 out.n225 vss 0.139f
C1806 out.t267 vss 0.255f
C1807 out.n226 vss 0.139f
C1808 out.t212 vss 0.255f
C1809 out.n227 vss 0.139f
C1810 out.t162 vss 0.255f
C1811 out.n228 vss 0.139f
C1812 out.t106 vss 0.255f
C1813 out.n229 vss 0.139f
C1814 out.t326 vss 0.255f
C1815 out.n230 vss 0.139f
C1816 out.t233 vss 0.255f
C1817 out.n231 vss 0.139f
C1818 out.t178 vss 0.255f
C1819 out.n232 vss 0.139f
C1820 out.t123 vss 0.255f
C1821 out.n233 vss 0.139f
C1822 out.t412 vss 0.255f
C1823 out.n234 vss 0.139f
C1824 out.t356 vss 0.255f
C1825 out.n235 vss 0.139f
C1826 out.t262 vss 0.255f
C1827 out.n236 vss 0.139f
C1828 out.t207 vss 0.255f
C1829 out.n237 vss 0.139f
C1830 out.t153 vss 0.255f
C1831 out.n238 vss 0.139f
C1832 out.t101 vss 0.255f
C1833 out.n239 vss 0.139f
C1834 out.t387 vss 0.255f
C1835 out.n240 vss 0.139f
C1836 out.t293 vss 0.255f
C1837 out.n241 vss 0.139f
C1838 out.t156 vss 0.255f
C1839 out.t309 vss 0.375f
C1840 out.t211 vss 0.255f
C1841 out.n242 vss 0.139f
C1842 out.t158 vss 0.255f
C1843 out.n243 vss 0.139f
C1844 out.t104 vss 0.255f
C1845 out.n244 vss 0.139f
C1846 out.t389 vss 0.255f
C1847 out.n245 vss 0.139f
C1848 out.t335 vss 0.255f
C1849 out.n246 vss 0.139f
C1850 out.t242 vss 0.255f
C1851 out.n247 vss 0.139f
C1852 out.t187 vss 0.255f
C1853 out.n248 vss 0.139f
C1854 out.t329 vss 0.255f
C1855 out.n249 vss 0.139f
C1856 out.t276 vss 0.255f
C1857 out.n250 vss 0.139f
C1858 out.t223 vss 0.255f
C1859 out.n251 vss 0.139f
C1860 out.t129 vss 0.255f
C1861 out.n252 vss 0.139f
C1862 out.t416 vss 0.255f
C1863 out.n253 vss 0.139f
C1864 out.t362 vss 0.255f
C1865 out.n254 vss 0.139f
C1866 out.t308 vss 0.255f
C1867 out.n255 vss 0.139f
C1868 out.t253 vss 0.255f
C1869 out.n256 vss 0.139f
C1870 out.t160 vss 0.255f
C1871 out.n257 vss 0.139f
C1872 out.t103 vss 0.255f
C1873 out.n258 vss 0.139f
C1874 out.t391 vss 0.255f
C1875 out.n259 vss 0.139f
C1876 out.t337 vss 0.255f
C1877 out.n260 vss 0.139f
C1878 out.t218 vss 0.255f
C1879 out.n261 vss 0.139f
C1880 out.t124 vss 0.255f
C1881 out.n262 vss 0.139f
C1882 out.t409 vss 0.255f
C1883 out.n263 vss 0.139f
C1884 out.t355 vss 0.255f
C1885 out.n264 vss 0.139f
C1886 out.t300 vss 0.255f
C1887 out.n265 vss 0.139f
C1888 out.t246 vss 0.255f
C1889 out.n266 vss 0.139f
C1890 out.t152 vss 0.255f
C1891 out.n267 vss 0.139f
C1892 out.t99 vss 0.255f
C1893 out.n268 vss 0.139f
C1894 out.t386 vss 0.255f
C1895 out.n269 vss 0.139f
C1896 out.t332 vss 0.255f
C1897 out.n270 vss 0.139f
C1898 out.t277 vss 0.255f
C1899 out.n271 vss 0.139f
C1900 out.t184 vss 0.255f
C1901 out.n272 vss 0.139f
C1902 out.t349 vss 0.255f
C1903 out.t294 vss 0.255f
C1904 out.t201 vss 0.255f
C1905 out.t147 vss 0.255f
C1906 out.t91 vss 0.255f
C1907 out.t380 vss 0.255f
C1908 out.t324 vss 0.255f
C1909 out.t230 vss 0.255f
C1910 out.t177 vss 0.255f
C1911 out.t316 vss 0.255f
C1912 out.t263 vss 0.255f
C1913 out.t210 vss 0.255f
C1914 out.t117 vss 0.255f
C1915 out.t402 vss 0.255f
C1916 out.t351 vss 0.255f
C1917 out.t295 vss 0.255f
C1918 out.t241 vss 0.255f
C1919 out.t148 vss 0.255f
C1920 out.t92 vss 0.255f
C1921 out.t383 vss 0.255f
C1922 out.t325 vss 0.255f
C1923 out.t206 vss 0.255f
C1924 out.t114 vss 0.255f
C1925 out.t398 vss 0.255f
C1926 out.t346 vss 0.255f
C1927 out.t291 vss 0.255f
C1928 out.t237 vss 0.255f
C1929 out.t142 vss 0.255f
C1930 out.t87 vss 0.255f
C1931 out.t373 vss 0.255f
C1932 out.t319 vss 0.255f
C1933 out.t265 vss 0.255f
C1934 out.t173 vss 0.255f
C1935 out.t146 vss 0.255f
C1936 out.t376 vss 0.255f
C1937 out.t185 vss 0.375f
C1938 out.t90 vss 0.255f
C1939 out.n273 vss 0.139f
C1940 out.t377 vss 0.255f
C1941 out.n274 vss 0.139f
C1942 out.t322 vss 0.255f
C1943 out.n275 vss 0.139f
C1944 out.t270 vss 0.255f
C1945 out.n276 vss 0.139f
C1946 out.t215 vss 0.255f
C1947 out.n277 vss 0.139f
C1948 out.t121 vss 0.255f
C1949 out.n278 vss 0.139f
C1950 out.t407 vss 0.255f
C1951 out.n279 vss 0.139f
C1952 out.t208 vss 0.255f
C1953 out.n280 vss 0.139f
C1954 out.t154 vss 0.255f
C1955 out.n281 vss 0.139f
C1956 out.t100 vss 0.255f
C1957 out.n282 vss 0.139f
C1958 out.t348 vss 0.255f
C1959 out.n283 vss 0.139f
C1960 out.t292 vss 0.255f
C1961 out.n284 vss 0.139f
C1962 out.t240 vss 0.255f
C1963 out.n285 vss 0.139f
C1964 out.t186 vss 0.255f
C1965 out.n286 vss 0.139f
C1966 out.t132 vss 0.255f
C1967 out.n287 vss 0.139f
C1968 out.t379 vss 0.255f
C1969 out.n288 vss 0.139f
C1970 out.t323 vss 0.255f
C1971 out.n289 vss 0.139f
C1972 out.t271 vss 0.255f
C1973 out.n290 vss 0.139f
C1974 out.t217 vss 0.255f
C1975 out.n291 vss 0.139f
C1976 out.t96 vss 0.255f
C1977 out.n292 vss 0.139f
C1978 out.t343 vss 0.255f
C1979 out.n293 vss 0.139f
C1980 out.t288 vss 0.255f
C1981 out.n294 vss 0.139f
C1982 out.t236 vss 0.255f
C1983 out.n295 vss 0.139f
C1984 out.t182 vss 0.255f
C1985 out.n296 vss 0.139f
C1986 out.t126 vss 0.255f
C1987 out.n297 vss 0.139f
C1988 out.t371 vss 0.255f
C1989 out.n298 vss 0.139f
C1990 out.t317 vss 0.255f
C1991 out.n299 vss 0.139f
C1992 out.t264 vss 0.255f
C1993 out.n300 vss 0.139f
C1994 out.t209 vss 0.255f
C1995 out.n301 vss 0.139f
C1996 out.t155 vss 0.255f
C1997 out.n302 vss 0.139f
C1998 out.t404 vss 0.255f
C1999 out.n303 vss 0.139f
C2000 out.n304 vss 0.0498f
C2001 out.n305 vss 0.111f
C2002 out.n306 vss 0.0556f
C2003 out.n307 vss 0.106f
C2004 out.n308 vss 0.139f
C2005 out.n309 vss 0.139f
C2006 out.n310 vss 0.139f
C2007 out.n311 vss 0.139f
C2008 out.n312 vss 0.139f
C2009 out.n313 vss 0.139f
C2010 out.n314 vss 0.139f
C2011 out.n315 vss 0.139f
C2012 out.n316 vss 0.139f
C2013 out.n317 vss 0.139f
C2014 out.n318 vss 0.139f
C2015 out.n319 vss 0.139f
C2016 out.n320 vss 0.139f
C2017 out.n321 vss 0.139f
C2018 out.n322 vss 0.139f
C2019 out.n323 vss 0.139f
C2020 out.n324 vss 0.139f
C2021 out.n325 vss 0.139f
C2022 out.n326 vss 0.139f
C2023 out.n327 vss 0.139f
C2024 out.n328 vss 0.139f
C2025 out.n329 vss 0.139f
C2026 out.n330 vss 0.139f
C2027 out.n331 vss 0.139f
C2028 out.n332 vss 0.139f
C2029 out.n333 vss 0.139f
C2030 out.n334 vss 0.139f
C2031 out.n335 vss 0.139f
C2032 out.n336 vss 0.139f
C2033 out.n337 vss 0.139f
C2034 out.n338 vss 0.139f
C2035 out.n339 vss 0.139f
C2036 out.n340 vss 0.138f
C2037 out.t239 vss 0.255f
C2038 out.n341 vss 0.118f
C2039 out.t311 vss 0.255f
C2040 out.n342 vss 0.118f
C2041 out.t203 vss 0.255f
C2042 out.n343 vss 0.118f
C2043 out.t274 vss 0.255f
C2044 out.n344 vss 0.118f
C2045 out.t167 vss 0.255f
C2046 out.n345 vss 0.118f
C2047 out.t396 vss 0.255f
C2048 out.n346 vss 0.118f
C2049 out.t128 vss 0.255f
C2050 out.n347 vss 0.118f
C2051 out.t359 vss 0.255f
C2052 out.n348 vss 0.118f
C2053 out.t94 vss 0.255f
C2054 out.n349 vss 0.0928f
C2055 out.n350 vss 0.0534f
C2056 out.t382 vss 0.255f
C2057 out.n351 vss 0.139f
C2058 out.t283 vss 0.255f
C2059 out.n352 vss 0.139f
C2060 out.t232 vss 0.255f
C2061 out.n353 vss 0.139f
C2062 out.t176 vss 0.255f
C2063 out.n354 vss 0.139f
C2064 out.t122 vss 0.255f
C2065 out.n355 vss 0.139f
C2066 out.t411 vss 0.255f
C2067 out.n356 vss 0.139f
C2068 out.t315 vss 0.255f
C2069 out.n357 vss 0.139f
C2070 out.t261 vss 0.255f
C2071 out.n358 vss 0.139f
C2072 out.t403 vss 0.255f
C2073 out.n359 vss 0.139f
C2074 out.t350 vss 0.255f
C2075 out.n360 vss 0.139f
C2076 out.t296 vss 0.255f
C2077 out.n361 vss 0.139f
C2078 out.t202 vss 0.255f
C2079 out.n362 vss 0.139f
C2080 out.t149 vss 0.255f
C2081 out.n363 vss 0.139f
C2082 out.t93 vss 0.255f
C2083 out.n364 vss 0.139f
C2084 out.t381 vss 0.255f
C2085 out.n365 vss 0.139f
C2086 out.t327 vss 0.255f
C2087 out.n366 vss 0.139f
C2088 out.t231 vss 0.255f
C2089 out.n367 vss 0.139f
C2090 out.t179 vss 0.255f
C2091 out.n368 vss 0.139f
C2092 out.t125 vss 0.255f
C2093 out.n369 vss 0.139f
C2094 out.t410 vss 0.255f
C2095 out.n370 vss 0.139f
C2096 out.t289 vss 0.255f
C2097 out.n371 vss 0.139f
C2098 out.t195 vss 0.255f
C2099 out.n372 vss 0.139f
C2100 out.t139 vss 0.255f
C2101 out.n373 vss 0.139f
C2102 out.t88 vss 0.255f
C2103 out.n374 vss 0.139f
C2104 out.t374 vss 0.255f
C2105 out.n375 vss 0.139f
C2106 out.t318 vss 0.255f
C2107 out.n376 vss 0.139f
C2108 out.t225 vss 0.255f
C2109 out.n377 vss 0.139f
C2110 out.t171 vss 0.255f
C2111 out.n378 vss 0.139f
C2112 out.t118 vss 0.255f
C2113 out.n379 vss 0.139f
C2114 out.t406 vss 0.255f
C2115 out.n380 vss 0.139f
C2116 out.t352 vss 0.255f
C2117 out.n381 vss 0.139f
C2118 out.t257 vss 0.255f
C2119 out.n382 vss 0.139f
C2120 out.t229 vss 0.255f
C2121 out.n383 vss 0.106f
C2122 out.n384 vss 0.0513f
C2123 out.n385 vss 0.0498f
C2124 out.n386 vss 0.11f
C2125 out.n387 vss 0.0498f
C2126 out.n388 vss 0.11f
C2127 out.n389 vss 0.0498f
C2128 out.n390 vss 0.108f
C2129 out.n391 vss 0.0498f
C2130 out.n392 vss 0.112f
C2131 out.n393 vss 0.0498f
C2132 out.n394 vss 0.112f
C2133 out.n395 vss 0.0498f
C2134 out.n396 vss 0.107f
C2135 out.n397 vss 0.0498f
C2136 out.n398 vss 0.139f
C2137 out.n399 vss 0.139f
C2138 out.n400 vss 0.139f
C2139 out.n401 vss 0.139f
C2140 out.n402 vss 0.125f
C2141 out.n403 vss 0.0712f
C2142 out.n404 vss 0.0621f
C2143 out.n405 vss 0.124f
C2144 out.n406 vss 0.121f
C2145 out.n407 vss 0.235f
C2146 out.n408 vss 0.0149f
C2147 vin.t7 vss 0.0293f
C2148 vin.t51 vss 0.0323f
C2149 vin.t6 vss 0.0243f
C2150 vin.t2 vss 0.0243f
C2151 vin.n0 vss 0.171f
C2152 vin.t56 vss 0.0243f
C2153 vin.t58 vss 0.0243f
C2154 vin.n1 vss 0.171f
C2155 vin.t5 vss 0.0243f
C2156 vin.t9 vss 0.0243f
C2157 vin.n2 vss 0.171f
C2158 vin.t50 vss 0.0243f
C2159 vin.t59 vss 0.0243f
C2160 vin.n3 vss 0.171f
C2161 vin.t8 vss 0.0243f
C2162 vin.t0 vss 0.0243f
C2163 vin.n4 vss 0.171f
C2164 vin.t54 vss 0.0243f
C2165 vin.t55 vss 0.0243f
C2166 vin.n5 vss 0.171f
C2167 vin.t1 vss 0.0243f
C2168 vin.t4 vss 0.0243f
C2169 vin.n6 vss 0.171f
C2170 vin.t57 vss 0.0243f
C2171 vin.t53 vss 0.0243f
C2172 vin.n7 vss 0.171f
C2173 vin.t3 vss 0.0293f
C2174 vin.t52 vss 0.0323f
C2175 vin.n8 vss 0.489f
C2176 vin.n9 vss 0.143f
C2177 vin.n10 vss 0.143f
C2178 vin.n11 vss 0.143f
C2179 vin.n12 vss 0.144f
C2180 vin.n13 vss 0.508f
C2181 vin.t70 vss 0.0293f
C2182 vin.t38 vss 0.0323f
C2183 vin.t75 vss 0.0243f
C2184 vin.t77 vss 0.0243f
C2185 vin.n14 vss 0.171f
C2186 vin.t37 vss 0.0243f
C2187 vin.t31 vss 0.0243f
C2188 vin.n15 vss 0.171f
C2189 vin.t74 vss 0.0243f
C2190 vin.t78 vss 0.0243f
C2191 vin.n16 vss 0.171f
C2192 vin.t36 vss 0.0243f
C2193 vin.t30 vss 0.0243f
C2194 vin.n17 vss 0.171f
C2195 vin.t72 vss 0.0243f
C2196 vin.t73 vss 0.0243f
C2197 vin.n18 vss 0.171f
C2198 vin.t33 vss 0.0243f
C2199 vin.t35 vss 0.0243f
C2200 vin.n19 vss 0.171f
C2201 vin.t71 vss 0.0243f
C2202 vin.t76 vss 0.0243f
C2203 vin.n20 vss 0.171f
C2204 vin.t39 vss 0.0243f
C2205 vin.t34 vss 0.0243f
C2206 vin.n21 vss 0.171f
C2207 vin.t79 vss 0.0293f
C2208 vin.t32 vss 0.0323f
C2209 vin.n22 vss 0.489f
C2210 vin.n23 vss 0.143f
C2211 vin.n24 vss 0.143f
C2212 vin.n25 vss 0.143f
C2213 vin.n26 vss 0.144f
C2214 vin.n27 vss 0.509f
C2215 vin.n28 vss 0.0764f
C2216 vin.t14 vss 0.0293f
C2217 vin.t46 vss 0.0323f
C2218 vin.t11 vss 0.0243f
C2219 vin.t18 vss 0.0243f
C2220 vin.n29 vss 0.171f
C2221 vin.t42 vss 0.0243f
C2222 vin.t47 vss 0.0243f
C2223 vin.n30 vss 0.171f
C2224 vin.t17 vss 0.0243f
C2225 vin.t13 vss 0.0243f
C2226 vin.n31 vss 0.171f
C2227 vin.t41 vss 0.0243f
C2228 vin.t45 vss 0.0243f
C2229 vin.n32 vss 0.171f
C2230 vin.t16 vss 0.0243f
C2231 vin.t19 vss 0.0243f
C2232 vin.n33 vss 0.171f
C2233 vin.t40 vss 0.0243f
C2234 vin.t44 vss 0.0243f
C2235 vin.n34 vss 0.171f
C2236 vin.t12 vss 0.0243f
C2237 vin.t10 vss 0.0243f
C2238 vin.n35 vss 0.171f
C2239 vin.t43 vss 0.0243f
C2240 vin.t49 vss 0.0243f
C2241 vin.n36 vss 0.171f
C2242 vin.t15 vss 0.0293f
C2243 vin.t48 vss 0.0323f
C2244 vin.n37 vss 0.489f
C2245 vin.n38 vss 0.143f
C2246 vin.n39 vss 0.143f
C2247 vin.n40 vss 0.143f
C2248 vin.n41 vss 0.144f
C2249 vin.n42 vss 0.509f
C2250 vin.n43 vss 0.0766f
C2251 vin.t23 vss 0.0293f
C2252 vin.t69 vss 0.0323f
C2253 vin.t20 vss 0.0243f
C2254 vin.t29 vss 0.0243f
C2255 vin.n44 vss 0.171f
C2256 vin.t68 vss 0.0243f
C2257 vin.t65 vss 0.0243f
C2258 vin.n45 vss 0.171f
C2259 vin.t28 vss 0.0243f
C2260 vin.t22 vss 0.0243f
C2261 vin.n46 vss 0.171f
C2262 vin.t62 vss 0.0243f
C2263 vin.t64 vss 0.0243f
C2264 vin.n47 vss 0.171f
C2265 vin.t24 vss 0.0243f
C2266 vin.t27 vss 0.0243f
C2267 vin.n48 vss 0.171f
C2268 vin.t61 vss 0.0243f
C2269 vin.t67 vss 0.0243f
C2270 vin.n49 vss 0.171f
C2271 vin.t21 vss 0.0243f
C2272 vin.t26 vss 0.0243f
C2273 vin.n50 vss 0.171f
C2274 vin.t60 vss 0.0243f
C2275 vin.t63 vss 0.0243f
C2276 vin.n51 vss 0.171f
C2277 vin.t25 vss 0.0293f
C2278 vin.t66 vss 0.0323f
C2279 vin.n52 vss 0.489f
C2280 vin.n53 vss 0.143f
C2281 vin.n54 vss 0.143f
C2282 vin.n55 vss 0.143f
C2283 vin.n56 vss 0.144f
C2284 vin.n57 vss 0.509f
C2285 vin.n58 vss 0.08f
C2286 vin.n59 vss 0.807f
C2287 vin.n60 vss 0.764f
C2288 vin.n61 vss 1.01f
C2289 vin.n62 vss 0.31f
.ends

