magic
tech sky130B
magscale 1 2
timestamp 1696887389
<< locali >>
rect 14183 4004 19393 4064
rect 14196 3724 14230 4004
rect 14816 3837 14851 4004
rect 14816 3811 14849 3837
rect 15431 3787 15491 4004
rect 16061 3772 16121 4004
rect 16704 3773 16764 4004
rect 17344 3772 17404 4004
rect 17989 3772 18049 4004
rect 18607 3770 18667 4004
rect 19239 3772 19299 4004
rect 20161 3933 20202 4145
rect 13889 2847 13930 3646
rect 9354 2784 13941 2847
rect 9354 2720 9417 2784
rect 14505 2723 14542 3642
rect 15151 2776 15191 3648
rect 15784 2886 15831 3649
rect 16424 2980 16473 3645
rect 17070 3055 17105 3642
rect 17707 3127 17744 3643
rect 18333 3197 18367 3627
rect 18962 3269 18997 3641
rect 18962 3234 22295 3269
rect 18333 3163 22151 3197
rect 17707 3090 21999 3127
rect 17070 3020 21824 3055
rect 16422 2947 21047 2980
rect 16422 2928 20985 2947
rect 20169 2886 20235 2889
rect 15778 2831 20235 2886
rect 21789 2839 21824 3020
rect 21962 2845 21999 3090
rect 15778 2827 20166 2831
rect 15151 2736 17394 2776
rect 22117 2840 22151 3163
rect 22260 2841 22295 3234
rect 10242 2664 14553 2723
<< viali >>
rect 9347 2643 9424 2720
rect 10178 2661 10242 2725
rect 20985 2875 21057 2947
rect 17394 2731 17445 2782
rect 20166 2759 20238 2831
rect 21772 2770 21841 2839
rect 21946 2776 22015 2845
rect 22098 2768 22170 2840
rect 22241 2769 22313 2841
<< metal1 >>
rect 20132 5580 20221 5812
rect 20677 5617 20772 5815
rect 20132 5207 20221 5213
rect 20132 5126 20138 5207
rect 20215 5126 20221 5207
rect 20132 5120 20221 5126
rect 13713 4106 14242 4199
rect 20979 2947 21063 2959
rect 20979 2875 20985 2947
rect 21057 2875 21063 2947
rect 20160 2831 20244 2843
rect 17382 2782 17457 2788
rect 9341 2720 9430 2732
rect 17382 2731 17394 2782
rect 17445 2731 17457 2782
rect 9341 2643 9347 2720
rect 9424 2643 9430 2720
rect 10166 2725 10254 2731
rect 17382 2725 17457 2731
rect 20160 2759 20166 2831
rect 20238 2759 20244 2831
rect 10166 2661 10178 2725
rect 10242 2661 10254 2725
rect 17388 2713 17451 2725
rect 20160 2723 20244 2759
rect 20979 2753 21063 2875
rect 21766 2839 21847 2851
rect 21766 2770 21772 2839
rect 21841 2770 21847 2839
rect 21766 2758 21847 2770
rect 21940 2845 22021 2857
rect 21940 2776 21946 2845
rect 22015 2776 22021 2845
rect 21940 2764 22021 2776
rect 22092 2840 22176 2846
rect 22092 2768 22098 2840
rect 22170 2768 22176 2840
rect 22092 2762 22176 2768
rect 22235 2841 22319 2853
rect 22235 2769 22241 2841
rect 22313 2769 22319 2841
rect 22957 2784 23005 4422
rect 22235 2757 22319 2769
rect 10166 2655 10254 2661
rect 9341 2631 9430 2643
use carray  carray_0
timestamp 1696461989
transform 1 0 -4081 0 1 2059
box 62 -5400 27110 802
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1693170804
transform 0 1 14289 1 0 3562
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1693170804
transform 0 1 18741 1 0 3560
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_2
timestamp 1693170804
transform 0 1 18109 1 0 3562
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_3
timestamp 1693170804
transform 0 1 17489 1 0 3562
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_4
timestamp 1693170804
transform 0 1 16849 1 0 3562
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_5
timestamp 1693170804
transform 0 1 16209 1 0 3562
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_6
timestamp 1693170804
transform 0 1 15569 1 0 3562
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_7
timestamp 1693170804
transform 0 1 14929 1 0 3562
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_8
timestamp 1693170804
transform 0 1 13365 1 0 3732
box -38 -48 314 592
use sw_top  sw_top_0
timestamp 1696887389
transform 1 0 20949 0 -1 3885
box -817 -1844 2074 554
<< end >>
