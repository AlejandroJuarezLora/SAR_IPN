magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect 0 269 812 590
<< pwell >>
rect 39 29 773 191
<< scnmos >>
rect 117 55 695 165
<< scpmoshvt >>
rect 117 331 695 505
<< ndiff >>
rect 65 120 117 165
rect 65 86 73 120
rect 107 86 117 120
rect 65 55 117 86
rect 695 120 747 165
rect 695 86 705 120
rect 739 86 747 120
rect 695 55 747 86
<< pdiff >>
rect 65 493 117 505
rect 65 459 73 493
rect 107 459 117 493
rect 65 391 117 459
rect 65 357 73 391
rect 107 357 117 391
rect 65 331 117 357
rect 695 493 747 505
rect 695 459 705 493
rect 739 459 747 493
rect 695 391 747 459
rect 695 357 705 391
rect 739 357 747 391
rect 695 331 747 357
<< ndiffc >>
rect 73 86 107 120
rect 705 86 739 120
<< pdiffc >>
rect 73 459 107 493
rect 73 357 107 391
rect 705 459 739 493
rect 705 357 739 391
<< poly >>
rect 117 505 695 531
rect 117 305 695 331
rect 117 283 381 305
rect 117 249 133 283
rect 167 249 232 283
rect 266 249 331 283
rect 365 249 381 283
rect 117 233 381 249
rect 423 247 695 263
rect 423 213 439 247
rect 473 213 542 247
rect 576 213 645 247
rect 679 213 695 247
rect 423 191 695 213
rect 117 165 695 191
rect 117 29 695 55
<< polycont >>
rect 133 249 167 283
rect 232 249 266 283
rect 331 249 365 283
rect 439 213 473 247
rect 542 213 576 247
rect 645 213 679 247
<< locali >>
rect 38 535 67 569
rect 101 535 159 569
rect 193 535 251 569
rect 285 535 343 569
rect 377 535 435 569
rect 469 535 527 569
rect 561 535 619 569
rect 653 535 711 569
rect 745 535 774 569
rect 55 493 757 535
rect 55 459 73 493
rect 107 459 705 493
rect 739 459 757 493
rect 55 391 757 459
rect 55 357 73 391
rect 107 357 705 391
rect 739 357 757 391
rect 55 317 757 357
rect 55 249 133 283
rect 167 249 232 283
rect 266 249 331 283
rect 365 249 385 283
rect 55 179 385 249
rect 419 247 757 317
rect 419 213 439 247
rect 473 213 542 247
rect 576 213 645 247
rect 679 213 757 247
rect 55 120 757 179
rect 55 86 73 120
rect 107 86 705 120
rect 739 86 757 120
rect 55 25 757 86
rect 38 -9 67 25
rect 101 -9 159 25
rect 193 -9 251 25
rect 285 -9 343 25
rect 377 -9 435 25
rect 469 -9 527 25
rect 561 -9 619 25
rect 653 -9 711 25
rect 745 -9 774 25
<< viali >>
rect 67 535 101 569
rect 159 535 193 569
rect 251 535 285 569
rect 343 535 377 569
rect 435 535 469 569
rect 527 535 561 569
rect 619 535 653 569
rect 711 535 745 569
rect 67 -9 101 25
rect 159 -9 193 25
rect 251 -9 285 25
rect 343 -9 377 25
rect 435 -9 469 25
rect 527 -9 561 25
rect 619 -9 653 25
rect 711 -9 745 25
<< metal1 >>
rect 38 569 774 600
rect 38 535 67 569
rect 101 535 159 569
rect 193 535 251 569
rect 285 535 343 569
rect 377 535 435 569
rect 469 535 527 569
rect 561 535 619 569
rect 653 535 711 569
rect 745 535 774 569
rect 38 504 774 535
rect 38 25 774 56
rect 38 -9 67 25
rect 101 -9 159 25
rect 193 -9 251 25
rect 285 -9 343 25
rect 377 -9 435 25
rect 469 -9 527 25
rect 561 -9 619 25
rect 653 -9 711 25
rect 745 -9 774 25
rect 38 -40 774 -9
<< labels >>
rlabel comment s 38 8 38 8 4 decap_8
<< properties >>
string FIXED_BBOX 38 8 774 552
string path 0.950 0.200 19.350 0.200 
<< end >>
