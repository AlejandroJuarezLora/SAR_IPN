magic
tech sky130B
magscale 1 2
timestamp 1696109480
<< metal1 >>
rect 176 1185 182 1295
rect 292 1185 298 1295
rect 179 405 185 512
rect 292 405 298 512
<< via1 >>
rect 182 1185 292 1295
rect 185 405 292 512
<< metal2 >>
rect 182 1295 292 1301
rect 178 1190 182 1290
rect 292 1190 296 1290
rect 182 1179 292 1185
rect 185 512 292 518
rect 181 410 185 507
rect 292 410 296 507
rect 185 399 292 405
<< via2 >>
rect 187 1190 287 1290
rect 190 410 287 507
<< metal3 >>
rect 182 1294 292 1295
rect 177 1186 183 1294
rect 291 1186 297 1294
rect 182 1185 292 1186
rect 185 507 292 892
rect 185 410 190 507
rect 287 410 292 507
rect 185 405 292 410
<< via3 >>
rect 183 1290 291 1294
rect 183 1190 187 1290
rect 187 1190 287 1290
rect 287 1190 291 1290
rect 183 1186 291 1190
<< metal4 >>
rect 182 1294 292 1295
rect 182 1186 183 1294
rect 291 1186 292 1294
rect 182 836 292 1186
use sky130_fd_pr__cap_mim_m3_1  XC2
timestamp 1695772557
transform 1 0 386 0 1 840
box -386 -240 90 240
<< labels >>
flabel space 152 376 320 526 0 FreeSans 800 0 0 0 cn
port 0 nsew
flabel space 154 1166 318 1324 0 FreeSans 800 0 0 0 cp
port 1 nsew
<< end >>
