magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 958 542
<< pwell >>
rect 1 -19 919 163
rect 30 -57 64 -19
<< scnmos >>
rect 79 7 109 137
rect 163 7 193 137
rect 247 7 277 137
rect 331 7 361 137
rect 519 7 549 137
rect 609 7 639 137
rect 711 7 741 137
rect 811 7 841 137
<< scpmoshvt >>
rect 79 257 109 457
rect 163 257 193 457
rect 247 257 277 457
rect 331 257 361 457
rect 415 257 445 457
rect 609 257 639 457
rect 711 257 741 457
rect 811 257 841 457
<< ndiff >>
rect 27 125 79 137
rect 27 91 35 125
rect 69 91 79 125
rect 27 7 79 91
rect 109 53 163 137
rect 109 19 119 53
rect 153 19 163 53
rect 109 7 163 19
rect 193 125 247 137
rect 193 91 203 125
rect 237 91 247 125
rect 193 7 247 91
rect 277 53 331 137
rect 277 19 287 53
rect 321 19 331 53
rect 277 7 331 19
rect 361 125 413 137
rect 361 91 371 125
rect 405 91 413 125
rect 361 7 413 91
rect 467 125 519 137
rect 467 91 475 125
rect 509 91 519 125
rect 467 7 519 91
rect 549 53 609 137
rect 549 19 565 53
rect 599 19 609 53
rect 549 7 609 19
rect 639 129 711 137
rect 639 95 651 129
rect 685 95 711 129
rect 639 61 711 95
rect 639 27 651 61
rect 685 27 711 61
rect 639 7 711 27
rect 741 53 811 137
rect 741 19 751 53
rect 785 19 811 53
rect 741 7 811 19
rect 841 125 893 137
rect 841 91 851 125
rect 885 91 893 125
rect 841 53 893 91
rect 841 19 851 53
rect 885 19 893 53
rect 841 7 893 19
<< pdiff >>
rect 27 437 79 457
rect 27 403 35 437
rect 69 403 79 437
rect 27 367 79 403
rect 27 333 35 367
rect 69 333 79 367
rect 27 257 79 333
rect 109 419 163 457
rect 109 385 119 419
rect 153 385 163 419
rect 109 257 163 385
rect 193 437 247 457
rect 193 403 203 437
rect 237 403 247 437
rect 193 367 247 403
rect 193 333 203 367
rect 237 333 247 367
rect 193 257 247 333
rect 277 419 331 457
rect 277 385 287 419
rect 321 385 331 419
rect 277 257 331 385
rect 361 437 415 457
rect 361 403 371 437
rect 405 403 415 437
rect 361 367 415 403
rect 361 333 371 367
rect 405 333 415 367
rect 361 257 415 333
rect 445 419 609 457
rect 445 385 478 419
rect 512 385 546 419
rect 580 385 609 419
rect 445 257 609 385
rect 639 437 711 457
rect 639 403 667 437
rect 701 403 711 437
rect 639 367 711 403
rect 639 333 667 367
rect 701 333 711 367
rect 639 257 711 333
rect 741 383 811 457
rect 741 349 767 383
rect 801 349 811 383
rect 741 303 811 349
rect 741 269 767 303
rect 801 269 811 303
rect 741 257 811 269
rect 841 437 893 457
rect 841 403 851 437
rect 885 403 893 437
rect 841 369 893 403
rect 841 335 851 369
rect 885 335 893 369
rect 841 257 893 335
<< ndiffc >>
rect 35 91 69 125
rect 119 19 153 53
rect 203 91 237 125
rect 287 19 321 53
rect 371 91 405 125
rect 475 91 509 125
rect 565 19 599 53
rect 651 95 685 129
rect 651 27 685 61
rect 751 19 785 53
rect 851 91 885 125
rect 851 19 885 53
<< pdiffc >>
rect 35 403 69 437
rect 35 333 69 367
rect 119 385 153 419
rect 203 403 237 437
rect 203 333 237 367
rect 287 385 321 419
rect 371 403 405 437
rect 371 333 405 367
rect 478 385 512 419
rect 546 385 580 419
rect 667 403 701 437
rect 667 333 701 367
rect 767 349 801 383
rect 767 269 801 303
rect 851 403 885 437
rect 851 335 885 369
<< poly >>
rect 79 457 109 483
rect 163 457 193 483
rect 247 457 277 483
rect 331 457 361 483
rect 415 457 445 483
rect 609 457 639 483
rect 711 457 741 483
rect 811 457 841 483
rect 79 225 109 257
rect 163 225 193 257
rect 247 225 277 257
rect 331 225 361 257
rect 415 225 445 257
rect 609 225 639 257
rect 22 209 193 225
rect 22 175 32 209
rect 66 175 104 209
rect 138 175 193 209
rect 22 159 193 175
rect 235 209 361 225
rect 235 175 245 209
rect 279 175 317 209
rect 351 175 361 209
rect 235 159 361 175
rect 403 209 639 225
rect 403 175 413 209
rect 447 175 499 209
rect 533 175 581 209
rect 615 175 639 209
rect 403 159 639 175
rect 79 137 109 159
rect 163 137 193 159
rect 247 137 277 159
rect 331 137 361 159
rect 519 137 549 159
rect 609 137 639 159
rect 711 225 741 257
rect 811 225 841 257
rect 711 209 898 225
rect 711 175 780 209
rect 814 175 848 209
rect 882 175 898 209
rect 711 159 898 175
rect 711 137 741 159
rect 811 137 841 159
rect 79 -19 109 7
rect 163 -19 193 7
rect 247 -19 277 7
rect 331 -19 361 7
rect 519 -19 549 7
rect 609 -19 639 7
rect 711 -19 741 7
rect 811 -19 841 7
<< polycont >>
rect 32 175 66 209
rect 104 175 138 209
rect 245 175 279 209
rect 317 175 351 209
rect 413 175 447 209
rect 499 175 533 209
rect 581 175 615 209
rect 780 175 814 209
rect 848 175 882 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 920 521
rect 35 437 69 453
rect 35 367 69 403
rect 103 419 169 487
rect 103 385 119 419
rect 153 385 169 419
rect 203 437 237 453
rect 203 367 237 403
rect 271 419 337 487
rect 271 385 287 419
rect 321 385 337 419
rect 371 437 405 453
rect 69 333 203 351
rect 371 367 405 403
rect 462 419 596 487
rect 462 385 478 419
rect 512 385 546 419
rect 580 385 596 419
rect 667 437 885 453
rect 701 419 851 437
rect 237 333 371 351
rect 667 367 701 403
rect 405 333 667 351
rect 35 317 701 333
rect 751 349 767 383
rect 801 349 817 383
rect 751 303 817 349
rect 851 369 885 403
rect 851 319 885 335
rect 751 283 767 303
rect 29 209 164 283
rect 29 175 32 209
rect 66 175 104 209
rect 138 175 164 209
rect 29 159 164 175
rect 210 209 351 283
rect 210 175 245 209
rect 279 175 317 209
rect 210 159 351 175
rect 391 209 533 283
rect 651 269 767 283
rect 801 269 817 303
rect 651 249 817 269
rect 391 175 413 209
rect 447 175 499 209
rect 391 159 533 175
rect 581 209 615 225
rect 581 159 615 175
rect 651 129 714 249
rect 853 215 898 285
rect 764 209 898 215
rect 764 175 780 209
rect 814 175 848 209
rect 882 175 898 209
rect 19 91 35 125
rect 69 91 203 125
rect 237 91 371 125
rect 405 91 421 125
rect 459 91 475 125
rect 509 95 651 125
rect 685 125 714 129
rect 685 95 851 125
rect 509 91 851 95
rect 885 91 901 125
rect 651 61 685 91
rect 103 19 119 53
rect 153 19 169 53
rect 271 19 287 53
rect 321 19 565 53
rect 599 19 615 53
rect 835 53 901 91
rect 103 -23 169 19
rect 651 11 685 27
rect 735 19 751 53
rect 785 19 801 53
rect 835 19 851 53
rect 885 19 901 53
rect 735 -23 801 19
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 920 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 857 487 891 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
rect 857 -57 891 -23
<< metal1 >>
rect 0 521 920 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 920 521
rect 0 456 920 487
rect 0 -23 920 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 920 -23
rect 0 -88 920 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 a31oi_2
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 122 181 156 215 0 FreeSans 200 0 0 0 A3
port 11 nsew
flabel locali s 764 181 798 215 0 FreeSans 200 0 0 0 B1
port 7 nsew
flabel locali s 856 181 890 215 0 FreeSans 200 0 0 0 B1
port 7 nsew
flabel locali s 672 181 706 215 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel locali s 672 249 706 283 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel locali s 856 249 890 283 0 FreeSans 200 0 0 0 B1
port 7 nsew
flabel locali s 494 249 528 283 0 FreeSans 200 0 0 0 A1
port 9 nsew
flabel locali s 398 249 432 283 0 FreeSans 200 0 0 0 A1
port 9 nsew
flabel locali s 398 181 432 215 0 FreeSans 200 0 0 0 A1
port 9 nsew
flabel locali s 672 113 706 147 0 FreeSans 200 0 0 0 Y
port 8 nsew
flabel locali s 306 249 340 283 0 FreeSans 200 0 0 0 A2
port 10 nsew
flabel locali s 214 181 248 215 0 FreeSans 200 0 0 0 A2
port 10 nsew
flabel locali s 214 249 248 283 0 FreeSans 200 0 0 0 A2
port 10 nsew
flabel locali s 494 181 528 215 0 FreeSans 200 0 0 0 A1
port 9 nsew
flabel locali s 122 249 156 283 0 FreeSans 200 0 0 0 A3
port 11 nsew
flabel locali s 30 249 64 283 0 FreeSans 200 0 0 0 A3
port 11 nsew
flabel locali s 30 181 64 215 0 FreeSans 200 0 0 0 A3
port 11 nsew
flabel locali s 306 181 340 215 0 FreeSans 200 0 0 0 A2
port 10 nsew
<< properties >>
string FIXED_BBOX 0 -40 920 504
string path 0.000 12.600 23.000 12.600 
<< end >>
