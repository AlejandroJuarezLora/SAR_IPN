magic
tech sky130B
timestamp 1696364841
<< pwell >>
rect 4016 1132 4432 1175
rect 4016 935 4059 1132
rect 4389 935 4432 1132
rect 4016 892 4432 935
<< psubdiff >>
rect 4029 1145 4132 1162
rect 4149 1145 4166 1162
rect 4183 1145 4200 1162
rect 4217 1145 4234 1162
rect 4251 1145 4268 1162
rect 4285 1145 4302 1162
rect 4319 1145 4419 1162
rect 4029 1062 4046 1145
rect 4029 1028 4046 1045
rect 4029 922 4046 1011
rect 4402 1062 4419 1145
rect 4402 1028 4419 1045
rect 4402 922 4419 1011
rect 4029 905 4132 922
rect 4149 905 4166 922
rect 4183 905 4200 922
rect 4217 905 4234 922
rect 4251 905 4268 922
rect 4285 905 4302 922
rect 4319 905 4419 922
<< psubdiffcont >>
rect 4132 1145 4149 1162
rect 4166 1145 4183 1162
rect 4200 1145 4217 1162
rect 4234 1145 4251 1162
rect 4268 1145 4285 1162
rect 4302 1145 4319 1162
rect 4029 1045 4046 1062
rect 4029 1011 4046 1028
rect 4402 1045 4419 1062
rect 4402 1011 4419 1028
rect 4132 905 4149 922
rect 4166 905 4183 922
rect 4200 905 4217 922
rect 4234 905 4251 922
rect 4268 905 4285 922
rect 4302 905 4319 922
<< locali >>
rect 4029 1145 4132 1162
rect 4149 1145 4166 1162
rect 4183 1145 4200 1162
rect 4217 1145 4234 1162
rect 4251 1145 4268 1162
rect 4285 1145 4302 1162
rect 4319 1145 4419 1162
rect 4029 1062 4046 1145
rect 4029 1028 4046 1045
rect 4029 922 4046 1011
rect 4402 1062 4419 1145
rect 4402 1028 4419 1045
rect 4402 922 4419 1011
rect 4029 905 4132 922
rect 4149 905 4166 922
rect 4183 905 4200 922
rect 4217 905 4234 922
rect 4251 905 4268 922
rect 4285 905 4302 922
rect 4319 905 4419 922
<< properties >>
string path 40.290 11.535 44.105 11.535 44.105 9.135 40.375 9.135 40.375 11.535 
<< end >>
