magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect 0 269 352 590
<< pwell >>
rect 39 29 313 191
<< scnmos >>
rect 117 55 235 165
<< scpmoshvt >>
rect 117 331 235 505
<< ndiff >>
rect 65 122 117 165
rect 65 88 73 122
rect 107 88 117 122
rect 65 55 117 88
rect 235 122 287 165
rect 235 88 245 122
rect 279 88 287 122
rect 235 55 287 88
<< pdiff >>
rect 65 493 117 505
rect 65 459 73 493
rect 107 459 117 493
rect 65 398 117 459
rect 65 364 73 398
rect 107 364 117 398
rect 65 331 117 364
rect 235 493 287 505
rect 235 459 245 493
rect 279 459 287 493
rect 235 398 287 459
rect 235 364 245 398
rect 279 364 287 398
rect 235 331 287 364
<< ndiffc >>
rect 73 88 107 122
rect 245 88 279 122
<< pdiffc >>
rect 73 459 107 493
rect 73 364 107 398
rect 245 459 279 493
rect 245 364 279 398
<< poly >>
rect 117 505 235 531
rect 117 301 235 331
rect 117 299 155 301
rect 89 283 155 299
rect 89 249 105 283
rect 139 249 155 283
rect 89 233 155 249
rect 197 243 263 259
rect 197 209 213 243
rect 247 209 263 243
rect 197 193 263 209
rect 197 191 235 193
rect 117 165 235 191
rect 117 29 235 55
<< polycont >>
rect 105 249 139 283
rect 213 209 247 243
<< locali >>
rect 38 535 67 569
rect 101 535 159 569
rect 193 535 251 569
rect 285 535 314 569
rect 55 493 297 535
rect 55 459 73 493
rect 107 459 245 493
rect 279 459 297 493
rect 55 398 297 459
rect 55 364 73 398
rect 107 364 245 398
rect 279 364 297 398
rect 55 317 297 364
rect 55 249 105 283
rect 139 249 159 283
rect 55 175 159 249
rect 193 243 297 317
rect 193 209 213 243
rect 247 209 297 243
rect 55 122 297 175
rect 55 88 73 122
rect 107 88 245 122
rect 279 88 297 122
rect 55 25 297 88
rect 38 -9 67 25
rect 101 -9 159 25
rect 193 -9 251 25
rect 285 -9 314 25
<< viali >>
rect 67 535 101 569
rect 159 535 193 569
rect 251 535 285 569
rect 67 -9 101 25
rect 159 -9 193 25
rect 251 -9 285 25
<< metal1 >>
rect 38 569 314 600
rect 38 535 67 569
rect 101 535 159 569
rect 193 535 251 569
rect 285 535 314 569
rect 38 504 314 535
rect 38 25 314 56
rect 38 -9 67 25
rect 101 -9 159 25
rect 193 -9 251 25
rect 285 -9 314 25
rect 38 -40 314 -9
<< labels >>
rlabel comment s 38 8 38 8 4 decap_3
<< properties >>
string FIXED_BBOX 38 8 314 552
string path 0.950 0.200 7.850 0.200 
<< end >>
