* SPICE3 file created from comp_temp.ext - technology: sky130B

.subckt comparator vn clk trim0 trim1 trim3 trimb0 trimb1 vp outp outn trim2 trimb4
+ trimb3 vdd trim4 trimb2 vss
X0 vdd.t4 clk.t0 outp.t2 sky130_fd_pr__pfet_01v8_2.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X1 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t4 trim3.t0 vss.t19 vss.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X2 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D trim2.t0 vss.t15 vss.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X3 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t1 IN.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 IN.t11 trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X5 diff clk.t1 vss.t23 vss.t22 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X6 trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D trim0.t0 vss.t1 vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X7 IP.t10 trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X8 vss.t5 trimb3.t0 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t4 vss.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X9 IN.t12 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t1 IP.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 vss.t25 trim4.t0 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t0 vss.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X12 IP.t11 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t2 IN.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t3 IN.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X15 IP.t9 vp.t0 diff vss.t26 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X16 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t0 trimb4.t0 vss.t12 vss.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X17 vss.t7 trimb1.t0 trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X18 vdd.t2 clk.t2 IN.t9 sky130_fd_pr__pfet_01v8_4.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X19 vdd.t5 outp.t3 outn.t1 sky130_fd_pr__pfet_01v8_1.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X20 IN.t13 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t4 IN.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 IP.t12 trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X23 outn.t2 outp.t4 IN.t10 vss.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X24 IP.t13 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t2 IP.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 IP.t14 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 vss.t17 trimb2.t0 trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D vss.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X28 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t5 IN.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X29 IN.t14 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t3 IP.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t4 IP.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t6 IN.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 IP.t15 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 IP.t16 trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t5 IP.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 IN.t15 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D trim1.t0 vss.t3 vss.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X38 vss.t9 trimb0.t0 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D vss.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X39 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t6 IP.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 outp.t0 outn.t3 IP vss.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X41 diff clk.t3 vss.t21 vss.t20 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X42 IN.t16 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 IP.t17 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t7 IN.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 IN.t17 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 vdd.t0 outn.t4 outp.t1 sky130_fd_pr__pfet_01v8_0.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X47 IN.t8 vn.t0 diff vss.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X48 IN.t18 trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X49 vdd.t3 clk.t4 outn.t0 sky130_fd_pr__pfet_01v8_3.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X50 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t8 IN.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t7 IP.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 vdd.t1 clk.t5 IP.t8 sky130_fd_pr__pfet_01v8_5.B sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.3
X53 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t8 IP.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 clk clk.t2 142.674
R1 clk clk.t4 142.674
R2 clk clk.t5 142.674
R3 clk.n1 clk.t0 138.101
R4 clk.n14 clk.t3 135.446
R5 clk.n9 clk.t1 135.445
R6 clk.n2 clk.n1 9.37697
R7 clk.n3 clk.n0 9.06819
R8 clk.n12 clk 9.0005
R9 clk.n5 clk 4.22973
R10 clk.n13 clk.n7 1.31023
R11 clk.n7 clk.n4 1.1896
R12 clk.n7 clk.n6 1.05722
R13 clk.n4 clk 0.666671
R14 clk.n6 clk.n5 0.63735
R15 clk.n14 clk.n13 0.391763
R16 clk.n13 clk.n12 0.217838
R17 clk clk.n14 0.06197
R18 clk clk.n11 0.0378839
R19 clk.n3 clk.n2 0.0320091
R20 clk.n6 clk 0.0187196
R21 clk.n11 clk.n10 0.0143459
R22 clk clk.n0 0.0112152
R23 clk.n5 clk 0.00793321
R24 clk.n12 clk.n8 0.00630322
R25 clk.n12 clk.n10 0.00285497
R26 clk.n2 clk 0.00258333
R27 clk.n10 clk.n9 0.00223611
R28 clk.n4 clk.n3 0.0016242
R29 outp outp.t3 142.75
R30 outp outp.t4 135.556
R31 outp.n0 outp.t1 28.5716
R32 outp.n6 outp.t2 28.5716
R33 outp.n2 outp.t0 17.4065
R34 outp.n3 outp.n1 12.1416
R35 outp.n5 outp 11.9327
R36 outp.n6 outp.n5 2.48232
R37 outp.n1 outp 1.96671
R38 outp.n1 outp 1.67658
R39 outp.n5 outp.n4 1.40229
R40 outp.n4 outp.n0 0.925267
R41 outp.n3 outp.n2 0.87748
R42 outp.n2 outp 0.223326
R43 outp.n4 outp.n3 0.1255
R44 outp.n0 outp 0.00593478
R45 outp outp.n6 0.00126219
R46 vdd vdd.t2 28.5765
R47 vdd vdd.t3 28.5764
R48 vdd vdd.t5 28.5764
R49 vdd vdd.t0 28.5764
R50 vdd vdd.t4 28.5764
R51 vdd vdd.t1 28.5764
R52 vdd vdd.n4 4.65558
R53 vdd.n0 vdd 4.63326
R54 vdd.n1 vdd.n0 3.42461
R55 vdd.n4 vdd.n3 3.3755
R56 vdd.n3 vdd.n2 2.5005
R57 vdd.n2 vdd.n1 2.01389
R58 vdd.n3 vdd 1.03505
R59 vdd.n4 vdd 1.03505
R60 vdd.n0 vdd 0.999332
R61 vdd.n1 vdd 0.999332
R62 vdd.n2 vdd 0.304071
R63 trim3.n0 trim3.t0 135.52
R64 trim3 trim3.n0 14.5581
R65 trim3.n1 trim3 0.143357
R66 trim3.n0 trim3 0.0588333
R67 trim3 trim3.n1 0.0551875
R68 trim3.n1 trim3 0.0551875
R69 vss.n16 vss 563.201
R70 vss.n17 vss.n16 299.421
R71 vss.n16 vss 231.439
R72 vss.n16 vss 187.733
R73 vss.n17 vss.n13 127.248
R74 vss.n35 vss.t24 116.466
R75 vss.n42 vss.t18 116.466
R76 vss.n32 vss.t14 116.466
R77 vss.n27 vss.t2 116.466
R78 vss.n22 vss.t0 116.466
R79 vss.n14 vss.n1 98.2576
R80 vss.n52 vss.n51 89.9979
R81 vss.n23 vss.n20 89.9979
R82 vss.n41 vss.n19 89.6005
R83 vss.n33 vss.n30 89.6005
R84 vss.n28 vss.n25 87.3417
R85 vss.n18 vss.n17 85.4593
R86 vss.n43 vss.t26 83.5656
R87 vss.n10 vss.n9 67.3887
R88 vss.n45 vss.n44 67.3887
R89 vss.n4 vss.n3 67.0332
R90 vss.n37 vss.n36 67.0332
R91 vss.n7 vss.n6 66.6358
R92 vss.n47 vss 57.2449
R93 vss.n50 vss.t27 55.2719
R94 vss.n56 vss.n8 46.3089
R95 vss.n57 vss.n5 46.3084
R96 vss.n55 vss.n11 44.1615
R97 vss.n51 vss 34.2593
R98 vss vss.n33 34.2593
R99 vss vss.n28 34.2593
R100 vss vss.n23 34.2593
R101 vss.n49 vss 28.2358
R102 vss.n48 vss 28.2358
R103 vss.n12 vss 28.2358
R104 vss.n18 vss 27.4829
R105 vss.n47 vss.n46 26.3534
R106 vss.n41 vss.n40 26.3534
R107 vss.n36 vss.n35 23.1984
R108 vss.n5 vss.n4 22.9652
R109 vss.n11 vss.n10 22.2123
R110 vss.n46 vss.n45 22.2123
R111 vss.n8 vss.n7 20.7064
R112 vss.n54 vss.n47 18.9589
R113 vss.n0 vss.t21 17.4428
R114 vss.n62 vss.t23 17.4102
R115 vss.n6 vss.t3 17.4063
R116 vss.n9 vss.t15 17.4063
R117 vss.n44 vss.t19 17.4063
R118 vss.n52 vss.t25 17.4063
R119 vss.n3 vss.t1 17.4063
R120 vss.n19 vss.t5 17.4063
R121 vss.n30 vss.t17 17.4063
R122 vss.n25 vss.t7 17.4063
R123 vss.n20 vss.t9 17.4063
R124 vss.n37 vss.t12 17.4063
R125 vss.n7 vss 13.5534
R126 vss.n61 vss.n60 12.4338
R127 vss.n29 vss 12.0501
R128 vss.n24 vss 12.0501
R129 vss.n10 vss 12.0476
R130 vss.n45 vss 12.0476
R131 vss.t24 vss.t11 11.8444
R132 vss.n43 vss.n42 11.8444
R133 vss.t18 vss.t4 11.8444
R134 vss.n32 vss.n31 11.8444
R135 vss.t14 vss.t16 11.8444
R136 vss.n27 vss.n26 11.8444
R137 vss.t2 vss.t6 11.8444
R138 vss.n22 vss.n21 11.8444
R139 vss.t0 vss.t8 11.8444
R140 vss vss.n39 11.4922
R141 vss.n4 vss 11.2946
R142 vss.n36 vss 11.2946
R143 vss.n34 vss 9.90264
R144 vss.n60 vss.n2 8.58383
R145 vss.n40 vss 7.90638
R146 vss.n55 vss.n54 7.6021
R147 vss.n39 vss.n34 7.6021
R148 vss.n40 vss 7.46717
R149 vss.n58 vss.n57 6.90727
R150 vss.n39 vss.n38 6.87685
R151 vss.n54 vss.n53 6.87685
R152 vss.n24 vss.n2 6.87163
R153 vss.n59 vss.n58 6.59633
R154 vss vss.n15 6.14104
R155 vss.n56 vss.n55 3.87142
R156 vss.n34 vss.n29 3.87142
R157 vss.t26 vss.t10 3.29047
R158 vss.t27 vss.t13 2.63247
R159 vss.n29 vss.n24 2.40865
R160 vss.n57 vss.n56 2.40717
R161 vss.n1 vss.n0 1.80424
R162 vss.n62 vss.n61 1.01843
R163 vss.n61 vss.n1 0.800069
R164 vss.n59 vss 0.429667
R165 vss.n15 vss.n14 0.346446
R166 vss.t13 vss.n48 0.233661
R167 vss.t27 vss.n49 0.233661
R168 vss.t26 vss.n18 0.233661
R169 vss.n42 vss.n41 0.233661
R170 vss.n33 vss.n32 0.233661
R171 vss.n28 vss.n27 0.233661
R172 vss.n23 vss.n22 0.233661
R173 vss.n21 vss.n5 0.233661
R174 vss.n26 vss.n8 0.233661
R175 vss.n31 vss.n11 0.233661
R176 vss.n46 vss.n43 0.233661
R177 vss.n51 vss.n50 0.233661
R178 vss.t10 vss.n12 0.233661
R179 vss.n14 vss.t20 0.233661
R180 vss.n15 vss.t22 0.233661
R181 vss.n6 vss 0.201423
R182 vss.n9 vss 0.201423
R183 vss.n44 vss 0.201423
R184 vss.n3 vss 0.201423
R185 vss.n19 vss 0.201423
R186 vss.n30 vss 0.201423
R187 vss.n25 vss 0.201423
R188 vss.n20 vss 0.201423
R189 vss.n53 vss 0.19887
R190 vss.n38 vss 0.19887
R191 vss vss.n62 0.17713
R192 vss.n0 vss 0.144522
R193 vss.n2 vss 0.0688594
R194 vss.n58 vss 0.0337031
R195 vss.n60 vss.n59 0.0171667
R196 vss.n53 vss.n52 0.00305354
R197 vss.n38 vss.n37 0.00305354
R198 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t4 17.4065
R199 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t3 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t1 1.43874
R200 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t0 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t2 1.4117
R201 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.n0 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t0 0.839436
R202 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.n0 0.774957
R203 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.n0 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D.t3 0.517943
R204 trim2 trim2.t0 135.587
R205 trim2.n0 trim2 0.143357
R206 trim2.n0 trim2 0.0551875
R207 trim2 trim2.n0 0.047375
R208 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t0 17.4065
R209 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t7 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t3 2.24615
R210 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t6 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t1 2.17052
R211 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t4 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t7 2.13604
R212 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t1 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t4 2.11449
R213 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t2 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t5 2.10156
R214 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t5 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t6 2.06707
R215 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.n0 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t8 1.05221
R216 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.n0 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.t2 1.00578
R217 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D.n0 0.815415
R218 IN IN.t9 28.5716
R219 IN IN.t8 17.556
R220 IN IN.t10 17.4323
R221 IN.n1 IN.t15 6.43651
R222 IN IN.n1 4.86211
R223 IN.t1 IN.t5 2.28931
R224 IN.t2 IN.n2 2.2568
R225 IN.t4 IN.t1 2.22109
R226 IN.t16 IN.t14 2.21178
R227 IN.n2 IN.t4 2.19877
R228 IN.t6 IN.t3 2.18538
R229 IN.t13 IN.t12 2.17606
R230 IN.t0 IN.t6 2.16752
R231 IN.t18 IN.t11 2.15937
R232 IN.t3 IN.t2 2.14966
R233 IN.t14 IN.t13 2.13833
R234 IN.t12 IN.t17 2.13142
R235 IN.t17 IN.t18 2.07368
R236 IN.n0 IN 1.36688
R237 IN.n0 IN.t16 1.18651
R238 IN.n1 IN 1.08946
R239 IN.t15 IN.n0 0.887375
R240 IN IN.t0 0.830136
R241 IN.n2 IN.t7 0.14958
R242 trim0.n0 trim0.t0 135.528
R243 trim0 trim0.n0 0.883312
R244 trim0.n1 trim0 0.143357
R245 trim0.n0 trim0 0.0597105
R246 trim0 trim0.n1 0.0551875
R247 trim0.n1 trim0 0.0551875
R248 IP IP.t8 28.5716
R249 IP IP.t9 17.4065
R250 IP.n0 IP.t6 6.12031
R251 IP IP.n0 5.21925
R252 IP.t5 IP.t3 2.28887
R253 IP.t1 IP.t2 2.2568
R254 IP.t4 IP.t5 2.22109
R255 IP.t15 IP.t17 2.21178
R256 IP.t2 IP.t4 2.19877
R257 IP.t7 IP.t0 2.18538
R258 IP.t13 IP.t10 2.17606
R259 IP.t6 IP.t7 2.16752
R260 IP.t12 IP.t14 2.15837
R261 IP.t0 IP.t1 2.14966
R262 IP.t17 IP.t13 2.13833
R263 IP.t10 IP.t16 2.13142
R264 IP.t16 IP.t12 2.07368
R265 IP IP.n1 1.91429
R266 IP.n1 IP.t15 1.20437
R267 IP.n0 IP 1.1341
R268 IP.n1 IP.t11 0.869517
R269 IP.t11 IP 0.789188
R270 trimb3.n0 trimb3.t0 135.52
R271 trimb3 trimb3.n0 14.6093
R272 trimb3.n1 trimb3 1.7505
R273 trimb3.n1 trimb3 0.147821
R274 trimb3.n0 trimb3 0.0662895
R275 trimb3 trimb3.n1 0.0551875
R276 trimb3.n1 trimb3 0.0239375
R277 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t4 17.4065
R278 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t1 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t3 1.4383
R279 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t0 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t2 1.41126
R280 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.n0 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t0 0.839436
R281 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.n0 0.774957
R282 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.n0 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D.t1 0.517943
R283 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t0 17.4065
R284 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t4 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t5 2.24515
R285 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t7 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t6 2.17052
R286 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t1 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t4 2.13604
R287 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t6 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t1 2.11449
R288 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t8 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t3 2.10156
R289 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t3 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t7 2.06707
R290 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.n0 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t2 1.05121
R291 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.n0 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.t8 1.00578
R292 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D.n0 0.811943
R293 trim4 trim4.t0 135.587
R294 trim4.n0 trim4 1.7505
R295 trim4.n0 trim4 0.147821
R296 trim4 trim4.n0 0.0551875
R297 trim4.n0 trim4 0.047375
R298 vp vp.t0 135.585
R299 vp.n1 vp 21.551
R300 vp.n1 vp.n0 4.563
R301 vp vp.n1 0.063
R302 trimb4.n0 trimb4.t0 135.52
R303 trimb4 trimb4.n0 16.1639
R304 trimb4.n1 trimb4 0.143357
R305 trimb4.n0 trimb4 0.0662895
R306 trimb4.n1 trimb4 0.0551875
R307 trimb4 trimb4.n1 0.016125
R308 trimb1.n0 trimb1.t0 135.52
R309 trimb1 trimb1.n0 3.6366
R310 trimb1.n1 trimb1 1.7505
R311 trimb1.n1 trimb1 0.147821
R312 trimb1.n0 trimb1 0.0662895
R313 trimb1 trimb1.n1 0.0551875
R314 trimb1.n1 trimb1 0.016125
R315 outn outn.t4 142.75
R316 outn outn.t3 135.583
R317 outn.n3 outn.t0 28.5716
R318 outn.n1 outn.t1 28.5716
R319 outn.n6 outn.t2 17.5179
R320 outn.n4 outn 11.9171
R321 outn.n2 outn.n0 11.5801
R322 outn.n0 outn 2.30064
R323 outn.n4 outn.n3 2.19828
R324 outn.n0 outn 1.96165
R325 outn.n5 outn.n4 1.56914
R326 outn.n6 outn.n5 1.11657
R327 outn.n2 outn.n1 0.75805
R328 outn outn.n6 0.111913
R329 outn.n5 outn.n2 0.0228214
R330 outn.n1 outn 0.00593478
R331 outn.n3 outn 0.00126219
R332 trimb2.n0 trimb2.t0 135.52
R333 trimb2 trimb2.n0 7.55066
R334 trimb2.n1 trimb2 1.7505
R335 trimb2.n1 trimb2 0.147821
R336 trimb2.n0 trimb2 0.0662895
R337 trimb2 trimb2.n1 0.0551875
R338 trimb2.n1 trimb2 0.016125
R339 trim1 trim1.t0 135.587
R340 trim1.n0 trim1 1.7505
R341 trim1.n0 trim1 0.147821
R342 trim1 trim1.n0 0.0551875
R343 trim1.n0 trim1 0.047375
R344 trimb0.n0 trimb0.t0 135.52
R345 trimb0 trimb0.n0 0.889891
R346 trimb0.n1 trimb0 0.143357
R347 trimb0.n0 trimb0 0.0662895
R348 trimb0.n1 trimb0 0.0551875
R349 trimb0 trimb0.n1 0.047375
R350 vn.n0 vn.t0 135.524
R351 vn.n2 vn.n0 20.9926
R352 vn.n2 vn.n1 4.563
R353 vn vn.n2 0.063
R354 vn.n0 vn 0.0609167
C0 vp sky130_fd_pr__pfet_01v8_0.B 4.75e-19
C1 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D 2.52f
C2 diff trim3 1.63e-20
C3 IP vp 0.403f
C4 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D vp 0.00303f
C5 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D trimb3 0.084f
C6 trimb0 trimb2 6.91e-19
C7 vp trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D 9.83e-19
C8 vp trimb3 2.49e-20
C9 trim0 trim4 3.47e-19
C10 trim1 trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D 0.00763f
C11 sky130_fd_pr__pfet_01v8_5.B outp 0.0109f
C12 clk outp 0.195f
C13 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D 0.0266f
C14 vn trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D 0.00697f
C15 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D trimb2 0.0106f
C16 sky130_fd_pr__pfet_01v8_5.B vdd 0.0991f
C17 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D vp 5.11e-19
C18 trim0 IN 0.00459f
C19 clk vdd 0.261f
C20 sky130_fd_pr__pfet_01v8_5.B sky130_fd_pr__pfet_01v8_0.B 3.52e-20
C21 clk sky130_fd_pr__pfet_01v8_0.B 0.0404f
C22 IP sky130_fd_pr__pfet_01v8_5.B 0.0928f
C23 vn outp 0.00223f
C24 vp trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D 0.00677f
C25 IP clk 0.108f
C26 sky130_fd_pr__pfet_01v8_5.B trimb3 2.83e-19
C27 trim4 trim3 1.96f
C28 vn vdd 2.83e-20
C29 clk trimb3 0.0013f
C30 trim2 trim4 3.38e-19
C31 outn sky130_fd_pr__pfet_01v8_1.B 0.123f
C32 trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D trim3 0.00112f
C33 IP vn 0.00193f
C34 trim3 IN 0.0362f
C35 trimb1 trimb4 3.47e-19
C36 sky130_fd_pr__pfet_01v8_3.B clk 0.156f
C37 trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D trim2 0.00594f
C38 sky130_fd_pr__pfet_01v8_5.B trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D 2.63e-21
C39 trim2 IN 0.0256f
C40 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D clk 0.0216f
C41 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D clk 0.175f
C42 sky130_fd_pr__pfet_01v8_4.B vdd 0.0952f
C43 vp clk 0.0398f
C44 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D trim3 0.084f
C45 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D vn 0.00375f
C46 trim1 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D 0.00694f
C47 trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D trimb2 0.0431f
C48 vn trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D 6.06e-21
C49 diff outn 0.0167f
C50 trim0 trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D 0.0175f
C51 vn vp 0.0219f
C52 trimb1 trimb0 0.1f
C53 sky130_fd_pr__pfet_01v8_2.B outn 0.00136f
C54 IP trimb2 0.0256f
C55 IN sky130_fd_pr__pfet_01v8_1.B 3.5e-20
C56 sky130_fd_pr__pfet_01v8_5.B clk 0.149f
C57 trimb1 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D 0.00694f
C58 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D trimb2 0.0014f
C59 sky130_fd_pr__pfet_01v8_3.B sky130_fd_pr__pfet_01v8_4.B 0.00281f
C60 trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D trimb2 0.00594f
C61 trimb2 trimb3 0.835f
C62 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D sky130_fd_pr__pfet_01v8_4.B 0.00457f
C63 trim3 trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D 0.00115f
C64 vn clk 0.028f
C65 trim2 trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D 0.0014f
C66 trim1 vn 0.00133f
C67 diff IN 0.101f
C68 vp trimb2 2.01e-20
C69 trim3 vdd 1.73e-20
C70 IN outn 0.391f
C71 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D trim0 0.00404f
C72 clk sky130_fd_pr__pfet_01v8_4.B 0.165f
C73 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D diff 0.0031f
C74 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D outn 0.00822f
C75 trimb0 trimb4 3.47e-19
C76 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D trim3 0.0222f
C77 trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D trim4 9.87e-19
C78 trim4 IN 0.0398f
C79 sky130_fd_pr__pfet_01v8_1.B outp 0.168f
C80 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D trimb4 1.21f
C81 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D trim2 0.0431f
C82 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D trim3 0.0258f
C83 IP trimb1 0.0187f
C84 sky130_fd_pr__pfet_01v8_1.B vdd 0.118f
C85 trimb1 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D 0.00763f
C86 trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D IN 0.601f
C87 trimb1 trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D 0.0172f
C88 trimb1 trimb3 4.63e-19
C89 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D trim2 0.0106f
C90 sky130_fd_pr__pfet_01v8_1.B sky130_fd_pr__pfet_01v8_0.B 8.91e-19
C91 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D trim4 0.0328f
C92 trim1 trim0 0.102f
C93 vn trim0 0.00391f
C94 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D IN 2.52f
C95 diff outp 0.0134f
C96 trimb0 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D 0.00404f
C97 outn outp 0.469f
C98 trimb1 vp 2e-20
C99 sky130_fd_pr__pfet_01v8_3.B sky130_fd_pr__pfet_01v8_1.B 0.0133f
C100 diff vdd 0.00601f
C101 trim3 clk 0.0014f
C102 sky130_fd_pr__pfet_01v8_2.B outp 0.0994f
C103 outn vdd 0.354f
C104 trim1 trim3 4.63e-19
C105 IP diff 0.0997f
C106 outn sky130_fd_pr__pfet_01v8_0.B 0.166f
C107 sky130_fd_pr__pfet_01v8_2.B vdd 0.13f
C108 trim4 trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D 0.00101f
C109 IP outn 0.0272f
C110 vn trim3 2.88e-20
C111 diff trimb3 1.55e-22
C112 sky130_fd_pr__pfet_01v8_2.B sky130_fd_pr__pfet_01v8_0.B 0.0133f
C113 trim1 trim2 0.366f
C114 trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D trimb4 0.00203f
C115 IP sky130_fd_pr__pfet_01v8_2.B 0.0388f
C116 vn trim2 4.13e-20
C117 trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D 0.254f
C118 trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D IN 0.575f
C119 IP trimb4 0.0395f
C120 trim4 vdd 4.01e-20
C121 sky130_fd_pr__pfet_01v8_3.B outn 0.103f
C122 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D trimb4 0.00101f
C123 diff trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D 0.00242f
C124 trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D trimb4 9.87e-19
C125 trim3 sky130_fd_pr__pfet_01v8_4.B 3.06e-19
C126 clk sky130_fd_pr__pfet_01v8_1.B 0.0413f
C127 trimb4 trimb3 1.96f
C128 IN outp 0.0292f
C129 vp diff 0.0941f
C130 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D outn 9.15e-19
C131 vp outn 0.00191f
C132 IN vdd 0.136f
C133 sky130_fd_pr__pfet_01v8_2.B trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D 0.0104f
C134 vn sky130_fd_pr__pfet_01v8_1.B 4.18e-19
C135 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D outp 0.00116f
C136 IP IN 0.0261f
C137 trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D 0.0266f
C138 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D trimb4 0.0328f
C139 IP trimb0 0.00459f
C140 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D trim4 0.00203f
C141 vp trimb4 1.01e-20
C142 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D vdd 6.95e-20
C143 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D trimb0 0.0175f
C144 trimb0 trimb3 4.63e-19
C145 diff clk 0.115f
C146 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D trim4 1.21f
C147 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D 4.97f
C148 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D 0.236f
C149 trim0 trim3 4.63e-19
C150 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D IN 1.22f
C151 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D 0.0161f
C152 clk outn 0.195f
C153 trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D 0.0162f
C154 sky130_fd_pr__pfet_01v8_5.B sky130_fd_pr__pfet_01v8_2.B 0.00281f
C155 sky130_fd_pr__pfet_01v8_3.B IN 0.0368f
C156 trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D trimb3 0.0258f
C157 sky130_fd_pr__pfet_01v8_1.B sky130_fd_pr__pfet_01v8_4.B 3.52e-20
C158 sky130_fd_pr__pfet_01v8_2.B clk 0.155f
C159 trim2 trim0 6.91e-19
C160 trimb1 trimb2 0.363f
C161 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D 0.0162f
C162 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D IN 4.97f
C163 vn diff 0.102f
C164 trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D vp 2.6e-19
C165 vp IN 0.00462f
C166 sky130_fd_pr__pfet_01v8_5.B trimb4 5.34e-19
C167 vn outn 6.16e-19
C168 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D 0.232f
C169 clk trimb4 0.00429f
C170 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D sky130_fd_pr__pfet_01v8_3.B 0.0142f
C171 vp trimb0 5.71e-20
C172 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D 0.0818f
C173 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D 0.0818f
C174 vp trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D 4.12e-19
C175 trim4 clk 0.00314f
C176 trim2 trim3 0.839f
C177 trim1 trim4 3.47e-19
C178 outp vdd 0.339f
C179 outn sky130_fd_pr__pfet_01v8_4.B 0.0118f
C180 clk IN 0.182f
C181 sky130_fd_pr__pfet_01v8_0.B outp 0.119f
C182 IP outp 0.359f
C183 trim1 trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D 0.0172f
C184 trim1 IN 0.0187f
C185 sky130_fd_pr__pfet_01v8_0.B vdd 0.121f
C186 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D 1.22f
C187 trim_1.sky130_fd_pr__nfet_01v8_lvt_0.D trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D 0.00134f
C188 vn trim_1.sky130_fd_pr__nfet_01v8_lvt_3.D 0.00195f
C189 IP vdd 0.136f
C190 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D 0.00134f
C191 clk trim_0.sky130_fd_pr__nfet_01v8_lvt_2.D 5.12e-19
C192 vn IN 0.711f
C193 trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D clk 0.194f
C194 trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D 0.236f
C195 trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D trimb3 0.0222f
C196 IP sky130_fd_pr__pfet_01v8_0.B 7.44e-19
C197 trim_1.sky130_fd_pr__nfet_01v8_lvt_2.D trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D 0.0161f
C198 trimb3 vdd 1.16e-20
C199 vp trim_1.sky130_fd_pr__nfet_01v8_lvt_1.D 3.91e-19
C200 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D 0.575f
C201 trim4 sky130_fd_pr__pfet_01v8_4.B 9.49e-19
C202 sky130_fd_pr__pfet_01v8_3.B outp 0.00119f
C203 IP trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D 0.601f
C204 IP trimb3 0.0362f
C205 trimb2 trimb4 3.38e-19
C206 vn trim_1.sky130_fd_pr__nfet_01v8_lvt_4.D 0.00752f
C207 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D 0.254f
C208 trim_0.sky130_fd_pr__nfet_01v8_lvt_1.D trimb3 0.00115f
C209 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D outp 0.00758f
C210 sky130_fd_pr__pfet_01v8_3.B vdd 0.127f
C211 trim_0.sky130_fd_pr__nfet_01v8_lvt_3.D trimb3 0.00112f
C212 vp outp 0.00127f
C213 IN sky130_fd_pr__pfet_01v8_4.B 0.0939f
C214 trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D 0.232f
C215 trim_0.sky130_fd_pr__nfet_01v8_lvt_4.D vdd 6.67e-20
C216 vp trim_0.sky130_fd_pr__nfet_01v8_lvt_0.D 0.0019f
C217 vp vdd 3.04e-20
.ends

