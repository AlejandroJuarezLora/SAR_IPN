magic
tech sky130B
magscale 1 2
timestamp 1696271643
<< metal1 >>
rect -390 920 -266 1036
rect -348 -52 -318 174
rect -204 -152 -146 -92
rect -372 -196 -286 -168
use sky130_fd_pr__nfet_01v8_lvt_E33R59  sky130_fd_pr__nfet_01v8_lvt_E33R59_0
timestamp 1696271506
transform 0 1 -299 -1 0 -122
box -226 -279 226 279
use trimcap  trimcap_1
timestamp 1696109480
transform 1 0 -566 0 1 -262
box 0 376 476 1324
<< labels >>
flabel metal1 -390 920 -266 1036 0 FreeSans 480 0 0 0 todrain
flabel metal1 -204 -152 -146 -92 0 FreeSans 480 0 0 0 d_i
flabel metal1 -372 -196 -286 -168 0 FreeSans 480 0 0 0 tovss
<< end >>
