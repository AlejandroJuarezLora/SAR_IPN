magic
tech sky130B
magscale 1 2
timestamp 1697663034
<< metal1 >>
rect 13417 -260 13506 -244
rect 13416 -349 13422 -260
rect 13511 -349 13517 -260
rect 14247 -339 14253 -263
rect 14329 -339 14335 -263
rect 22670 -1288 23032 -1225
rect 23095 -1288 27211 -1225
rect 24241 -1805 24325 -1799
rect 24325 -1889 27237 -1805
rect 24241 -1895 24325 -1889
rect 25060 -2424 25144 -2418
rect 25144 -2508 27223 -2424
rect 25060 -2514 25144 -2508
<< via1 >>
rect 13422 -349 13511 -260
rect 14253 -339 14329 -263
rect 23032 -1288 23095 -1225
rect 24241 -1889 24325 -1805
rect 25060 -2508 25144 -2424
<< metal2 >>
rect 13422 -1 13511 0
rect 13417 -90 27222 -1
rect 13422 -260 13511 -90
rect 13422 -355 13511 -349
rect 14253 -263 14329 -257
rect 14253 -628 14329 -339
rect 14253 -704 27217 -628
rect 23032 -1225 23095 -1219
rect 22670 -1288 22679 -1225
rect 22742 -1288 23032 -1225
rect 23032 -1294 23095 -1288
rect 24246 -1805 24320 -1801
rect 24235 -1889 24241 -1805
rect 24325 -1889 24331 -1805
rect 25852 -1826 25923 -1821
rect 25847 -1830 26616 -1826
rect 24246 -1893 24320 -1889
rect 25847 -1905 25852 -1830
rect 25923 -1905 26616 -1830
rect 25847 -1907 26616 -1905
rect 25852 -1914 25923 -1907
rect 25065 -2424 25139 -2420
rect 25054 -2508 25060 -2424
rect 25144 -2508 25150 -2424
rect 25065 -2512 25139 -2508
rect 26535 -2999 26616 -1907
rect 26529 -3005 26623 -2999
rect 25847 -3035 26349 -3029
rect 25843 -3106 25852 -3035
rect 25923 -3106 26349 -3035
rect 26529 -3087 27237 -3005
rect 26529 -3093 26623 -3087
rect 25847 -3110 26349 -3106
rect 26268 -3599 26349 -3110
rect 26268 -3680 27238 -3599
rect 26267 -3822 26341 -3818
rect 26256 -3827 26352 -3822
rect 26256 -3901 26267 -3827
rect 26341 -3901 26352 -3827
rect 26256 -3906 26352 -3901
rect 26261 -3910 26341 -3906
rect 26261 -4233 26334 -3910
rect 26261 -4306 27229 -4233
rect 26270 -4427 26354 -4416
rect 26270 -4501 26275 -4427
rect 26349 -4501 26354 -4427
rect 26270 -4512 26354 -4501
rect 26280 -4812 26343 -4512
rect 26280 -4875 27212 -4812
<< via2 >>
rect 13427 -344 13506 -265
rect 14258 -334 14324 -268
rect 22679 -1288 22742 -1225
rect 24246 -1884 24320 -1810
rect 25852 -1905 25923 -1830
rect 25065 -2503 25139 -2429
rect 25852 -3106 25923 -3035
rect 26267 -3901 26341 -3827
rect 26275 -4501 26349 -4427
<< metal3 >>
rect 1056 -265 13511 -260
rect 1056 -344 13427 -265
rect 13506 -344 13511 -265
rect 1056 -349 13511 -344
rect 13833 -268 14329 -263
rect 13833 -334 14258 -268
rect 14324 -334 14329 -268
rect 13833 -339 14329 -334
rect 14623 -290 15522 -214
rect 1056 -874 1145 -349
rect 1056 -963 13160 -874
rect 13071 -1466 13160 -963
rect 1007 -1555 13160 -1466
rect 1007 -2123 1096 -1555
rect 1007 -2212 13127 -2123
rect 13038 -2732 13127 -2212
rect 1024 -2821 13127 -2732
rect 1024 -3323 1113 -2821
rect 1024 -3412 13111 -3323
rect 13022 -3849 13111 -3412
rect 991 -3938 13111 -3849
rect 991 -4474 1080 -3938
rect 991 -4563 13111 -4474
rect 13833 -4487 13909 -339
rect 14623 -4487 14699 -290
rect 13833 -4563 14699 -4487
rect 15446 -4471 15522 -290
rect 16236 -306 17102 -230
rect 24241 -247 24325 -222
rect 16236 -4471 16312 -306
rect 15446 -4547 16312 -4471
rect 17026 -4454 17102 -306
rect 17864 -323 18714 -247
rect 22679 -254 22742 -253
rect 17864 -4454 17940 -323
rect 17026 -4530 17940 -4454
rect 18638 -4487 18714 -323
rect 19434 -333 19526 -257
rect 19436 -4487 19512 -333
rect 18638 -4563 19512 -4487
rect 20237 -4526 20300 -296
rect 21069 -368 21901 -305
rect 22660 -317 22761 -254
rect 21069 -4526 21132 -368
rect 20237 -4589 21132 -4526
rect 21838 -4526 21901 -368
rect 22679 -1158 22742 -317
rect 23462 -331 24325 -247
rect 22614 -1225 22809 -1158
rect 22614 -1288 22679 -1225
rect 22742 -1288 22809 -1225
rect 22614 -1353 22809 -1288
rect 22679 -4526 22742 -1353
rect 21838 -4589 22742 -4526
rect 23462 -4475 23546 -331
rect 24241 -1810 24325 -331
rect 24241 -1884 24246 -1810
rect 24320 -1884 24325 -1810
rect 24241 -4475 24325 -1884
rect 23462 -4559 24325 -4475
rect 25060 -2429 25144 -222
rect 25847 -1830 25928 -329
rect 25847 -1905 25852 -1830
rect 25923 -1905 25928 -1830
rect 25847 -2400 25928 -1905
rect 25060 -2503 25065 -2429
rect 25139 -2503 25144 -2429
rect 25060 -4645 25144 -2503
rect 25847 -3035 25928 -2521
rect 25847 -3106 25852 -3035
rect 25923 -3106 25928 -3035
rect 25847 -3450 25928 -3106
rect 25945 -3827 26346 -3822
rect 25945 -3901 26267 -3827
rect 26341 -3901 26346 -3827
rect 25945 -3906 26346 -3901
rect 25958 -4427 26354 -4422
rect 25958 -4501 26275 -4427
rect 26349 -4501 26354 -4427
rect 25958 -4506 26354 -4501
<< metal4 >>
rect 257 198 26743 258
rect 257 -408 317 198
rect 257 -468 25856 -408
rect 257 -1022 317 -468
rect 257 -1082 25934 -1022
rect 257 -1590 317 -1082
rect 257 -1650 25914 -1590
rect 257 -2210 317 -1650
rect 257 -2270 25934 -2210
rect 257 -2810 317 -2270
rect 257 -2870 25904 -2810
rect 257 -3392 317 -2870
rect 257 -3452 25934 -3392
rect 257 -4002 317 -3452
rect 257 -4062 25944 -4002
rect 257 -4602 317 -4062
rect 257 -4662 25914 -4602
rect 257 -5134 317 -4662
rect 26683 -5134 26743 198
rect 257 -5194 26743 -5134
rect 257 -5215 317 -5194
use unitcap  unitcap_0
timestamp 1696453761
transform 1 0 2462 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_1
timestamp 1696453761
transform 1 0 2462 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_2
timestamp 1696453761
transform 1 0 2462 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_3
timestamp 1696453761
transform 1 0 2462 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_4
timestamp 1696453761
transform 1 0 2462 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_5
timestamp 1696453761
transform 1 0 2462 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_6
timestamp 1696453761
transform 1 0 2462 0 1 -600
box 0 0 486 480
use unitcap  unitcap_7
timestamp 1696453761
transform 1 0 2462 0 1 0
box 0 0 486 480
use unitcap  unitcap_8
timestamp 1696453761
transform 1 0 62 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_9
timestamp 1696453761
transform 1 0 62 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_10
timestamp 1696453761
transform 1 0 62 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_11
timestamp 1696453761
transform 1 0 62 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_12
timestamp 1696453761
transform 1 0 62 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_13
timestamp 1696453761
transform 1 0 62 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_14
timestamp 1696453761
transform 1 0 62 0 1 -600
box 0 0 486 480
use unitcap  unitcap_15
timestamp 1696453761
transform 1 0 62 0 1 0
box 0 0 486 480
use unitcap  unitcap_16
timestamp 1696453761
transform 1 0 862 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_17
timestamp 1696453761
transform 1 0 862 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_18
timestamp 1696453761
transform 1 0 862 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_19
timestamp 1696453761
transform 1 0 862 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_20
timestamp 1696453761
transform 1 0 862 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_21
timestamp 1696453761
transform 1 0 862 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_22
timestamp 1696453761
transform 1 0 862 0 1 -600
box 0 0 486 480
use unitcap  unitcap_23
timestamp 1696453761
transform 1 0 862 0 1 0
box 0 0 486 480
use unitcap  unitcap_24
timestamp 1696453761
transform 1 0 1662 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_25
timestamp 1696453761
transform 1 0 1662 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_26
timestamp 1696453761
transform 1 0 1662 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_27
timestamp 1696453761
transform 1 0 1662 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_28
timestamp 1696453761
transform 1 0 1662 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_29
timestamp 1696453761
transform 1 0 1662 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_30
timestamp 1696453761
transform 1 0 1662 0 1 -600
box 0 0 486 480
use unitcap  unitcap_31
timestamp 1696453761
transform 1 0 1662 0 1 0
box 0 0 486 480
use unitcap  unitcap_32
timestamp 1696453761
transform 1 0 4062 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_33
timestamp 1696453761
transform 1 0 4062 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_34
timestamp 1696453761
transform 1 0 4062 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_35
timestamp 1696453761
transform 1 0 4062 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_36
timestamp 1696453761
transform 1 0 4062 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_37
timestamp 1696453761
transform 1 0 4062 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_38
timestamp 1696453761
transform 1 0 4062 0 1 -600
box 0 0 486 480
use unitcap  unitcap_39
timestamp 1696453761
transform 1 0 4062 0 1 0
box 0 0 486 480
use unitcap  unitcap_40
timestamp 1696453761
transform 1 0 3262 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_41
timestamp 1696453761
transform 1 0 3262 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_42
timestamp 1696453761
transform 1 0 3262 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_43
timestamp 1696453761
transform 1 0 3262 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_44
timestamp 1696453761
transform 1 0 3262 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_45
timestamp 1696453761
transform 1 0 3262 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_46
timestamp 1696453761
transform 1 0 3262 0 1 -600
box 0 0 486 480
use unitcap  unitcap_47
timestamp 1696453761
transform 1 0 3262 0 1 0
box 0 0 486 480
use unitcap  unitcap_48
timestamp 1696453761
transform 1 0 5662 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_49
timestamp 1696453761
transform 1 0 5662 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_50
timestamp 1696453761
transform 1 0 5662 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_51
timestamp 1696453761
transform 1 0 5662 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_52
timestamp 1696453761
transform 1 0 5662 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_53
timestamp 1696453761
transform 1 0 5662 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_54
timestamp 1696453761
transform 1 0 5662 0 1 -600
box 0 0 486 480
use unitcap  unitcap_55
timestamp 1696453761
transform 1 0 5662 0 1 0
box 0 0 486 480
use unitcap  unitcap_56
timestamp 1696453761
transform 1 0 4862 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_57
timestamp 1696453761
transform 1 0 4862 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_58
timestamp 1696453761
transform 1 0 4862 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_59
timestamp 1696453761
transform 1 0 4862 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_60
timestamp 1696453761
transform 1 0 4862 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_61
timestamp 1696453761
transform 1 0 4862 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_62
timestamp 1696453761
transform 1 0 4862 0 1 -600
box 0 0 486 480
use unitcap  unitcap_63
timestamp 1696453761
transform 1 0 4862 0 1 0
box 0 0 486 480
use unitcap  unitcap_64
timestamp 1696453761
transform 1 0 8062 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_65
timestamp 1696453761
transform 1 0 8062 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_66
timestamp 1696453761
transform 1 0 8062 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_67
timestamp 1696453761
transform 1 0 8062 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_68
timestamp 1696453761
transform 1 0 8062 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_69
timestamp 1696453761
transform 1 0 8062 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_70
timestamp 1696453761
transform 1 0 8062 0 1 -600
box 0 0 486 480
use unitcap  unitcap_71
timestamp 1696453761
transform 1 0 8062 0 1 0
box 0 0 486 480
use unitcap  unitcap_72
timestamp 1696453761
transform 1 0 6462 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_73
timestamp 1696453761
transform 1 0 6462 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_74
timestamp 1696453761
transform 1 0 6462 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_75
timestamp 1696453761
transform 1 0 6462 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_76
timestamp 1696453761
transform 1 0 6462 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_77
timestamp 1696453761
transform 1 0 6462 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_78
timestamp 1696453761
transform 1 0 6462 0 1 -600
box 0 0 486 480
use unitcap  unitcap_79
timestamp 1696453761
transform 1 0 6462 0 1 0
box 0 0 486 480
use unitcap  unitcap_80
timestamp 1696453761
transform 1 0 7262 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_81
timestamp 1696453761
transform 1 0 7262 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_82
timestamp 1696453761
transform 1 0 7262 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_83
timestamp 1696453761
transform 1 0 7262 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_84
timestamp 1696453761
transform 1 0 7262 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_85
timestamp 1696453761
transform 1 0 7262 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_86
timestamp 1696453761
transform 1 0 7262 0 1 -600
box 0 0 486 480
use unitcap  unitcap_87
timestamp 1696453761
transform 1 0 7262 0 1 0
box 0 0 486 480
use unitcap  unitcap_88
timestamp 1696453761
transform 1 0 8862 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_89
timestamp 1696453761
transform 1 0 8862 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_90
timestamp 1696453761
transform 1 0 8862 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_91
timestamp 1696453761
transform 1 0 8862 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_92
timestamp 1696453761
transform 1 0 8862 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_93
timestamp 1696453761
transform 1 0 8862 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_94
timestamp 1696453761
transform 1 0 8862 0 1 -600
box 0 0 486 480
use unitcap  unitcap_95
timestamp 1696453761
transform 1 0 8862 0 1 0
box 0 0 486 480
use unitcap  unitcap_96
timestamp 1696453761
transform 1 0 10462 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_97
timestamp 1696453761
transform 1 0 10462 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_98
timestamp 1696453761
transform 1 0 10462 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_99
timestamp 1696453761
transform 1 0 10462 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_100
timestamp 1696453761
transform 1 0 10462 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_101
timestamp 1696453761
transform 1 0 10462 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_102
timestamp 1696453761
transform 1 0 10462 0 1 -600
box 0 0 486 480
use unitcap  unitcap_103
timestamp 1696453761
transform 1 0 10462 0 1 0
box 0 0 486 480
use unitcap  unitcap_104
timestamp 1696453761
transform 1 0 9662 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_105
timestamp 1696453761
transform 1 0 9662 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_106
timestamp 1696453761
transform 1 0 9662 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_107
timestamp 1696453761
transform 1 0 9662 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_108
timestamp 1696453761
transform 1 0 9662 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_109
timestamp 1696453761
transform 1 0 9662 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_110
timestamp 1696453761
transform 1 0 9662 0 1 -600
box 0 0 486 480
use unitcap  unitcap_111
timestamp 1696453761
transform 1 0 9662 0 1 0
box 0 0 486 480
use unitcap  unitcap_112
timestamp 1696453761
transform 1 0 12062 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_113
timestamp 1696453761
transform 1 0 12062 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_114
timestamp 1696453761
transform 1 0 12062 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_115
timestamp 1696453761
transform 1 0 12062 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_116
timestamp 1696453761
transform 1 0 12062 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_117
timestamp 1696453761
transform 1 0 12062 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_118
timestamp 1696453761
transform 1 0 12062 0 1 -600
box 0 0 486 480
use unitcap  unitcap_119
timestamp 1696453761
transform 1 0 12062 0 1 0
box 0 0 486 480
use unitcap  unitcap_120
timestamp 1696453761
transform 1 0 11262 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_121
timestamp 1696453761
transform 1 0 11262 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_122
timestamp 1696453761
transform 1 0 11262 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_123
timestamp 1696453761
transform 1 0 11262 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_124
timestamp 1696453761
transform 1 0 11262 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_125
timestamp 1696453761
transform 1 0 11262 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_126
timestamp 1696453761
transform 1 0 11262 0 1 -600
box 0 0 486 480
use unitcap  unitcap_127
timestamp 1696453761
transform 1 0 11262 0 1 0
box 0 0 486 480
use unitcap  unitcap_128
timestamp 1696453761
transform 1 0 13662 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_129
timestamp 1696453761
transform 1 0 13662 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_130
timestamp 1696453761
transform 1 0 13662 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_131
timestamp 1696453761
transform 1 0 13662 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_132
timestamp 1696453761
transform 1 0 13662 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_133
timestamp 1696453761
transform 1 0 13662 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_134
timestamp 1696453761
transform 1 0 13662 0 1 -600
box 0 0 486 480
use unitcap  unitcap_135
timestamp 1696453761
transform 1 0 13662 0 1 0
box 0 0 486 480
use unitcap  unitcap_136
timestamp 1696453761
transform 1 0 12862 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_137
timestamp 1696453761
transform 1 0 12862 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_138
timestamp 1696453761
transform 1 0 12862 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_139
timestamp 1696453761
transform 1 0 12862 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_140
timestamp 1696453761
transform 1 0 12862 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_141
timestamp 1696453761
transform 1 0 12862 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_142
timestamp 1696453761
transform 1 0 12862 0 1 -600
box 0 0 486 480
use unitcap  unitcap_143
timestamp 1696453761
transform 1 0 12862 0 1 0
box 0 0 486 480
use unitcap  unitcap_144
timestamp 1696453761
transform 1 0 15262 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_145
timestamp 1696453761
transform 1 0 15262 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_146
timestamp 1696453761
transform 1 0 15262 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_147
timestamp 1696453761
transform 1 0 15262 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_148
timestamp 1696453761
transform 1 0 15262 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_149
timestamp 1696453761
transform 1 0 15262 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_150
timestamp 1696453761
transform 1 0 15262 0 1 -600
box 0 0 486 480
use unitcap  unitcap_151
timestamp 1696453761
transform 1 0 15262 0 1 0
box 0 0 486 480
use unitcap  unitcap_152
timestamp 1696453761
transform 1 0 14462 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_153
timestamp 1696453761
transform 1 0 14462 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_154
timestamp 1696453761
transform 1 0 14462 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_155
timestamp 1696453761
transform 1 0 14462 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_156
timestamp 1696453761
transform 1 0 14462 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_157
timestamp 1696453761
transform 1 0 14462 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_158
timestamp 1696453761
transform 1 0 14462 0 1 -600
box 0 0 486 480
use unitcap  unitcap_159
timestamp 1696453761
transform 1 0 14462 0 1 0
box 0 0 486 480
use unitcap  unitcap_160
timestamp 1696453761
transform 1 0 16062 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_161
timestamp 1696453761
transform 1 0 16062 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_162
timestamp 1696453761
transform 1 0 16062 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_163
timestamp 1696453761
transform 1 0 16062 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_164
timestamp 1696453761
transform 1 0 16062 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_165
timestamp 1696453761
transform 1 0 16062 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_166
timestamp 1696453761
transform 1 0 16062 0 1 -600
box 0 0 486 480
use unitcap  unitcap_167
timestamp 1696453761
transform 1 0 16062 0 1 0
box 0 0 486 480
use unitcap  unitcap_168
timestamp 1696453761
transform 1 0 17662 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_169
timestamp 1696453761
transform 1 0 17662 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_170
timestamp 1696453761
transform 1 0 17662 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_171
timestamp 1696453761
transform 1 0 17662 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_172
timestamp 1696453761
transform 1 0 17662 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_173
timestamp 1696453761
transform 1 0 17662 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_174
timestamp 1696453761
transform 1 0 17662 0 1 -600
box 0 0 486 480
use unitcap  unitcap_175
timestamp 1696453761
transform 1 0 17662 0 1 0
box 0 0 486 480
use unitcap  unitcap_176
timestamp 1696453761
transform 1 0 16862 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_177
timestamp 1696453761
transform 1 0 16862 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_178
timestamp 1696453761
transform 1 0 16862 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_179
timestamp 1696453761
transform 1 0 16862 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_180
timestamp 1696453761
transform 1 0 16862 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_181
timestamp 1696453761
transform 1 0 16862 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_182
timestamp 1696453761
transform 1 0 16862 0 1 -600
box 0 0 486 480
use unitcap  unitcap_183
timestamp 1696453761
transform 1 0 16862 0 1 0
box 0 0 486 480
use unitcap  unitcap_184
timestamp 1696453761
transform 1 0 20062 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_185
timestamp 1696453761
transform 1 0 20062 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_186
timestamp 1696453761
transform 1 0 20062 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_187
timestamp 1696453761
transform 1 0 20062 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_188
timestamp 1696453761
transform 1 0 20062 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_189
timestamp 1696453761
transform 1 0 20062 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_190
timestamp 1696453761
transform 1 0 20062 0 1 -600
box 0 0 486 480
use unitcap  unitcap_191
timestamp 1696453761
transform 1 0 20062 0 1 0
box 0 0 486 480
use unitcap  unitcap_192
timestamp 1696453761
transform 1 0 18462 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_193
timestamp 1696453761
transform 1 0 18462 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_194
timestamp 1696453761
transform 1 0 18462 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_195
timestamp 1696453761
transform 1 0 18462 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_196
timestamp 1696453761
transform 1 0 18462 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_197
timestamp 1696453761
transform 1 0 18462 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_198
timestamp 1696453761
transform 1 0 18462 0 1 -600
box 0 0 486 480
use unitcap  unitcap_199
timestamp 1696453761
transform 1 0 18462 0 1 0
box 0 0 486 480
use unitcap  unitcap_200
timestamp 1696453761
transform 1 0 19262 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_201
timestamp 1696453761
transform 1 0 19262 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_202
timestamp 1696453761
transform 1 0 19262 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_203
timestamp 1696453761
transform 1 0 19262 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_204
timestamp 1696453761
transform 1 0 19262 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_205
timestamp 1696453761
transform 1 0 19262 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_206
timestamp 1696453761
transform 1 0 19262 0 1 -600
box 0 0 486 480
use unitcap  unitcap_207
timestamp 1696453761
transform 1 0 19262 0 1 0
box 0 0 486 480
use unitcap  unitcap_208
timestamp 1696453761
transform 1 0 20862 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_209
timestamp 1696453761
transform 1 0 20862 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_210
timestamp 1696453761
transform 1 0 20862 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_211
timestamp 1696453761
transform 1 0 20862 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_212
timestamp 1696453761
transform 1 0 20862 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_213
timestamp 1696453761
transform 1 0 20862 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_214
timestamp 1696453761
transform 1 0 20862 0 1 -600
box 0 0 486 480
use unitcap  unitcap_215
timestamp 1696453761
transform 1 0 20862 0 1 0
box 0 0 486 480
use unitcap  unitcap_216
timestamp 1696453761
transform 1 0 22462 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_217
timestamp 1696453761
transform 1 0 22462 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_218
timestamp 1696453761
transform 1 0 22462 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_219
timestamp 1696453761
transform 1 0 22462 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_220
timestamp 1696453761
transform 1 0 22462 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_221
timestamp 1696453761
transform 1 0 22462 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_222
timestamp 1696453761
transform 1 0 22462 0 1 -600
box 0 0 486 480
use unitcap  unitcap_223
timestamp 1696453761
transform 1 0 22462 0 1 0
box 0 0 486 480
use unitcap  unitcap_224
timestamp 1696453761
transform 1 0 21662 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_225
timestamp 1696453761
transform 1 0 21662 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_226
timestamp 1696453761
transform 1 0 21662 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_227
timestamp 1696453761
transform 1 0 21662 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_228
timestamp 1696453761
transform 1 0 21662 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_229
timestamp 1696453761
transform 1 0 21662 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_230
timestamp 1696453761
transform 1 0 21662 0 1 -600
box 0 0 486 480
use unitcap  unitcap_231
timestamp 1696453761
transform 1 0 21662 0 1 0
box 0 0 486 480
use unitcap  unitcap_232
timestamp 1696453761
transform 1 0 24062 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_233
timestamp 1696453761
transform 1 0 24062 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_234
timestamp 1696453761
transform 1 0 24062 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_235
timestamp 1696453761
transform 1 0 24062 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_236
timestamp 1696453761
transform 1 0 24062 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_237
timestamp 1696453761
transform 1 0 24062 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_238
timestamp 1696453761
transform 1 0 24062 0 1 -600
box 0 0 486 480
use unitcap  unitcap_239
timestamp 1696453761
transform 1 0 24062 0 1 0
box 0 0 486 480
use unitcap  unitcap_240
timestamp 1696453761
transform 1 0 23262 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_241
timestamp 1696453761
transform 1 0 23262 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_242
timestamp 1696453761
transform 1 0 23262 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_243
timestamp 1696453761
transform 1 0 23262 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_244
timestamp 1696453761
transform 1 0 23262 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_245
timestamp 1696453761
transform 1 0 23262 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_246
timestamp 1696453761
transform 1 0 23262 0 1 -600
box 0 0 486 480
use unitcap  unitcap_247
timestamp 1696453761
transform 1 0 23262 0 1 0
box 0 0 486 480
use unitcap  unitcap_248
timestamp 1696453761
transform 1 0 24862 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_249
timestamp 1696453761
transform 1 0 24862 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_250
timestamp 1696453761
transform 1 0 24862 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_251
timestamp 1696453761
transform 1 0 24862 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_252
timestamp 1696453761
transform 1 0 24862 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_253
timestamp 1696453761
transform 1 0 24862 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_254
timestamp 1696453761
transform 1 0 24862 0 1 -600
box 0 0 486 480
use unitcap  unitcap_255
timestamp 1696453761
transform 1 0 24862 0 1 0
box 0 0 486 480
use unitcap  unitcap_256
timestamp 1696453761
transform 1 0 62 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_257
timestamp 1696453761
transform 1 0 862 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_258
timestamp 1696453761
transform 1 0 1662 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_259
timestamp 1696453761
transform 1 0 2462 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_260
timestamp 1696453761
transform 1 0 3262 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_261
timestamp 1696453761
transform 1 0 4062 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_262
timestamp 1696453761
transform 1 0 4862 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_263
timestamp 1696453761
transform 1 0 5662 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_264
timestamp 1696453761
transform 1 0 6462 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_265
timestamp 1696453761
transform 1 0 7262 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_266
timestamp 1696453761
transform 1 0 8062 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_267
timestamp 1696453761
transform 1 0 8862 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_268
timestamp 1696453761
transform 1 0 9662 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_269
timestamp 1696453761
transform 1 0 10462 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_270
timestamp 1696453761
transform 1 0 11262 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_271
timestamp 1696453761
transform 1 0 12062 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_272
timestamp 1696453761
transform 1 0 12862 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_273
timestamp 1696453761
transform 1 0 13662 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_274
timestamp 1696453761
transform 1 0 14462 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_275
timestamp 1696453761
transform 1 0 15262 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_276
timestamp 1696453761
transform 1 0 16062 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_277
timestamp 1696453761
transform 1 0 16862 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_278
timestamp 1696453761
transform 1 0 17662 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_279
timestamp 1696453761
transform 1 0 18462 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_280
timestamp 1696453761
transform 1 0 20062 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_281
timestamp 1696453761
transform 1 0 19262 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_282
timestamp 1696453761
transform 1 0 20862 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_283
timestamp 1696453761
transform 1 0 22462 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_284
timestamp 1696453761
transform 1 0 21662 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_285
timestamp 1696453761
transform 1 0 24062 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_286
timestamp 1696453761
transform 1 0 23262 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_287
timestamp 1696453761
transform 1 0 24862 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_288
timestamp 1696453761
transform 1 0 62 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_289
timestamp 1696453761
transform 1 0 862 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_290
timestamp 1696453761
transform 1 0 1662 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_291
timestamp 1696453761
transform 1 0 2462 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_292
timestamp 1696453761
transform 1 0 3262 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_293
timestamp 1696453761
transform 1 0 4062 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_294
timestamp 1696453761
transform 1 0 4862 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_295
timestamp 1696453761
transform 1 0 5662 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_296
timestamp 1696453761
transform 1 0 6462 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_297
timestamp 1696453761
transform 1 0 7262 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_298
timestamp 1696453761
transform 1 0 8062 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_299
timestamp 1696453761
transform 1 0 8862 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_300
timestamp 1696453761
transform 1 0 9662 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_301
timestamp 1696453761
transform 1 0 10462 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_302
timestamp 1696453761
transform 1 0 11262 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_303
timestamp 1696453761
transform 1 0 12062 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_304
timestamp 1696453761
transform 1 0 12862 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_305
timestamp 1696453761
transform 1 0 13662 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_306
timestamp 1696453761
transform 1 0 14462 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_307
timestamp 1696453761
transform 1 0 15262 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_308
timestamp 1696453761
transform 1 0 16062 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_309
timestamp 1696453761
transform 1 0 16862 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_310
timestamp 1696453761
transform 1 0 17662 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_311
timestamp 1696453761
transform 1 0 18462 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_312
timestamp 1696453761
transform 1 0 20062 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_313
timestamp 1696453761
transform 1 0 19262 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_314
timestamp 1696453761
transform 1 0 20862 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_315
timestamp 1696453761
transform 1 0 22462 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_316
timestamp 1696453761
transform 1 0 21662 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_317
timestamp 1696453761
transform 1 0 24062 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_318
timestamp 1696453761
transform 1 0 23262 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_319
timestamp 1696453761
transform 1 0 24862 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_320
timestamp 1696453761
transform 1 0 26462 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_321
timestamp 1696453761
transform 1 0 25662 0 1 -5400
box 0 0 486 480
use unitcap  unitcap_322
timestamp 1696453761
transform 1 0 26462 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_323
timestamp 1696453761
transform 1 0 25662 0 1 -4200
box 0 0 486 480
use unitcap  unitcap_324
timestamp 1696453761
transform 1 0 26462 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_325
timestamp 1696453761
transform 1 0 25662 0 1 -4800
box 0 0 486 480
use unitcap  unitcap_326
timestamp 1696453761
transform 1 0 26462 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_327
timestamp 1696453761
transform 1 0 25662 0 1 -3000
box 0 0 486 480
use unitcap  unitcap_328
timestamp 1696453761
transform 1 0 26462 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_329
timestamp 1696453761
transform 1 0 25662 0 1 -3600
box 0 0 486 480
use unitcap  unitcap_330
timestamp 1696453761
transform 1 0 26462 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_331
timestamp 1696453761
transform 1 0 26462 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_332
timestamp 1696453761
transform 1 0 25662 0 1 -1200
box 0 0 486 480
use unitcap  unitcap_333
timestamp 1696453761
transform 1 0 25662 0 1 -1800
box 0 0 486 480
use unitcap  unitcap_334
timestamp 1696453761
transform 1 0 26462 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_335
timestamp 1696453761
transform 1 0 25662 0 1 -2400
box 0 0 486 480
use unitcap  unitcap_336
timestamp 1696453761
transform 1 0 26462 0 1 0
box 0 0 486 480
use unitcap  unitcap_337
timestamp 1696453761
transform 1 0 26462 0 1 -600
box 0 0 486 480
use unitcap  unitcap_338
timestamp 1696453761
transform 1 0 25662 0 1 0
box 0 0 486 480
use unitcap  unitcap_339
timestamp 1696453761
transform 1 0 25662 0 1 -600
box 0 0 486 480
<< labels >>
flabel metal1 s 27132 -2508 27216 -2424 0 FreeSans 640 90 0 0 n3
flabel metal1 s 27153 -1889 27237 -1805 0 FreeSans 640 90 0 0 n4
flabel metal1 s 27148 -1288 27211 -1225 0 FreeSans 640 90 0 0 n5
flabel metal2 s 27155 -3087 27237 -3005 0 FreeSans 640 0 0 0 n2
flabel metal2 27149 -4875 27212 -4812 0 FreeSans 640 0 0 0 ndum
flabel metal2 s 27156 -4306 27229 -4233 0 FreeSans 640 0 0 0 n0
flabel metal2 27157 -3680 27238 -3599 0 FreeSans 640 0 0 0 n1
flabel metal2 27133 -90 27222 -1 0 FreeSans 640 0 0 0 n7
flabel metal2 27136 -704 27212 -628 0 FreeSans 640 0 0 0 n6
flabel metal4 257 -5215 317 258 0 FreeSans 800 0 0 0 top
<< end >>
