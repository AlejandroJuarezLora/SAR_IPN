magic
tech sky130B
magscale 1 2
timestamp 1697836898
<< locali >>
rect 33137 9133 33183 9149
rect 28817 9087 33183 9133
rect 33137 7445 33183 9087
rect 33804 7445 33850 7456
rect 32443 7399 33850 7445
rect 32443 6075 32489 7399
rect 33804 7264 33850 7399
rect 32156 6024 32489 6075
rect 32156 6023 32428 6024
rect 28147 4501 28279 4535
rect 33145 4526 33179 5083
rect 28147 2897 28181 4501
rect 32501 4492 33179 4526
rect 28147 2863 28299 2897
<< metal1 >>
rect 28235 12072 31318 12167
rect 31413 12072 31419 12167
rect 28235 11909 28330 12072
rect 28781 11964 32208 12006
rect 28781 11912 28986 11964
rect 29038 11912 32208 11964
rect 28781 11911 32208 11912
rect 32303 11911 32309 12006
rect -305 11847 -211 11853
rect -861 11781 -767 11787
rect -861 9874 -767 11687
rect -305 10412 -211 11753
rect -305 10318 94 10412
rect -861 9780 173 9874
rect 29444 9037 29490 9236
rect 30686 9042 30730 9236
rect 31774 9055 31820 9236
rect 32293 9022 32337 9236
rect 33027 8873 33077 9236
rect -1106 8526 160 8562
rect 32762 7546 32814 7552
rect 32814 7504 33776 7536
rect 32762 7488 32814 7494
rect 33744 7234 33776 7504
rect 31190 6510 31242 6516
rect 31190 6452 31242 6458
rect 31200 6295 31232 6452
rect 34399 6139 34502 6199
rect 29992 6079 29998 6131
rect 30050 6079 30056 6131
rect 29984 5958 29990 6018
rect 30050 5958 30056 6018
rect 31182 5588 31214 5795
rect 31172 5582 31224 5588
rect 31172 5524 31224 5530
rect 33732 5064 33738 5116
rect 33790 5064 33796 5116
rect -1072 3444 220 3480
rect 29467 2727 29513 2936
rect 30709 2712 30753 2937
rect 31797 2721 31843 2963
rect 32316 2718 32360 2976
rect 33050 2701 33100 3031
rect -869 2132 177 2226
rect -869 755 -775 2132
rect -869 655 -775 661
rect -307 1594 94 1688
rect -307 755 -213 1594
rect -307 655 -213 661
rect 28235 -44 28330 97
rect 31956 95 32051 101
rect 28781 0 31956 95
rect 31956 -6 32051 0
rect 31398 -44 31493 -38
rect 28235 -70 31398 -44
rect 28235 -122 28938 -70
rect 28990 -122 31398 -70
rect 28235 -139 31398 -122
rect 31398 -145 31493 -139
<< via1 >>
rect 31318 12072 31413 12167
rect 28986 11912 29038 11964
rect 32208 11911 32303 12006
rect -861 11687 -767 11781
rect -305 11753 -211 11847
rect 32762 7494 32814 7546
rect 31190 6458 31242 6510
rect 29998 6079 30050 6131
rect 29990 5958 30050 6018
rect 31172 5530 31224 5582
rect 33738 5064 33790 5116
rect -869 661 -775 755
rect -307 661 -213 755
rect 31956 0 32051 95
rect 28938 -122 28990 -70
rect 31398 -139 31493 -44
<< metal2 >>
rect 31318 12167 31413 12173
rect 31309 12072 31318 12167
rect 31413 12072 31422 12167
rect 31318 12066 31413 12072
rect 32208 12006 32303 12012
rect 28986 11964 29038 11970
rect 28986 11906 29038 11912
rect 32199 11911 32208 12006
rect 32303 11911 32312 12006
rect -305 11847 -211 11856
rect -870 11687 -861 11781
rect -767 11687 -758 11781
rect -311 11753 -305 11847
rect -211 11753 -205 11847
rect -305 11744 -211 11753
rect 28995 11707 29028 11906
rect 32208 11905 32303 11911
rect 28951 11674 29028 11707
rect 28923 11395 29047 11429
rect 28929 11124 29045 11158
rect 28937 10847 29045 10881
rect 28931 10573 29045 10607
rect 48 1528 89 10480
rect 28927 10298 29045 10332
rect 28929 10022 29047 10056
rect 28935 9747 29039 9781
rect 28941 9473 29033 9507
rect 32756 7536 32762 7546
rect 31200 7504 32762 7536
rect 31200 6510 31232 7504
rect 32756 7494 32762 7504
rect 32814 7494 32820 7546
rect 32982 7460 34476 7488
rect 29152 6460 29208 6469
rect 31184 6458 31190 6510
rect 31242 6458 31248 6510
rect 29208 6415 30041 6450
rect 29152 6395 29208 6404
rect 30006 6137 30041 6415
rect 29998 6131 30050 6137
rect 29998 6073 30050 6079
rect 29990 6018 30050 6024
rect 29990 5954 30050 5958
rect 29983 5898 29992 5954
rect 30048 5898 30057 5954
rect 29990 5896 30050 5898
rect 32982 5646 33010 7460
rect 32228 5616 33011 5646
rect 31166 5530 31172 5582
rect 31224 5530 31230 5582
rect 31182 4932 31214 5530
rect 33738 5116 33790 5122
rect 33738 5058 33790 5064
rect 33748 4932 33780 5058
rect 31182 4900 33780 4932
rect 28933 2499 29043 2533
rect 28925 2225 29043 2259
rect 28927 1950 29043 1984
rect 28931 1674 29041 1708
rect 28939 1399 29037 1433
rect 28925 1125 29031 1159
rect 28935 848 29029 882
rect -869 755 -775 764
rect -307 755 -213 764
rect -875 661 -869 755
rect -775 661 -769 755
rect -313 661 -307 755
rect -213 661 -207 755
rect -869 652 -775 661
rect -307 652 -213 661
rect 28927 577 29033 611
rect 28947 -64 28981 333
rect 31956 95 32051 104
rect 31950 0 31956 95
rect 32051 0 32057 95
rect 31956 -9 32051 0
rect 31398 -44 31493 -35
rect 28938 -70 28990 -64
rect 28938 -128 28990 -122
rect 31392 -139 31398 -44
rect 31493 -139 31499 -44
rect 31398 -148 31493 -139
<< via2 >>
rect 31318 12072 31413 12167
rect 32208 11911 32303 12006
rect -861 11687 -767 11781
rect -305 11753 -211 11847
rect 29152 6404 29208 6460
rect 29992 5898 30048 5954
rect -869 661 -775 755
rect -307 661 -213 755
rect 31956 0 32051 95
rect 31398 -139 31493 -44
<< metal3 >>
rect 31313 12167 31323 12172
rect 31313 12072 31318 12167
rect 31313 12067 31323 12072
rect 31418 12067 31424 12172
rect 32203 12006 32213 12011
rect 32203 11911 32208 12006
rect 32203 11906 32213 11911
rect 32308 11906 32314 12011
rect -310 11852 -206 11858
rect -866 11786 -762 11792
rect -310 11753 -305 11758
rect -211 11753 -206 11758
rect -310 11748 -206 11753
rect -866 11687 -861 11692
rect -767 11687 -762 11692
rect -866 11682 -762 11687
rect 29126 6464 29224 6478
rect 29126 6400 29148 6464
rect 29212 6400 29224 6464
rect 29126 6380 29224 6400
rect 29980 5958 30056 6018
rect 29980 5894 29988 5958
rect 30052 5894 30056 5958
rect 29980 5888 30056 5894
rect -874 755 -770 760
rect -874 750 -869 755
rect -775 750 -770 755
rect -874 650 -770 656
rect -312 755 -208 760
rect -312 750 -307 755
rect -213 750 -208 755
rect -312 650 -208 656
rect 31951 100 32056 106
rect 31951 0 31956 5
rect 32051 0 32056 5
rect 31951 -5 32056 0
rect 31393 -39 31498 -33
rect 31393 -139 31398 -134
rect 31493 -139 31498 -134
rect 31393 -144 31498 -139
<< via3 >>
rect 31323 12167 31418 12172
rect 31323 12072 31413 12167
rect 31413 12072 31418 12167
rect 31323 12067 31418 12072
rect 32213 12006 32308 12011
rect 32213 11911 32303 12006
rect 32303 11911 32308 12006
rect 32213 11906 32308 11911
rect -310 11847 -206 11852
rect -866 11781 -762 11786
rect -866 11692 -861 11781
rect -861 11692 -767 11781
rect -767 11692 -762 11781
rect -310 11758 -305 11847
rect -305 11758 -211 11847
rect -211 11758 -206 11847
rect 29148 6460 29212 6464
rect 29148 6404 29152 6460
rect 29152 6404 29208 6460
rect 29208 6404 29212 6460
rect 29148 6400 29212 6404
rect 29988 5954 30052 5958
rect 29988 5898 29992 5954
rect 29992 5898 30048 5954
rect 30048 5898 30052 5954
rect 29988 5894 30052 5898
rect -874 661 -869 750
rect -869 661 -775 750
rect -775 661 -770 750
rect -874 656 -770 661
rect -312 661 -307 750
rect -307 661 -213 750
rect -213 661 -208 750
rect -312 656 -208 661
rect 31951 95 32056 100
rect 31951 5 31956 95
rect 31956 5 32051 95
rect 32051 5 32056 95
rect 31393 -44 31498 -39
rect 31393 -134 31398 -44
rect 31398 -134 31493 -44
rect 31493 -134 31498 -44
<< metal4 >>
rect -934 12706 -694 17670
rect -934 11786 -694 12386
rect -934 11692 -866 11786
rect -762 11692 -694 11786
rect -934 750 -694 11692
rect -934 656 -874 750
rect -770 656 -694 750
rect -934 -320 -694 656
rect -370 11852 -130 15054
rect 31252 12172 31492 15094
rect 32138 12744 32378 17660
rect 31252 12067 31323 12172
rect 31418 12067 31492 12172
rect 31252 12046 31492 12067
rect -370 11758 -310 11852
rect -206 11758 -130 11852
rect 32138 12011 32378 12424
rect 32138 11906 32213 12011
rect 32308 11906 32378 12011
rect 32138 11850 32378 11906
rect -370 750 -130 11758
rect 29147 6464 29213 6465
rect 29147 6400 29148 6464
rect 29212 6400 29213 6464
rect 29147 6399 29213 6400
rect 26536 6098 26596 6386
rect 29150 6098 29210 6399
rect 26536 6038 29212 6098
rect 29987 5958 30053 5959
rect 29987 5956 29988 5958
rect 26536 5896 29988 5956
rect 26536 5620 26596 5896
rect 29987 5894 29988 5896
rect 30052 5894 30053 5958
rect 29987 5893 30053 5894
rect -370 656 -312 750
rect -208 656 -130 750
rect -974 -5462 -654 -640
rect -370 -2904 -130 656
rect 31890 100 32130 176
rect 31890 5 31951 100
rect 32056 5 32130 100
rect 31338 -39 31578 2
rect 31338 -134 31393 -39
rect 31498 -134 31578 -39
rect 31338 -2960 31578 -134
rect 31890 -368 32130 5
rect 31890 -5532 32130 -688
<< via4 >>
rect -974 17670 -654 17990
rect 32098 17660 32418 17980
rect -410 15054 -90 15374
rect 31212 15094 31532 15414
rect -974 12386 -654 12706
rect 32098 12424 32418 12744
rect -974 -640 -654 -320
rect -410 -3224 -90 -2904
rect 31850 -688 32170 -368
rect 31298 -3280 31618 -2960
rect -974 -5782 -654 -5462
rect 31850 -5852 32170 -5532
<< metal5 >>
rect -1257 17990 32567 18180
rect -1257 17670 -974 17990
rect -654 17980 32567 17990
rect -654 17670 32098 17980
rect -1257 17660 32098 17670
rect 32418 17660 32567 17980
rect -1257 17518 32567 17660
rect -591 15414 31685 15558
rect -591 15374 31212 15414
rect -591 15054 -410 15374
rect -90 15094 31212 15374
rect 31532 15094 31685 15414
rect -90 15054 31685 15094
rect -591 14896 31685 15054
rect -1143 12744 32607 12928
rect -1143 12706 32098 12744
rect -1143 12386 -974 12706
rect -654 12424 32098 12706
rect 32418 12424 32607 12744
rect -654 12386 32607 12424
rect -1143 12266 32607 12386
rect -1097 -320 32251 -182
rect -1097 -640 -974 -320
rect -654 -368 32251 -320
rect -654 -640 31850 -368
rect -1097 -688 31850 -640
rect 32170 -688 32251 -368
rect -1097 -844 32251 -688
rect -526 -2904 31651 -2758
rect -526 -3224 -410 -2904
rect -90 -2960 31651 -2904
rect -90 -3224 31298 -2960
rect -526 -3280 31298 -3224
rect 31618 -3280 31651 -2960
rect -526 -3420 31651 -3280
rect -1139 -5462 32313 -5320
rect -1139 -5782 -974 -5462
rect -654 -5532 32313 -5462
rect -654 -5782 31850 -5532
rect -1139 -5852 31850 -5782
rect 32170 -5852 32313 -5532
rect -1139 -5982 32313 -5852
use comparator  comparator_0 comparator
timestamp 1697741630
transform 0 1 30094 1 0 4665
box -1805 -1948 4495 3006
use dac  dac_0 dac
timestamp 1697762684
transform 1 0 280 0 -1 11984
box -280 -22 28705 5880
use dac  dac_1
timestamp 1697762684
transform 1 0 280 0 1 22
box -280 -22 28705 5880
use latch  latch_0 latch
timestamp 1697130564
transform 0 1 33111 -1 0 7322
box 0 -41 2306 1348
use vpp_cap  vpp_cap_0
timestamp 1697748102
transform 1 0 28848 0 1 -2942
box 4 4 2286 2342
use vpp_cap  vpp_cap_1
timestamp 1697748102
transform 1 0 28854 0 -1 -3254
box 4 4 2286 2342
use vpp_cap  vpp_cap_2
timestamp 1697748102
transform 1 0 26230 0 1 -2942
box 4 4 2286 2342
use vpp_cap  vpp_cap_3
timestamp 1697748102
transform 1 0 26236 0 -1 -3254
box 4 4 2286 2342
use vpp_cap  vpp_cap_4
timestamp 1697748102
transform 1 0 23618 0 -1 -3258
box 4 4 2286 2342
use vpp_cap  vpp_cap_5
timestamp 1697748102
transform 1 0 23612 0 1 -2938
box 4 4 2286 2342
use vpp_cap  vpp_cap_6
timestamp 1697748102
transform 1 0 20994 0 1 -2938
box 4 4 2286 2342
use vpp_cap  vpp_cap_7
timestamp 1697748102
transform 1 0 21000 0 -1 -3258
box 4 4 2286 2342
use vpp_cap  vpp_cap_8
timestamp 1697748102
transform 1 0 5300 0 -1 -3262
box 4 4 2286 2342
use vpp_cap  vpp_cap_9
timestamp 1697748102
transform 1 0 7918 0 -1 -3262
box 4 4 2286 2342
use vpp_cap  vpp_cap_10
timestamp 1697748102
transform 1 0 64 0 -1 -3266
box 4 4 2286 2342
use vpp_cap  vpp_cap_11
timestamp 1697748102
transform 1 0 2682 0 -1 -3266
box 4 4 2286 2342
use vpp_cap  vpp_cap_12
timestamp 1697748102
transform 1 0 5294 0 1 -2934
box 4 4 2286 2342
use vpp_cap  vpp_cap_13
timestamp 1697748102
transform 1 0 7912 0 1 -2934
box 4 4 2286 2342
use vpp_cap  vpp_cap_14
timestamp 1697748102
transform 1 0 58 0 1 -2930
box 4 4 2286 2342
use vpp_cap  vpp_cap_15
timestamp 1697748102
transform 1 0 2676 0 1 -2930
box 4 4 2286 2342
use vpp_cap  vpp_cap_16
timestamp 1697748102
transform 1 0 10528 0 -1 -3262
box 4 4 2286 2342
use vpp_cap  vpp_cap_17
timestamp 1697748102
transform 1 0 13146 0 -1 -3262
box 4 4 2286 2342
use vpp_cap  vpp_cap_18
timestamp 1697748102
transform 1 0 15764 0 -1 -3258
box 4 4 2286 2342
use vpp_cap  vpp_cap_19
timestamp 1697748102
transform 1 0 18382 0 -1 -3258
box 4 4 2286 2342
use vpp_cap  vpp_cap_20
timestamp 1697748102
transform 1 0 10522 0 1 -2934
box 4 4 2286 2342
use vpp_cap  vpp_cap_21
timestamp 1697748102
transform 1 0 13140 0 1 -2934
box 4 4 2286 2342
use vpp_cap  vpp_cap_22
timestamp 1697748102
transform 1 0 15758 0 1 -2938
box 4 4 2286 2342
use vpp_cap  vpp_cap_23
timestamp 1697748102
transform 1 0 18376 0 1 -2938
box 4 4 2286 2342
use vpp_cap  vpp_cap_24
timestamp 1697748102
transform 1 0 10440 0 -1 15066
box 4 4 2286 2342
use vpp_cap  vpp_cap_25
timestamp 1697748102
transform 1 0 7830 0 -1 15066
box 4 4 2286 2342
use vpp_cap  vpp_cap_26
timestamp 1697748102
transform 1 0 5212 0 -1 15066
box 4 4 2286 2342
use vpp_cap  vpp_cap_27
timestamp 1697748102
transform 1 0 2594 0 -1 15062
box 4 4 2286 2342
use vpp_cap  vpp_cap_28
timestamp 1697748102
transform 1 0 -24 0 -1 15062
box 4 4 2286 2342
use vpp_cap  vpp_cap_29
timestamp 1697748102
transform 1 0 28766 0 -1 15074
box 4 4 2286 2342
use vpp_cap  vpp_cap_30
timestamp 1697748102
transform 1 0 26148 0 -1 15074
box 4 4 2286 2342
use vpp_cap  vpp_cap_31
timestamp 1697748102
transform 1 0 23530 0 -1 15070
box 4 4 2286 2342
use vpp_cap  vpp_cap_32
timestamp 1697748102
transform 1 0 20912 0 -1 15070
box 4 4 2286 2342
use vpp_cap  vpp_cap_33
timestamp 1697748102
transform 1 0 18294 0 -1 15070
box 4 4 2286 2342
use vpp_cap  vpp_cap_34
timestamp 1697748102
transform 1 0 15676 0 -1 15070
box 4 4 2286 2342
use vpp_cap  vpp_cap_35
timestamp 1697748102
transform 1 0 13058 0 -1 15066
box 4 4 2286 2342
use vpp_cap  vpp_cap_36
timestamp 1697748102
transform 1 0 10434 0 1 15394
box 4 4 2286 2342
use vpp_cap  vpp_cap_37
timestamp 1697748102
transform 1 0 7824 0 1 15394
box 4 4 2286 2342
use vpp_cap  vpp_cap_38
timestamp 1697748102
transform 1 0 5206 0 1 15394
box 4 4 2286 2342
use vpp_cap  vpp_cap_39
timestamp 1697748102
transform 1 0 2588 0 1 15398
box 4 4 2286 2342
use vpp_cap  vpp_cap_40
timestamp 1697748102
transform 1 0 -30 0 1 15398
box 4 4 2286 2342
use vpp_cap  vpp_cap_41
timestamp 1697748102
transform 1 0 28760 0 1 15386
box 4 4 2286 2342
use vpp_cap  vpp_cap_42
timestamp 1697748102
transform 1 0 26142 0 1 15386
box 4 4 2286 2342
use vpp_cap  vpp_cap_43
timestamp 1697748102
transform 1 0 23524 0 1 15390
box 4 4 2286 2342
use vpp_cap  vpp_cap_44
timestamp 1697748102
transform 1 0 20906 0 1 15390
box 4 4 2286 2342
use vpp_cap  vpp_cap_45
timestamp 1697748102
transform 1 0 18288 0 1 15390
box 4 4 2286 2342
use vpp_cap  vpp_cap_46
timestamp 1697748102
transform 1 0 15670 0 1 15390
box 4 4 2286 2342
use vpp_cap  vpp_cap_47
timestamp 1697748102
transform 1 0 13052 0 1 15394
box 4 4 2286 2342
<< labels >>
flabel metal1 34442 6139 34502 6199 0 FreeSans 1280 0 0 0 comp
port 30 nsew
flabel metal2 34448 7460 34476 7488 0 FreeSans 1280 0 0 0 clkc
port 31 nsew
flabel metal4 -370 750 -130 11758 0 FreeSans 1280 90 0 0 avss
port 33 nsew
flabel metal4 -934 750 -694 11692 0 FreeSans 1280 90 0 0 avdd
port 32 nsew
flabel metal1 -1106 8526 -1070 8562 0 FreeSans 1280 0 0 0 vinp
port 27 nsew
flabel metal1 -1072 3444 -1036 3480 0 FreeSans 1280 0 0 0 vinn
port 28 nsew
flabel metal2 28999 9473 29033 9507 0 FreeSans 1280 0 0 0 ctlp7
port 1 nsew
flabel metal2 29005 9747 29039 9781 0 FreeSans 1280 0 0 0 ctlp6
port 2 nsew
flabel metal2 29013 10022 29047 10056 0 FreeSans 1280 0 0 0 ctlp5
port 3 nsew
flabel metal2 29011 10298 29045 10332 0 FreeSans 1280 0 0 0 ctlp4
port 4 nsew
flabel metal2 29011 10573 29045 10607 0 FreeSans 1280 0 0 0 ctlp3
port 5 nsew
flabel metal2 29011 10847 29045 10881 0 FreeSans 1280 0 0 0 ctlp2
port 6 nsew
flabel metal2 29011 11124 29045 11158 0 FreeSans 1280 0 0 0 ctlp1
port 7 nsew
flabel metal2 29013 11395 29047 11429 0 FreeSans 1280 0 0 0 ctlp0
port 8 nsew
flabel metal2 28999 577 29033 611 0 FreeSans 1280 0 0 0 ctln0
port 16 nsew
flabel metal2 28995 848 29029 882 0 FreeSans 1280 0 0 0 ctln1
port 15 nsew
flabel metal2 28997 1125 29031 1159 0 FreeSans 1280 0 0 0 ctln2
port 14 nsew
flabel metal2 29003 1399 29037 1433 0 FreeSans 1280 0 0 0 ctln3
port 13 nsew
flabel metal2 29007 1674 29041 1708 0 FreeSans 1280 0 0 0 ctln4
port 12 nsew
flabel metal2 29009 1950 29043 1984 0 FreeSans 1280 0 0 0 ctln5
port 11 nsew
flabel metal2 29009 2225 29043 2259 0 FreeSans 1280 0 0 0 ctln6
port 10 nsew
flabel metal2 29009 2499 29043 2533 0 FreeSans 1280 0 0 0 ctln7
port 9 nsew
flabel metal1 29467 2727 29513 3014 0 FreeSans 1280 90 0 0 trim4
port 17 nsew
flabel metal1 30709 2712 30753 3014 0 FreeSans 1280 90 0 0 trim3
port 18 nsew
flabel metal1 31797 2721 31843 3018 0 FreeSans 1280 90 0 0 trim2
port 19 nsew
flabel metal1 32316 2718 32360 3023 0 FreeSans 1280 90 0 0 trim1
port 20 nsew
flabel metal1 33050 2701 33100 2751 0 FreeSans 1280 90 0 0 trim0
port 21 nsew
flabel metal1 33027 9186 33077 9236 0 FreeSans 1280 90 0 0 trimb0
port 26 nsew
flabel metal1 32293 9192 32337 9236 0 FreeSans 1280 90 0 0 trimb1
port 25 nsew
flabel metal1 31774 9190 31820 9236 0 FreeSans 1280 90 0 0 trimb2
port 24 nsew
flabel metal1 30686 9192 30730 9236 0 FreeSans 1280 90 0 0 trimb3
port 23 nsew
flabel metal1 29444 9190 29490 9236 0 FreeSans 1280 90 0 0 trimb4
port 22 nsew
flabel metal2 48 1528 89 10480 0 FreeSans 1280 90 0 0 sample
port 29 nsew
<< end >>
