magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 1142 542
<< pwell >>
rect 1 -19 1103 143
rect 29 -57 63 -19
<< scnmos >>
rect 79 7 1025 117
<< scpmoshvt >>
rect 79 283 1025 457
<< ndiff >>
rect 27 72 79 117
rect 27 38 35 72
rect 69 38 79 72
rect 27 7 79 38
rect 1025 72 1077 117
rect 1025 38 1035 72
rect 1069 38 1077 72
rect 1025 7 1077 38
<< pdiff >>
rect 27 445 79 457
rect 27 411 35 445
rect 69 411 79 445
rect 27 343 79 411
rect 27 309 35 343
rect 69 309 79 343
rect 27 283 79 309
rect 1025 445 1077 457
rect 1025 411 1035 445
rect 1069 411 1077 445
rect 1025 343 1077 411
rect 1025 309 1035 343
rect 1069 309 1077 343
rect 1025 283 1077 309
<< ndiffc >>
rect 35 38 69 72
rect 1035 38 1069 72
<< pdiffc >>
rect 35 411 69 445
rect 35 309 69 343
rect 1035 411 1069 445
rect 1035 309 1069 343
<< poly >>
rect 79 457 1025 483
rect 79 257 1025 283
rect 79 235 529 257
rect 79 201 95 235
rect 129 201 223 235
rect 257 201 351 235
rect 385 201 479 235
rect 513 201 529 235
rect 79 185 529 201
rect 571 199 1025 215
rect 571 165 587 199
rect 621 165 715 199
rect 749 165 843 199
rect 877 165 971 199
rect 1005 165 1025 199
rect 571 143 1025 165
rect 79 117 1025 143
rect 79 -19 1025 7
<< polycont >>
rect 95 201 129 235
rect 223 201 257 235
rect 351 201 385 235
rect 479 201 513 235
rect 587 165 621 199
rect 715 165 749 199
rect 843 165 877 199
rect 971 165 1005 199
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1104 521
rect 17 445 1086 487
rect 17 411 35 445
rect 69 411 1035 445
rect 1069 411 1086 445
rect 17 343 1086 411
rect 17 309 35 343
rect 69 309 1035 343
rect 1069 309 1086 343
rect 17 269 1086 309
rect 17 201 95 235
rect 129 201 223 235
rect 257 201 351 235
rect 385 201 479 235
rect 513 201 533 235
rect 17 131 533 201
rect 567 199 1086 269
rect 567 165 587 199
rect 621 165 715 199
rect 749 165 843 199
rect 877 165 971 199
rect 1005 165 1086 199
rect 17 72 1086 131
rect 17 38 35 72
rect 69 38 1035 72
rect 1069 38 1086 72
rect 17 -23 1086 38
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1104 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 857 487 891 521
rect 949 487 983 521
rect 1041 487 1075 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
rect 857 -57 891 -23
rect 949 -57 983 -23
rect 1041 -57 1075 -23
<< metal1 >>
rect 0 521 1104 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1104 521
rect 0 456 1104 487
rect 0 -23 1104 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1104 -23
rect 0 -88 1104 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 decap_12
flabel metal1 s 29 -57 63 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 29 487 63 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 29 487 63 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 29 -57 63 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
<< properties >>
string FIXED_BBOX 0 -40 1104 504
string path 0.000 -1.000 27.600 -1.000 
<< end >>
