magic
tech sky130B
magscale 1 2
timestamp 1696032376
<< metal1 >>
rect 9 3051 499 3081
rect 1755 3051 4279 3081
rect 15 110 45 3051
rect 997 2301 1191 2331
rect 200 1790 207 1800
rect 237 1699 267 1816
rect 2511 1699 2541 1825
rect 3675 1699 3705 1819
rect 4255 1699 4285 1805
rect 4934 1699 4964 3118
rect 5190 1800 5302 1812
rect 5190 1740 5210 1800
rect 5280 1740 5302 1800
rect 5190 1728 5302 1740
rect 237 1669 4964 1699
rect 5190 1680 5300 1692
rect 237 1357 267 1669
rect 5190 1620 5210 1680
rect 5280 1620 5300 1680
rect 5190 1610 5300 1620
rect 5190 1570 5300 1580
rect 5190 1510 5210 1570
rect 5280 1510 5300 1570
rect 5190 1498 5300 1510
rect 5190 1460 5300 1470
rect 5190 1400 5210 1460
rect 5280 1400 5300 1460
rect 5190 1390 5300 1400
rect 5190 1340 5300 1350
rect 5190 1280 5210 1340
rect 5280 1280 5300 1340
rect 5190 1270 5300 1280
rect 15 80 265 110
<< via1 >>
rect 5210 1740 5280 1800
rect 5210 1620 5280 1680
rect 5210 1510 5280 1570
rect 5210 1400 5280 1460
rect 5210 1280 5280 1340
<< metal2 >>
rect 377 1457 411 1880
rect 2676 1562 2710 1884
rect 3835 1669 3869 1870
rect 4398 1850 4448 1887
rect 4390 1844 4450 1850
rect 4398 1787 4448 1844
rect 5190 1800 5302 1812
rect 5190 1787 5210 1800
rect 4398 1753 5210 1787
rect 4722 1750 4756 1753
rect 5190 1740 5210 1753
rect 5280 1740 5302 1800
rect 5190 1728 5302 1740
rect 5190 1680 5300 1692
rect 5190 1669 5210 1680
rect 3833 1635 5210 1669
rect 4719 1632 4753 1635
rect 5190 1620 5210 1635
rect 5280 1620 5300 1680
rect 5190 1610 5300 1620
rect 5190 1570 5300 1580
rect 4719 1562 4753 1564
rect 5190 1562 5210 1570
rect 2676 1528 5210 1562
rect 4719 1525 4753 1528
rect 5190 1510 5210 1528
rect 5280 1510 5300 1570
rect 5190 1498 5300 1510
rect 5190 1460 5300 1470
rect 5190 1457 5210 1460
rect 377 1423 5210 1457
rect 4719 1422 4753 1423
rect 5190 1400 5210 1423
rect 5280 1400 5300 1460
rect 5190 1390 5300 1400
rect 4719 1340 4753 1341
rect 5190 1340 5300 1350
rect 414 1306 5210 1340
rect 5190 1280 5210 1306
rect 5280 1280 5300 1340
rect 5190 1270 5300 1280
use nfet_2mimcap_combo  nfet_2mimcap_combo_0
timestamp 1696029511
transform 1 0 2290 0 1 1782
box 0 0 1046 1330
use nfet_4mimcap_combo  nfet_4mimcap_combo_0
timestamp 1696029615
transform 1 0 -10 0 1 1780
box 0 0 2196 1334
use nfet_8mimcap_combo  nfet_8mimcap_combo_0
timestamp 1696029713
transform 1 0 0 0 -1 1394
box 0 0 5050 1334
use nfet_mimcap_combo  nfet_mimcap_combo_0
timestamp 1696029511
transform 1 0 4624 0 1 2274
box -604 -494 -128 836
use nfet_mimcap_combo  nfet_mimcap_combo_1
timestamp 1696029511
transform 1 0 4054 0 1 2274
box -604 -494 -128 836
<< labels >>
rlabel metal1 5300 1770 5300 1770 3 d0
port 3 e
rlabel metal1 5300 1650 5300 1650 3 d1
port 4 e
rlabel metal1 5300 1540 5300 1540 3 d2
port 5 e
rlabel metal1 5300 1430 5300 1430 3 d3
port 6 e
rlabel metal1 5300 1310 5300 1310 3 d4
port 7 e
rlabel metal1 4934 3088 4964 3118 1 VSS
port 1 n
rlabel metal1 16 1736 16 1736 7 drain
port 2 w
<< end >>
