magic
tech sky130B
magscale 1 2
timestamp 1696112986
<< metal1 >>
rect 1944 1276 5976 1304
rect 2148 520 2176 522
rect 1942 492 5974 520
rect 2148 310 2176 492
rect 2339 223 2397 283
rect 2171 177 2251 207
use sky130_fd_pr__nfet_01v8_lvt_E33R59  sky130_fd_pr__nfet_01v8_lvt_E33R59_0
timestamp 1696108744
transform 0 1 2245 -1 0 250
box -226 -279 226 279
use trimcap  trimcap_0
timestamp 1696109480
transform 1 0 1722 0 1 60
box 0 376 476 1324
use trimcap  trimcap_1
timestamp 1696109480
transform 1 0 2294 0 1 58
box 0 376 476 1324
use trimcap  trimcap_2
timestamp 1696109480
transform 1 0 4574 0 1 68
box 0 376 476 1324
use trimcap  trimcap_3
timestamp 1696109480
transform 1 0 5142 0 1 68
box 0 376 476 1324
use trimcap  trimcap_4
timestamp 1696109480
transform 1 0 5710 0 1 68
box 0 376 476 1324
use trimcap  trimcap_5
timestamp 1696109480
transform 1 0 2864 0 1 58
box 0 376 476 1324
use trimcap  trimcap_6
timestamp 1696109480
transform 1 0 3432 0 1 58
box 0 376 476 1324
use trimcap  trimcap_7
timestamp 1696109480
transform 1 0 4000 0 1 58
box 0 376 476 1324
<< labels >>
flabel metal1 1944 1276 5976 1304 0 FreeSans 480 0 0 0 todrain
flabel metal1 2339 223 2397 283 0 FreeSans 480 0 0 0 d_i
flabel metal1 2171 177 2251 207 0 FreeSans 480 0 0 0 tovss
<< end >>
