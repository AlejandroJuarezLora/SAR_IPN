magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 1142 542
<< pwell >>
rect 1 -19 1065 163
rect 30 -57 64 -19
<< scnmos >>
rect 81 7 111 137
rect 165 7 195 137
rect 353 7 383 137
rect 437 7 467 137
rect 521 7 551 137
rect 605 7 635 137
rect 705 7 735 137
rect 789 7 819 137
rect 873 7 903 137
rect 957 7 987 137
<< scpmoshvt >>
rect 81 257 111 457
rect 165 257 195 457
rect 353 257 383 457
rect 437 257 467 457
rect 521 257 551 457
rect 605 257 635 457
rect 705 257 735 457
rect 789 257 819 457
rect 873 257 903 457
rect 957 257 987 457
<< ndiff >>
rect 27 123 81 137
rect 27 89 37 123
rect 71 89 81 123
rect 27 55 81 89
rect 27 21 37 55
rect 71 21 81 55
rect 27 7 81 21
rect 111 123 165 137
rect 111 89 121 123
rect 155 89 165 123
rect 111 55 165 89
rect 111 21 121 55
rect 155 21 165 55
rect 111 7 165 21
rect 195 55 353 137
rect 195 21 205 55
rect 239 21 309 55
rect 343 21 353 55
rect 195 7 353 21
rect 383 55 437 137
rect 383 21 393 55
rect 427 21 437 55
rect 383 7 437 21
rect 467 123 521 137
rect 467 89 477 123
rect 511 89 521 123
rect 467 7 521 89
rect 551 55 605 137
rect 551 21 561 55
rect 595 21 605 55
rect 551 7 605 21
rect 635 55 705 137
rect 635 21 654 55
rect 688 21 705 55
rect 635 7 705 21
rect 735 55 789 137
rect 735 21 745 55
rect 779 21 789 55
rect 735 7 789 21
rect 819 123 873 137
rect 819 89 829 123
rect 863 89 873 123
rect 819 7 873 89
rect 903 123 957 137
rect 903 89 913 123
rect 947 89 957 123
rect 903 55 957 89
rect 903 21 913 55
rect 947 21 957 55
rect 903 7 957 21
rect 987 123 1039 137
rect 987 89 997 123
rect 1031 89 1039 123
rect 987 55 1039 89
rect 987 21 997 55
rect 1031 21 1039 55
rect 987 7 1039 21
<< pdiff >>
rect 27 443 81 457
rect 27 409 37 443
rect 71 409 81 443
rect 27 353 81 409
rect 27 319 37 353
rect 71 319 81 353
rect 27 257 81 319
rect 111 369 165 457
rect 111 335 121 369
rect 155 335 165 369
rect 111 301 165 335
rect 111 267 121 301
rect 155 267 165 301
rect 111 257 165 267
rect 195 437 247 457
rect 195 403 205 437
rect 239 403 247 437
rect 195 309 247 403
rect 195 275 205 309
rect 239 275 247 309
rect 195 257 247 275
rect 301 437 353 457
rect 301 403 309 437
rect 343 403 353 437
rect 301 257 353 403
rect 383 369 437 457
rect 383 335 393 369
rect 427 335 437 369
rect 383 257 437 335
rect 467 437 521 457
rect 467 403 477 437
rect 511 403 521 437
rect 467 257 521 403
rect 551 369 605 457
rect 551 335 561 369
rect 595 335 605 369
rect 551 257 605 335
rect 635 437 705 457
rect 635 403 653 437
rect 687 403 705 437
rect 635 367 705 403
rect 635 333 653 367
rect 687 333 705 367
rect 635 257 705 333
rect 735 437 789 457
rect 735 403 745 437
rect 779 403 789 437
rect 735 257 789 403
rect 819 437 873 457
rect 819 403 829 437
rect 863 403 873 437
rect 819 369 873 403
rect 819 335 829 369
rect 863 335 873 369
rect 819 257 873 335
rect 903 437 957 457
rect 903 403 913 437
rect 947 403 957 437
rect 903 257 957 403
rect 987 437 1044 457
rect 987 403 998 437
rect 1032 403 1044 437
rect 987 369 1044 403
rect 987 335 998 369
rect 1032 335 1044 369
rect 987 301 1044 335
rect 987 267 998 301
rect 1032 267 1044 301
rect 987 257 1044 267
<< ndiffc >>
rect 37 89 71 123
rect 37 21 71 55
rect 121 89 155 123
rect 121 21 155 55
rect 205 21 239 55
rect 309 21 343 55
rect 393 21 427 55
rect 477 89 511 123
rect 561 21 595 55
rect 654 21 688 55
rect 745 21 779 55
rect 829 89 863 123
rect 913 89 947 123
rect 913 21 947 55
rect 997 89 1031 123
rect 997 21 1031 55
<< pdiffc >>
rect 37 409 71 443
rect 37 319 71 353
rect 121 335 155 369
rect 121 267 155 301
rect 205 403 239 437
rect 205 275 239 309
rect 309 403 343 437
rect 393 335 427 369
rect 477 403 511 437
rect 561 335 595 369
rect 653 403 687 437
rect 653 333 687 367
rect 745 403 779 437
rect 829 403 863 437
rect 829 335 863 369
rect 913 403 947 437
rect 998 403 1032 437
rect 998 335 1032 369
rect 998 267 1032 301
<< poly >>
rect 81 457 111 483
rect 165 457 195 483
rect 353 457 383 483
rect 437 457 467 483
rect 521 457 551 483
rect 605 457 635 483
rect 705 457 735 483
rect 789 457 819 483
rect 873 457 903 483
rect 957 457 987 483
rect 81 225 111 257
rect 165 225 195 257
rect 353 225 383 257
rect 437 225 467 257
rect 521 225 551 257
rect 605 225 635 257
rect 705 225 735 257
rect 789 225 819 257
rect 873 225 903 257
rect 957 225 987 257
rect 22 209 195 225
rect 22 175 34 209
rect 68 175 195 209
rect 22 159 195 175
rect 341 209 395 225
rect 341 175 351 209
rect 385 175 395 209
rect 341 159 395 175
rect 437 209 551 225
rect 437 175 477 209
rect 511 175 551 209
rect 437 159 551 175
rect 593 209 647 225
rect 593 175 603 209
rect 637 175 647 209
rect 593 159 647 175
rect 693 209 747 225
rect 693 175 703 209
rect 737 175 747 209
rect 693 159 747 175
rect 789 209 903 225
rect 789 175 829 209
rect 863 175 903 209
rect 789 159 903 175
rect 945 209 999 225
rect 945 175 955 209
rect 989 175 999 209
rect 945 159 999 175
rect 81 137 111 159
rect 165 137 195 159
rect 353 137 383 159
rect 437 137 467 159
rect 521 137 551 159
rect 605 137 635 159
rect 705 137 735 159
rect 789 137 819 159
rect 873 137 903 159
rect 957 137 987 159
rect 81 -19 111 7
rect 165 -19 195 7
rect 353 -19 383 7
rect 437 -19 467 7
rect 521 -19 551 7
rect 605 -19 635 7
rect 705 -19 735 7
rect 789 -19 819 7
rect 873 -19 903 7
rect 957 -19 987 7
<< polycont >>
rect 34 175 68 209
rect 351 175 385 209
rect 477 175 511 209
rect 603 175 637 209
rect 703 175 737 209
rect 829 175 863 209
rect 955 175 989 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1104 521
rect 18 443 255 453
rect 18 409 37 443
rect 71 437 255 443
rect 71 419 205 437
rect 71 409 87 419
rect 18 353 87 409
rect 239 403 255 437
rect 18 319 37 353
rect 71 319 87 353
rect 121 369 171 385
rect 155 335 171 369
rect 121 301 171 335
rect 18 209 84 283
rect 18 175 34 209
rect 68 175 84 209
rect 155 267 171 301
rect 121 141 171 267
rect 205 351 255 403
rect 301 437 695 453
rect 301 403 309 437
rect 343 419 477 437
rect 343 403 351 419
rect 301 385 351 403
rect 469 403 477 419
rect 511 419 653 437
rect 511 403 519 419
rect 469 385 519 403
rect 645 403 653 419
rect 687 403 695 437
rect 385 369 435 385
rect 385 351 393 369
rect 205 335 393 351
rect 427 351 435 369
rect 553 369 603 385
rect 553 351 561 369
rect 427 335 561 351
rect 595 335 603 369
rect 205 317 603 335
rect 645 367 695 403
rect 737 437 787 487
rect 737 403 745 437
rect 779 403 787 437
rect 737 385 787 403
rect 821 437 871 453
rect 821 403 829 437
rect 863 403 871 437
rect 645 333 653 367
rect 687 351 695 367
rect 821 369 871 403
rect 905 437 955 487
rect 905 403 913 437
rect 947 403 955 437
rect 905 385 955 403
rect 998 437 1039 453
rect 1032 403 1039 437
rect 821 351 829 369
rect 687 335 829 351
rect 863 351 871 369
rect 998 369 1039 403
rect 863 335 998 351
rect 1032 335 1039 369
rect 687 333 1039 335
rect 645 317 1039 333
rect 205 309 255 317
rect 239 275 255 309
rect 998 301 1039 317
rect 205 259 255 275
rect 301 249 653 283
rect 301 209 408 249
rect 301 175 351 209
rect 385 175 408 209
rect 442 209 553 215
rect 442 175 477 209
rect 511 175 553 209
rect 587 209 653 249
rect 587 175 603 209
rect 637 175 653 209
rect 687 249 964 283
rect 1032 267 1039 301
rect 998 251 1039 267
rect 687 209 753 249
rect 930 215 964 249
rect 687 175 703 209
rect 737 175 753 209
rect 797 209 896 215
rect 797 175 829 209
rect 863 175 896 209
rect 930 209 1087 215
rect 930 175 955 209
rect 989 175 1087 209
rect 21 123 71 139
rect 121 133 879 141
rect 21 89 37 123
rect 21 55 71 89
rect 21 21 37 55
rect 105 123 879 133
rect 105 89 121 123
rect 155 105 477 123
rect 155 89 171 105
rect 457 89 477 105
rect 511 105 829 123
rect 511 89 527 105
rect 813 89 829 105
rect 863 89 879 123
rect 913 123 963 141
rect 947 89 963 123
rect 105 55 171 89
rect 105 21 121 55
rect 155 21 171 55
rect 205 55 343 71
rect 654 55 688 71
rect 913 55 963 89
rect 239 21 309 55
rect 21 -23 71 21
rect 205 -23 343 21
rect 377 21 393 55
rect 427 21 561 55
rect 595 21 611 55
rect 377 11 611 21
rect 654 -23 688 21
rect 729 21 745 55
rect 779 21 913 55
rect 947 21 963 55
rect 729 11 963 21
rect 997 123 1031 141
rect 997 55 1031 89
rect 997 -23 1031 21
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1104 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 765 487 799 521
rect 857 487 891 521
rect 949 487 983 521
rect 1041 487 1075 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
rect 765 -57 799 -23
rect 857 -57 891 -23
rect 949 -57 983 -23
rect 1041 -57 1075 -23
<< metal1 >>
rect 0 521 1104 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 765 521
rect 799 487 857 521
rect 891 487 949 521
rect 983 487 1041 521
rect 1075 487 1104 521
rect 0 456 1104 487
rect 0 -23 1104 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 765 -23
rect 799 -57 857 -23
rect 891 -57 949 -23
rect 983 -57 1041 -23
rect 1075 -57 1104 -23
rect 0 -88 1104 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 a221oi_2
flabel metal1 s 30 -57 64 -23 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 30 487 64 521 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 30 487 64 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 30 -57 64 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 310 249 344 283 0 FreeSans 400 0 0 0 B2
port 10 nsew
flabel locali s 30 181 64 215 0 FreeSans 400 0 0 0 C1
port 13 nsew
flabel locali s 1046 181 1080 215 0 FreeSans 400 180 0 0 A2
port 7 nsew
flabel locali s 862 181 896 215 0 FreeSans 400 180 0 0 A1
port 8 nsew
flabel locali s 494 181 528 215 0 FreeSans 400 0 0 0 B1
port 9 nsew
flabel locali s 310 181 344 215 0 FreeSans 400 0 0 0 B2
port 10 nsew
flabel locali s 122 181 156 215 0 FreeSans 400 0 0 0 Y
port 12 nsew
flabel locali s 30 249 64 283 0 FreeSans 400 0 0 0 C1
port 13 nsew
<< properties >>
string FIXED_BBOX 0 -40 1104 504
string path 0.000 -1.000 27.600 -1.000 
<< end >>
