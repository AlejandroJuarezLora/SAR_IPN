* SPICE3 file created from latch.ext - technology: sky130B

.subckt M2_1 a_n98_n109# a_n40_n197# a_40_n109# VSUBS
X0 a_40_n109# a_n40_n197# a_n98_n109# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
C0 a_40_n109# a_n40_n197# 0.0145f
C1 a_n98_n109# a_40_n109# 0.104f
C2 a_n98_n109# a_n40_n197# 0.0145f
C3 a_40_n109# VSUBS 0.122f
C4 a_n98_n109# VSUBS 0.122f
C5 a_n40_n197# VSUBS 0.259f
.ends

.subckt M2_inv a_n40_n201# a_40_n104# w_n236_n324# a_n98_n104# VSUBS
X0 a_40_n104# a_n40_n201# a_n98_n104# w_n236_n324# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
C0 a_40_n104# a_n40_n201# 0.0145f
C1 a_40_n104# w_n236_n324# 0.0219f
C2 w_n236_n324# a_n40_n201# 0.12f
C3 a_40_n104# a_n98_n104# 0.104f
C4 a_n40_n201# a_n98_n104# 0.0145f
C5 w_n236_n324# a_n98_n104# 0.0219f
C6 a_40_n104# VSUBS 0.1f
C7 a_n98_n104# VSUBS 0.1f
C8 a_n40_n201# VSUBS 0.146f
C9 w_n236_n324# VSUBS 0.804f
.ends

.subckt M1_inv a_40_n171# a_n40_n197# a_n98_n171# VSUBS
X0 a_40_n171# a_n40_n197# a_n98_n171# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
C0 a_40_n171# a_n98_n171# 0.104f
C1 a_40_n171# a_n40_n197# 0.0145f
C2 a_n40_n197# a_n98_n171# 0.0145f
C3 a_40_n171# VSUBS 0.122f
C4 a_n98_n171# VSUBS 0.122f
C5 a_n40_n197# VSUBS 0.259f
.ends

.subckt inv_lvt M2_inv_0/a_n98_n104# M2_inv_0/w_n236_n324# M1_inv_0/a_n98_n171# m1_170_505#
+ m2_289_257# VSUBS
XM2_inv_0 m1_170_505# m2_289_257# M2_inv_0/w_n236_n324# M2_inv_0/a_n98_n104# VSUBS
+ M2_inv
XM1_inv_0 m2_289_257# m1_170_505# M1_inv_0/a_n98_n171# VSUBS M1_inv
C0 M2_inv_0/a_n98_n104# m1_170_505# 0.0037f
C1 M2_inv_0/a_n98_n104# M2_inv_0/w_n236_n324# -1.52e-20
C2 M2_inv_0/w_n236_n324# m1_170_505# 0.0237f
C3 m2_289_257# M2_inv_0/a_n98_n104# 0.00406f
C4 m2_289_257# m1_170_505# 0.086f
C5 m2_289_257# M2_inv_0/w_n236_n324# 0.046f
C6 M2_inv_0/a_n98_n104# M1_inv_0/a_n98_n171# 0.00387f
C7 M1_inv_0/a_n98_n171# m1_170_505# 0.00383f
C8 M2_inv_0/w_n236_n324# M1_inv_0/a_n98_n171# 0.00225f
C9 m2_289_257# M1_inv_0/a_n98_n171# 0.00406f
C10 m2_289_257# VSUBS 0.547f
C11 M1_inv_0/a_n98_n171# VSUBS 0.122f
C12 M2_inv_0/a_n98_n104# VSUBS 0.1f
C13 m1_170_505# VSUBS 0.453f
C14 M2_inv_0/w_n236_n324# VSUBS 0.804f
.ends

.subckt M1_2 a_n98_n109# a_n40_n197# a_40_n109# VSUBS
X0 a_40_n109# a_n40_n197# a_n98_n109# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.4
C0 a_40_n109# a_n40_n197# 0.0145f
C1 a_40_n109# a_n98_n109# 0.104f
C2 a_n98_n109# a_n40_n197# 0.0145f
C3 a_40_n109# VSUBS 0.122f
C4 a_n98_n109# VSUBS 0.122f
C5 a_n40_n197# VSUBS 0.259f
.ends

.subckt latch vdd vss Qn S R Q
XM2_1_0 vss m1_1673_493# Q vss M2_1
Xinv_lvt_0 vdd vdd vss R m1_1673_493# vss inv_lvt
Xinv_lvt_1 vdd vdd vss S m1_458_623# vss inv_lvt
Xinv_lvt_2 vdd vdd vss Qn Q vss inv_lvt
Xinv_lvt_3 vdd vdd vss Q Qn vss inv_lvt
XM1_2_0 Qn m1_458_623# vss vss M1_2
X0 Q Qn.t0 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X1 Qn Q.t1 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X2 m1_1673_493# R.t1 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X3 m1_458_623# S.t1 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X4 Q Qn.t1 vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X5 Qn Q.t0 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X6 m1_1673_493# R.t0 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
X7 m1_458_623# S.t0 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=0 l=0
R0 vss.n33 vss.n32 403.438
R1 vss.n147 vss.n146 403.438
R2 vss.n35 vss.n34 394
R3 vss.n151 vss.n148 394
R4 vss.n286 vss.n285 371.921
R5 vss.n244 vss.n243 359.312
R6 vss.n208 vss.n207 346.705
R7 vss.n55 vss.n51 334.098
R8 vss.n10 vss.n6 334.098
R9 vss.n128 vss.n127 334.098
R10 vss.n171 vss.n170 334.098
R11 vss.n313 vss.n312 334.098
R12 vss.n83 vss.n82 292.5
R13 vss.n81 vss.n80 292.5
R14 vss.n77 vss.n76 292.5
R15 vss.n75 vss.n74 292.5
R16 vss.n73 vss.n72 292.5
R17 vss.n71 vss.n70 292.5
R18 vss.n69 vss.n68 292.5
R19 vss.n51 vss.n50 292.5
R20 vss.n54 vss.n53 292.5
R21 vss.n36 vss.n35 292.5
R22 vss.n6 vss.n5 292.5
R23 vss.n9 vss.n8 292.5
R24 vss.n124 vss.n123 292.5
R25 vss.n125 vss.n124 292.5
R26 vss.n127 vss.n126 292.5
R27 vss.n151 vss.n150 292.5
R28 vss.n152 vss.n151 292.5
R29 vss.n167 vss.n166 292.5
R30 vss.n168 vss.n167 292.5
R31 vss.n170 vss.n169 292.5
R32 vss.n188 vss.n187 292.5
R33 vss.n189 vss.n188 292.5
R34 vss.n205 vss.n204 292.5
R35 vss.n207 vss.n206 292.5
R36 vss.n226 vss.n225 292.5
R37 vss.n241 vss.n240 292.5
R38 vss.n243 vss.n242 292.5
R39 vss.n262 vss.n261 292.5
R40 vss.n283 vss.n282 292.5
R41 vss.n285 vss.n284 292.5
R42 vss.n301 vss.n300 292.5
R43 vss.n303 vss.n302 292.5
R44 vss.n306 vss.n305 292.5
R45 vss.n305 vss.n304 292.5
R46 vss.n309 vss.n308 292.5
R47 vss.n311 vss.n310 292.5
R48 vss.n316 vss.n315 292.5
R49 vss.n319 vss.n318 292.5
R50 vss.n318 vss.n317 292.5
R51 vss.n322 vss.n321 292.5
R52 vss.n321 vss.n320 292.5
R53 vss.n324 vss.n323 292.5
R54 vss.n251 vss.n250 292.5
R55 vss.n137 vss.n136 292.5
R56 vss.n25 vss.n24 292.5
R57 vss.n23 vss.n22 292.5
R58 vss.n139 vss.n138 292.5
R59 vss.n178 vss.n177 292.5
R60 vss.n216 vss.n215 292.5
R61 vss.n97 vss.n96 292.5
R62 vss.n95 vss.n94 292.5
R63 vss.n94 vss.n93 292.5
R64 vss.n92 vss.n91 292.5
R65 vss.n91 vss.n90 292.5
R66 vss.n89 vss.n88 292.5
R67 vss.n88 vss.n87 292.5
R68 vss.n86 vss.n85 292.5
R69 vss.n85 vss.n84 292.5
R70 vss.n77 vss.n75 156.236
R71 vss.n319 vss.n316 156.236
R72 vss.n86 vss.n83 144.189
R73 vss.n309 vss.n306 142.683
R74 vss.n314 vss.n313 134.577
R75 vss.n80 vss.n79 117.719
R76 vss.n55 vss.n54 94.5564
R77 vss.n10 vss.n9 94.5564
R78 vss.n128 vss.n125 94.5564
R79 vss.n171 vss.n168 94.5564
R80 vss.n308 vss.n307 90.6381
R81 vss.n315 vss.n314 90.6381
R82 vss.n79 vss.n78 87.3925
R83 vss.n56 vss.n49 86.9123
R84 vss.n11 vss.n4 86.9123
R85 vss.n129 vss.n120 86.9123
R86 vss.n172 vss.n164 86.9123
R87 vss.n37 vss.n36 81.9489
R88 vss.n153 vss.n152 81.9489
R89 vss.n208 vss.n205 81.9489
R90 vss.n38 vss.n31 75.324
R91 vss.n154 vss.n145 75.324
R92 vss.n209 vss.n202 75.324
R93 vss.n190 vss.n189 69.3415
R94 vss.n244 vss.n241 69.3415
R95 vss.n191 vss.n184 63.7358
R96 vss.n245 vss.n238 63.7358
R97 vss.n262 vss.n260 63.0378
R98 vss.n259 vss.n258 57.9417
R99 vss.n227 vss.n226 56.734
R100 vss.n286 vss.n283 56.734
R101 vss.n228 vss.n223 52.1476
R102 vss.n287 vss.n280 52.1476
R103 vss.n226 vss.n224 50.4303
R104 vss.n283 vss.n281 50.4303
R105 vss.n223 vss.n222 46.3534
R106 vss.n280 vss.n279 46.3534
R107 vss.n263 vss.n262 44.1266
R108 vss.n264 vss.n259 40.5593
R109 vss.n189 vss.n185 37.8228
R110 vss.n241 vss.n239 37.8228
R111 vss.n184 vss.n183 34.7652
R112 vss.n238 vss.n237 34.7652
R113 vss.n81 vss.n77 25.6005
R114 vss.n83 vss.n81 25.6005
R115 vss.n75 vss.n73 25.6005
R116 vss.n73 vss.n71 25.6005
R117 vss.n71 vss.n69 25.6005
R118 vss.n69 vss.n67 25.6005
R119 vss.n67 vss.n66 25.6005
R120 vss.n66 vss.n65 25.6005
R121 vss.n65 vss.n64 25.6005
R122 vss.n64 vss.n63 25.6005
R123 vss.n63 vss.n62 25.6005
R124 vss.n123 vss.n122 25.6005
R125 vss.n150 vss.n149 25.6005
R126 vss.n187 vss.n186 25.6005
R127 vss.n293 vss.n292 25.6005
R128 vss.n294 vss.n293 25.6005
R129 vss.n295 vss.n294 25.6005
R130 vss.n296 vss.n295 25.6005
R131 vss.n297 vss.n296 25.6005
R132 vss.n298 vss.n297 25.6005
R133 vss.n299 vss.n298 25.6005
R134 vss.n301 vss.n299 25.6005
R135 vss.n303 vss.n301 25.6005
R136 vss.n306 vss.n303 25.6005
R137 vss.n311 vss.n309 25.6005
R138 vss.n316 vss.n311 25.6005
R139 vss.n89 vss.n86 25.6005
R140 vss.n92 vss.n89 25.6005
R141 vss.n95 vss.n92 25.6005
R142 vss.n97 vss.n95 25.6005
R143 vss.n324 vss.n322 25.6005
R144 vss.n322 vss.n319 25.6005
R145 vss.n36 vss.n33 25.2154
R146 vss.n152 vss.n147 25.2154
R147 vss.n205 vss.n203 25.2154
R148 vss.n31 vss.n30 23.177
R149 vss.n145 vss.n144 23.177
R150 vss.n202 vss.n201 23.177
R151 vss.n325 vss.n324 15.8123
R152 vss.n252 vss.n251 15.0593
R153 vss.n217 vss.n216 14.3064
R154 vss.n98 vss.n97 13.5534
R155 vss.n179 vss.n178 13.5534
R156 vss.n26 vss.n23 12.8005
R157 vss.n26 vss.n25 12.8005
R158 vss.n140 vss.n137 12.8005
R159 vss.n140 vss.n139 12.8005
R160 vss.n54 vss.n52 12.608
R161 vss.n9 vss.n7 12.608
R162 vss.n125 vss.n121 12.608
R163 vss.n168 vss.n165 12.608
R164 vss.n49 vss.n48 11.5887
R165 vss.n4 vss.n3 11.5887
R166 vss.n120 vss.n119 11.5887
R167 vss.n164 vss.n163 11.5887
R168 vss.n99 vss.n98 9.30167
R169 vss.n270 vss.n269 9.3005
R170 vss.n268 vss.n267 9.3005
R171 vss.n234 vss.n233 9.3005
R172 vss.n218 vss.n217 9.3005
R173 vss.n174 vss.n173 9.3005
R174 vss.n173 vss.n172 9.3005
R175 vss.n172 vss.n171 9.3005
R176 vss.n17 vss.n16 9.3005
R177 vss.n44 vss.n43 9.3005
R178 vss.n42 vss.n41 9.3005
R179 vss.n40 vss.n39 9.3005
R180 vss.n39 vss.n38 9.3005
R181 vss.n38 vss.n37 9.3005
R182 vss.n15 vss.n14 9.3005
R183 vss.n13 vss.n12 9.3005
R184 vss.n12 vss.n11 9.3005
R185 vss.n11 vss.n10 9.3005
R186 vss.n131 vss.n130 9.3005
R187 vss.n130 vss.n129 9.3005
R188 vss.n129 vss.n128 9.3005
R189 vss.n135 vss.n134 9.3005
R190 vss.n133 vss.n132 9.3005
R191 vss.n156 vss.n155 9.3005
R192 vss.n155 vss.n154 9.3005
R193 vss.n154 vss.n153 9.3005
R194 vss.n160 vss.n159 9.3005
R195 vss.n158 vss.n157 9.3005
R196 vss.n176 vss.n175 9.3005
R197 vss.n180 vss.n179 9.3005
R198 vss.n193 vss.n192 9.3005
R199 vss.n192 vss.n191 9.3005
R200 vss.n191 vss.n190 9.3005
R201 vss.n197 vss.n196 9.3005
R202 vss.n195 vss.n194 9.3005
R203 vss.n211 vss.n210 9.3005
R204 vss.n210 vss.n209 9.3005
R205 vss.n209 vss.n208 9.3005
R206 vss.n232 vss.n231 9.3005
R207 vss.n230 vss.n229 9.3005
R208 vss.n229 vss.n228 9.3005
R209 vss.n228 vss.n227 9.3005
R210 vss.n247 vss.n246 9.3005
R211 vss.n246 vss.n245 9.3005
R212 vss.n245 vss.n244 9.3005
R213 vss.n253 vss.n252 9.3005
R214 vss.n249 vss.n248 9.3005
R215 vss.n265 vss.n264 9.3005
R216 vss.n264 vss.n263 9.3005
R217 vss.n289 vss.n288 9.3005
R218 vss.n288 vss.n287 9.3005
R219 vss.n287 vss.n286 9.3005
R220 vss.n326 vss.n325 9.3005
R221 vss.n291 vss.n290 9.3005
R222 vss.n58 vss.n57 9.3005
R223 vss.n57 vss.n56 9.3005
R224 vss.n56 vss.n55 9.3005
R225 vss.n278 vss.n277 9.0005
R226 vss.n272 vss.n271 9.0005
R227 vss.n19 vss.n18 9.0005
R228 vss.n214 vss.n213 9.0005
R229 vss.n61 vss.n60 9.0005
R230 vss.n57 vss.n47 5.64756
R231 vss.n12 vss.n2 5.64756
R232 vss.n130 vss.n118 5.64756
R233 vss.n173 vss.n162 5.64756
R234 vss.n39 vss.n29 4.89462
R235 vss.n155 vss.n143 4.89462
R236 vss.n210 vss.n200 4.89462
R237 vss.n27 vss.n26 4.6505
R238 vss.n141 vss.n140 4.6505
R239 vss.n266 vss.n265 4.57427
R240 vss.n192 vss.n182 4.14168
R241 vss.n246 vss.n236 4.14168
R242 vss.n257 vss.n256 3.76521
R243 vss.n229 vss.n221 3.38874
R244 vss.n221 vss.n220 3.01226
R245 vss.n276 vss.n275 3.01226
R246 vss.n327 vss.n326 2.69871
R247 vss.n265 vss.n257 2.63579
R248 vss.n277 vss.n276 2.63579
R249 vss.n182 vss.n181 2.25932
R250 vss.n236 vss.n235 2.25932
R251 vss.n29 vss.n28 1.50638
R252 vss.n143 vss.n142 1.50638
R253 vss.n200 vss.n199 1.50638
R254 vss.n100 vss.n99 1.45154
R255 vss.n106 vss.n105 0.827063
R256 vss.n47 vss.n46 0.753441
R257 vss.n2 vss.n1 0.753441
R258 vss.n118 vss.n117 0.753441
R259 vss.n162 vss.n161 0.753441
R260 vss.n327 vss.n116 0.409111
R261 vss.n110 vss.n109 0.3755
R262 vss.n102 vss.n101 0.341125
R263 vss.n40 vss.n27 0.240083
R264 vss.n156 vss.n141 0.240083
R265 vss.n193 vss.n180 0.240083
R266 vss.n254 vss.n253 0.185917
R267 vss.n141 vss.n135 0.146333
R268 vss.n230 vss.n219 0.133833
R269 vss.n174 vss.n160 0.110917
R270 vss.n247 vss.n234 0.110917
R271 vss.n219 vss.n218 0.10675
R272 vss vss.n327 0.0949305
R273 vss.n45 vss.n44 0.09425
R274 vss.n109 vss.n108 0.0864375
R275 vss.n27 vss.n21 0.0859167
R276 vss.n198 vss.n197 0.0838333
R277 vss.n105 vss.n104 0.078625
R278 vss.n13 vss.n0 0.063
R279 vss.n273 vss.n272 0.0421667
R280 vss.n278 vss.n274 0.0421667
R281 vss.n113 vss.n112 0.0364375
R282 vss.n266 vss.n255 0.0338333
R283 vss.n268 vss.n266 0.0338333
R284 vss.n133 vss.n131 0.03175
R285 vss.n176 vss.n174 0.03175
R286 vss.n291 vss.n289 0.03175
R287 vss.n101 vss.n100 0.03175
R288 vss.n114 vss.n113 0.03175
R289 vss.n116 vss.n115 0.03175
R290 vss.n20 vss.n19 0.0296667
R291 vss.n17 vss.n15 0.0296667
R292 vss.n42 vss.n40 0.0275833
R293 vss.n158 vss.n156 0.0275833
R294 vss.n211 vss.n198 0.0275833
R295 vss.n107 vss.n106 0.0270625
R296 vss.n59 vss.n58 0.0255
R297 vss.n21 vss.n20 0.0255
R298 vss.n112 vss.n111 0.0255
R299 vss.n195 vss.n193 0.0234167
R300 vss.n249 vss.n247 0.0234167
R301 vss.n104 vss.n103 0.022375
R302 vss.n255 vss.n254 0.0213333
R303 vss.n214 vss.n212 0.01925
R304 vss.n232 vss.n230 0.01925
R305 vss.n103 vss.n102 0.01925
R306 vss.n58 vss.n45 0.0171667
R307 vss.n234 vss.n232 0.0171667
R308 vss.n111 vss.n110 0.016125
R309 vss.n108 vss.n107 0.0145625
R310 vss.n197 vss.n195 0.013
R311 vss.n253 vss.n249 0.013
R312 vss.n272 vss.n270 0.013
R313 vss.n274 vss.n273 0.0109167
R314 vss.n44 vss.n42 0.00883333
R315 vss.n160 vss.n158 0.00883333
R316 vss.n212 vss.n211 0.00883333
R317 vss.n218 vss.n214 0.00883333
R318 vss.n115 vss.n114 0.0083125
R319 vss.n61 vss.n59 0.00675
R320 vss.n19 vss.n17 0.00675
R321 vss.n15 vss.n13 0.00675
R322 vss.n135 vss.n133 0.00466667
R323 vss.n180 vss.n176 0.00466667
R324 vss.n289 vss.n278 0.00466667
R325 vss.n326 vss.n291 0.00466667
R326 vss.n99 vss.n61 0.00449567
R327 vss.n270 vss.n268 0.00258333
R328 Q.n16 Q.n15 185.683
R329 Q.n49 Q.t0 112.225
R330 Q.n49 Q.t1 107.438
R331 Q.n35 Q.n34 92.5005
R332 Q.n11 Q.n10 13.177
R333 Q.n36 Q.n35 13.177
R334 Q.n17 Q.n16 9.32733
R335 Q.n41 Q.n40 9.32596
R336 Q.n12 Q.n11 9.3005
R337 Q.n5 Q.n4 9.3005
R338 Q.n2 Q.n1 9.3005
R339 Q.n25 Q.n24 9.3005
R340 Q.n37 Q.n36 9.3005
R341 Q.n29 Q.n28 9.3005
R342 Q.n3 Q.n0 9.0005
R343 Q.n14 Q.n13 9.0005
R344 Q.n39 Q.n38 9.0005
R345 Q.n27 Q.n26 9.0005
R346 Q.n50 Q.n48 2.77388
R347 Q.n42 Q.n41 2.2535
R348 Q.n18 Q.n17 2.25346
R349 Q Q.n50 1.00467
R350 Q.n48 Q.n23 0.682942
R351 Q.n48 Q.n47 0.660969
R352 Q.n50 Q.n49 0.462457
R353 Q.n8 Q.n7 0.0525833
R354 Q.n32 Q.n31 0.0525833
R355 Q.n9 Q.n8 0.0421667
R356 Q.n31 Q.n30 0.0421667
R357 Q.n7 Q.n6 0.0400833
R358 Q.n33 Q.n32 0.0400833
R359 Q.n20 Q.n19 0.0395625
R360 Q.n44 Q.n43 0.0395625
R361 Q.n3 Q.n2 0.0338333
R362 Q.n27 Q.n25 0.0338333
R363 Q.n19 Q.n18 0.03175
R364 Q.n23 Q.n22 0.03175
R365 Q.n45 Q.n44 0.03175
R366 Q.n21 Q.n20 0.0301875
R367 Q.n47 Q.n46 0.0301875
R368 Q.n43 Q.n42 0.0301875
R369 Q.n17 Q.n14 0.00990809
R370 Q.n41 Q.n39 0.009283
R371 Q.n12 Q.n9 0.00675
R372 Q.n6 Q.n5 0.00675
R373 Q.n22 Q.n21 0.00675
R374 Q.n30 Q.n29 0.00675
R375 Q.n37 Q.n33 0.00675
R376 Q.n46 Q.n45 0.00675
R377 Q.n14 Q.n12 0.00258333
R378 Q.n5 Q.n3 0.00258333
R379 Q.n29 Q.n27 0.00258333
R380 Q.n39 Q.n37 0.00258333
R381 R.n0 R.t0 112.543
R382 R.n0 R.t1 107.12
R383 R R.n0 0.354667
R384 vdd.n18 vdd.n14 99.0123
R385 vdd.n38 vdd.n36 95.8462
R386 vdd.n127 vdd.n125 95.8462
R387 vdd.n163 vdd.n161 95.8462
R388 vdd.n230 vdd.n228 95.8462
R389 vdd.n164 vdd.n163 93.0272
R390 vdd.n249 vdd.n239 92.5005
R391 vdd.n239 vdd.n238 92.5005
R392 vdd.n248 vdd.n247 92.5005
R393 vdd.n245 vdd.n244 92.5005
R394 vdd.n243 vdd.n242 92.5005
R395 vdd.n241 vdd.n240 92.5005
R396 vdd.n254 vdd.n253 92.5005
R397 vdd.n228 vdd.n227 92.5005
R398 vdd.n230 vdd.n229 92.5005
R399 vdd.n225 vdd.n224 92.5005
R400 vdd.n226 vdd.n225 92.5005
R401 vdd.n206 vdd.n205 92.5005
R402 vdd.n207 vdd.n206 92.5005
R403 vdd.n188 vdd.n187 92.5005
R404 vdd.n185 vdd.n184 92.5005
R405 vdd.n186 vdd.n185 92.5005
R406 vdd.n172 vdd.n171 92.5005
R407 vdd.n173 vdd.n172 92.5005
R408 vdd.n163 vdd.n162 92.5005
R409 vdd.n161 vdd.n160 92.5005
R410 vdd.n149 vdd.n148 92.5005
R411 vdd.n145 vdd.n144 92.5005
R412 vdd.n141 vdd.n140 92.5005
R413 vdd.n137 vdd.n136 92.5005
R414 vdd.n93 vdd.n92 92.5005
R415 vdd.n97 vdd.n96 92.5005
R416 vdd.n101 vdd.n100 92.5005
R417 vdd.n105 vdd.n104 92.5005
R418 vdd.n125 vdd.n124 92.5005
R419 vdd.n127 vdd.n126 92.5005
R420 vdd.n123 vdd.n122 92.5005
R421 vdd.n129 vdd.n123 92.5005
R422 vdd.n81 vdd.n80 92.5005
R423 vdd.n83 vdd.n81 92.5005
R424 vdd.n79 vdd.n78 92.5005
R425 vdd.n61 vdd.n60 92.5005
R426 vdd.n63 vdd.n61 92.5005
R427 vdd.n44 vdd.n43 92.5005
R428 vdd.n46 vdd.n44 92.5005
R429 vdd.n38 vdd.n37 92.5005
R430 vdd.n36 vdd.n35 92.5005
R431 vdd.n20 vdd.n19 92.5005
R432 vdd.n16 vdd.n15 92.5005
R433 vdd.n1 vdd.n0 92.5005
R434 vdd.n3 vdd.n2 92.5005
R435 vdd.n6 vdd.n5 92.5005
R436 vdd.n9 vdd.n8 92.5005
R437 vdd.n14 vdd.n13 92.5005
R438 vdd.n18 vdd.n17 92.5005
R439 vdd.n17 vdd.n16 92.5005
R440 vdd.n22 vdd.n21 92.5005
R441 vdd.n21 vdd.n20 92.5005
R442 vdd.n24 vdd.n23 92.5005
R443 vdd.n26 vdd.n25 92.5005
R444 vdd.n69 vdd.n68 92.5005
R445 vdd.n111 vdd.n110 92.5005
R446 vdd.n109 vdd.n108 92.5005
R447 vdd.n107 vdd.n106 92.5005
R448 vdd.n106 vdd.n105 92.5005
R449 vdd.n103 vdd.n102 92.5005
R450 vdd.n102 vdd.n101 92.5005
R451 vdd.n99 vdd.n98 92.5005
R452 vdd.n98 vdd.n97 92.5005
R453 vdd.n95 vdd.n94 92.5005
R454 vdd.n94 vdd.n93 92.5005
R455 vdd.n139 vdd.n138 92.5005
R456 vdd.n138 vdd.n137 92.5005
R457 vdd.n143 vdd.n142 92.5005
R458 vdd.n142 vdd.n141 92.5005
R459 vdd.n147 vdd.n146 92.5005
R460 vdd.n146 vdd.n145 92.5005
R461 vdd.n151 vdd.n150 92.5005
R462 vdd.n150 vdd.n149 92.5005
R463 vdd.n153 vdd.n152 92.5005
R464 vdd.n155 vdd.n154 92.5005
R465 vdd.n196 vdd.n195 92.5005
R466 vdd.n260 vdd.n259 92.5005
R467 vdd.n258 vdd.n257 92.5005
R468 vdd.n256 vdd.n255 92.5005
R469 vdd.n255 vdd.n254 92.5005
R470 vdd.n252 vdd.n251 92.5005
R471 vdd.n251 vdd.n250 92.5005
R472 vdd.n47 vdd.n38 85.9797
R473 vdd.n84 vdd.n79 83.1607
R474 vdd.n128 vdd.n127 81.7512
R475 vdd.n252 vdd.n249 79.4358
R476 vdd.n231 vdd.n230 74.7038
R477 vdd.n5 vdd.n4 72.7879
R478 vdd.n8 vdd.n7 72.7879
R479 vdd.n189 vdd.n188 71.8848
R480 vdd.n190 vdd.n183 60.0005
R481 vdd.n175 vdd.n159 52.9417
R482 vdd.n232 vdd.n219 52.9417
R483 vdd.n247 vdd.n246 52.2363
R484 vdd.n209 vdd.n202 45.8829
R485 vdd.n13 vdd.n12 42.8997
R486 vdd.n58 vdd.n57 42.3534
R487 vdd.n34 vdd.n33 35.2946
R488 vdd.n115 vdd.n114 35.2946
R489 vdd.n12 vdd.n11 33.0688
R490 vdd.n11 vdd.n10 33.0686
R491 vdd.n85 vdd.n77 31.7652
R492 vdd.n77 vdd.n76 28.2358
R493 vdd.n249 vdd.n248 25.6005
R494 vdd.n248 vdd.n245 25.6005
R495 vdd.n245 vdd.n243 25.6005
R496 vdd.n243 vdd.n241 25.6005
R497 vdd.n40 vdd.n39 25.6005
R498 vdd.n41 vdd.n40 25.6005
R499 vdd.n42 vdd.n41 25.6005
R500 vdd.n43 vdd.n42 25.6005
R501 vdd.n60 vdd.n59 25.6005
R502 vdd.n122 vdd.n121 25.6005
R503 vdd.n121 vdd.n120 25.6005
R504 vdd.n120 vdd.n119 25.6005
R505 vdd.n119 vdd.n118 25.6005
R506 vdd.n118 vdd.n117 25.6005
R507 vdd.n117 vdd.n116 25.6005
R508 vdd.n166 vdd.n165 25.6005
R509 vdd.n167 vdd.n166 25.6005
R510 vdd.n168 vdd.n167 25.6005
R511 vdd.n169 vdd.n168 25.6005
R512 vdd.n170 vdd.n169 25.6005
R513 vdd.n171 vdd.n170 25.6005
R514 vdd.n205 vdd.n204 25.6005
R515 vdd.n224 vdd.n223 25.6005
R516 vdd.n223 vdd.n222 25.6005
R517 vdd.n222 vdd.n221 25.6005
R518 vdd.n14 vdd.n9 25.6005
R519 vdd.n9 vdd.n6 25.6005
R520 vdd.n6 vdd.n3 25.6005
R521 vdd.n3 vdd.n1 25.6005
R522 vdd.n22 vdd.n18 25.6005
R523 vdd.n24 vdd.n22 25.6005
R524 vdd.n26 vdd.n24 25.6005
R525 vdd.n111 vdd.n109 25.6005
R526 vdd.n109 vdd.n107 25.6005
R527 vdd.n107 vdd.n103 25.6005
R528 vdd.n103 vdd.n99 25.6005
R529 vdd.n99 vdd.n95 25.6005
R530 vdd.n143 vdd.n139 25.6005
R531 vdd.n147 vdd.n143 25.6005
R532 vdd.n151 vdd.n147 25.6005
R533 vdd.n153 vdd.n151 25.6005
R534 vdd.n155 vdd.n153 25.6005
R535 vdd.n260 vdd.n258 25.6005
R536 vdd.n258 vdd.n256 25.6005
R537 vdd.n256 vdd.n252 25.6005
R538 vdd.n156 vdd.n155 24.8476
R539 vdd.n48 vdd.n34 24.7064
R540 vdd.n131 vdd.n115 24.7064
R541 vdd.n189 vdd.n186 23.9619
R542 vdd.n112 vdd.n111 21.8358
R543 vdd.n174 vdd.n173 21.1429
R544 vdd.n231 vdd.n226 21.1429
R545 vdd.n238 vdd.n237 20.1334
R546 vdd.n208 vdd.n207 18.3239
R547 vdd.n65 vdd.n58 17.6476
R548 vdd.n63 vdd.n62 16.9144
R549 vdd.n27 vdd.n26 16.5652
R550 vdd.n70 vdd.n69 15.8123
R551 vdd.n202 vdd.n201 14.1181
R552 vdd.n46 vdd.n45 14.0955
R553 vdd.n129 vdd.n128 14.0955
R554 vdd.n261 vdd.n260 13.5534
R555 vdd.n197 vdd.n196 12.8005
R556 vdd.n84 vdd.n83 12.686
R557 vdd.n83 vdd.n82 11.2765
R558 vdd.n47 vdd.n46 9.86697
R559 vdd.n130 vdd.n129 9.86697
R560 vdd.n262 vdd.n261 9.3005
R561 vdd.n192 vdd.n191 9.3005
R562 vdd.n191 vdd.n190 9.3005
R563 vdd.n190 vdd.n189 9.3005
R564 vdd.n177 vdd.n176 9.3005
R565 vdd.n176 vdd.n175 9.3005
R566 vdd.n175 vdd.n174 9.3005
R567 vdd.n181 vdd.n180 9.3005
R568 vdd.n179 vdd.n178 9.3005
R569 vdd.n194 vdd.n193 9.3005
R570 vdd.n198 vdd.n197 9.3005
R571 vdd.n211 vdd.n210 9.3005
R572 vdd.n210 vdd.n209 9.3005
R573 vdd.n209 vdd.n208 9.3005
R574 vdd.n215 vdd.n214 9.3005
R575 vdd.n213 vdd.n212 9.3005
R576 vdd.n236 vdd.n235 9.3005
R577 vdd.n234 vdd.n233 9.3005
R578 vdd.n233 vdd.n232 9.3005
R579 vdd.n232 vdd.n231 9.3005
R580 vdd.n89 vdd.n88 9.3005
R581 vdd.n71 vdd.n70 9.3005
R582 vdd.n67 vdd.n66 9.3005
R583 vdd.n66 vdd.n65 9.3005
R584 vdd.n65 vdd.n64 9.3005
R585 vdd.n52 vdd.n51 9.3005
R586 vdd.n28 vdd.n27 9.3005
R587 vdd.n54 vdd.n53 9.3005
R588 vdd.n30 vdd.n29 9.3005
R589 vdd.n50 vdd.n49 9.3005
R590 vdd.n49 vdd.n48 9.3005
R591 vdd.n48 vdd.n47 9.3005
R592 vdd.n87 vdd.n86 9.3005
R593 vdd.n86 vdd.n85 9.3005
R594 vdd.n85 vdd.n84 9.3005
R595 vdd.n73 vdd.n72 9.3005
R596 vdd.n91 vdd.n90 9.3005
R597 vdd.n133 vdd.n132 9.3005
R598 vdd.n132 vdd.n131 9.3005
R599 vdd.n131 vdd.n130 9.3005
R600 vdd.n159 vdd.n158 7.05932
R601 vdd.n219 vdd.n218 7.05932
R602 vdd.n64 vdd.n63 7.04798
R603 vdd.n191 vdd.n182 6.4005
R604 vdd.n176 vdd.n157 5.64756
R605 vdd.n233 vdd.n217 5.64756
R606 vdd.n207 vdd.n203 5.63848
R607 vdd.n210 vdd.n200 4.89462
R608 vdd.n56 vdd.n55 4.51815
R609 vdd.n32 vdd.n31 3.76521
R610 vdd.n113 vdd.n112 3.76521
R611 vdd.n86 vdd.n75 3.38874
R612 vdd.n75 vdd.n74 3.01226
R613 vdd.n173 vdd.n164 2.81949
R614 vdd.n226 vdd.n220 2.81949
R615 vdd.n49 vdd.n32 2.63579
R616 vdd.n132 vdd.n113 2.63579
R617 vdd.n263 vdd.n262 2.52787
R618 vdd.n134 vdd.n133 2.43829
R619 vdd.n66 vdd.n56 1.88285
R620 vdd.n200 vdd.n199 1.50638
R621 vdd.n263 vdd.n135 0.980223
R622 vdd.n135 vdd.n134 0.954986
R623 vdd.n157 vdd.n156 0.753441
R624 vdd.n217 vdd.n216 0.753441
R625 vdd.n211 vdd.n198 0.240083
R626 vdd.n71 vdd.n67 0.240083
R627 vdd.n192 vdd.n181 0.110917
R628 vdd.n234 vdd.n215 0.110917
R629 vdd.n52 vdd.n50 0.110917
R630 vdd.n89 vdd.n87 0.110917
R631 vdd vdd.n263 0.0949305
R632 vdd.n194 vdd.n192 0.0338333
R633 vdd.n179 vdd.n177 0.0296667
R634 vdd.n236 vdd.n234 0.0296667
R635 vdd.n213 vdd.n211 0.0255
R636 vdd.n54 vdd.n52 0.0234167
R637 vdd.n87 vdd.n73 0.0213333
R638 vdd.n30 vdd.n28 0.01925
R639 vdd.n91 vdd.n89 0.01925
R640 vdd.n50 vdd.n30 0.0171667
R641 vdd.n133 vdd.n91 0.0171667
R642 vdd.n73 vdd.n71 0.0150833
R643 vdd.n67 vdd.n54 0.013
R644 vdd.n215 vdd.n213 0.0109167
R645 vdd.n181 vdd.n179 0.00675
R646 vdd.n262 vdd.n236 0.00675
R647 vdd.n198 vdd.n194 0.00258333
R648 S.n0 S.t0 112.543
R649 S.n0 S.t1 107.12
R650 S S.n0 0.417167
R651 Qn.n16 Qn.n15 185.683
R652 Qn.n49 Qn.t0 112.859
R653 Qn.n49 Qn.t1 106.802
R654 Qn.n35 Qn.n34 92.5005
R655 Qn.n11 Qn.n10 13.177
R656 Qn.n36 Qn.n35 13.177
R657 Qn.n17 Qn.n16 9.32733
R658 Qn.n41 Qn.n40 9.32596
R659 Qn.n12 Qn.n11 9.3005
R660 Qn.n5 Qn.n4 9.3005
R661 Qn.n2 Qn.n1 9.3005
R662 Qn.n25 Qn.n24 9.3005
R663 Qn.n37 Qn.n36 9.3005
R664 Qn.n29 Qn.n28 9.3005
R665 Qn.n3 Qn.n0 9.0005
R666 Qn.n14 Qn.n13 9.0005
R667 Qn.n39 Qn.n38 9.0005
R668 Qn.n27 Qn.n26 9.0005
R669 Qn Qn.n48 2.98602
R670 Qn.n42 Qn.n41 2.2535
R671 Qn.n18 Qn.n17 2.25346
R672 Qn.n48 Qn.n23 0.68449
R673 Qn.n48 Qn.n47 0.660418
R674 Qn Qn.n49 0.410826
R675 Qn.n8 Qn.n7 0.0525833
R676 Qn.n32 Qn.n31 0.0525833
R677 Qn.n9 Qn.n8 0.0421667
R678 Qn.n31 Qn.n30 0.0421667
R679 Qn.n7 Qn.n6 0.0400833
R680 Qn.n33 Qn.n32 0.0400833
R681 Qn.n20 Qn.n19 0.0395625
R682 Qn.n44 Qn.n43 0.0395625
R683 Qn.n3 Qn.n2 0.0338333
R684 Qn.n27 Qn.n25 0.0338333
R685 Qn.n19 Qn.n18 0.03175
R686 Qn.n23 Qn.n22 0.03175
R687 Qn.n45 Qn.n44 0.03175
R688 Qn.n21 Qn.n20 0.0301875
R689 Qn.n47 Qn.n46 0.0301875
R690 Qn.n43 Qn.n42 0.0301875
R691 Qn.n17 Qn.n14 0.00990809
R692 Qn.n41 Qn.n39 0.009283
R693 Qn.n12 Qn.n9 0.00675
R694 Qn.n6 Qn.n5 0.00675
R695 Qn.n22 Qn.n21 0.00675
R696 Qn.n30 Qn.n29 0.00675
R697 Qn.n37 Qn.n33 0.00675
R698 Qn.n46 Qn.n45 0.00675
R699 Qn.n14 Qn.n12 0.00258333
R700 Qn.n5 Qn.n3 0.00258333
R701 Qn.n29 Qn.n27 0.00258333
R702 Qn.n39 Qn.n37 0.00258333
C0 Qn S 0.0154f
C1 vdd m1_458_623# 0.205f
C2 Qn Q 0.597f
C3 Q R 0.0155f
C4 vdd S 0.16f
C5 Q vdd 0.478f
C6 Qn vdd 0.213f
C7 Q m1_1673_493# 0.102f
C8 vdd R 0.157f
C9 Qn m1_1673_493# 0.0695f
C10 m1_1673_493# R 0.0341f
C11 S m1_458_623# 0.0341f
C12 m1_1673_493# vdd 0.206f
C13 Q m1_458_623# 0.0695f
C14 Qn m1_458_623# 0.102f
C15 Q S 1.46e-19
C16 Q vss 0.819f
C17 Qn vss 0.884f
C18 m1_458_623# vss 0.663f
C19 S vss 0.479f
C20 m1_1673_493# vss 0.66f
C21 R vss 0.478f
C22 vdd vss 6.99f
.ends

