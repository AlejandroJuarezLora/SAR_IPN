magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_p >>
rect -743 1183 1687 1245
rect -743 1077 -681 1183
rect -575 677 -513 1077
rect -575 615 1519 677
rect 1625 615 1687 1183
<< nwell >>
rect -681 1077 1625 1183
rect -681 615 -575 1077
rect 1519 615 1625 1077
rect -681 509 1625 615
<< nsubdiff >>
rect -645 1113 -557 1147
rect -523 1113 -489 1147
rect -455 1113 -421 1147
rect -387 1113 -353 1147
rect -319 1113 -285 1147
rect -251 1113 -217 1147
rect -183 1113 -149 1147
rect -115 1113 -81 1147
rect -47 1113 -13 1147
rect 21 1113 55 1147
rect 89 1113 123 1147
rect 157 1113 191 1147
rect 225 1113 259 1147
rect 293 1113 327 1147
rect 361 1113 395 1147
rect 429 1113 463 1147
rect 497 1113 531 1147
rect 565 1113 599 1147
rect 633 1113 667 1147
rect 701 1113 735 1147
rect 769 1113 803 1147
rect 837 1113 871 1147
rect 905 1113 939 1147
rect 973 1113 1007 1147
rect 1041 1113 1075 1147
rect 1109 1113 1143 1147
rect 1177 1113 1211 1147
rect 1245 1113 1279 1147
rect 1313 1113 1347 1147
rect 1381 1113 1415 1147
rect 1449 1113 1589 1147
rect -645 1007 -611 1113
rect -645 939 -611 973
rect -645 871 -611 905
rect -645 803 -611 837
rect -645 735 -611 769
rect -645 579 -611 701
rect 1555 1007 1589 1113
rect 1555 939 1589 973
rect 1555 871 1589 905
rect 1555 803 1589 837
rect 1555 735 1589 769
rect 1555 579 1589 701
rect -645 545 -489 579
rect -455 545 -421 579
rect -387 545 -353 579
rect -319 545 -285 579
rect -251 545 -217 579
rect -183 545 -149 579
rect -115 545 -81 579
rect -47 545 -13 579
rect 21 545 55 579
rect 89 545 123 579
rect 157 545 191 579
rect 225 545 259 579
rect 293 545 327 579
rect 361 545 395 579
rect 429 545 463 579
rect 497 545 531 579
rect 565 545 599 579
rect 633 545 667 579
rect 701 545 735 579
rect 769 545 803 579
rect 837 545 871 579
rect 905 545 939 579
rect 973 545 1007 579
rect 1041 545 1075 579
rect 1109 545 1143 579
rect 1177 545 1211 579
rect 1245 545 1279 579
rect 1313 545 1347 579
rect 1381 545 1415 579
rect 1449 545 1589 579
<< nsubdiffcont >>
rect -557 1113 -523 1147
rect -489 1113 -455 1147
rect -421 1113 -387 1147
rect -353 1113 -319 1147
rect -285 1113 -251 1147
rect -217 1113 -183 1147
rect -149 1113 -115 1147
rect -81 1113 -47 1147
rect -13 1113 21 1147
rect 55 1113 89 1147
rect 123 1113 157 1147
rect 191 1113 225 1147
rect 259 1113 293 1147
rect 327 1113 361 1147
rect 395 1113 429 1147
rect 463 1113 497 1147
rect 531 1113 565 1147
rect 599 1113 633 1147
rect 667 1113 701 1147
rect 735 1113 769 1147
rect 803 1113 837 1147
rect 871 1113 905 1147
rect 939 1113 973 1147
rect 1007 1113 1041 1147
rect 1075 1113 1109 1147
rect 1143 1113 1177 1147
rect 1211 1113 1245 1147
rect 1279 1113 1313 1147
rect 1347 1113 1381 1147
rect 1415 1113 1449 1147
rect -645 973 -611 1007
rect -645 905 -611 939
rect -645 837 -611 871
rect -645 769 -611 803
rect -645 701 -611 735
rect 1555 973 1589 1007
rect 1555 905 1589 939
rect 1555 837 1589 871
rect 1555 769 1589 803
rect 1555 701 1589 735
rect -489 545 -455 579
rect -421 545 -387 579
rect -353 545 -319 579
rect -285 545 -251 579
rect -217 545 -183 579
rect -149 545 -115 579
rect -81 545 -47 579
rect -13 545 21 579
rect 55 545 89 579
rect 123 545 157 579
rect 191 545 225 579
rect 259 545 293 579
rect 327 545 361 579
rect 395 545 429 579
rect 463 545 497 579
rect 531 545 565 579
rect 599 545 633 579
rect 667 545 701 579
rect 735 545 769 579
rect 803 545 837 579
rect 871 545 905 579
rect 939 545 973 579
rect 1007 545 1041 579
rect 1075 545 1109 579
rect 1143 545 1177 579
rect 1211 545 1245 579
rect 1279 545 1313 579
rect 1347 545 1381 579
rect 1415 545 1449 579
<< locali >>
rect -645 1113 -557 1147
rect -523 1113 -489 1147
rect -455 1113 -421 1147
rect -387 1113 -353 1147
rect -319 1113 -285 1147
rect -251 1113 -217 1147
rect -183 1113 -149 1147
rect -115 1113 -81 1147
rect -47 1113 -13 1147
rect 21 1113 55 1147
rect 89 1113 123 1147
rect 157 1113 191 1147
rect 225 1113 259 1147
rect 293 1113 327 1147
rect 361 1113 395 1147
rect 429 1113 463 1147
rect 497 1113 531 1147
rect 565 1113 599 1147
rect 633 1113 667 1147
rect 701 1113 735 1147
rect 769 1113 803 1147
rect 837 1113 871 1147
rect 905 1113 939 1147
rect 973 1113 1007 1147
rect 1041 1113 1075 1147
rect 1109 1113 1143 1147
rect 1177 1113 1211 1147
rect 1245 1113 1279 1147
rect 1313 1113 1347 1147
rect 1381 1113 1415 1147
rect 1449 1113 1589 1147
rect -645 1007 -611 1113
rect -645 939 -611 973
rect -645 871 -611 905
rect -645 803 -611 837
rect -645 735 -611 769
rect -645 579 -611 701
rect 1555 1007 1589 1113
rect 1555 939 1589 973
rect 1555 871 1589 905
rect 1555 803 1589 837
rect 1555 735 1589 769
rect 1555 579 1589 701
rect -645 545 -489 579
rect -455 545 -421 579
rect -387 545 -353 579
rect -319 545 -285 579
rect -251 545 -217 579
rect -183 545 -149 579
rect -115 545 -81 579
rect -47 545 -13 579
rect 21 545 55 579
rect 89 545 123 579
rect 157 545 191 579
rect 225 545 259 579
rect 293 545 327 579
rect 361 545 395 579
rect 429 545 463 579
rect 497 545 531 579
rect 565 545 599 579
rect 633 545 667 579
rect 701 545 735 579
rect 769 545 803 579
rect 837 545 871 579
rect 905 545 939 579
rect 973 545 1007 579
rect 1041 545 1075 579
rect 1109 545 1143 579
rect 1177 545 1211 579
rect 1245 545 1279 579
rect 1313 545 1347 579
rect 1381 545 1415 579
rect 1449 545 1589 579
<< properties >>
string path -17.025 28.250 39.300 28.250 39.300 14.050 -15.700 14.050 -15.700 28.250 
<< end >>
