magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< nwell >>
rect -38 221 774 542
<< pwell >>
rect 35 -19 735 163
rect 35 -23 62 -19
rect 28 -57 62 -23
<< scnmos >>
rect 113 7 143 137
rect 197 7 227 137
rect 293 7 323 137
rect 401 7 431 137
rect 509 7 539 137
rect 621 7 651 137
<< scpmoshvt >>
rect 113 257 143 457
rect 197 257 227 457
rect 293 257 323 457
rect 401 257 431 457
rect 509 257 539 457
rect 621 257 651 457
<< ndiff >>
rect 61 121 113 137
rect 61 87 69 121
rect 103 87 113 121
rect 61 53 113 87
rect 61 19 69 53
rect 103 19 113 53
rect 61 7 113 19
rect 143 53 197 137
rect 143 19 153 53
rect 187 19 197 53
rect 143 7 197 19
rect 227 121 293 137
rect 227 87 244 121
rect 278 87 293 121
rect 227 53 293 87
rect 227 19 244 53
rect 278 19 293 53
rect 227 7 293 19
rect 323 53 401 137
rect 323 19 345 53
rect 379 19 401 53
rect 323 7 401 19
rect 431 121 509 137
rect 431 87 458 121
rect 492 87 509 121
rect 431 53 509 87
rect 431 19 458 53
rect 492 19 509 53
rect 431 7 509 19
rect 539 121 621 137
rect 539 87 558 121
rect 592 87 621 121
rect 539 7 621 87
rect 651 53 709 137
rect 651 19 661 53
rect 695 19 709 53
rect 651 7 709 19
<< pdiff >>
rect 46 435 113 457
rect 46 401 60 435
rect 94 401 113 435
rect 46 329 113 401
rect 46 295 60 329
rect 94 295 113 329
rect 46 257 113 295
rect 143 445 197 457
rect 143 411 153 445
rect 187 411 197 445
rect 143 377 197 411
rect 143 343 153 377
rect 187 343 197 377
rect 143 257 197 343
rect 227 257 293 457
rect 323 257 401 457
rect 431 445 509 457
rect 431 411 452 445
rect 486 411 509 445
rect 431 377 509 411
rect 431 343 452 377
rect 486 343 509 377
rect 431 257 509 343
rect 539 257 621 457
rect 651 445 709 457
rect 651 411 661 445
rect 695 411 709 445
rect 651 377 709 411
rect 651 343 661 377
rect 695 343 709 377
rect 651 309 709 343
rect 651 275 661 309
rect 695 275 709 309
rect 651 257 709 275
<< ndiffc >>
rect 69 87 103 121
rect 69 19 103 53
rect 153 19 187 53
rect 244 87 278 121
rect 244 19 278 53
rect 345 19 379 53
rect 458 87 492 121
rect 458 19 492 53
rect 558 87 592 121
rect 661 19 695 53
<< pdiffc >>
rect 60 401 94 435
rect 60 295 94 329
rect 153 411 187 445
rect 153 343 187 377
rect 452 411 486 445
rect 452 343 486 377
rect 661 411 695 445
rect 661 343 695 377
rect 661 275 695 309
<< poly >>
rect 113 457 143 483
rect 197 457 227 483
rect 293 457 323 483
rect 401 457 431 483
rect 509 457 539 483
rect 621 457 651 483
rect 113 225 143 257
rect 197 225 227 257
rect 293 225 323 257
rect 401 225 431 257
rect 509 225 539 257
rect 621 225 651 257
rect 77 209 143 225
rect 77 175 93 209
rect 127 175 143 209
rect 77 159 143 175
rect 185 209 251 225
rect 185 175 201 209
rect 235 175 251 209
rect 185 159 251 175
rect 293 209 359 225
rect 293 175 309 209
rect 343 175 359 209
rect 293 159 359 175
rect 401 209 467 225
rect 401 175 417 209
rect 451 175 467 209
rect 401 159 467 175
rect 509 209 575 225
rect 509 175 525 209
rect 559 175 575 209
rect 509 159 575 175
rect 621 209 714 225
rect 621 175 664 209
rect 698 175 714 209
rect 621 159 714 175
rect 113 137 143 159
rect 197 137 227 159
rect 293 137 323 159
rect 401 137 431 159
rect 509 137 539 159
rect 621 137 651 159
rect 113 -19 143 7
rect 197 -19 227 7
rect 293 -19 323 7
rect 401 -19 431 7
rect 509 -19 539 7
rect 621 -19 651 7
<< polycont >>
rect 93 175 127 209
rect 201 175 235 209
rect 309 175 343 209
rect 417 175 451 209
rect 525 175 559 209
rect 664 175 698 209
<< locali >>
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 17 435 94 451
rect 17 401 60 435
rect 17 329 94 401
rect 17 295 60 329
rect 137 445 195 487
rect 137 411 153 445
rect 187 411 195 445
rect 137 377 195 411
rect 137 343 153 377
rect 187 343 195 377
rect 137 327 195 343
rect 229 445 502 453
rect 229 419 452 445
rect 17 259 94 295
rect 229 293 263 419
rect 436 411 452 419
rect 486 411 502 445
rect 128 259 263 293
rect 17 125 52 259
rect 128 225 162 259
rect 297 225 362 385
rect 436 377 502 411
rect 661 445 719 487
rect 695 411 719 445
rect 661 377 719 411
rect 436 343 452 377
rect 486 343 627 377
rect 436 327 627 343
rect 89 209 162 225
rect 89 175 93 209
rect 127 175 162 209
rect 201 209 251 225
rect 235 175 251 209
rect 293 209 362 225
rect 293 175 309 209
rect 343 175 362 209
rect 89 159 127 175
rect 201 159 235 175
rect 293 159 362 175
rect 396 209 451 292
rect 396 175 417 209
rect 396 159 451 175
rect 488 209 559 292
rect 488 175 525 209
rect 488 159 559 175
rect 593 125 627 327
rect 695 343 719 377
rect 661 309 719 343
rect 695 275 719 309
rect 661 259 719 275
rect 664 209 719 225
rect 698 175 719 209
rect 664 159 719 175
rect 17 121 119 125
rect 17 87 69 121
rect 103 87 119 121
rect 228 121 508 125
rect 17 53 119 87
rect 17 19 69 53
rect 103 19 119 53
rect 17 11 119 19
rect 153 53 187 89
rect 153 -23 187 19
rect 228 87 244 121
rect 278 91 458 121
rect 278 87 294 91
rect 228 53 294 87
rect 442 87 458 91
rect 492 87 508 121
rect 542 121 627 125
rect 542 87 558 121
rect 592 87 627 121
rect 228 19 244 53
rect 278 19 294 53
rect 228 11 294 19
rect 329 53 395 57
rect 329 19 345 53
rect 379 19 395 53
rect 329 -23 395 19
rect 442 53 508 87
rect 661 53 719 107
rect 442 19 458 53
rect 492 19 661 53
rect 695 19 719 53
rect 442 11 719 19
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
<< viali >>
rect 29 487 63 521
rect 121 487 155 521
rect 213 487 247 521
rect 305 487 339 521
rect 397 487 431 521
rect 489 487 523 521
rect 581 487 615 521
rect 673 487 707 521
rect 29 -57 63 -23
rect 121 -57 155 -23
rect 213 -57 247 -23
rect 305 -57 339 -23
rect 397 -57 431 -23
rect 489 -57 523 -23
rect 581 -57 615 -23
rect 673 -57 707 -23
<< metal1 >>
rect 0 521 736 552
rect 0 487 29 521
rect 63 487 121 521
rect 155 487 213 521
rect 247 487 305 521
rect 339 487 397 521
rect 431 487 489 521
rect 523 487 581 521
rect 615 487 673 521
rect 707 487 736 521
rect 0 456 736 487
rect 0 -23 736 8
rect 0 -57 29 -23
rect 63 -57 121 -23
rect 155 -57 213 -23
rect 247 -57 305 -23
rect 339 -57 397 -23
rect 431 -57 489 -23
rect 523 -57 581 -23
rect 615 -57 673 -23
rect 707 -57 736 -23
rect 0 -88 736 -57
<< labels >>
rlabel comment s 0 -40 0 -40 4 o32a_1
flabel metal1 s 28 487 62 521 0 FreeSans 200 0 0 0 VPWR
port 2 nsew
flabel metal1 s 28 -57 62 -23 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel nwell s 28 487 62 521 0 FreeSans 200 0 0 0 VPB
port 5 nsew
flabel pwell s 28 -57 62 -23 0 FreeSans 200 0 0 0 VNB
port 6 nsew
flabel locali s 28 45 62 79 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 28 385 62 419 0 FreeSans 250 0 0 0 X
port 7 nsew
flabel locali s 396 249 430 283 0 FreeSans 250 0 0 0 A3
port 10 nsew
flabel locali s 212 181 246 215 0 FreeSans 250 0 0 0 A1
port 8 nsew
flabel locali s 304 181 338 215 0 FreeSans 250 0 0 0 A2
port 9 nsew
flabel locali s 396 181 430 215 0 FreeSans 250 0 0 0 A3
port 10 nsew
flabel locali s 672 181 706 215 0 FreeSans 250 0 0 0 B1
port 12 nsew
flabel locali s 488 181 522 215 0 FreeSans 250 0 0 0 B2
port 11 nsew
flabel locali s 304 249 338 283 0 FreeSans 250 0 0 0 A2
port 9 nsew
flabel locali s 304 317 338 351 0 FreeSans 250 0 0 0 A2
port 9 nsew
flabel locali s 488 249 522 283 0 FreeSans 250 0 0 0 B2
port 11 nsew
flabel locali s 28 317 62 351 0 FreeSans 250 0 0 0 X
port 7 nsew
<< properties >>
string FIXED_BBOX 0 -40 736 504
string path 0.000 -1.000 18.400 -1.000 
<< end >>
