magic
tech sky130B
magscale 1 2
timestamp 1696364841
<< error_p >>
rect -36 -151 36 -145
rect -36 -185 -17 -151
rect -36 -191 36 -185
<< nwell >>
rect -236 -324 236 244
<< pmoslvt >>
rect -40 -104 40 96
<< pdiff >>
rect -98 81 -40 96
rect -98 47 -86 81
rect -52 47 -40 81
rect -98 13 -40 47
rect -98 -21 -86 13
rect -52 -21 -40 13
rect -98 -55 -40 -21
rect -98 -89 -86 -55
rect -52 -89 -40 -55
rect -98 -104 -40 -89
rect 40 81 98 96
rect 40 47 52 81
rect 86 47 98 81
rect 40 13 98 47
rect 40 -21 52 13
rect 86 -21 98 13
rect 40 -55 98 -21
rect 40 -89 52 -55
rect 86 -89 98 -55
rect 40 -104 98 -89
<< pdiffc >>
rect -86 47 -52 81
rect -86 -21 -52 13
rect -86 -89 -52 -55
rect 52 47 86 81
rect 52 -21 86 13
rect 52 -89 86 -55
<< poly >>
rect -40 96 40 122
rect -40 -151 40 -104
rect -40 -185 -17 -151
rect 17 -185 40 -151
rect -40 -201 40 -185
<< polycont >>
rect -17 -185 17 -151
<< locali >>
rect -86 81 -52 100
rect -86 13 -52 15
rect -86 -23 -52 -21
rect -86 -108 -52 -89
rect 52 81 86 100
rect 52 13 86 15
rect 52 -23 86 -21
rect 52 -108 86 -89
rect -40 -185 -17 -151
rect 17 -185 40 -151
<< viali >>
rect -86 47 -52 49
rect -86 15 -52 47
rect -86 -55 -52 -23
rect -86 -57 -52 -55
rect 52 47 86 49
rect 52 15 86 47
rect 52 -55 86 -23
rect 52 -57 86 -55
rect -17 -185 17 -151
<< metal1 >>
rect -92 49 -46 96
rect -92 15 -86 49
rect -52 15 -46 49
rect -92 -23 -46 15
rect -92 -57 -86 -23
rect -52 -57 -46 -23
rect -92 -104 -46 -57
rect 46 49 92 96
rect 46 15 52 49
rect 86 15 92 49
rect 46 -23 92 15
rect 46 -57 52 -23
rect 86 -57 92 -23
rect 46 -104 92 -57
rect -36 -151 36 -145
rect -36 -185 -17 -151
rect 17 -185 36 -151
rect -36 -191 36 -185
<< end >>
