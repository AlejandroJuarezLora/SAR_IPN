magic
tech sky130B
magscale 1 2
timestamp 1697748102
<< metal1 >>
rect 4 2335 2286 2342
rect 4 2283 72 2335
rect 124 2283 136 2335
rect 188 2283 296 2335
rect 348 2283 360 2335
rect 412 2283 520 2335
rect 572 2283 584 2335
rect 636 2283 744 2335
rect 796 2283 808 2335
rect 860 2283 968 2335
rect 1020 2283 1032 2335
rect 1084 2283 1192 2335
rect 1244 2283 1256 2335
rect 1308 2283 1416 2335
rect 1468 2283 1480 2335
rect 1532 2283 1640 2335
rect 1692 2283 1704 2335
rect 1756 2283 1864 2335
rect 1916 2283 1928 2335
rect 1980 2283 2088 2335
rect 2140 2283 2152 2335
rect 2204 2283 2286 2335
rect 4 2276 2286 2283
rect 4 98 32 2276
rect 60 70 88 2248
rect 116 98 144 2276
rect 172 70 200 2248
rect 228 98 256 2276
rect 284 70 312 2248
rect 340 98 368 2276
rect 396 70 424 2248
rect 452 98 480 2276
rect 508 70 536 2248
rect 564 98 592 2276
rect 620 70 648 2248
rect 676 98 704 2276
rect 732 70 760 2248
rect 788 98 816 2276
rect 844 70 872 2248
rect 900 98 928 2276
rect 956 70 984 2248
rect 1012 98 1040 2276
rect 1068 70 1096 2248
rect 1124 98 1152 2276
rect 1180 70 1208 2248
rect 1236 98 1264 2276
rect 1292 70 1320 2248
rect 1348 98 1376 2276
rect 1404 70 1432 2248
rect 1460 98 1488 2276
rect 1516 70 1544 2248
rect 1572 98 1600 2276
rect 1628 70 1656 2248
rect 1684 98 1712 2276
rect 1740 70 1768 2248
rect 1796 98 1824 2276
rect 1852 70 1880 2248
rect 1908 98 1936 2276
rect 1964 70 1992 2248
rect 2020 98 2048 2276
rect 2076 70 2104 2248
rect 2132 98 2160 2276
rect 2188 70 2216 2248
rect 2244 98 2286 2276
rect 4 63 2286 70
rect 4 11 28 63
rect 80 11 92 63
rect 144 11 240 63
rect 292 11 304 63
rect 356 11 464 63
rect 516 11 528 63
rect 580 11 688 63
rect 740 11 752 63
rect 804 11 912 63
rect 964 11 976 63
rect 1028 11 1136 63
rect 1188 11 1200 63
rect 1252 11 1360 63
rect 1412 11 1424 63
rect 1476 11 1584 63
rect 1636 11 1648 63
rect 1700 11 1808 63
rect 1860 11 1872 63
rect 1924 11 2032 63
rect 2084 11 2096 63
rect 2148 11 2286 63
rect 4 4 2286 11
<< via1 >>
rect 72 2283 124 2335
rect 136 2283 188 2335
rect 296 2283 348 2335
rect 360 2283 412 2335
rect 520 2283 572 2335
rect 584 2283 636 2335
rect 744 2283 796 2335
rect 808 2283 860 2335
rect 968 2283 1020 2335
rect 1032 2283 1084 2335
rect 1192 2283 1244 2335
rect 1256 2283 1308 2335
rect 1416 2283 1468 2335
rect 1480 2283 1532 2335
rect 1640 2283 1692 2335
rect 1704 2283 1756 2335
rect 1864 2283 1916 2335
rect 1928 2283 1980 2335
rect 2088 2283 2140 2335
rect 2152 2283 2204 2335
rect 28 11 80 63
rect 92 11 144 63
rect 240 11 292 63
rect 304 11 356 63
rect 464 11 516 63
rect 528 11 580 63
rect 688 11 740 63
rect 752 11 804 63
rect 912 11 964 63
rect 976 11 1028 63
rect 1136 11 1188 63
rect 1200 11 1252 63
rect 1360 11 1412 63
rect 1424 11 1476 63
rect 1584 11 1636 63
rect 1648 11 1700 63
rect 1808 11 1860 63
rect 1872 11 1924 63
rect 2032 11 2084 63
rect 2096 11 2148 63
<< metal2 >>
rect 4 70 32 2342
rect 60 2337 200 2342
rect 60 2335 102 2337
rect 158 2335 200 2337
rect 60 2283 72 2335
rect 188 2283 200 2335
rect 60 2281 102 2283
rect 158 2281 200 2283
rect 60 2276 200 2281
rect 60 98 88 2276
rect 116 70 144 2248
rect 4 65 144 70
rect 4 63 46 65
rect 102 63 144 65
rect 4 11 28 63
rect 4 9 46 11
rect 102 9 144 11
rect 4 4 144 9
rect 172 4 200 2276
rect 228 70 256 2342
rect 284 2337 424 2342
rect 284 2335 326 2337
rect 382 2335 424 2337
rect 284 2283 296 2335
rect 412 2283 424 2335
rect 284 2281 326 2283
rect 382 2281 424 2283
rect 284 2276 424 2281
rect 284 98 312 2276
rect 340 70 368 2248
rect 228 65 368 70
rect 228 63 270 65
rect 326 63 368 65
rect 228 11 240 63
rect 356 11 368 63
rect 228 9 270 11
rect 326 9 368 11
rect 228 4 368 9
rect 396 4 424 2276
rect 452 70 480 2342
rect 508 2337 648 2342
rect 508 2335 550 2337
rect 606 2335 648 2337
rect 508 2283 520 2335
rect 636 2283 648 2335
rect 508 2281 550 2283
rect 606 2281 648 2283
rect 508 2276 648 2281
rect 508 98 536 2276
rect 564 70 592 2248
rect 452 65 592 70
rect 452 63 494 65
rect 550 63 592 65
rect 452 11 464 63
rect 580 11 592 63
rect 452 9 494 11
rect 550 9 592 11
rect 452 4 592 9
rect 620 4 648 2276
rect 676 70 704 2342
rect 732 2337 872 2342
rect 732 2335 774 2337
rect 830 2335 872 2337
rect 732 2283 744 2335
rect 860 2283 872 2335
rect 732 2281 774 2283
rect 830 2281 872 2283
rect 732 2276 872 2281
rect 732 98 760 2276
rect 788 70 816 2248
rect 676 65 816 70
rect 676 63 718 65
rect 774 63 816 65
rect 676 11 688 63
rect 804 11 816 63
rect 676 9 718 11
rect 774 9 816 11
rect 676 4 816 9
rect 844 4 872 2276
rect 900 70 928 2342
rect 956 2337 1096 2342
rect 956 2335 998 2337
rect 1054 2335 1096 2337
rect 956 2283 968 2335
rect 1084 2283 1096 2335
rect 956 2281 998 2283
rect 1054 2281 1096 2283
rect 956 2276 1096 2281
rect 956 98 984 2276
rect 1012 70 1040 2248
rect 900 65 1040 70
rect 900 63 942 65
rect 998 63 1040 65
rect 900 11 912 63
rect 1028 11 1040 63
rect 900 9 942 11
rect 998 9 1040 11
rect 900 4 1040 9
rect 1068 4 1096 2276
rect 1124 70 1152 2342
rect 1180 2337 1320 2342
rect 1180 2335 1222 2337
rect 1278 2335 1320 2337
rect 1180 2283 1192 2335
rect 1308 2283 1320 2335
rect 1180 2281 1222 2283
rect 1278 2281 1320 2283
rect 1180 2276 1320 2281
rect 1180 98 1208 2276
rect 1236 70 1264 2248
rect 1124 65 1264 70
rect 1124 63 1166 65
rect 1222 63 1264 65
rect 1124 11 1136 63
rect 1252 11 1264 63
rect 1124 9 1166 11
rect 1222 9 1264 11
rect 1124 4 1264 9
rect 1292 4 1320 2276
rect 1348 70 1376 2342
rect 1404 2337 1544 2342
rect 1404 2335 1446 2337
rect 1502 2335 1544 2337
rect 1404 2283 1416 2335
rect 1532 2283 1544 2335
rect 1404 2281 1446 2283
rect 1502 2281 1544 2283
rect 1404 2276 1544 2281
rect 1404 98 1432 2276
rect 1460 70 1488 2248
rect 1348 65 1488 70
rect 1348 63 1390 65
rect 1446 63 1488 65
rect 1348 11 1360 63
rect 1476 11 1488 63
rect 1348 9 1390 11
rect 1446 9 1488 11
rect 1348 4 1488 9
rect 1516 4 1544 2276
rect 1572 70 1600 2342
rect 1628 2337 1768 2342
rect 1628 2335 1670 2337
rect 1726 2335 1768 2337
rect 1628 2283 1640 2335
rect 1756 2283 1768 2335
rect 1628 2281 1670 2283
rect 1726 2281 1768 2283
rect 1628 2276 1768 2281
rect 1628 98 1656 2276
rect 1684 70 1712 2248
rect 1572 65 1712 70
rect 1572 63 1614 65
rect 1670 63 1712 65
rect 1572 11 1584 63
rect 1700 11 1712 63
rect 1572 9 1614 11
rect 1670 9 1712 11
rect 1572 4 1712 9
rect 1740 4 1768 2276
rect 1796 70 1824 2342
rect 1852 2337 2286 2342
rect 1852 2335 1894 2337
rect 1950 2335 2118 2337
rect 2174 2335 2286 2337
rect 1852 2283 1864 2335
rect 1980 2283 2088 2335
rect 2204 2283 2286 2335
rect 1852 2281 1894 2283
rect 1950 2281 2118 2283
rect 2174 2281 2286 2283
rect 1852 2276 2286 2281
rect 1852 98 1880 2276
rect 1908 70 1936 2248
rect 1796 65 1936 70
rect 1796 63 1838 65
rect 1894 63 1936 65
rect 1796 11 1808 63
rect 1924 11 1936 63
rect 1796 9 1838 11
rect 1894 9 1936 11
rect 1796 4 1936 9
rect 1964 4 1992 2276
rect 2020 70 2048 2248
rect 2076 98 2104 2276
rect 2132 70 2160 2248
rect 2188 98 2216 2276
rect 2244 70 2286 2248
rect 2020 65 2286 70
rect 2020 63 2062 65
rect 2118 63 2286 65
rect 2020 11 2032 63
rect 2148 11 2286 63
rect 2020 9 2062 11
rect 2118 9 2286 11
rect 2020 4 2286 9
<< via2 >>
rect 102 2335 158 2337
rect 102 2283 124 2335
rect 124 2283 136 2335
rect 136 2283 158 2335
rect 102 2281 158 2283
rect 46 63 102 65
rect 46 11 80 63
rect 80 11 92 63
rect 92 11 102 63
rect 46 9 102 11
rect 326 2335 382 2337
rect 326 2283 348 2335
rect 348 2283 360 2335
rect 360 2283 382 2335
rect 326 2281 382 2283
rect 270 63 326 65
rect 270 11 292 63
rect 292 11 304 63
rect 304 11 326 63
rect 270 9 326 11
rect 550 2335 606 2337
rect 550 2283 572 2335
rect 572 2283 584 2335
rect 584 2283 606 2335
rect 550 2281 606 2283
rect 494 63 550 65
rect 494 11 516 63
rect 516 11 528 63
rect 528 11 550 63
rect 494 9 550 11
rect 774 2335 830 2337
rect 774 2283 796 2335
rect 796 2283 808 2335
rect 808 2283 830 2335
rect 774 2281 830 2283
rect 718 63 774 65
rect 718 11 740 63
rect 740 11 752 63
rect 752 11 774 63
rect 718 9 774 11
rect 998 2335 1054 2337
rect 998 2283 1020 2335
rect 1020 2283 1032 2335
rect 1032 2283 1054 2335
rect 998 2281 1054 2283
rect 942 63 998 65
rect 942 11 964 63
rect 964 11 976 63
rect 976 11 998 63
rect 942 9 998 11
rect 1222 2335 1278 2337
rect 1222 2283 1244 2335
rect 1244 2283 1256 2335
rect 1256 2283 1278 2335
rect 1222 2281 1278 2283
rect 1166 63 1222 65
rect 1166 11 1188 63
rect 1188 11 1200 63
rect 1200 11 1222 63
rect 1166 9 1222 11
rect 1446 2335 1502 2337
rect 1446 2283 1468 2335
rect 1468 2283 1480 2335
rect 1480 2283 1502 2335
rect 1446 2281 1502 2283
rect 1390 63 1446 65
rect 1390 11 1412 63
rect 1412 11 1424 63
rect 1424 11 1446 63
rect 1390 9 1446 11
rect 1670 2335 1726 2337
rect 1670 2283 1692 2335
rect 1692 2283 1704 2335
rect 1704 2283 1726 2335
rect 1670 2281 1726 2283
rect 1614 63 1670 65
rect 1614 11 1636 63
rect 1636 11 1648 63
rect 1648 11 1670 63
rect 1614 9 1670 11
rect 1894 2335 1950 2337
rect 2118 2335 2174 2337
rect 1894 2283 1916 2335
rect 1916 2283 1928 2335
rect 1928 2283 1950 2335
rect 2118 2283 2140 2335
rect 2140 2283 2152 2335
rect 2152 2283 2174 2335
rect 1894 2281 1950 2283
rect 2118 2281 2174 2283
rect 1838 63 1894 65
rect 1838 11 1860 63
rect 1860 11 1872 63
rect 1872 11 1894 63
rect 1838 9 1894 11
rect 2062 63 2118 65
rect 2062 11 2084 63
rect 2084 11 2096 63
rect 2096 11 2118 63
rect 2062 9 2118 11
<< metal3 >>
rect 4 2341 2286 2342
rect 4 2277 32 2341
rect 96 2337 112 2341
rect 96 2281 102 2337
rect 96 2277 112 2281
rect 176 2277 192 2341
rect 256 2277 272 2341
rect 336 2337 352 2341
rect 336 2277 352 2281
rect 416 2277 432 2341
rect 496 2277 512 2341
rect 576 2337 592 2341
rect 576 2277 592 2281
rect 656 2277 672 2341
rect 736 2277 752 2341
rect 816 2337 832 2341
rect 830 2281 832 2337
rect 816 2277 832 2281
rect 896 2277 912 2341
rect 976 2277 992 2341
rect 1056 2277 1072 2341
rect 1136 2277 1152 2341
rect 1216 2337 1232 2341
rect 1216 2281 1222 2337
rect 1216 2277 1232 2281
rect 1296 2277 1312 2341
rect 1376 2277 1392 2341
rect 1456 2337 1472 2341
rect 1456 2277 1472 2281
rect 1536 2277 1552 2341
rect 1616 2277 1632 2341
rect 1696 2337 1712 2341
rect 1696 2277 1712 2281
rect 1776 2277 1792 2341
rect 1856 2277 1872 2341
rect 1936 2337 1952 2341
rect 1950 2281 1952 2337
rect 1936 2277 1952 2281
rect 2016 2277 2032 2341
rect 2096 2277 2112 2341
rect 2176 2277 2192 2341
rect 2256 2277 2286 2341
rect 4 2276 2286 2277
rect 4 130 64 2276
rect 124 70 184 2216
rect 244 130 304 2276
rect 364 70 424 2216
rect 484 130 544 2276
rect 604 70 664 2216
rect 724 130 784 2276
rect 844 70 904 2216
rect 964 130 1024 2276
rect 1084 70 1144 2216
rect 1204 130 1264 2276
rect 1324 70 1384 2216
rect 1444 130 1504 2276
rect 1564 70 1624 2216
rect 1684 130 1744 2276
rect 1804 70 1864 2216
rect 1924 130 1984 2276
rect 2044 70 2104 2216
rect 2164 130 2286 2276
rect 4 69 2286 70
rect 4 5 32 69
rect 96 65 112 69
rect 102 9 112 65
rect 96 5 112 9
rect 176 5 192 69
rect 256 65 272 69
rect 256 9 270 65
rect 256 5 272 9
rect 336 5 352 69
rect 416 5 432 69
rect 496 65 512 69
rect 496 5 512 9
rect 576 5 592 69
rect 656 5 672 69
rect 736 65 752 69
rect 736 5 752 9
rect 816 5 832 69
rect 896 5 912 69
rect 976 65 992 69
rect 976 5 992 9
rect 1056 5 1072 69
rect 1136 5 1152 69
rect 1216 65 1232 69
rect 1222 9 1232 65
rect 1216 5 1232 9
rect 1296 5 1312 69
rect 1376 65 1392 69
rect 1376 9 1390 65
rect 1376 5 1392 9
rect 1456 5 1472 69
rect 1536 5 1552 69
rect 1616 65 1632 69
rect 1616 5 1632 9
rect 1696 5 1712 69
rect 1776 5 1792 69
rect 1856 65 1872 69
rect 1856 5 1872 9
rect 1936 5 1952 69
rect 2016 5 2032 69
rect 2096 65 2112 69
rect 2096 5 2112 9
rect 2176 5 2192 69
rect 2256 5 2286 69
rect 4 4 2286 5
<< via3 >>
rect 32 2277 96 2341
rect 112 2337 176 2341
rect 112 2281 158 2337
rect 158 2281 176 2337
rect 112 2277 176 2281
rect 192 2277 256 2341
rect 272 2337 336 2341
rect 352 2337 416 2341
rect 272 2281 326 2337
rect 326 2281 336 2337
rect 352 2281 382 2337
rect 382 2281 416 2337
rect 272 2277 336 2281
rect 352 2277 416 2281
rect 432 2277 496 2341
rect 512 2337 576 2341
rect 592 2337 656 2341
rect 512 2281 550 2337
rect 550 2281 576 2337
rect 592 2281 606 2337
rect 606 2281 656 2337
rect 512 2277 576 2281
rect 592 2277 656 2281
rect 672 2277 736 2341
rect 752 2337 816 2341
rect 752 2281 774 2337
rect 774 2281 816 2337
rect 752 2277 816 2281
rect 832 2277 896 2341
rect 912 2277 976 2341
rect 992 2337 1056 2341
rect 992 2281 998 2337
rect 998 2281 1054 2337
rect 1054 2281 1056 2337
rect 992 2277 1056 2281
rect 1072 2277 1136 2341
rect 1152 2277 1216 2341
rect 1232 2337 1296 2341
rect 1232 2281 1278 2337
rect 1278 2281 1296 2337
rect 1232 2277 1296 2281
rect 1312 2277 1376 2341
rect 1392 2337 1456 2341
rect 1472 2337 1536 2341
rect 1392 2281 1446 2337
rect 1446 2281 1456 2337
rect 1472 2281 1502 2337
rect 1502 2281 1536 2337
rect 1392 2277 1456 2281
rect 1472 2277 1536 2281
rect 1552 2277 1616 2341
rect 1632 2337 1696 2341
rect 1712 2337 1776 2341
rect 1632 2281 1670 2337
rect 1670 2281 1696 2337
rect 1712 2281 1726 2337
rect 1726 2281 1776 2337
rect 1632 2277 1696 2281
rect 1712 2277 1776 2281
rect 1792 2277 1856 2341
rect 1872 2337 1936 2341
rect 1872 2281 1894 2337
rect 1894 2281 1936 2337
rect 1872 2277 1936 2281
rect 1952 2277 2016 2341
rect 2032 2277 2096 2341
rect 2112 2337 2176 2341
rect 2112 2281 2118 2337
rect 2118 2281 2174 2337
rect 2174 2281 2176 2337
rect 2112 2277 2176 2281
rect 2192 2277 2256 2341
rect 32 65 96 69
rect 32 9 46 65
rect 46 9 96 65
rect 32 5 96 9
rect 112 5 176 69
rect 192 5 256 69
rect 272 65 336 69
rect 272 9 326 65
rect 326 9 336 65
rect 272 5 336 9
rect 352 5 416 69
rect 432 65 496 69
rect 512 65 576 69
rect 432 9 494 65
rect 494 9 496 65
rect 512 9 550 65
rect 550 9 576 65
rect 432 5 496 9
rect 512 5 576 9
rect 592 5 656 69
rect 672 65 736 69
rect 752 65 816 69
rect 672 9 718 65
rect 718 9 736 65
rect 752 9 774 65
rect 774 9 816 65
rect 672 5 736 9
rect 752 5 816 9
rect 832 5 896 69
rect 912 65 976 69
rect 992 65 1056 69
rect 912 9 942 65
rect 942 9 976 65
rect 992 9 998 65
rect 998 9 1056 65
rect 912 5 976 9
rect 992 5 1056 9
rect 1072 5 1136 69
rect 1152 65 1216 69
rect 1152 9 1166 65
rect 1166 9 1216 65
rect 1152 5 1216 9
rect 1232 5 1296 69
rect 1312 5 1376 69
rect 1392 65 1456 69
rect 1392 9 1446 65
rect 1446 9 1456 65
rect 1392 5 1456 9
rect 1472 5 1536 69
rect 1552 65 1616 69
rect 1632 65 1696 69
rect 1552 9 1614 65
rect 1614 9 1616 65
rect 1632 9 1670 65
rect 1670 9 1696 65
rect 1552 5 1616 9
rect 1632 5 1696 9
rect 1712 5 1776 69
rect 1792 65 1856 69
rect 1872 65 1936 69
rect 1792 9 1838 65
rect 1838 9 1856 65
rect 1872 9 1894 65
rect 1894 9 1936 65
rect 1792 5 1856 9
rect 1872 5 1936 9
rect 1952 5 2016 69
rect 2032 65 2096 69
rect 2112 65 2176 69
rect 2032 9 2062 65
rect 2062 9 2096 65
rect 2112 9 2118 65
rect 2118 9 2176 65
rect 2032 5 2096 9
rect 2112 5 2176 9
rect 2192 5 2256 69
<< metal4 >>
rect 4 2341 2286 2342
rect 4 2277 32 2341
rect 96 2277 112 2341
rect 176 2277 192 2341
rect 256 2277 272 2341
rect 336 2277 352 2341
rect 416 2277 432 2341
rect 496 2277 512 2341
rect 576 2277 592 2341
rect 656 2277 672 2341
rect 736 2277 752 2341
rect 816 2277 832 2341
rect 896 2277 912 2341
rect 976 2277 992 2341
rect 1056 2277 1072 2341
rect 1136 2277 1152 2341
rect 1216 2277 1232 2341
rect 1296 2277 1312 2341
rect 1376 2277 1392 2341
rect 1456 2277 1472 2341
rect 1536 2277 1552 2341
rect 1616 2277 1632 2341
rect 1696 2277 1712 2341
rect 1776 2277 1792 2341
rect 1856 2277 1872 2341
rect 1936 2277 1952 2341
rect 2016 2277 2032 2341
rect 2096 2277 2112 2341
rect 2176 2277 2192 2341
rect 2256 2277 2286 2341
rect 4 2276 2286 2277
rect 124 2267 424 2276
rect 4 70 64 2216
rect 124 2031 156 2267
rect 392 2031 424 2267
rect 124 130 184 2031
rect 244 315 304 1971
rect 364 375 424 2031
rect 484 315 544 2216
rect 244 79 276 315
rect 512 79 544 315
rect 604 130 664 2276
rect 244 70 544 79
rect 724 70 784 2216
rect 844 130 904 2276
rect 964 70 1024 2216
rect 1084 130 1144 2276
rect 1204 70 1264 2216
rect 1324 130 1384 2276
rect 1564 2267 1864 2276
rect 1444 70 1504 2216
rect 1564 2031 1596 2267
rect 1832 2031 1864 2267
rect 1564 130 1624 2031
rect 1684 315 1744 1971
rect 1804 375 1864 2031
rect 1924 315 1984 2216
rect 1684 79 1716 315
rect 1952 79 1984 315
rect 2044 130 2104 2276
rect 1684 70 1984 79
rect 2164 70 2286 2216
rect 4 69 2286 70
rect 4 5 32 69
rect 96 5 112 69
rect 176 5 192 69
rect 256 5 272 69
rect 336 5 352 69
rect 416 5 432 69
rect 496 5 512 69
rect 576 5 592 69
rect 656 5 672 69
rect 736 5 752 69
rect 816 5 832 69
rect 896 5 912 69
rect 976 5 992 69
rect 1056 5 1072 69
rect 1136 5 1152 69
rect 1216 5 1232 69
rect 1296 5 1312 69
rect 1376 5 1392 69
rect 1456 5 1472 69
rect 1536 5 1552 69
rect 1616 5 1632 69
rect 1696 5 1712 69
rect 1776 5 1792 69
rect 1856 5 1872 69
rect 1936 5 1952 69
rect 2016 5 2032 69
rect 2096 5 2112 69
rect 2176 5 2192 69
rect 2256 5 2286 69
rect 4 4 2286 5
<< via4 >>
rect 156 2031 392 2267
rect 276 79 512 315
rect 1596 2031 1832 2267
rect 1716 79 1952 315
<< metal5 >>
rect 4 2267 2286 2342
rect 4 2031 156 2267
rect 392 2031 1596 2267
rect 1832 2031 2286 2267
rect 4 2007 2286 2031
rect 4 659 324 2007
rect 644 339 964 1687
rect 1284 659 1604 2007
rect 1924 339 2286 1687
rect 4 315 2286 339
rect 4 79 276 315
rect 512 79 1716 315
rect 1952 79 2286 315
rect 4 4 2286 79
<< end >>
