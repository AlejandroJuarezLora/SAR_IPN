** sch_path: /home/alex/Desktop/SAR_IPN/xschem/user_analog_project_wrapper.sch
.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i_3_,wbs_sel_i_2_,wbs_sel_i_1_,wbs_sel_i_0_
+ wbs_dat_i_31_,wbs_dat_i_30_,wbs_dat_i_29_,wbs_dat_i_28_,wbs_dat_i_27_,wbs_dat_i_26_,wbs_dat_i_25_,wbs_dat_i_24_,wbs_dat_i_23_,wbs_dat_i_22_,wbs_dat_i_21_,wbs_dat_i_20_,wbs_dat_i_19_,wbs_dat_i_18_,wbs_dat_i_17_,wbs_dat_i_16_,wbs_dat_i_15_,wbs_dat_i_14_,wbs_dat_i_13_,wbs_dat_i_12_,wbs_dat_i_11_,wbs_dat_i_10_,wbs_dat_i_9_,wbs_dat_i_8_,wbs_dat_i_7_,wbs_dat_i_6_,wbs_dat_i_5_,wbs_dat_i_4_,wbs_dat_i_3_,wbs_dat_i_2_,wbs_dat_i_1_,wbs_dat_i_0_
+ wbs_adr_i_31_,wbs_adr_i_30_,wbs_adr_i_29_,wbs_adr_i_28_,wbs_adr_i_27_,wbs_adr_i_26_,wbs_adr_i_25_,wbs_adr_i_24_,wbs_adr_i_23_,wbs_adr_i_22_,wbs_adr_i_21_,wbs_adr_i_20_,wbs_adr_i_19_,wbs_adr_i_18_,wbs_adr_i_17_,wbs_adr_i_16_,wbs_adr_i_15_,wbs_adr_i_14_,wbs_adr_i_13_,wbs_adr_i_12_,wbs_adr_i_11_,wbs_adr_i_10_,wbs_adr_i_9_,wbs_adr_i_8_,wbs_adr_i_7_,wbs_adr_i_6_,wbs_adr_i_5_,wbs_adr_i_4_,wbs_adr_i_3_,wbs_adr_i_2_,wbs_adr_i_1_,wbs_adr_i_0_ wbs_ack_o
+ wbs_dat_o_31_,wbs_dat_o_30_,wbs_dat_o_29_,wbs_dat_o_28_,wbs_dat_o_27_,wbs_dat_o_26_,wbs_dat_o_25_,wbs_dat_o_24_,wbs_dat_o_23_,wbs_dat_o_22_,wbs_dat_o_21_,wbs_dat_o_20_,wbs_dat_o_19_,wbs_dat_o_18_,wbs_dat_o_17_,wbs_dat_o_16_,wbs_dat_o_15_,wbs_dat_o_14_,wbs_dat_o_13_,wbs_dat_o_12_,wbs_dat_o_11_,wbs_dat_o_10_,wbs_dat_o_9_,wbs_dat_o_8_,wbs_dat_o_7_,wbs_dat_o_6_,wbs_dat_o_5_,wbs_dat_o_4_,wbs_dat_o_3_,wbs_dat_o_2_,wbs_dat_o_1_,wbs_dat_o_0_
+ la_data_in_127_,la_data_in_126_,la_data_in_125_,la_data_in_124_,la_data_in_123_,la_data_in_122_,la_data_in_121_,la_data_in_120_,la_data_in_119_,la_data_in_118_,la_data_in_117_,la_data_in_116_,la_data_in_115_,la_data_in_114_,la_data_in_113_,la_data_in_112_,la_data_in_111_,la_data_in_110_,la_data_in_109_,la_data_in_108_,la_data_in_107_,la_data_in_106_,la_data_in_105_,la_data_in_104_,la_data_in_103_,la_data_in_102_,la_data_in_101_,la_data_in_100_,la_data_in_99_,la_data_in_98_,la_data_in_97_,la_data_in_96_,la_data_in_95_,la_data_in_94_,la_data_in_93_,la_data_in_92_,la_data_in_91_,la_data_in_90_,la_data_in_89_,la_data_in_88_,la_data_in_87_,la_data_in_86_,la_data_in_85_,la_data_in_84_,la_data_in_83_,la_data_in_82_,la_data_in_81_,la_data_in_80_,la_data_in_79_,la_data_in_78_,la_data_in_77_,la_data_in_76_,la_data_in_75_,la_data_in_74_,la_data_in_73_,la_data_in_72_,la_data_in_71_,la_data_in_70_,la_data_in_69_,la_data_in_68_,la_data_in_67_,la_data_in_66_,la_data_in_65_,la_data_in_64_,la_data_in_63_,la_data_in_62_,la_data_in_61_,la_data_in_60_,la_data_in_59_,la_data_in_58_,la_data_in_57_,la_data_in_56_,la_data_in_55_,la_data_in_54_,la_data_in_53_,la_data_in_52_,la_data_in_51_,la_data_in_50_,la_data_in_49_,la_data_in_48_,la_data_in_47_,la_data_in_46_,la_data_in_45_,la_data_in_44_,la_data_in_43_,la_data_in_42_,la_data_in_41_,la_data_in_40_,la_data_in_39_,la_data_in_38_,la_data_in_37_,la_data_in_36_,la_data_in_35_,la_data_in_34_,la_data_in_33_,la_data_in_32_,la_data_in_31_,la_data_in_30_,la_data_in_29_,la_data_in_28_,la_data_in_27_,la_data_in_26_,la_data_in_25_,la_data_in_24_,la_data_in_23_,la_data_in_22_,la_data_in_21_,la_data_in_20_,la_data_in_19_,la_data_in_18_,la_data_in_17_,la_data_in_16_,la_data_in_15_,la_data_in_14_,la_data_in_13_,la_data_in_12_,la_data_in_11_,la_data_in_10_,la_data_in_9_,la_data_in_8_,la_data_in_7_,la_data_in_6_,la_data_in_5_,la_data_in_4_,la_data_in_3_,la_data_in_2_,la_data_in_1_,la_data_in_0_
+ la_data_out_127_,la_data_out_126_,la_data_out_125_,la_data_out_124_,la_data_out_123_,la_data_out_122_,la_data_out_121_,la_data_out_120_,la_data_out_119_,la_data_out_118_,la_data_out_117_,la_data_out_116_,la_data_out_115_,la_data_out_114_,la_data_out_113_,la_data_out_112_,la_data_out_111_,la_data_out_110_,la_data_out_109_,la_data_out_108_,la_data_out_107_,la_data_out_106_,la_data_out_105_,la_data_out_104_,la_data_out_103_,la_data_out_102_,la_data_out_101_,la_data_out_100_,la_data_out_99_,la_data_out_98_,la_data_out_97_,la_data_out_96_,la_data_out_95_,la_data_out_94_,la_data_out_93_,la_data_out_92_,la_data_out_91_,la_data_out_90_,la_data_out_89_,la_data_out_88_,la_data_out_87_,la_data_out_86_,la_data_out_85_,la_data_out_84_,la_data_out_83_,la_data_out_82_,la_data_out_81_,la_data_out_80_,la_data_out_79_,la_data_out_78_,la_data_out_77_,la_data_out_76_,la_data_out_75_,la_data_out_74_,la_data_out_73_,la_data_out_72_,la_data_out_71_,la_data_out_70_,la_data_out_69_,la_data_out_68_,la_data_out_67_,la_data_out_66_,la_data_out_65_,la_data_out_64_,la_data_out_63_,la_data_out_62_,la_data_out_61_,la_data_out_60_,la_data_out_59_,la_data_out_58_,la_data_out_57_,la_data_out_56_,la_data_out_55_,la_data_out_54_,la_data_out_53_,la_data_out_52_,la_data_out_51_,la_data_out_50_,la_data_out_49_,la_data_out_48_,la_data_out_47_,la_data_out_46_,la_data_out_45_,la_data_out_44_,la_data_out_43_,la_data_out_42_,la_data_out_41_,la_data_out_40_,la_data_out_39_,la_data_out_38_,la_data_out_37_,la_data_out_36_,la_data_out_35_,la_data_out_34_,la_data_out_33_,la_data_out_32_,la_data_out_31_,la_data_out_30_,la_data_out_29_,la_data_out_28_,la_data_out_27_,la_data_out_26_,la_data_out_25_,la_data_out_24_,la_data_out_23_,la_data_out_22_,la_data_out_21_,la_data_out_20_,la_data_out_19_,la_data_out_18_,la_data_out_17_,la_data_out_16_,la_data_out_15_,la_data_out_14_,la_data_out_13_,la_data_out_12_,la_data_out_11_,la_data_out_10_,la_data_out_9_,la_data_out_8_,la_data_out_7_,la_data_out_6_,la_data_out_5_,la_data_out_4_,la_data_out_3_,la_data_out_2_,la_data_out_1_,la_data_out_0_
+ io_in_26_,io_in_25_,io_in_24_,io_in_23_,io_in_22_,io_in_21_,io_in_20_,io_in_19_,io_in_18_,io_in_17_,io_in_16_,io_in_15_,io_in_14_,io_in_13_,io_in_12_,io_in_11_,io_in_10_,io_in_9_,io_in_8_,io_in_7_,io_in_6_,io_in_5_,io_in_4_,io_in_3_,io_in_2_,io_in_1_,io_in_0_
+ io_in_3v3_26_,io_in_3v3_25_,io_in_3v3_24_,io_in_3v3_23_,io_in_3v3_22_,io_in_3v3_21_,io_in_3v3_20_,io_in_3v3_19_,io_in_3v3_18_,io_in_3v3_17_,io_in_3v3_16_,io_in_3v3_15_,io_in_3v3_14_,io_in_3v3_13_,io_in_3v3_12_,io_in_3v3_11_,io_in_3v3_10_,io_in_3v3_9_,io_in_3v3_8_,io_in_3v3_7_,io_in_3v3_6_,io_in_3v3_5_,io_in_3v3_4_,io_in_3v3_3_,io_in_3v3_2_,io_in_3v3_1_,io_in_3v3_0_ user_clock2
+ io_out_26_,io_out_25_,io_out_24_,io_out_23_,io_out_22_,io_out_21_,io_out_20_,io_out_19_,io_out_18_,io_out_17_,io_out_16_,io_out_15_,io_out_14_,io_out_13_,io_out_12_,io_out_11_,io_out_10_,io_out_9_,io_out_8_,io_out_7_,io_out_6_,io_out_5_,io_out_4_,io_out_3_,io_out_2_,io_out_1_,io_out_0_
+ io_oeb_26_,io_oeb_25_,io_oeb_24_,io_oeb_23_,io_oeb_22_,io_oeb_21_,io_oeb_20_,io_oeb_19_,io_oeb_18_,io_oeb_17_,io_oeb_16_,io_oeb_15_,io_oeb_14_,io_oeb_13_,io_oeb_12_,io_oeb_11_,io_oeb_10_,io_oeb_9_,io_oeb_8_,io_oeb_7_,io_oeb_6_,io_oeb_5_,io_oeb_4_,io_oeb_3_,io_oeb_2_,io_oeb_1_,io_oeb_0_
+ gpio_analog_17_,gpio_analog_16_,gpio_analog_15_,gpio_analog_14_,gpio_analog_13_,gpio_analog_12_,gpio_analog_11_,gpio_analog_10_,gpio_analog_9_,gpio_analog_8_,gpio_analog_7_,gpio_analog_6_,gpio_analog_5_,gpio_analog_4_,gpio_analog_3_,gpio_analog_2_,gpio_analog_1_,gpio_analog_0_
+ gpio_noesd_17_,gpio_noesd_16_,gpio_noesd_15_,gpio_noesd_14_,gpio_noesd_13_,gpio_noesd_12_,gpio_noesd_11_,gpio_noesd_10_,gpio_noesd_9_,gpio_noesd_8_,gpio_noesd_7_,gpio_noesd_6_,gpio_noesd_5_,gpio_noesd_4_,gpio_noesd_3_,gpio_noesd_2_,gpio_noesd_1_,gpio_noesd_0_
+ io_analog_10_,io_analog_9_,io_analog_8_,io_analog_7_,io_analog_6_,io_analog_5_,io_analog_4_,io_analog_3_,io_analog_2_,io_analog_1_,io_analog_0_ io_clamp_high_2_,io_clamp_high_1_,io_clamp_high_0_ io_clamp_low_2_,io_clamp_low_1_,io_clamp_low_0_
+ user_irq_2_,user_irq_1_,user_irq_0_
+ la_oenb_127_,la_oenb_126_,la_oenb_125_,la_oenb_124_,la_oenb_123_,la_oenb_122_,la_oenb_121_,la_oenb_120_,la_oenb_119_,la_oenb_118_,la_oenb_117_,la_oenb_116_,la_oenb_115_,la_oenb_114_,la_oenb_113_,la_oenb_112_,la_oenb_111_,la_oenb_110_,la_oenb_109_,la_oenb_108_,la_oenb_107_,la_oenb_106_,la_oenb_105_,la_oenb_104_,la_oenb_103_,la_oenb_102_,la_oenb_101_,la_oenb_100_,la_oenb_99_,la_oenb_98_,la_oenb_97_,la_oenb_96_,la_oenb_95_,la_oenb_94_,la_oenb_93_,la_oenb_92_,la_oenb_91_,la_oenb_90_,la_oenb_89_,la_oenb_88_,la_oenb_87_,la_oenb_86_,la_oenb_85_,la_oenb_84_,la_oenb_83_,la_oenb_82_,la_oenb_81_,la_oenb_80_,la_oenb_79_,la_oenb_78_,la_oenb_77_,la_oenb_76_,la_oenb_75_,la_oenb_74_,la_oenb_73_,la_oenb_72_,la_oenb_71_,la_oenb_70_,la_oenb_69_,la_oenb_68_,la_oenb_67_,la_oenb_66_,la_oenb_65_,la_oenb_64_,la_oenb_63_,la_oenb_62_,la_oenb_61_,la_oenb_60_,la_oenb_59_,la_oenb_58_,la_oenb_57_,la_oenb_56_,la_oenb_55_,la_oenb_54_,la_oenb_53_,la_oenb_52_,la_oenb_51_,la_oenb_50_,la_oenb_49_,la_oenb_48_,la_oenb_47_,la_oenb_46_,la_oenb_45_,la_oenb_44_,la_oenb_43_,la_oenb_42_,la_oenb_41_,la_oenb_40_,la_oenb_39_,la_oenb_38_,la_oenb_37_,la_oenb_36_,la_oenb_35_,la_oenb_34_,la_oenb_33_,la_oenb_32_,la_oenb_31_,la_oenb_30_,la_oenb_29_,la_oenb_28_,la_oenb_27_,la_oenb_26_,la_oenb_25_,la_oenb_24_,la_oenb_23_,la_oenb_22_,la_oenb_21_,la_oenb_20_,la_oenb_19_,la_oenb_18_,la_oenb_17_,la_oenb_16_,la_oenb_15_,la_oenb_14_,la_oenb_13_,la_oenb_12_,la_oenb_11_,la_oenb_10_,la_oenb_9_,la_oenb_8_,la_oenb_7_,la_oenb_6_,la_oenb_5_,la_oenb_4_,la_oenb_3_,la_oenb_2_,la_oenb_1_,la_oenb_0_
*.iopin vdda1
*.iopin vdda2
*.iopin vssa1
*.iopin vssa2
*.iopin vccd1
*.iopin vccd2
*.iopin vssd1
*.iopin vssd2
*.ipin wb_clk_i
*.ipin wb_rst_i
*.ipin wbs_stb_i
*.ipin wbs_cyc_i
*.ipin wbs_we_i
*.ipin wbs_sel_i_3_,wbs_sel_i_2_,wbs_sel_i_1_,wbs_sel_i_0_
*.ipin
*+ wbs_dat_i_31_,wbs_dat_i_30_,wbs_dat_i_29_,wbs_dat_i_28_,wbs_dat_i_27_,wbs_dat_i_26_,wbs_dat_i_25_,wbs_dat_i_24_,wbs_dat_i_23_,wbs_dat_i_22_,wbs_dat_i_21_,wbs_dat_i_20_,wbs_dat_i_19_,wbs_dat_i_18_,wbs_dat_i_17_,wbs_dat_i_16_,wbs_dat_i_15_,wbs_dat_i_14_,wbs_dat_i_13_,wbs_dat_i_12_,wbs_dat_i_11_,wbs_dat_i_10_,wbs_dat_i_9_,wbs_dat_i_8_,wbs_dat_i_7_,wbs_dat_i_6_,wbs_dat_i_5_,wbs_dat_i_4_,wbs_dat_i_3_,wbs_dat_i_2_,wbs_dat_i_1_,wbs_dat_i_0_
*.ipin
*+ wbs_adr_i_31_,wbs_adr_i_30_,wbs_adr_i_29_,wbs_adr_i_28_,wbs_adr_i_27_,wbs_adr_i_26_,wbs_adr_i_25_,wbs_adr_i_24_,wbs_adr_i_23_,wbs_adr_i_22_,wbs_adr_i_21_,wbs_adr_i_20_,wbs_adr_i_19_,wbs_adr_i_18_,wbs_adr_i_17_,wbs_adr_i_16_,wbs_adr_i_15_,wbs_adr_i_14_,wbs_adr_i_13_,wbs_adr_i_12_,wbs_adr_i_11_,wbs_adr_i_10_,wbs_adr_i_9_,wbs_adr_i_8_,wbs_adr_i_7_,wbs_adr_i_6_,wbs_adr_i_5_,wbs_adr_i_4_,wbs_adr_i_3_,wbs_adr_i_2_,wbs_adr_i_1_,wbs_adr_i_0_
*.opin wbs_ack_o
*.opin
*+ wbs_dat_o_31_,wbs_dat_o_30_,wbs_dat_o_29_,wbs_dat_o_28_,wbs_dat_o_27_,wbs_dat_o_26_,wbs_dat_o_25_,wbs_dat_o_24_,wbs_dat_o_23_,wbs_dat_o_22_,wbs_dat_o_21_,wbs_dat_o_20_,wbs_dat_o_19_,wbs_dat_o_18_,wbs_dat_o_17_,wbs_dat_o_16_,wbs_dat_o_15_,wbs_dat_o_14_,wbs_dat_o_13_,wbs_dat_o_12_,wbs_dat_o_11_,wbs_dat_o_10_,wbs_dat_o_9_,wbs_dat_o_8_,wbs_dat_o_7_,wbs_dat_o_6_,wbs_dat_o_5_,wbs_dat_o_4_,wbs_dat_o_3_,wbs_dat_o_2_,wbs_dat_o_1_,wbs_dat_o_0_
*.ipin
*+ la_data_in_127_,la_data_in_126_,la_data_in_125_,la_data_in_124_,la_data_in_123_,la_data_in_122_,la_data_in_121_,la_data_in_120_,la_data_in_119_,la_data_in_118_,la_data_in_117_,la_data_in_116_,la_data_in_115_,la_data_in_114_,la_data_in_113_,la_data_in_112_,la_data_in_111_,la_data_in_110_,la_data_in_109_,la_data_in_108_,la_data_in_107_,la_data_in_106_,la_data_in_105_,la_data_in_104_,la_data_in_103_,la_data_in_102_,la_data_in_101_,la_data_in_100_,la_data_in_99_,la_data_in_98_,la_data_in_97_,la_data_in_96_,la_data_in_95_,la_data_in_94_,la_data_in_93_,la_data_in_92_,la_data_in_91_,la_data_in_90_,la_data_in_89_,la_data_in_88_,la_data_in_87_,la_data_in_86_,la_data_in_85_,la_data_in_84_,la_data_in_83_,la_data_in_82_,la_data_in_81_,la_data_in_80_,la_data_in_79_,la_data_in_78_,la_data_in_77_,la_data_in_76_,la_data_in_75_,la_data_in_74_,la_data_in_73_,la_data_in_72_,la_data_in_71_,la_data_in_70_,la_data_in_69_,la_data_in_68_,la_data_in_67_,la_data_in_66_,la_data_in_65_,la_data_in_64_,la_data_in_63_,la_data_in_62_,la_data_in_61_,la_data_in_60_,la_data_in_59_,la_data_in_58_,la_data_in_57_,la_data_in_56_,la_data_in_55_,la_data_in_54_,la_data_in_53_,la_data_in_52_,la_data_in_51_,la_data_in_50_,la_data_in_49_,la_data_in_48_,la_data_in_47_,la_data_in_46_,la_data_in_45_,la_data_in_44_,la_data_in_43_,la_data_in_42_,la_data_in_41_,la_data_in_40_,la_data_in_39_,la_data_in_38_,la_data_in_37_,la_data_in_36_,la_data_in_35_,la_data_in_34_,la_data_in_33_,la_data_in_32_,la_data_in_31_,la_data_in_30_,la_data_in_29_,la_data_in_28_,la_data_in_27_,la_data_in_26_,la_data_in_25_,la_data_in_24_,la_data_in_23_,la_data_in_22_,la_data_in_21_,la_data_in_20_,la_data_in_19_,la_data_in_18_,la_data_in_17_,la_data_in_16_,la_data_in_15_,la_data_in_14_,la_data_in_13_,la_data_in_12_,la_data_in_11_,la_data_in_10_,la_data_in_9_,la_data_in_8_,la_data_in_7_,la_data_in_6_,la_data_in_5_,la_data_in_4_,la_data_in_3_,la_data_in_2_,la_data_in_1_,la_data_in_0_
*.opin
*+ la_data_out_127_,la_data_out_126_,la_data_out_125_,la_data_out_124_,la_data_out_123_,la_data_out_122_,la_data_out_121_,la_data_out_120_,la_data_out_119_,la_data_out_118_,la_data_out_117_,la_data_out_116_,la_data_out_115_,la_data_out_114_,la_data_out_113_,la_data_out_112_,la_data_out_111_,la_data_out_110_,la_data_out_109_,la_data_out_108_,la_data_out_107_,la_data_out_106_,la_data_out_105_,la_data_out_104_,la_data_out_103_,la_data_out_102_,la_data_out_101_,la_data_out_100_,la_data_out_99_,la_data_out_98_,la_data_out_97_,la_data_out_96_,la_data_out_95_,la_data_out_94_,la_data_out_93_,la_data_out_92_,la_data_out_91_,la_data_out_90_,la_data_out_89_,la_data_out_88_,la_data_out_87_,la_data_out_86_,la_data_out_85_,la_data_out_84_,la_data_out_83_,la_data_out_82_,la_data_out_81_,la_data_out_80_,la_data_out_79_,la_data_out_78_,la_data_out_77_,la_data_out_76_,la_data_out_75_,la_data_out_74_,la_data_out_73_,la_data_out_72_,la_data_out_71_,la_data_out_70_,la_data_out_69_,la_data_out_68_,la_data_out_67_,la_data_out_66_,la_data_out_65_,la_data_out_64_,la_data_out_63_,la_data_out_62_,la_data_out_61_,la_data_out_60_,la_data_out_59_,la_data_out_58_,la_data_out_57_,la_data_out_56_,la_data_out_55_,la_data_out_54_,la_data_out_53_,la_data_out_52_,la_data_out_51_,la_data_out_50_,la_data_out_49_,la_data_out_48_,la_data_out_47_,la_data_out_46_,la_data_out_45_,la_data_out_44_,la_data_out_43_,la_data_out_42_,la_data_out_41_,la_data_out_40_,la_data_out_39_,la_data_out_38_,la_data_out_37_,la_data_out_36_,la_data_out_35_,la_data_out_34_,la_data_out_33_,la_data_out_32_,la_data_out_31_,la_data_out_30_,la_data_out_29_,la_data_out_28_,la_data_out_27_,la_data_out_26_,la_data_out_25_,la_data_out_24_,la_data_out_23_,la_data_out_22_,la_data_out_21_,la_data_out_20_,la_data_out_19_,la_data_out_18_,la_data_out_17_,la_data_out_16_,la_data_out_15_,la_data_out_14_,la_data_out_13_,la_data_out_12_,la_data_out_11_,la_data_out_10_,la_data_out_9_,la_data_out_8_,la_data_out_7_,la_data_out_6_,la_data_out_5_,la_data_out_4_,la_data_out_3_,la_data_out_2_,la_data_out_1_,la_data_out_0_
*.ipin
*+ io_in_26_,io_in_25_,io_in_24_,io_in_23_,io_in_22_,io_in_21_,io_in_20_,io_in_19_,io_in_18_,io_in_17_,io_in_16_,io_in_15_,io_in_14_,io_in_13_,io_in_12_,io_in_11_,io_in_10_,io_in_9_,io_in_8_,io_in_7_,io_in_6_,io_in_5_,io_in_4_,io_in_3_,io_in_2_,io_in_1_,io_in_0_
*.ipin
*+ io_in_3v3_26_,io_in_3v3_25_,io_in_3v3_24_,io_in_3v3_23_,io_in_3v3_22_,io_in_3v3_21_,io_in_3v3_20_,io_in_3v3_19_,io_in_3v3_18_,io_in_3v3_17_,io_in_3v3_16_,io_in_3v3_15_,io_in_3v3_14_,io_in_3v3_13_,io_in_3v3_12_,io_in_3v3_11_,io_in_3v3_10_,io_in_3v3_9_,io_in_3v3_8_,io_in_3v3_7_,io_in_3v3_6_,io_in_3v3_5_,io_in_3v3_4_,io_in_3v3_3_,io_in_3v3_2_,io_in_3v3_1_,io_in_3v3_0_
*.ipin user_clock2
*.opin
*+ io_out_26_,io_out_25_,io_out_24_,io_out_23_,io_out_22_,io_out_21_,io_out_20_,io_out_19_,io_out_18_,io_out_17_,io_out_16_,io_out_15_,io_out_14_,io_out_13_,io_out_12_,io_out_11_,io_out_10_,io_out_9_,io_out_8_,io_out_7_,io_out_6_,io_out_5_,io_out_4_,io_out_3_,io_out_2_,io_out_1_,io_out_0_
*.opin
*+ io_oeb_26_,io_oeb_25_,io_oeb_24_,io_oeb_23_,io_oeb_22_,io_oeb_21_,io_oeb_20_,io_oeb_19_,io_oeb_18_,io_oeb_17_,io_oeb_16_,io_oeb_15_,io_oeb_14_,io_oeb_13_,io_oeb_12_,io_oeb_11_,io_oeb_10_,io_oeb_9_,io_oeb_8_,io_oeb_7_,io_oeb_6_,io_oeb_5_,io_oeb_4_,io_oeb_3_,io_oeb_2_,io_oeb_1_,io_oeb_0_
*.iopin
*+ gpio_analog_17_,gpio_analog_16_,gpio_analog_15_,gpio_analog_14_,gpio_analog_13_,gpio_analog_12_,gpio_analog_11_,gpio_analog_10_,gpio_analog_9_,gpio_analog_8_,gpio_analog_7_,gpio_analog_6_,gpio_analog_5_,gpio_analog_4_,gpio_analog_3_,gpio_analog_2_,gpio_analog_1_,gpio_analog_0_
*.iopin
*+ gpio_noesd_17_,gpio_noesd_16_,gpio_noesd_15_,gpio_noesd_14_,gpio_noesd_13_,gpio_noesd_12_,gpio_noesd_11_,gpio_noesd_10_,gpio_noesd_9_,gpio_noesd_8_,gpio_noesd_7_,gpio_noesd_6_,gpio_noesd_5_,gpio_noesd_4_,gpio_noesd_3_,gpio_noesd_2_,gpio_noesd_1_,gpio_noesd_0_
*.iopin
*+ io_analog_10_,io_analog_9_,io_analog_8_,io_analog_7_,io_analog_6_,io_analog_5_,io_analog_4_,io_analog_3_,io_analog_2_,io_analog_1_,io_analog_0_
*.iopin io_clamp_high_2_,io_clamp_high_1_,io_clamp_high_0_
*.iopin io_clamp_low_2_,io_clamp_low_1_,io_clamp_low_0_
*.opin user_irq_2_,user_irq_1_,user_irq_0_
*.ipin
*+ la_oenb_127_,la_oenb_126_,la_oenb_125_,la_oenb_124_,la_oenb_123_,la_oenb_122_,la_oenb_121_,la_oenb_120_,la_oenb_119_,la_oenb_118_,la_oenb_117_,la_oenb_116_,la_oenb_115_,la_oenb_114_,la_oenb_113_,la_oenb_112_,la_oenb_111_,la_oenb_110_,la_oenb_109_,la_oenb_108_,la_oenb_107_,la_oenb_106_,la_oenb_105_,la_oenb_104_,la_oenb_103_,la_oenb_102_,la_oenb_101_,la_oenb_100_,la_oenb_99_,la_oenb_98_,la_oenb_97_,la_oenb_96_,la_oenb_95_,la_oenb_94_,la_oenb_93_,la_oenb_92_,la_oenb_91_,la_oenb_90_,la_oenb_89_,la_oenb_88_,la_oenb_87_,la_oenb_86_,la_oenb_85_,la_oenb_84_,la_oenb_83_,la_oenb_82_,la_oenb_81_,la_oenb_80_,la_oenb_79_,la_oenb_78_,la_oenb_77_,la_oenb_76_,la_oenb_75_,la_oenb_74_,la_oenb_73_,la_oenb_72_,la_oenb_71_,la_oenb_70_,la_oenb_69_,la_oenb_68_,la_oenb_67_,la_oenb_66_,la_oenb_65_,la_oenb_64_,la_oenb_63_,la_oenb_62_,la_oenb_61_,la_oenb_60_,la_oenb_59_,la_oenb_58_,la_oenb_57_,la_oenb_56_,la_oenb_55_,la_oenb_54_,la_oenb_53_,la_oenb_52_,la_oenb_51_,la_oenb_50_,la_oenb_49_,la_oenb_48_,la_oenb_47_,la_oenb_46_,la_oenb_45_,la_oenb_44_,la_oenb_43_,la_oenb_42_,la_oenb_41_,la_oenb_40_,la_oenb_39_,la_oenb_38_,la_oenb_37_,la_oenb_36_,la_oenb_35_,la_oenb_34_,la_oenb_33_,la_oenb_32_,la_oenb_31_,la_oenb_30_,la_oenb_29_,la_oenb_28_,la_oenb_27_,la_oenb_26_,la_oenb_25_,la_oenb_24_,la_oenb_23_,la_oenb_22_,la_oenb_21_,la_oenb_20_,la_oenb_19_,la_oenb_18_,la_oenb_17_,la_oenb_16_,la_oenb_15_,la_oenb_14_,la_oenb_13_,la_oenb_12_,la_oenb_11_,la_oenb_10_,la_oenb_9_,la_oenb_8_,la_oenb_7_,la_oenb_6_,la_oenb_5_,la_oenb_4_,la_oenb_3_,la_oenb_2_,la_oenb_1_,la_oenb_0_
xsar vdda1 vccd2 vssd2 la_data_out_29_ la_data_out_30_ la_data_out_31_ la_data_out_32_
+ la_data_out_33_ la_data_out_34_ la_data_out_35_ la_data_out_36_ io_analog_4_ vssa1 io_in_20_ io_analog_5_ io_in_19_
+ io_out_17_ io_in_18_ io_in_23_ sar
.ends

* expanding   symbol:  sar/sar/sar.sym # of pins=12
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/sar/sar.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/sar/sar.sch
.subckt sar avdd dvdd dvss result_7_ result_6_ result_5_ result_4_ result_3_ result_2_ result_1_
+ result_0_ vinn avss clk vinp en valid cal rstn
*.iopin avss
*.iopin avdd
*.iopin dvss
*.iopin dvdd
*.ipin vinp
*.ipin vinn
*.opin result_7_,result_6_,result_5_,result_4_,result_3_,result_2_,result_1_,result_0_
*.ipin clk
*.ipin en
*.opin valid
*.ipin cal
*.ipin rstn
xlat avdd comp net1 avss outn outp latch
**** begin user architecture code

.include /home/alex/Desktop/SAR_IPN/xschem/sar/control/cmos_cells_digital.sp
.include /home/alex/Desktop/SAR_IPN/xschem/sar/control/sar_logic.sp
*.include /home/alex/Desktop/SAR_IPN/xschem/sar/control/sar_logic_sky.sp

**** end user architecture code
xdn vn sample avdd avss vinn ctln_7_ ctln_6_ ctln_5_ ctln_4_ ctln_3_ ctln_2_ ctln_1_ ctln_0_ avss
+ dac
xdp vp sample avdd avss vinp ctlp_7_ ctlp_6_ ctlp_5_ ctlp_4_ ctlp_3_ ctlp_2_ ctlp_1_ ctlp_0_ avdd
+ dac
xcom avss avdd clkc outp vp outn vn trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ trimb_4_ trimb_3_
+ trimb_2_ trimb_1_ trimb_0_ comparator
**** begin user architecture code


Xuut dclk drstn den dcomp dcal dvalid dres0 dres1 dres2 dres3 dres4 dres5 dres6 dres7 dsamp dctlp0
+ dctlp1 dctlp2 dctlp3 dctlp4 dctlp5 dctlp6 dctlp7 dctln0 dctln1 dctln2 dctln3 dctln4 dctln5 dctln6 dctln7
+ dtrim0 dtrim1 dtrim2 dtrim3 dtrim4 dtrimb0 dtrimb1 dtrimb2 dtrimb3 dtrimb4 dclkc sar_logic

.model adc_buff adc_bridge(in_low = 0.2 in_high=0.8)
.model dac_buff dac_bridge(out_high = 1.2)

Aad [clk rstn en comp cal] [dclk drstn den dcomp dcal] adc_buff
Ada [dctlp0 dctlp1 dctlp2 dctlp3 dctlp4 dctlp5 dctlp6 dctlp7 dctln0 dctln1 dctln2 dctln3 dctln4
+ dctln5 dctln6 dctln7 dres0 dres1 dres2 dres3 dres4 dres5 dres6 dres7 dsamp dclkc] [ctlp_0_ ctlp_1_ ctlp_2_
+ ctlp_3_ ctlp_4_ ctlp_5_ ctlp_6_ ctlp_7_ ctln_0_ ctln_1_ ctln_2_ ctln_3_ ctln_4_ ctln_5_ ctln_6_ ctln_7_
+ res0 res1 res2 res3 res4 res5 res6 res7 sample clkc] dac_buff
Ada2 [dtrim4 dtrim3 dtrim2 dtrim1 dtrim0 dtrimb4 dtrimb3 dtrimb2 dtrimb1 dtrimb0] [trim_4_ trim_3_
+ trim_2_ trim_1_ trim_0_ trimb_4_ trimb_3_ trimb_2_ trimb_1_ trimb_0_ ] dac_buff



**** end user architecture code
.ends


* expanding   symbol:  sar/latch/latch.sym # of pins=6
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/latch/latch.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/latch/latch.sch
.subckt latch vdd Q Qn vss R S
*.ipin S
*.ipin R
*.iopin vss
*.iopin vdd
*.opin Q
*.opin Qn
x1 vdd Qn Q vss inv_lvt
x2 vdd Q Qn vss inv_lvt
x3 vdd R net2 vss inv_lvt
x4 vdd S net1 vss inv_lvt
XM4 Q net2 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 Qn net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sar/dac/dac.sym # of pins=7
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/dac/dac.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/dac/dac.sch
.subckt dac out sample vdd vss vin ctl_7_ ctl_6_ ctl_5_ ctl_4_ ctl_3_ ctl_2_ ctl_1_ ctl_0_ dum
*.ipin vin
*.ipin sample
*.opin out
*.ipin ctl_7_,ctl_6_,ctl_5_,ctl_4_,ctl_3_,ctl_2_,ctl_1_,ctl_0_
*.ipin dum
*.iopin vdd
*.iopin vss
xca out n6 n0 n5 n4 n2 ndum n3 n1 n7 carray
xi6 ctl_6_ vss vss vdd vdd n6 sky130_fd_sc_hd__inv_2
xi5 ctl_5_ vss vss vdd vdd n5 sky130_fd_sc_hd__inv_2
xi4 ctl_4_ vss vss vdd vdd n4 sky130_fd_sc_hd__inv_2
xi3 ctl_3_ vss vss vdd vdd n3 sky130_fd_sc_hd__inv_2
xi2 ctl_2_ vss vss vdd vdd n2 sky130_fd_sc_hd__inv_2
xi1 ctl_1_ vss vss vdd vdd n1 sky130_fd_sc_hd__inv_2
xi0 ctl_0_ vss vss vdd vdd n0 sky130_fd_sc_hd__inv_2
xidum dum vss vss vdd vdd ndum sky130_fd_sc_hd__inv_2
xi7 ctl_7_ vss vss vdd vdd n7 sky130_fd_sc_hd__inv_2
xswt out sample vdd vin vss sw_top
.ends


* expanding   symbol:  sar/comparator/comparator.sym # of pins=9
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/comparator.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/comparator.sch
.subckt comparator vss vdd clk outp vp outn vn trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ trimb_4_
+ trimb_3_ trimb_2_ trimb_1_ trimb_0_
*.ipin vn
*.ipin vp
*.ipin clk
*.iopin vdd
*.iopin vss
*.opin outp
*.opin outn
*.ipin trim_4_,trim_3_,trim_2_,trim_1_,trim_0_
*.ipin trimb_4_,trimb_3_,trimb_2_,trimb_1_,trimb_0_
x2 in trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ vss trim
x3 ip trimb_4_ trimb_3_ trimb_2_ trimb_1_ trimb_0_ vss trim
XM1 in clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 outn clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 outn outp vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMl4 outp outn vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 outp clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 ip clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMl2 outp outn ip vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMl1 outn outp in vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMinn in vn diff vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMinp ip vp diff vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMdiff diff clk vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  logic/inv_lvt.sym # of pins=4
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/logic/inv_lvt.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/logic/inv_lvt.sch
.subckt inv_lvt vdd in out vss
*.iopin vdd
*.iopin vss
*.ipin in
*.opin out
XM3 out in vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 out in vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sar/dac/carray.sym # of pins=10
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/dac/carray.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/dac/carray.sch
.subckt carray top n6 n0 n5 n4 n2 ndum n3 n1 n7
*.iopin top
*.iopin n7
*.iopin n6
*.iopin n5
*.iopin n4
*.iopin n2
*.iopin n0
*.iopin ndum
*.iopin n3
*.iopin n1
xcdum top ndum unitcap
xc0 top n0 unitcap
xc1_1_ top n1 unitcap
xc1_0_ top n1 unitcap
xc2_3_ top n2 unitcap
xc2_2_ top n2 unitcap
xc2_1_ top n2 unitcap
xc2_0_ top n2 unitcap
xc3_7_ top n3 unitcap
xc3_6_ top n3 unitcap
xc3_5_ top n3 unitcap
xc3_4_ top n3 unitcap
xc3_3_ top n3 unitcap
xc3_2_ top n3 unitcap
xc3_1_ top n3 unitcap
xc3_0_ top n3 unitcap
xc4_15_ top n4 unitcap
xc4_14_ top n4 unitcap
xc4_13_ top n4 unitcap
xc4_12_ top n4 unitcap
xc4_11_ top n4 unitcap
xc4_10_ top n4 unitcap
xc4_9_ top n4 unitcap
xc4_8_ top n4 unitcap
xc4_7_ top n4 unitcap
xc4_6_ top n4 unitcap
xc4_5_ top n4 unitcap
xc4_4_ top n4 unitcap
xc4_3_ top n4 unitcap
xc4_2_ top n4 unitcap
xc4_1_ top n4 unitcap
xc4_0_ top n4 unitcap
xc5_31_ top n5 unitcap
xc5_30_ top n5 unitcap
xc5_29_ top n5 unitcap
xc5_28_ top n5 unitcap
xc5_27_ top n5 unitcap
xc5_26_ top n5 unitcap
xc5_25_ top n5 unitcap
xc5_24_ top n5 unitcap
xc5_23_ top n5 unitcap
xc5_22_ top n5 unitcap
xc5_21_ top n5 unitcap
xc5_20_ top n5 unitcap
xc5_19_ top n5 unitcap
xc5_18_ top n5 unitcap
xc5_17_ top n5 unitcap
xc5_16_ top n5 unitcap
xc5_15_ top n5 unitcap
xc5_14_ top n5 unitcap
xc5_13_ top n5 unitcap
xc5_12_ top n5 unitcap
xc5_11_ top n5 unitcap
xc5_10_ top n5 unitcap
xc5_9_ top n5 unitcap
xc5_8_ top n5 unitcap
xc5_7_ top n5 unitcap
xc5_6_ top n5 unitcap
xc5_5_ top n5 unitcap
xc5_4_ top n5 unitcap
xc5_3_ top n5 unitcap
xc5_2_ top n5 unitcap
xc5_1_ top n5 unitcap
xc5_0_ top n5 unitcap
xc6_63_ top n6 unitcap
xc6_62_ top n6 unitcap
xc6_61_ top n6 unitcap
xc6_60_ top n6 unitcap
xc6_59_ top n6 unitcap
xc6_58_ top n6 unitcap
xc6_57_ top n6 unitcap
xc6_56_ top n6 unitcap
xc6_55_ top n6 unitcap
xc6_54_ top n6 unitcap
xc6_53_ top n6 unitcap
xc6_52_ top n6 unitcap
xc6_51_ top n6 unitcap
xc6_50_ top n6 unitcap
xc6_49_ top n6 unitcap
xc6_48_ top n6 unitcap
xc6_47_ top n6 unitcap
xc6_46_ top n6 unitcap
xc6_45_ top n6 unitcap
xc6_44_ top n6 unitcap
xc6_43_ top n6 unitcap
xc6_42_ top n6 unitcap
xc6_41_ top n6 unitcap
xc6_40_ top n6 unitcap
xc6_39_ top n6 unitcap
xc6_38_ top n6 unitcap
xc6_37_ top n6 unitcap
xc6_36_ top n6 unitcap
xc6_35_ top n6 unitcap
xc6_34_ top n6 unitcap
xc6_33_ top n6 unitcap
xc6_32_ top n6 unitcap
xc6_31_ top n6 unitcap
xc6_30_ top n6 unitcap
xc6_29_ top n6 unitcap
xc6_28_ top n6 unitcap
xc6_27_ top n6 unitcap
xc6_26_ top n6 unitcap
xc6_25_ top n6 unitcap
xc6_24_ top n6 unitcap
xc6_23_ top n6 unitcap
xc6_22_ top n6 unitcap
xc6_21_ top n6 unitcap
xc6_20_ top n6 unitcap
xc6_19_ top n6 unitcap
xc6_18_ top n6 unitcap
xc6_17_ top n6 unitcap
xc6_16_ top n6 unitcap
xc6_15_ top n6 unitcap
xc6_14_ top n6 unitcap
xc6_13_ top n6 unitcap
xc6_12_ top n6 unitcap
xc6_11_ top n6 unitcap
xc6_10_ top n6 unitcap
xc6_9_ top n6 unitcap
xc6_8_ top n6 unitcap
xc6_7_ top n6 unitcap
xc6_6_ top n6 unitcap
xc6_5_ top n6 unitcap
xc6_4_ top n6 unitcap
xc6_3_ top n6 unitcap
xc6_2_ top n6 unitcap
xc6_1_ top n6 unitcap
xc6_0_ top n6 unitcap
xc7_127_ top n7 unitcap
xc7_126_ top n7 unitcap
xc7_125_ top n7 unitcap
xc7_124_ top n7 unitcap
xc7_123_ top n7 unitcap
xc7_122_ top n7 unitcap
xc7_121_ top n7 unitcap
xc7_120_ top n7 unitcap
xc7_119_ top n7 unitcap
xc7_118_ top n7 unitcap
xc7_117_ top n7 unitcap
xc7_116_ top n7 unitcap
xc7_115_ top n7 unitcap
xc7_114_ top n7 unitcap
xc7_113_ top n7 unitcap
xc7_112_ top n7 unitcap
xc7_111_ top n7 unitcap
xc7_110_ top n7 unitcap
xc7_109_ top n7 unitcap
xc7_108_ top n7 unitcap
xc7_107_ top n7 unitcap
xc7_106_ top n7 unitcap
xc7_105_ top n7 unitcap
xc7_104_ top n7 unitcap
xc7_103_ top n7 unitcap
xc7_102_ top n7 unitcap
xc7_101_ top n7 unitcap
xc7_100_ top n7 unitcap
xc7_99_ top n7 unitcap
xc7_98_ top n7 unitcap
xc7_97_ top n7 unitcap
xc7_96_ top n7 unitcap
xc7_95_ top n7 unitcap
xc7_94_ top n7 unitcap
xc7_93_ top n7 unitcap
xc7_92_ top n7 unitcap
xc7_91_ top n7 unitcap
xc7_90_ top n7 unitcap
xc7_89_ top n7 unitcap
xc7_88_ top n7 unitcap
xc7_87_ top n7 unitcap
xc7_86_ top n7 unitcap
xc7_85_ top n7 unitcap
xc7_84_ top n7 unitcap
xc7_83_ top n7 unitcap
xc7_82_ top n7 unitcap
xc7_81_ top n7 unitcap
xc7_80_ top n7 unitcap
xc7_79_ top n7 unitcap
xc7_78_ top n7 unitcap
xc7_77_ top n7 unitcap
xc7_76_ top n7 unitcap
xc7_75_ top n7 unitcap
xc7_74_ top n7 unitcap
xc7_73_ top n7 unitcap
xc7_72_ top n7 unitcap
xc7_71_ top n7 unitcap
xc7_70_ top n7 unitcap
xc7_69_ top n7 unitcap
xc7_68_ top n7 unitcap
xc7_67_ top n7 unitcap
xc7_66_ top n7 unitcap
xc7_65_ top n7 unitcap
xc7_64_ top n7 unitcap
xc7_63_ top n7 unitcap
xc7_62_ top n7 unitcap
xc7_61_ top n7 unitcap
xc7_60_ top n7 unitcap
xc7_59_ top n7 unitcap
xc7_58_ top n7 unitcap
xc7_57_ top n7 unitcap
xc7_56_ top n7 unitcap
xc7_55_ top n7 unitcap
xc7_54_ top n7 unitcap
xc7_53_ top n7 unitcap
xc7_52_ top n7 unitcap
xc7_51_ top n7 unitcap
xc7_50_ top n7 unitcap
xc7_49_ top n7 unitcap
xc7_48_ top n7 unitcap
xc7_47_ top n7 unitcap
xc7_46_ top n7 unitcap
xc7_45_ top n7 unitcap
xc7_44_ top n7 unitcap
xc7_43_ top n7 unitcap
xc7_42_ top n7 unitcap
xc7_41_ top n7 unitcap
xc7_40_ top n7 unitcap
xc7_39_ top n7 unitcap
xc7_38_ top n7 unitcap
xc7_37_ top n7 unitcap
xc7_36_ top n7 unitcap
xc7_35_ top n7 unitcap
xc7_34_ top n7 unitcap
xc7_33_ top n7 unitcap
xc7_32_ top n7 unitcap
xc7_31_ top n7 unitcap
xc7_30_ top n7 unitcap
xc7_29_ top n7 unitcap
xc7_28_ top n7 unitcap
xc7_27_ top n7 unitcap
xc7_26_ top n7 unitcap
xc7_25_ top n7 unitcap
xc7_24_ top n7 unitcap
xc7_23_ top n7 unitcap
xc7_22_ top n7 unitcap
xc7_21_ top n7 unitcap
xc7_20_ top n7 unitcap
xc7_19_ top n7 unitcap
xc7_18_ top n7 unitcap
xc7_17_ top n7 unitcap
xc7_16_ top n7 unitcap
xc7_15_ top n7 unitcap
xc7_14_ top n7 unitcap
xc7_13_ top n7 unitcap
xc7_12_ top n7 unitcap
xc7_11_ top n7 unitcap
xc7_10_ top n7 unitcap
xc7_9_ top n7 unitcap
xc7_8_ top n7 unitcap
xc7_7_ top n7 unitcap
xc7_6_ top n7 unitcap
xc7_5_ top n7 unitcap
xc7_4_ top n7 unitcap
xc7_3_ top n7 unitcap
xc7_2_ top n7 unitcap
xc7_1_ top n7 unitcap
xc7_0_ top n7 unitcap
xdummy_83_ top dum_bot_83_ unitcap
xdummy_82_ top dum_bot_82_ unitcap
xdummy_81_ top dum_bot_81_ unitcap
xdummy_80_ top dum_bot_80_ unitcap
xdummy_79_ top dum_bot_79_ unitcap
xdummy_78_ top dum_bot_78_ unitcap
xdummy_77_ top dum_bot_77_ unitcap
xdummy_76_ top dum_bot_76_ unitcap
xdummy_75_ top dum_bot_75_ unitcap
xdummy_74_ top dum_bot_74_ unitcap
xdummy_73_ top dum_bot_73_ unitcap
xdummy_72_ top dum_bot_72_ unitcap
xdummy_71_ top dum_bot_71_ unitcap
xdummy_70_ top dum_bot_70_ unitcap
xdummy_69_ top dum_bot_69_ unitcap
xdummy_68_ top dum_bot_68_ unitcap
xdummy_67_ top dum_bot_67_ unitcap
xdummy_66_ top dum_bot_66_ unitcap
xdummy_65_ top dum_bot_65_ unitcap
xdummy_64_ top dum_bot_64_ unitcap
xdummy_63_ top dum_bot_63_ unitcap
xdummy_62_ top dum_bot_62_ unitcap
xdummy_61_ top dum_bot_61_ unitcap
xdummy_60_ top dum_bot_60_ unitcap
xdummy_59_ top dum_bot_59_ unitcap
xdummy_58_ top dum_bot_58_ unitcap
xdummy_57_ top dum_bot_57_ unitcap
xdummy_56_ top dum_bot_56_ unitcap
xdummy_55_ top dum_bot_55_ unitcap
xdummy_54_ top dum_bot_54_ unitcap
xdummy_53_ top dum_bot_53_ unitcap
xdummy_52_ top dum_bot_52_ unitcap
xdummy_51_ top dum_bot_51_ unitcap
xdummy_50_ top dum_bot_50_ unitcap
xdummy_49_ top dum_bot_49_ unitcap
xdummy_48_ top dum_bot_48_ unitcap
xdummy_47_ top dum_bot_47_ unitcap
xdummy_46_ top dum_bot_46_ unitcap
xdummy_45_ top dum_bot_45_ unitcap
xdummy_44_ top dum_bot_44_ unitcap
xdummy_43_ top dum_bot_43_ unitcap
xdummy_42_ top dum_bot_42_ unitcap
xdummy_41_ top dum_bot_41_ unitcap
xdummy_40_ top dum_bot_40_ unitcap
xdummy_39_ top dum_bot_39_ unitcap
xdummy_38_ top dum_bot_38_ unitcap
xdummy_37_ top dum_bot_37_ unitcap
xdummy_36_ top dum_bot_36_ unitcap
xdummy_35_ top dum_bot_35_ unitcap
xdummy_34_ top dum_bot_34_ unitcap
xdummy_33_ top dum_bot_33_ unitcap
xdummy_32_ top dum_bot_32_ unitcap
xdummy_31_ top dum_bot_31_ unitcap
xdummy_30_ top dum_bot_30_ unitcap
xdummy_29_ top dum_bot_29_ unitcap
xdummy_28_ top dum_bot_28_ unitcap
xdummy_27_ top dum_bot_27_ unitcap
xdummy_26_ top dum_bot_26_ unitcap
xdummy_25_ top dum_bot_25_ unitcap
xdummy_24_ top dum_bot_24_ unitcap
xdummy_23_ top dum_bot_23_ unitcap
xdummy_22_ top dum_bot_22_ unitcap
xdummy_21_ top dum_bot_21_ unitcap
xdummy_20_ top dum_bot_20_ unitcap
xdummy_19_ top dum_bot_19_ unitcap
xdummy_18_ top dum_bot_18_ unitcap
xdummy_17_ top dum_bot_17_ unitcap
xdummy_16_ top dum_bot_16_ unitcap
xdummy_15_ top dum_bot_15_ unitcap
xdummy_14_ top dum_bot_14_ unitcap
xdummy_13_ top dum_bot_13_ unitcap
xdummy_12_ top dum_bot_12_ unitcap
xdummy_11_ top dum_bot_11_ unitcap
xdummy_10_ top dum_bot_10_ unitcap
xdummy_9_ top dum_bot_9_ unitcap
xdummy_8_ top dum_bot_8_ unitcap
xdummy_7_ top dum_bot_7_ unitcap
xdummy_6_ top dum_bot_6_ unitcap
xdummy_5_ top dum_bot_5_ unitcap
xdummy_4_ top dum_bot_4_ unitcap
xdummy_3_ top dum_bot_3_ unitcap
xdummy_2_ top dum_bot_2_ unitcap
xdummy_1_ top dum_bot_1_ unitcap
xdummy_0_ top dum_bot_0_ unitcap
.ends


* expanding   symbol:  sar/sw/sw_top.sym # of pins=5
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/sw/sw_top.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/sw/sw_top.sch
.subckt sw_top out en vdd in vss
*.iopin out
*.ipin en
*.iopin vss
*.iopin vdd
*.iopin in
x2 vss vss vdd vdd sky130_fd_sc_hd__decap_8
x4 en vss vss vdd vdd en_buf sky130_fd_sc_hd__inv_4
x1 VGND VNB VPB VPWR sky130_fd_sc_hd__decap_3
XM1 in en out vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
XM2 in en_buf out vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=10 m=10
.ends


* expanding   symbol:  sar/comparator/trim.sym # of pins=3
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/trim.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/trim.sch
.subckt trim drain d_4_ d_3_ d_2_ d_1_ d_0_ vss
*.iopin vss
*.ipin d_4_,d_3_,d_2_,d_1_,d_0_
*.opin drain
x4_7_ drain n4 trimcap
x4_6_ drain n4 trimcap
x4_5_ drain n4 trimcap
x4_4_ drain n4 trimcap
x4_3_ drain n4 trimcap
x4_2_ drain n4 trimcap
x4_1_ drain n4 trimcap
x4_0_ drain n4 trimcap
x3_3_ drain n3 trimcap
x3_2_ drain n3 trimcap
x3_1_ drain n3 trimcap
x3_0_ drain n3 trimcap
x2_1_ drain n2 trimcap
x2_0_ drain n2 trimcap
x1 drain n1 trimcap
x0 drain n0 trimcap
XM4_7_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_6_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_5_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_4_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_3_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_2_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_1_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4_0_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3_3_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3_2_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3_1_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3_0_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2_1_ n2 d_2_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2_0_ n2 d_2_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 n1 d_1_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 n0 d_0_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sar/unitcap/unitcap.sym # of pins=2
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/unitcap/unitcap.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/unitcap/unitcap.sch
.subckt unitcap cp cn
*.iopin cp
*.iopin cn
XC2 cp cn sky130_fd_pr__cap_mim_m3_1 W=2 L=2 MF=1 m=1
.ends


* expanding   symbol:  sar/comparator/trimcap.sym # of pins=2
** sym_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/trimcap.sym
** sch_path: /home/alex/Desktop/SAR_IPN/xschem/sar/comparator/trimcap.sch
.subckt trimcap cp cn
*.iopin cp
*.iopin cn
C1 cp cn 2f m=1
.ends

.end
